module Benchmark_testing35000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2859,I2866,I22708,I22720,I22729,I22732,I22717,I22726,I22714,I22723,I22711,I69771,I69747,I69759,I69753,I69768,I69762,I69756,I69750,I69765,I143020,I143044,I143026,I143029,I143017,I143035,I143038,I143023,I143032,I143041,I160435,I160414,I160408,I160423,I160411,I160426,I160417,I160420,I160432,I160429,I210259,I210256,I210241,I210253,I210247,I210235,I210244,I210250,I210238,I255082,I255079,I255070,I255073,I255067,I255076,I255064,I255088,I255085,I292649,I292652,I292634,I292643,I292655,I292646,I292637,I292640,I292658,I350758,I350761,I350752,I350743,I350746,I350755,I350740,I350749,I392836,I392839,I392815,I392827,I392842,I392830,I392824,I392818,I392821,I392833,I398004,I398007,I397983,I397995,I398010,I397998,I397992,I397986,I397989,I398001,I455101,I455089,I455110,I455086,I455107,I455098,I455104,I455095,I455092,I473019,I473007,I473028,I473004,I473025,I473016,I473022,I473013,I473010,I483423,I483411,I483432,I483408,I483429,I483420,I483426,I483417,I483414,I484001,I483989,I484010,I483986,I484007,I483998,I484004,I483995,I483992,I496717,I496705,I496726,I496702,I496723,I496714,I496720,I496711,I496708,I521240,I521219,I521225,I521234,I521237,I521216,I521231,I521228,I521222,I558823,I558838,I558820,I558832,I558847,I558844,I558841,I558835,I558829,I558826);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2859,I2866;
output I22708,I22720,I22729,I22732,I22717,I22726,I22714,I22723,I22711,I69771,I69747,I69759,I69753,I69768,I69762,I69756,I69750,I69765,I143020,I143044,I143026,I143029,I143017,I143035,I143038,I143023,I143032,I143041,I160435,I160414,I160408,I160423,I160411,I160426,I160417,I160420,I160432,I160429,I210259,I210256,I210241,I210253,I210247,I210235,I210244,I210250,I210238,I255082,I255079,I255070,I255073,I255067,I255076,I255064,I255088,I255085,I292649,I292652,I292634,I292643,I292655,I292646,I292637,I292640,I292658,I350758,I350761,I350752,I350743,I350746,I350755,I350740,I350749,I392836,I392839,I392815,I392827,I392842,I392830,I392824,I392818,I392821,I392833,I398004,I398007,I397983,I397995,I398010,I397998,I397992,I397986,I397989,I398001,I455101,I455089,I455110,I455086,I455107,I455098,I455104,I455095,I455092,I473019,I473007,I473028,I473004,I473025,I473016,I473022,I473013,I473010,I483423,I483411,I483432,I483408,I483429,I483420,I483426,I483417,I483414,I484001,I483989,I484010,I483986,I484007,I483998,I484004,I483995,I483992,I496717,I496705,I496726,I496702,I496723,I496714,I496720,I496711,I496708,I521240,I521219,I521225,I521234,I521237,I521216,I521231,I521228,I521222,I558823,I558838,I558820,I558832,I558847,I558844,I558841,I558835,I558829,I558826;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2859,I2866,I2898,I92955,I2924,I2932,I2949,I2890,I92961,I2989,I2997,I3014,I92970,I3031,I92964,I3048,I3065,I2869,I3096,I3113,I3130,I92967,I92973,I2872,I3161,I3178,I92976,I3195,I92952,I3212,I3229,I3246,I2881,I3277,I92958,I3294,I3311,I2887,I3342,I2884,I3373,I3399,I3407,I3424,I2878,I2875,I3493,I411570,I3519,I3527,I411561,I3544,I3485,I411564,I3584,I3592,I3609,I411576,I3626,I411555,I3643,I3660,I3464,I3691,I3708,I3725,I411567,I411573,I3467,I3756,I3773,I411558,I3790,I411549,I3807,I3824,I3841,I3476,I3872,I3889,I3906,I3482,I3937,I3479,I3968,I411552,I3994,I4002,I4019,I3473,I3470,I4088,I536225,I4114,I4122,I536216,I4139,I4080,I536219,I4179,I4187,I4204,I536231,I4221,I536222,I4238,I4255,I4059,I4286,I4303,I4320,I536210,I4062,I4351,I4368,I536234,I4385,I536213,I4402,I4419,I4436,I4071,I4467,I536228,I4484,I4501,I4077,I4532,I4074,I4563,I536237,I4589,I4597,I4614,I4068,I4065,I4683,I176749,I4709,I4717,I176731,I4734,I4675,I176743,I4774,I4782,I4799,I176728,I4816,I176737,I4833,I4850,I4654,I4881,I4898,I4915,I176734,I176755,I4657,I4946,I4963,I176746,I4980,I176752,I4997,I5014,I5031,I4666,I5062,I5079,I5096,I4672,I5127,I4669,I5158,I176740,I5184,I5192,I5209,I4663,I4660,I5278,I184909,I5304,I5312,I184891,I5329,I5270,I184903,I5369,I5377,I5394,I184888,I5411,I184897,I5428,I5445,I5249,I5476,I5493,I5510,I184894,I184915,I5252,I5541,I5558,I184906,I5575,I184912,I5592,I5609,I5626,I5261,I5657,I5674,I5691,I5267,I5722,I5264,I5753,I184900,I5779,I5787,I5804,I5258,I5255,I5876,I529323,I5902,I5919,I5927,I5944,I529326,I529320,I5961,I529329,I5987,I5868,I5859,I529317,I6032,I6040,I529332,I6057,I5856,I529308,I6097,I6105,I5862,I5850,I6150,I529311,I6167,I6193,I6201,I5844,I6232,I6249,I529314,I6266,I6283,I6300,I5865,I6331,I5853,I5847,I6403,I288016,I6429,I6446,I6454,I6471,I288031,I288034,I6488,I288013,I6514,I6395,I6386,I288019,I6559,I6567,I288025,I6584,I6383,I6624,I6632,I6389,I6377,I6677,I288028,I288010,I6694,I288022,I6720,I6728,I6371,I6759,I6776,I6793,I6810,I6827,I6392,I6858,I6380,I6374,I6930,I195768,I6956,I6973,I6981,I6998,I195771,I7015,I195792,I7041,I6922,I6913,I195780,I7086,I7094,I195783,I7111,I6910,I195789,I7151,I7159,I6916,I6904,I7204,I195786,I195774,I7221,I195777,I7247,I7255,I6898,I7286,I7303,I195795,I7320,I7337,I7354,I6919,I7385,I6907,I6901,I7457,I496148,I7483,I7500,I7508,I7525,I496136,I496127,I7542,I496124,I7568,I7449,I7440,I496130,I7613,I7621,I496142,I7638,I7437,I496139,I7678,I7686,I7443,I7431,I7731,I496133,I7748,I496145,I7774,I7782,I7425,I7813,I7830,I7847,I7864,I7881,I7446,I7912,I7434,I7428,I7984,I207864,I8010,I8027,I8035,I8052,I207870,I207858,I8069,I207855,I8095,I7976,I7967,I207867,I8140,I8148,I207861,I8165,I7964,I207879,I8205,I8213,I7970,I7958,I8258,I207873,I207876,I8275,I8301,I8309,I7952,I8340,I8357,I8374,I8391,I8408,I7973,I8439,I7961,I7955,I8511,I281658,I8537,I8554,I8562,I8579,I281673,I281676,I8596,I281655,I8622,I8503,I8494,I281661,I8667,I8675,I281667,I8692,I8491,I8732,I8740,I8497,I8485,I8785,I281670,I281652,I8802,I281664,I8828,I8836,I8479,I8867,I8884,I8901,I8918,I8935,I8500,I8966,I8488,I8482,I9038,I101883,I9064,I9081,I9089,I9106,I101901,I101886,I9123,I101889,I9149,I9030,I9021,I101877,I9194,I9202,I101880,I9219,I9018,I101892,I9259,I9267,I9024,I9012,I9312,I101898,I101895,I9329,I9355,I9363,I9006,I9394,I9411,I9428,I9445,I9462,I9027,I9493,I9015,I9009,I9565,I253923,I9591,I9608,I9616,I9633,I253908,I253926,I9650,I253920,I9676,I9557,I9548,I253917,I9721,I9729,I9746,I9545,I253911,I9786,I9794,I9551,I9539,I9839,I253932,I253914,I9856,I253929,I9882,I9890,I9533,I9921,I9938,I9955,I9972,I9989,I9554,I10020,I9542,I9536,I10092,I331777,I10118,I10135,I10143,I10160,I331768,I331789,I10177,I331771,I10203,I10084,I10075,I10248,I10256,I331786,I10273,I10072,I331780,I10313,I10321,I10078,I10066,I10366,I331774,I331783,I10383,I10409,I10417,I10060,I10448,I10465,I10482,I10499,I10516,I10081,I10547,I10069,I10063,I10619,I535615,I10645,I10662,I10670,I10687,I535618,I535624,I10704,I535633,I10730,I10611,I10602,I535636,I10775,I10783,I535627,I10800,I10599,I10840,I10848,I10605,I10593,I10893,I535642,I535621,I10910,I535630,I10936,I10944,I10587,I10975,I10992,I535639,I11009,I11026,I11043,I10608,I11074,I10596,I10590,I11146,I456844,I11172,I11189,I11197,I11214,I456832,I456823,I11231,I456820,I11257,I11138,I11129,I456826,I11302,I11310,I456838,I11327,I11126,I456835,I11367,I11375,I11132,I11120,I11420,I456829,I11437,I456841,I11463,I11471,I11114,I11502,I11519,I11536,I11553,I11570,I11135,I11601,I11123,I11117,I11673,I341790,I11699,I11716,I11724,I11741,I341781,I341802,I11758,I341784,I11784,I11665,I11656,I11829,I11837,I341799,I11854,I11653,I341793,I11894,I11902,I11659,I11647,I11947,I341787,I341796,I11964,I11990,I11998,I11641,I12029,I12046,I12063,I12080,I12097,I11662,I12128,I11650,I11644,I12200,I206674,I12226,I12243,I12251,I12268,I206680,I206668,I12285,I206665,I12311,I12192,I12183,I206677,I12356,I12364,I206671,I12381,I12180,I206689,I12421,I12429,I12186,I12174,I12474,I206683,I206686,I12491,I12517,I12525,I12168,I12556,I12573,I12590,I12607,I12624,I12189,I12655,I12177,I12171,I12727,I163672,I12753,I12770,I12778,I12795,I163675,I12812,I163696,I12838,I12719,I12710,I163684,I12883,I12891,I163687,I12908,I12707,I163693,I12948,I12956,I12713,I12701,I13001,I163690,I163678,I13018,I163681,I13044,I13052,I12695,I13083,I13100,I163699,I13117,I13134,I13151,I12716,I13182,I12704,I12698,I13254,I338628,I13280,I13297,I13305,I13322,I338619,I338640,I13339,I338622,I13365,I13246,I13237,I13410,I13418,I338637,I13435,I13234,I338631,I13475,I13483,I13240,I13228,I13528,I338625,I338634,I13545,I13571,I13579,I13222,I13610,I13627,I13644,I13661,I13678,I13243,I13709,I13231,I13225,I13781,I272988,I13807,I13824,I13832,I13849,I273003,I273006,I13866,I272985,I13892,I13773,I13764,I272991,I13937,I13945,I272997,I13962,I13761,I14002,I14010,I13767,I13755,I14055,I273000,I272982,I14072,I272994,I14098,I14106,I13749,I14137,I14154,I14171,I14188,I14205,I13770,I14236,I13758,I13752,I14308,I188152,I14334,I14351,I14359,I14376,I188155,I14393,I188176,I14419,I14300,I14291,I188164,I14464,I14472,I188167,I14489,I14288,I188173,I14529,I14537,I14294,I14282,I14582,I188170,I188158,I14599,I188161,I14625,I14633,I14276,I14664,I14681,I188179,I14698,I14715,I14732,I14297,I14763,I14285,I14279,I14835,I404467,I14861,I14878,I14886,I14903,I404443,I404470,I14920,I404455,I14946,I14827,I14818,I404461,I14991,I14999,I404446,I15016,I14815,I404464,I15056,I15064,I14821,I14809,I15109,I404449,I404452,I15126,I15152,I15160,I14803,I15191,I15208,I404458,I15225,I15242,I15259,I14824,I15290,I14812,I14806,I15362,I256235,I15388,I15405,I15413,I15430,I256220,I256238,I15447,I256232,I15473,I15354,I15345,I256229,I15518,I15526,I15543,I15342,I256223,I15583,I15591,I15348,I15336,I15636,I256244,I256226,I15653,I256241,I15679,I15687,I15330,I15718,I15735,I15752,I15769,I15786,I15351,I15817,I15339,I15333,I15889,I353384,I15915,I15932,I15940,I15957,I353375,I353396,I15974,I353378,I16000,I15881,I15872,I16045,I16053,I353393,I16070,I15869,I353387,I16110,I16118,I15875,I15863,I16163,I353381,I353390,I16180,I16206,I16214,I15857,I16245,I16262,I16279,I16296,I16313,I15878,I16344,I15866,I15860,I16416,I16442,I16459,I16467,I16484,I16501,I16527,I16408,I16399,I16572,I16580,I16597,I16396,I16637,I16645,I16402,I16390,I16690,I16707,I16733,I16741,I16384,I16772,I16789,I16806,I16823,I16840,I16405,I16871,I16393,I16387,I16943,I524121,I16969,I16986,I16994,I17011,I524124,I524118,I17028,I524127,I17054,I16935,I16926,I524115,I17099,I17107,I524130,I17124,I16923,I524106,I17164,I17172,I16929,I16917,I17217,I524109,I17234,I17260,I17268,I16911,I17299,I17316,I524112,I17333,I17350,I17367,I16932,I17398,I16920,I16914,I17470,I96528,I17496,I17513,I17521,I17538,I96546,I96531,I17555,I96534,I17581,I17462,I17453,I96522,I17626,I17634,I96525,I17651,I17450,I96537,I17691,I17699,I17456,I17444,I17744,I96543,I96540,I17761,I17787,I17795,I17438,I17826,I17843,I17860,I17877,I17894,I17459,I17925,I17447,I17441,I17997,I227913,I18023,I18040,I18048,I18065,I227898,I227916,I18082,I227910,I18108,I17989,I17980,I227907,I18153,I18161,I18178,I17977,I227901,I18218,I18226,I17983,I17971,I18271,I227922,I227904,I18288,I227919,I18314,I18322,I17965,I18353,I18370,I18387,I18404,I18421,I17986,I18452,I17974,I17968,I18524,I222127,I18550,I18558,I18575,I222139,I222124,I18592,I222118,I18618,I222133,I18635,I18643,I222121,I18660,I18492,I18691,I18708,I18504,I222130,I18748,I18513,I18770,I222136,I222142,I18787,I18813,I18830,I18516,I18852,I18501,I18883,I18900,I18917,I18934,I18510,I18965,I18498,I18507,I18495,I19051,I19077,I19085,I19102,I19119,I19145,I19162,I19170,I19187,I19019,I19218,I19235,I19031,I19275,I19040,I19297,I19314,I19340,I19357,I19043,I19379,I19028,I19410,I19427,I19444,I19461,I19037,I19492,I19025,I19034,I19022,I19578,I328615,I19604,I19612,I19629,I328612,I328627,I19646,I328609,I19672,I328606,I19689,I19697,I19714,I19546,I19745,I19762,I19558,I19802,I19567,I19824,I328621,I19841,I328624,I19867,I19884,I19570,I19906,I19555,I19937,I328618,I19954,I19971,I19988,I19564,I20019,I19552,I19561,I19549,I20105,I564782,I20131,I20139,I20156,I564776,I564797,I20173,I564773,I20199,I564794,I20216,I20224,I564791,I20241,I20073,I20272,I20289,I20085,I564779,I20329,I20094,I20351,I564788,I564785,I20368,I564770,I20394,I20411,I20097,I20433,I20082,I20464,I20481,I20498,I20515,I20091,I20546,I20079,I20088,I20076,I20632,I142517,I20658,I20666,I20683,I142499,I142514,I20700,I142490,I20726,I142493,I20743,I20751,I142508,I20768,I20600,I20799,I20816,I20612,I142511,I20856,I20621,I20878,I142502,I20895,I142496,I20921,I20938,I20624,I20960,I20609,I20991,I142505,I21008,I21025,I21042,I20618,I21073,I20606,I20615,I20603,I21159,I367630,I21185,I21193,I21210,I367648,I367642,I21227,I367621,I21253,I367639,I21270,I21278,I367624,I21295,I21127,I21326,I21343,I21139,I367636,I21383,I21148,I21405,I367645,I367633,I21422,I367627,I21448,I21465,I21151,I21487,I21136,I21518,I21535,I21552,I21569,I21145,I21600,I21133,I21142,I21130,I21686,I471854,I21712,I21720,I21737,I471869,I471848,I21754,I471851,I21780,I471872,I21797,I21805,I21822,I21654,I21853,I21870,I21666,I21910,I21675,I21932,I471860,I471857,I21949,I471863,I21975,I21992,I21678,I22014,I21663,I22045,I471866,I22062,I22079,I22096,I21672,I22127,I21660,I21669,I21657,I22213,I320183,I22239,I22247,I22264,I320180,I320195,I22281,I320177,I22307,I320174,I22324,I22332,I22349,I22181,I22380,I22397,I22193,I22437,I22202,I22459,I320189,I22476,I320192,I22502,I22519,I22205,I22541,I22190,I22572,I320186,I22589,I22606,I22623,I22199,I22654,I22187,I22196,I22184,I22740,I420392,I22766,I22774,I22791,I420389,I420395,I22808,I22834,I22851,I22859,I22876,I22907,I22924,I420398,I22964,I22986,I420401,I420410,I23003,I420404,I23029,I23046,I23068,I23099,I420407,I23116,I23133,I23150,I23181,I23267,I139882,I23293,I23301,I23318,I139864,I139879,I23335,I139855,I23361,I139858,I23378,I23386,I139873,I23403,I23235,I23434,I23451,I23247,I139876,I23491,I23256,I23513,I139867,I23530,I139861,I23556,I23573,I23259,I23595,I23244,I23626,I139870,I23643,I23660,I23677,I23253,I23708,I23241,I23250,I23238,I23794,I245825,I23820,I23828,I23845,I245837,I245822,I23862,I245816,I23888,I245831,I23905,I23913,I245819,I23930,I23762,I23961,I23978,I23774,I245828,I24018,I23783,I24040,I245834,I245840,I24057,I24083,I24100,I23786,I24122,I23771,I24153,I24170,I24187,I24204,I23780,I24235,I23768,I23777,I23765,I24321,I476478,I24347,I24355,I24372,I476493,I476472,I24389,I476475,I24415,I476496,I24432,I24440,I24457,I24289,I24488,I24505,I24301,I24545,I24310,I24567,I476484,I476481,I24584,I476487,I24610,I24627,I24313,I24649,I24298,I24680,I476490,I24697,I24714,I24731,I24307,I24762,I24295,I24304,I24292,I24848,I460294,I24874,I24882,I24899,I460309,I460288,I24916,I460291,I24942,I460312,I24959,I24967,I24984,I24816,I25015,I25032,I24828,I25072,I24837,I25094,I460300,I460297,I25111,I460303,I25137,I25154,I24840,I25176,I24825,I25207,I460306,I25224,I25241,I25258,I24834,I25289,I24822,I24831,I24819,I25375,I333358,I25401,I25409,I25426,I333355,I333370,I25443,I333352,I25469,I333349,I25486,I25494,I25511,I25343,I25542,I25559,I25355,I25599,I25364,I25621,I333364,I25638,I333367,I25664,I25681,I25367,I25703,I25352,I25734,I333361,I25751,I25768,I25785,I25361,I25816,I25349,I25358,I25346,I25902,I374736,I25928,I25936,I25953,I374754,I374748,I25970,I374727,I25996,I374745,I26013,I26021,I374730,I26038,I25870,I26069,I26086,I25882,I374742,I26126,I25891,I26148,I374751,I374739,I26165,I374733,I26191,I26208,I25894,I26230,I25879,I26261,I26278,I26295,I26312,I25888,I26343,I25876,I25885,I25873,I26429,I391532,I26455,I26463,I26480,I391550,I391544,I26497,I391523,I26523,I391541,I26540,I26548,I391526,I26565,I26397,I26596,I26613,I26409,I391538,I26653,I26418,I26675,I391547,I391535,I26692,I391529,I26718,I26735,I26421,I26757,I26406,I26788,I26805,I26822,I26839,I26415,I26870,I26403,I26412,I26400,I26956,I505208,I26982,I26990,I27007,I505202,I505223,I27024,I505214,I27050,I505205,I27067,I27075,I505217,I27092,I26924,I27123,I27140,I26936,I27180,I26945,I27202,I505226,I505211,I27219,I27245,I27262,I26948,I27284,I26933,I27315,I505220,I27332,I27349,I27366,I26942,I27397,I26930,I26939,I26927,I27483,I120910,I27509,I27517,I27534,I120892,I120907,I27551,I120883,I27577,I120886,I27594,I27602,I120901,I27619,I27451,I27650,I27667,I27463,I120904,I27707,I27472,I27729,I120895,I27746,I120889,I27772,I27789,I27475,I27811,I27460,I27842,I120898,I27859,I27876,I27893,I27469,I27924,I27457,I27466,I27454,I28010,I403160,I28036,I28044,I28061,I403178,I403172,I28078,I403151,I28104,I403169,I28121,I28129,I403154,I28146,I27978,I28177,I28194,I27990,I403166,I28234,I27999,I28256,I403175,I403163,I28273,I403157,I28299,I28316,I28002,I28338,I27987,I28369,I28386,I28403,I28420,I27996,I28451,I27984,I27993,I27981,I28537,I255651,I28563,I28571,I28588,I255663,I255648,I28605,I255642,I28631,I255657,I28648,I28656,I255645,I28673,I28505,I28704,I28721,I28517,I255654,I28761,I28526,I28783,I255660,I255666,I28800,I28826,I28843,I28529,I28865,I28514,I28896,I28913,I28930,I28947,I28523,I28978,I28511,I28520,I28508,I29064,I171306,I29090,I29098,I29115,I171300,I171291,I29132,I171312,I29158,I171294,I29175,I29183,I171288,I29200,I29032,I29231,I29248,I29044,I29288,I29053,I29310,I171315,I171297,I29327,I171303,I29353,I29370,I29056,I29392,I29041,I29423,I171309,I29440,I29457,I29474,I29050,I29505,I29038,I29047,I29035,I29591,I59644,I29617,I29625,I29642,I59638,I59632,I29659,I59653,I29685,I59650,I29702,I29710,I59647,I29727,I29559,I29758,I29775,I29571,I29815,I29580,I29837,I59635,I29854,I59656,I29880,I29897,I29583,I29919,I29568,I29950,I59641,I29967,I29984,I30001,I29577,I30032,I29565,I29574,I29562,I30118,I94154,I30144,I30152,I30169,I94148,I94142,I30186,I94163,I30212,I94160,I30229,I30237,I94157,I30254,I30086,I30285,I30302,I30098,I30342,I30107,I30364,I94145,I30381,I94166,I30407,I30424,I30110,I30446,I30095,I30477,I94151,I30494,I30511,I30528,I30104,I30559,I30092,I30101,I30089,I30645,I67974,I30671,I30679,I30696,I67968,I67962,I30713,I67983,I30739,I67980,I30756,I30764,I67977,I30781,I30613,I30812,I30829,I30625,I30869,I30634,I30891,I67965,I30908,I67986,I30934,I30951,I30637,I30973,I30622,I31004,I67971,I31021,I31038,I31055,I30631,I31086,I30619,I30628,I30616,I31172,I145679,I31198,I31206,I31223,I145661,I145676,I31240,I145652,I31266,I145655,I31283,I31291,I145670,I31308,I31140,I31339,I31356,I31152,I145673,I31396,I31161,I31418,I145664,I31435,I145658,I31461,I31478,I31164,I31500,I31149,I31531,I145667,I31548,I31565,I31582,I31158,I31613,I31146,I31155,I31143,I31699,I335466,I31725,I31733,I31750,I335463,I335478,I31767,I335460,I31793,I335457,I31810,I31818,I31835,I31667,I31866,I31883,I31679,I31923,I31688,I31945,I335472,I31962,I335475,I31988,I32005,I31691,I32027,I31676,I32058,I335469,I32075,I32092,I32109,I31685,I32140,I31673,I31682,I31670,I32226,I166410,I32252,I32260,I32277,I166404,I166395,I32294,I166416,I32320,I166398,I32337,I32345,I166392,I32362,I32194,I32393,I32410,I32206,I32450,I32215,I32472,I166419,I166401,I32489,I166407,I32515,I32532,I32218,I32554,I32203,I32585,I166413,I32602,I32619,I32636,I32212,I32667,I32200,I32209,I32197,I32753,I563592,I32779,I32787,I32804,I563586,I563607,I32821,I563583,I32847,I563604,I32864,I32872,I563601,I32889,I32721,I32920,I32937,I32733,I563589,I32977,I32742,I32999,I563598,I563595,I33016,I563580,I33042,I33059,I32745,I33081,I32730,I33112,I33129,I33146,I33163,I32739,I33194,I32727,I32736,I32724,I33280,I445266,I33306,I33314,I33331,I445281,I445260,I33348,I445263,I33374,I445284,I33391,I33399,I33416,I33248,I33447,I33464,I33260,I33504,I33269,I33526,I445272,I445269,I33543,I445275,I33569,I33586,I33272,I33608,I33257,I33639,I445278,I33656,I33673,I33690,I33266,I33721,I33254,I33263,I33251,I33807,I564187,I33833,I33841,I33858,I564181,I564202,I33875,I564178,I33901,I564199,I33918,I33926,I564196,I33943,I33775,I33974,I33991,I33787,I564184,I34031,I33796,I34053,I564193,I564190,I34070,I564175,I34096,I34113,I33799,I34135,I33784,I34166,I34183,I34200,I34217,I33793,I34248,I33781,I33790,I33778,I34334,I306518,I34360,I34368,I34385,I306509,I306527,I34402,I306506,I34428,I34445,I34453,I306512,I34470,I34302,I34501,I34518,I34314,I34558,I34323,I34580,I306524,I306515,I34597,I306530,I34623,I34640,I34326,I34662,I34311,I34693,I306521,I34710,I34727,I34744,I34320,I34775,I34308,I34317,I34305,I34861,I535032,I34887,I34895,I34912,I535026,I535047,I34929,I535023,I34955,I535044,I34972,I34980,I535041,I34997,I34829,I35028,I35045,I34841,I535029,I35085,I34850,I35107,I535038,I535035,I35124,I535020,I35150,I35167,I34853,I35189,I34838,I35220,I35237,I35254,I35271,I34847,I35302,I34835,I34844,I34832,I35388,I451046,I35414,I35422,I35439,I451061,I451040,I35456,I451043,I35482,I451064,I35499,I35507,I35524,I35356,I35555,I35572,I35368,I35612,I35377,I35634,I451052,I451049,I35651,I451055,I35677,I35694,I35380,I35716,I35365,I35747,I451058,I35764,I35781,I35798,I35374,I35829,I35362,I35371,I35359,I35915,I109029,I35941,I35949,I35966,I109023,I109017,I35983,I109038,I36009,I109035,I36026,I36034,I109032,I36051,I35883,I36082,I36099,I35895,I36139,I35904,I36161,I109020,I36178,I109041,I36204,I36221,I35907,I36243,I35892,I36274,I109026,I36291,I36308,I36325,I35901,I36356,I35889,I35898,I35886,I36442,I155165,I36468,I36476,I36493,I155147,I155162,I36510,I155138,I36536,I155141,I36553,I36561,I155156,I36578,I36410,I36609,I36626,I36422,I155159,I36666,I36431,I36688,I155150,I36705,I155144,I36731,I36748,I36434,I36770,I36419,I36801,I155153,I36818,I36835,I36852,I36428,I36883,I36416,I36425,I36413,I36969,I198506,I36995,I37003,I37020,I198500,I198491,I37037,I198512,I37063,I198494,I37080,I37088,I198488,I37105,I36937,I37136,I37153,I36949,I37193,I36958,I37215,I198515,I198497,I37232,I198503,I37258,I37275,I36961,I37297,I36946,I37328,I198509,I37345,I37362,I37379,I36955,I37410,I36943,I36952,I36940,I37496,I203693,I37522,I37530,I37547,I203714,I203708,I37564,I203690,I37590,I37607,I37615,I203702,I37632,I37464,I37663,I37680,I37476,I203699,I37720,I37485,I37742,I203705,I203696,I37759,I37785,I37802,I37488,I37824,I37473,I37855,I203711,I37872,I37889,I37906,I37482,I37937,I37470,I37479,I37467,I38023,I319129,I38049,I38057,I38074,I319126,I319141,I38091,I319123,I38117,I319120,I38134,I38142,I38159,I37991,I38190,I38207,I38003,I38247,I38012,I38269,I319135,I38286,I319138,I38312,I38329,I38015,I38351,I38000,I38382,I319132,I38399,I38416,I38433,I38009,I38464,I37997,I38006,I37994,I38550,I531620,I38576,I38584,I38601,I531626,I531644,I38618,I531641,I38644,I531638,I38661,I38669,I531632,I38686,I38518,I38717,I38734,I38530,I38774,I38539,I38796,I531635,I531623,I38813,I531647,I38839,I38856,I38542,I38878,I38527,I38909,I531629,I38926,I38943,I38960,I38536,I38991,I38524,I38533,I38521,I39077,I98319,I39103,I39111,I39128,I98313,I98307,I39145,I98328,I39171,I98325,I39188,I39196,I98322,I39213,I39045,I39244,I39261,I39057,I39301,I39066,I39323,I98310,I39340,I98331,I39366,I39383,I39069,I39405,I39054,I39436,I98316,I39453,I39470,I39487,I39063,I39518,I39051,I39060,I39048,I39604,I69164,I39630,I39638,I39655,I69158,I69152,I39672,I69173,I39698,I69170,I39715,I39723,I69167,I39740,I39572,I39771,I39788,I39584,I39828,I39593,I39850,I69155,I39867,I69176,I39893,I39910,I39596,I39932,I39581,I39963,I69161,I39980,I39997,I40014,I39590,I40045,I39578,I39587,I39575,I40131,I530485,I40157,I40165,I40182,I530488,I530482,I40199,I530479,I40225,I530464,I40242,I40250,I530473,I40267,I40099,I40298,I40315,I40111,I40355,I40120,I40377,I530467,I530470,I40394,I530476,I40420,I40437,I40123,I40459,I40108,I40490,I40507,I40524,I40541,I40117,I40572,I40105,I40114,I40102,I40658,I517769,I40684,I40692,I40709,I517772,I517766,I40726,I517763,I40752,I517748,I40769,I40777,I517757,I40794,I40626,I40825,I40842,I40638,I40882,I40647,I40904,I517751,I517754,I40921,I517760,I40947,I40964,I40650,I40986,I40635,I41017,I41034,I41051,I41068,I40644,I41099,I40632,I40641,I40629,I41185,I293224,I41211,I41219,I41236,I293215,I293233,I41253,I293212,I41279,I41296,I41304,I293218,I41321,I41153,I41352,I41369,I41165,I41409,I41174,I41431,I293230,I293221,I41448,I293236,I41474,I41491,I41177,I41513,I41162,I41544,I293227,I41561,I41578,I41595,I41171,I41626,I41159,I41168,I41156,I41712,I387656,I41738,I41746,I41763,I387674,I387668,I41780,I387647,I41806,I387665,I41823,I41831,I387650,I41848,I41680,I41879,I41896,I41692,I387662,I41936,I41701,I41958,I387671,I387659,I41975,I387653,I42001,I42018,I41704,I42040,I41689,I42071,I42088,I42105,I42122,I41698,I42153,I41686,I41695,I41683,I42239,I321237,I42265,I42273,I42290,I321234,I321249,I42307,I321231,I42333,I321228,I42350,I42358,I42375,I42207,I42406,I42423,I42219,I42463,I42228,I42485,I321243,I42502,I321246,I42528,I42545,I42231,I42567,I42216,I42598,I321240,I42615,I42632,I42649,I42225,I42680,I42213,I42222,I42210,I42766,I423758,I42792,I42800,I42817,I423755,I423761,I42834,I42860,I42877,I42885,I42902,I42734,I42933,I42950,I42746,I423764,I42990,I42755,I43012,I423767,I423776,I43029,I423770,I43055,I43072,I42758,I43094,I42743,I43125,I423773,I43142,I43159,I43176,I42752,I43207,I42740,I42749,I42737,I43293,I316922,I43319,I43327,I43344,I316913,I316931,I43361,I316910,I43387,I43404,I43412,I316916,I43429,I43261,I43460,I43477,I43273,I43517,I43282,I43539,I316928,I316919,I43556,I316934,I43582,I43599,I43285,I43621,I43270,I43652,I316925,I43669,I43686,I43703,I43279,I43734,I43267,I43276,I43264,I43820,I89394,I43846,I43854,I43871,I89388,I89382,I43888,I89403,I43914,I89400,I43931,I43939,I89397,I43956,I43788,I43987,I44004,I43800,I44044,I43809,I44066,I89385,I44083,I89406,I44109,I44126,I43812,I44148,I43797,I44179,I89391,I44196,I44213,I44230,I43806,I44261,I43794,I43803,I43791,I44347,I463184,I44373,I44381,I44398,I463199,I463178,I44415,I463181,I44441,I463202,I44458,I44466,I44483,I44315,I44514,I44531,I44327,I44571,I44336,I44593,I463190,I463187,I44610,I463193,I44636,I44653,I44339,I44675,I44324,I44706,I463196,I44723,I44740,I44757,I44333,I44788,I44321,I44330,I44318,I44874,I428807,I44900,I44908,I44925,I428804,I428810,I44942,I44968,I44985,I44993,I45010,I44842,I45041,I45058,I44854,I428813,I45098,I44863,I45120,I428816,I428825,I45137,I428819,I45163,I45180,I44866,I45202,I44851,I45233,I428822,I45250,I45267,I45284,I44860,I45315,I44848,I44857,I44845,I45401,I220948,I45427,I45435,I45452,I220969,I220963,I45469,I220945,I45495,I45512,I45520,I220957,I45537,I45369,I45568,I45585,I45381,I220954,I45625,I45390,I45647,I220960,I220951,I45664,I45690,I45707,I45393,I45729,I45378,I45760,I220966,I45777,I45794,I45811,I45387,I45842,I45375,I45384,I45372,I45928,I532742,I45954,I45962,I45979,I532748,I532766,I45996,I532763,I46022,I532760,I46039,I46047,I532754,I46064,I45896,I46095,I46112,I45908,I46152,I45917,I46174,I532757,I532745,I46191,I532769,I46217,I46234,I45920,I46256,I45905,I46287,I532751,I46304,I46321,I46338,I45914,I46369,I45902,I45911,I45899,I46455,I81659,I46481,I46489,I46506,I81653,I81647,I46523,I81668,I46549,I81665,I46566,I46574,I81662,I46591,I46423,I46622,I46639,I46435,I46679,I46444,I46701,I81650,I46718,I81671,I46744,I46761,I46447,I46783,I46432,I46814,I81656,I46831,I46848,I46865,I46441,I46896,I46429,I46438,I46426,I46982,I311720,I47008,I47016,I47033,I311711,I311729,I47050,I311708,I47076,I47093,I47101,I311714,I47118,I46950,I47149,I47166,I46962,I47206,I46971,I47228,I311726,I311717,I47245,I311732,I47271,I47288,I46974,I47310,I46959,I47341,I311723,I47358,I47375,I47392,I46968,I47423,I46956,I46965,I46953,I47509,I396700,I47535,I47543,I47560,I396718,I396712,I47577,I396691,I47603,I396709,I47620,I47628,I396694,I47645,I47477,I47676,I47693,I47489,I396706,I47733,I47498,I47755,I396715,I396703,I47772,I396697,I47798,I47815,I47501,I47837,I47486,I47868,I47885,I47902,I47919,I47495,I47950,I47483,I47492,I47480,I48036,I566567,I48062,I48070,I48087,I566561,I566582,I48104,I566558,I48130,I566579,I48147,I48155,I566576,I48172,I48004,I48203,I48220,I48016,I566564,I48260,I48025,I48282,I566573,I566570,I48299,I566555,I48325,I48342,I48028,I48364,I48013,I48395,I48412,I48429,I48446,I48022,I48477,I48010,I48019,I48007,I48563,I274150,I48589,I48597,I48614,I274141,I274159,I48631,I274138,I48657,I48674,I48682,I274144,I48699,I48531,I48730,I48747,I48543,I48787,I48552,I48809,I274156,I274147,I48826,I274162,I48852,I48869,I48555,I48891,I48540,I48922,I274153,I48939,I48956,I48973,I48549,I49004,I48537,I48546,I48534,I49090,I550502,I49116,I49124,I49141,I550496,I550517,I49158,I550493,I49184,I550514,I49201,I49209,I550511,I49226,I49058,I49257,I49274,I49070,I550499,I49314,I49079,I49336,I550508,I550505,I49353,I550490,I49379,I49396,I49082,I49418,I49067,I49449,I49466,I49483,I49500,I49076,I49531,I49064,I49073,I49061,I49617,I486882,I49643,I49651,I49668,I486897,I486876,I49685,I486879,I49711,I486900,I49728,I49736,I49753,I49585,I49784,I49801,I49597,I49841,I49606,I49863,I486888,I486885,I49880,I486891,I49906,I49923,I49609,I49945,I49594,I49976,I486894,I49993,I50010,I50027,I49603,I50058,I49591,I49600,I49588,I50147,I112460,I50173,I50181,I112457,I50207,I50215,I112454,I50232,I112466,I50249,I50124,I50280,I112475,I50118,I50311,I112472,I50328,I50345,I112451,I50362,I50379,I50396,I50133,I50130,I50136,I50455,I50472,I50489,I112463,I112478,I50515,I50115,I50546,I50554,I112469,I50139,I50585,I50602,I50619,I50121,I50650,I50667,I50112,I50127,I50742,I216197,I50768,I50776,I216203,I50802,I50810,I216185,I50827,I216209,I50844,I50719,I50875,I216200,I50713,I50906,I216191,I50923,I50940,I216194,I216188,I50957,I50974,I50991,I50728,I50725,I50731,I51050,I51067,I51084,I216206,I51110,I50710,I51141,I51149,I50734,I51180,I51197,I51214,I50716,I51245,I51262,I50707,I50722,I51337,I135121,I51363,I51371,I135118,I51397,I51405,I135115,I51422,I135127,I51439,I51314,I51470,I135136,I51308,I51501,I135133,I51518,I51535,I135112,I51552,I51569,I51586,I51323,I51320,I51326,I51645,I51662,I51679,I135124,I135139,I51705,I51305,I51736,I51744,I135130,I51329,I51775,I51792,I51809,I51311,I51840,I51857,I51302,I51317,I51932,I377963,I51958,I51966,I377984,I51992,I52000,I377966,I52017,I377957,I52034,I51909,I52065,I377969,I51903,I52096,I377960,I52113,I52130,I377978,I377981,I52147,I52164,I52181,I51918,I51915,I51921,I52240,I52257,I52274,I377972,I377975,I52300,I51900,I52331,I52339,I51924,I52370,I52387,I52404,I51906,I52435,I52452,I51897,I51912,I52527,I442373,I52553,I52561,I442370,I52587,I52595,I442379,I52612,I52629,I52504,I52660,I442382,I52498,I52691,I442376,I52708,I52725,I442391,I52742,I52759,I52776,I52513,I52510,I52516,I52835,I52852,I52869,I442394,I442388,I52895,I52495,I52926,I52934,I442385,I52519,I52965,I52982,I52999,I52501,I53030,I53047,I52492,I52507,I53122,I53148,I53156,I53182,I53190,I53207,I53224,I53099,I53255,I53093,I53286,I53303,I53320,I53337,I53354,I53371,I53108,I53105,I53111,I53430,I53447,I53464,I53490,I53090,I53521,I53529,I53114,I53560,I53577,I53594,I53096,I53625,I53642,I53087,I53102,I53717,I499595,I53743,I53751,I499592,I53777,I53785,I499601,I53802,I53819,I53694,I53850,I499604,I53688,I53881,I499598,I53898,I53915,I499613,I53932,I53949,I53966,I53703,I53700,I53706,I54025,I54042,I54059,I499616,I499610,I54085,I53685,I54116,I54124,I499607,I53709,I54155,I54172,I54189,I53691,I54220,I54237,I53682,I53697,I54309,I320707,I54335,I54352,I54301,I54374,I320701,I54400,I54408,I54425,I320719,I54442,I54459,I54476,I54493,I320713,I54510,I320704,I54527,I54277,I54558,I54575,I54592,I54609,I54289,I54283,I54654,I320716,I54298,I54292,I54699,I54716,I320722,I54733,I54750,I320710,I54776,I54784,I54286,I54280,I54838,I54846,I54295,I54904,I384432,I54930,I54947,I54896,I54969,I384441,I54995,I55003,I55020,I384429,I55037,I384420,I55054,I55071,I384426,I55088,I384444,I55105,I384417,I55122,I54872,I55153,I55170,I55187,I55204,I54884,I54878,I55249,I384423,I54893,I54887,I55294,I55311,I384435,I55328,I55345,I384438,I55371,I55379,I54881,I54875,I55433,I55441,I54890,I55499,I492656,I55525,I55542,I55491,I55564,I55590,I55598,I55615,I492659,I55632,I492671,I55649,I55666,I492677,I55683,I492668,I55700,I492674,I55717,I55467,I55748,I55765,I55782,I55799,I55479,I55473,I55844,I492665,I55488,I55482,I55889,I55906,I492662,I55923,I492680,I55940,I55966,I55974,I55476,I55470,I56028,I56036,I55485,I56094,I540396,I56120,I56137,I56086,I56159,I540387,I56185,I56193,I56210,I540381,I56227,I540375,I56244,I56261,I540402,I56278,I56295,I540399,I56312,I56062,I56343,I56360,I56377,I56394,I56074,I56068,I56439,I540384,I56083,I56077,I56484,I56501,I540390,I56518,I540393,I56535,I540378,I56561,I56569,I56071,I56065,I56623,I56631,I56080,I56689,I549321,I56715,I56732,I56681,I56754,I549312,I56780,I56788,I56805,I549306,I56822,I549300,I56839,I56856,I549327,I56873,I56890,I549324,I56907,I56657,I56938,I56955,I56972,I56989,I56669,I56663,I57034,I549309,I56678,I56672,I57079,I57096,I549315,I57113,I549318,I57130,I549303,I57156,I57164,I56666,I56660,I57218,I57226,I56675,I57284,I57310,I57327,I57276,I57349,I57375,I57383,I57400,I57417,I57434,I57451,I57468,I57485,I57502,I57252,I57533,I57550,I57567,I57584,I57264,I57258,I57629,I57273,I57267,I57674,I57691,I57708,I57725,I57751,I57759,I57261,I57255,I57813,I57821,I57270,I57879,I57905,I57922,I57871,I57944,I57970,I57978,I57995,I58012,I58029,I58046,I58063,I58080,I58097,I57847,I58128,I58145,I58162,I58179,I57859,I57853,I58224,I57868,I57862,I58269,I58286,I58303,I58320,I58346,I58354,I57856,I57850,I58408,I58416,I57865,I58474,I188720,I58500,I58517,I58466,I58539,I188708,I58565,I58573,I58590,I188717,I58607,I188714,I58624,I58641,I188705,I58658,I188711,I58675,I188696,I58692,I58442,I58723,I58740,I58757,I58774,I58454,I58448,I58819,I58463,I58457,I58864,I58881,I188702,I58898,I188699,I58915,I188723,I58941,I58949,I58451,I58445,I59003,I59011,I58460,I59069,I439480,I59095,I59112,I59061,I59134,I59160,I59168,I59185,I439483,I59202,I439495,I59219,I59236,I439501,I59253,I439492,I59270,I439498,I59287,I59037,I59318,I59335,I59352,I59369,I59049,I59043,I59414,I439489,I59058,I59052,I59459,I59476,I439486,I59493,I439504,I59510,I59536,I59544,I59046,I59040,I59598,I59606,I59055,I59664,I478206,I59690,I59707,I59729,I59755,I59763,I59780,I478209,I59797,I478221,I59814,I59831,I478227,I59848,I478218,I59865,I478224,I59882,I59913,I59930,I59947,I59964,I60009,I478215,I60054,I60071,I478212,I60088,I478230,I60105,I60131,I60139,I60193,I60201,I60259,I392184,I60285,I60302,I60251,I60324,I392193,I60350,I60358,I60375,I392181,I60392,I392172,I60409,I60426,I392178,I60443,I392196,I60460,I392169,I60477,I60227,I60508,I60525,I60542,I60559,I60239,I60233,I60604,I392175,I60248,I60242,I60649,I60666,I392187,I60683,I60700,I392190,I60726,I60734,I60236,I60230,I60788,I60796,I60245,I60854,I60880,I60897,I60846,I60919,I60945,I60953,I60970,I60987,I61004,I61021,I61038,I61055,I61072,I60822,I61103,I61120,I61137,I61154,I60834,I60828,I61199,I60843,I60837,I61244,I61261,I61278,I61295,I61321,I61329,I60831,I60825,I61383,I61391,I60840,I61449,I210842,I61475,I61492,I61441,I61514,I210836,I61540,I61548,I61565,I210851,I61582,I210848,I61599,I61616,I210839,I61633,I210830,I61650,I210833,I61667,I61417,I61698,I61715,I61732,I61749,I61429,I61423,I61794,I210854,I61438,I61432,I61839,I61856,I210845,I61873,I61890,I61916,I61924,I61426,I61420,I61978,I61986,I61435,I62044,I522375,I62070,I62087,I62036,I62109,I522387,I62135,I62143,I62160,I522381,I62177,I522393,I62194,I62211,I522378,I62228,I522390,I62245,I522372,I62262,I62012,I62293,I62310,I62327,I62344,I62024,I62018,I62389,I522384,I62033,I62027,I62434,I62451,I62468,I62485,I522396,I62511,I62519,I62021,I62015,I62573,I62581,I62030,I62639,I168048,I62665,I62682,I62631,I62704,I168036,I62730,I62738,I62755,I168045,I62772,I168042,I62789,I62806,I168033,I62823,I168039,I62840,I168024,I62857,I62607,I62888,I62905,I62922,I62939,I62619,I62613,I62984,I62628,I62622,I63029,I63046,I168030,I63063,I168027,I63080,I168051,I63106,I63114,I62616,I62610,I63168,I63176,I62625,I63234,I512292,I63260,I63277,I63226,I63299,I512277,I63325,I63333,I63350,I512295,I63367,I63384,I63401,I512298,I63418,I512289,I63435,I512286,I63452,I63202,I63483,I63500,I63517,I63534,I63214,I63208,I63579,I512283,I63223,I63217,I63624,I63641,I512274,I63658,I512280,I63675,I63701,I63709,I63211,I63205,I63763,I63771,I63220,I63829,I218577,I63855,I63872,I63821,I63894,I218571,I63920,I63928,I63945,I218586,I63962,I218583,I63979,I63996,I218574,I64013,I218565,I64030,I218568,I64047,I63797,I64078,I64095,I64112,I64129,I63809,I63803,I64174,I218589,I63818,I63812,I64219,I64236,I218580,I64253,I64270,I64296,I64304,I63806,I63800,I64358,I64366,I63815,I64424,I146706,I64450,I64467,I64416,I64489,I146721,I64515,I64523,I64540,I146718,I64557,I64574,I64591,I146715,I64608,I146730,I64625,I146727,I64642,I64392,I64673,I64690,I64707,I64724,I64404,I64398,I64769,I146724,I64413,I64407,I64814,I64831,I146712,I64848,I146733,I64865,I146709,I64891,I64899,I64401,I64395,I64953,I64961,I64410,I65019,I372804,I65045,I65062,I65011,I65084,I372813,I65110,I65118,I65135,I372801,I65152,I372792,I65169,I65186,I372798,I65203,I372816,I65220,I372789,I65237,I64987,I65268,I65285,I65302,I65319,I64999,I64993,I65364,I372795,I65008,I65002,I65409,I65426,I372807,I65443,I65460,I372810,I65486,I65494,I64996,I64990,I65548,I65556,I65005,I65614,I461444,I65640,I65657,I65606,I65679,I65705,I65713,I65730,I461447,I65747,I461459,I65764,I65781,I461465,I65798,I461456,I65815,I461462,I65832,I65582,I65863,I65880,I65897,I65914,I65594,I65588,I65959,I461453,I65603,I65597,I66004,I66021,I461450,I66038,I461468,I66055,I66081,I66089,I65591,I65585,I66143,I66151,I65600,I66209,I66235,I66252,I66201,I66274,I66300,I66308,I66325,I66342,I66359,I66376,I66393,I66410,I66427,I66177,I66458,I66475,I66492,I66509,I66189,I66183,I66554,I66198,I66192,I66599,I66616,I66633,I66650,I66676,I66684,I66186,I66180,I66738,I66746,I66195,I66804,I66830,I66847,I66796,I66869,I66895,I66903,I66920,I66937,I66954,I66971,I66988,I67005,I67022,I66772,I67053,I67070,I67087,I67104,I66784,I66778,I67149,I66793,I66787,I67194,I67211,I67228,I67245,I67271,I67279,I66781,I66775,I67333,I67341,I66790,I67399,I565981,I67425,I67442,I67391,I67464,I565972,I67490,I67498,I67515,I565966,I67532,I565960,I67549,I67566,I565987,I67583,I67600,I565984,I67617,I67367,I67648,I67665,I67682,I67699,I67379,I67373,I67744,I565969,I67388,I67382,I67789,I67806,I565975,I67823,I565978,I67840,I565963,I67866,I67874,I67376,I67370,I67928,I67936,I67385,I67994,I180560,I68020,I68037,I68059,I180548,I68085,I68093,I68110,I180557,I68127,I180554,I68144,I68161,I180545,I68178,I180551,I68195,I180536,I68212,I68243,I68260,I68277,I68294,I68339,I68384,I68401,I180542,I68418,I180539,I68435,I180563,I68461,I68469,I68523,I68531,I68589,I537421,I68615,I68632,I68581,I68654,I537412,I68680,I68688,I68705,I537406,I68722,I537400,I68739,I68756,I537427,I68773,I68790,I537424,I68807,I68557,I68838,I68855,I68872,I68889,I68569,I68563,I68934,I537409,I68578,I68572,I68979,I68996,I537415,I69013,I537418,I69030,I537403,I69056,I69064,I68566,I68560,I69118,I69126,I68575,I69184,I429929,I69210,I69227,I69249,I429938,I69275,I69283,I69300,I429932,I69317,I429926,I69334,I69351,I429941,I69368,I69385,I429935,I69402,I69433,I69450,I69467,I69484,I69529,I69574,I69591,I429947,I69608,I429944,I69625,I69651,I69659,I69713,I69721,I69779,I153030,I69805,I69822,I69844,I153045,I69870,I69878,I69895,I153042,I69912,I69929,I69946,I153039,I69963,I153054,I69980,I153051,I69997,I70028,I70045,I70062,I70079,I70124,I153048,I70169,I70186,I153036,I70203,I153057,I70220,I153033,I70246,I70254,I70308,I70316,I70374,I373450,I70400,I70417,I70366,I70439,I373459,I70465,I70473,I70490,I373447,I70507,I373438,I70524,I70541,I373444,I70558,I373462,I70575,I373435,I70592,I70342,I70623,I70640,I70657,I70674,I70354,I70348,I70719,I373441,I70363,I70357,I70764,I70781,I373453,I70798,I70815,I373456,I70841,I70849,I70351,I70345,I70903,I70911,I70360,I70969,I70995,I71012,I70961,I71034,I71060,I71068,I71085,I71102,I71119,I71136,I71153,I71170,I71187,I70937,I71218,I71235,I71252,I71269,I70949,I70943,I71314,I70958,I70952,I71359,I71376,I71393,I71410,I71436,I71444,I70946,I70940,I71498,I71506,I70955,I71564,I71590,I71607,I71556,I71629,I71655,I71663,I71680,I71697,I71714,I71731,I71748,I71765,I71782,I71532,I71813,I71830,I71847,I71864,I71544,I71538,I71909,I71553,I71547,I71954,I71971,I71988,I72005,I72031,I72039,I71541,I71535,I72093,I72101,I71550,I72159,I500170,I72185,I72202,I72151,I72224,I72250,I72258,I72275,I500173,I72292,I500185,I72309,I72326,I500191,I72343,I500182,I72360,I500188,I72377,I72127,I72408,I72425,I72442,I72459,I72139,I72133,I72504,I500179,I72148,I72142,I72549,I72566,I500176,I72583,I500194,I72600,I72626,I72634,I72136,I72130,I72688,I72696,I72145,I72754,I383140,I72780,I72797,I72746,I72819,I383149,I72845,I72853,I72870,I383137,I72887,I383128,I72904,I72921,I383134,I72938,I383152,I72955,I383125,I72972,I72722,I73003,I73020,I73037,I73054,I72734,I72728,I73099,I383131,I72743,I72737,I73144,I73161,I383143,I73178,I73195,I383146,I73221,I73229,I72731,I72725,I73283,I73291,I72740,I73349,I567766,I73375,I73392,I73341,I73414,I567757,I73440,I73448,I73465,I567751,I73482,I567745,I73499,I73516,I567772,I73533,I73550,I567769,I73567,I73317,I73598,I73615,I73632,I73649,I73329,I73323,I73694,I567754,I73338,I73332,I73739,I73756,I567760,I73773,I567763,I73790,I567748,I73816,I73824,I73326,I73320,I73878,I73886,I73335,I73944,I444104,I73970,I73987,I73936,I74009,I74035,I74043,I74060,I444107,I74077,I444119,I74094,I74111,I444125,I74128,I444116,I74145,I444122,I74162,I73912,I74193,I74210,I74227,I74244,I73924,I73918,I74289,I444113,I73933,I73927,I74334,I74351,I444110,I74368,I444128,I74385,I74411,I74419,I73921,I73915,I74473,I74481,I73930,I74539,I155665,I74565,I74582,I74531,I74604,I155680,I74630,I74638,I74655,I155677,I74672,I74689,I74706,I155674,I74723,I155689,I74740,I155686,I74757,I74507,I74788,I74805,I74822,I74839,I74519,I74513,I74884,I155683,I74528,I74522,I74929,I74946,I155671,I74963,I155692,I74980,I155668,I75006,I75014,I74516,I74510,I75068,I75076,I74525,I75134,I211437,I75160,I75177,I75126,I75199,I211431,I75225,I75233,I75250,I211446,I75267,I211443,I75284,I75301,I211434,I75318,I211425,I75335,I211428,I75352,I75102,I75383,I75400,I75417,I75434,I75114,I75108,I75479,I211449,I75123,I75117,I75524,I75541,I211440,I75558,I75575,I75601,I75609,I75111,I75105,I75663,I75671,I75120,I75729,I231381,I75755,I75772,I75721,I75794,I231372,I75820,I75828,I75845,I231390,I75862,I231387,I75879,I75896,I231366,I75913,I231369,I75930,I231378,I75947,I75697,I75978,I75995,I76012,I76029,I75709,I75703,I76074,I231384,I75718,I75712,I76119,I76136,I76153,I231375,I76170,I76196,I76204,I75706,I75700,I76258,I76266,I75715,I76324,I202512,I76350,I76367,I76316,I76389,I202506,I76415,I76423,I76440,I202521,I76457,I202518,I76474,I76491,I202509,I76508,I202500,I76525,I202503,I76542,I76292,I76573,I76590,I76607,I76624,I76304,I76298,I76669,I202524,I76313,I76307,I76714,I76731,I202515,I76748,I76765,I76791,I76799,I76301,I76295,I76853,I76861,I76310,I76919,I181104,I76945,I76962,I76911,I76984,I181092,I77010,I77018,I77035,I181101,I77052,I181098,I77069,I77086,I181089,I77103,I181095,I77120,I181080,I77137,I76887,I77168,I77185,I77202,I77219,I76899,I76893,I77264,I76908,I76902,I77309,I77326,I181086,I77343,I181083,I77360,I181107,I77386,I77394,I76896,I76890,I77448,I77456,I76905,I77514,I502500,I77540,I77557,I77506,I77579,I502485,I77605,I77613,I77630,I502503,I77647,I77664,I77681,I502506,I77698,I502497,I77715,I502494,I77732,I77482,I77763,I77780,I77797,I77814,I77494,I77488,I77859,I502491,I77503,I77497,I77904,I77921,I502482,I77938,I502488,I77955,I77981,I77989,I77491,I77485,I78043,I78051,I77500,I78109,I78135,I78152,I78101,I78174,I78200,I78208,I78225,I78242,I78259,I78276,I78293,I78310,I78327,I78077,I78358,I78375,I78392,I78409,I78089,I78083,I78454,I78098,I78092,I78499,I78516,I78533,I78550,I78576,I78584,I78086,I78080,I78638,I78646,I78095,I78704,I127734,I78730,I78747,I78696,I78769,I127749,I78795,I78803,I78820,I127746,I78837,I78854,I78871,I127743,I78888,I127758,I78905,I127755,I78922,I78672,I78953,I78970,I78987,I79004,I78684,I78678,I79049,I127752,I78693,I78687,I79094,I79111,I127740,I79128,I127761,I79145,I127737,I79171,I79179,I78681,I78675,I79233,I79241,I78690,I79299,I369574,I79325,I79342,I79291,I79364,I369583,I79390,I79398,I79415,I369571,I79432,I369562,I79449,I79466,I369568,I79483,I369586,I79500,I369559,I79517,I79267,I79548,I79565,I79582,I79599,I79279,I79273,I79644,I369565,I79288,I79282,I79689,I79706,I369577,I79723,I79740,I369580,I79766,I79774,I79276,I79270,I79828,I79836,I79285,I79894,I358651,I79920,I79937,I79886,I79959,I358645,I79985,I79993,I80010,I358663,I80027,I80044,I80061,I80078,I358657,I80095,I358648,I80112,I79862,I80143,I80160,I80177,I80194,I79874,I79868,I80239,I358660,I79883,I79877,I80284,I80301,I358666,I80318,I80335,I358654,I80361,I80369,I79871,I79865,I80423,I80431,I79880,I80489,I219767,I80515,I80532,I80481,I80554,I219761,I80580,I80588,I80605,I219776,I80622,I219773,I80639,I80656,I219764,I80673,I219755,I80690,I219758,I80707,I80457,I80738,I80755,I80772,I80789,I80469,I80463,I80834,I219779,I80478,I80472,I80879,I80896,I219770,I80913,I80930,I80956,I80964,I80466,I80460,I81018,I81026,I80475,I81084,I304784,I81110,I81127,I81076,I81149,I304781,I81175,I81183,I81200,I304787,I81217,I304772,I81234,I81251,I304775,I81268,I304796,I81285,I304793,I81302,I81052,I81333,I81350,I81367,I81384,I81064,I81058,I81429,I81073,I81067,I81474,I81491,I304778,I81508,I304790,I81525,I81551,I81559,I81061,I81055,I81613,I81621,I81070,I81679,I377326,I81705,I81722,I81744,I377335,I81770,I81778,I81795,I377323,I81812,I377314,I81829,I81846,I377320,I81863,I377338,I81880,I377311,I81897,I81928,I81945,I81962,I81979,I82024,I377317,I82069,I82086,I377329,I82103,I82120,I377332,I82146,I82154,I82208,I82216,I82274,I187088,I82300,I82317,I82266,I82339,I187076,I82365,I82373,I82390,I187085,I82407,I187082,I82424,I82441,I187073,I82458,I187079,I82475,I187064,I82492,I82242,I82523,I82540,I82557,I82574,I82254,I82248,I82619,I82263,I82257,I82664,I82681,I187070,I82698,I187067,I82715,I187091,I82741,I82749,I82251,I82245,I82803,I82811,I82260,I82869,I448150,I82895,I82912,I82861,I82934,I82960,I82968,I82985,I448153,I83002,I448165,I83019,I83036,I448171,I83053,I448162,I83070,I448168,I83087,I82837,I83118,I83135,I83152,I83169,I82849,I82843,I83214,I448159,I82858,I82852,I83259,I83276,I448156,I83293,I448174,I83310,I83336,I83344,I82846,I82840,I83398,I83406,I82855,I83464,I233115,I83490,I83507,I83456,I83529,I233106,I83555,I83563,I83580,I233124,I83597,I233121,I83614,I83631,I233100,I83648,I233103,I83665,I233112,I83682,I83432,I83713,I83730,I83747,I83764,I83444,I83438,I83809,I233118,I83453,I83447,I83854,I83871,I83888,I233109,I83905,I83931,I83939,I83441,I83435,I83993,I84001,I83450,I84059,I243519,I84085,I84102,I84051,I84124,I243510,I84150,I84158,I84175,I243528,I84192,I243525,I84209,I84226,I243504,I84243,I243507,I84260,I243516,I84277,I84027,I84308,I84325,I84342,I84359,I84039,I84033,I84404,I243522,I84048,I84042,I84449,I84466,I84483,I243513,I84500,I84526,I84534,I84036,I84030,I84588,I84596,I84045,I84654,I532208,I84680,I84697,I84646,I84719,I532181,I84745,I84753,I84770,I532205,I84787,I532202,I84804,I84821,I84838,I532199,I84855,I532187,I84872,I84622,I84903,I84920,I84937,I84954,I84634,I84628,I84999,I532193,I84643,I84637,I85044,I85061,I532196,I85078,I532184,I85095,I532190,I85121,I85129,I84631,I84625,I85183,I85191,I84640,I85249,I468958,I85275,I85292,I85241,I85314,I85340,I85348,I85365,I468961,I85382,I468973,I85399,I85416,I468979,I85433,I468970,I85450,I468976,I85467,I85217,I85498,I85515,I85532,I85549,I85229,I85223,I85594,I468967,I85238,I85232,I85639,I85656,I468964,I85673,I468982,I85690,I85716,I85724,I85226,I85220,I85778,I85786,I85235,I85844,I514468,I85870,I85887,I85836,I85909,I514453,I85935,I85943,I85960,I514471,I85977,I85994,I86011,I514474,I86028,I514465,I86045,I514462,I86062,I85812,I86093,I86110,I86127,I86144,I85824,I85818,I86189,I514459,I85833,I85827,I86234,I86251,I514450,I86268,I514456,I86285,I86311,I86319,I85821,I85815,I86373,I86381,I85830,I86439,I150395,I86465,I86482,I86431,I86504,I150410,I86530,I86538,I86555,I150407,I86572,I86589,I86606,I150404,I86623,I150419,I86640,I150416,I86657,I86407,I86688,I86705,I86722,I86739,I86419,I86413,I86784,I150413,I86428,I86422,I86829,I86846,I150401,I86863,I150422,I86880,I150398,I86906,I86914,I86416,I86410,I86968,I86976,I86425,I87034,I206082,I87060,I87077,I87026,I87099,I206076,I87125,I87133,I87150,I206091,I87167,I206088,I87184,I87201,I206079,I87218,I206070,I87235,I206073,I87252,I87002,I87283,I87300,I87317,I87334,I87014,I87008,I87379,I206094,I87023,I87017,I87424,I87441,I206085,I87458,I87475,I87501,I87509,I87011,I87005,I87563,I87571,I87020,I87629,I87655,I87672,I87621,I87694,I87720,I87728,I87745,I87762,I87779,I87796,I87813,I87830,I87847,I87597,I87878,I87895,I87912,I87929,I87609,I87603,I87974,I87618,I87612,I88019,I88036,I88053,I88070,I88096,I88104,I87606,I87600,I88158,I88166,I87615,I88224,I395414,I88250,I88267,I88216,I88289,I395423,I88315,I88323,I88340,I395411,I88357,I395402,I88374,I88391,I395408,I88408,I395426,I88425,I395399,I88442,I88192,I88473,I88490,I88507,I88524,I88204,I88198,I88569,I395405,I88213,I88207,I88614,I88631,I395417,I88648,I88665,I395420,I88691,I88699,I88201,I88195,I88753,I88761,I88210,I88819,I288600,I88845,I88862,I88811,I88884,I288597,I88910,I88918,I88935,I288603,I88952,I288588,I88969,I88986,I288591,I89003,I288612,I89020,I288609,I89037,I88787,I89068,I89085,I89102,I89119,I88799,I88793,I89164,I88808,I88802,I89209,I89226,I288594,I89243,I288606,I89260,I89286,I89294,I88796,I88790,I89348,I89356,I88805,I89414,I170224,I89440,I89457,I89479,I170212,I89505,I89513,I89530,I170221,I89547,I170218,I89564,I89581,I170209,I89598,I170215,I89615,I170200,I89632,I89663,I89680,I89697,I89714,I89759,I89804,I89821,I170206,I89838,I170203,I89855,I170227,I89881,I89889,I89943,I89951,I90009,I442948,I90035,I90052,I90001,I90074,I90100,I90108,I90125,I442951,I90142,I442963,I90159,I90176,I442969,I90193,I442960,I90210,I442966,I90227,I89977,I90258,I90275,I90292,I90309,I89989,I89983,I90354,I442957,I89998,I89992,I90399,I90416,I442954,I90433,I442972,I90450,I90476,I90484,I89986,I89980,I90538,I90546,I89995,I90604,I90630,I90647,I90596,I90669,I90695,I90703,I90720,I90737,I90754,I90771,I90788,I90805,I90822,I90572,I90853,I90870,I90887,I90904,I90584,I90578,I90949,I90593,I90587,I90994,I91011,I91028,I91045,I91071,I91079,I90581,I90575,I91133,I91141,I90590,I91199,I330193,I91225,I91242,I91191,I91264,I330187,I91290,I91298,I91315,I330205,I91332,I91349,I91366,I91383,I330199,I91400,I330190,I91417,I91167,I91448,I91465,I91482,I91499,I91179,I91173,I91544,I330202,I91188,I91182,I91589,I91606,I330208,I91623,I91640,I330196,I91666,I91674,I91176,I91170,I91728,I91736,I91185,I91794,I91820,I91837,I91786,I91859,I91885,I91893,I91910,I91927,I91944,I91961,I91978,I91995,I92012,I91762,I92043,I92060,I92077,I92094,I91774,I91768,I92139,I91783,I91777,I92184,I92201,I92218,I92235,I92261,I92269,I91771,I91765,I92323,I92331,I91780,I92389,I323869,I92415,I92432,I92381,I92454,I323863,I92480,I92488,I92505,I323881,I92522,I92539,I92556,I92573,I323875,I92590,I323866,I92607,I92357,I92638,I92655,I92672,I92689,I92369,I92363,I92734,I323878,I92378,I92372,I92779,I92796,I323884,I92813,I92830,I323872,I92856,I92864,I92366,I92360,I92918,I92926,I92375,I92984,I366990,I93010,I93027,I93049,I366999,I93075,I93083,I93100,I366987,I93117,I366978,I93134,I93151,I366984,I93168,I367002,I93185,I366975,I93202,I93233,I93250,I93267,I93284,I93329,I366981,I93374,I93391,I366993,I93408,I93425,I366996,I93451,I93459,I93513,I93521,I93579,I475316,I93605,I93622,I93571,I93644,I93670,I93678,I93695,I475319,I93712,I475331,I93729,I93746,I475337,I93763,I475328,I93780,I475334,I93797,I93547,I93828,I93845,I93862,I93879,I93559,I93553,I93924,I475325,I93568,I93562,I93969,I93986,I475322,I94003,I475340,I94020,I94046,I94054,I93556,I93550,I94108,I94116,I93565,I94174,I418709,I94200,I94217,I94239,I418718,I94265,I94273,I94290,I418712,I94307,I418706,I94324,I94341,I418721,I94358,I94375,I418715,I94392,I94423,I94440,I94457,I94474,I94519,I94564,I94581,I418727,I94598,I418724,I94615,I94641,I94649,I94703,I94711,I94769,I131423,I94795,I94812,I94761,I94834,I131438,I94860,I94868,I94885,I131435,I94902,I94919,I94936,I131432,I94953,I131447,I94970,I131444,I94987,I94737,I95018,I95035,I95052,I95069,I94749,I94743,I95114,I131441,I94758,I94752,I95159,I95176,I131429,I95193,I131450,I95210,I131426,I95236,I95244,I94746,I94740,I95298,I95306,I94755,I95364,I321761,I95390,I95407,I95356,I95429,I321755,I95455,I95463,I95480,I321773,I95497,I95514,I95531,I95548,I321767,I95565,I321758,I95582,I95332,I95613,I95630,I95647,I95664,I95344,I95338,I95709,I321770,I95353,I95347,I95754,I95771,I321776,I95788,I95805,I321764,I95831,I95839,I95341,I95335,I95893,I95901,I95350,I95959,I213222,I95985,I96002,I95951,I96024,I213216,I96050,I96058,I96075,I213231,I96092,I213228,I96109,I96126,I213219,I96143,I213210,I96160,I213213,I96177,I95927,I96208,I96225,I96242,I96259,I95939,I95933,I96304,I213234,I95948,I95942,I96349,I96366,I213225,I96383,I96400,I96426,I96434,I95936,I95930,I96488,I96496,I95945,I96554,I96580,I96597,I96619,I96645,I96653,I96670,I96687,I96704,I96721,I96738,I96755,I96772,I96803,I96820,I96837,I96854,I96899,I96944,I96961,I96978,I96995,I97021,I97029,I97083,I97091,I97149,I486298,I97175,I97192,I97141,I97214,I97240,I97248,I97265,I486301,I97282,I486313,I97299,I97316,I486319,I97333,I486310,I97350,I486316,I97367,I97117,I97398,I97415,I97432,I97449,I97129,I97123,I97494,I486307,I97138,I97132,I97539,I97556,I486304,I97573,I486322,I97590,I97616,I97624,I97126,I97120,I97678,I97686,I97135,I97744,I174032,I97770,I97787,I97736,I97809,I174020,I97835,I97843,I97860,I174029,I97877,I174026,I97894,I97911,I174017,I97928,I174023,I97945,I174008,I97962,I97712,I97993,I98010,I98027,I98044,I97724,I97718,I98089,I97733,I97727,I98134,I98151,I174014,I98168,I174011,I98185,I174035,I98211,I98219,I97721,I97715,I98273,I98281,I97730,I98339,I98365,I98382,I98404,I98430,I98438,I98455,I98472,I98489,I98506,I98523,I98540,I98557,I98588,I98605,I98622,I98639,I98684,I98729,I98746,I98763,I98780,I98806,I98814,I98868,I98876,I98934,I98960,I98977,I98926,I98999,I99025,I99033,I99050,I99067,I99084,I99101,I99118,I99135,I99152,I98902,I99183,I99200,I99217,I99234,I98914,I98908,I99279,I98923,I98917,I99324,I99341,I99358,I99375,I99401,I99409,I98911,I98905,I99463,I99471,I98920,I99529,I513380,I99555,I99572,I99521,I99594,I513365,I99620,I99628,I99645,I513383,I99662,I99679,I99696,I513386,I99713,I513377,I99730,I513374,I99747,I99497,I99778,I99795,I99812,I99829,I99509,I99503,I99874,I513371,I99518,I99512,I99919,I99936,I513362,I99953,I513368,I99970,I99996,I100004,I99506,I99500,I100058,I100066,I99515,I100124,I111924,I100150,I100167,I100116,I100189,I111939,I100215,I100223,I100240,I111936,I100257,I100274,I100291,I111933,I100308,I111948,I100325,I111945,I100342,I100092,I100373,I100390,I100407,I100424,I100104,I100098,I100469,I111942,I100113,I100107,I100514,I100531,I111930,I100548,I111951,I100565,I111927,I100591,I100599,I100101,I100095,I100653,I100661,I100110,I100719,I100745,I100762,I100711,I100784,I100810,I100818,I100835,I100852,I100869,I100886,I100903,I100920,I100937,I100687,I100968,I100985,I101002,I101019,I100699,I100693,I101064,I100708,I100702,I101109,I101126,I101143,I101160,I101186,I101194,I100696,I100690,I101248,I101256,I100705,I101314,I134058,I101340,I101357,I101306,I101379,I134073,I101405,I101413,I101430,I134070,I101447,I101464,I101481,I134067,I101498,I134082,I101515,I134079,I101532,I101282,I101563,I101580,I101597,I101614,I101294,I101288,I101659,I134076,I101303,I101297,I101704,I101721,I134064,I101738,I134085,I101755,I134061,I101781,I101789,I101291,I101285,I101843,I101851,I101300,I101909,I493234,I101935,I101952,I101974,I102000,I102008,I102025,I493237,I102042,I493249,I102059,I102076,I493255,I102093,I493246,I102110,I493252,I102127,I102158,I102175,I102192,I102209,I102254,I493243,I102299,I102316,I493240,I102333,I493258,I102350,I102376,I102384,I102438,I102446,I102504,I494390,I102530,I102547,I102496,I102569,I102595,I102603,I102620,I494393,I102637,I494405,I102654,I102671,I494411,I102688,I494402,I102705,I494408,I102722,I102472,I102753,I102770,I102787,I102804,I102484,I102478,I102849,I494399,I102493,I102487,I102894,I102911,I494396,I102928,I494414,I102945,I102971,I102979,I102481,I102475,I103033,I103041,I102490,I103099,I516100,I103125,I103142,I103091,I103164,I516085,I103190,I103198,I103215,I516103,I103232,I103249,I103266,I516106,I103283,I516097,I103300,I516094,I103317,I103067,I103348,I103365,I103382,I103399,I103079,I103073,I103444,I516091,I103088,I103082,I103489,I103506,I516082,I103523,I516088,I103540,I103566,I103574,I103076,I103070,I103628,I103636,I103085,I103694,I407042,I103720,I103737,I103686,I103759,I407051,I103785,I103793,I103810,I407039,I103827,I407030,I103844,I103861,I407036,I103878,I407054,I103895,I407027,I103912,I103662,I103943,I103960,I103977,I103994,I103674,I103668,I104039,I407033,I103683,I103677,I104084,I104101,I407045,I104118,I104135,I407048,I104161,I104169,I103671,I103665,I104223,I104231,I103680,I104289,I167504,I104315,I104332,I104281,I104354,I167492,I104380,I104388,I104405,I167501,I104422,I167498,I104439,I104456,I167489,I104473,I167495,I104490,I167480,I104507,I104257,I104538,I104555,I104572,I104589,I104269,I104263,I104634,I104278,I104272,I104679,I104696,I167486,I104713,I167483,I104730,I167507,I104756,I104764,I104266,I104260,I104818,I104826,I104275,I104884,I448728,I104910,I104927,I104876,I104949,I104975,I104983,I105000,I448731,I105017,I448743,I105034,I105051,I448749,I105068,I448740,I105085,I448746,I105102,I104852,I105133,I105150,I105167,I105184,I104864,I104858,I105229,I448737,I104873,I104867,I105274,I105291,I448734,I105308,I448752,I105325,I105351,I105359,I104861,I104855,I105413,I105421,I104870,I105479,I339679,I105505,I105522,I105471,I105544,I339673,I105570,I105578,I105595,I339691,I105612,I105629,I105646,I105663,I339685,I105680,I339676,I105697,I105447,I105728,I105745,I105762,I105779,I105459,I105453,I105824,I339688,I105468,I105462,I105869,I105886,I339694,I105903,I105920,I339682,I105946,I105954,I105456,I105450,I106008,I106016,I105465,I106074,I282242,I106100,I106117,I106066,I106139,I282239,I106165,I106173,I106190,I282245,I106207,I282230,I106224,I106241,I282233,I106258,I282254,I106275,I282251,I106292,I106042,I106323,I106340,I106357,I106374,I106054,I106048,I106419,I106063,I106057,I106464,I106481,I282236,I106498,I282248,I106515,I106541,I106549,I106051,I106045,I106603,I106611,I106060,I106669,I315188,I106695,I106712,I106661,I106734,I315185,I106760,I106768,I106785,I315191,I106802,I315176,I106819,I106836,I315179,I106853,I315200,I106870,I315197,I106887,I106637,I106918,I106935,I106952,I106969,I106649,I106643,I107014,I106658,I106652,I107059,I107076,I315182,I107093,I315194,I107110,I107136,I107144,I106646,I106640,I107198,I107206,I106655,I107264,I279930,I107290,I107307,I107256,I107329,I279927,I107355,I107363,I107380,I279933,I107397,I279918,I107414,I107431,I279921,I107448,I279942,I107465,I279939,I107482,I107232,I107513,I107530,I107547,I107564,I107244,I107238,I107609,I107253,I107247,I107654,I107671,I279924,I107688,I279936,I107705,I107731,I107739,I107241,I107235,I107793,I107801,I107250,I107859,I173488,I107885,I107902,I107851,I107924,I173476,I107950,I107958,I107975,I173485,I107992,I173482,I108009,I108026,I173473,I108043,I173479,I108060,I173464,I108077,I107827,I108108,I108125,I108142,I108159,I107839,I107833,I108204,I107848,I107842,I108249,I108266,I173470,I108283,I173467,I108300,I173491,I108326,I108334,I107836,I107830,I108388,I108396,I107845,I108454,I432173,I108480,I108497,I108446,I108519,I432182,I108545,I108553,I108570,I432176,I108587,I432170,I108604,I108621,I432185,I108638,I108655,I432179,I108672,I108422,I108703,I108720,I108737,I108754,I108434,I108428,I108799,I108443,I108437,I108844,I108861,I432191,I108878,I432188,I108895,I108921,I108929,I108431,I108425,I108983,I108991,I108440,I109049,I548131,I109075,I109092,I109114,I548122,I109140,I109148,I109165,I548116,I109182,I548110,I109199,I109216,I548137,I109233,I109250,I548134,I109267,I109298,I109315,I109332,I109349,I109394,I548119,I109439,I109456,I548125,I109473,I548128,I109490,I548113,I109516,I109524,I109578,I109586,I109644,I398644,I109670,I109687,I109636,I109709,I398653,I109735,I109743,I109760,I398641,I109777,I398632,I109794,I109811,I398638,I109828,I398656,I109845,I398629,I109862,I109612,I109893,I109910,I109927,I109944,I109624,I109618,I109989,I398635,I109633,I109627,I110034,I110051,I398647,I110068,I110085,I398650,I110111,I110119,I109621,I109615,I110173,I110181,I109630,I110239,I234271,I110265,I110282,I110231,I110304,I234262,I110330,I110338,I110355,I234280,I110372,I234277,I110389,I110406,I234256,I110423,I234259,I110440,I234268,I110457,I110207,I110488,I110505,I110522,I110539,I110219,I110213,I110584,I234274,I110228,I110222,I110629,I110646,I110663,I234265,I110680,I110706,I110714,I110216,I110210,I110768,I110776,I110225,I110834,I168592,I110860,I110877,I110826,I110899,I168580,I110925,I110933,I110950,I168589,I110967,I168586,I110984,I111001,I168577,I111018,I168583,I111035,I168568,I111052,I110802,I111083,I111100,I111117,I111134,I110814,I110808,I111179,I110823,I110817,I111224,I111241,I168574,I111258,I168571,I111275,I168595,I111301,I111309,I110811,I110805,I111363,I111371,I110820,I111432,I265480,I111458,I111466,I265471,I265486,I111483,I265492,I111509,I111400,I111531,I265477,I111557,I111565,I111582,I111608,I111424,I111630,I111406,I265474,I111670,I111687,I111695,I111712,I111409,I111743,I265468,I265483,I111760,I111786,I111794,I111397,I111415,I111839,I265489,I111856,I111418,I111403,I111412,I111421,I111959,I217378,I111985,I111993,I217390,I112010,I217375,I112036,I112058,I217399,I112084,I112092,I217396,I112109,I112135,I112157,I217387,I112197,I112214,I112222,I112239,I112270,I217384,I112287,I217393,I112313,I112321,I112366,I217381,I112383,I112486,I426563,I112512,I112520,I426560,I112537,I426572,I112563,I112585,I112611,I112619,I426578,I112636,I112662,I112684,I426566,I112724,I112741,I112749,I112766,I112797,I426575,I426581,I112814,I112840,I112848,I112893,I426569,I112910,I113013,I113039,I113047,I113064,I113090,I112981,I113112,I113138,I113146,I113163,I113189,I113005,I113211,I112987,I113251,I113268,I113276,I113293,I112990,I113324,I113341,I113367,I113375,I112978,I112996,I113420,I113437,I112999,I112984,I112993,I113002,I113540,I162596,I113566,I113574,I162608,I162587,I113591,I162611,I113617,I113508,I113639,I162602,I113665,I113673,I162584,I113690,I113716,I113532,I113738,I113514,I162599,I113778,I113795,I113803,I113820,I113517,I113851,I162590,I113868,I162593,I113894,I113902,I113505,I113523,I113947,I162605,I113964,I113526,I113511,I113520,I113529,I114067,I342838,I114093,I114101,I342841,I342835,I114118,I342847,I114144,I114035,I114166,I342850,I114192,I114200,I114217,I114243,I114059,I114265,I114041,I342853,I114305,I114322,I114330,I114347,I114044,I114378,I342844,I114395,I114421,I114429,I114032,I114050,I114474,I342856,I114491,I114053,I114038,I114047,I114056,I114594,I317500,I114620,I114628,I317491,I317506,I114645,I317512,I114671,I114562,I114693,I317497,I114719,I114727,I114744,I114770,I114586,I114792,I114568,I317494,I114832,I114849,I114857,I114874,I114571,I114905,I317488,I317503,I114922,I114948,I114956,I114559,I114577,I115001,I317509,I115018,I114580,I114565,I114574,I114583,I115121,I415343,I115147,I115155,I415340,I115172,I415352,I115198,I115089,I115220,I115246,I115254,I415358,I115271,I115297,I115113,I115319,I115095,I415346,I115359,I115376,I115384,I115401,I115098,I115432,I415355,I415361,I115449,I115475,I115483,I115086,I115104,I115528,I415349,I115545,I115107,I115092,I115101,I115110,I115648,I251611,I115674,I115682,I251596,I251599,I115699,I251614,I115725,I115616,I115747,I251608,I115773,I115781,I115798,I115824,I115640,I115846,I115622,I251605,I115886,I115903,I115911,I115928,I115625,I115959,I251620,I115976,I251617,I116002,I116010,I115613,I115631,I116055,I251602,I116072,I115634,I115619,I115628,I115637,I116175,I412844,I116201,I116209,I412841,I412859,I116226,I412850,I116252,I116143,I116274,I412865,I116300,I116308,I412847,I116325,I116351,I116167,I116373,I116149,I412853,I116413,I116430,I116438,I116455,I116152,I116486,I412868,I116503,I412856,I116529,I116537,I116140,I116158,I116582,I412862,I116599,I116161,I116146,I116155,I116164,I116702,I239473,I116728,I116736,I239458,I239461,I116753,I239476,I116779,I116670,I116801,I239470,I116827,I116835,I116852,I116878,I116694,I116900,I116676,I239467,I116940,I116957,I116965,I116982,I116679,I117013,I239482,I117030,I239479,I117056,I117064,I116667,I116685,I117109,I239464,I117126,I116688,I116673,I116682,I116691,I117229,I394110,I117255,I117263,I394107,I394125,I117280,I394116,I117306,I117197,I117328,I394131,I117354,I117362,I394113,I117379,I117405,I117221,I117427,I117203,I394119,I117467,I117484,I117492,I117509,I117206,I117540,I394134,I117557,I394122,I117583,I117591,I117194,I117212,I117636,I394128,I117653,I117215,I117200,I117209,I117218,I117756,I567171,I117782,I117790,I567150,I117807,I567177,I117833,I117724,I117855,I567165,I117881,I117889,I567168,I117906,I117932,I117748,I117954,I117730,I567159,I117994,I118011,I118019,I118036,I117733,I118067,I567156,I567153,I118084,I567174,I118110,I118118,I117721,I117739,I118163,I567162,I118180,I117742,I117727,I117736,I117745,I118283,I541586,I118309,I118317,I541565,I118334,I541592,I118360,I118251,I118382,I541580,I118408,I118416,I541583,I118433,I118459,I118275,I118481,I118257,I541574,I118521,I118538,I118546,I118563,I118260,I118594,I541571,I541568,I118611,I541589,I118637,I118645,I118248,I118266,I118690,I541577,I118707,I118269,I118254,I118263,I118272,I118810,I182180,I118836,I118844,I182192,I182171,I118861,I182195,I118887,I118778,I118909,I182186,I118935,I118943,I182168,I118960,I118986,I118802,I119008,I118784,I182183,I119048,I119065,I119073,I119090,I118787,I119121,I182174,I119138,I182177,I119164,I119172,I118775,I118793,I119217,I182189,I119234,I118796,I118781,I118790,I118799,I119337,I119363,I119371,I119388,I119414,I119305,I119436,I119462,I119470,I119487,I119513,I119329,I119535,I119311,I119575,I119592,I119600,I119617,I119314,I119648,I119665,I119691,I119699,I119302,I119320,I119744,I119761,I119323,I119308,I119317,I119326,I119864,I249299,I119890,I119898,I249284,I249287,I119915,I249302,I119941,I119832,I119963,I249296,I119989,I119997,I120014,I120040,I119856,I120062,I119838,I249293,I120102,I120119,I120127,I120144,I119841,I120175,I249308,I120192,I249305,I120218,I120226,I119829,I119847,I120271,I249290,I120288,I119850,I119835,I119844,I119853,I120391,I333879,I120417,I120425,I333882,I333876,I120442,I333888,I120468,I120359,I120490,I333891,I120516,I120524,I120541,I120567,I120383,I120589,I120365,I333894,I120629,I120646,I120654,I120671,I120368,I120702,I333885,I120719,I120745,I120753,I120356,I120374,I120798,I333897,I120815,I120377,I120362,I120371,I120380,I120918,I522965,I120944,I120952,I522962,I522953,I120969,I522950,I120995,I121017,I522959,I121043,I121051,I522968,I121068,I121094,I121116,I522971,I121156,I121173,I121181,I121198,I121229,I522956,I121246,I522974,I121272,I121280,I121325,I121342,I121445,I121471,I121479,I121496,I121522,I121413,I121544,I121570,I121578,I121595,I121621,I121437,I121643,I121419,I121683,I121700,I121708,I121725,I121422,I121756,I121773,I121799,I121807,I121410,I121428,I121852,I121869,I121431,I121416,I121425,I121434,I121972,I481096,I121998,I122006,I481111,I122023,I481114,I122049,I121940,I122071,I481120,I122097,I122105,I481102,I122122,I122148,I121964,I122170,I121946,I481099,I122210,I122227,I122235,I122252,I121949,I122283,I481105,I122300,I481117,I122326,I122334,I121937,I121955,I122379,I481108,I122396,I121958,I121943,I121952,I121961,I122499,I350216,I122525,I122533,I350219,I350213,I122550,I350225,I122576,I122467,I122598,I350228,I122624,I122632,I122649,I122675,I122491,I122697,I122473,I350231,I122737,I122754,I122762,I122779,I122476,I122810,I350222,I122827,I122853,I122861,I122464,I122482,I122906,I350234,I122923,I122485,I122470,I122479,I122488,I123026,I204883,I123052,I123060,I204895,I123077,I204880,I123103,I122994,I123125,I204904,I123151,I123159,I204901,I123176,I123202,I123018,I123224,I123000,I204892,I123264,I123281,I123289,I123306,I123003,I123337,I204889,I123354,I204898,I123380,I123388,I122991,I123009,I123433,I204886,I123450,I123012,I122997,I123006,I123015,I123553,I510116,I123579,I123587,I510098,I510122,I123604,I510113,I123630,I123521,I123652,I510119,I123678,I123686,I510107,I123703,I123729,I123545,I123751,I123527,I123791,I123808,I123816,I123833,I123530,I123864,I510104,I510101,I123881,I510110,I123907,I123915,I123518,I123536,I123960,I123977,I123539,I123524,I123533,I123542,I124080,I325447,I124106,I124114,I325450,I325444,I124131,I325456,I124157,I124048,I124179,I325459,I124205,I124213,I124230,I124256,I124072,I124278,I124054,I325462,I124318,I124335,I124343,I124360,I124057,I124391,I325453,I124408,I124434,I124442,I124045,I124063,I124487,I325465,I124504,I124066,I124051,I124060,I124069,I124607,I343892,I124633,I124641,I343895,I343889,I124658,I343901,I124684,I124575,I124706,I343904,I124732,I124740,I124757,I124783,I124599,I124805,I124581,I343907,I124845,I124862,I124870,I124887,I124584,I124918,I343898,I124935,I124961,I124969,I124572,I124590,I125014,I343910,I125031,I124593,I124578,I124587,I124596,I125134,I529901,I125160,I125168,I529898,I529889,I125185,I529886,I125211,I125102,I125233,I529895,I125259,I125267,I529904,I125284,I125310,I125126,I125332,I125108,I529907,I125372,I125389,I125397,I125414,I125111,I125445,I529892,I125462,I529910,I125488,I125496,I125099,I125117,I125541,I125558,I125120,I125105,I125114,I125123,I125661,I328082,I125687,I125695,I328085,I328079,I125712,I328091,I125738,I125629,I125760,I328094,I125786,I125794,I125811,I125837,I125653,I125859,I125635,I328097,I125899,I125916,I125924,I125941,I125638,I125972,I328088,I125989,I126015,I126023,I125626,I125644,I126068,I328100,I126085,I125647,I125632,I125641,I125650,I126188,I551701,I126214,I126222,I551680,I126239,I551707,I126265,I126156,I126287,I551695,I126313,I126321,I551698,I126338,I126364,I126180,I126386,I126162,I551689,I126426,I126443,I126451,I126468,I126165,I126499,I551686,I551683,I126516,I551704,I126542,I126550,I126153,I126171,I126595,I551692,I126612,I126174,I126159,I126168,I126177,I126715,I161508,I126741,I126749,I161520,I161499,I126766,I161523,I126792,I126683,I126814,I161514,I126840,I126848,I161496,I126865,I126891,I126707,I126913,I126689,I161511,I126953,I126970,I126978,I126995,I126692,I127026,I161502,I127043,I161505,I127069,I127077,I126680,I126698,I127122,I161517,I127139,I126701,I126686,I126695,I126704,I127242,I205478,I127268,I127276,I205490,I127293,I205475,I127319,I127210,I127341,I205499,I127367,I127375,I205496,I127392,I127418,I127234,I127440,I127216,I205487,I127480,I127497,I127505,I127522,I127219,I127553,I205484,I127570,I205493,I127596,I127604,I127207,I127225,I127649,I205481,I127666,I127228,I127213,I127222,I127231,I127769,I127795,I127803,I127820,I127846,I127868,I127894,I127902,I127919,I127945,I127967,I128007,I128024,I128032,I128049,I128080,I128097,I128123,I128131,I128176,I128193,I128296,I177284,I128322,I128330,I177296,I177275,I128347,I177299,I128373,I128264,I128395,I177290,I128421,I128429,I177272,I128446,I128472,I128288,I128494,I128270,I177287,I128534,I128551,I128559,I128576,I128273,I128607,I177278,I128624,I177281,I128650,I128658,I128261,I128279,I128703,I177293,I128720,I128282,I128267,I128276,I128285,I128823,I356013,I128849,I128857,I356016,I356010,I128874,I356022,I128900,I128791,I128922,I356025,I128948,I128956,I128973,I128999,I128815,I129021,I128797,I356028,I129061,I129078,I129086,I129103,I128800,I129134,I356019,I129151,I129177,I129185,I128788,I128806,I129230,I356031,I129247,I128809,I128794,I128803,I128812,I129350,I129376,I129384,I129401,I129427,I129318,I129449,I129475,I129483,I129500,I129526,I129342,I129548,I129324,I129588,I129605,I129613,I129630,I129327,I129661,I129678,I129704,I129712,I129315,I129333,I129757,I129774,I129336,I129321,I129330,I129339,I129877,I129903,I129911,I129928,I129954,I129845,I129976,I130002,I130010,I130027,I130053,I129869,I130075,I129851,I130115,I130132,I130140,I130157,I129854,I130188,I130205,I130231,I130239,I129842,I129860,I130284,I130301,I129863,I129848,I129857,I129866,I130404,I433295,I130430,I130438,I433292,I130455,I433304,I130481,I130372,I130503,I130529,I130537,I433310,I130554,I130580,I130396,I130602,I130378,I433298,I130642,I130659,I130667,I130684,I130381,I130715,I433307,I433313,I130732,I130758,I130766,I130369,I130387,I130811,I433301,I130828,I130390,I130375,I130384,I130393,I130931,I341257,I130957,I130965,I341260,I341254,I130982,I341266,I131008,I130899,I131030,I341269,I131056,I131064,I131081,I131107,I130923,I131129,I130905,I341272,I131169,I131186,I131194,I131211,I130908,I131242,I341263,I131259,I131285,I131293,I130896,I130914,I131338,I341275,I131355,I130917,I130902,I130911,I130920,I131458,I362456,I131484,I131492,I362453,I362471,I131509,I362462,I131535,I131557,I362477,I131583,I131591,I362459,I131608,I131634,I131656,I362465,I131696,I131713,I131721,I131738,I131769,I362480,I131786,I362468,I131812,I131820,I131865,I362474,I131882,I131985,I381836,I132011,I132019,I381833,I381851,I132036,I381842,I132062,I131953,I132084,I381857,I132110,I132118,I381839,I132135,I132161,I131977,I132183,I131959,I381845,I132223,I132240,I132248,I132265,I131962,I132296,I381860,I132313,I381848,I132339,I132347,I131950,I131968,I132392,I381854,I132409,I131971,I131956,I131965,I131974,I132512,I551106,I132538,I132546,I551085,I132563,I551112,I132589,I132480,I132611,I551100,I132637,I132645,I551103,I132662,I132688,I132504,I132710,I132486,I551094,I132750,I132767,I132775,I132792,I132489,I132823,I551091,I551088,I132840,I551109,I132866,I132874,I132477,I132495,I132919,I551097,I132936,I132498,I132483,I132492,I132501,I133039,I452196,I133065,I133073,I452211,I133090,I452214,I133116,I133007,I133138,I452220,I133164,I133172,I452202,I133189,I133215,I133031,I133237,I133013,I452199,I133277,I133294,I133302,I133319,I133016,I133350,I452205,I133367,I452217,I133393,I133401,I133004,I133022,I133446,I452208,I133463,I133025,I133010,I133019,I133028,I133566,I133592,I133600,I133617,I133643,I133534,I133665,I133691,I133699,I133716,I133742,I133558,I133764,I133540,I133804,I133821,I133829,I133846,I133543,I133877,I133894,I133920,I133928,I133531,I133549,I133973,I133990,I133552,I133537,I133546,I133555,I134093,I214403,I134119,I134127,I214415,I134144,I214400,I134170,I134192,I214424,I134218,I134226,I214421,I134243,I134269,I134291,I214412,I134331,I134348,I134356,I134373,I134404,I214409,I134421,I214418,I134447,I134455,I134500,I214406,I134517,I134620,I190884,I134646,I134654,I190896,I190875,I134671,I190899,I134697,I134588,I134719,I190890,I134745,I134753,I190872,I134770,I134796,I134612,I134818,I134594,I190887,I134858,I134875,I134883,I134900,I134597,I134931,I190878,I134948,I190881,I134974,I134982,I134585,I134603,I135027,I190893,I135044,I134606,I134591,I134600,I134609,I135147,I462022,I135173,I135181,I462037,I135198,I462040,I135224,I135246,I462046,I135272,I135280,I462028,I135297,I135323,I135345,I462025,I135385,I135402,I135410,I135427,I135458,I462031,I135475,I462043,I135501,I135509,I135554,I462034,I135571,I135674,I135700,I135708,I135725,I135751,I135642,I135773,I135799,I135807,I135824,I135850,I135666,I135872,I135648,I135912,I135929,I135937,I135954,I135651,I135985,I136002,I136028,I136036,I135639,I135657,I136081,I136098,I135660,I135645,I135654,I135663,I136201,I376668,I136227,I136235,I376665,I376683,I136252,I376674,I136278,I136169,I136300,I376689,I136326,I136334,I376671,I136351,I136377,I136193,I136399,I136175,I376677,I136439,I136456,I136464,I136481,I136178,I136512,I376692,I136529,I376680,I136555,I136563,I136166,I136184,I136608,I376686,I136625,I136187,I136172,I136181,I136190,I136728,I241207,I136754,I136762,I241192,I241195,I136779,I241210,I136805,I136696,I136827,I241204,I136853,I136861,I136878,I136904,I136720,I136926,I136702,I241201,I136966,I136983,I136991,I137008,I136705,I137039,I241216,I137056,I241213,I137082,I137090,I136693,I136711,I137135,I241198,I137152,I136714,I136699,I136708,I136717,I137255,I137281,I137289,I137306,I137332,I137223,I137354,I137380,I137388,I137405,I137431,I137247,I137453,I137229,I137493,I137510,I137518,I137535,I137232,I137566,I137583,I137609,I137617,I137220,I137238,I137662,I137679,I137241,I137226,I137235,I137244,I137782,I137808,I137816,I137833,I137859,I137750,I137881,I137907,I137915,I137932,I137958,I137774,I137980,I137756,I138020,I138037,I138045,I138062,I137759,I138093,I138110,I138136,I138144,I137747,I137765,I138189,I138206,I137768,I137753,I137762,I137771,I138309,I249877,I138335,I138343,I249862,I249865,I138360,I249880,I138386,I138277,I138408,I249874,I138434,I138442,I138459,I138485,I138301,I138507,I138283,I249871,I138547,I138564,I138572,I138589,I138286,I138620,I249886,I138637,I249883,I138663,I138671,I138274,I138292,I138716,I249868,I138733,I138295,I138280,I138289,I138298,I138836,I138862,I138870,I138887,I138913,I138804,I138935,I138961,I138969,I138986,I139012,I138828,I139034,I138810,I139074,I139091,I139099,I139116,I138813,I139147,I139164,I139190,I139198,I138801,I138819,I139243,I139260,I138822,I138807,I138816,I138825,I139363,I256813,I139389,I139397,I256798,I256801,I139414,I256816,I139440,I139331,I139462,I256810,I139488,I139496,I139513,I139539,I139355,I139561,I139337,I256807,I139601,I139618,I139626,I139643,I139340,I139674,I256822,I139691,I256819,I139717,I139725,I139328,I139346,I139770,I256804,I139787,I139349,I139334,I139343,I139352,I139890,I494968,I139916,I139924,I494983,I139941,I494986,I139967,I139989,I494992,I140015,I140023,I494974,I140040,I140066,I140088,I494971,I140128,I140145,I140153,I140170,I140201,I494977,I140218,I494989,I140244,I140252,I140297,I494980,I140314,I140417,I260856,I140443,I140451,I260847,I260862,I140468,I260868,I140494,I140385,I140516,I260853,I140542,I140550,I140567,I140593,I140409,I140615,I140391,I260850,I140655,I140672,I140680,I140697,I140394,I140728,I260844,I260859,I140745,I140771,I140779,I140382,I140400,I140824,I260865,I140841,I140403,I140388,I140397,I140406,I140944,I432734,I140970,I140978,I432731,I140995,I432743,I141021,I140912,I141043,I141069,I141077,I432749,I141094,I141120,I140936,I141142,I140918,I432737,I141182,I141199,I141207,I141224,I140921,I141255,I432746,I432752,I141272,I141298,I141306,I140909,I140927,I141351,I432740,I141368,I140930,I140915,I140924,I140933,I141471,I363748,I141497,I141505,I363745,I363763,I141522,I363754,I141548,I141439,I141570,I363769,I141596,I141604,I363751,I141621,I141647,I141463,I141669,I141445,I363757,I141709,I141726,I141734,I141751,I141448,I141782,I363772,I141799,I363760,I141825,I141833,I141436,I141454,I141878,I363766,I141895,I141457,I141442,I141451,I141460,I141998,I142024,I142032,I142049,I142075,I141966,I142097,I142123,I142131,I142148,I142174,I141990,I142196,I141972,I142236,I142253,I142261,I142278,I141975,I142309,I142326,I142352,I142360,I141963,I141981,I142405,I142422,I141984,I141969,I141978,I141987,I142525,I142551,I142559,I142576,I142602,I142624,I142650,I142658,I142675,I142701,I142723,I142763,I142780,I142788,I142805,I142836,I142853,I142879,I142887,I142932,I142949,I143052,I379252,I143078,I143086,I379249,I379267,I143103,I379258,I143129,I143151,I379273,I143177,I143185,I379255,I143202,I143228,I143250,I379261,I143290,I143307,I143315,I143332,I143363,I379276,I143380,I379264,I143406,I143414,I143459,I379270,I143476,I143579,I509572,I143605,I143613,I509554,I509578,I143630,I509569,I143656,I143547,I143678,I509575,I143704,I143712,I509563,I143729,I143755,I143571,I143777,I143553,I143817,I143834,I143842,I143859,I143556,I143890,I509560,I509557,I143907,I509566,I143933,I143941,I143544,I143562,I143986,I144003,I143565,I143550,I143559,I143568,I144106,I312298,I144132,I144140,I312289,I312304,I144157,I312310,I144183,I144074,I144205,I312295,I144231,I144239,I144256,I144282,I144098,I144304,I144080,I312292,I144344,I144361,I144369,I144386,I144083,I144417,I312286,I312301,I144434,I144460,I144468,I144071,I144089,I144513,I312307,I144530,I144092,I144077,I144086,I144095,I144633,I332825,I144659,I144667,I332828,I332822,I144684,I332834,I144710,I144601,I144732,I332837,I144758,I144766,I144783,I144809,I144625,I144831,I144607,I332840,I144871,I144888,I144896,I144913,I144610,I144944,I332831,I144961,I144987,I144995,I144598,I144616,I145040,I332843,I145057,I144619,I144604,I144613,I144622,I145160,I209048,I145186,I145194,I209060,I145211,I209045,I145237,I145128,I145259,I209069,I145285,I145293,I209066,I145310,I145336,I145152,I145358,I145134,I209057,I145398,I145415,I145423,I145440,I145137,I145471,I209054,I145488,I209063,I145514,I145522,I145125,I145143,I145567,I209051,I145584,I145146,I145131,I145140,I145149,I145687,I308830,I145713,I145721,I308821,I308836,I145738,I308842,I145764,I145786,I308827,I145812,I145820,I145837,I145863,I145885,I308824,I145925,I145942,I145950,I145967,I145998,I308818,I308833,I146015,I146041,I146049,I146094,I308839,I146111,I146214,I146240,I146248,I146265,I146291,I146182,I146313,I146339,I146347,I146364,I146390,I146206,I146412,I146188,I146452,I146469,I146477,I146494,I146191,I146525,I146542,I146568,I146576,I146179,I146197,I146621,I146638,I146200,I146185,I146194,I146203,I146741,I556461,I146767,I146775,I556440,I146792,I556467,I146818,I146840,I556455,I146866,I146874,I556458,I146891,I146917,I146939,I556449,I146979,I146996,I147004,I147021,I147052,I556446,I556443,I147069,I556464,I147095,I147103,I147148,I556452,I147165,I147268,I254501,I147294,I147302,I254486,I254489,I147319,I254504,I147345,I147236,I147367,I254498,I147393,I147401,I147418,I147444,I147260,I147466,I147242,I254495,I147506,I147523,I147531,I147548,I147245,I147579,I254510,I147596,I254507,I147622,I147630,I147233,I147251,I147675,I254492,I147692,I147254,I147239,I147248,I147257,I147795,I270682,I147821,I147829,I270673,I270688,I147846,I270694,I147872,I147763,I147894,I270679,I147920,I147928,I147945,I147971,I147787,I147993,I147769,I270676,I148033,I148050,I148058,I148075,I147772,I148106,I270670,I270685,I148123,I148149,I148157,I147760,I147778,I148202,I270691,I148219,I147781,I147766,I147775,I147784,I148322,I148348,I148356,I148373,I148399,I148290,I148421,I148447,I148455,I148472,I148498,I148314,I148520,I148296,I148560,I148577,I148585,I148602,I148299,I148633,I148650,I148676,I148684,I148287,I148305,I148729,I148746,I148308,I148293,I148302,I148311,I148849,I148875,I148883,I148900,I148926,I148817,I148948,I148974,I148982,I148999,I149025,I148841,I149047,I148823,I149087,I149104,I149112,I149129,I148826,I149160,I149177,I149203,I149211,I148814,I148832,I149256,I149273,I148835,I148820,I148829,I148838,I149376,I324920,I149402,I149410,I324923,I324917,I149427,I324929,I149453,I149344,I149475,I324932,I149501,I149509,I149526,I149552,I149368,I149574,I149350,I324935,I149614,I149631,I149639,I149656,I149353,I149687,I324926,I149704,I149730,I149738,I149341,I149359,I149783,I324938,I149800,I149362,I149347,I149356,I149365,I149903,I374084,I149929,I149937,I374081,I374099,I149954,I374090,I149980,I149871,I150002,I374105,I150028,I150036,I374087,I150053,I150079,I149895,I150101,I149877,I374093,I150141,I150158,I150166,I150183,I149880,I150214,I374108,I150231,I374096,I150257,I150265,I149868,I149886,I150310,I374102,I150327,I149889,I149874,I149883,I149892,I150430,I353905,I150456,I150464,I353908,I353902,I150481,I353914,I150507,I150529,I353917,I150555,I150563,I150580,I150606,I150628,I353920,I150668,I150685,I150693,I150710,I150741,I353911,I150758,I150784,I150792,I150837,I353923,I150854,I150957,I478784,I150983,I150991,I478799,I151008,I478802,I151034,I150925,I151056,I478808,I151082,I151090,I478790,I151107,I151133,I150949,I151155,I150931,I478787,I151195,I151212,I151220,I151237,I150934,I151268,I478793,I151285,I478805,I151311,I151319,I150922,I150940,I151364,I478796,I151381,I150943,I150928,I150937,I150946,I151484,I264324,I151510,I151518,I264315,I264330,I151535,I264336,I151561,I151452,I151583,I264321,I151609,I151617,I151634,I151660,I151476,I151682,I151458,I264318,I151722,I151739,I151747,I151764,I151461,I151795,I264312,I264327,I151812,I151838,I151846,I151449,I151467,I151891,I264333,I151908,I151470,I151455,I151464,I151473,I152011,I169668,I152037,I152045,I169680,I169659,I152062,I169683,I152088,I151979,I152110,I169674,I152136,I152144,I169656,I152161,I152187,I152003,I152209,I151985,I169671,I152249,I152266,I152274,I152291,I151988,I152322,I169662,I152339,I169665,I152365,I152373,I151976,I151994,I152418,I169677,I152435,I151997,I151982,I151991,I152000,I152538,I229069,I152564,I152572,I229054,I229057,I152589,I229072,I152615,I152506,I152637,I229066,I152663,I152671,I152688,I152714,I152530,I152736,I152512,I229063,I152776,I152793,I152801,I152818,I152515,I152849,I229078,I152866,I229075,I152892,I152900,I152503,I152521,I152945,I229060,I152962,I152524,I152509,I152518,I152527,I153065,I153091,I153099,I153116,I153142,I153164,I153190,I153198,I153215,I153241,I153263,I153303,I153320,I153328,I153345,I153376,I153393,I153419,I153427,I153472,I153489,I153592,I465490,I153618,I153626,I465505,I153643,I465508,I153669,I153560,I153691,I465514,I153717,I153725,I465496,I153742,I153768,I153584,I153790,I153566,I465493,I153830,I153847,I153855,I153872,I153569,I153903,I465499,I153920,I465511,I153946,I153954,I153557,I153575,I153999,I465502,I154016,I153578,I153563,I153572,I153581,I154119,I449306,I154145,I154153,I449321,I154170,I449324,I154196,I154087,I154218,I449330,I154244,I154252,I449312,I154269,I154295,I154111,I154317,I154093,I449309,I154357,I154374,I154382,I154399,I154096,I154430,I449315,I154447,I449327,I154473,I154481,I154084,I154102,I154526,I449318,I154543,I154105,I154090,I154099,I154108,I154646,I338095,I154672,I154680,I338098,I338092,I154697,I338104,I154723,I154614,I154745,I338107,I154771,I154779,I154796,I154822,I154638,I154844,I154620,I338110,I154884,I154901,I154909,I154926,I154623,I154957,I338101,I154974,I155000,I155008,I154611,I154629,I155053,I338113,I155070,I154632,I154617,I154626,I154635,I155173,I155199,I155207,I155224,I155250,I155272,I155298,I155306,I155323,I155349,I155371,I155411,I155428,I155436,I155453,I155484,I155501,I155527,I155535,I155580,I155597,I155700,I467224,I155726,I155734,I467239,I155751,I467242,I155777,I155799,I467248,I155825,I155833,I467230,I155850,I155876,I155898,I467227,I155938,I155955,I155963,I155980,I156011,I467233,I156028,I467245,I156054,I156062,I156107,I467236,I156124,I156227,I441792,I156253,I156261,I441807,I156278,I441810,I156304,I156195,I156326,I441816,I156352,I156360,I441798,I156377,I156403,I156219,I156425,I156201,I441795,I156465,I156482,I156490,I156507,I156204,I156538,I441801,I156555,I441813,I156581,I156589,I156192,I156210,I156634,I441804,I156651,I156213,I156198,I156207,I156216,I156754,I156780,I156788,I156805,I156831,I156722,I156853,I156879,I156887,I156904,I156930,I156746,I156952,I156728,I156992,I157009,I157017,I157034,I156731,I157065,I157082,I157108,I157116,I156719,I156737,I157161,I157178,I156740,I156725,I156734,I156743,I157281,I310564,I157307,I157315,I310555,I310570,I157332,I310576,I157358,I157249,I157380,I310561,I157406,I157414,I157431,I157457,I157273,I157479,I157255,I310558,I157519,I157536,I157544,I157561,I157258,I157592,I310552,I310567,I157609,I157635,I157643,I157246,I157264,I157688,I310573,I157705,I157267,I157252,I157261,I157270,I157808,I458554,I157834,I157842,I458569,I157859,I458572,I157885,I157776,I157907,I458578,I157933,I157941,I458560,I157958,I157984,I157800,I158006,I157782,I458557,I158046,I158063,I158071,I158088,I157785,I158119,I458563,I158136,I458575,I158162,I158170,I157773,I157791,I158215,I458566,I158232,I157794,I157779,I157788,I157797,I158335,I257388,I158361,I158369,I257379,I257394,I158386,I257400,I158412,I158303,I158434,I257385,I158460,I158468,I158485,I158511,I158327,I158533,I158309,I257382,I158573,I158590,I158598,I158615,I158312,I158646,I257376,I257391,I158663,I158689,I158697,I158300,I158318,I158742,I257397,I158759,I158321,I158306,I158315,I158324,I158862,I434978,I158888,I158896,I434975,I158913,I434987,I158939,I158830,I158961,I158987,I158995,I434993,I159012,I159038,I158854,I159060,I158836,I434981,I159100,I159117,I159125,I159142,I158839,I159173,I434990,I434996,I159190,I159216,I159224,I158827,I158845,I159269,I434984,I159286,I158848,I158833,I158842,I158851,I159389,I253345,I159415,I159423,I253330,I253333,I159440,I253348,I159466,I159357,I159488,I253342,I159514,I159522,I159539,I159565,I159381,I159587,I159363,I253339,I159627,I159644,I159652,I159669,I159366,I159700,I253354,I159717,I253351,I159743,I159751,I159354,I159372,I159796,I253336,I159813,I159375,I159360,I159369,I159378,I159916,I160964,I159942,I159950,I160976,I160955,I159967,I160979,I159993,I159884,I160015,I160970,I160041,I160049,I160952,I160066,I160092,I159908,I160114,I159890,I160967,I160154,I160171,I160179,I160196,I159893,I160227,I160958,I160244,I160961,I160270,I160278,I159881,I159899,I160323,I160973,I160340,I159902,I159887,I159896,I159905,I160443,I501907,I160469,I160486,I160508,I160525,I501919,I160542,I501910,I160568,I160576,I501928,I160602,I160610,I501904,I160627,I501922,I160667,I160675,I160720,I501916,I501913,I160737,I501925,I160763,I160785,I160802,I160819,I160850,I160867,I160898,I160987,I501329,I161013,I161030,I161052,I161069,I501341,I161086,I501332,I161112,I161120,I501350,I161146,I161154,I501326,I161171,I501344,I161211,I161219,I161264,I501338,I501335,I161281,I501347,I161307,I161329,I161346,I161363,I161394,I161411,I161442,I161531,I294371,I161557,I161574,I161596,I161613,I294392,I294383,I161630,I161656,I161664,I294377,I161690,I161698,I294374,I161715,I294368,I161755,I161763,I161808,I294380,I161825,I294389,I161851,I161873,I161890,I161907,I161938,I161955,I294386,I161986,I162075,I162101,I162118,I162067,I162140,I162157,I162174,I162200,I162208,I162234,I162242,I162259,I162046,I162299,I162307,I162040,I162055,I162352,I162369,I162395,I162043,I162417,I162434,I162451,I162058,I162482,I162499,I162049,I162530,I162052,I162064,I162061,I162619,I162645,I162662,I162684,I162701,I162718,I162744,I162752,I162778,I162786,I162803,I162843,I162851,I162896,I162913,I162939,I162961,I162978,I162995,I163026,I163043,I163074,I163163,I232525,I163189,I163206,I163155,I163228,I163245,I232522,I232543,I163262,I232546,I163288,I163296,I232531,I163322,I163330,I232534,I163347,I163134,I232537,I163387,I163395,I163128,I163143,I163440,I232528,I163457,I232540,I163483,I163131,I163505,I163522,I163539,I163146,I163570,I163587,I163137,I163618,I163140,I163152,I163149,I163707,I163733,I163750,I163772,I163789,I163806,I163832,I163840,I163866,I163874,I163891,I163931,I163939,I163984,I164001,I164027,I164049,I164066,I164083,I164114,I164131,I164162,I164251,I368273,I164277,I164294,I164243,I164316,I164333,I368288,I368276,I164350,I368267,I164376,I164384,I368279,I164410,I164418,I368270,I164435,I164222,I368285,I164475,I164483,I164216,I164231,I164528,I368294,I368282,I164545,I368291,I164571,I164219,I164593,I164610,I164627,I164234,I164658,I164675,I164225,I164706,I164228,I164240,I164237,I164795,I164821,I164838,I164787,I164860,I164877,I164894,I164920,I164928,I164954,I164962,I164979,I164766,I165019,I165027,I164760,I164775,I165072,I165089,I165115,I164763,I165137,I165154,I165171,I164778,I165202,I165219,I164769,I165250,I164772,I164784,I164781,I165339,I352860,I165365,I165382,I165331,I165404,I165421,I352854,I352851,I165438,I352866,I165464,I165472,I165498,I165506,I352848,I165523,I165310,I165563,I165571,I165304,I165319,I165616,I352863,I352857,I165633,I165659,I165307,I165681,I165698,I165715,I165322,I165746,I165763,I352869,I165313,I165794,I165316,I165328,I165325,I165883,I425438,I165909,I165926,I165875,I165948,I165965,I425456,I165982,I425450,I166008,I166016,I425444,I166042,I166050,I425453,I166067,I165854,I425441,I166107,I166115,I165848,I165863,I166160,I425459,I166177,I166203,I165851,I166225,I166242,I166259,I165866,I166290,I166307,I425447,I165857,I166338,I165860,I165872,I165869,I166427,I368919,I166453,I166470,I166492,I166509,I368934,I368922,I166526,I368913,I166552,I166560,I368925,I166586,I166594,I368916,I166611,I368931,I166651,I166659,I166704,I368940,I368928,I166721,I368937,I166747,I166769,I166786,I166803,I166834,I166851,I166882,I166971,I166997,I167014,I166963,I167036,I167053,I167070,I167096,I167104,I167130,I167138,I167155,I166942,I167195,I167203,I166936,I166951,I167248,I167265,I167291,I166939,I167313,I167330,I167347,I166954,I167378,I167395,I166945,I167426,I166948,I166960,I166957,I167515,I351806,I167541,I167558,I167580,I167597,I351800,I351797,I167614,I351812,I167640,I167648,I167674,I167682,I351794,I167699,I167739,I167747,I167792,I351809,I351803,I167809,I167835,I167857,I167874,I167891,I167922,I167939,I351815,I167970,I168059,I298995,I168085,I168102,I168124,I168141,I299016,I299007,I168158,I168184,I168192,I299001,I168218,I168226,I298998,I168243,I298992,I168283,I168291,I168336,I299004,I168353,I299013,I168379,I168401,I168418,I168435,I168466,I168483,I299010,I168514,I168603,I444685,I168629,I168646,I168668,I168685,I444697,I168702,I444688,I168728,I168736,I444706,I168762,I168770,I444682,I168787,I444700,I168827,I168835,I168880,I444694,I444691,I168897,I444703,I168923,I168945,I168962,I168979,I169010,I169027,I169058,I169147,I511733,I169173,I169190,I169139,I169212,I169229,I511745,I511748,I169246,I511751,I169272,I169280,I511736,I169306,I169314,I511742,I169331,I169118,I511730,I169371,I169379,I169112,I169127,I169424,I511754,I169441,I511739,I169467,I169115,I169489,I169506,I169523,I169130,I169554,I169571,I169121,I169602,I169124,I169136,I169133,I169691,I481677,I169717,I169734,I169756,I169773,I481689,I169790,I481680,I169816,I169824,I481698,I169850,I169858,I481674,I169875,I481692,I169915,I169923,I169968,I481686,I481683,I169985,I481695,I170011,I170033,I170050,I170067,I170098,I170115,I170146,I170235,I539807,I170261,I170278,I170300,I170317,I539783,I539804,I170334,I539801,I170360,I170368,I539780,I170394,I170402,I539792,I170419,I539795,I170459,I170467,I170512,I539798,I539786,I170529,I539789,I170555,I170577,I170594,I170611,I170642,I170659,I170690,I170779,I412201,I170805,I170822,I170771,I170844,I170861,I412216,I412204,I170878,I412195,I170904,I170912,I412207,I170938,I170946,I412198,I170963,I170750,I412213,I171003,I171011,I170744,I170759,I171056,I412222,I412210,I171073,I412219,I171099,I170747,I171121,I171138,I171155,I170762,I171186,I171203,I170753,I171234,I170756,I170768,I170765,I171323,I406387,I171349,I171366,I171388,I171405,I406402,I406390,I171422,I406381,I171448,I171456,I406393,I171482,I171490,I406384,I171507,I406399,I171547,I171555,I171600,I406408,I406396,I171617,I406405,I171643,I171665,I171682,I171699,I171730,I171747,I171778,I171867,I414779,I171893,I171910,I171859,I171932,I171949,I414797,I171966,I414791,I171992,I172000,I414785,I172026,I172034,I414794,I172051,I171838,I414782,I172091,I172099,I171832,I171847,I172144,I414800,I172161,I172187,I171835,I172209,I172226,I172243,I171850,I172274,I172291,I414788,I171841,I172322,I171844,I171856,I171853,I172411,I172437,I172454,I172403,I172476,I172493,I172510,I172536,I172544,I172570,I172578,I172595,I172382,I172635,I172643,I172376,I172391,I172688,I172705,I172731,I172379,I172753,I172770,I172787,I172394,I172818,I172835,I172385,I172866,I172388,I172400,I172397,I172955,I382485,I172981,I172998,I172947,I173020,I173037,I382500,I382488,I173054,I382479,I173080,I173088,I382491,I173114,I173122,I382482,I173139,I172926,I382497,I173179,I173187,I172920,I172935,I173232,I382506,I382494,I173249,I382503,I173275,I172923,I173297,I173314,I173331,I172938,I173362,I173379,I172929,I173410,I172932,I172944,I172941,I173499,I173525,I173542,I173564,I173581,I173598,I173624,I173632,I173658,I173666,I173683,I173723,I173731,I173776,I173793,I173819,I173841,I173858,I173875,I173906,I173923,I173954,I174043,I348644,I174069,I174086,I174108,I174125,I348638,I348635,I174142,I348650,I174168,I174176,I174202,I174210,I348632,I174227,I174267,I174275,I174320,I348647,I348641,I174337,I174363,I174385,I174402,I174419,I174450,I174467,I348653,I174498,I174587,I500751,I174613,I174630,I174579,I174652,I174669,I500763,I174686,I500754,I174712,I174720,I500772,I174746,I174754,I500748,I174771,I174558,I500766,I174811,I174819,I174552,I174567,I174864,I500760,I500757,I174881,I500769,I174907,I174555,I174929,I174946,I174963,I174570,I174994,I175011,I174561,I175042,I174564,I174576,I174573,I175131,I175157,I175174,I175123,I175196,I175213,I175230,I175256,I175264,I175290,I175298,I175315,I175102,I175355,I175363,I175096,I175111,I175408,I175425,I175451,I175099,I175473,I175490,I175507,I175114,I175538,I175555,I175105,I175586,I175108,I175120,I175117,I175675,I446997,I175701,I175718,I175667,I175740,I175757,I447009,I175774,I447000,I175800,I175808,I447018,I175834,I175842,I446994,I175859,I175646,I447012,I175899,I175907,I175640,I175655,I175952,I447006,I447003,I175969,I447015,I175995,I175643,I176017,I176034,I176051,I175658,I176082,I176099,I175649,I176130,I175652,I175664,I175661,I176219,I545162,I176245,I176262,I176211,I176284,I176301,I545138,I545159,I176318,I545156,I176344,I176352,I545135,I176378,I176386,I545147,I176403,I176190,I545150,I176443,I176451,I176184,I176199,I176496,I545153,I545141,I176513,I545144,I176539,I176187,I176561,I176578,I176595,I176202,I176626,I176643,I176193,I176674,I176196,I176208,I176205,I176763,I176789,I176806,I176828,I176845,I176862,I176888,I176896,I176922,I176930,I176947,I176987,I176995,I177040,I177057,I177083,I177105,I177122,I177139,I177170,I177187,I177218,I177307,I177333,I177350,I177372,I177389,I177406,I177432,I177440,I177466,I177474,I177491,I177531,I177539,I177584,I177601,I177627,I177649,I177666,I177683,I177714,I177731,I177762,I177851,I296683,I177877,I177894,I177843,I177916,I177933,I296704,I296695,I177950,I177976,I177984,I296689,I178010,I178018,I296686,I178035,I177822,I296680,I178075,I178083,I177816,I177831,I178128,I296692,I178145,I296701,I178171,I177819,I178193,I178210,I178227,I177834,I178258,I178275,I296698,I177825,I178306,I177828,I177840,I177837,I178395,I178421,I178438,I178387,I178460,I178477,I178494,I178520,I178528,I178554,I178562,I178579,I178366,I178619,I178627,I178360,I178375,I178672,I178689,I178715,I178363,I178737,I178754,I178771,I178378,I178802,I178819,I178369,I178850,I178372,I178384,I178381,I178939,I290325,I178965,I178982,I178931,I179004,I179021,I290346,I290337,I179038,I179064,I179072,I290331,I179098,I179106,I290328,I179123,I178910,I290322,I179163,I179171,I178904,I178919,I179216,I290334,I179233,I290343,I179259,I178907,I179281,I179298,I179315,I178922,I179346,I179363,I290340,I178913,I179394,I178916,I178928,I178925,I179483,I179509,I179526,I179475,I179548,I179565,I179582,I179608,I179616,I179642,I179650,I179667,I179454,I179707,I179715,I179448,I179463,I179760,I179777,I179803,I179451,I179825,I179842,I179859,I179466,I179890,I179907,I179457,I179938,I179460,I179472,I179469,I180027,I542782,I180053,I180070,I180019,I180092,I180109,I542758,I542779,I180126,I542776,I180152,I180160,I542755,I180186,I180194,I542767,I180211,I179998,I542770,I180251,I180259,I179992,I180007,I180304,I542773,I542761,I180321,I542764,I180347,I179995,I180369,I180386,I180403,I180010,I180434,I180451,I180001,I180482,I180004,I180016,I180013,I180571,I360238,I180597,I180614,I180636,I180653,I360232,I360229,I180670,I360244,I180696,I180704,I180730,I180738,I360226,I180755,I180795,I180803,I180848,I360241,I360235,I180865,I180891,I180913,I180930,I180947,I180978,I180995,I360247,I181026,I181115,I181141,I181158,I181180,I181197,I181214,I181240,I181248,I181274,I181282,I181299,I181339,I181347,I181392,I181409,I181435,I181457,I181474,I181491,I181522,I181539,I181570,I181659,I446419,I181685,I181702,I181651,I181724,I181741,I446431,I181758,I446422,I181784,I181792,I446440,I181818,I181826,I446416,I181843,I181630,I446434,I181883,I181891,I181624,I181639,I181936,I446428,I446425,I181953,I446437,I181979,I181627,I182001,I182018,I182035,I181642,I182066,I182083,I181633,I182114,I181636,I181648,I181645,I182203,I364397,I182229,I182246,I182268,I182285,I364412,I364400,I182302,I364391,I182328,I182336,I364403,I182362,I182370,I364394,I182387,I364409,I182427,I182435,I182480,I364418,I364406,I182497,I364415,I182523,I182545,I182562,I182579,I182610,I182627,I182658,I182747,I497861,I182773,I182790,I182739,I182812,I182829,I497873,I182846,I497864,I182872,I182880,I497882,I182906,I182914,I497858,I182931,I182718,I497876,I182971,I182979,I182712,I182727,I183024,I497870,I497867,I183041,I497879,I183067,I182715,I183089,I183106,I183123,I182730,I183154,I183171,I182721,I183202,I182724,I182736,I182733,I183291,I492081,I183317,I183334,I183283,I183356,I183373,I492093,I183390,I492084,I183416,I183424,I492102,I183450,I183458,I492078,I183475,I183262,I492096,I183515,I183523,I183256,I183271,I183568,I492090,I492087,I183585,I492099,I183611,I183259,I183633,I183650,I183667,I183274,I183698,I183715,I183265,I183746,I183268,I183280,I183277,I183835,I488035,I183861,I183878,I183827,I183900,I183917,I488047,I183934,I488038,I183960,I183968,I488056,I183994,I184002,I488032,I184019,I183806,I488050,I184059,I184067,I183800,I183815,I184112,I488044,I488041,I184129,I488053,I184155,I183803,I184177,I184194,I184211,I183818,I184242,I184259,I183809,I184290,I183812,I183824,I183821,I184379,I569557,I184405,I184422,I184371,I184444,I184461,I569533,I569554,I184478,I569551,I184504,I184512,I569530,I184538,I184546,I569542,I184563,I184350,I569545,I184603,I184611,I184344,I184359,I184656,I569548,I569536,I184673,I569539,I184699,I184347,I184721,I184738,I184755,I184362,I184786,I184803,I184353,I184834,I184356,I184368,I184365,I184923,I184949,I184966,I184988,I185005,I185022,I185048,I185056,I185082,I185090,I185107,I185147,I185155,I185200,I185217,I185243,I185265,I185282,I185299,I185330,I185347,I185378,I185467,I248131,I185493,I185510,I185459,I185532,I185549,I248128,I248149,I185566,I248152,I185592,I185600,I248137,I185626,I185634,I248140,I185651,I185438,I248143,I185691,I185699,I185432,I185447,I185744,I248134,I185761,I248146,I185787,I185435,I185809,I185826,I185843,I185450,I185874,I185891,I185441,I185922,I185444,I185456,I185453,I186011,I186037,I186054,I186003,I186076,I186093,I186110,I186136,I186144,I186170,I186178,I186195,I185982,I186235,I186243,I185976,I185991,I186288,I186305,I186331,I185979,I186353,I186370,I186387,I185994,I186418,I186435,I185985,I186466,I185988,I186000,I185997,I186555,I186581,I186598,I186547,I186620,I186637,I186654,I186680,I186688,I186714,I186722,I186739,I186526,I186779,I186787,I186520,I186535,I186832,I186849,I186875,I186523,I186897,I186914,I186931,I186538,I186962,I186979,I186529,I187010,I186532,I186544,I186541,I187099,I238883,I187125,I187142,I187164,I187181,I238880,I238901,I187198,I238904,I187224,I187232,I238889,I187258,I187266,I238892,I187283,I238895,I187323,I187331,I187376,I238886,I187393,I238898,I187419,I187441,I187458,I187475,I187506,I187523,I187554,I187643,I507381,I187669,I187686,I187635,I187708,I187725,I507393,I507396,I187742,I507399,I187768,I187776,I507384,I187802,I187810,I507390,I187827,I187614,I507378,I187867,I187875,I187608,I187623,I187920,I507402,I187937,I507387,I187963,I187611,I187985,I188002,I188019,I187626,I188050,I188067,I187617,I188098,I187620,I187632,I187629,I188187,I413493,I188213,I188230,I188252,I188269,I413508,I413496,I188286,I413487,I188312,I188320,I413499,I188346,I188354,I413490,I188371,I413505,I188411,I188419,I188464,I413514,I413502,I188481,I413511,I188507,I188529,I188546,I188563,I188594,I188611,I188642,I188731,I390883,I188757,I188774,I188796,I188813,I390898,I390886,I188830,I390877,I188856,I188864,I390889,I188890,I188898,I390880,I188915,I390895,I188955,I188963,I189008,I390904,I390892,I189025,I390901,I189051,I189073,I189090,I189107,I189138,I189155,I189186,I189275,I189301,I189318,I189267,I189340,I189357,I189374,I189400,I189408,I189434,I189442,I189459,I189246,I189499,I189507,I189240,I189255,I189552,I189569,I189595,I189243,I189617,I189634,I189651,I189258,I189682,I189699,I189249,I189730,I189252,I189264,I189261,I189819,I528170,I189845,I189862,I189811,I189884,I189901,I528167,I528164,I189918,I528152,I189944,I189952,I528176,I189978,I189986,I528161,I190003,I189790,I528155,I190043,I190051,I189784,I189799,I190096,I528158,I190113,I528173,I190139,I189787,I190161,I190178,I190195,I189802,I190226,I190243,I189793,I190274,I189796,I189808,I189805,I190363,I312867,I190389,I190406,I190355,I190428,I190445,I312888,I312879,I190462,I190488,I190496,I312873,I190522,I190530,I312870,I190547,I190334,I312864,I190587,I190595,I190328,I190343,I190640,I312876,I190657,I312885,I190683,I190331,I190705,I190722,I190739,I190346,I190770,I190787,I312882,I190337,I190818,I190340,I190352,I190349,I190907,I571342,I190933,I190950,I190972,I190989,I571318,I571339,I191006,I571336,I191032,I191040,I571315,I191066,I191074,I571327,I191091,I571330,I191131,I191139,I191184,I571333,I571321,I191201,I571324,I191227,I191249,I191266,I191283,I191314,I191331,I191362,I191451,I191477,I191494,I191443,I191516,I191533,I191550,I191576,I191584,I191610,I191618,I191635,I191422,I191675,I191683,I191416,I191431,I191728,I191745,I191771,I191419,I191793,I191810,I191827,I191434,I191858,I191875,I191425,I191906,I191428,I191440,I191437,I191995,I192021,I192038,I191987,I192060,I192077,I192094,I192120,I192128,I192154,I192162,I192179,I191966,I192219,I192227,I191960,I191975,I192272,I192289,I192315,I191963,I192337,I192354,I192371,I191978,I192402,I192419,I191969,I192450,I191972,I191984,I191981,I192539,I479365,I192565,I192582,I192531,I192604,I192621,I479377,I192638,I479368,I192664,I192672,I479386,I192698,I192706,I479362,I192723,I192510,I479380,I192763,I192771,I192504,I192519,I192816,I479374,I479371,I192833,I479383,I192859,I192507,I192881,I192898,I192915,I192522,I192946,I192963,I192513,I192994,I192516,I192528,I192525,I193083,I305353,I193109,I193126,I193075,I193148,I193165,I305374,I305365,I193182,I193208,I193216,I305359,I193242,I193250,I305356,I193267,I193054,I305350,I193307,I193315,I193048,I193063,I193360,I305362,I193377,I305371,I193403,I193051,I193425,I193442,I193459,I193066,I193490,I193507,I305368,I193057,I193538,I193060,I193072,I193069,I193627,I193653,I193670,I193619,I193692,I193709,I193726,I193752,I193760,I193786,I193794,I193811,I193598,I193851,I193859,I193592,I193607,I193904,I193921,I193947,I193595,I193969,I193986,I194003,I193610,I194034,I194051,I193601,I194082,I193604,I193616,I193613,I194171,I194197,I194214,I194163,I194236,I194253,I194270,I194296,I194304,I194330,I194338,I194355,I194142,I194395,I194403,I194136,I194151,I194448,I194465,I194491,I194139,I194513,I194530,I194547,I194154,I194578,I194595,I194145,I194626,I194148,I194160,I194157,I194715,I360765,I194741,I194758,I194707,I194780,I194797,I360759,I360756,I194814,I360771,I194840,I194848,I194874,I194882,I360753,I194899,I194686,I194939,I194947,I194680,I194695,I194992,I360768,I360762,I195009,I195035,I194683,I195057,I195074,I195091,I194698,I195122,I195139,I360774,I194689,I195170,I194692,I194704,I194701,I195259,I348117,I195285,I195302,I195251,I195324,I195341,I348111,I348108,I195358,I348123,I195384,I195392,I195418,I195426,I348105,I195443,I195230,I195483,I195491,I195224,I195239,I195536,I348120,I348114,I195553,I195579,I195227,I195601,I195618,I195635,I195242,I195666,I195683,I348126,I195233,I195714,I195236,I195248,I195245,I195803,I294949,I195829,I195846,I195868,I195885,I294970,I294961,I195902,I195928,I195936,I294955,I195962,I195970,I294952,I195987,I294946,I196027,I196035,I196080,I294958,I196097,I294967,I196123,I196145,I196162,I196179,I196210,I196227,I294964,I196258,I196347,I493815,I196373,I196390,I196339,I196412,I196429,I493827,I196446,I493818,I196472,I196480,I493836,I196506,I196514,I493812,I196531,I196318,I493830,I196571,I196579,I196312,I196327,I196624,I493824,I493821,I196641,I493833,I196667,I196315,I196689,I196706,I196723,I196330,I196754,I196771,I196321,I196802,I196324,I196336,I196333,I196891,I196917,I196934,I196883,I196956,I196973,I196990,I197016,I197024,I197050,I197058,I197075,I196862,I197115,I197123,I196856,I196871,I197168,I197185,I197211,I196859,I197233,I197250,I197267,I196874,I197298,I197315,I196865,I197346,I196868,I196880,I196877,I197435,I237149,I197461,I197478,I197427,I197500,I197517,I237146,I237167,I197534,I237170,I197560,I197568,I237155,I197594,I197602,I237158,I197619,I197406,I237161,I197659,I197667,I197400,I197415,I197712,I237152,I197729,I237164,I197755,I197403,I197777,I197794,I197811,I197418,I197842,I197859,I197409,I197890,I197412,I197424,I197421,I197979,I198005,I198022,I197971,I198044,I198061,I198078,I198104,I198112,I198138,I198146,I198163,I197950,I198203,I198211,I197944,I197959,I198256,I198273,I198299,I197947,I198321,I198338,I198355,I197962,I198386,I198403,I197953,I198434,I197956,I197968,I197965,I198523,I495549,I198549,I198566,I198588,I198605,I495561,I198622,I495552,I198648,I198656,I495570,I198682,I198690,I495546,I198707,I495564,I198747,I198755,I198800,I495558,I495555,I198817,I495567,I198843,I198865,I198882,I198899,I198930,I198947,I198978,I199067,I199093,I199110,I199059,I199132,I199149,I199166,I199192,I199200,I199226,I199234,I199251,I199038,I199291,I199299,I199032,I199047,I199344,I199361,I199387,I199035,I199409,I199426,I199443,I199050,I199474,I199491,I199041,I199522,I199044,I199056,I199053,I199611,I199637,I199654,I199603,I199676,I199693,I199710,I199736,I199744,I199770,I199778,I199795,I199582,I199835,I199843,I199576,I199591,I199888,I199905,I199931,I199579,I199953,I199970,I199987,I199594,I200018,I200035,I199585,I200066,I199588,I199600,I199597,I200152,I200178,I200195,I200144,I200226,I200234,I200251,I200268,I200285,I200302,I200319,I200336,I200141,I200367,I200384,I200401,I200126,I200138,I200446,I200463,I200132,I200494,I200511,I200120,I200542,I200559,I200576,I200602,I200610,I200129,I200641,I200658,I200135,I200689,I200123,I200747,I200773,I200790,I200739,I200821,I200829,I200846,I200863,I200880,I200897,I200914,I200931,I200736,I200962,I200979,I200996,I200721,I200733,I201041,I201058,I200727,I201089,I201106,I200715,I201137,I201154,I201171,I201197,I201205,I200724,I201236,I201253,I200730,I201284,I200718,I201342,I201368,I201385,I201334,I201416,I201424,I201441,I201458,I201475,I201492,I201509,I201526,I201331,I201557,I201574,I201591,I201316,I201328,I201636,I201653,I201322,I201684,I201701,I201310,I201732,I201749,I201766,I201792,I201800,I201319,I201831,I201848,I201325,I201879,I201313,I201937,I201963,I201980,I201929,I202011,I202019,I202036,I202053,I202070,I202087,I202104,I202121,I201926,I202152,I202169,I202186,I201911,I201923,I202231,I202248,I201917,I202279,I202296,I201905,I202327,I202344,I202361,I202387,I202395,I201914,I202426,I202443,I201920,I202474,I201908,I202532,I423194,I202558,I202575,I423197,I202606,I202614,I423200,I202631,I202648,I423212,I202665,I423203,I202682,I202699,I202716,I202747,I423209,I202764,I202781,I202826,I202843,I202874,I202891,I202922,I423206,I202939,I202956,I423215,I202982,I202990,I203021,I203038,I203069,I203127,I454526,I203153,I203170,I203119,I454508,I203201,I203209,I454514,I203226,I203243,I454529,I203260,I454520,I203277,I203294,I203311,I203116,I203342,I454532,I203359,I454511,I203376,I203101,I203113,I203421,I203438,I203107,I203469,I454517,I203486,I203095,I203517,I454523,I203534,I203551,I203577,I203585,I203104,I203616,I203633,I203110,I203664,I203098,I203722,I357600,I203748,I203765,I357597,I203796,I203804,I203821,I203838,I357594,I203855,I357609,I203872,I203889,I203906,I203937,I357603,I203954,I357591,I203971,I204016,I204033,I204064,I357612,I204081,I204112,I204129,I357606,I204146,I204172,I204180,I204211,I204228,I204259,I204317,I525271,I204343,I204360,I204309,I525277,I204391,I204399,I525265,I204416,I204433,I525268,I204450,I525274,I204467,I204484,I204501,I204306,I204532,I204549,I525283,I204566,I204291,I204303,I204611,I204628,I204297,I204659,I525262,I204676,I204285,I204707,I525286,I204724,I204741,I525280,I204767,I204775,I204294,I204806,I204823,I204300,I204854,I204288,I204912,I204938,I204955,I204986,I204994,I205011,I205028,I205045,I205062,I205079,I205096,I205127,I205144,I205161,I205206,I205223,I205254,I205271,I205302,I205319,I205336,I205362,I205370,I205401,I205418,I205449,I205507,I506290,I205533,I205550,I506305,I205581,I205589,I506314,I205606,I205623,I506293,I205640,I506299,I205657,I205674,I205691,I205722,I506311,I205739,I506308,I205756,I205801,I205818,I205849,I205866,I205897,I506302,I205914,I506296,I205931,I205957,I205965,I205996,I206013,I206044,I206102,I206128,I206145,I206176,I206184,I206201,I206218,I206235,I206252,I206269,I206286,I206317,I206334,I206351,I206396,I206413,I206444,I206461,I206492,I206509,I206526,I206552,I206560,I206591,I206608,I206639,I206697,I206723,I206740,I206771,I206779,I206796,I206813,I206830,I206847,I206864,I206881,I206912,I206929,I206946,I206991,I207008,I207039,I207056,I207087,I207104,I207121,I207147,I207155,I207186,I207203,I207234,I207292,I207318,I207335,I207284,I207366,I207374,I207391,I207408,I207425,I207442,I207459,I207476,I207281,I207507,I207524,I207541,I207266,I207278,I207586,I207603,I207272,I207634,I207651,I207260,I207682,I207699,I207716,I207742,I207750,I207269,I207781,I207798,I207275,I207829,I207263,I207887,I207913,I207930,I207961,I207969,I207986,I208003,I208020,I208037,I208054,I208071,I208102,I208119,I208136,I208181,I208198,I208229,I208246,I208277,I208294,I208311,I208337,I208345,I208376,I208393,I208424,I208482,I554655,I208508,I208525,I208474,I554661,I208556,I208564,I554676,I208581,I208598,I554667,I208615,I554664,I208632,I208649,I208666,I208471,I208697,I208714,I554679,I208731,I208456,I208468,I208776,I208793,I208462,I208824,I554673,I208841,I208450,I208872,I554658,I208889,I554670,I208906,I554682,I208932,I208940,I208459,I208971,I208988,I208465,I209019,I208453,I209077,I359181,I209103,I209120,I359178,I209151,I209159,I209176,I209193,I359175,I209210,I359190,I209227,I209244,I209261,I209292,I359184,I209309,I359172,I209326,I209371,I209388,I209419,I359193,I209436,I209467,I209484,I359187,I209501,I209527,I209535,I209566,I209583,I209614,I209672,I242351,I209698,I209715,I209664,I242363,I209746,I209754,I242348,I209771,I209788,I242366,I209805,I242357,I209822,I209839,I209856,I209661,I209887,I242369,I209904,I242372,I209921,I209646,I209658,I209966,I209983,I209652,I210014,I210031,I209640,I210062,I242360,I210079,I242354,I210096,I210122,I210130,I209649,I210161,I210178,I209655,I210209,I209643,I210267,I210293,I210310,I210341,I210349,I210366,I210383,I210400,I210417,I210434,I210451,I210482,I210499,I210516,I210561,I210578,I210609,I210626,I210657,I210674,I210691,I210717,I210725,I210756,I210773,I210804,I210862,I469554,I210888,I210905,I469536,I210936,I210944,I469542,I210961,I210978,I469557,I210995,I469548,I211012,I211029,I211046,I211077,I469560,I211094,I469539,I211111,I211156,I211173,I211204,I469545,I211221,I211252,I469551,I211269,I211286,I211312,I211320,I211351,I211368,I211399,I211457,I479958,I211483,I211500,I479940,I211531,I211539,I479946,I211556,I211573,I479961,I211590,I479952,I211607,I211624,I211641,I211672,I479964,I211689,I479943,I211706,I211751,I211768,I211799,I479949,I211816,I211847,I479955,I211864,I211881,I211907,I211915,I211946,I211963,I211994,I212052,I267789,I212078,I212095,I212044,I267783,I212126,I212134,I267780,I212151,I212168,I267792,I212185,I267795,I212202,I212219,I212236,I212041,I212267,I267804,I212284,I267798,I212301,I212026,I212038,I212346,I212363,I212032,I212394,I267786,I212411,I212020,I212442,I267801,I212459,I212476,I212502,I212510,I212029,I212541,I212558,I212035,I212589,I212023,I212647,I212673,I212690,I212639,I212721,I212729,I212746,I212763,I212780,I212797,I212814,I212831,I212636,I212862,I212879,I212896,I212621,I212633,I212941,I212958,I212627,I212989,I213006,I212615,I213037,I213054,I213071,I213097,I213105,I212624,I213136,I213153,I212630,I213184,I212618,I213242,I351276,I213268,I213285,I351273,I213316,I213324,I213341,I213358,I351270,I213375,I351285,I213392,I213409,I213426,I213457,I351279,I213474,I351267,I213491,I213536,I213553,I213584,I351288,I213601,I213632,I213649,I351282,I213666,I213692,I213700,I213731,I213748,I213779,I213837,I420950,I213863,I213880,I213829,I420953,I213911,I213919,I420956,I213936,I213953,I420968,I213970,I420959,I213987,I214004,I214021,I213826,I214052,I420965,I214069,I214086,I213811,I213823,I214131,I214148,I213817,I214179,I214196,I213805,I214227,I420962,I214244,I214261,I420971,I214287,I214295,I213814,I214326,I214343,I213820,I214374,I213808,I214432,I514994,I214458,I214475,I515009,I214506,I214514,I515018,I214531,I214548,I514997,I214565,I515003,I214582,I214599,I214616,I214647,I515015,I214664,I515012,I214681,I214726,I214743,I214774,I214791,I214822,I515006,I214839,I515000,I214856,I214882,I214890,I214921,I214938,I214969,I215027,I536805,I215053,I215070,I215019,I536811,I215101,I215109,I536826,I215126,I215143,I536817,I215160,I536814,I215177,I215194,I215211,I215016,I215242,I215259,I536829,I215276,I215001,I215013,I215321,I215338,I215007,I215369,I536823,I215386,I214995,I215417,I536808,I215434,I536820,I215451,I536832,I215477,I215485,I215004,I215516,I215533,I215010,I215564,I214998,I215622,I215648,I215665,I215614,I215696,I215704,I215721,I215738,I215755,I215772,I215789,I215806,I215611,I215837,I215854,I215871,I215596,I215608,I215916,I215933,I215602,I215964,I215981,I215590,I216012,I216029,I216046,I216072,I216080,I215599,I216111,I216128,I215605,I216159,I215593,I216217,I468398,I216243,I216260,I468380,I216291,I216299,I468386,I216316,I216333,I468401,I216350,I468392,I216367,I216384,I216401,I216432,I468404,I216449,I468383,I216466,I216511,I216528,I216559,I468389,I216576,I216607,I468395,I216624,I216641,I216667,I216675,I216706,I216723,I216754,I216812,I322818,I216838,I216855,I216804,I322815,I216886,I216894,I216911,I216928,I322812,I216945,I322827,I216962,I216979,I216996,I216801,I217027,I322821,I217044,I322809,I217061,I216786,I216798,I217106,I217123,I216792,I217154,I322830,I217171,I216780,I217202,I217219,I322824,I217236,I217262,I217270,I216789,I217301,I217318,I216795,I217349,I216783,I217407,I217433,I217450,I217481,I217489,I217506,I217523,I217540,I217557,I217574,I217591,I217622,I217639,I217656,I217701,I217718,I217749,I217766,I217797,I217814,I217831,I217857,I217865,I217896,I217913,I217944,I218002,I218028,I218045,I217994,I218076,I218084,I218101,I218118,I218135,I218152,I218169,I218186,I217991,I218217,I218234,I218251,I217976,I217988,I218296,I218313,I217982,I218344,I218361,I217970,I218392,I218409,I218426,I218452,I218460,I217979,I218491,I218508,I217985,I218539,I217973,I218597,I434414,I218623,I218640,I434417,I218671,I218679,I434420,I218696,I218713,I434432,I218730,I434423,I218747,I218764,I218781,I218812,I434429,I218829,I218846,I218891,I218908,I218939,I218956,I218987,I434426,I219004,I219021,I434435,I219047,I219055,I219086,I219103,I219134,I219192,I354438,I219218,I219235,I219184,I354435,I219266,I219274,I219291,I219308,I354432,I219325,I354447,I219342,I219359,I219376,I219181,I219407,I354441,I219424,I354429,I219441,I219166,I219178,I219486,I219503,I219172,I219534,I354450,I219551,I219160,I219582,I219599,I354444,I219616,I219642,I219650,I219169,I219681,I219698,I219175,I219729,I219163,I219787,I568340,I219813,I219830,I568346,I219861,I219869,I568361,I219886,I219903,I568352,I219920,I568349,I219937,I219954,I219971,I220002,I220019,I568364,I220036,I220081,I220098,I220129,I568358,I220146,I220177,I568343,I220194,I568355,I220211,I568367,I220237,I220245,I220276,I220293,I220324,I220382,I470710,I220408,I220425,I220374,I470692,I220456,I220464,I470698,I220481,I220498,I470713,I220515,I470704,I220532,I220549,I220566,I220371,I220597,I470716,I220614,I470695,I220631,I220356,I220368,I220676,I220693,I220362,I220724,I470701,I220741,I220350,I220772,I470707,I220789,I220806,I220832,I220840,I220359,I220871,I220888,I220365,I220919,I220353,I220977,I221003,I221020,I221051,I221059,I221076,I221093,I221110,I221127,I221144,I221161,I221192,I221209,I221226,I221271,I221288,I221319,I221336,I221367,I221384,I221401,I221427,I221435,I221466,I221483,I221514,I221572,I276450,I221598,I221606,I276462,I221632,I221640,I276453,I221657,I276456,I221674,I221691,I276459,I221708,I221558,I221739,I221756,I221773,I221790,I276465,I221555,I221546,I221835,I221549,I221543,I221880,I276471,I221897,I221914,I221552,I221945,I221962,I276468,I221979,I276474,I222005,I222013,I221540,I221564,I222058,I222075,I222092,I221561,I222150,I415922,I222176,I222184,I415913,I222210,I222218,I415907,I222235,I415919,I222252,I222269,I415910,I222286,I222317,I222334,I222351,I415916,I222368,I415901,I222413,I222458,I222475,I222492,I222523,I415904,I222540,I222557,I222583,I222591,I222636,I222653,I222670,I222728,I222754,I222762,I222788,I222796,I222813,I222830,I222847,I222864,I222714,I222895,I222912,I222929,I222946,I222711,I222702,I222991,I222705,I222699,I223036,I223053,I223070,I222708,I223101,I223118,I223135,I223161,I223169,I222696,I222720,I223214,I223231,I223248,I222717,I223306,I527008,I223332,I223340,I527020,I223366,I223374,I527011,I223391,I526999,I223408,I223425,I526996,I223442,I223292,I223473,I223490,I223507,I527002,I223524,I223289,I223280,I223569,I223283,I223277,I223614,I527017,I223631,I223648,I223286,I223679,I527005,I223696,I223713,I527014,I223739,I223747,I223274,I223298,I223792,I223809,I223826,I223295,I223884,I387007,I223910,I223918,I387004,I223944,I223952,I387001,I223969,I387028,I223986,I224003,I387016,I224020,I223870,I224051,I224068,I224085,I387022,I224102,I387013,I223867,I223858,I224147,I223861,I223855,I224192,I387010,I224209,I224226,I223864,I224257,I387025,I224274,I387019,I224291,I224317,I224325,I223852,I223876,I224370,I224387,I224404,I223873,I224462,I224488,I224496,I224522,I224530,I224547,I224564,I224581,I224598,I224448,I224629,I224646,I224663,I224680,I224445,I224436,I224725,I224439,I224433,I224770,I224787,I224804,I224442,I224835,I224852,I224869,I224895,I224903,I224430,I224454,I224948,I224965,I224982,I224451,I225040,I277028,I225066,I225074,I277040,I225100,I225108,I277031,I225125,I277034,I225142,I225159,I277037,I225176,I225026,I225207,I225224,I225241,I225258,I277043,I225023,I225014,I225303,I225017,I225011,I225348,I277049,I225365,I225382,I225020,I225413,I225430,I277046,I225447,I277052,I225473,I225481,I225008,I225032,I225526,I225543,I225560,I225029,I225618,I325977,I225644,I225652,I225678,I225686,I325974,I225703,I325989,I225720,I225737,I325983,I225754,I225604,I225785,I225802,I225819,I325980,I225836,I325971,I225601,I225592,I225881,I225595,I225589,I225926,I325992,I225943,I225960,I225598,I225991,I226008,I226025,I325986,I226051,I226059,I225586,I225610,I226104,I226121,I226138,I225607,I226196,I336517,I226222,I226230,I226256,I226264,I336514,I226281,I336529,I226298,I226315,I336523,I226332,I226182,I226363,I226380,I226397,I336520,I226414,I336511,I226179,I226170,I226459,I226173,I226167,I226504,I336532,I226521,I226538,I226176,I226569,I226586,I226603,I336526,I226629,I226637,I226164,I226188,I226682,I226699,I226716,I226185,I226774,I441214,I226800,I226808,I441220,I226834,I226842,I226859,I441217,I226876,I226893,I441235,I226910,I226760,I226941,I226958,I226975,I441238,I226992,I226757,I226748,I227037,I226751,I226745,I227082,I441223,I227099,I227116,I226754,I227147,I441229,I227164,I441226,I227181,I441232,I227207,I227215,I226742,I226766,I227260,I227277,I227294,I226763,I227352,I296102,I227378,I227386,I296114,I227412,I227420,I296105,I227437,I296108,I227454,I227471,I296111,I227488,I227338,I227519,I227536,I227553,I227570,I296117,I227335,I227326,I227615,I227329,I227323,I227660,I296123,I227677,I227694,I227332,I227725,I227742,I296120,I227759,I296126,I227785,I227793,I227320,I227344,I227838,I227855,I227872,I227341,I227930,I227956,I227964,I227990,I227998,I228015,I228032,I228049,I228066,I228097,I228114,I228131,I228148,I228193,I228238,I228255,I228272,I228303,I228320,I228337,I228363,I228371,I228416,I228433,I228450,I228508,I307084,I228534,I228542,I307096,I228568,I228576,I307087,I228593,I307090,I228610,I228627,I307093,I228644,I228494,I228675,I228692,I228709,I228726,I307099,I228491,I228482,I228771,I228485,I228479,I228816,I307105,I228833,I228850,I228488,I228881,I228898,I307102,I228915,I307108,I228941,I228949,I228476,I228500,I228994,I229011,I229028,I228497,I229086,I309396,I229112,I229120,I309408,I229146,I229154,I309399,I229171,I309402,I229188,I229205,I309405,I229222,I229253,I229270,I229287,I229304,I309411,I229349,I229394,I309417,I229411,I229428,I229459,I229476,I309414,I229493,I309420,I229519,I229527,I229572,I229589,I229606,I229664,I327558,I229690,I229698,I229724,I229732,I327555,I229749,I327570,I229766,I229783,I327564,I229800,I229650,I229831,I229848,I229865,I327561,I229882,I327552,I229647,I229638,I229927,I229641,I229635,I229972,I327573,I229989,I230006,I229644,I230037,I230054,I230071,I327567,I230097,I230105,I229632,I229656,I230150,I230167,I230184,I229653,I230242,I459710,I230268,I230276,I459716,I230302,I230310,I230327,I459713,I230344,I230361,I459731,I230378,I230228,I230409,I230426,I230443,I459734,I230460,I230225,I230216,I230505,I230219,I230213,I230550,I459719,I230567,I230584,I230222,I230615,I459725,I230632,I459722,I230649,I459728,I230675,I230683,I230210,I230234,I230728,I230745,I230762,I230231,I230820,I230846,I230854,I230880,I230888,I230905,I230922,I230939,I230956,I230806,I230987,I231004,I231021,I231038,I230803,I230794,I231083,I230797,I230791,I231128,I231145,I231162,I230800,I231193,I231210,I231227,I231253,I231261,I230788,I230812,I231306,I231323,I231340,I230809,I231398,I231424,I231432,I231458,I231466,I231483,I231500,I231517,I231534,I231565,I231582,I231599,I231616,I231661,I231706,I231723,I231740,I231771,I231788,I231805,I231831,I231839,I231884,I231901,I231918,I231976,I438362,I232002,I232010,I438353,I232036,I232044,I438347,I232061,I438359,I232078,I232095,I438350,I232112,I231962,I232143,I232160,I232177,I438356,I232194,I438341,I231959,I231950,I232239,I231953,I231947,I232284,I232301,I232318,I231956,I232349,I438344,I232366,I232383,I232409,I232417,I231944,I231968,I232462,I232479,I232496,I231965,I232554,I311130,I232580,I232588,I311142,I232614,I232622,I311133,I232639,I311136,I232656,I232673,I311139,I232690,I232721,I232738,I232755,I232772,I311145,I232817,I232862,I311151,I232879,I232896,I232927,I232944,I311148,I232961,I311154,I232987,I232995,I233040,I233057,I233074,I233132,I233158,I233166,I233192,I233200,I233217,I233234,I233251,I233268,I233299,I233316,I233333,I233350,I233395,I233440,I233457,I233474,I233505,I233522,I233539,I233565,I233573,I233618,I233635,I233652,I233710,I233736,I233744,I233770,I233778,I233795,I233812,I233829,I233846,I233696,I233877,I233894,I233911,I233928,I233693,I233684,I233973,I233687,I233681,I234018,I234035,I234052,I233690,I234083,I234100,I234117,I234143,I234151,I233678,I233702,I234196,I234213,I234230,I233699,I234288,I234314,I234322,I234348,I234356,I234373,I234390,I234407,I234424,I234455,I234472,I234489,I234506,I234551,I234596,I234613,I234630,I234661,I234678,I234695,I234721,I234729,I234774,I234791,I234808,I234866,I234892,I234900,I234926,I234934,I234951,I234968,I234985,I235002,I234852,I235033,I235050,I235067,I235084,I234849,I234840,I235129,I234843,I234837,I235174,I235191,I235208,I234846,I235239,I235256,I235273,I235299,I235307,I234834,I234858,I235352,I235369,I235386,I234855,I235444,I235470,I235478,I235504,I235512,I235529,I235546,I235563,I235580,I235430,I235611,I235628,I235645,I235662,I235427,I235418,I235707,I235421,I235415,I235752,I235769,I235786,I235424,I235817,I235834,I235851,I235877,I235885,I235412,I235436,I235930,I235947,I235964,I235433,I236022,I474738,I236048,I236056,I474744,I236082,I236090,I236107,I474741,I236124,I236141,I474759,I236158,I236008,I236189,I236206,I236223,I474762,I236240,I236005,I235996,I236285,I235999,I235993,I236330,I474747,I236347,I236364,I236002,I236395,I474753,I236412,I474750,I236429,I474756,I236455,I236463,I235990,I236014,I236508,I236525,I236542,I236011,I236600,I511204,I236626,I236634,I511198,I236660,I236668,I511207,I236685,I511186,I236702,I236719,I511195,I236736,I236586,I236767,I236784,I236801,I511210,I236818,I511189,I236583,I236574,I236863,I236577,I236571,I236908,I511192,I236925,I236942,I236580,I236973,I511201,I236990,I237007,I237033,I237041,I236568,I236592,I237086,I237103,I237120,I236589,I237178,I237204,I237212,I237238,I237246,I237263,I237280,I237297,I237314,I237345,I237362,I237379,I237396,I237441,I237486,I237503,I237520,I237551,I237568,I237585,I237611,I237619,I237664,I237681,I237698,I237756,I528742,I237782,I237790,I528754,I237816,I237824,I528745,I237841,I528733,I237858,I237875,I528730,I237892,I237742,I237923,I237940,I237957,I528736,I237974,I237739,I237730,I238019,I237733,I237727,I238064,I528751,I238081,I238098,I237736,I238129,I528739,I238146,I238163,I528748,I238189,I238197,I237724,I237748,I238242,I238259,I238276,I237745,I238334,I315754,I238360,I238368,I315766,I238394,I238402,I315757,I238419,I315760,I238436,I238453,I315763,I238470,I238320,I238501,I238518,I238535,I238552,I315769,I238317,I238308,I238597,I238311,I238305,I238642,I315775,I238659,I238676,I238314,I238707,I238724,I315772,I238741,I315778,I238767,I238775,I238302,I238326,I238820,I238837,I238854,I238323,I238912,I238938,I238946,I238972,I238980,I238997,I239014,I239031,I239048,I239079,I239096,I239113,I239130,I239175,I239220,I239237,I239254,I239285,I239302,I239319,I239345,I239353,I239398,I239415,I239432,I239490,I239516,I239524,I239550,I239558,I239575,I239592,I239609,I239626,I239657,I239674,I239691,I239708,I239753,I239798,I239815,I239832,I239863,I239880,I239897,I239923,I239931,I239976,I239993,I240010,I240068,I262578,I240094,I240102,I262590,I240128,I240136,I262581,I240153,I262584,I240170,I240187,I262587,I240204,I240054,I240235,I240252,I240269,I240286,I262593,I240051,I240042,I240331,I240045,I240039,I240376,I262599,I240393,I240410,I240048,I240441,I240458,I262596,I240475,I262602,I240501,I240509,I240036,I240060,I240554,I240571,I240588,I240057,I240646,I240672,I240680,I240706,I240714,I240731,I240748,I240765,I240782,I240632,I240813,I240830,I240847,I240864,I240629,I240620,I240909,I240623,I240617,I240954,I240971,I240988,I240626,I241019,I241036,I241053,I241079,I241087,I240614,I240638,I241132,I241149,I241166,I240635,I241224,I291478,I241250,I241258,I291490,I241284,I241292,I291481,I241309,I291484,I241326,I241343,I291487,I241360,I241391,I241408,I241425,I241442,I291493,I241487,I241532,I291499,I241549,I241566,I241597,I241614,I291496,I241631,I291502,I241657,I241665,I241710,I241727,I241744,I241802,I487454,I241828,I241836,I487460,I241862,I241870,I241887,I487457,I241904,I241921,I487475,I241938,I241788,I241969,I241986,I242003,I487478,I242020,I241785,I241776,I242065,I241779,I241773,I242110,I487463,I242127,I242144,I241782,I242175,I487469,I242192,I487466,I242209,I487472,I242235,I242243,I241770,I241794,I242288,I242305,I242322,I241791,I242380,I447572,I242406,I242414,I447578,I242440,I242448,I242465,I447575,I242482,I242499,I447593,I242516,I242547,I242564,I242581,I447596,I242598,I242643,I242688,I447581,I242705,I242722,I242753,I447587,I242770,I447584,I242787,I447590,I242813,I242821,I242866,I242883,I242900,I242958,I349692,I242984,I242992,I243018,I243026,I349689,I243043,I349704,I243060,I243077,I349698,I243094,I242944,I243125,I243142,I243159,I349695,I243176,I349686,I242941,I242932,I243221,I242935,I242929,I243266,I349707,I243283,I243300,I242938,I243331,I243348,I243365,I349701,I243391,I243399,I242926,I242950,I243444,I243461,I243478,I242947,I243536,I243562,I243570,I243596,I243604,I243621,I243638,I243655,I243672,I243703,I243720,I243737,I243754,I243799,I243844,I243861,I243878,I243909,I243926,I243943,I243969,I243977,I244022,I244039,I244056,I244114,I244140,I244148,I244174,I244182,I244199,I244216,I244233,I244250,I244100,I244281,I244298,I244315,I244332,I244097,I244088,I244377,I244091,I244085,I244422,I244439,I244456,I244094,I244487,I244504,I244521,I244547,I244555,I244082,I244106,I244600,I244617,I244634,I244103,I244692,I568935,I244718,I244726,I244752,I244760,I568959,I244777,I568941,I244794,I244811,I568956,I244828,I244678,I244859,I244876,I244893,I568938,I244910,I568947,I244675,I244666,I244955,I244669,I244663,I245000,I568944,I245017,I245034,I244672,I245065,I568953,I245082,I568962,I245099,I568950,I245125,I245133,I244660,I244684,I245178,I245195,I245212,I244681,I245270,I245296,I245304,I245330,I245338,I245355,I245372,I245389,I245406,I245256,I245437,I245454,I245471,I245488,I245253,I245244,I245533,I245247,I245241,I245578,I245595,I245612,I245250,I245643,I245660,I245677,I245703,I245711,I245238,I245262,I245756,I245773,I245790,I245259,I245848,I308240,I245874,I245882,I308252,I245908,I245916,I308243,I245933,I308246,I245950,I245967,I308249,I245984,I246015,I246032,I246049,I246066,I308255,I246111,I246156,I308261,I246173,I246190,I246221,I246238,I308258,I246255,I308264,I246281,I246289,I246334,I246351,I246368,I246426,I513924,I246452,I246460,I513918,I246486,I246494,I513927,I246511,I513906,I246528,I246545,I513915,I246562,I246412,I246593,I246610,I246627,I513930,I246644,I513909,I246409,I246400,I246689,I246403,I246397,I246734,I513912,I246751,I246768,I246406,I246799,I513921,I246816,I246833,I246859,I246867,I246394,I246418,I246912,I246929,I246946,I246415,I247004,I264890,I247030,I247038,I264902,I247064,I247072,I264893,I247089,I264896,I247106,I247123,I264899,I247140,I246990,I247171,I247188,I247205,I247222,I264905,I246987,I246978,I247267,I246981,I246975,I247312,I264911,I247329,I247346,I246984,I247377,I247394,I264908,I247411,I264914,I247437,I247445,I246972,I246996,I247490,I247507,I247524,I246993,I247582,I277606,I247608,I247616,I277618,I247642,I247650,I277609,I247667,I277612,I247684,I247701,I277615,I247718,I247568,I247749,I247766,I247783,I247800,I277621,I247565,I247556,I247845,I247559,I247553,I247890,I277627,I247907,I247924,I247562,I247955,I247972,I277624,I247989,I277630,I248015,I248023,I247550,I247574,I248068,I248085,I248102,I247571,I248160,I508484,I248186,I248194,I508478,I248220,I248228,I508487,I248245,I508466,I248262,I248279,I508475,I248296,I248327,I248344,I248361,I508490,I248378,I508469,I248423,I248468,I508472,I248485,I248502,I248533,I508481,I248550,I248567,I248593,I248601,I248646,I248663,I248680,I248738,I499014,I248764,I248772,I499020,I248798,I248806,I248823,I499017,I248840,I248857,I499035,I248874,I248724,I248905,I248922,I248939,I499038,I248956,I248721,I248712,I249001,I248715,I248709,I249046,I499023,I249063,I249080,I248718,I249111,I499029,I249128,I499026,I249145,I499032,I249171,I249179,I248706,I248730,I249224,I249241,I249258,I248727,I249316,I249342,I249350,I249376,I249384,I249401,I249418,I249435,I249452,I249483,I249500,I249517,I249534,I249579,I249624,I249641,I249658,I249689,I249706,I249723,I249749,I249757,I249802,I249819,I249836,I249894,I249920,I249928,I249954,I249962,I249979,I249996,I250013,I250030,I250061,I250078,I250095,I250112,I250157,I250202,I250219,I250236,I250267,I250284,I250301,I250327,I250335,I250380,I250397,I250414,I250472,I533864,I250498,I250506,I533882,I250532,I250540,I533879,I250557,I533870,I250574,I250591,I533867,I250608,I250458,I250639,I250656,I250673,I533873,I250690,I533888,I250455,I250446,I250735,I250449,I250443,I250780,I250797,I250814,I250452,I250845,I533885,I250862,I533876,I250879,I533891,I250905,I250913,I250440,I250464,I250958,I250975,I250992,I250461,I251050,I251076,I251084,I251110,I251118,I251135,I251152,I251169,I251186,I251036,I251217,I251234,I251251,I251268,I251033,I251024,I251313,I251027,I251021,I251358,I251375,I251392,I251030,I251423,I251440,I251457,I251483,I251491,I251018,I251042,I251536,I251553,I251570,I251039,I251628,I302460,I251654,I251662,I302472,I251688,I251696,I302463,I251713,I302466,I251730,I251747,I302469,I251764,I251795,I251812,I251829,I251846,I302475,I251891,I251936,I302481,I251953,I251970,I252001,I252018,I302478,I252035,I302484,I252061,I252069,I252114,I252131,I252148,I252206,I552870,I252232,I252240,I252266,I252274,I552894,I252291,I552876,I252308,I252325,I552891,I252342,I252192,I252373,I252390,I252407,I552873,I252424,I552882,I252189,I252180,I252469,I252183,I252177,I252514,I552879,I252531,I252548,I252186,I252579,I552888,I252596,I552897,I252613,I552885,I252639,I252647,I252174,I252198,I252692,I252709,I252726,I252195,I252784,I431630,I252810,I252818,I431621,I252844,I252852,I431615,I252869,I431627,I252886,I252903,I431618,I252920,I252770,I252951,I252968,I252985,I431624,I253002,I431609,I252767,I252758,I253047,I252761,I252755,I253092,I253109,I253126,I252764,I253157,I431612,I253174,I253191,I253217,I253225,I252752,I252776,I253270,I253287,I253304,I252773,I253362,I253388,I253396,I253422,I253430,I253447,I253464,I253481,I253498,I253529,I253546,I253563,I253580,I253625,I253670,I253687,I253704,I253735,I253752,I253769,I253795,I253803,I253848,I253865,I253882,I253940,I267202,I253966,I253974,I267214,I254000,I254008,I267205,I254025,I267208,I254042,I254059,I267211,I254076,I254107,I254124,I254141,I254158,I267217,I254203,I254248,I267223,I254265,I254282,I254313,I254330,I267220,I254347,I267226,I254373,I254381,I254426,I254443,I254460,I254518,I405095,I254544,I254552,I405092,I254578,I254586,I405089,I254603,I405116,I254620,I254637,I405104,I254654,I254685,I254702,I254719,I405110,I254736,I405101,I254781,I254826,I405098,I254843,I254860,I254891,I405113,I254908,I405107,I254925,I254951,I254959,I255004,I255021,I255038,I255096,I427142,I255122,I255130,I427133,I255156,I255164,I427127,I255181,I427139,I255198,I255215,I427130,I255232,I255263,I255280,I255297,I427136,I255314,I427121,I255359,I255404,I255421,I255438,I255469,I427124,I255486,I255503,I255529,I255537,I255582,I255599,I255616,I255674,I279340,I255700,I255708,I279352,I255734,I255742,I279343,I255759,I279346,I255776,I255793,I279349,I255810,I255841,I255858,I255875,I255892,I279355,I255937,I255982,I279361,I255999,I256016,I256047,I256064,I279358,I256081,I279364,I256107,I256115,I256160,I256177,I256194,I256252,I256278,I256286,I256312,I256320,I256337,I256354,I256371,I256388,I256419,I256436,I256453,I256470,I256515,I256560,I256577,I256594,I256625,I256642,I256659,I256685,I256693,I256738,I256755,I256772,I256830,I410909,I256856,I256864,I410906,I256890,I256898,I410903,I256915,I410930,I256932,I256949,I410918,I256966,I256997,I257014,I257031,I410924,I257048,I410915,I257093,I257138,I410912,I257155,I257172,I257203,I410927,I257220,I410921,I257237,I257263,I257271,I257316,I257333,I257350,I257408,I518904,I257434,I257442,I257459,I518928,I518910,I257476,I518916,I257502,I257510,I518922,I518907,I257536,I257544,I257561,I257578,I257595,I518919,I257635,I257643,I257660,I257677,I257694,I257725,I518925,I518913,I257742,I257768,I257776,I257807,I257838,I257855,I257886,I257986,I543972,I258012,I258020,I258037,I543957,I543945,I258054,I543960,I258080,I258088,I543963,I258114,I258122,I258139,I258156,I258173,I257969,I543951,I258213,I258221,I258238,I258255,I258272,I257972,I258303,I543948,I543954,I258320,I543969,I258346,I258354,I257954,I258385,I257963,I258416,I258433,I257975,I258464,I543966,I257966,I257957,I257960,I257978,I258564,I258590,I258598,I258615,I258632,I258658,I258666,I258692,I258700,I258717,I258734,I258751,I258547,I258791,I258799,I258816,I258833,I258850,I258550,I258881,I258898,I258924,I258932,I258532,I258963,I258541,I258994,I259011,I258553,I259042,I258544,I258535,I258538,I258556,I259142,I410281,I259168,I259176,I259193,I410257,I410272,I259210,I410284,I259236,I259244,I410269,I410260,I259270,I259278,I259295,I259312,I259329,I259125,I259369,I259377,I259394,I259411,I259428,I259128,I259459,I410275,I410266,I259476,I410278,I259502,I259510,I259110,I259541,I259119,I259572,I259589,I259131,I259620,I410263,I259122,I259113,I259116,I259134,I259720,I431054,I259746,I259754,I259771,I431051,I431069,I259788,I431066,I259814,I259822,I431048,I259848,I259856,I259873,I259890,I259907,I259703,I431060,I259947,I259955,I259972,I259989,I260006,I259706,I260037,I431063,I260054,I260080,I260088,I259688,I260119,I259697,I260150,I260167,I259709,I260198,I431057,I259700,I259691,I259694,I259712,I260298,I260324,I260332,I260349,I260366,I260392,I260400,I260426,I260434,I260451,I260468,I260485,I260281,I260525,I260533,I260550,I260567,I260584,I260284,I260615,I260632,I260658,I260666,I260266,I260697,I260275,I260728,I260745,I260287,I260776,I260278,I260269,I260272,I260290,I260876,I260902,I260910,I260927,I260944,I260970,I260978,I261004,I261012,I261029,I261046,I261063,I261103,I261111,I261128,I261145,I261162,I261193,I261210,I261236,I261244,I261275,I261306,I261323,I261354,I261454,I261480,I261488,I261505,I261522,I261548,I261556,I261582,I261590,I261607,I261624,I261641,I261437,I261681,I261689,I261706,I261723,I261740,I261440,I261771,I261788,I261814,I261822,I261422,I261853,I261431,I261884,I261901,I261443,I261932,I261434,I261425,I261428,I261446,I262032,I262058,I262066,I262083,I262100,I262126,I262134,I262160,I262168,I262185,I262202,I262219,I262015,I262259,I262267,I262284,I262301,I262318,I262018,I262349,I262366,I262392,I262400,I262000,I262431,I262009,I262462,I262479,I262021,I262510,I262012,I262003,I262006,I262024,I262610,I262636,I262644,I262661,I262678,I262704,I262712,I262738,I262746,I262763,I262780,I262797,I262837,I262845,I262862,I262879,I262896,I262927,I262944,I262970,I262978,I263009,I263040,I263057,I263088,I263188,I365061,I263214,I263222,I263239,I365037,I365052,I263256,I365064,I263282,I263290,I365049,I365040,I263316,I263324,I263341,I263358,I263375,I263171,I263415,I263423,I263440,I263457,I263474,I263174,I263505,I365055,I365046,I263522,I365058,I263548,I263556,I263156,I263587,I263165,I263618,I263635,I263177,I263666,I365043,I263168,I263159,I263162,I263180,I263766,I453370,I263792,I263800,I263817,I453352,I453364,I263834,I453367,I263860,I263868,I453361,I453358,I263894,I263902,I263919,I263936,I263953,I263749,I453376,I263993,I264001,I264018,I264035,I264052,I263752,I264083,I453355,I264100,I264126,I264134,I263734,I264165,I263743,I264196,I264213,I263755,I264244,I453373,I263746,I263737,I263740,I263758,I264344,I264370,I264378,I264395,I264412,I264438,I264446,I264472,I264480,I264497,I264514,I264531,I264571,I264579,I264596,I264613,I264630,I264661,I264678,I264704,I264712,I264743,I264774,I264791,I264822,I264922,I450480,I264948,I264956,I264973,I450462,I450474,I264990,I450477,I265016,I265024,I450471,I450468,I265050,I265058,I265075,I265092,I265109,I450486,I265149,I265157,I265174,I265191,I265208,I265239,I450465,I265256,I265282,I265290,I265321,I265352,I265369,I265400,I450483,I265500,I265526,I265534,I265551,I265568,I265594,I265602,I265628,I265636,I265653,I265670,I265687,I265727,I265735,I265752,I265769,I265786,I265817,I265834,I265860,I265868,I265899,I265930,I265947,I265978,I266078,I266104,I266112,I266129,I266146,I266172,I266180,I266206,I266214,I266231,I266248,I266265,I266061,I266305,I266313,I266330,I266347,I266364,I266064,I266395,I266412,I266438,I266446,I266046,I266477,I266055,I266508,I266525,I266067,I266556,I266058,I266049,I266052,I266070,I266656,I266682,I266690,I266707,I266724,I266750,I266758,I266784,I266792,I266809,I266826,I266843,I266639,I266883,I266891,I266908,I266925,I266942,I266642,I266973,I266990,I267016,I267024,I266624,I267055,I266633,I267086,I267103,I266645,I267134,I266636,I266627,I266630,I266648,I267234,I388963,I267260,I267268,I267285,I388939,I388954,I267302,I388966,I267328,I267336,I388951,I388942,I267362,I267370,I267387,I267404,I267421,I267461,I267469,I267486,I267503,I267520,I267551,I388957,I388948,I267568,I388960,I267594,I267602,I267633,I267664,I267681,I267712,I388945,I267812,I443544,I267838,I267846,I267863,I443526,I443538,I267880,I443541,I267906,I267914,I443535,I443532,I267940,I267948,I267965,I267982,I267999,I443550,I268039,I268047,I268064,I268081,I268098,I268129,I443529,I268146,I268172,I268180,I268211,I268242,I268259,I268290,I443547,I268390,I268416,I268424,I268441,I268458,I268484,I268492,I268518,I268526,I268543,I268560,I268577,I268373,I268617,I268625,I268642,I268659,I268676,I268376,I268707,I268724,I268750,I268758,I268358,I268789,I268367,I268820,I268837,I268379,I268868,I268370,I268361,I268364,I268382,I268968,I548732,I268994,I269002,I269019,I548717,I548705,I269036,I548720,I269062,I269070,I548723,I269096,I269104,I269121,I269138,I269155,I268951,I548711,I269195,I269203,I269220,I269237,I269254,I268954,I269285,I548708,I548714,I269302,I548729,I269328,I269336,I268936,I269367,I268945,I269398,I269415,I268957,I269446,I548726,I268948,I268939,I268942,I268960,I269546,I426005,I269572,I269580,I269597,I426002,I426020,I269614,I426017,I269640,I269648,I425999,I269674,I269682,I269699,I269716,I269733,I269529,I426011,I269773,I269781,I269798,I269815,I269832,I269532,I269863,I426014,I269880,I269906,I269914,I269514,I269945,I269523,I269976,I269993,I269535,I270024,I426008,I269526,I269517,I269520,I269538,I270124,I270150,I270158,I270175,I270192,I270218,I270226,I270252,I270260,I270277,I270294,I270311,I270107,I270351,I270359,I270376,I270393,I270410,I270110,I270441,I270458,I270484,I270492,I270092,I270523,I270101,I270554,I270571,I270113,I270602,I270104,I270095,I270098,I270116,I270702,I546947,I270728,I270736,I270753,I546932,I546920,I270770,I546935,I270796,I270804,I546938,I270830,I270838,I270855,I270872,I270889,I546926,I270929,I270937,I270954,I270971,I270988,I271019,I546923,I546929,I271036,I546944,I271062,I271070,I271101,I271132,I271149,I271180,I546941,I271280,I363123,I271306,I271314,I271331,I363099,I363114,I271348,I363126,I271374,I271382,I363111,I363102,I271408,I271416,I271433,I271450,I271467,I271263,I271507,I271515,I271532,I271549,I271566,I271266,I271597,I363117,I363108,I271614,I363120,I271640,I271648,I271248,I271679,I271257,I271710,I271727,I271269,I271758,I363105,I271260,I271251,I271254,I271272,I271858,I271884,I271892,I271909,I271926,I271952,I271960,I271986,I271994,I272011,I272028,I272045,I271841,I272085,I272093,I272110,I272127,I272144,I271844,I272175,I272192,I272218,I272226,I271826,I272257,I271835,I272288,I272305,I271847,I272336,I271838,I271829,I271832,I271850,I272436,I272462,I272470,I272487,I272504,I272530,I272538,I272564,I272572,I272589,I272606,I272623,I272419,I272663,I272671,I272688,I272705,I272722,I272422,I272753,I272770,I272796,I272804,I272404,I272835,I272413,I272866,I272883,I272425,I272914,I272416,I272407,I272410,I272428,I273014,I390255,I273040,I273048,I273065,I390231,I390246,I273082,I390258,I273108,I273116,I390243,I390234,I273142,I273150,I273167,I273184,I273201,I273241,I273249,I273266,I273283,I273300,I273331,I390249,I390240,I273348,I390252,I273374,I273382,I273413,I273444,I273461,I273492,I390237,I273592,I366353,I273618,I273626,I273643,I366329,I366344,I273660,I366356,I273686,I273694,I366341,I366332,I273720,I273728,I273745,I273762,I273779,I273575,I273819,I273827,I273844,I273861,I273878,I273578,I273909,I366347,I366338,I273926,I366350,I273952,I273960,I273560,I273991,I273569,I274022,I274039,I273581,I274070,I366335,I273572,I273563,I273566,I273584,I274170,I517170,I274196,I274204,I274221,I517194,I517176,I274238,I517182,I274264,I274272,I517188,I517173,I274298,I274306,I274323,I274340,I274357,I517185,I274397,I274405,I274422,I274439,I274456,I274487,I517191,I517179,I274504,I274530,I274538,I274569,I274600,I274617,I274648,I274748,I466664,I274774,I274782,I274799,I466646,I466658,I274816,I466661,I274842,I274850,I466655,I466652,I274876,I274884,I274901,I274918,I274935,I274731,I466670,I274975,I274983,I275000,I275017,I275034,I274734,I275065,I466649,I275082,I275108,I275116,I274716,I275147,I274725,I275178,I275195,I274737,I275226,I466667,I274728,I274719,I274722,I274740,I275326,I389609,I275352,I275360,I275377,I389585,I389600,I275394,I389612,I275420,I275428,I389597,I389588,I275454,I275462,I275479,I275496,I275513,I275309,I275553,I275561,I275578,I275595,I275612,I275312,I275643,I389603,I389594,I275660,I389606,I275686,I275694,I275294,I275725,I275303,I275756,I275773,I275315,I275804,I389591,I275306,I275297,I275300,I275318,I275904,I275930,I275938,I275955,I275972,I275998,I276006,I276032,I276040,I276057,I276074,I276091,I275887,I276131,I276139,I276156,I276173,I276190,I275890,I276221,I276238,I276264,I276272,I275872,I276303,I275881,I276334,I276351,I275893,I276382,I275884,I275875,I275878,I275896,I276482,I276508,I276516,I276533,I276550,I276576,I276584,I276610,I276618,I276635,I276652,I276669,I276709,I276717,I276734,I276751,I276768,I276799,I276816,I276842,I276850,I276881,I276912,I276929,I276960,I277060,I323351,I277086,I277094,I277111,I323339,I323357,I277128,I323354,I277154,I277162,I323345,I323342,I277188,I277196,I277213,I277230,I277247,I323336,I277287,I277295,I277312,I277329,I277346,I277377,I277394,I277420,I277428,I277459,I277490,I277507,I277538,I323348,I277638,I277664,I277672,I277689,I277706,I277732,I277740,I277766,I277774,I277791,I277808,I277825,I277865,I277873,I277890,I277907,I277924,I277955,I277972,I277998,I278006,I278037,I278068,I278085,I278116,I278216,I357079,I278242,I278250,I278267,I357067,I357085,I278284,I357082,I278310,I278318,I357073,I357070,I278344,I278352,I278369,I278386,I278403,I278199,I357064,I278443,I278451,I278468,I278485,I278502,I278202,I278533,I278550,I278576,I278584,I278184,I278615,I278193,I278646,I278663,I278205,I278694,I357076,I278196,I278187,I278190,I278208,I278794,I519482,I278820,I278828,I278845,I519506,I519488,I278862,I519494,I278888,I278896,I519500,I519485,I278922,I278930,I278947,I278964,I278981,I278777,I519497,I279021,I279029,I279046,I279063,I279080,I278780,I279111,I519503,I519491,I279128,I279154,I279162,I278762,I279193,I278771,I279224,I279241,I278783,I279272,I278774,I278765,I278768,I278786,I279372,I527574,I279398,I279406,I279423,I527598,I527580,I279440,I527586,I279466,I279474,I527592,I527577,I279500,I279508,I279525,I279542,I279559,I527589,I279599,I279607,I279624,I279641,I279658,I279689,I527595,I527583,I279706,I279732,I279740,I279771,I279802,I279819,I279850,I279950,I346539,I279976,I279984,I280001,I346527,I346545,I280018,I346542,I280044,I280052,I346533,I346530,I280078,I280086,I280103,I280120,I280137,I346524,I280177,I280185,I280202,I280219,I280236,I280267,I280284,I280310,I280318,I280349,I280380,I280397,I280428,I346536,I280528,I280554,I280562,I280579,I280596,I280622,I280630,I280656,I280664,I280681,I280698,I280715,I280511,I280755,I280763,I280780,I280797,I280814,I280514,I280845,I280862,I280888,I280896,I280496,I280927,I280505,I280958,I280975,I280517,I281006,I280508,I280499,I280502,I280520,I281106,I408343,I281132,I281140,I281157,I408319,I408334,I281174,I408346,I281200,I281208,I408331,I408322,I281234,I281242,I281259,I281276,I281293,I281089,I281333,I281341,I281358,I281375,I281392,I281092,I281423,I408337,I408328,I281440,I408340,I281466,I281474,I281074,I281505,I281083,I281536,I281553,I281095,I281584,I408325,I281086,I281077,I281080,I281098,I281684,I281710,I281718,I281735,I281752,I281778,I281786,I281812,I281820,I281837,I281854,I281871,I281911,I281919,I281936,I281953,I281970,I282001,I282018,I282044,I282052,I282083,I282114,I282131,I282162,I282262,I485738,I282288,I282296,I282313,I485720,I485732,I282330,I485735,I282356,I282364,I485729,I485726,I282390,I282398,I282415,I282432,I282449,I485744,I282489,I282497,I282514,I282531,I282548,I282579,I485723,I282596,I282622,I282630,I282661,I282692,I282709,I282740,I485741,I282840,I282866,I282874,I282891,I282908,I282934,I282942,I282968,I282976,I282993,I283010,I283027,I282823,I283067,I283075,I283092,I283109,I283126,I282826,I283157,I283174,I283200,I283208,I282808,I283239,I282817,I283270,I283287,I282829,I283318,I282820,I282811,I282814,I282832,I283418,I283444,I283452,I283469,I283486,I283512,I283520,I283546,I283554,I283571,I283588,I283605,I283401,I283645,I283653,I283670,I283687,I283704,I283404,I283735,I283752,I283778,I283786,I283386,I283817,I283395,I283848,I283865,I283407,I283896,I283398,I283389,I283392,I283410,I283996,I284022,I284030,I284047,I284064,I284090,I284098,I284124,I284132,I284149,I284166,I284183,I283979,I284223,I284231,I284248,I284265,I284282,I283982,I284313,I284330,I284356,I284364,I283964,I284395,I283973,I284426,I284443,I283985,I284474,I283976,I283967,I283970,I283988,I284574,I375397,I284600,I284608,I284625,I375373,I375388,I284642,I375400,I284668,I284676,I375385,I375376,I284702,I284710,I284727,I284744,I284761,I284557,I284801,I284809,I284826,I284843,I284860,I284560,I284891,I375391,I375382,I284908,I375394,I284934,I284942,I284542,I284973,I284551,I285004,I285021,I284563,I285052,I375379,I284554,I284545,I284548,I284566,I285152,I285178,I285186,I285203,I285220,I285246,I285254,I285280,I285288,I285305,I285322,I285339,I285135,I285379,I285387,I285404,I285421,I285438,I285138,I285469,I285486,I285512,I285520,I285120,I285551,I285129,I285582,I285599,I285141,I285630,I285132,I285123,I285126,I285144,I285730,I285756,I285764,I285781,I285798,I285824,I285832,I285858,I285866,I285883,I285900,I285917,I285713,I285957,I285965,I285982,I285999,I286016,I285716,I286047,I286064,I286090,I286098,I285698,I286129,I285707,I286160,I286177,I285719,I286208,I285710,I285701,I285704,I285722,I286308,I383795,I286334,I286342,I286359,I383771,I383786,I286376,I383798,I286402,I286410,I383783,I383774,I286436,I286444,I286461,I286478,I286495,I286291,I286535,I286543,I286560,I286577,I286594,I286294,I286625,I383789,I383780,I286642,I383792,I286668,I286676,I286276,I286707,I286285,I286738,I286755,I286297,I286786,I383777,I286288,I286279,I286282,I286300,I286886,I286912,I286920,I286937,I286954,I286980,I286988,I287014,I287022,I287039,I287056,I287073,I286869,I287113,I287121,I287138,I287155,I287172,I286872,I287203,I287220,I287246,I287254,I286854,I287285,I286863,I287316,I287333,I286875,I287364,I286866,I286857,I286860,I286878,I287464,I287490,I287498,I287515,I287532,I287558,I287566,I287592,I287600,I287617,I287634,I287651,I287447,I287691,I287699,I287716,I287733,I287750,I287450,I287781,I287798,I287824,I287832,I287432,I287863,I287441,I287894,I287911,I287453,I287942,I287444,I287435,I287438,I287456,I288042,I288068,I288076,I288093,I288110,I288136,I288144,I288170,I288178,I288195,I288212,I288229,I288269,I288277,I288294,I288311,I288328,I288359,I288376,I288402,I288410,I288441,I288472,I288489,I288520,I288620,I464352,I288646,I288654,I288671,I464334,I464346,I288688,I464349,I288714,I288722,I464343,I464340,I288748,I288756,I288773,I288790,I288807,I464358,I288847,I288855,I288872,I288889,I288906,I288937,I464337,I288954,I288980,I288988,I289019,I289050,I289067,I289098,I464355,I289198,I289224,I289232,I289249,I289266,I289292,I289300,I289326,I289334,I289351,I289368,I289385,I289181,I289425,I289433,I289450,I289467,I289484,I289184,I289515,I289532,I289558,I289566,I289166,I289597,I289175,I289628,I289645,I289187,I289676,I289178,I289169,I289172,I289190,I289776,I397361,I289802,I289810,I289827,I397337,I397352,I289844,I397364,I289870,I289878,I397349,I397340,I289904,I289912,I289929,I289946,I289963,I289759,I290003,I290011,I290028,I290045,I290062,I289762,I290093,I397355,I397346,I290110,I397358,I290136,I290144,I289744,I290175,I289753,I290206,I290223,I289765,I290254,I397343,I289756,I289747,I289750,I289768,I290354,I347066,I290380,I290388,I290405,I347054,I347072,I290422,I347069,I290448,I290456,I347060,I347057,I290482,I290490,I290507,I290524,I290541,I347051,I290581,I290589,I290606,I290623,I290640,I290671,I290688,I290714,I290722,I290753,I290784,I290801,I290832,I347063,I290932,I331256,I290958,I290966,I290983,I331244,I331262,I291000,I331259,I291026,I291034,I331250,I331247,I291060,I291068,I291085,I291102,I291119,I290915,I331241,I291159,I291167,I291184,I291201,I291218,I290918,I291249,I291266,I291292,I291300,I290900,I291331,I290909,I291362,I291379,I290921,I291410,I331253,I290912,I290903,I290906,I290924,I291510,I456260,I291536,I291544,I291561,I456242,I456254,I291578,I456257,I291604,I291612,I456251,I456248,I291638,I291646,I291663,I291680,I291697,I456266,I291737,I291745,I291762,I291779,I291796,I291827,I456245,I291844,I291870,I291878,I291909,I291940,I291957,I291988,I456263,I292088,I376043,I292114,I292122,I292139,I376019,I376034,I292156,I376046,I292182,I292190,I376031,I376022,I292216,I292224,I292241,I292258,I292275,I292071,I292315,I292323,I292340,I292357,I292374,I292074,I292405,I376037,I376028,I292422,I376040,I292448,I292456,I292056,I292487,I292065,I292518,I292535,I292077,I292566,I376025,I292068,I292059,I292062,I292080,I292666,I422078,I292692,I292700,I292717,I422075,I422093,I292734,I422090,I292760,I292768,I422072,I292794,I292802,I292819,I292836,I292853,I422084,I292893,I292901,I292918,I292935,I292952,I292983,I422087,I293000,I293026,I293034,I293065,I293096,I293113,I293144,I422081,I293244,I293270,I293278,I293295,I293312,I293338,I293346,I293372,I293380,I293397,I293414,I293431,I293471,I293479,I293496,I293513,I293530,I293561,I293578,I293604,I293612,I293643,I293674,I293691,I293722,I293822,I505746,I293848,I293856,I293873,I505749,I505758,I293890,I505761,I293916,I293924,I505770,I505752,I293950,I293958,I293975,I293992,I294009,I293805,I294049,I294057,I294074,I294091,I294108,I293808,I294139,I505767,I294156,I505764,I294182,I294190,I293790,I294221,I293799,I294252,I294269,I293811,I294300,I505755,I293802,I293793,I293796,I293814,I294400,I294426,I294434,I294451,I294468,I294494,I294502,I294528,I294536,I294553,I294570,I294587,I294627,I294635,I294652,I294669,I294686,I294717,I294734,I294760,I294768,I294799,I294830,I294847,I294878,I294978,I295004,I295012,I295029,I295046,I295072,I295080,I295106,I295114,I295131,I295148,I295165,I295205,I295213,I295230,I295247,I295264,I295295,I295312,I295338,I295346,I295377,I295408,I295425,I295456,I295556,I295582,I295590,I295607,I295624,I295650,I295658,I295684,I295692,I295709,I295726,I295743,I295539,I295783,I295791,I295808,I295825,I295842,I295542,I295873,I295890,I295916,I295924,I295524,I295955,I295533,I295986,I296003,I295545,I296034,I295536,I295527,I295530,I295548,I296134,I557062,I296160,I296168,I296185,I557047,I557035,I296202,I557050,I296228,I296236,I557053,I296262,I296270,I296287,I296304,I296321,I557041,I296361,I296369,I296386,I296403,I296420,I296451,I557038,I557044,I296468,I557059,I296494,I296502,I296533,I296564,I296581,I296612,I557056,I296712,I424322,I296738,I296746,I296763,I424319,I424337,I296780,I424334,I296806,I296814,I424316,I296840,I296848,I296865,I296882,I296899,I424328,I296939,I296947,I296964,I296981,I296998,I297029,I424331,I297046,I297072,I297080,I297111,I297142,I297159,I297190,I424325,I297290,I340215,I297316,I297324,I297341,I340203,I340221,I297358,I340218,I297384,I297392,I340209,I340206,I297418,I297426,I297443,I297460,I297477,I297273,I340200,I297517,I297525,I297542,I297559,I297576,I297276,I297607,I297624,I297650,I297658,I297258,I297689,I297267,I297720,I297737,I297279,I297768,I340212,I297270,I297261,I297264,I297282,I297868,I297894,I297902,I297919,I297936,I297962,I297970,I297996,I298004,I298021,I298038,I298055,I297851,I298095,I298103,I298120,I298137,I298154,I297854,I298185,I298202,I298228,I298236,I297836,I298267,I297845,I298298,I298315,I297857,I298346,I297848,I297839,I297842,I297860,I298446,I298472,I298480,I298497,I298514,I298540,I298548,I298574,I298582,I298599,I298616,I298633,I298429,I298673,I298681,I298698,I298715,I298732,I298432,I298763,I298780,I298806,I298814,I298414,I298845,I298423,I298876,I298893,I298435,I298924,I298426,I298417,I298420,I298438,I299024,I299050,I299058,I299075,I299092,I299118,I299126,I299152,I299160,I299177,I299194,I299211,I299251,I299259,I299276,I299293,I299310,I299341,I299358,I299384,I299392,I299423,I299454,I299471,I299502,I299602,I559442,I299628,I299636,I299653,I559427,I559415,I299670,I559430,I299696,I299704,I559433,I299730,I299738,I299755,I299772,I299789,I299585,I559421,I299829,I299837,I299854,I299871,I299888,I299588,I299919,I559418,I559424,I299936,I559439,I299962,I299970,I299570,I300001,I299579,I300032,I300049,I299591,I300080,I559436,I299582,I299573,I299576,I299594,I300180,I300206,I300214,I300231,I300248,I300274,I300282,I300308,I300316,I300333,I300350,I300367,I300163,I300407,I300415,I300432,I300449,I300466,I300166,I300497,I300514,I300540,I300548,I300148,I300579,I300157,I300610,I300627,I300169,I300658,I300160,I300151,I300154,I300172,I300758,I334945,I300784,I300792,I300809,I334933,I334951,I300826,I334948,I300852,I300860,I334939,I334936,I300886,I300894,I300911,I300928,I300945,I300741,I334930,I300985,I300993,I301010,I301027,I301044,I300744,I301075,I301092,I301118,I301126,I300726,I301157,I300735,I301188,I301205,I300747,I301236,I334942,I300738,I300729,I300732,I300750,I301336,I301362,I301370,I301387,I301404,I301430,I301438,I301464,I301472,I301489,I301506,I301523,I301319,I301563,I301571,I301588,I301605,I301622,I301322,I301653,I301670,I301696,I301704,I301304,I301735,I301313,I301766,I301783,I301325,I301814,I301316,I301307,I301310,I301328,I301914,I301940,I301948,I301965,I301982,I302008,I302016,I302042,I302050,I302067,I302084,I302101,I301897,I302141,I302149,I302166,I302183,I302200,I301900,I302231,I302248,I302274,I302282,I301882,I302313,I301891,I302344,I302361,I301903,I302392,I301894,I301885,I301888,I301906,I302492,I302518,I302526,I302543,I302560,I302586,I302594,I302620,I302628,I302645,I302662,I302679,I302719,I302727,I302744,I302761,I302778,I302809,I302826,I302852,I302860,I302891,I302922,I302939,I302970,I303070,I422639,I303096,I303104,I303121,I422636,I422654,I303138,I422651,I303164,I303172,I422633,I303198,I303206,I303223,I303240,I303257,I303053,I422645,I303297,I303305,I303322,I303339,I303356,I303056,I303387,I422648,I303404,I303430,I303438,I303038,I303469,I303047,I303500,I303517,I303059,I303548,I422642,I303050,I303041,I303044,I303062,I303648,I386379,I303674,I303682,I303699,I386355,I386370,I303716,I386382,I303742,I303750,I386367,I386358,I303776,I303784,I303801,I303818,I303835,I303631,I303875,I303883,I303900,I303917,I303934,I303634,I303965,I386373,I386364,I303982,I386376,I304008,I304016,I303616,I304047,I303625,I304078,I304095,I303637,I304126,I386361,I303628,I303619,I303622,I303640,I304226,I304252,I304260,I304277,I304294,I304320,I304328,I304354,I304362,I304379,I304396,I304413,I304209,I304453,I304461,I304478,I304495,I304512,I304212,I304543,I304560,I304586,I304594,I304194,I304625,I304203,I304656,I304673,I304215,I304704,I304206,I304197,I304200,I304218,I304804,I449902,I304830,I304838,I304855,I449884,I449896,I304872,I449899,I304898,I304906,I449893,I449890,I304932,I304940,I304957,I304974,I304991,I449908,I305031,I305039,I305056,I305073,I305090,I305121,I449887,I305138,I305164,I305172,I305203,I305234,I305251,I305282,I449905,I305382,I305408,I305416,I305433,I305450,I305476,I305484,I305510,I305518,I305535,I305552,I305569,I305609,I305617,I305634,I305651,I305668,I305699,I305716,I305742,I305750,I305781,I305812,I305829,I305860,I305960,I305986,I305994,I306011,I306028,I306054,I306062,I306088,I306096,I306113,I306130,I306147,I305943,I306187,I306195,I306212,I306229,I306246,I305946,I306277,I306294,I306320,I306328,I305928,I306359,I305937,I306390,I306407,I305949,I306438,I305940,I305931,I305934,I305952,I306538,I352336,I306564,I306572,I306589,I352324,I352342,I306606,I352339,I306632,I306640,I352330,I352327,I306666,I306674,I306691,I306708,I306725,I352321,I306765,I306773,I306790,I306807,I306824,I306855,I306872,I306898,I306906,I306937,I306968,I306985,I307016,I352333,I307116,I307142,I307150,I307167,I307184,I307210,I307218,I307244,I307252,I307269,I307286,I307303,I307343,I307351,I307368,I307385,I307402,I307433,I307450,I307476,I307484,I307515,I307546,I307563,I307594,I307694,I334418,I307720,I307728,I307745,I334406,I334424,I307762,I334421,I307788,I307796,I334412,I334409,I307822,I307830,I307847,I307864,I307881,I307677,I334403,I307921,I307929,I307946,I307963,I307980,I307680,I308011,I308028,I308054,I308062,I307662,I308093,I307671,I308124,I308141,I307683,I308172,I334415,I307674,I307665,I307668,I307686,I308272,I308298,I308306,I308323,I308340,I308366,I308374,I308400,I308408,I308425,I308442,I308459,I308499,I308507,I308524,I308541,I308558,I308589,I308606,I308632,I308640,I308671,I308702,I308719,I308750,I308850,I329675,I308876,I308884,I308901,I329663,I329681,I308918,I329678,I308944,I308952,I329669,I329666,I308978,I308986,I309003,I309020,I309037,I329660,I309077,I309085,I309102,I309119,I309136,I309167,I309184,I309210,I309218,I309249,I309280,I309297,I309328,I329672,I309428,I309454,I309462,I309479,I309496,I309522,I309530,I309556,I309564,I309581,I309598,I309615,I309655,I309663,I309680,I309697,I309714,I309745,I309762,I309788,I309796,I309827,I309858,I309875,I309906,I310006,I417590,I310032,I310040,I310057,I417587,I417605,I310074,I417602,I310100,I310108,I417584,I310134,I310142,I310159,I310176,I310193,I309989,I417596,I310233,I310241,I310258,I310275,I310292,I309992,I310323,I417599,I310340,I310366,I310374,I309974,I310405,I309983,I310436,I310453,I309995,I310484,I417593,I309986,I309977,I309980,I309998,I310584,I561227,I310610,I310618,I310635,I561212,I561200,I310652,I561215,I310678,I310686,I561218,I310712,I310720,I310737,I310754,I310771,I561206,I310811,I310819,I310836,I310853,I310870,I310901,I561203,I561209,I310918,I561224,I310944,I310952,I310983,I311014,I311031,I311062,I561221,I311162,I311188,I311196,I311213,I311230,I311256,I311264,I311290,I311298,I311315,I311332,I311349,I311389,I311397,I311414,I311431,I311448,I311479,I311496,I311522,I311530,I311561,I311592,I311609,I311640,I311740,I311766,I311774,I311791,I311808,I311834,I311842,I311868,I311876,I311893,I311910,I311927,I311967,I311975,I311992,I312009,I312026,I312057,I312074,I312100,I312108,I312139,I312170,I312187,I312218,I312318,I312344,I312352,I312369,I312386,I312412,I312420,I312446,I312454,I312471,I312488,I312505,I312545,I312553,I312570,I312587,I312604,I312635,I312652,I312678,I312686,I312717,I312748,I312765,I312796,I312896,I312922,I312930,I312947,I312964,I312990,I312998,I313024,I313032,I313049,I313066,I313083,I313123,I313131,I313148,I313165,I313182,I313213,I313230,I313256,I313264,I313295,I313326,I313343,I313374,I313474,I506834,I313500,I313508,I313525,I506837,I506846,I313542,I506849,I313568,I313576,I506858,I506840,I313602,I313610,I313627,I313644,I313661,I313457,I313701,I313709,I313726,I313743,I313760,I313460,I313791,I506855,I313808,I506852,I313834,I313842,I313442,I313873,I313451,I313904,I313921,I313463,I313952,I506843,I313454,I313445,I313448,I313466,I314052,I361831,I314078,I314086,I314103,I361807,I361822,I314120,I361834,I314146,I314154,I361819,I361810,I314180,I314188,I314205,I314222,I314239,I314035,I314279,I314287,I314304,I314321,I314338,I314038,I314369,I361825,I361816,I314386,I361828,I314412,I314420,I314020,I314451,I314029,I314482,I314499,I314041,I314530,I361813,I314032,I314023,I314026,I314044,I314630,I314656,I314664,I314681,I314698,I314724,I314732,I314758,I314766,I314783,I314800,I314817,I314613,I314857,I314865,I314882,I314899,I314916,I314616,I314947,I314964,I314990,I314998,I314598,I315029,I314607,I315060,I315077,I314619,I315108,I314610,I314601,I314604,I314622,I315208,I401883,I315234,I315242,I315259,I401859,I401874,I315276,I401886,I315302,I315310,I401871,I401862,I315336,I315344,I315361,I315378,I315395,I315435,I315443,I315460,I315477,I315494,I315525,I401877,I401868,I315542,I401880,I315568,I315576,I315607,I315638,I315655,I315686,I401865,I315786,I430493,I315812,I315820,I315837,I430490,I430508,I315854,I430505,I315880,I315888,I430487,I315914,I315922,I315939,I315956,I315973,I430499,I316013,I316021,I316038,I316055,I316072,I316103,I430502,I316120,I316146,I316154,I316185,I316216,I316233,I316264,I430496,I316364,I316390,I316398,I316415,I316432,I316458,I316466,I316492,I316500,I316517,I316534,I316551,I316347,I316591,I316599,I316616,I316633,I316650,I316350,I316681,I316698,I316724,I316732,I316332,I316763,I316341,I316794,I316811,I316353,I316842,I316344,I316335,I316338,I316356,I316942,I316968,I316976,I316993,I317010,I317036,I317044,I317070,I317078,I317095,I317112,I317129,I317169,I317177,I317194,I317211,I317228,I317259,I317276,I317302,I317310,I317341,I317372,I317389,I317420,I317520,I322297,I317546,I317554,I317571,I322285,I322303,I317588,I322300,I317614,I317622,I322291,I322288,I317648,I317656,I317673,I317690,I317707,I322282,I317747,I317755,I317772,I317789,I317806,I317837,I317854,I317880,I317888,I317919,I317950,I317967,I317998,I322294,I318095,I497298,I318121,I318129,I318146,I497280,I318163,I497286,I318189,I318084,I497283,I318220,I318228,I497292,I318245,I318271,I318279,I318087,I497304,I318319,I318078,I318069,I318355,I497295,I497289,I318372,I318398,I318406,I318423,I318072,I318454,I497301,I318471,I318488,I318081,I318519,I318066,I318550,I318567,I318075,I318622,I396048,I318648,I318656,I318673,I396063,I396045,I318690,I318716,I318611,I396054,I318747,I318755,I396072,I318772,I318798,I318806,I318614,I396069,I318846,I318605,I318596,I318882,I396066,I396057,I318899,I396051,I318925,I318933,I318950,I318599,I318981,I396060,I318998,I319015,I318608,I319046,I318593,I319077,I319094,I318602,I319149,I319175,I319183,I319200,I319217,I319243,I319274,I319282,I319299,I319325,I319333,I319373,I319409,I319426,I319452,I319460,I319477,I319508,I319525,I319542,I319573,I319604,I319621,I319676,I319702,I319710,I319727,I319744,I319770,I319665,I319801,I319809,I319826,I319852,I319860,I319668,I319900,I319659,I319650,I319936,I319953,I319979,I319987,I320004,I319653,I320035,I320052,I320069,I319662,I320100,I319647,I320131,I320148,I319656,I320203,I320229,I320237,I320254,I320271,I320297,I320328,I320336,I320353,I320379,I320387,I320427,I320463,I320480,I320506,I320514,I320531,I320562,I320579,I320596,I320627,I320658,I320675,I320730,I419837,I320756,I320764,I320781,I419846,I419834,I320798,I419831,I320824,I320855,I320863,I419828,I320880,I320906,I320914,I320954,I320990,I419849,I419840,I321007,I419843,I321033,I321041,I321058,I321089,I321106,I321123,I321154,I321185,I321202,I321257,I321283,I321291,I321308,I321325,I321351,I321382,I321390,I321407,I321433,I321441,I321481,I321517,I321534,I321560,I321568,I321585,I321616,I321633,I321650,I321681,I321712,I321729,I321784,I321810,I321818,I321835,I321852,I321878,I321909,I321917,I321934,I321960,I321968,I322008,I322044,I322061,I322087,I322095,I322112,I322143,I322160,I322177,I322208,I322239,I322256,I322311,I322337,I322345,I322362,I322379,I322405,I322436,I322444,I322461,I322487,I322495,I322535,I322571,I322588,I322614,I322622,I322639,I322670,I322687,I322704,I322735,I322766,I322783,I322838,I542175,I322864,I322872,I322889,I542172,I542181,I322906,I542160,I322932,I542163,I322963,I322971,I542178,I322988,I323014,I323022,I542184,I323062,I323098,I542166,I542187,I323115,I542169,I323141,I323149,I323166,I323197,I323214,I323231,I323262,I323293,I323310,I323365,I323391,I323399,I323416,I323433,I323459,I323490,I323498,I323515,I323541,I323549,I323589,I323625,I323642,I323668,I323676,I323693,I323724,I323741,I323758,I323789,I323820,I323837,I323892,I323918,I323926,I323943,I323960,I323986,I324017,I324025,I324042,I324068,I324076,I324116,I324152,I324169,I324195,I324203,I324220,I324251,I324268,I324285,I324316,I324347,I324364,I324419,I324445,I324453,I324470,I324487,I324513,I324408,I324544,I324552,I324569,I324595,I324603,I324411,I324643,I324402,I324393,I324679,I324696,I324722,I324730,I324747,I324396,I324778,I324795,I324812,I324405,I324843,I324390,I324874,I324891,I324399,I324946,I473600,I324972,I324980,I324997,I473582,I325014,I473588,I325040,I473585,I325071,I325079,I473594,I325096,I325122,I325130,I473606,I325170,I325206,I473597,I473591,I325223,I325249,I325257,I325274,I325305,I473603,I325322,I325339,I325370,I325401,I325418,I325473,I565380,I325499,I325507,I325524,I565377,I565386,I325541,I565365,I325567,I565368,I325598,I325606,I565383,I325623,I325649,I325657,I565389,I325697,I325733,I565371,I565392,I325750,I565374,I325776,I325784,I325801,I325832,I325849,I325866,I325897,I325928,I325945,I326000,I326026,I326034,I326051,I326068,I326094,I326125,I326133,I326150,I326176,I326184,I326224,I326260,I326277,I326303,I326311,I326328,I326359,I326376,I326393,I326424,I326455,I326472,I326527,I326553,I326561,I326578,I326595,I326621,I326516,I326652,I326660,I326677,I326703,I326711,I326519,I326751,I326510,I326501,I326787,I326804,I326830,I326838,I326855,I326504,I326886,I326903,I326920,I326513,I326951,I326498,I326982,I326999,I326507,I327054,I327080,I327088,I327105,I327122,I327148,I327043,I327179,I327187,I327204,I327230,I327238,I327046,I327278,I327037,I327028,I327314,I327331,I327357,I327365,I327382,I327031,I327413,I327430,I327447,I327040,I327478,I327025,I327509,I327526,I327034,I327581,I563000,I327607,I327615,I327632,I562997,I563006,I327649,I562985,I327675,I562988,I327706,I327714,I563003,I327731,I327757,I327765,I563009,I327805,I327841,I562991,I563012,I327858,I562994,I327884,I327892,I327909,I327940,I327957,I327974,I328005,I328036,I328053,I328108,I385712,I328134,I328142,I328159,I385727,I385709,I328176,I328202,I385718,I328233,I328241,I385736,I328258,I328284,I328292,I385733,I328332,I328368,I385730,I385721,I328385,I385715,I328411,I328419,I328436,I328467,I385724,I328484,I328501,I328532,I328563,I328580,I328635,I547530,I328661,I328669,I328686,I547527,I547536,I328703,I547515,I328729,I547518,I328760,I328768,I547533,I328785,I328811,I328819,I547539,I328859,I328895,I547521,I547542,I328912,I547524,I328938,I328946,I328963,I328994,I329011,I329028,I329059,I329090,I329107,I329162,I329188,I329196,I329213,I329230,I329256,I329151,I329287,I329295,I329312,I329338,I329346,I329154,I329386,I329145,I329136,I329422,I329439,I329465,I329473,I329490,I329139,I329521,I329538,I329555,I329148,I329586,I329133,I329617,I329634,I329142,I329689,I329715,I329723,I329740,I329757,I329783,I329814,I329822,I329839,I329865,I329873,I329913,I329949,I329966,I329992,I330000,I330017,I330048,I330065,I330082,I330113,I330144,I330161,I330216,I427691,I330242,I330250,I330267,I427700,I427688,I330284,I427685,I330310,I330341,I330349,I427682,I330366,I330392,I330400,I330440,I330476,I427703,I427694,I330493,I427697,I330519,I330527,I330544,I330575,I330592,I330609,I330640,I330671,I330688,I330743,I330769,I330777,I330794,I330811,I330837,I330732,I330868,I330876,I330893,I330919,I330927,I330735,I330967,I330726,I330717,I331003,I331020,I331046,I331054,I331071,I330720,I331102,I331119,I331136,I330729,I331167,I330714,I331198,I331215,I330723,I331270,I331296,I331304,I331321,I331338,I331364,I331395,I331403,I331420,I331446,I331454,I331494,I331530,I331547,I331573,I331581,I331598,I331629,I331646,I331663,I331694,I331725,I331742,I331797,I573115,I331823,I331831,I331848,I573112,I573121,I331865,I573100,I331891,I573103,I331922,I331930,I573118,I331947,I331973,I331981,I573124,I332021,I332057,I573106,I573127,I332074,I573109,I332100,I332108,I332125,I332156,I332173,I332190,I332221,I332252,I332269,I332324,I332350,I332358,I332375,I332392,I332418,I332313,I332449,I332457,I332474,I332500,I332508,I332316,I332548,I332307,I332298,I332584,I332601,I332627,I332635,I332652,I332301,I332683,I332700,I332717,I332310,I332748,I332295,I332779,I332796,I332304,I332851,I332877,I332885,I332902,I332919,I332945,I332976,I332984,I333001,I333027,I333035,I333075,I333111,I333128,I333154,I333162,I333179,I333210,I333227,I333244,I333275,I333306,I333323,I333378,I480536,I333404,I333412,I333429,I480518,I333446,I480524,I333472,I480521,I333503,I333511,I480530,I333528,I333554,I333562,I480542,I333602,I333638,I480533,I480527,I333655,I333681,I333689,I333706,I333737,I480539,I333754,I333771,I333802,I333833,I333850,I333905,I546340,I333931,I333939,I333956,I546337,I546346,I333973,I546325,I333999,I546328,I334030,I334038,I546343,I334055,I334081,I334089,I546349,I334129,I334165,I546331,I546352,I334182,I546334,I334208,I334216,I334233,I334264,I334281,I334298,I334329,I334360,I334377,I334432,I379898,I334458,I334466,I334483,I379913,I379895,I334500,I334526,I379904,I334557,I334565,I379922,I334582,I334608,I334616,I379919,I334656,I334692,I379916,I379907,I334709,I379901,I334735,I334743,I334760,I334791,I379910,I334808,I334825,I334856,I334887,I334904,I334959,I334985,I334993,I335010,I335027,I335053,I335084,I335092,I335109,I335135,I335143,I335183,I335219,I335236,I335262,I335270,I335287,I335318,I335335,I335352,I335383,I335414,I335431,I335486,I408968,I335512,I335520,I335537,I408983,I408965,I335554,I335580,I408974,I335611,I335619,I408992,I335636,I335662,I335670,I408989,I335710,I335746,I408986,I408977,I335763,I408971,I335789,I335797,I335814,I335845,I408980,I335862,I335879,I335910,I335941,I335958,I336013,I336039,I336047,I336064,I336081,I336107,I336002,I336138,I336146,I336163,I336189,I336197,I336005,I336237,I335996,I335987,I336273,I336290,I336316,I336324,I336341,I335990,I336372,I336389,I336406,I335999,I336437,I335984,I336468,I336485,I335993,I336540,I336566,I336574,I336591,I336608,I336634,I336665,I336673,I336690,I336716,I336724,I336764,I336800,I336817,I336843,I336851,I336868,I336899,I336916,I336933,I336964,I336995,I337012,I337067,I525858,I337093,I337101,I337118,I525840,I525843,I337135,I525855,I337161,I337056,I525864,I337192,I337200,I525849,I337217,I337243,I337251,I337059,I525861,I337291,I337050,I337041,I337327,I525852,I525846,I337344,I337370,I337378,I337395,I337044,I337426,I337443,I337460,I337053,I337491,I337038,I337522,I337539,I337047,I337594,I337620,I337628,I337645,I337662,I337688,I337583,I337719,I337727,I337744,I337770,I337778,I337586,I337818,I337577,I337568,I337854,I337871,I337897,I337905,I337922,I337571,I337953,I337970,I337987,I337580,I338018,I337565,I338049,I338066,I337574,I338121,I490362,I338147,I338155,I338172,I490344,I338189,I490350,I338215,I490347,I338246,I338254,I490356,I338271,I338297,I338305,I490368,I338345,I338381,I490359,I490353,I338398,I338424,I338432,I338449,I338480,I490365,I338497,I338514,I338545,I338576,I338593,I338648,I388296,I338674,I338682,I338699,I388311,I388293,I338716,I338742,I388302,I338773,I338781,I388320,I338798,I338824,I338832,I388317,I338872,I338908,I388314,I388305,I338925,I388299,I338951,I338959,I338976,I339007,I388308,I339024,I339041,I339072,I339103,I339120,I339175,I339201,I339209,I339226,I339243,I339269,I339164,I339300,I339308,I339325,I339351,I339359,I339167,I339399,I339158,I339149,I339435,I339452,I339478,I339486,I339503,I339152,I339534,I339551,I339568,I339161,I339599,I339146,I339630,I339647,I339155,I339702,I339728,I339736,I339753,I339770,I339796,I339827,I339835,I339852,I339878,I339886,I339926,I339962,I339979,I340005,I340013,I340030,I340061,I340078,I340095,I340126,I340157,I340174,I340229,I471288,I340255,I340263,I340280,I471270,I340297,I471276,I340323,I471273,I340354,I340362,I471282,I340379,I340405,I340413,I471294,I340453,I340489,I471285,I471279,I340506,I340532,I340540,I340557,I340588,I471291,I340605,I340622,I340653,I340684,I340701,I340756,I419276,I340782,I340790,I340807,I419285,I419273,I340824,I419270,I340850,I340745,I340881,I340889,I419267,I340906,I340932,I340940,I340748,I340980,I340739,I340730,I341016,I419288,I419279,I341033,I419282,I341059,I341067,I341084,I340733,I341115,I341132,I341149,I340742,I341180,I340727,I341211,I341228,I340736,I341283,I341309,I341317,I341334,I341351,I341377,I341408,I341416,I341433,I341459,I341467,I341507,I341543,I341560,I341586,I341594,I341611,I341642,I341659,I341676,I341707,I341738,I341755,I341810,I436667,I341836,I341844,I341861,I436676,I436664,I341878,I436661,I341904,I341935,I341943,I436658,I341960,I341986,I341994,I342034,I342070,I436679,I436670,I342087,I436673,I342113,I342121,I342138,I342169,I342186,I342203,I342234,I342265,I342282,I342337,I342363,I342371,I342388,I342405,I342431,I342326,I342462,I342470,I342487,I342513,I342521,I342329,I342561,I342320,I342311,I342597,I342614,I342640,I342648,I342665,I342314,I342696,I342713,I342730,I342323,I342761,I342308,I342792,I342809,I342317,I342864,I342890,I342898,I342915,I342932,I342958,I342989,I342997,I343014,I343040,I343048,I343088,I343124,I343141,I343167,I343175,I343192,I343223,I343240,I343257,I343288,I343319,I343336,I343391,I343417,I343425,I343442,I343459,I343485,I343380,I343516,I343524,I343541,I343567,I343575,I343383,I343615,I343374,I343365,I343651,I343668,I343694,I343702,I343719,I343368,I343750,I343767,I343784,I343377,I343815,I343362,I343846,I343863,I343371,I343918,I343944,I343952,I343969,I343986,I344012,I344043,I344051,I344068,I344094,I344102,I344142,I344178,I344195,I344221,I344229,I344246,I344277,I344294,I344311,I344342,I344373,I344390,I344445,I344471,I344479,I344496,I344513,I344539,I344434,I344570,I344578,I344595,I344621,I344629,I344437,I344669,I344428,I344419,I344705,I344722,I344748,I344756,I344773,I344422,I344804,I344821,I344838,I344431,I344869,I344416,I344900,I344917,I344425,I344972,I344998,I345006,I345023,I345040,I345066,I344961,I345097,I345105,I345122,I345148,I345156,I344964,I345196,I344955,I344946,I345232,I345249,I345275,I345283,I345300,I344949,I345331,I345348,I345365,I344958,I345396,I344943,I345427,I345444,I344952,I345499,I345525,I345533,I345550,I345567,I345593,I345488,I345624,I345632,I345649,I345675,I345683,I345491,I345723,I345482,I345473,I345759,I345776,I345802,I345810,I345827,I345476,I345858,I345875,I345892,I345485,I345923,I345470,I345954,I345971,I345479,I346026,I466086,I346052,I346060,I346077,I466068,I346094,I466074,I346120,I346015,I466071,I346151,I346159,I466080,I346176,I346202,I346210,I346018,I466092,I346250,I346009,I346000,I346286,I466083,I466077,I346303,I346329,I346337,I346354,I346003,I346385,I466089,I346402,I346419,I346012,I346450,I345997,I346481,I346498,I346006,I346553,I346579,I346587,I346604,I346621,I346647,I346678,I346686,I346703,I346729,I346737,I346777,I346813,I346830,I346856,I346864,I346881,I346912,I346929,I346946,I346977,I347008,I347025,I347080,I543365,I347106,I347114,I347131,I543362,I543371,I347148,I543350,I347174,I543353,I347205,I347213,I543368,I347230,I347256,I347264,I543374,I347304,I347340,I543356,I543377,I347357,I543359,I347383,I347391,I347408,I347439,I347456,I347473,I347504,I347535,I347552,I347607,I475912,I347633,I347641,I347658,I475894,I347675,I475900,I347701,I347596,I475897,I347732,I347740,I475906,I347757,I347783,I347791,I347599,I475918,I347831,I347590,I347581,I347867,I475909,I475903,I347884,I347910,I347918,I347935,I347584,I347966,I475915,I347983,I348000,I347593,I348031,I347578,I348062,I348079,I347587,I348134,I348160,I348168,I348185,I348202,I348228,I348259,I348267,I348284,I348310,I348318,I348358,I348394,I348411,I348437,I348445,I348462,I348493,I348510,I348527,I348558,I348589,I348606,I348661,I460884,I348687,I348695,I348712,I460866,I348729,I460872,I348755,I460869,I348786,I348794,I460878,I348811,I348837,I348845,I460890,I348885,I348921,I460881,I460875,I348938,I348964,I348972,I348989,I349020,I460887,I349037,I349054,I349085,I349116,I349133,I349188,I470132,I349214,I349222,I349239,I470114,I349256,I470120,I349282,I349177,I470117,I349313,I349321,I470126,I349338,I349364,I349372,I349180,I470138,I349412,I349171,I349162,I349448,I470129,I470123,I349465,I349491,I349499,I349516,I349165,I349547,I470135,I349564,I349581,I349174,I349612,I349159,I349643,I349660,I349168,I349715,I349741,I349749,I349766,I349783,I349809,I349840,I349848,I349865,I349891,I349899,I349939,I349975,I349992,I350018,I350026,I350043,I350074,I350091,I350108,I350139,I350170,I350187,I350242,I380544,I350268,I350276,I350293,I380559,I380541,I350310,I350336,I380550,I350367,I350375,I380568,I350392,I350418,I350426,I380565,I350466,I350502,I380562,I380553,I350519,I380547,I350545,I350553,I350570,I350601,I380556,I350618,I350635,I350666,I350697,I350714,I350769,I350795,I350803,I350820,I350837,I350863,I350894,I350902,I350919,I350945,I350953,I350993,I351029,I351046,I351072,I351080,I351097,I351128,I351145,I351162,I351193,I351224,I351241,I351296,I351322,I351330,I351347,I351364,I351390,I351421,I351429,I351446,I351472,I351480,I351520,I351556,I351573,I351599,I351607,I351624,I351655,I351672,I351689,I351720,I351751,I351768,I351823,I351849,I351857,I351874,I351891,I351917,I351948,I351956,I351973,I351999,I352007,I352047,I352083,I352100,I352126,I352134,I352151,I352182,I352199,I352216,I352247,I352278,I352295,I352350,I352376,I352384,I352401,I352418,I352444,I352475,I352483,I352500,I352526,I352534,I352574,I352610,I352627,I352653,I352661,I352678,I352709,I352726,I352743,I352774,I352805,I352822,I352877,I538010,I352903,I352911,I352928,I538007,I538016,I352945,I537995,I352971,I537998,I353002,I353010,I538013,I353027,I353053,I353061,I538019,I353101,I353137,I538001,I538022,I353154,I538004,I353180,I353188,I353205,I353236,I353253,I353270,I353301,I353332,I353349,I353404,I353430,I353438,I353455,I353472,I353498,I353529,I353537,I353554,I353580,I353588,I353628,I353664,I353681,I353707,I353715,I353732,I353763,I353780,I353797,I353828,I353859,I353876,I353931,I353957,I353965,I353982,I353999,I354025,I354056,I354064,I354081,I354107,I354115,I354155,I354191,I354208,I354234,I354242,I354259,I354290,I354307,I354324,I354355,I354386,I354403,I354458,I354484,I354492,I354509,I354526,I354552,I354583,I354591,I354608,I354634,I354642,I354682,I354718,I354735,I354761,I354769,I354786,I354817,I354834,I354851,I354882,I354913,I354930,I354985,I355011,I355019,I355036,I355053,I355079,I354974,I355110,I355118,I355135,I355161,I355169,I354977,I355209,I354968,I354959,I355245,I355262,I355288,I355296,I355313,I354962,I355344,I355361,I355378,I354971,I355409,I354956,I355440,I355457,I354965,I355512,I355538,I355546,I355563,I355580,I355606,I355501,I355637,I355645,I355662,I355688,I355696,I355504,I355736,I355495,I355486,I355772,I355789,I355815,I355823,I355840,I355489,I355871,I355888,I355905,I355498,I355936,I355483,I355967,I355984,I355492,I356039,I356065,I356073,I356090,I356107,I356133,I356164,I356172,I356189,I356215,I356223,I356263,I356299,I356316,I356342,I356350,I356367,I356398,I356415,I356432,I356463,I356494,I356511,I356566,I544555,I356592,I356600,I356617,I544552,I544561,I356634,I544540,I356660,I356555,I544543,I356691,I356699,I544558,I356716,I356742,I356750,I356558,I544564,I356790,I356549,I356540,I356826,I544546,I544567,I356843,I544549,I356869,I356877,I356894,I356543,I356925,I356942,I356959,I356552,I356990,I356537,I357021,I357038,I356546,I357093,I357119,I357127,I357144,I357161,I357187,I357218,I357226,I357243,I357269,I357277,I357317,I357353,I357370,I357396,I357404,I357421,I357452,I357469,I357486,I357517,I357548,I357565,I357620,I357646,I357654,I357671,I357688,I357714,I357745,I357753,I357770,I357796,I357804,I357844,I357880,I357897,I357923,I357931,I357948,I357979,I357996,I358013,I358044,I358075,I358092,I358147,I358173,I358181,I358198,I358215,I358241,I358136,I358272,I358280,I358297,I358323,I358331,I358139,I358371,I358130,I358121,I358407,I358424,I358450,I358458,I358475,I358124,I358506,I358523,I358540,I358133,I358571,I358118,I358602,I358619,I358127,I358674,I474178,I358700,I358708,I358725,I474160,I358742,I474166,I358768,I474163,I358799,I358807,I474172,I358824,I358850,I358858,I474184,I358898,I358934,I474175,I474169,I358951,I358977,I358985,I359002,I359033,I474181,I359050,I359067,I359098,I359129,I359146,I359201,I457416,I359227,I359235,I359252,I457398,I359269,I457404,I359295,I457401,I359326,I359334,I457410,I359351,I359377,I359385,I457422,I359425,I359461,I457413,I457407,I359478,I359504,I359512,I359529,I359560,I457419,I359577,I359594,I359625,I359656,I359673,I359728,I359754,I359762,I359779,I359796,I359822,I359717,I359853,I359861,I359878,I359904,I359912,I359720,I359952,I359711,I359702,I359988,I360005,I360031,I360039,I360056,I359705,I360087,I360104,I360121,I359714,I360152,I359699,I360183,I360200,I359708,I360255,I381190,I360281,I360289,I360306,I381205,I381187,I360323,I360349,I381196,I360380,I360388,I381214,I360405,I360431,I360439,I381211,I360479,I360515,I381208,I381199,I360532,I381193,I360558,I360566,I360583,I360614,I381202,I360631,I360648,I360679,I360710,I360727,I360782,I503582,I360808,I360816,I360833,I503588,I503570,I360850,I503579,I360876,I503585,I360907,I360915,I503573,I360932,I360958,I360966,I503591,I361006,I361042,I503576,I361059,I503594,I361085,I361093,I361110,I361141,I361158,I361175,I361206,I361237,I361254,I361309,I361335,I361343,I361360,I361377,I361403,I361298,I361434,I361442,I361459,I361485,I361493,I361301,I361533,I361292,I361283,I361569,I361586,I361612,I361620,I361637,I361286,I361668,I361685,I361702,I361295,I361733,I361280,I361764,I361781,I361289,I361842,I361868,I361885,I361893,I361910,I361927,I361944,I361961,I361978,I362009,I362026,I362057,I362074,I362091,I362122,I362162,I362170,I362187,I362204,I362221,I362252,I362269,I362286,I362312,I362334,I362351,I362382,I362427,I362488,I362514,I362531,I362539,I362556,I362573,I362590,I362607,I362624,I362655,I362672,I362703,I362720,I362737,I362768,I362808,I362816,I362833,I362850,I362867,I362898,I362915,I362932,I362958,I362980,I362997,I363028,I363073,I363134,I467820,I363160,I467802,I363177,I363185,I363202,I467811,I363219,I467823,I363236,I467805,I363253,I467814,I363270,I363301,I363318,I363349,I363366,I467826,I363383,I363414,I363454,I363462,I363479,I363496,I363513,I363544,I467808,I363561,I467817,I363578,I363604,I363626,I363643,I363674,I363719,I363780,I363806,I363823,I363831,I363848,I363865,I363882,I363899,I363916,I363947,I363964,I363995,I364012,I364029,I364060,I364100,I364108,I364125,I364142,I364159,I364190,I364207,I364224,I364250,I364272,I364289,I364320,I364365,I364426,I364452,I364469,I364477,I364494,I364511,I364528,I364545,I364562,I364593,I364610,I364641,I364658,I364675,I364706,I364746,I364754,I364771,I364788,I364805,I364836,I364853,I364870,I364896,I364918,I364935,I364966,I365011,I365072,I365098,I365115,I365123,I365140,I365157,I365174,I365191,I365208,I365239,I365256,I365287,I365304,I365321,I365352,I365392,I365400,I365417,I365434,I365451,I365482,I365499,I365516,I365542,I365564,I365581,I365612,I365657,I365718,I365744,I365761,I365769,I365786,I365803,I365820,I365837,I365854,I365704,I365885,I365902,I365707,I365933,I365950,I365967,I365683,I365998,I365695,I366038,I366046,I366063,I366080,I366097,I365710,I366128,I366145,I366162,I366188,I365698,I366210,I366227,I365692,I366258,I365686,I365689,I366303,I365701,I366364,I366390,I366407,I366415,I366432,I366449,I366466,I366483,I366500,I366531,I366548,I366579,I366596,I366613,I366644,I366684,I366692,I366709,I366726,I366743,I366774,I366791,I366808,I366834,I366856,I366873,I366904,I366949,I367010,I367036,I367053,I367061,I367078,I367095,I367112,I367129,I367146,I367177,I367194,I367225,I367242,I367259,I367290,I367330,I367338,I367355,I367372,I367389,I367420,I367437,I367454,I367480,I367502,I367519,I367550,I367595,I367656,I367682,I367699,I367707,I367724,I367741,I367758,I367775,I367792,I367823,I367840,I367871,I367888,I367905,I367936,I367976,I367984,I368001,I368018,I368035,I368066,I368083,I368100,I368126,I368148,I368165,I368196,I368241,I368302,I368328,I368345,I368353,I368370,I368387,I368404,I368421,I368438,I368469,I368486,I368517,I368534,I368551,I368582,I368622,I368630,I368647,I368664,I368681,I368712,I368729,I368746,I368772,I368794,I368811,I368842,I368887,I368948,I453948,I368974,I453930,I368991,I368999,I369016,I453939,I369033,I453951,I369050,I453933,I369067,I453942,I369084,I369115,I369132,I369163,I369180,I453954,I369197,I369228,I369268,I369276,I369293,I369310,I369327,I369358,I453936,I369375,I453945,I369392,I369418,I369440,I369457,I369488,I369533,I369594,I369620,I369637,I369645,I369662,I369679,I369696,I369713,I369730,I369761,I369778,I369809,I369826,I369843,I369874,I369914,I369922,I369939,I369956,I369973,I370004,I370021,I370038,I370064,I370086,I370103,I370134,I370179,I370240,I370266,I370283,I370291,I370308,I370325,I370342,I370359,I370376,I370226,I370407,I370424,I370229,I370455,I370472,I370489,I370205,I370520,I370217,I370560,I370568,I370585,I370602,I370619,I370232,I370650,I370667,I370684,I370710,I370220,I370732,I370749,I370214,I370780,I370208,I370211,I370825,I370223,I370886,I462618,I370912,I462600,I370929,I370937,I370954,I462609,I370971,I462621,I370988,I462603,I371005,I462612,I371022,I370872,I371053,I371070,I370875,I371101,I371118,I462624,I371135,I370851,I371166,I370863,I371206,I371214,I371231,I371248,I371265,I370878,I371296,I462606,I371313,I462615,I371330,I371356,I370866,I371378,I371395,I370860,I371426,I370854,I370857,I371471,I370869,I371532,I371558,I371575,I371583,I371600,I371617,I371634,I371651,I371668,I371518,I371699,I371716,I371521,I371747,I371764,I371781,I371497,I371812,I371509,I371852,I371860,I371877,I371894,I371911,I371524,I371942,I371959,I371976,I372002,I371512,I372024,I372041,I371506,I372072,I371500,I371503,I372117,I371515,I372178,I372204,I372221,I372229,I372246,I372263,I372280,I372297,I372314,I372164,I372345,I372362,I372167,I372393,I372410,I372427,I372143,I372458,I372155,I372498,I372506,I372523,I372540,I372557,I372170,I372588,I372605,I372622,I372648,I372158,I372670,I372687,I372152,I372718,I372146,I372149,I372763,I372161,I372824,I372850,I372867,I372875,I372892,I372909,I372926,I372943,I372960,I372991,I373008,I373039,I373056,I373073,I373104,I373144,I373152,I373169,I373186,I373203,I373234,I373251,I373268,I373294,I373316,I373333,I373364,I373409,I373470,I373496,I373513,I373521,I373538,I373555,I373572,I373589,I373606,I373637,I373654,I373685,I373702,I373719,I373750,I373790,I373798,I373815,I373832,I373849,I373880,I373897,I373914,I373940,I373962,I373979,I374010,I374055,I374116,I374142,I374159,I374167,I374184,I374201,I374218,I374235,I374252,I374283,I374300,I374331,I374348,I374365,I374396,I374436,I374444,I374461,I374478,I374495,I374526,I374543,I374560,I374586,I374608,I374625,I374656,I374701,I374762,I374788,I374805,I374813,I374830,I374847,I374864,I374881,I374898,I374929,I374946,I374977,I374994,I375011,I375042,I375082,I375090,I375107,I375124,I375141,I375172,I375189,I375206,I375232,I375254,I375271,I375302,I375347,I375408,I375434,I375451,I375459,I375476,I375493,I375510,I375527,I375544,I375575,I375592,I375623,I375640,I375657,I375688,I375728,I375736,I375753,I375770,I375787,I375818,I375835,I375852,I375878,I375900,I375917,I375948,I375993,I376054,I376080,I376097,I376105,I376122,I376139,I376156,I376173,I376190,I376221,I376238,I376269,I376286,I376303,I376334,I376374,I376382,I376399,I376416,I376433,I376464,I376481,I376498,I376524,I376546,I376563,I376594,I376639,I376700,I515556,I376726,I515562,I376743,I376751,I376768,I515559,I376785,I515538,I376802,I515541,I376819,I515547,I376836,I376867,I376884,I376915,I376932,I376949,I376980,I377020,I377028,I377045,I377062,I515550,I377079,I377110,I377127,I515544,I377144,I515553,I377170,I377192,I377209,I377240,I377285,I377346,I377372,I377389,I377397,I377414,I377431,I377448,I377465,I377482,I377513,I377530,I377561,I377578,I377595,I377626,I377666,I377674,I377691,I377708,I377725,I377756,I377773,I377790,I377816,I377838,I377855,I377886,I377931,I377992,I378018,I378035,I378043,I378060,I378077,I378094,I378111,I378128,I378159,I378176,I378207,I378224,I378241,I378272,I378312,I378320,I378337,I378354,I378371,I378402,I378419,I378436,I378462,I378484,I378501,I378532,I378577,I378638,I378664,I378681,I378689,I378706,I378723,I378740,I378757,I378774,I378624,I378805,I378822,I378627,I378853,I378870,I378887,I378603,I378918,I378615,I378958,I378966,I378983,I379000,I379017,I378630,I379048,I379065,I379082,I379108,I378618,I379130,I379147,I378612,I379178,I378606,I378609,I379223,I378621,I379284,I379310,I379327,I379335,I379352,I379369,I379386,I379403,I379420,I379451,I379468,I379499,I379516,I379533,I379564,I379604,I379612,I379629,I379646,I379663,I379694,I379711,I379728,I379754,I379776,I379793,I379824,I379869,I379930,I379956,I379973,I379981,I379998,I380015,I380032,I380049,I380066,I380097,I380114,I380145,I380162,I380179,I380210,I380250,I380258,I380275,I380292,I380309,I380340,I380357,I380374,I380400,I380422,I380439,I380470,I380515,I380576,I380602,I380619,I380627,I380644,I380661,I380678,I380695,I380712,I380743,I380760,I380791,I380808,I380825,I380856,I380896,I380904,I380921,I380938,I380955,I380986,I381003,I381020,I381046,I381068,I381085,I381116,I381161,I381222,I381248,I381265,I381273,I381290,I381307,I381324,I381341,I381358,I381389,I381406,I381437,I381454,I381471,I381502,I381542,I381550,I381567,I381584,I381601,I381632,I381649,I381666,I381692,I381714,I381731,I381762,I381807,I381868,I381894,I381911,I381919,I381936,I381953,I381970,I381987,I382004,I382035,I382052,I382083,I382100,I382117,I382148,I382188,I382196,I382213,I382230,I382247,I382278,I382295,I382312,I382338,I382360,I382377,I382408,I382453,I382514,I382540,I382557,I382565,I382582,I382599,I382616,I382633,I382650,I382681,I382698,I382729,I382746,I382763,I382794,I382834,I382842,I382859,I382876,I382893,I382924,I382941,I382958,I382984,I383006,I383023,I383054,I383099,I383160,I383186,I383203,I383211,I383228,I383245,I383262,I383279,I383296,I383327,I383344,I383375,I383392,I383409,I383440,I383480,I383488,I383505,I383522,I383539,I383570,I383587,I383604,I383630,I383652,I383669,I383700,I383745,I383806,I383832,I383849,I383857,I383874,I383891,I383908,I383925,I383942,I383973,I383990,I384021,I384038,I384055,I384086,I384126,I384134,I384151,I384168,I384185,I384216,I384233,I384250,I384276,I384298,I384315,I384346,I384391,I384452,I440654,I384478,I440636,I384495,I384503,I384520,I440645,I384537,I440657,I384554,I440639,I384571,I440648,I384588,I384619,I384636,I384667,I384684,I440660,I384701,I384732,I384772,I384780,I384797,I384814,I384831,I384862,I440642,I384879,I440651,I384896,I384922,I384944,I384961,I384992,I385037,I385098,I463774,I385124,I463756,I385141,I385149,I385166,I463765,I385183,I463777,I385200,I463759,I385217,I463768,I385234,I385084,I385265,I385282,I385087,I385313,I385330,I463780,I385347,I385063,I385378,I385075,I385418,I385426,I385443,I385460,I385477,I385090,I385508,I463762,I385525,I463771,I385542,I385568,I385078,I385590,I385607,I385072,I385638,I385066,I385069,I385683,I385081,I385744,I385770,I385787,I385795,I385812,I385829,I385846,I385863,I385880,I385911,I385928,I385959,I385976,I385993,I386024,I386064,I386072,I386089,I386106,I386123,I386154,I386171,I386188,I386214,I386236,I386253,I386284,I386329,I386390,I484582,I386416,I484564,I386433,I386441,I386458,I484573,I386475,I484585,I386492,I484567,I386509,I484576,I386526,I386557,I386574,I386605,I386622,I484588,I386639,I386670,I386710,I386718,I386735,I386752,I386769,I386800,I484570,I386817,I484579,I386834,I386860,I386882,I386899,I386930,I386975,I387036,I387062,I387079,I387087,I387104,I387121,I387138,I387155,I387172,I387203,I387220,I387251,I387268,I387285,I387316,I387356,I387364,I387381,I387398,I387415,I387446,I387463,I387480,I387506,I387528,I387545,I387576,I387621,I387682,I387708,I387725,I387733,I387750,I387767,I387784,I387801,I387818,I387849,I387866,I387897,I387914,I387931,I387962,I388002,I388010,I388027,I388044,I388061,I388092,I388109,I388126,I388152,I388174,I388191,I388222,I388267,I388328,I489206,I388354,I489188,I388371,I388379,I388396,I489197,I388413,I489209,I388430,I489191,I388447,I489200,I388464,I388495,I388512,I388543,I388560,I489212,I388577,I388608,I388648,I388656,I388673,I388690,I388707,I388738,I489194,I388755,I489203,I388772,I388798,I388820,I388837,I388868,I388913,I388974,I389000,I389017,I389025,I389042,I389059,I389076,I389093,I389110,I389141,I389158,I389189,I389206,I389223,I389254,I389294,I389302,I389319,I389336,I389353,I389384,I389401,I389418,I389444,I389466,I389483,I389514,I389559,I389620,I554060,I389646,I554084,I389663,I389671,I389688,I554066,I389705,I554075,I389722,I389739,I554081,I389756,I389787,I389804,I389835,I389852,I554078,I389869,I389900,I389940,I389948,I389965,I389982,I554072,I389999,I390030,I554063,I390047,I554087,I390064,I554069,I390090,I390112,I390129,I390160,I390205,I390266,I390292,I390309,I390317,I390334,I390351,I390368,I390385,I390402,I390433,I390450,I390481,I390498,I390515,I390546,I390586,I390594,I390611,I390628,I390645,I390676,I390693,I390710,I390736,I390758,I390775,I390806,I390851,I390912,I504676,I390938,I504682,I390955,I390963,I390980,I504679,I390997,I504658,I391014,I504661,I391031,I504667,I391048,I391079,I391096,I391127,I391144,I391161,I391192,I391232,I391240,I391257,I391274,I504670,I391291,I391322,I391339,I504664,I391356,I504673,I391382,I391404,I391421,I391452,I391497,I391558,I391584,I391601,I391609,I391626,I391643,I391660,I391677,I391694,I391725,I391742,I391773,I391790,I391807,I391838,I391878,I391886,I391903,I391920,I391937,I391968,I391985,I392002,I392028,I392050,I392067,I392098,I392143,I392204,I392230,I392247,I392255,I392272,I392289,I392306,I392323,I392340,I392371,I392388,I392419,I392436,I392453,I392484,I392524,I392532,I392549,I392566,I392583,I392614,I392631,I392648,I392674,I392696,I392713,I392744,I392789,I392850,I392876,I392893,I392901,I392918,I392935,I392952,I392969,I392986,I393017,I393034,I393065,I393082,I393099,I393130,I393170,I393178,I393195,I393212,I393229,I393260,I393277,I393294,I393320,I393342,I393359,I393390,I393435,I393496,I393522,I393539,I393547,I393564,I393581,I393598,I393615,I393632,I393482,I393663,I393680,I393485,I393711,I393728,I393745,I393461,I393776,I393473,I393816,I393824,I393841,I393858,I393875,I393488,I393906,I393923,I393940,I393966,I393476,I393988,I394005,I393470,I394036,I393464,I393467,I394081,I393479,I394142,I394168,I394185,I394193,I394210,I394227,I394244,I394261,I394278,I394309,I394326,I394357,I394374,I394391,I394422,I394462,I394470,I394487,I394504,I394521,I394552,I394569,I394586,I394612,I394634,I394651,I394682,I394727,I394788,I394814,I394831,I394839,I394856,I394873,I394890,I394907,I394924,I394774,I394955,I394972,I394777,I395003,I395020,I395037,I394753,I395068,I394765,I395108,I395116,I395133,I395150,I395167,I394780,I395198,I395215,I395232,I395258,I394768,I395280,I395297,I394762,I395328,I394756,I394759,I395373,I394771,I395434,I395460,I395477,I395485,I395502,I395519,I395536,I395553,I395570,I395601,I395618,I395649,I395666,I395683,I395714,I395754,I395762,I395779,I395796,I395813,I395844,I395861,I395878,I395904,I395926,I395943,I395974,I396019,I396080,I396106,I396123,I396131,I396148,I396165,I396182,I396199,I396216,I396247,I396264,I396295,I396312,I396329,I396360,I396400,I396408,I396425,I396442,I396459,I396490,I396507,I396524,I396550,I396572,I396589,I396620,I396665,I396726,I396752,I396769,I396777,I396794,I396811,I396828,I396845,I396862,I396893,I396910,I396941,I396958,I396975,I397006,I397046,I397054,I397071,I397088,I397105,I397136,I397153,I397170,I397196,I397218,I397235,I397266,I397311,I397372,I397398,I397415,I397423,I397440,I397457,I397474,I397491,I397508,I397539,I397556,I397587,I397604,I397621,I397652,I397692,I397700,I397717,I397734,I397751,I397782,I397799,I397816,I397842,I397864,I397881,I397912,I397957,I398018,I398044,I398061,I398069,I398086,I398103,I398120,I398137,I398154,I398185,I398202,I398233,I398250,I398267,I398298,I398338,I398346,I398363,I398380,I398397,I398428,I398445,I398462,I398488,I398510,I398527,I398558,I398603,I398664,I398690,I398707,I398715,I398732,I398749,I398766,I398783,I398800,I398831,I398848,I398879,I398896,I398913,I398944,I398984,I398992,I399009,I399026,I399043,I399074,I399091,I399108,I399134,I399156,I399173,I399204,I399249,I399310,I399336,I399353,I399361,I399378,I399395,I399412,I399429,I399446,I399296,I399477,I399494,I399299,I399525,I399542,I399559,I399275,I399590,I399287,I399630,I399638,I399655,I399672,I399689,I399302,I399720,I399737,I399754,I399780,I399290,I399802,I399819,I399284,I399850,I399278,I399281,I399895,I399293,I399956,I399982,I399999,I400007,I400024,I400041,I400058,I400075,I400092,I399942,I400123,I400140,I399945,I400171,I400188,I400205,I399921,I400236,I399933,I400276,I400284,I400301,I400318,I400335,I399948,I400366,I400383,I400400,I400426,I399936,I400448,I400465,I399930,I400496,I399924,I399927,I400541,I399939,I400602,I400628,I400645,I400653,I400670,I400687,I400704,I400721,I400738,I400588,I400769,I400786,I400591,I400817,I400834,I400851,I400567,I400882,I400579,I400922,I400930,I400947,I400964,I400981,I400594,I401012,I401029,I401046,I401072,I400582,I401094,I401111,I400576,I401142,I400570,I400573,I401187,I400585,I401248,I401274,I401291,I401299,I401316,I401333,I401350,I401367,I401384,I401234,I401415,I401432,I401237,I401463,I401480,I401497,I401213,I401528,I401225,I401568,I401576,I401593,I401610,I401627,I401240,I401658,I401675,I401692,I401718,I401228,I401740,I401757,I401222,I401788,I401216,I401219,I401833,I401231,I401894,I455682,I401920,I455664,I401937,I401945,I401962,I455673,I401979,I455685,I401996,I455667,I402013,I455676,I402030,I402061,I402078,I402109,I402126,I455688,I402143,I402174,I402214,I402222,I402239,I402256,I402273,I402304,I455670,I402321,I455679,I402338,I402364,I402386,I402403,I402434,I402479,I402540,I402566,I402583,I402591,I402608,I402625,I402642,I402659,I402676,I402526,I402707,I402724,I402529,I402755,I402772,I402789,I402505,I402820,I402517,I402860,I402868,I402885,I402902,I402919,I402532,I402950,I402967,I402984,I403010,I402520,I403032,I403049,I402514,I403080,I402508,I402511,I403125,I402523,I403186,I403212,I403229,I403237,I403254,I403271,I403288,I403305,I403322,I403353,I403370,I403401,I403418,I403435,I403466,I403506,I403514,I403531,I403548,I403565,I403596,I403613,I403630,I403656,I403678,I403695,I403726,I403771,I403832,I403858,I403875,I403883,I403900,I403917,I403934,I403951,I403968,I403818,I403999,I404016,I403821,I404047,I404064,I404081,I403797,I404112,I403809,I404152,I404160,I404177,I404194,I404211,I403824,I404242,I404259,I404276,I404302,I403812,I404324,I404341,I403806,I404372,I403800,I403803,I404417,I403815,I404478,I488628,I404504,I488610,I404521,I404529,I404546,I488619,I404563,I488631,I404580,I488613,I404597,I488622,I404614,I404645,I404662,I404693,I404710,I488634,I404727,I404758,I404798,I404806,I404823,I404840,I404857,I404888,I488616,I404905,I488625,I404922,I404948,I404970,I404987,I405018,I405063,I405124,I405150,I405167,I405175,I405192,I405209,I405226,I405243,I405260,I405291,I405308,I405339,I405356,I405373,I405404,I405444,I405452,I405469,I405486,I405503,I405534,I405551,I405568,I405594,I405616,I405633,I405664,I405709,I405770,I405796,I405813,I405821,I405838,I405855,I405872,I405889,I405906,I405756,I405937,I405954,I405759,I405985,I406002,I406019,I405735,I406050,I405747,I406090,I406098,I406115,I406132,I406149,I405762,I406180,I406197,I406214,I406240,I405750,I406262,I406279,I405744,I406310,I405738,I405741,I406355,I405753,I406416,I406442,I406459,I406467,I406484,I406501,I406518,I406535,I406552,I406583,I406600,I406631,I406648,I406665,I406696,I406736,I406744,I406761,I406778,I406795,I406826,I406843,I406860,I406886,I406908,I406925,I406956,I407001,I407062,I407088,I407105,I407113,I407130,I407147,I407164,I407181,I407198,I407229,I407246,I407277,I407294,I407311,I407342,I407382,I407390,I407407,I407424,I407441,I407472,I407489,I407506,I407532,I407554,I407571,I407602,I407647,I407708,I407734,I407751,I407759,I407776,I407793,I407810,I407827,I407844,I407694,I407875,I407892,I407697,I407923,I407940,I407957,I407673,I407988,I407685,I408028,I408036,I408053,I408070,I408087,I407700,I408118,I408135,I408152,I408178,I407688,I408200,I408217,I407682,I408248,I407676,I407679,I408293,I407691,I408354,I408380,I408397,I408405,I408422,I408439,I408456,I408473,I408490,I408521,I408538,I408569,I408586,I408603,I408634,I408674,I408682,I408699,I408716,I408733,I408764,I408781,I408798,I408824,I408846,I408863,I408894,I408939,I409000,I438920,I409026,I438902,I409043,I409051,I409068,I438911,I409085,I438923,I409102,I438905,I409119,I438914,I409136,I409167,I409184,I409215,I409232,I438926,I409249,I409280,I409320,I409328,I409345,I409362,I409379,I409410,I438908,I409427,I438917,I409444,I409470,I409492,I409509,I409540,I409585,I409646,I409672,I409689,I409697,I409714,I409731,I409748,I409765,I409782,I409632,I409813,I409830,I409635,I409861,I409878,I409895,I409611,I409926,I409623,I409966,I409974,I409991,I410008,I410025,I409638,I410056,I410073,I410090,I410116,I409626,I410138,I410155,I409620,I410186,I409614,I409617,I410231,I409629,I410292,I418145,I410318,I418148,I410335,I410343,I410360,I410377,I418157,I410394,I418166,I410411,I418154,I410428,I410459,I410476,I410507,I410524,I418160,I410541,I410572,I410612,I410620,I410637,I410654,I418151,I410671,I410702,I418163,I410719,I410736,I410762,I410784,I410801,I410832,I410877,I410938,I410964,I410981,I410989,I411006,I411023,I411040,I411057,I411074,I411105,I411122,I411153,I411170,I411187,I411218,I411258,I411266,I411283,I411300,I411317,I411348,I411365,I411382,I411408,I411430,I411447,I411478,I411523,I411584,I518335,I411610,I518329,I411627,I411635,I411652,I518338,I411669,I518350,I411686,I518332,I411703,I411720,I411751,I411768,I411799,I411816,I518326,I411833,I411864,I411904,I411912,I411929,I411946,I518347,I411963,I411994,I518341,I412011,I412028,I518344,I412054,I412076,I412093,I412124,I412169,I412230,I412256,I412273,I412281,I412298,I412315,I412332,I412349,I412366,I412397,I412414,I412445,I412462,I412479,I412510,I412550,I412558,I412575,I412592,I412609,I412640,I412657,I412674,I412700,I412722,I412739,I412770,I412815,I412876,I412902,I412919,I412927,I412944,I412961,I412978,I412995,I413012,I413043,I413060,I413091,I413108,I413125,I413156,I413196,I413204,I413221,I413238,I413255,I413286,I413303,I413320,I413346,I413368,I413385,I413416,I413461,I413522,I413548,I413565,I413573,I413590,I413607,I413624,I413641,I413658,I413689,I413706,I413737,I413754,I413771,I413802,I413842,I413850,I413867,I413884,I413901,I413932,I413949,I413966,I413992,I414014,I414031,I414062,I414107,I414168,I414194,I414211,I414219,I414236,I414253,I414270,I414287,I414304,I414154,I414335,I414352,I414157,I414383,I414400,I414417,I414133,I414448,I414145,I414488,I414496,I414513,I414530,I414547,I414160,I414578,I414595,I414612,I414638,I414148,I414660,I414677,I414142,I414708,I414136,I414139,I414753,I414151,I414808,I414834,I414851,I414873,I414899,I414907,I414924,I414941,I414958,I414975,I414992,I415009,I415040,I415071,I415088,I415105,I415122,I415153,I415198,I415215,I415232,I415258,I415266,I415297,I415314,I415369,I415395,I415412,I415434,I415460,I415468,I415485,I415502,I415519,I415536,I415553,I415570,I415601,I415632,I415649,I415666,I415683,I415714,I415759,I415776,I415793,I415819,I415827,I415858,I415875,I415930,I415956,I415973,I415995,I416021,I416029,I416046,I416063,I416080,I416097,I416114,I416131,I416162,I416193,I416210,I416227,I416244,I416275,I416320,I416337,I416354,I416380,I416388,I416419,I416436,I416491,I416517,I416534,I416483,I416556,I416582,I416590,I416607,I416624,I416641,I416658,I416675,I416692,I416465,I416723,I416468,I416754,I416771,I416788,I416805,I416477,I416836,I416480,I416474,I416881,I416898,I416915,I416941,I416949,I416462,I416980,I416997,I416471,I417052,I417078,I417095,I417044,I417117,I417143,I417151,I417168,I417185,I417202,I417219,I417236,I417253,I417026,I417284,I417029,I417315,I417332,I417349,I417366,I417038,I417397,I417041,I417035,I417442,I417459,I417476,I417502,I417510,I417023,I417541,I417558,I417032,I417613,I560620,I417639,I417656,I417678,I560614,I417704,I417712,I560605,I417729,I417746,I560632,I417763,I560617,I560626,I417780,I417797,I560611,I417814,I417845,I417876,I560629,I417893,I417910,I417927,I417958,I418003,I560623,I418020,I418037,I560608,I418063,I418071,I418102,I418119,I418174,I418200,I418217,I418239,I418265,I418273,I418290,I418307,I418324,I418341,I418358,I418375,I418406,I418437,I418454,I418471,I418488,I418519,I418564,I418581,I418598,I418624,I418632,I418663,I418680,I418735,I418761,I418778,I418800,I418826,I418834,I418851,I418868,I418885,I418902,I418919,I418936,I418967,I418998,I419015,I419032,I419049,I419080,I419125,I419142,I419159,I419185,I419193,I419224,I419241,I419296,I419322,I419339,I419361,I419387,I419395,I419412,I419429,I419446,I419463,I419480,I419497,I419528,I419559,I419576,I419593,I419610,I419641,I419686,I419703,I419720,I419746,I419754,I419785,I419802,I419857,I459147,I419883,I419900,I419922,I459138,I419948,I419956,I459135,I419973,I419990,I459144,I420007,I459153,I420024,I420041,I459132,I420058,I420089,I420120,I459141,I420137,I420154,I420171,I420202,I420247,I459156,I420264,I420281,I459150,I420307,I420315,I420346,I420363,I420418,I420444,I420461,I420483,I420509,I420517,I420534,I420551,I420568,I420585,I420602,I420619,I420650,I420681,I420698,I420715,I420732,I420763,I420808,I420825,I420842,I420868,I420876,I420907,I420924,I420979,I464927,I421005,I421022,I421044,I464918,I421070,I421078,I464915,I421095,I421112,I464924,I421129,I464933,I421146,I421163,I464912,I421180,I421211,I421242,I464921,I421259,I421276,I421293,I421324,I421369,I464936,I421386,I421403,I464930,I421429,I421437,I421468,I421485,I421540,I421566,I421583,I421532,I421605,I421631,I421639,I421656,I421673,I421690,I421707,I421724,I421741,I421514,I421772,I421517,I421803,I421820,I421837,I421854,I421526,I421885,I421529,I421523,I421930,I421947,I421964,I421990,I421998,I421511,I422029,I422046,I421520,I422101,I422127,I422144,I422166,I422192,I422200,I422217,I422234,I422251,I422268,I422285,I422302,I422333,I422364,I422381,I422398,I422415,I422446,I422491,I422508,I422525,I422551,I422559,I422590,I422607,I422662,I422688,I422705,I422727,I422753,I422761,I422778,I422795,I422812,I422829,I422846,I422863,I422894,I422925,I422942,I422959,I422976,I423007,I423052,I423069,I423086,I423112,I423120,I423151,I423168,I423223,I482845,I423249,I423266,I423288,I482836,I423314,I423322,I482833,I423339,I423356,I482842,I423373,I482851,I423390,I423407,I482830,I423424,I423455,I423486,I482839,I423503,I423520,I423537,I423568,I423613,I482854,I423630,I423647,I482848,I423673,I423681,I423712,I423729,I423784,I423810,I423827,I423849,I423875,I423883,I423900,I423917,I423934,I423951,I423968,I423985,I424016,I424047,I424064,I424081,I424098,I424129,I424174,I424191,I424208,I424234,I424242,I424273,I424290,I424345,I491515,I424371,I424388,I424410,I491506,I424436,I424444,I491503,I424461,I424478,I491512,I424495,I491521,I424512,I424529,I491500,I424546,I424577,I424608,I491509,I424625,I424642,I424659,I424690,I424735,I491524,I424752,I424769,I491518,I424795,I424803,I424834,I424851,I424906,I424932,I424949,I424898,I424971,I424997,I425005,I425022,I425039,I425056,I425073,I425090,I425107,I424880,I425138,I424883,I425169,I425186,I425203,I425220,I424892,I425251,I424895,I424889,I425296,I425313,I425330,I425356,I425364,I424877,I425395,I425412,I424886,I425467,I425493,I425510,I425532,I425558,I425566,I425583,I425600,I425617,I425634,I425651,I425668,I425699,I425730,I425747,I425764,I425781,I425812,I425857,I425874,I425891,I425917,I425925,I425956,I425973,I426028,I426054,I426071,I426093,I426119,I426127,I426144,I426161,I426178,I426195,I426212,I426229,I426260,I426291,I426308,I426325,I426342,I426373,I426418,I426435,I426452,I426478,I426486,I426517,I426534,I426589,I426615,I426632,I426654,I426680,I426688,I426705,I426722,I426739,I426756,I426773,I426790,I426821,I426852,I426869,I426886,I426903,I426934,I426979,I426996,I427013,I427039,I427047,I427078,I427095,I427150,I452789,I427176,I427193,I427215,I452780,I427241,I427249,I452777,I427266,I427283,I452786,I427300,I452795,I427317,I427334,I452774,I427351,I427382,I427413,I452783,I427430,I427447,I427464,I427495,I427540,I452798,I427557,I427574,I452792,I427600,I427608,I427639,I427656,I427711,I485157,I427737,I427754,I427776,I485148,I427802,I427810,I485145,I427827,I427844,I485154,I427861,I485163,I427878,I427895,I485142,I427912,I427943,I427974,I485151,I427991,I428008,I428025,I428056,I428101,I485166,I428118,I428135,I485160,I428161,I428169,I428200,I428217,I428272,I428298,I428315,I428264,I428337,I428363,I428371,I428388,I428405,I428422,I428439,I428456,I428473,I428246,I428504,I428249,I428535,I428552,I428569,I428586,I428258,I428617,I428261,I428255,I428662,I428679,I428696,I428722,I428730,I428243,I428761,I428778,I428252,I428833,I428859,I428876,I428898,I428924,I428932,I428949,I428966,I428983,I429000,I429017,I429034,I429065,I429096,I429113,I429130,I429147,I429178,I429223,I429240,I429257,I429283,I429291,I429322,I429339,I429394,I429420,I429437,I429386,I429459,I429485,I429493,I429510,I429527,I429544,I429561,I429578,I429595,I429368,I429626,I429371,I429657,I429674,I429691,I429708,I429380,I429739,I429383,I429377,I429784,I429801,I429818,I429844,I429852,I429365,I429883,I429900,I429374,I429955,I489781,I429981,I429998,I430020,I489772,I430046,I430054,I489769,I430071,I430088,I489778,I430105,I489787,I430122,I430139,I489766,I430156,I430187,I430218,I489775,I430235,I430252,I430269,I430300,I430345,I489790,I430362,I430379,I489784,I430405,I430413,I430444,I430461,I430516,I520063,I430542,I430559,I430581,I520060,I430607,I430615,I520066,I430632,I430649,I520075,I430666,I520069,I430683,I430700,I520081,I430717,I430748,I430779,I520078,I430796,I430813,I430830,I430861,I430906,I520072,I430923,I520084,I430940,I430966,I430974,I431005,I431022,I431077,I431103,I431120,I431142,I431168,I431176,I431193,I431210,I431227,I431244,I431261,I431278,I431309,I431340,I431357,I431374,I431391,I431422,I431467,I431484,I431501,I431527,I431535,I431566,I431583,I431638,I526421,I431664,I431681,I431703,I526418,I431729,I431737,I526424,I431754,I431771,I526433,I431788,I526427,I431805,I431822,I526439,I431839,I431870,I431901,I526436,I431918,I431935,I431952,I431983,I432028,I526430,I432045,I526442,I432062,I432088,I432096,I432127,I432144,I432199,I432225,I432242,I432264,I432290,I432298,I432315,I432332,I432349,I432366,I432383,I432400,I432431,I432462,I432479,I432496,I432513,I432544,I432589,I432606,I432623,I432649,I432657,I432688,I432705,I432760,I432786,I432803,I432825,I432851,I432859,I432876,I432893,I432910,I432927,I432944,I432961,I432992,I433023,I433040,I433057,I433074,I433105,I433150,I433167,I433184,I433210,I433218,I433249,I433266,I433321,I433347,I433364,I433386,I433412,I433420,I433437,I433454,I433471,I433488,I433505,I433522,I433553,I433584,I433601,I433618,I433635,I433666,I433711,I433728,I433745,I433771,I433779,I433810,I433827,I433882,I433908,I433925,I433874,I433947,I433973,I433981,I433998,I434015,I434032,I434049,I434066,I434083,I433856,I434114,I433859,I434145,I434162,I434179,I434196,I433868,I434227,I433871,I433865,I434272,I434289,I434306,I434332,I434340,I433853,I434371,I434388,I433862,I434443,I434469,I434486,I434508,I434534,I434542,I434559,I434576,I434593,I434610,I434627,I434644,I434675,I434706,I434723,I434740,I434757,I434788,I434833,I434850,I434867,I434893,I434901,I434932,I434949,I435004,I435030,I435047,I435069,I435095,I435103,I435120,I435137,I435154,I435171,I435188,I435205,I435236,I435267,I435284,I435301,I435318,I435349,I435394,I435411,I435428,I435454,I435462,I435493,I435510,I435565,I435591,I435608,I435557,I435630,I435656,I435664,I435681,I435698,I435715,I435732,I435749,I435766,I435539,I435797,I435542,I435828,I435845,I435862,I435879,I435551,I435910,I435554,I435548,I435955,I435972,I435989,I436015,I436023,I435536,I436054,I436071,I435545,I436126,I451633,I436152,I436169,I436118,I436191,I451624,I436217,I436225,I451621,I436242,I436259,I451630,I436276,I451639,I436293,I436310,I451618,I436327,I436100,I436358,I436103,I436389,I451627,I436406,I436423,I436440,I436112,I436471,I436115,I436109,I436516,I451642,I436533,I436550,I451636,I436576,I436584,I436097,I436615,I436632,I436106,I436687,I570140,I436713,I436730,I436752,I570134,I436778,I436786,I570125,I436803,I436820,I570152,I436837,I570137,I570146,I436854,I436871,I570131,I436888,I436919,I436950,I570149,I436967,I436984,I437001,I437032,I437077,I570143,I437094,I437111,I570128,I437137,I437145,I437176,I437193,I437248,I437274,I437291,I437240,I437313,I437339,I437347,I437364,I437381,I437398,I437415,I437432,I437449,I437222,I437480,I437225,I437511,I437528,I437545,I437562,I437234,I437593,I437237,I437231,I437638,I437655,I437672,I437698,I437706,I437219,I437737,I437754,I437228,I437809,I437835,I437852,I437801,I437874,I437900,I437908,I437925,I437942,I437959,I437976,I437993,I438010,I437783,I438041,I437786,I438072,I438089,I438106,I438123,I437795,I438154,I437798,I437792,I438199,I438216,I438233,I438259,I438267,I437780,I438298,I438315,I437789,I438370,I438396,I438413,I438435,I438461,I438469,I438486,I438503,I438520,I438537,I438554,I438571,I438602,I438633,I438650,I438667,I438684,I438715,I438760,I438777,I438794,I438820,I438828,I438859,I438876,I438934,I438960,I438968,I439008,I439016,I439033,I439050,I439090,I439112,I439129,I439155,I439163,I439180,I439197,I439214,I439231,I439276,I439307,I439324,I439350,I439358,I439389,I439406,I439423,I439440,I439512,I439538,I439546,I439586,I439594,I439611,I439628,I439668,I439690,I439707,I439733,I439741,I439758,I439775,I439792,I439809,I439854,I439885,I439902,I439928,I439936,I439967,I439984,I440001,I440018,I440090,I440116,I440124,I440073,I440164,I440172,I440189,I440206,I440061,I440246,I440082,I440268,I440285,I440311,I440319,I440336,I440353,I440370,I440387,I440058,I440079,I440432,I440070,I440463,I440480,I440506,I440514,I440076,I440545,I440562,I440579,I440596,I440067,I440064,I440668,I440694,I440702,I440742,I440750,I440767,I440784,I440824,I440846,I440863,I440889,I440897,I440914,I440931,I440948,I440965,I441010,I441041,I441058,I441084,I441092,I441123,I441140,I441157,I441174,I441246,I441272,I441280,I441320,I441328,I441345,I441362,I441402,I441424,I441441,I441467,I441475,I441492,I441509,I441526,I441543,I441588,I441619,I441636,I441662,I441670,I441701,I441718,I441735,I441752,I441824,I441850,I441858,I441898,I441906,I441923,I441940,I441980,I442002,I442019,I442045,I442053,I442070,I442087,I442104,I442121,I442166,I442197,I442214,I442240,I442248,I442279,I442296,I442313,I442330,I442402,I552302,I442428,I442436,I552284,I552275,I442476,I442484,I552290,I442501,I552278,I442518,I442558,I442580,I552287,I442597,I442623,I442631,I442648,I552296,I442665,I442682,I442699,I442744,I552299,I442775,I442792,I552293,I552281,I442818,I442826,I442857,I442874,I442891,I442908,I442980,I443006,I443014,I443054,I443062,I443079,I443096,I443136,I443158,I443175,I443201,I443209,I443226,I443243,I443260,I443277,I443322,I443353,I443370,I443396,I443404,I443435,I443452,I443469,I443486,I443558,I443584,I443592,I443632,I443640,I443657,I443674,I443714,I443736,I443753,I443779,I443787,I443804,I443821,I443838,I443855,I443900,I443931,I443948,I443974,I443982,I444013,I444030,I444047,I444064,I444136,I444162,I444170,I444210,I444218,I444235,I444252,I444292,I444314,I444331,I444357,I444365,I444382,I444399,I444416,I444433,I444478,I444509,I444526,I444552,I444560,I444591,I444608,I444625,I444642,I444714,I561822,I444740,I444748,I561804,I561795,I444788,I444796,I561810,I444813,I561798,I444830,I444870,I444892,I561807,I444909,I444935,I444943,I444960,I561816,I444977,I444994,I445011,I445056,I561819,I445087,I445104,I561813,I561801,I445130,I445138,I445169,I445186,I445203,I445220,I445292,I445318,I445326,I445366,I445374,I445391,I445408,I445448,I445470,I445487,I445513,I445521,I445538,I445555,I445572,I445589,I445634,I445665,I445682,I445708,I445716,I445747,I445764,I445781,I445798,I445870,I445896,I445904,I445853,I445944,I445952,I445969,I445986,I445841,I446026,I445862,I446048,I446065,I446091,I446099,I446116,I446133,I446150,I446167,I445838,I445859,I446212,I445850,I446243,I446260,I446286,I446294,I445856,I446325,I446342,I446359,I446376,I445847,I445844,I446448,I446474,I446482,I446522,I446530,I446547,I446564,I446604,I446626,I446643,I446669,I446677,I446694,I446711,I446728,I446745,I446790,I446821,I446838,I446864,I446872,I446903,I446920,I446937,I446954,I447026,I447052,I447060,I447100,I447108,I447125,I447142,I447182,I447204,I447221,I447247,I447255,I447272,I447289,I447306,I447323,I447368,I447399,I447416,I447442,I447450,I447481,I447498,I447515,I447532,I447604,I447630,I447638,I447678,I447686,I447703,I447720,I447760,I447782,I447799,I447825,I447833,I447850,I447867,I447884,I447901,I447946,I447977,I447994,I448020,I448028,I448059,I448076,I448093,I448110,I448182,I448208,I448216,I448256,I448264,I448281,I448298,I448338,I448360,I448377,I448403,I448411,I448428,I448445,I448462,I448479,I448524,I448555,I448572,I448598,I448606,I448637,I448654,I448671,I448688,I448760,I448786,I448794,I448834,I448842,I448859,I448876,I448916,I448938,I448955,I448981,I448989,I449006,I449023,I449040,I449057,I449102,I449133,I449150,I449176,I449184,I449215,I449232,I449249,I449266,I449338,I449364,I449372,I449412,I449420,I449437,I449454,I449494,I449516,I449533,I449559,I449567,I449584,I449601,I449618,I449635,I449680,I449711,I449728,I449754,I449762,I449793,I449810,I449827,I449844,I449916,I449942,I449950,I449990,I449998,I450015,I450032,I450072,I450094,I450111,I450137,I450145,I450162,I450179,I450196,I450213,I450258,I450289,I450306,I450332,I450340,I450371,I450388,I450405,I450422,I450494,I450520,I450528,I450568,I450576,I450593,I450610,I450650,I450672,I450689,I450715,I450723,I450740,I450757,I450774,I450791,I450836,I450867,I450884,I450910,I450918,I450949,I450966,I450983,I451000,I451072,I451098,I451106,I451146,I451154,I451171,I451188,I451228,I451250,I451267,I451293,I451301,I451318,I451335,I451352,I451369,I451414,I451445,I451462,I451488,I451496,I451527,I451544,I451561,I451578,I451650,I555872,I451676,I451684,I555854,I555845,I451724,I451732,I555860,I451749,I555848,I451766,I451806,I451828,I555857,I451845,I451871,I451879,I451896,I555866,I451913,I451930,I451947,I451992,I555869,I452023,I452040,I555863,I555851,I452066,I452074,I452105,I452122,I452139,I452156,I452228,I452254,I452262,I452302,I452310,I452327,I452344,I452384,I452406,I452423,I452449,I452457,I452474,I452491,I452508,I452525,I452570,I452601,I452618,I452644,I452652,I452683,I452700,I452717,I452734,I452806,I452832,I452840,I452880,I452888,I452905,I452922,I452962,I452984,I453001,I453027,I453035,I453052,I453069,I453086,I453103,I453148,I453179,I453196,I453222,I453230,I453261,I453278,I453295,I453312,I453384,I453410,I453418,I453458,I453466,I453483,I453500,I453540,I453562,I453579,I453605,I453613,I453630,I453647,I453664,I453681,I453726,I453757,I453774,I453800,I453808,I453839,I453856,I453873,I453890,I453962,I453988,I453996,I454036,I454044,I454061,I454078,I454118,I454140,I454157,I454183,I454191,I454208,I454225,I454242,I454259,I454304,I454335,I454352,I454378,I454386,I454417,I454434,I454451,I454468,I454540,I454566,I454574,I454614,I454622,I454639,I454656,I454696,I454718,I454735,I454761,I454769,I454786,I454803,I454820,I454837,I454882,I454913,I454930,I454956,I454964,I454995,I455012,I455029,I455046,I455118,I455144,I455152,I455192,I455200,I455217,I455234,I455274,I455296,I455313,I455339,I455347,I455364,I455381,I455398,I455415,I455460,I455491,I455508,I455534,I455542,I455573,I455590,I455607,I455624,I455696,I455722,I455730,I455770,I455778,I455795,I455812,I455852,I455874,I455891,I455917,I455925,I455942,I455959,I455976,I455993,I456038,I456069,I456086,I456112,I456120,I456151,I456168,I456185,I456202,I456274,I456300,I456308,I456348,I456356,I456373,I456390,I456430,I456452,I456469,I456495,I456503,I456520,I456537,I456554,I456571,I456616,I456647,I456664,I456690,I456698,I456729,I456746,I456763,I456780,I456852,I456878,I456886,I456926,I456934,I456951,I456968,I457008,I457030,I457047,I457073,I457081,I457098,I457115,I457132,I457149,I457194,I457225,I457242,I457268,I457276,I457307,I457324,I457341,I457358,I457430,I457456,I457464,I457504,I457512,I457529,I457546,I457586,I457608,I457625,I457651,I457659,I457676,I457693,I457710,I457727,I457772,I457803,I457820,I457846,I457854,I457885,I457902,I457919,I457936,I458008,I458034,I458042,I457991,I458082,I458090,I458107,I458124,I457979,I458164,I458000,I458186,I458203,I458229,I458237,I458254,I458271,I458288,I458305,I457976,I457997,I458350,I457988,I458381,I458398,I458424,I458432,I457994,I458463,I458480,I458497,I458514,I457985,I457982,I458586,I516647,I458612,I458620,I516641,I516626,I458660,I458668,I516632,I458685,I516644,I458702,I458742,I458764,I458781,I458807,I458815,I458832,I516650,I458849,I516638,I458866,I458883,I458928,I516629,I458959,I458976,I516635,I459002,I459010,I459041,I459058,I459075,I459092,I459164,I459190,I459198,I459238,I459246,I459263,I459280,I459320,I459342,I459359,I459385,I459393,I459410,I459427,I459444,I459461,I459506,I459537,I459554,I459580,I459588,I459619,I459636,I459653,I459670,I459742,I459768,I459776,I459816,I459824,I459841,I459858,I459898,I459920,I459937,I459963,I459971,I459988,I460005,I460022,I460039,I460084,I460115,I460132,I460158,I460166,I460197,I460214,I460231,I460248,I460320,I460346,I460354,I460394,I460402,I460419,I460436,I460476,I460498,I460515,I460541,I460549,I460566,I460583,I460600,I460617,I460662,I460693,I460710,I460736,I460744,I460775,I460792,I460809,I460826,I460898,I460924,I460932,I460972,I460980,I460997,I461014,I461054,I461076,I461093,I461119,I461127,I461144,I461161,I461178,I461195,I461240,I461271,I461288,I461314,I461322,I461353,I461370,I461387,I461404,I461476,I461502,I461510,I461550,I461558,I461575,I461592,I461632,I461654,I461671,I461697,I461705,I461722,I461739,I461756,I461773,I461818,I461849,I461866,I461892,I461900,I461931,I461948,I461965,I461982,I462054,I462080,I462088,I462128,I462136,I462153,I462170,I462210,I462232,I462249,I462275,I462283,I462300,I462317,I462334,I462351,I462396,I462427,I462444,I462470,I462478,I462509,I462526,I462543,I462560,I462632,I462658,I462666,I462706,I462714,I462731,I462748,I462788,I462810,I462827,I462853,I462861,I462878,I462895,I462912,I462929,I462974,I463005,I463022,I463048,I463056,I463087,I463104,I463121,I463138,I463210,I463236,I463244,I463284,I463292,I463309,I463326,I463366,I463388,I463405,I463431,I463439,I463456,I463473,I463490,I463507,I463552,I463583,I463600,I463626,I463634,I463665,I463682,I463699,I463716,I463788,I572532,I463814,I463822,I572514,I572505,I463862,I463870,I572520,I463887,I572508,I463904,I463944,I463966,I572517,I463983,I464009,I464017,I464034,I572526,I464051,I464068,I464085,I464130,I572529,I464161,I464178,I572523,I572511,I464204,I464212,I464243,I464260,I464277,I464294,I464366,I464392,I464400,I464440,I464448,I464465,I464482,I464522,I464544,I464561,I464587,I464595,I464612,I464629,I464646,I464663,I464708,I464739,I464756,I464782,I464790,I464821,I464838,I464855,I464872,I464944,I464970,I464978,I465018,I465026,I465043,I465060,I465100,I465122,I465139,I465165,I465173,I465190,I465207,I465224,I465241,I465286,I465317,I465334,I465360,I465368,I465399,I465416,I465433,I465450,I465522,I465548,I465556,I465596,I465604,I465621,I465638,I465678,I465700,I465717,I465743,I465751,I465768,I465785,I465802,I465819,I465864,I465895,I465912,I465938,I465946,I465977,I465994,I466011,I466028,I466100,I466126,I466134,I466174,I466182,I466199,I466216,I466256,I466278,I466295,I466321,I466329,I466346,I466363,I466380,I466397,I466442,I466473,I466490,I466516,I466524,I466555,I466572,I466589,I466606,I466678,I466704,I466712,I466752,I466760,I466777,I466794,I466834,I466856,I466873,I466899,I466907,I466924,I466941,I466958,I466975,I467020,I467051,I467068,I467094,I467102,I467133,I467150,I467167,I467184,I467256,I467282,I467290,I467330,I467338,I467355,I467372,I467412,I467434,I467451,I467477,I467485,I467502,I467519,I467536,I467553,I467598,I467629,I467646,I467672,I467680,I467711,I467728,I467745,I467762,I467834,I467860,I467868,I467908,I467916,I467933,I467950,I467990,I468012,I468029,I468055,I468063,I468080,I468097,I468114,I468131,I468176,I468207,I468224,I468250,I468258,I468289,I468306,I468323,I468340,I468412,I468438,I468446,I468486,I468494,I468511,I468528,I468568,I468590,I468607,I468633,I468641,I468658,I468675,I468692,I468709,I468754,I468785,I468802,I468828,I468836,I468867,I468884,I468901,I468918,I468990,I469016,I469024,I469064,I469072,I469089,I469106,I469146,I469168,I469185,I469211,I469219,I469236,I469253,I469270,I469287,I469332,I469363,I469380,I469406,I469414,I469445,I469462,I469479,I469496,I469568,I469594,I469602,I469642,I469650,I469667,I469684,I469724,I469746,I469763,I469789,I469797,I469814,I469831,I469848,I469865,I469910,I469941,I469958,I469984,I469992,I470023,I470040,I470057,I470074,I470146,I470172,I470180,I470220,I470228,I470245,I470262,I470302,I470324,I470341,I470367,I470375,I470392,I470409,I470426,I470443,I470488,I470519,I470536,I470562,I470570,I470601,I470618,I470635,I470652,I470724,I534452,I470750,I470758,I534434,I534425,I470798,I470806,I534440,I470823,I534428,I470840,I470880,I470902,I534437,I470919,I470945,I470953,I470970,I534446,I470987,I471004,I471021,I471066,I534449,I471097,I471114,I534443,I534431,I471140,I471148,I471179,I471196,I471213,I471230,I471302,I538617,I471328,I471336,I538599,I538590,I471376,I471384,I538605,I471401,I538593,I471418,I471458,I471480,I538602,I471497,I471523,I471531,I471548,I538611,I471565,I471582,I471599,I471644,I538614,I471675,I471692,I538608,I538596,I471718,I471726,I471757,I471774,I471791,I471808,I471880,I471906,I471914,I471954,I471962,I471979,I471996,I472036,I472058,I472075,I472101,I472109,I472126,I472143,I472160,I472177,I472222,I472253,I472270,I472296,I472304,I472335,I472352,I472369,I472386,I472458,I472484,I472492,I472441,I472532,I472540,I472557,I472574,I472429,I472614,I472450,I472636,I472653,I472679,I472687,I472704,I472721,I472738,I472755,I472426,I472447,I472800,I472438,I472831,I472848,I472874,I472882,I472444,I472913,I472930,I472947,I472964,I472435,I472432,I473036,I473062,I473070,I473110,I473118,I473135,I473152,I473192,I473214,I473231,I473257,I473265,I473282,I473299,I473316,I473333,I473378,I473409,I473426,I473452,I473460,I473491,I473508,I473525,I473542,I473614,I473640,I473648,I473688,I473696,I473713,I473730,I473770,I473792,I473809,I473835,I473843,I473860,I473877,I473894,I473911,I473956,I473987,I474004,I474030,I474038,I474069,I474086,I474103,I474120,I474192,I474218,I474226,I474266,I474274,I474291,I474308,I474348,I474370,I474387,I474413,I474421,I474438,I474455,I474472,I474489,I474534,I474565,I474582,I474608,I474616,I474647,I474664,I474681,I474698,I474770,I474796,I474804,I474844,I474852,I474869,I474886,I474926,I474948,I474965,I474991,I474999,I475016,I475033,I475050,I475067,I475112,I475143,I475160,I475186,I475194,I475225,I475242,I475259,I475276,I475348,I475374,I475382,I475422,I475430,I475447,I475464,I475504,I475526,I475543,I475569,I475577,I475594,I475611,I475628,I475645,I475690,I475721,I475738,I475764,I475772,I475803,I475820,I475837,I475854,I475926,I553492,I475952,I475960,I553474,I553465,I476000,I476008,I553480,I476025,I553468,I476042,I476082,I476104,I553477,I476121,I476147,I476155,I476172,I553486,I476189,I476206,I476223,I476268,I553489,I476299,I476316,I553483,I553471,I476342,I476350,I476381,I476398,I476415,I476432,I476504,I503047,I476530,I476538,I503041,I503026,I476578,I476586,I503032,I476603,I503044,I476620,I476660,I476682,I476699,I476725,I476733,I476750,I503050,I476767,I503038,I476784,I476801,I476846,I503029,I476877,I476894,I503035,I476920,I476928,I476959,I476976,I476993,I477010,I477082,I477108,I477116,I477065,I477156,I477164,I477181,I477198,I477053,I477238,I477074,I477260,I477277,I477303,I477311,I477328,I477345,I477362,I477379,I477050,I477071,I477424,I477062,I477455,I477472,I477498,I477506,I477068,I477537,I477554,I477571,I477588,I477059,I477056,I477660,I477686,I477694,I477643,I477734,I477742,I477759,I477776,I477631,I477816,I477652,I477838,I477855,I477881,I477889,I477906,I477923,I477940,I477957,I477628,I477649,I478002,I477640,I478033,I478050,I478076,I478084,I477646,I478115,I478132,I478149,I478166,I477637,I477634,I478238,I478264,I478272,I478312,I478320,I478337,I478354,I478394,I478416,I478433,I478459,I478467,I478484,I478501,I478518,I478535,I478580,I478611,I478628,I478654,I478662,I478693,I478710,I478727,I478744,I478816,I478842,I478850,I478890,I478898,I478915,I478932,I478972,I478994,I479011,I479037,I479045,I479062,I479079,I479096,I479113,I479158,I479189,I479206,I479232,I479240,I479271,I479288,I479305,I479322,I479394,I479420,I479428,I479468,I479476,I479493,I479510,I479550,I479572,I479589,I479615,I479623,I479640,I479657,I479674,I479691,I479736,I479767,I479784,I479810,I479818,I479849,I479866,I479883,I479900,I479972,I479998,I480006,I480046,I480054,I480071,I480088,I480128,I480150,I480167,I480193,I480201,I480218,I480235,I480252,I480269,I480314,I480345,I480362,I480388,I480396,I480427,I480444,I480461,I480478,I480550,I480576,I480584,I480624,I480632,I480649,I480666,I480706,I480728,I480745,I480771,I480779,I480796,I480813,I480830,I480847,I480892,I480923,I480940,I480966,I480974,I481005,I481022,I481039,I481056,I481128,I549922,I481154,I481162,I549904,I549895,I481202,I481210,I549910,I481227,I549898,I481244,I481284,I481306,I549907,I481323,I481349,I481357,I481374,I549916,I481391,I481408,I481425,I481470,I549919,I481501,I481518,I549913,I549901,I481544,I481552,I481583,I481600,I481617,I481634,I481706,I481732,I481740,I481780,I481788,I481805,I481822,I481862,I481884,I481901,I481927,I481935,I481952,I481969,I481986,I482003,I482048,I482079,I482096,I482122,I482130,I482161,I482178,I482195,I482212,I482284,I545757,I482310,I482318,I545739,I482267,I545730,I482358,I482366,I545745,I482383,I545733,I482400,I482255,I482440,I482276,I482462,I545742,I482479,I482505,I482513,I482530,I545751,I482547,I482564,I482581,I482252,I482273,I482626,I545754,I482264,I482657,I482674,I545748,I545736,I482700,I482708,I482270,I482739,I482756,I482773,I482790,I482261,I482258,I482862,I482888,I482896,I482936,I482944,I482961,I482978,I483018,I483040,I483057,I483083,I483091,I483108,I483125,I483142,I483159,I483204,I483235,I483252,I483278,I483286,I483317,I483334,I483351,I483368,I483440,I483466,I483474,I483514,I483522,I483539,I483556,I483596,I483618,I483635,I483661,I483669,I483686,I483703,I483720,I483737,I483782,I483813,I483830,I483856,I483864,I483895,I483912,I483929,I483946,I484018,I484044,I484052,I484092,I484100,I484117,I484134,I484174,I484196,I484213,I484239,I484247,I484264,I484281,I484298,I484315,I484360,I484391,I484408,I484434,I484442,I484473,I484490,I484507,I484524,I484596,I555277,I484622,I484630,I555259,I555250,I484670,I484678,I555265,I484695,I555253,I484712,I484752,I484774,I555262,I484791,I484817,I484825,I484842,I555271,I484859,I484876,I484893,I484938,I555274,I484969,I484986,I555268,I555256,I485012,I485020,I485051,I485068,I485085,I485102,I485174,I485200,I485208,I485248,I485256,I485273,I485290,I485330,I485352,I485369,I485395,I485403,I485420,I485437,I485454,I485471,I485516,I485547,I485564,I485590,I485598,I485629,I485646,I485663,I485680,I485752,I485778,I485786,I485826,I485834,I485851,I485868,I485908,I485930,I485947,I485973,I485981,I485998,I486015,I486032,I486049,I486094,I486125,I486142,I486168,I486176,I486207,I486224,I486241,I486258,I486330,I486356,I486364,I486404,I486412,I486429,I486446,I486486,I486508,I486525,I486551,I486559,I486576,I486593,I486610,I486627,I486672,I486703,I486720,I486746,I486754,I486785,I486802,I486819,I486836,I486908,I486934,I486942,I486982,I486990,I487007,I487024,I487064,I487086,I487103,I487129,I487137,I487154,I487171,I487188,I487205,I487250,I487281,I487298,I487324,I487332,I487363,I487380,I487397,I487414,I487486,I487512,I487520,I487560,I487568,I487585,I487602,I487642,I487664,I487681,I487707,I487715,I487732,I487749,I487766,I487783,I487828,I487859,I487876,I487902,I487910,I487941,I487958,I487975,I487992,I488064,I507943,I488090,I488098,I507937,I507922,I488138,I488146,I507928,I488163,I507940,I488180,I488220,I488242,I488259,I488285,I488293,I488310,I507946,I488327,I507934,I488344,I488361,I488406,I507925,I488437,I488454,I507931,I488480,I488488,I488519,I488536,I488553,I488570,I488642,I488668,I488676,I488716,I488724,I488741,I488758,I488798,I488820,I488837,I488863,I488871,I488888,I488905,I488922,I488939,I488984,I489015,I489032,I489058,I489066,I489097,I489114,I489131,I489148,I489220,I489246,I489254,I489294,I489302,I489319,I489336,I489376,I489398,I489415,I489441,I489449,I489466,I489483,I489500,I489517,I489562,I489593,I489610,I489636,I489644,I489675,I489692,I489709,I489726,I489798,I489824,I489832,I489872,I489880,I489897,I489914,I489954,I489976,I489993,I490019,I490027,I490044,I490061,I490078,I490095,I490140,I490171,I490188,I490214,I490222,I490253,I490270,I490287,I490304,I490376,I490402,I490410,I490450,I490458,I490475,I490492,I490532,I490554,I490571,I490597,I490605,I490622,I490639,I490656,I490673,I490718,I490749,I490766,I490792,I490800,I490831,I490848,I490865,I490882,I490954,I490980,I490988,I490937,I491028,I491036,I491053,I491070,I490925,I491110,I490946,I491132,I491149,I491175,I491183,I491200,I491217,I491234,I491251,I490922,I490943,I491296,I490934,I491327,I491344,I491370,I491378,I490940,I491409,I491426,I491443,I491460,I490931,I490928,I491532,I491558,I491566,I491606,I491614,I491631,I491648,I491688,I491710,I491727,I491753,I491761,I491778,I491795,I491812,I491829,I491874,I491905,I491922,I491948,I491956,I491987,I492004,I492021,I492038,I492110,I492136,I492144,I492184,I492192,I492209,I492226,I492266,I492288,I492305,I492331,I492339,I492356,I492373,I492390,I492407,I492452,I492483,I492500,I492526,I492534,I492565,I492582,I492599,I492616,I492688,I509031,I492714,I492722,I509025,I509010,I492762,I492770,I509016,I492787,I509028,I492804,I492844,I492866,I492883,I492909,I492917,I492934,I509034,I492951,I509022,I492968,I492985,I493030,I509013,I493061,I493078,I509019,I493104,I493112,I493143,I493160,I493177,I493194,I493266,I493292,I493300,I493340,I493348,I493365,I493382,I493422,I493444,I493461,I493487,I493495,I493512,I493529,I493546,I493563,I493608,I493639,I493656,I493682,I493690,I493721,I493738,I493755,I493772,I493844,I521818,I493870,I493878,I521800,I521809,I493918,I493926,I521794,I493943,I521806,I493960,I494000,I494022,I521797,I494039,I494065,I494073,I494090,I494107,I494124,I494141,I494186,I521815,I494217,I494234,I521803,I521812,I494260,I494268,I494299,I494316,I494333,I494350,I494422,I562417,I494448,I494456,I562399,I562390,I494496,I494504,I562405,I494521,I562393,I494538,I494578,I494600,I562402,I494617,I494643,I494651,I494668,I562411,I494685,I494702,I494719,I494764,I562414,I494795,I494812,I562408,I562396,I494838,I494846,I494877,I494894,I494911,I494928,I495000,I495026,I495034,I495074,I495082,I495099,I495116,I495156,I495178,I495195,I495221,I495229,I495246,I495263,I495280,I495297,I495342,I495373,I495390,I495416,I495424,I495455,I495472,I495489,I495506,I495578,I495604,I495612,I495652,I495660,I495677,I495694,I495734,I495756,I495773,I495799,I495807,I495824,I495841,I495858,I495875,I495920,I495951,I495968,I495994,I496002,I496033,I496050,I496067,I496084,I496156,I496182,I496190,I496230,I496238,I496255,I496272,I496312,I496334,I496351,I496377,I496385,I496402,I496419,I496436,I496453,I496498,I496529,I496546,I496572,I496580,I496611,I496628,I496645,I496662,I496734,I496760,I496768,I496808,I496816,I496833,I496850,I496890,I496912,I496929,I496955,I496963,I496980,I496997,I497014,I497031,I497076,I497107,I497124,I497150,I497158,I497189,I497206,I497223,I497240,I497312,I497338,I497346,I497386,I497394,I497411,I497428,I497468,I497490,I497507,I497533,I497541,I497558,I497575,I497592,I497609,I497654,I497685,I497702,I497728,I497736,I497767,I497784,I497801,I497818,I497890,I497916,I497924,I497964,I497972,I497989,I498006,I498046,I498068,I498085,I498111,I498119,I498136,I498153,I498170,I498187,I498232,I498263,I498280,I498306,I498314,I498345,I498362,I498379,I498396,I498468,I510663,I498494,I498502,I510657,I498451,I510642,I498542,I498550,I510648,I498567,I510660,I498584,I498439,I498624,I498460,I498646,I498663,I498689,I498697,I498714,I510666,I498731,I510654,I498748,I498765,I498436,I498457,I498810,I510645,I498448,I498841,I498858,I510651,I498884,I498892,I498454,I498923,I498940,I498957,I498974,I498445,I498442,I499046,I499072,I499080,I499120,I499128,I499145,I499162,I499202,I499224,I499241,I499267,I499275,I499292,I499309,I499326,I499343,I499388,I499419,I499436,I499462,I499470,I499501,I499518,I499535,I499552,I499624,I499650,I499658,I499698,I499706,I499723,I499740,I499780,I499802,I499819,I499845,I499853,I499870,I499887,I499904,I499921,I499966,I499997,I500014,I500040,I500048,I500079,I500096,I500113,I500130,I500202,I500228,I500236,I500276,I500284,I500301,I500318,I500358,I500380,I500397,I500423,I500431,I500448,I500465,I500482,I500499,I500544,I500575,I500592,I500618,I500626,I500657,I500674,I500691,I500708,I500780,I500806,I500814,I500854,I500862,I500879,I500896,I500936,I500958,I500975,I501001,I501009,I501026,I501043,I501060,I501077,I501122,I501153,I501170,I501196,I501204,I501235,I501252,I501269,I501286,I501358,I501384,I501392,I501432,I501440,I501457,I501474,I501514,I501536,I501553,I501579,I501587,I501604,I501621,I501638,I501655,I501700,I501731,I501748,I501774,I501782,I501813,I501830,I501847,I501864,I501936,I501962,I501970,I502010,I502018,I502035,I502052,I502092,I502114,I502131,I502157,I502165,I502182,I502199,I502216,I502233,I502278,I502309,I502326,I502352,I502360,I502391,I502408,I502425,I502442,I502514,I502540,I502548,I502574,I502591,I502613,I502630,I502647,I502664,I502681,I502712,I502729,I502746,I502763,I502808,I502825,I502842,I502901,I502927,I502935,I502952,I502969,I503000,I503058,I531051,I503084,I503092,I531060,I531063,I503118,I503135,I503157,I531057,I503174,I531054,I503191,I531048,I503208,I503225,I503256,I531045,I503273,I531042,I503290,I503307,I503352,I503369,I503386,I503445,I531066,I503471,I503479,I503496,I503513,I503544,I503602,I503628,I503636,I503662,I503679,I503701,I503718,I503735,I503752,I503769,I503800,I503817,I503834,I503851,I503896,I503913,I503930,I503989,I504015,I504023,I504040,I504057,I504088,I504146,I557657,I504172,I504180,I557642,I557636,I504206,I504223,I504138,I504245,I557630,I504262,I557651,I504279,I557639,I504296,I504313,I504117,I504344,I557648,I504361,I557654,I504378,I557645,I504395,I504120,I504135,I504440,I557633,I504457,I504474,I504132,I504129,I504126,I504533,I504559,I504567,I504584,I504601,I504114,I504632,I504123,I504690,I504716,I504724,I504750,I504767,I504789,I504806,I504823,I504840,I504857,I504888,I504905,I504922,I504939,I504984,I505001,I505018,I505077,I505103,I505111,I505128,I505145,I505176,I505234,I505260,I505268,I505294,I505311,I505333,I505350,I505367,I505384,I505401,I505432,I505449,I505466,I505483,I505528,I505545,I505562,I505621,I505647,I505655,I505672,I505689,I505720,I505778,I540997,I505804,I505812,I540982,I540976,I505838,I505855,I505877,I540970,I505894,I540991,I505911,I540979,I505928,I505945,I505976,I540988,I505993,I540994,I506010,I540985,I506027,I506072,I540973,I506089,I506106,I506165,I506191,I506199,I506216,I506233,I506264,I506322,I573722,I506348,I506356,I573707,I573701,I506382,I506399,I506421,I573695,I506438,I573716,I506455,I573704,I506472,I506489,I506520,I573713,I506537,I573719,I506554,I573710,I506571,I506616,I573698,I506633,I506650,I506709,I506735,I506743,I506760,I506777,I506808,I506866,I539212,I506892,I506900,I539197,I539191,I506926,I506943,I506965,I539185,I506982,I539206,I506999,I539194,I507016,I507033,I507064,I539203,I507081,I539209,I507098,I539200,I507115,I507160,I539188,I507177,I507194,I507253,I507279,I507287,I507304,I507321,I507352,I507410,I507436,I507444,I507470,I507487,I507509,I507526,I507543,I507560,I507577,I507608,I507625,I507642,I507659,I507704,I507721,I507738,I507797,I507823,I507831,I507848,I507865,I507896,I507954,I507980,I507988,I508014,I508031,I508053,I508070,I508087,I508104,I508121,I508152,I508169,I508186,I508203,I508248,I508265,I508282,I508341,I508367,I508375,I508392,I508409,I508440,I508498,I508524,I508532,I508558,I508575,I508597,I508614,I508631,I508648,I508665,I508696,I508713,I508730,I508747,I508792,I508809,I508826,I508885,I508911,I508919,I508936,I508953,I508984,I509042,I509068,I509076,I509102,I509119,I509141,I509158,I509175,I509192,I509209,I509240,I509257,I509274,I509291,I509336,I509353,I509370,I509429,I509455,I509463,I509480,I509497,I509528,I509586,I509612,I509620,I509646,I509663,I509685,I509702,I509719,I509736,I509753,I509784,I509801,I509818,I509835,I509880,I509897,I509914,I509973,I509999,I510007,I510024,I510041,I510072,I510130,I510156,I510164,I510190,I510207,I510229,I510246,I510263,I510280,I510297,I510328,I510345,I510362,I510379,I510424,I510441,I510458,I510517,I510543,I510551,I510568,I510585,I510616,I510674,I510700,I510708,I510734,I510751,I510773,I510790,I510807,I510824,I510841,I510872,I510889,I510906,I510923,I510968,I510985,I511002,I511061,I511087,I511095,I511112,I511129,I511160,I511218,I511244,I511252,I511278,I511295,I511317,I511334,I511351,I511368,I511385,I511416,I511433,I511450,I511467,I511512,I511529,I511546,I511605,I511631,I511639,I511656,I511673,I511704,I511762,I558252,I511788,I511796,I558237,I558231,I511822,I511839,I511861,I558225,I511878,I558246,I511895,I558234,I511912,I511929,I511960,I558243,I511977,I558249,I511994,I558240,I512011,I512056,I558228,I512073,I512090,I512149,I512175,I512183,I512200,I512217,I512248,I512306,I512332,I512340,I512366,I512383,I512405,I512422,I512439,I512456,I512473,I512504,I512521,I512538,I512555,I512600,I512617,I512634,I512693,I512719,I512727,I512744,I512761,I512792,I512850,I512876,I512884,I512910,I512927,I512842,I512949,I512966,I512983,I513000,I513017,I512821,I513048,I513065,I513082,I513099,I512824,I512839,I513144,I513161,I513178,I512836,I512833,I512830,I513237,I513263,I513271,I513288,I513305,I512818,I513336,I512827,I513394,I513420,I513428,I513454,I513471,I513493,I513510,I513527,I513544,I513561,I513592,I513609,I513626,I513643,I513688,I513705,I513722,I513781,I513807,I513815,I513832,I513849,I513880,I513938,I513964,I513972,I513998,I514015,I514037,I514054,I514071,I514088,I514105,I514136,I514153,I514170,I514187,I514232,I514249,I514266,I514325,I514351,I514359,I514376,I514393,I514424,I514482,I514508,I514516,I514542,I514559,I514581,I514598,I514615,I514632,I514649,I514680,I514697,I514714,I514731,I514776,I514793,I514810,I514869,I514895,I514903,I514920,I514937,I514968,I515026,I515052,I515060,I515086,I515103,I515125,I515142,I515159,I515176,I515193,I515224,I515241,I515258,I515275,I515320,I515337,I515354,I515413,I515439,I515447,I515464,I515481,I515512,I515570,I515596,I515604,I515630,I515647,I515669,I515686,I515703,I515720,I515737,I515768,I515785,I515802,I515819,I515864,I515881,I515898,I515957,I515983,I515991,I516008,I516025,I516056,I516114,I516140,I516148,I516174,I516191,I516213,I516230,I516247,I516264,I516281,I516312,I516329,I516346,I516363,I516408,I516425,I516442,I516501,I516527,I516535,I516552,I516569,I516600,I516658,I516684,I516692,I516718,I516735,I516757,I516774,I516791,I516808,I516825,I516856,I516873,I516890,I516907,I516952,I516969,I516986,I517045,I517071,I517079,I517096,I517113,I517144,I517202,I517228,I517236,I517253,I517279,I517287,I517304,I517321,I517338,I517355,I517386,I517403,I517420,I517451,I517468,I517508,I517516,I517547,I517564,I517581,I517598,I517629,I517660,I517686,I517708,I517780,I517806,I517814,I517831,I517857,I517865,I517882,I517899,I517916,I517933,I517964,I517981,I517998,I518029,I518046,I518086,I518094,I518125,I518142,I518159,I518176,I518207,I518238,I518264,I518286,I518358,I518384,I518392,I518409,I518435,I518443,I518460,I518477,I518494,I518511,I518542,I518559,I518576,I518607,I518624,I518664,I518672,I518703,I518720,I518737,I518754,I518785,I518816,I518842,I518864,I518936,I518962,I518970,I518987,I519013,I519021,I519038,I519055,I519072,I519089,I519120,I519137,I519154,I519185,I519202,I519242,I519250,I519281,I519298,I519315,I519332,I519363,I519394,I519420,I519442,I519514,I519540,I519548,I519565,I519591,I519599,I519616,I519633,I519650,I519667,I519698,I519715,I519732,I519763,I519780,I519820,I519828,I519859,I519876,I519893,I519910,I519941,I519972,I519998,I520020,I520092,I520118,I520126,I520143,I520169,I520177,I520194,I520211,I520228,I520245,I520276,I520293,I520310,I520341,I520358,I520398,I520406,I520437,I520454,I520471,I520488,I520519,I520550,I520576,I520598,I520670,I520696,I520704,I520721,I520747,I520755,I520772,I520789,I520806,I520823,I520662,I520854,I520871,I520888,I520641,I520919,I520936,I520647,I520976,I520984,I520656,I521015,I521032,I521049,I521066,I520659,I521097,I520638,I521128,I521154,I520653,I521176,I520650,I520644,I521248,I521274,I521282,I521299,I521325,I521333,I521350,I521367,I521384,I521401,I521432,I521449,I521466,I521497,I521514,I521554,I521562,I521593,I521610,I521627,I521644,I521675,I521706,I521732,I521754,I521826,I521852,I521860,I521877,I521903,I521911,I521928,I521945,I521962,I521979,I522010,I522027,I522044,I522075,I522092,I522132,I522140,I522171,I522188,I522205,I522222,I522253,I522284,I522310,I522332,I522404,I522430,I522438,I522455,I522481,I522489,I522506,I522523,I522540,I522557,I522588,I522605,I522622,I522653,I522670,I522710,I522718,I522749,I522766,I522783,I522800,I522831,I522862,I522888,I522910,I522982,I523008,I523016,I523033,I523059,I523067,I523084,I523101,I523118,I523135,I523166,I523183,I523200,I523231,I523248,I523288,I523296,I523327,I523344,I523361,I523378,I523409,I523440,I523466,I523488,I523560,I523586,I523594,I523611,I523637,I523645,I523662,I523679,I523696,I523713,I523552,I523744,I523761,I523778,I523531,I523809,I523826,I523537,I523866,I523874,I523546,I523905,I523922,I523939,I523956,I523549,I523987,I523528,I524018,I524044,I523543,I524066,I523540,I523534,I524138,I524164,I524172,I524189,I524215,I524223,I524240,I524257,I524274,I524291,I524322,I524339,I524356,I524387,I524404,I524444,I524452,I524483,I524500,I524517,I524534,I524565,I524596,I524622,I524644,I524716,I524742,I524750,I524767,I524793,I524801,I524818,I524835,I524852,I524869,I524708,I524900,I524917,I524934,I524687,I524965,I524982,I524693,I525022,I525030,I524702,I525061,I525078,I525095,I525112,I524705,I525143,I524684,I525174,I525200,I524699,I525222,I524696,I524690,I525294,I525320,I525328,I525345,I525371,I525379,I525396,I525413,I525430,I525447,I525478,I525495,I525512,I525543,I525560,I525600,I525608,I525639,I525656,I525673,I525690,I525721,I525752,I525778,I525800,I525872,I560034,I525898,I525906,I560025,I525923,I560010,I525949,I525957,I525974,I560013,I525991,I560022,I526008,I526025,I560019,I526056,I560031,I526073,I526090,I526121,I560016,I526138,I526178,I526186,I526217,I560037,I526234,I526251,I526268,I526299,I526330,I560028,I526356,I526378,I526450,I526476,I526484,I526501,I526527,I526535,I526552,I526569,I526586,I526603,I526634,I526651,I526668,I526699,I526716,I526756,I526764,I526795,I526812,I526829,I526846,I526877,I526908,I526934,I526956,I527028,I527054,I527062,I527079,I527105,I527113,I527130,I527147,I527164,I527181,I527212,I527229,I527246,I527277,I527294,I527334,I527342,I527373,I527390,I527407,I527424,I527455,I527486,I527512,I527534,I527606,I527632,I527640,I527657,I527683,I527691,I527708,I527725,I527742,I527759,I527790,I527807,I527824,I527855,I527872,I527912,I527920,I527951,I527968,I527985,I528002,I528033,I528064,I528090,I528112,I528184,I528210,I528218,I528235,I528261,I528269,I528286,I528303,I528320,I528337,I528368,I528385,I528402,I528433,I528450,I528490,I528498,I528529,I528546,I528563,I528580,I528611,I528642,I528668,I528690,I528762,I528788,I528796,I528813,I528839,I528847,I528864,I528881,I528898,I528915,I528946,I528963,I528980,I529011,I529028,I529068,I529076,I529107,I529124,I529141,I529158,I529189,I529220,I529246,I529268,I529340,I529366,I529374,I529391,I529417,I529425,I529442,I529459,I529476,I529493,I529524,I529541,I529558,I529589,I529606,I529646,I529654,I529685,I529702,I529719,I529736,I529767,I529798,I529824,I529846,I529918,I529944,I529952,I529969,I529995,I530003,I530020,I530037,I530054,I530071,I530102,I530119,I530136,I530167,I530184,I530224,I530232,I530263,I530280,I530297,I530314,I530345,I530376,I530402,I530424,I530496,I530522,I530530,I530547,I530573,I530581,I530598,I530615,I530632,I530649,I530680,I530697,I530714,I530745,I530762,I530802,I530810,I530841,I530858,I530875,I530892,I530923,I530954,I530980,I531002,I531074,I570744,I531100,I531108,I570735,I531125,I570720,I531151,I531159,I531176,I570723,I531193,I570732,I531210,I531227,I570729,I531258,I570741,I531275,I531292,I531323,I570726,I531340,I531380,I531388,I531419,I570747,I531436,I531453,I531470,I531501,I531532,I570738,I531558,I531580,I531655,I531681,I531689,I531706,I531732,I531740,I531757,I531774,I531805,I531836,I531853,I531870,I531887,I531904,I531935,I531994,I532011,I532037,I532059,I532085,I532093,I532110,I532141,I532216,I571925,I532242,I532250,I571919,I532267,I571937,I532293,I532301,I532318,I571922,I571913,I532335,I532366,I571928,I532397,I571931,I532414,I571934,I532431,I532448,I571916,I532465,I532496,I532555,I571910,I532572,I532598,I532620,I532646,I532654,I532671,I532702,I532777,I532803,I532811,I532828,I532854,I532862,I532879,I532896,I532927,I532958,I532975,I532992,I533009,I533026,I533057,I533116,I533133,I533159,I533181,I533207,I533215,I533232,I533263,I533338,I533364,I533372,I533389,I533415,I533423,I533440,I533457,I533324,I533488,I533327,I533519,I533536,I533553,I533570,I533587,I533312,I533618,I533315,I533309,I533306,I533677,I533694,I533720,I533330,I533742,I533768,I533776,I533793,I533321,I533824,I533303,I533318,I533899,I533925,I533933,I533950,I533976,I533984,I534001,I534018,I534049,I534080,I534097,I534114,I534131,I534148,I534179,I534238,I534255,I534281,I534303,I534329,I534337,I534354,I534385,I534460,I534486,I534503,I534511,I534556,I534573,I534590,I534607,I534624,I534641,I534658,I534689,I534706,I534751,I534768,I534785,I534816,I534842,I534850,I534881,I534898,I534915,I534941,I534949,I534966,I535055,I535081,I535098,I535106,I535151,I535168,I535185,I535202,I535219,I535236,I535253,I535284,I535301,I535346,I535363,I535380,I535411,I535437,I535445,I535476,I535493,I535510,I535536,I535544,I535561,I535650,I535676,I535693,I535701,I535746,I535763,I535780,I535797,I535814,I535831,I535848,I535879,I535896,I535941,I535958,I535975,I536006,I536032,I536040,I536071,I536088,I536105,I536131,I536139,I536156,I536245,I536271,I536288,I536296,I536341,I536358,I536375,I536392,I536409,I536426,I536443,I536474,I536491,I536536,I536553,I536570,I536601,I536627,I536635,I536666,I536683,I536700,I536726,I536734,I536751,I536840,I536866,I536883,I536891,I536936,I536953,I536970,I536987,I537004,I537021,I537038,I537069,I537086,I537131,I537148,I537165,I537196,I537222,I537230,I537261,I537278,I537295,I537321,I537329,I537346,I537435,I537461,I537478,I537486,I537531,I537548,I537565,I537582,I537599,I537616,I537633,I537664,I537681,I537726,I537743,I537760,I537791,I537817,I537825,I537856,I537873,I537890,I537916,I537924,I537941,I538030,I538056,I538073,I538081,I538126,I538143,I538160,I538177,I538194,I538211,I538228,I538259,I538276,I538321,I538338,I538355,I538386,I538412,I538420,I538451,I538468,I538485,I538511,I538519,I538536,I538625,I538651,I538668,I538676,I538721,I538738,I538755,I538772,I538789,I538806,I538823,I538854,I538871,I538916,I538933,I538950,I538981,I539007,I539015,I539046,I539063,I539080,I539106,I539114,I539131,I539220,I539246,I539263,I539271,I539316,I539333,I539350,I539367,I539384,I539401,I539418,I539449,I539466,I539511,I539528,I539545,I539576,I539602,I539610,I539641,I539658,I539675,I539701,I539709,I539726,I539815,I539841,I539858,I539866,I539911,I539928,I539945,I539962,I539979,I539996,I540013,I540044,I540061,I540106,I540123,I540140,I540171,I540197,I540205,I540236,I540253,I540270,I540296,I540304,I540321,I540410,I540436,I540453,I540461,I540506,I540523,I540540,I540557,I540574,I540591,I540608,I540639,I540656,I540701,I540718,I540735,I540766,I540792,I540800,I540831,I540848,I540865,I540891,I540899,I540916,I541005,I541031,I541048,I541056,I541101,I541118,I541135,I541152,I541169,I541186,I541203,I541234,I541251,I541296,I541313,I541330,I541361,I541387,I541395,I541426,I541443,I541460,I541486,I541494,I541511,I541600,I541626,I541643,I541651,I541696,I541713,I541730,I541747,I541764,I541781,I541798,I541829,I541846,I541891,I541908,I541925,I541956,I541982,I541990,I542021,I542038,I542055,I542081,I542089,I542106,I542195,I542221,I542238,I542246,I542291,I542308,I542325,I542342,I542359,I542376,I542393,I542424,I542441,I542486,I542503,I542520,I542551,I542577,I542585,I542616,I542633,I542650,I542676,I542684,I542701,I542790,I542816,I542833,I542841,I542886,I542903,I542920,I542937,I542954,I542971,I542988,I543019,I543036,I543081,I543098,I543115,I543146,I543172,I543180,I543211,I543228,I543245,I543271,I543279,I543296,I543385,I543411,I543428,I543436,I543481,I543498,I543515,I543532,I543549,I543566,I543583,I543614,I543631,I543676,I543693,I543710,I543741,I543767,I543775,I543806,I543823,I543840,I543866,I543874,I543891,I543980,I544006,I544023,I544031,I544076,I544093,I544110,I544127,I544144,I544161,I544178,I544209,I544226,I544271,I544288,I544305,I544336,I544362,I544370,I544401,I544418,I544435,I544461,I544469,I544486,I544575,I544601,I544618,I544626,I544671,I544688,I544705,I544722,I544739,I544756,I544773,I544804,I544821,I544866,I544883,I544900,I544931,I544957,I544965,I544996,I545013,I545030,I545056,I545064,I545081,I545170,I545196,I545213,I545221,I545266,I545283,I545300,I545317,I545334,I545351,I545368,I545399,I545416,I545461,I545478,I545495,I545526,I545552,I545560,I545591,I545608,I545625,I545651,I545659,I545676,I545765,I545791,I545808,I545816,I545861,I545878,I545895,I545912,I545929,I545946,I545963,I545994,I546011,I546056,I546073,I546090,I546121,I546147,I546155,I546186,I546203,I546220,I546246,I546254,I546271,I546360,I546386,I546403,I546411,I546456,I546473,I546490,I546507,I546524,I546541,I546558,I546589,I546606,I546651,I546668,I546685,I546716,I546742,I546750,I546781,I546798,I546815,I546841,I546849,I546866,I546955,I546981,I546998,I547006,I547051,I547068,I547085,I547102,I547119,I547136,I547153,I547184,I547201,I547246,I547263,I547280,I547311,I547337,I547345,I547376,I547393,I547410,I547436,I547444,I547461,I547550,I547576,I547593,I547601,I547646,I547663,I547680,I547697,I547714,I547731,I547748,I547779,I547796,I547841,I547858,I547875,I547906,I547932,I547940,I547971,I547988,I548005,I548031,I548039,I548056,I548145,I548171,I548188,I548196,I548241,I548258,I548275,I548292,I548309,I548326,I548343,I548374,I548391,I548436,I548453,I548470,I548501,I548527,I548535,I548566,I548583,I548600,I548626,I548634,I548651,I548740,I548766,I548783,I548791,I548836,I548853,I548870,I548887,I548904,I548921,I548938,I548969,I548986,I549031,I549048,I549065,I549096,I549122,I549130,I549161,I549178,I549195,I549221,I549229,I549246,I549335,I549361,I549378,I549386,I549431,I549448,I549465,I549482,I549499,I549516,I549533,I549564,I549581,I549626,I549643,I549660,I549691,I549717,I549725,I549756,I549773,I549790,I549816,I549824,I549841,I549930,I549956,I549973,I549981,I550026,I550043,I550060,I550077,I550094,I550111,I550128,I550159,I550176,I550221,I550238,I550255,I550286,I550312,I550320,I550351,I550368,I550385,I550411,I550419,I550436,I550525,I550551,I550568,I550576,I550621,I550638,I550655,I550672,I550689,I550706,I550723,I550754,I550771,I550816,I550833,I550850,I550881,I550907,I550915,I550946,I550963,I550980,I551006,I551014,I551031,I551120,I551146,I551163,I551171,I551216,I551233,I551250,I551267,I551284,I551301,I551318,I551349,I551366,I551411,I551428,I551445,I551476,I551502,I551510,I551541,I551558,I551575,I551601,I551609,I551626,I551715,I551741,I551758,I551766,I551811,I551828,I551845,I551862,I551879,I551896,I551913,I551944,I551961,I552006,I552023,I552040,I552071,I552097,I552105,I552136,I552153,I552170,I552196,I552204,I552221,I552310,I552336,I552353,I552361,I552406,I552423,I552440,I552457,I552474,I552491,I552508,I552539,I552556,I552601,I552618,I552635,I552666,I552692,I552700,I552731,I552748,I552765,I552791,I552799,I552816,I552905,I552931,I552948,I552956,I553001,I553018,I553035,I553052,I553069,I553086,I553103,I553134,I553151,I553196,I553213,I553230,I553261,I553287,I553295,I553326,I553343,I553360,I553386,I553394,I553411,I553500,I553526,I553543,I553551,I553596,I553613,I553630,I553647,I553664,I553681,I553698,I553729,I553746,I553791,I553808,I553825,I553856,I553882,I553890,I553921,I553938,I553955,I553981,I553989,I554006,I554095,I554121,I554138,I554146,I554191,I554208,I554225,I554242,I554259,I554276,I554293,I554324,I554341,I554386,I554403,I554420,I554451,I554477,I554485,I554516,I554533,I554550,I554576,I554584,I554601,I554690,I554716,I554733,I554741,I554786,I554803,I554820,I554837,I554854,I554871,I554888,I554919,I554936,I554981,I554998,I555015,I555046,I555072,I555080,I555111,I555128,I555145,I555171,I555179,I555196,I555285,I555311,I555328,I555336,I555381,I555398,I555415,I555432,I555449,I555466,I555483,I555514,I555531,I555576,I555593,I555610,I555641,I555667,I555675,I555706,I555723,I555740,I555766,I555774,I555791,I555880,I555906,I555923,I555931,I555976,I555993,I556010,I556027,I556044,I556061,I556078,I556109,I556126,I556171,I556188,I556205,I556236,I556262,I556270,I556301,I556318,I556335,I556361,I556369,I556386,I556475,I556501,I556518,I556526,I556571,I556588,I556605,I556622,I556639,I556656,I556673,I556704,I556721,I556766,I556783,I556800,I556831,I556857,I556865,I556896,I556913,I556930,I556956,I556964,I556981,I557070,I557096,I557113,I557121,I557166,I557183,I557200,I557217,I557234,I557251,I557268,I557299,I557316,I557361,I557378,I557395,I557426,I557452,I557460,I557491,I557508,I557525,I557551,I557559,I557576,I557665,I557691,I557708,I557716,I557761,I557778,I557795,I557812,I557829,I557846,I557863,I557894,I557911,I557956,I557973,I557990,I558021,I558047,I558055,I558086,I558103,I558120,I558146,I558154,I558171,I558260,I558286,I558303,I558311,I558356,I558373,I558390,I558407,I558424,I558441,I558458,I558489,I558506,I558551,I558568,I558585,I558616,I558642,I558650,I558681,I558698,I558715,I558741,I558749,I558766,I558855,I558881,I558898,I558906,I558951,I558968,I558985,I559002,I559019,I559036,I559053,I559084,I559101,I559146,I559163,I559180,I559211,I559237,I559245,I559276,I559293,I559310,I559336,I559344,I559361,I559450,I559476,I559493,I559501,I559546,I559563,I559580,I559597,I559614,I559631,I559648,I559679,I559696,I559741,I559758,I559775,I559806,I559832,I559840,I559871,I559888,I559905,I559931,I559939,I559956,I560045,I560071,I560088,I560096,I560141,I560158,I560175,I560192,I560209,I560226,I560243,I560274,I560291,I560336,I560353,I560370,I560401,I560427,I560435,I560466,I560483,I560500,I560526,I560534,I560551,I560640,I560666,I560683,I560691,I560736,I560753,I560770,I560787,I560804,I560821,I560838,I560869,I560886,I560931,I560948,I560965,I560996,I561022,I561030,I561061,I561078,I561095,I561121,I561129,I561146,I561235,I561261,I561278,I561286,I561331,I561348,I561365,I561382,I561399,I561416,I561433,I561464,I561481,I561526,I561543,I561560,I561591,I561617,I561625,I561656,I561673,I561690,I561716,I561724,I561741,I561830,I561856,I561873,I561881,I561926,I561943,I561960,I561977,I561994,I562011,I562028,I562059,I562076,I562121,I562138,I562155,I562186,I562212,I562220,I562251,I562268,I562285,I562311,I562319,I562336,I562425,I562451,I562468,I562476,I562521,I562538,I562555,I562572,I562589,I562606,I562623,I562654,I562671,I562716,I562733,I562750,I562781,I562807,I562815,I562846,I562863,I562880,I562906,I562914,I562931,I563020,I563046,I563063,I563071,I563116,I563133,I563150,I563167,I563184,I563201,I563218,I563249,I563266,I563311,I563328,I563345,I563376,I563402,I563410,I563441,I563458,I563475,I563501,I563509,I563526,I563615,I563641,I563658,I563666,I563711,I563728,I563745,I563762,I563779,I563796,I563813,I563844,I563861,I563906,I563923,I563940,I563971,I563997,I564005,I564036,I564053,I564070,I564096,I564104,I564121,I564210,I564236,I564253,I564261,I564306,I564323,I564340,I564357,I564374,I564391,I564408,I564439,I564456,I564501,I564518,I564535,I564566,I564592,I564600,I564631,I564648,I564665,I564691,I564699,I564716,I564805,I564831,I564848,I564856,I564901,I564918,I564935,I564952,I564969,I564986,I565003,I565034,I565051,I565096,I565113,I565130,I565161,I565187,I565195,I565226,I565243,I565260,I565286,I565294,I565311,I565400,I565426,I565443,I565451,I565496,I565513,I565530,I565547,I565564,I565581,I565598,I565629,I565646,I565691,I565708,I565725,I565756,I565782,I565790,I565821,I565838,I565855,I565881,I565889,I565906,I565995,I566021,I566038,I566046,I566091,I566108,I566125,I566142,I566159,I566176,I566193,I566224,I566241,I566286,I566303,I566320,I566351,I566377,I566385,I566416,I566433,I566450,I566476,I566484,I566501,I566590,I566616,I566633,I566641,I566686,I566703,I566720,I566737,I566754,I566771,I566788,I566819,I566836,I566881,I566898,I566915,I566946,I566972,I566980,I567011,I567028,I567045,I567071,I567079,I567096,I567185,I567211,I567228,I567236,I567281,I567298,I567315,I567332,I567349,I567366,I567383,I567414,I567431,I567476,I567493,I567510,I567541,I567567,I567575,I567606,I567623,I567640,I567666,I567674,I567691,I567780,I567806,I567823,I567831,I567876,I567893,I567910,I567927,I567944,I567961,I567978,I568009,I568026,I568071,I568088,I568105,I568136,I568162,I568170,I568201,I568218,I568235,I568261,I568269,I568286,I568375,I568401,I568418,I568426,I568471,I568488,I568505,I568522,I568539,I568556,I568573,I568604,I568621,I568666,I568683,I568700,I568731,I568757,I568765,I568796,I568813,I568830,I568856,I568864,I568881,I568970,I568996,I569013,I569021,I569066,I569083,I569100,I569117,I569134,I569151,I569168,I569199,I569216,I569261,I569278,I569295,I569326,I569352,I569360,I569391,I569408,I569425,I569451,I569459,I569476,I569565,I569591,I569608,I569616,I569661,I569678,I569695,I569712,I569729,I569746,I569763,I569794,I569811,I569856,I569873,I569890,I569921,I569947,I569955,I569986,I570003,I570020,I570046,I570054,I570071,I570160,I570186,I570203,I570211,I570256,I570273,I570290,I570307,I570324,I570341,I570358,I570389,I570406,I570451,I570468,I570485,I570516,I570542,I570550,I570581,I570598,I570615,I570641,I570649,I570666,I570755,I570781,I570798,I570806,I570851,I570868,I570885,I570902,I570919,I570936,I570953,I570984,I571001,I571046,I571063,I571080,I571111,I571137,I571145,I571176,I571193,I571210,I571236,I571244,I571261,I571350,I571376,I571393,I571401,I571446,I571463,I571480,I571497,I571514,I571531,I571548,I571579,I571596,I571641,I571658,I571675,I571706,I571732,I571740,I571771,I571788,I571805,I571831,I571839,I571856,I571945,I571971,I571988,I571996,I572041,I572058,I572075,I572092,I572109,I572126,I572143,I572174,I572191,I572236,I572253,I572270,I572301,I572327,I572335,I572366,I572383,I572400,I572426,I572434,I572451,I572540,I572566,I572583,I572591,I572636,I572653,I572670,I572687,I572704,I572721,I572738,I572769,I572786,I572831,I572848,I572865,I572896,I572922,I572930,I572961,I572978,I572995,I573021,I573029,I573046,I573135,I573161,I573178,I573186,I573231,I573248,I573265,I573282,I573299,I573316,I573333,I573364,I573381,I573426,I573443,I573460,I573491,I573517,I573525,I573556,I573573,I573590,I573616,I573624,I573641,I573730,I573756,I573773,I573781,I573826,I573843,I573860,I573877,I573894,I573911,I573928,I573959,I573976,I574021,I574038,I574055,I574086,I574112,I574120,I574151,I574168,I574185,I574211,I574219,I574236;
not I_0 (I2898,I2866);
DFFARX1 I_1 (I92955,I2859,I2898,I2924,);
nand I_2 (I2932,I2924,I92955);
not I_3 (I2949,I2932);
DFFARX1 I_4 (I2949,I2859,I2898,I2890,);
DFFARX1 I_5 (I92961,I2859,I2898,I2989,);
not I_6 (I2997,I2989);
not I_7 (I3014,I92970);
not I_8 (I3031,I92964);
nand I_9 (I3048,I2997,I3031);
nor I_10 (I3065,I3048,I92970);
DFFARX1 I_11 (I3065,I2859,I2898,I2869,);
nor I_12 (I3096,I92964,I92970);
nand I_13 (I3113,I2989,I3096);
nor I_14 (I3130,I92967,I92973);
nor I_15 (I2872,I3048,I92967);
not I_16 (I3161,I92967);
not I_17 (I3178,I92976);
nand I_18 (I3195,I3178,I92952);
nand I_19 (I3212,I3014,I3195);
not I_20 (I3229,I3212);
nor I_21 (I3246,I92976,I92973);
nor I_22 (I2881,I3229,I3246);
nor I_23 (I3277,I92958,I92976);
and I_24 (I3294,I3277,I3130);
nor I_25 (I3311,I3212,I3294);
DFFARX1 I_26 (I3311,I2859,I2898,I2887,);
nor I_27 (I3342,I2932,I3294);
DFFARX1 I_28 (I3342,I2859,I2898,I2884,);
nor I_29 (I3373,I92958,I92952);
DFFARX1 I_30 (I3373,I2859,I2898,I3399,);
nor I_31 (I3407,I3399,I92964);
nand I_32 (I3424,I3407,I3014);
nand I_33 (I2878,I3424,I3113);
nand I_34 (I2875,I3407,I3161);
not I_35 (I3493,I2866);
DFFARX1 I_36 (I411570,I2859,I3493,I3519,);
nand I_37 (I3527,I3519,I411561);
not I_38 (I3544,I3527);
DFFARX1 I_39 (I3544,I2859,I3493,I3485,);
DFFARX1 I_40 (I411564,I2859,I3493,I3584,);
not I_41 (I3592,I3584);
not I_42 (I3609,I411576);
not I_43 (I3626,I411555);
nand I_44 (I3643,I3592,I3626);
nor I_45 (I3660,I3643,I411576);
DFFARX1 I_46 (I3660,I2859,I3493,I3464,);
nor I_47 (I3691,I411555,I411576);
nand I_48 (I3708,I3584,I3691);
nor I_49 (I3725,I411567,I411573);
nor I_50 (I3467,I3643,I411567);
not I_51 (I3756,I411567);
not I_52 (I3773,I411558);
nand I_53 (I3790,I3773,I411549);
nand I_54 (I3807,I3609,I3790);
not I_55 (I3824,I3807);
nor I_56 (I3841,I411558,I411573);
nor I_57 (I3476,I3824,I3841);
nor I_58 (I3872,I411549,I411558);
and I_59 (I3889,I3872,I3725);
nor I_60 (I3906,I3807,I3889);
DFFARX1 I_61 (I3906,I2859,I3493,I3482,);
nor I_62 (I3937,I3527,I3889);
DFFARX1 I_63 (I3937,I2859,I3493,I3479,);
nor I_64 (I3968,I411549,I411552);
DFFARX1 I_65 (I3968,I2859,I3493,I3994,);
nor I_66 (I4002,I3994,I411555);
nand I_67 (I4019,I4002,I3609);
nand I_68 (I3473,I4019,I3708);
nand I_69 (I3470,I4002,I3756);
not I_70 (I4088,I2866);
DFFARX1 I_71 (I536225,I2859,I4088,I4114,);
nand I_72 (I4122,I4114,I536216);
not I_73 (I4139,I4122);
DFFARX1 I_74 (I4139,I2859,I4088,I4080,);
DFFARX1 I_75 (I536219,I2859,I4088,I4179,);
not I_76 (I4187,I4179);
not I_77 (I4204,I536231);
not I_78 (I4221,I536222);
nand I_79 (I4238,I4187,I4221);
nor I_80 (I4255,I4238,I536231);
DFFARX1 I_81 (I4255,I2859,I4088,I4059,);
nor I_82 (I4286,I536222,I536231);
nand I_83 (I4303,I4179,I4286);
nor I_84 (I4320,I536210,I536210);
nor I_85 (I4062,I4238,I536210);
not I_86 (I4351,I536210);
not I_87 (I4368,I536234);
nand I_88 (I4385,I4368,I536213);
nand I_89 (I4402,I4204,I4385);
not I_90 (I4419,I4402);
nor I_91 (I4436,I536234,I536210);
nor I_92 (I4071,I4419,I4436);
nor I_93 (I4467,I536228,I536234);
and I_94 (I4484,I4467,I4320);
nor I_95 (I4501,I4402,I4484);
DFFARX1 I_96 (I4501,I2859,I4088,I4077,);
nor I_97 (I4532,I4122,I4484);
DFFARX1 I_98 (I4532,I2859,I4088,I4074,);
nor I_99 (I4563,I536228,I536237);
DFFARX1 I_100 (I4563,I2859,I4088,I4589,);
nor I_101 (I4597,I4589,I536222);
nand I_102 (I4614,I4597,I4204);
nand I_103 (I4068,I4614,I4303);
nand I_104 (I4065,I4597,I4351);
not I_105 (I4683,I2866);
DFFARX1 I_106 (I176749,I2859,I4683,I4709,);
nand I_107 (I4717,I4709,I176731);
not I_108 (I4734,I4717);
DFFARX1 I_109 (I4734,I2859,I4683,I4675,);
DFFARX1 I_110 (I176743,I2859,I4683,I4774,);
not I_111 (I4782,I4774);
not I_112 (I4799,I176728);
not I_113 (I4816,I176737);
nand I_114 (I4833,I4782,I4816);
nor I_115 (I4850,I4833,I176728);
DFFARX1 I_116 (I4850,I2859,I4683,I4654,);
nor I_117 (I4881,I176737,I176728);
nand I_118 (I4898,I4774,I4881);
nor I_119 (I4915,I176734,I176755);
nor I_120 (I4657,I4833,I176734);
not I_121 (I4946,I176734);
not I_122 (I4963,I176746);
nand I_123 (I4980,I4963,I176752);
nand I_124 (I4997,I4799,I4980);
not I_125 (I5014,I4997);
nor I_126 (I5031,I176746,I176755);
nor I_127 (I4666,I5014,I5031);
nor I_128 (I5062,I176728,I176746);
and I_129 (I5079,I5062,I4915);
nor I_130 (I5096,I4997,I5079);
DFFARX1 I_131 (I5096,I2859,I4683,I4672,);
nor I_132 (I5127,I4717,I5079);
DFFARX1 I_133 (I5127,I2859,I4683,I4669,);
nor I_134 (I5158,I176728,I176740);
DFFARX1 I_135 (I5158,I2859,I4683,I5184,);
nor I_136 (I5192,I5184,I176737);
nand I_137 (I5209,I5192,I4799);
nand I_138 (I4663,I5209,I4898);
nand I_139 (I4660,I5192,I4946);
not I_140 (I5278,I2866);
DFFARX1 I_141 (I184909,I2859,I5278,I5304,);
nand I_142 (I5312,I5304,I184891);
not I_143 (I5329,I5312);
DFFARX1 I_144 (I5329,I2859,I5278,I5270,);
DFFARX1 I_145 (I184903,I2859,I5278,I5369,);
not I_146 (I5377,I5369);
not I_147 (I5394,I184888);
not I_148 (I5411,I184897);
nand I_149 (I5428,I5377,I5411);
nor I_150 (I5445,I5428,I184888);
DFFARX1 I_151 (I5445,I2859,I5278,I5249,);
nor I_152 (I5476,I184897,I184888);
nand I_153 (I5493,I5369,I5476);
nor I_154 (I5510,I184894,I184915);
nor I_155 (I5252,I5428,I184894);
not I_156 (I5541,I184894);
not I_157 (I5558,I184906);
nand I_158 (I5575,I5558,I184912);
nand I_159 (I5592,I5394,I5575);
not I_160 (I5609,I5592);
nor I_161 (I5626,I184906,I184915);
nor I_162 (I5261,I5609,I5626);
nor I_163 (I5657,I184888,I184906);
and I_164 (I5674,I5657,I5510);
nor I_165 (I5691,I5592,I5674);
DFFARX1 I_166 (I5691,I2859,I5278,I5267,);
nor I_167 (I5722,I5312,I5674);
DFFARX1 I_168 (I5722,I2859,I5278,I5264,);
nor I_169 (I5753,I184888,I184900);
DFFARX1 I_170 (I5753,I2859,I5278,I5779,);
nor I_171 (I5787,I5779,I184897);
nand I_172 (I5804,I5787,I5394);
nand I_173 (I5258,I5804,I5493);
nand I_174 (I5255,I5787,I5541);
not I_175 (I5876,I2866);
DFFARX1 I_176 (I529323,I2859,I5876,I5902,);
DFFARX1 I_177 (I5902,I2859,I5876,I5919,);
not I_178 (I5927,I5919);
nand I_179 (I5944,I529326,I529320);
and I_180 (I5961,I5944,I529329);
DFFARX1 I_181 (I5961,I2859,I5876,I5987,);
DFFARX1 I_182 (I5987,I2859,I5876,I5868,);
DFFARX1 I_183 (I5987,I2859,I5876,I5859,);
DFFARX1 I_184 (I529317,I2859,I5876,I6032,);
nand I_185 (I6040,I6032,I529332);
not I_186 (I6057,I6040);
nor I_187 (I5856,I5902,I6057);
DFFARX1 I_188 (I529308,I2859,I5876,I6097,);
not I_189 (I6105,I6097);
nor I_190 (I5862,I6105,I5927);
nand I_191 (I5850,I6105,I6040);
nand I_192 (I6150,I529311,I529311);
and I_193 (I6167,I6150,I529308);
DFFARX1 I_194 (I6167,I2859,I5876,I6193,);
nor I_195 (I6201,I6193,I5902);
DFFARX1 I_196 (I6201,I2859,I5876,I5844,);
not I_197 (I6232,I6193);
nor I_198 (I6249,I529314,I529311);
not I_199 (I6266,I6249);
nor I_200 (I6283,I6040,I6266);
nor I_201 (I6300,I6232,I6283);
DFFARX1 I_202 (I6300,I2859,I5876,I5865,);
nor I_203 (I6331,I6193,I6266);
nor I_204 (I5853,I6057,I6331);
nor I_205 (I5847,I6193,I6249);
not I_206 (I6403,I2866);
DFFARX1 I_207 (I288016,I2859,I6403,I6429,);
DFFARX1 I_208 (I6429,I2859,I6403,I6446,);
not I_209 (I6454,I6446);
nand I_210 (I6471,I288031,I288034);
and I_211 (I6488,I6471,I288013);
DFFARX1 I_212 (I6488,I2859,I6403,I6514,);
DFFARX1 I_213 (I6514,I2859,I6403,I6395,);
DFFARX1 I_214 (I6514,I2859,I6403,I6386,);
DFFARX1 I_215 (I288019,I2859,I6403,I6559,);
nand I_216 (I6567,I6559,I288025);
not I_217 (I6584,I6567);
nor I_218 (I6383,I6429,I6584);
DFFARX1 I_219 (I288013,I2859,I6403,I6624,);
not I_220 (I6632,I6624);
nor I_221 (I6389,I6632,I6454);
nand I_222 (I6377,I6632,I6567);
nand I_223 (I6677,I288028,I288010);
and I_224 (I6694,I6677,I288022);
DFFARX1 I_225 (I6694,I2859,I6403,I6720,);
nor I_226 (I6728,I6720,I6429);
DFFARX1 I_227 (I6728,I2859,I6403,I6371,);
not I_228 (I6759,I6720);
nor I_229 (I6776,I288010,I288010);
not I_230 (I6793,I6776);
nor I_231 (I6810,I6567,I6793);
nor I_232 (I6827,I6759,I6810);
DFFARX1 I_233 (I6827,I2859,I6403,I6392,);
nor I_234 (I6858,I6720,I6793);
nor I_235 (I6380,I6584,I6858);
nor I_236 (I6374,I6720,I6776);
not I_237 (I6930,I2866);
DFFARX1 I_238 (I195768,I2859,I6930,I6956,);
DFFARX1 I_239 (I6956,I2859,I6930,I6973,);
not I_240 (I6981,I6973);
nand I_241 (I6998,I195768,I195771);
and I_242 (I7015,I6998,I195792);
DFFARX1 I_243 (I7015,I2859,I6930,I7041,);
DFFARX1 I_244 (I7041,I2859,I6930,I6922,);
DFFARX1 I_245 (I7041,I2859,I6930,I6913,);
DFFARX1 I_246 (I195780,I2859,I6930,I7086,);
nand I_247 (I7094,I7086,I195783);
not I_248 (I7111,I7094);
nor I_249 (I6910,I6956,I7111);
DFFARX1 I_250 (I195789,I2859,I6930,I7151,);
not I_251 (I7159,I7151);
nor I_252 (I6916,I7159,I6981);
nand I_253 (I6904,I7159,I7094);
nand I_254 (I7204,I195786,I195774);
and I_255 (I7221,I7204,I195777);
DFFARX1 I_256 (I7221,I2859,I6930,I7247,);
nor I_257 (I7255,I7247,I6956);
DFFARX1 I_258 (I7255,I2859,I6930,I6898,);
not I_259 (I7286,I7247);
nor I_260 (I7303,I195795,I195774);
not I_261 (I7320,I7303);
nor I_262 (I7337,I7094,I7320);
nor I_263 (I7354,I7286,I7337);
DFFARX1 I_264 (I7354,I2859,I6930,I6919,);
nor I_265 (I7385,I7247,I7320);
nor I_266 (I6907,I7111,I7385);
nor I_267 (I6901,I7247,I7303);
not I_268 (I7457,I2866);
DFFARX1 I_269 (I496148,I2859,I7457,I7483,);
DFFARX1 I_270 (I7483,I2859,I7457,I7500,);
not I_271 (I7508,I7500);
nand I_272 (I7525,I496136,I496127);
and I_273 (I7542,I7525,I496124);
DFFARX1 I_274 (I7542,I2859,I7457,I7568,);
DFFARX1 I_275 (I7568,I2859,I7457,I7449,);
DFFARX1 I_276 (I7568,I2859,I7457,I7440,);
DFFARX1 I_277 (I496130,I2859,I7457,I7613,);
nand I_278 (I7621,I7613,I496142);
not I_279 (I7638,I7621);
nor I_280 (I7437,I7483,I7638);
DFFARX1 I_281 (I496139,I2859,I7457,I7678,);
not I_282 (I7686,I7678);
nor I_283 (I7443,I7686,I7508);
nand I_284 (I7431,I7686,I7621);
nand I_285 (I7731,I496133,I496127);
and I_286 (I7748,I7731,I496145);
DFFARX1 I_287 (I7748,I2859,I7457,I7774,);
nor I_288 (I7782,I7774,I7483);
DFFARX1 I_289 (I7782,I2859,I7457,I7425,);
not I_290 (I7813,I7774);
nor I_291 (I7830,I496124,I496127);
not I_292 (I7847,I7830);
nor I_293 (I7864,I7621,I7847);
nor I_294 (I7881,I7813,I7864);
DFFARX1 I_295 (I7881,I2859,I7457,I7446,);
nor I_296 (I7912,I7774,I7847);
nor I_297 (I7434,I7638,I7912);
nor I_298 (I7428,I7774,I7830);
not I_299 (I7984,I2866);
DFFARX1 I_300 (I207864,I2859,I7984,I8010,);
DFFARX1 I_301 (I8010,I2859,I7984,I8027,);
not I_302 (I8035,I8027);
nand I_303 (I8052,I207870,I207858);
and I_304 (I8069,I8052,I207855);
DFFARX1 I_305 (I8069,I2859,I7984,I8095,);
DFFARX1 I_306 (I8095,I2859,I7984,I7976,);
DFFARX1 I_307 (I8095,I2859,I7984,I7967,);
DFFARX1 I_308 (I207867,I2859,I7984,I8140,);
nand I_309 (I8148,I8140,I207861);
not I_310 (I8165,I8148);
nor I_311 (I7964,I8010,I8165);
DFFARX1 I_312 (I207879,I2859,I7984,I8205,);
not I_313 (I8213,I8205);
nor I_314 (I7970,I8213,I8035);
nand I_315 (I7958,I8213,I8148);
nand I_316 (I8258,I207873,I207876);
and I_317 (I8275,I8258,I207858);
DFFARX1 I_318 (I8275,I2859,I7984,I8301,);
nor I_319 (I8309,I8301,I8010);
DFFARX1 I_320 (I8309,I2859,I7984,I7952,);
not I_321 (I8340,I8301);
nor I_322 (I8357,I207855,I207876);
not I_323 (I8374,I8357);
nor I_324 (I8391,I8148,I8374);
nor I_325 (I8408,I8340,I8391);
DFFARX1 I_326 (I8408,I2859,I7984,I7973,);
nor I_327 (I8439,I8301,I8374);
nor I_328 (I7961,I8165,I8439);
nor I_329 (I7955,I8301,I8357);
not I_330 (I8511,I2866);
DFFARX1 I_331 (I281658,I2859,I8511,I8537,);
DFFARX1 I_332 (I8537,I2859,I8511,I8554,);
not I_333 (I8562,I8554);
nand I_334 (I8579,I281673,I281676);
and I_335 (I8596,I8579,I281655);
DFFARX1 I_336 (I8596,I2859,I8511,I8622,);
DFFARX1 I_337 (I8622,I2859,I8511,I8503,);
DFFARX1 I_338 (I8622,I2859,I8511,I8494,);
DFFARX1 I_339 (I281661,I2859,I8511,I8667,);
nand I_340 (I8675,I8667,I281667);
not I_341 (I8692,I8675);
nor I_342 (I8491,I8537,I8692);
DFFARX1 I_343 (I281655,I2859,I8511,I8732,);
not I_344 (I8740,I8732);
nor I_345 (I8497,I8740,I8562);
nand I_346 (I8485,I8740,I8675);
nand I_347 (I8785,I281670,I281652);
and I_348 (I8802,I8785,I281664);
DFFARX1 I_349 (I8802,I2859,I8511,I8828,);
nor I_350 (I8836,I8828,I8537);
DFFARX1 I_351 (I8836,I2859,I8511,I8479,);
not I_352 (I8867,I8828);
nor I_353 (I8884,I281652,I281652);
not I_354 (I8901,I8884);
nor I_355 (I8918,I8675,I8901);
nor I_356 (I8935,I8867,I8918);
DFFARX1 I_357 (I8935,I2859,I8511,I8500,);
nor I_358 (I8966,I8828,I8901);
nor I_359 (I8488,I8692,I8966);
nor I_360 (I8482,I8828,I8884);
not I_361 (I9038,I2866);
DFFARX1 I_362 (I101883,I2859,I9038,I9064,);
DFFARX1 I_363 (I9064,I2859,I9038,I9081,);
not I_364 (I9089,I9081);
nand I_365 (I9106,I101901,I101886);
and I_366 (I9123,I9106,I101889);
DFFARX1 I_367 (I9123,I2859,I9038,I9149,);
DFFARX1 I_368 (I9149,I2859,I9038,I9030,);
DFFARX1 I_369 (I9149,I2859,I9038,I9021,);
DFFARX1 I_370 (I101877,I2859,I9038,I9194,);
nand I_371 (I9202,I9194,I101880);
not I_372 (I9219,I9202);
nor I_373 (I9018,I9064,I9219);
DFFARX1 I_374 (I101892,I2859,I9038,I9259,);
not I_375 (I9267,I9259);
nor I_376 (I9024,I9267,I9089);
nand I_377 (I9012,I9267,I9202);
nand I_378 (I9312,I101898,I101895);
and I_379 (I9329,I9312,I101880);
DFFARX1 I_380 (I9329,I2859,I9038,I9355,);
nor I_381 (I9363,I9355,I9064);
DFFARX1 I_382 (I9363,I2859,I9038,I9006,);
not I_383 (I9394,I9355);
nor I_384 (I9411,I101877,I101895);
not I_385 (I9428,I9411);
nor I_386 (I9445,I9202,I9428);
nor I_387 (I9462,I9394,I9445);
DFFARX1 I_388 (I9462,I2859,I9038,I9027,);
nor I_389 (I9493,I9355,I9428);
nor I_390 (I9015,I9219,I9493);
nor I_391 (I9009,I9355,I9411);
not I_392 (I9565,I2866);
DFFARX1 I_393 (I253923,I2859,I9565,I9591,);
DFFARX1 I_394 (I9591,I2859,I9565,I9608,);
not I_395 (I9616,I9608);
nand I_396 (I9633,I253908,I253926);
and I_397 (I9650,I9633,I253920);
DFFARX1 I_398 (I9650,I2859,I9565,I9676,);
DFFARX1 I_399 (I9676,I2859,I9565,I9557,);
DFFARX1 I_400 (I9676,I2859,I9565,I9548,);
DFFARX1 I_401 (I253917,I2859,I9565,I9721,);
nand I_402 (I9729,I9721,I253908);
not I_403 (I9746,I9729);
nor I_404 (I9545,I9591,I9746);
DFFARX1 I_405 (I253911,I2859,I9565,I9786,);
not I_406 (I9794,I9786);
nor I_407 (I9551,I9794,I9616);
nand I_408 (I9539,I9794,I9729);
nand I_409 (I9839,I253932,I253914);
and I_410 (I9856,I9839,I253929);
DFFARX1 I_411 (I9856,I2859,I9565,I9882,);
nor I_412 (I9890,I9882,I9591);
DFFARX1 I_413 (I9890,I2859,I9565,I9533,);
not I_414 (I9921,I9882);
nor I_415 (I9938,I253911,I253914);
not I_416 (I9955,I9938);
nor I_417 (I9972,I9729,I9955);
nor I_418 (I9989,I9921,I9972);
DFFARX1 I_419 (I9989,I2859,I9565,I9554,);
nor I_420 (I10020,I9882,I9955);
nor I_421 (I9542,I9746,I10020);
nor I_422 (I9536,I9882,I9938);
not I_423 (I10092,I2866);
DFFARX1 I_424 (I331777,I2859,I10092,I10118,);
DFFARX1 I_425 (I10118,I2859,I10092,I10135,);
not I_426 (I10143,I10135);
nand I_427 (I10160,I331768,I331789);
and I_428 (I10177,I10160,I331771);
DFFARX1 I_429 (I10177,I2859,I10092,I10203,);
DFFARX1 I_430 (I10203,I2859,I10092,I10084,);
DFFARX1 I_431 (I10203,I2859,I10092,I10075,);
DFFARX1 I_432 (I331771,I2859,I10092,I10248,);
nand I_433 (I10256,I10248,I331786);
not I_434 (I10273,I10256);
nor I_435 (I10072,I10118,I10273);
DFFARX1 I_436 (I331780,I2859,I10092,I10313,);
not I_437 (I10321,I10313);
nor I_438 (I10078,I10321,I10143);
nand I_439 (I10066,I10321,I10256);
nand I_440 (I10366,I331774,I331783);
and I_441 (I10383,I10366,I331768);
DFFARX1 I_442 (I10383,I2859,I10092,I10409,);
nor I_443 (I10417,I10409,I10118);
DFFARX1 I_444 (I10417,I2859,I10092,I10060,);
not I_445 (I10448,I10409);
nor I_446 (I10465,I331774,I331783);
not I_447 (I10482,I10465);
nor I_448 (I10499,I10256,I10482);
nor I_449 (I10516,I10448,I10499);
DFFARX1 I_450 (I10516,I2859,I10092,I10081,);
nor I_451 (I10547,I10409,I10482);
nor I_452 (I10069,I10273,I10547);
nor I_453 (I10063,I10409,I10465);
not I_454 (I10619,I2866);
DFFARX1 I_455 (I535615,I2859,I10619,I10645,);
DFFARX1 I_456 (I10645,I2859,I10619,I10662,);
not I_457 (I10670,I10662);
nand I_458 (I10687,I535618,I535624);
and I_459 (I10704,I10687,I535633);
DFFARX1 I_460 (I10704,I2859,I10619,I10730,);
DFFARX1 I_461 (I10730,I2859,I10619,I10611,);
DFFARX1 I_462 (I10730,I2859,I10619,I10602,);
DFFARX1 I_463 (I535636,I2859,I10619,I10775,);
nand I_464 (I10783,I10775,I535627);
not I_465 (I10800,I10783);
nor I_466 (I10599,I10645,I10800);
DFFARX1 I_467 (I535615,I2859,I10619,I10840,);
not I_468 (I10848,I10840);
nor I_469 (I10605,I10848,I10670);
nand I_470 (I10593,I10848,I10783);
nand I_471 (I10893,I535642,I535621);
and I_472 (I10910,I10893,I535630);
DFFARX1 I_473 (I10910,I2859,I10619,I10936,);
nor I_474 (I10944,I10936,I10645);
DFFARX1 I_475 (I10944,I2859,I10619,I10587,);
not I_476 (I10975,I10936);
nor I_477 (I10992,I535639,I535621);
not I_478 (I11009,I10992);
nor I_479 (I11026,I10783,I11009);
nor I_480 (I11043,I10975,I11026);
DFFARX1 I_481 (I11043,I2859,I10619,I10608,);
nor I_482 (I11074,I10936,I11009);
nor I_483 (I10596,I10800,I11074);
nor I_484 (I10590,I10936,I10992);
not I_485 (I11146,I2866);
DFFARX1 I_486 (I456844,I2859,I11146,I11172,);
DFFARX1 I_487 (I11172,I2859,I11146,I11189,);
not I_488 (I11197,I11189);
nand I_489 (I11214,I456832,I456823);
and I_490 (I11231,I11214,I456820);
DFFARX1 I_491 (I11231,I2859,I11146,I11257,);
DFFARX1 I_492 (I11257,I2859,I11146,I11138,);
DFFARX1 I_493 (I11257,I2859,I11146,I11129,);
DFFARX1 I_494 (I456826,I2859,I11146,I11302,);
nand I_495 (I11310,I11302,I456838);
not I_496 (I11327,I11310);
nor I_497 (I11126,I11172,I11327);
DFFARX1 I_498 (I456835,I2859,I11146,I11367,);
not I_499 (I11375,I11367);
nor I_500 (I11132,I11375,I11197);
nand I_501 (I11120,I11375,I11310);
nand I_502 (I11420,I456829,I456823);
and I_503 (I11437,I11420,I456841);
DFFARX1 I_504 (I11437,I2859,I11146,I11463,);
nor I_505 (I11471,I11463,I11172);
DFFARX1 I_506 (I11471,I2859,I11146,I11114,);
not I_507 (I11502,I11463);
nor I_508 (I11519,I456820,I456823);
not I_509 (I11536,I11519);
nor I_510 (I11553,I11310,I11536);
nor I_511 (I11570,I11502,I11553);
DFFARX1 I_512 (I11570,I2859,I11146,I11135,);
nor I_513 (I11601,I11463,I11536);
nor I_514 (I11123,I11327,I11601);
nor I_515 (I11117,I11463,I11519);
not I_516 (I11673,I2866);
DFFARX1 I_517 (I341790,I2859,I11673,I11699,);
DFFARX1 I_518 (I11699,I2859,I11673,I11716,);
not I_519 (I11724,I11716);
nand I_520 (I11741,I341781,I341802);
and I_521 (I11758,I11741,I341784);
DFFARX1 I_522 (I11758,I2859,I11673,I11784,);
DFFARX1 I_523 (I11784,I2859,I11673,I11665,);
DFFARX1 I_524 (I11784,I2859,I11673,I11656,);
DFFARX1 I_525 (I341784,I2859,I11673,I11829,);
nand I_526 (I11837,I11829,I341799);
not I_527 (I11854,I11837);
nor I_528 (I11653,I11699,I11854);
DFFARX1 I_529 (I341793,I2859,I11673,I11894,);
not I_530 (I11902,I11894);
nor I_531 (I11659,I11902,I11724);
nand I_532 (I11647,I11902,I11837);
nand I_533 (I11947,I341787,I341796);
and I_534 (I11964,I11947,I341781);
DFFARX1 I_535 (I11964,I2859,I11673,I11990,);
nor I_536 (I11998,I11990,I11699);
DFFARX1 I_537 (I11998,I2859,I11673,I11641,);
not I_538 (I12029,I11990);
nor I_539 (I12046,I341787,I341796);
not I_540 (I12063,I12046);
nor I_541 (I12080,I11837,I12063);
nor I_542 (I12097,I12029,I12080);
DFFARX1 I_543 (I12097,I2859,I11673,I11662,);
nor I_544 (I12128,I11990,I12063);
nor I_545 (I11650,I11854,I12128);
nor I_546 (I11644,I11990,I12046);
not I_547 (I12200,I2866);
DFFARX1 I_548 (I206674,I2859,I12200,I12226,);
DFFARX1 I_549 (I12226,I2859,I12200,I12243,);
not I_550 (I12251,I12243);
nand I_551 (I12268,I206680,I206668);
and I_552 (I12285,I12268,I206665);
DFFARX1 I_553 (I12285,I2859,I12200,I12311,);
DFFARX1 I_554 (I12311,I2859,I12200,I12192,);
DFFARX1 I_555 (I12311,I2859,I12200,I12183,);
DFFARX1 I_556 (I206677,I2859,I12200,I12356,);
nand I_557 (I12364,I12356,I206671);
not I_558 (I12381,I12364);
nor I_559 (I12180,I12226,I12381);
DFFARX1 I_560 (I206689,I2859,I12200,I12421,);
not I_561 (I12429,I12421);
nor I_562 (I12186,I12429,I12251);
nand I_563 (I12174,I12429,I12364);
nand I_564 (I12474,I206683,I206686);
and I_565 (I12491,I12474,I206668);
DFFARX1 I_566 (I12491,I2859,I12200,I12517,);
nor I_567 (I12525,I12517,I12226);
DFFARX1 I_568 (I12525,I2859,I12200,I12168,);
not I_569 (I12556,I12517);
nor I_570 (I12573,I206665,I206686);
not I_571 (I12590,I12573);
nor I_572 (I12607,I12364,I12590);
nor I_573 (I12624,I12556,I12607);
DFFARX1 I_574 (I12624,I2859,I12200,I12189,);
nor I_575 (I12655,I12517,I12590);
nor I_576 (I12177,I12381,I12655);
nor I_577 (I12171,I12517,I12573);
not I_578 (I12727,I2866);
DFFARX1 I_579 (I163672,I2859,I12727,I12753,);
DFFARX1 I_580 (I12753,I2859,I12727,I12770,);
not I_581 (I12778,I12770);
nand I_582 (I12795,I163672,I163675);
and I_583 (I12812,I12795,I163696);
DFFARX1 I_584 (I12812,I2859,I12727,I12838,);
DFFARX1 I_585 (I12838,I2859,I12727,I12719,);
DFFARX1 I_586 (I12838,I2859,I12727,I12710,);
DFFARX1 I_587 (I163684,I2859,I12727,I12883,);
nand I_588 (I12891,I12883,I163687);
not I_589 (I12908,I12891);
nor I_590 (I12707,I12753,I12908);
DFFARX1 I_591 (I163693,I2859,I12727,I12948,);
not I_592 (I12956,I12948);
nor I_593 (I12713,I12956,I12778);
nand I_594 (I12701,I12956,I12891);
nand I_595 (I13001,I163690,I163678);
and I_596 (I13018,I13001,I163681);
DFFARX1 I_597 (I13018,I2859,I12727,I13044,);
nor I_598 (I13052,I13044,I12753);
DFFARX1 I_599 (I13052,I2859,I12727,I12695,);
not I_600 (I13083,I13044);
nor I_601 (I13100,I163699,I163678);
not I_602 (I13117,I13100);
nor I_603 (I13134,I12891,I13117);
nor I_604 (I13151,I13083,I13134);
DFFARX1 I_605 (I13151,I2859,I12727,I12716,);
nor I_606 (I13182,I13044,I13117);
nor I_607 (I12704,I12908,I13182);
nor I_608 (I12698,I13044,I13100);
not I_609 (I13254,I2866);
DFFARX1 I_610 (I338628,I2859,I13254,I13280,);
DFFARX1 I_611 (I13280,I2859,I13254,I13297,);
not I_612 (I13305,I13297);
nand I_613 (I13322,I338619,I338640);
and I_614 (I13339,I13322,I338622);
DFFARX1 I_615 (I13339,I2859,I13254,I13365,);
DFFARX1 I_616 (I13365,I2859,I13254,I13246,);
DFFARX1 I_617 (I13365,I2859,I13254,I13237,);
DFFARX1 I_618 (I338622,I2859,I13254,I13410,);
nand I_619 (I13418,I13410,I338637);
not I_620 (I13435,I13418);
nor I_621 (I13234,I13280,I13435);
DFFARX1 I_622 (I338631,I2859,I13254,I13475,);
not I_623 (I13483,I13475);
nor I_624 (I13240,I13483,I13305);
nand I_625 (I13228,I13483,I13418);
nand I_626 (I13528,I338625,I338634);
and I_627 (I13545,I13528,I338619);
DFFARX1 I_628 (I13545,I2859,I13254,I13571,);
nor I_629 (I13579,I13571,I13280);
DFFARX1 I_630 (I13579,I2859,I13254,I13222,);
not I_631 (I13610,I13571);
nor I_632 (I13627,I338625,I338634);
not I_633 (I13644,I13627);
nor I_634 (I13661,I13418,I13644);
nor I_635 (I13678,I13610,I13661);
DFFARX1 I_636 (I13678,I2859,I13254,I13243,);
nor I_637 (I13709,I13571,I13644);
nor I_638 (I13231,I13435,I13709);
nor I_639 (I13225,I13571,I13627);
not I_640 (I13781,I2866);
DFFARX1 I_641 (I272988,I2859,I13781,I13807,);
DFFARX1 I_642 (I13807,I2859,I13781,I13824,);
not I_643 (I13832,I13824);
nand I_644 (I13849,I273003,I273006);
and I_645 (I13866,I13849,I272985);
DFFARX1 I_646 (I13866,I2859,I13781,I13892,);
DFFARX1 I_647 (I13892,I2859,I13781,I13773,);
DFFARX1 I_648 (I13892,I2859,I13781,I13764,);
DFFARX1 I_649 (I272991,I2859,I13781,I13937,);
nand I_650 (I13945,I13937,I272997);
not I_651 (I13962,I13945);
nor I_652 (I13761,I13807,I13962);
DFFARX1 I_653 (I272985,I2859,I13781,I14002,);
not I_654 (I14010,I14002);
nor I_655 (I13767,I14010,I13832);
nand I_656 (I13755,I14010,I13945);
nand I_657 (I14055,I273000,I272982);
and I_658 (I14072,I14055,I272994);
DFFARX1 I_659 (I14072,I2859,I13781,I14098,);
nor I_660 (I14106,I14098,I13807);
DFFARX1 I_661 (I14106,I2859,I13781,I13749,);
not I_662 (I14137,I14098);
nor I_663 (I14154,I272982,I272982);
not I_664 (I14171,I14154);
nor I_665 (I14188,I13945,I14171);
nor I_666 (I14205,I14137,I14188);
DFFARX1 I_667 (I14205,I2859,I13781,I13770,);
nor I_668 (I14236,I14098,I14171);
nor I_669 (I13758,I13962,I14236);
nor I_670 (I13752,I14098,I14154);
not I_671 (I14308,I2866);
DFFARX1 I_672 (I188152,I2859,I14308,I14334,);
DFFARX1 I_673 (I14334,I2859,I14308,I14351,);
not I_674 (I14359,I14351);
nand I_675 (I14376,I188152,I188155);
and I_676 (I14393,I14376,I188176);
DFFARX1 I_677 (I14393,I2859,I14308,I14419,);
DFFARX1 I_678 (I14419,I2859,I14308,I14300,);
DFFARX1 I_679 (I14419,I2859,I14308,I14291,);
DFFARX1 I_680 (I188164,I2859,I14308,I14464,);
nand I_681 (I14472,I14464,I188167);
not I_682 (I14489,I14472);
nor I_683 (I14288,I14334,I14489);
DFFARX1 I_684 (I188173,I2859,I14308,I14529,);
not I_685 (I14537,I14529);
nor I_686 (I14294,I14537,I14359);
nand I_687 (I14282,I14537,I14472);
nand I_688 (I14582,I188170,I188158);
and I_689 (I14599,I14582,I188161);
DFFARX1 I_690 (I14599,I2859,I14308,I14625,);
nor I_691 (I14633,I14625,I14334);
DFFARX1 I_692 (I14633,I2859,I14308,I14276,);
not I_693 (I14664,I14625);
nor I_694 (I14681,I188179,I188158);
not I_695 (I14698,I14681);
nor I_696 (I14715,I14472,I14698);
nor I_697 (I14732,I14664,I14715);
DFFARX1 I_698 (I14732,I2859,I14308,I14297,);
nor I_699 (I14763,I14625,I14698);
nor I_700 (I14285,I14489,I14763);
nor I_701 (I14279,I14625,I14681);
not I_702 (I14835,I2866);
DFFARX1 I_703 (I404467,I2859,I14835,I14861,);
DFFARX1 I_704 (I14861,I2859,I14835,I14878,);
not I_705 (I14886,I14878);
nand I_706 (I14903,I404443,I404470);
and I_707 (I14920,I14903,I404455);
DFFARX1 I_708 (I14920,I2859,I14835,I14946,);
DFFARX1 I_709 (I14946,I2859,I14835,I14827,);
DFFARX1 I_710 (I14946,I2859,I14835,I14818,);
DFFARX1 I_711 (I404461,I2859,I14835,I14991,);
nand I_712 (I14999,I14991,I404446);
not I_713 (I15016,I14999);
nor I_714 (I14815,I14861,I15016);
DFFARX1 I_715 (I404464,I2859,I14835,I15056,);
not I_716 (I15064,I15056);
nor I_717 (I14821,I15064,I14886);
nand I_718 (I14809,I15064,I14999);
nand I_719 (I15109,I404449,I404452);
and I_720 (I15126,I15109,I404443);
DFFARX1 I_721 (I15126,I2859,I14835,I15152,);
nor I_722 (I15160,I15152,I14861);
DFFARX1 I_723 (I15160,I2859,I14835,I14803,);
not I_724 (I15191,I15152);
nor I_725 (I15208,I404458,I404452);
not I_726 (I15225,I15208);
nor I_727 (I15242,I14999,I15225);
nor I_728 (I15259,I15191,I15242);
DFFARX1 I_729 (I15259,I2859,I14835,I14824,);
nor I_730 (I15290,I15152,I15225);
nor I_731 (I14812,I15016,I15290);
nor I_732 (I14806,I15152,I15208);
not I_733 (I15362,I2866);
DFFARX1 I_734 (I256235,I2859,I15362,I15388,);
DFFARX1 I_735 (I15388,I2859,I15362,I15405,);
not I_736 (I15413,I15405);
nand I_737 (I15430,I256220,I256238);
and I_738 (I15447,I15430,I256232);
DFFARX1 I_739 (I15447,I2859,I15362,I15473,);
DFFARX1 I_740 (I15473,I2859,I15362,I15354,);
DFFARX1 I_741 (I15473,I2859,I15362,I15345,);
DFFARX1 I_742 (I256229,I2859,I15362,I15518,);
nand I_743 (I15526,I15518,I256220);
not I_744 (I15543,I15526);
nor I_745 (I15342,I15388,I15543);
DFFARX1 I_746 (I256223,I2859,I15362,I15583,);
not I_747 (I15591,I15583);
nor I_748 (I15348,I15591,I15413);
nand I_749 (I15336,I15591,I15526);
nand I_750 (I15636,I256244,I256226);
and I_751 (I15653,I15636,I256241);
DFFARX1 I_752 (I15653,I2859,I15362,I15679,);
nor I_753 (I15687,I15679,I15388);
DFFARX1 I_754 (I15687,I2859,I15362,I15330,);
not I_755 (I15718,I15679);
nor I_756 (I15735,I256223,I256226);
not I_757 (I15752,I15735);
nor I_758 (I15769,I15526,I15752);
nor I_759 (I15786,I15718,I15769);
DFFARX1 I_760 (I15786,I2859,I15362,I15351,);
nor I_761 (I15817,I15679,I15752);
nor I_762 (I15339,I15543,I15817);
nor I_763 (I15333,I15679,I15735);
not I_764 (I15889,I2866);
DFFARX1 I_765 (I353384,I2859,I15889,I15915,);
DFFARX1 I_766 (I15915,I2859,I15889,I15932,);
not I_767 (I15940,I15932);
nand I_768 (I15957,I353375,I353396);
and I_769 (I15974,I15957,I353378);
DFFARX1 I_770 (I15974,I2859,I15889,I16000,);
DFFARX1 I_771 (I16000,I2859,I15889,I15881,);
DFFARX1 I_772 (I16000,I2859,I15889,I15872,);
DFFARX1 I_773 (I353378,I2859,I15889,I16045,);
nand I_774 (I16053,I16045,I353393);
not I_775 (I16070,I16053);
nor I_776 (I15869,I15915,I16070);
DFFARX1 I_777 (I353387,I2859,I15889,I16110,);
not I_778 (I16118,I16110);
nor I_779 (I15875,I16118,I15940);
nand I_780 (I15863,I16118,I16053);
nand I_781 (I16163,I353381,I353390);
and I_782 (I16180,I16163,I353375);
DFFARX1 I_783 (I16180,I2859,I15889,I16206,);
nor I_784 (I16214,I16206,I15915);
DFFARX1 I_785 (I16214,I2859,I15889,I15857,);
not I_786 (I16245,I16206);
nor I_787 (I16262,I353381,I353390);
not I_788 (I16279,I16262);
nor I_789 (I16296,I16053,I16279);
nor I_790 (I16313,I16245,I16296);
DFFARX1 I_791 (I16313,I2859,I15889,I15878,);
nor I_792 (I16344,I16206,I16279);
nor I_793 (I15866,I16070,I16344);
nor I_794 (I15860,I16206,I16262);
not I_795 (I16416,I2866);
DFFARX1 I_796 (I4080,I2859,I16416,I16442,);
DFFARX1 I_797 (I16442,I2859,I16416,I16459,);
not I_798 (I16467,I16459);
nand I_799 (I16484,I4074,I4068);
and I_800 (I16501,I16484,I4065);
DFFARX1 I_801 (I16501,I2859,I16416,I16527,);
DFFARX1 I_802 (I16527,I2859,I16416,I16408,);
DFFARX1 I_803 (I16527,I2859,I16416,I16399,);
DFFARX1 I_804 (I4071,I2859,I16416,I16572,);
nand I_805 (I16580,I16572,I4065);
not I_806 (I16597,I16580);
nor I_807 (I16396,I16442,I16597);
DFFARX1 I_808 (I4062,I2859,I16416,I16637,);
not I_809 (I16645,I16637);
nor I_810 (I16402,I16645,I16467);
nand I_811 (I16390,I16645,I16580);
nand I_812 (I16690,I4059,I4059);
and I_813 (I16707,I16690,I4077);
DFFARX1 I_814 (I16707,I2859,I16416,I16733,);
nor I_815 (I16741,I16733,I16442);
DFFARX1 I_816 (I16741,I2859,I16416,I16384,);
not I_817 (I16772,I16733);
nor I_818 (I16789,I4062,I4059);
not I_819 (I16806,I16789);
nor I_820 (I16823,I16580,I16806);
nor I_821 (I16840,I16772,I16823);
DFFARX1 I_822 (I16840,I2859,I16416,I16405,);
nor I_823 (I16871,I16733,I16806);
nor I_824 (I16393,I16597,I16871);
nor I_825 (I16387,I16733,I16789);
not I_826 (I16943,I2866);
DFFARX1 I_827 (I524121,I2859,I16943,I16969,);
DFFARX1 I_828 (I16969,I2859,I16943,I16986,);
not I_829 (I16994,I16986);
nand I_830 (I17011,I524124,I524118);
and I_831 (I17028,I17011,I524127);
DFFARX1 I_832 (I17028,I2859,I16943,I17054,);
DFFARX1 I_833 (I17054,I2859,I16943,I16935,);
DFFARX1 I_834 (I17054,I2859,I16943,I16926,);
DFFARX1 I_835 (I524115,I2859,I16943,I17099,);
nand I_836 (I17107,I17099,I524130);
not I_837 (I17124,I17107);
nor I_838 (I16923,I16969,I17124);
DFFARX1 I_839 (I524106,I2859,I16943,I17164,);
not I_840 (I17172,I17164);
nor I_841 (I16929,I17172,I16994);
nand I_842 (I16917,I17172,I17107);
nand I_843 (I17217,I524109,I524109);
and I_844 (I17234,I17217,I524106);
DFFARX1 I_845 (I17234,I2859,I16943,I17260,);
nor I_846 (I17268,I17260,I16969);
DFFARX1 I_847 (I17268,I2859,I16943,I16911,);
not I_848 (I17299,I17260);
nor I_849 (I17316,I524112,I524109);
not I_850 (I17333,I17316);
nor I_851 (I17350,I17107,I17333);
nor I_852 (I17367,I17299,I17350);
DFFARX1 I_853 (I17367,I2859,I16943,I16932,);
nor I_854 (I17398,I17260,I17333);
nor I_855 (I16920,I17124,I17398);
nor I_856 (I16914,I17260,I17316);
not I_857 (I17470,I2866);
DFFARX1 I_858 (I96528,I2859,I17470,I17496,);
DFFARX1 I_859 (I17496,I2859,I17470,I17513,);
not I_860 (I17521,I17513);
nand I_861 (I17538,I96546,I96531);
and I_862 (I17555,I17538,I96534);
DFFARX1 I_863 (I17555,I2859,I17470,I17581,);
DFFARX1 I_864 (I17581,I2859,I17470,I17462,);
DFFARX1 I_865 (I17581,I2859,I17470,I17453,);
DFFARX1 I_866 (I96522,I2859,I17470,I17626,);
nand I_867 (I17634,I17626,I96525);
not I_868 (I17651,I17634);
nor I_869 (I17450,I17496,I17651);
DFFARX1 I_870 (I96537,I2859,I17470,I17691,);
not I_871 (I17699,I17691);
nor I_872 (I17456,I17699,I17521);
nand I_873 (I17444,I17699,I17634);
nand I_874 (I17744,I96543,I96540);
and I_875 (I17761,I17744,I96525);
DFFARX1 I_876 (I17761,I2859,I17470,I17787,);
nor I_877 (I17795,I17787,I17496);
DFFARX1 I_878 (I17795,I2859,I17470,I17438,);
not I_879 (I17826,I17787);
nor I_880 (I17843,I96522,I96540);
not I_881 (I17860,I17843);
nor I_882 (I17877,I17634,I17860);
nor I_883 (I17894,I17826,I17877);
DFFARX1 I_884 (I17894,I2859,I17470,I17459,);
nor I_885 (I17925,I17787,I17860);
nor I_886 (I17447,I17651,I17925);
nor I_887 (I17441,I17787,I17843);
not I_888 (I17997,I2866);
DFFARX1 I_889 (I227913,I2859,I17997,I18023,);
DFFARX1 I_890 (I18023,I2859,I17997,I18040,);
not I_891 (I18048,I18040);
nand I_892 (I18065,I227898,I227916);
and I_893 (I18082,I18065,I227910);
DFFARX1 I_894 (I18082,I2859,I17997,I18108,);
DFFARX1 I_895 (I18108,I2859,I17997,I17989,);
DFFARX1 I_896 (I18108,I2859,I17997,I17980,);
DFFARX1 I_897 (I227907,I2859,I17997,I18153,);
nand I_898 (I18161,I18153,I227898);
not I_899 (I18178,I18161);
nor I_900 (I17977,I18023,I18178);
DFFARX1 I_901 (I227901,I2859,I17997,I18218,);
not I_902 (I18226,I18218);
nor I_903 (I17983,I18226,I18048);
nand I_904 (I17971,I18226,I18161);
nand I_905 (I18271,I227922,I227904);
and I_906 (I18288,I18271,I227919);
DFFARX1 I_907 (I18288,I2859,I17997,I18314,);
nor I_908 (I18322,I18314,I18023);
DFFARX1 I_909 (I18322,I2859,I17997,I17965,);
not I_910 (I18353,I18314);
nor I_911 (I18370,I227901,I227904);
not I_912 (I18387,I18370);
nor I_913 (I18404,I18161,I18387);
nor I_914 (I18421,I18353,I18404);
DFFARX1 I_915 (I18421,I2859,I17997,I17986,);
nor I_916 (I18452,I18314,I18387);
nor I_917 (I17974,I18178,I18452);
nor I_918 (I17968,I18314,I18370);
not I_919 (I18524,I2866);
DFFARX1 I_920 (I222127,I2859,I18524,I18550,);
not I_921 (I18558,I18550);
nand I_922 (I18575,I222139,I222124);
and I_923 (I18592,I18575,I222118);
DFFARX1 I_924 (I18592,I2859,I18524,I18618,);
DFFARX1 I_925 (I222133,I2859,I18524,I18635,);
and I_926 (I18643,I18635,I222121);
nor I_927 (I18660,I18618,I18643);
DFFARX1 I_928 (I18660,I2859,I18524,I18492,);
nand I_929 (I18691,I18635,I222121);
nand I_930 (I18708,I18558,I18691);
not I_931 (I18504,I18708);
DFFARX1 I_932 (I222130,I2859,I18524,I18748,);
DFFARX1 I_933 (I18748,I2859,I18524,I18513,);
nand I_934 (I18770,I222136,I222142);
and I_935 (I18787,I18770,I222118);
DFFARX1 I_936 (I18787,I2859,I18524,I18813,);
DFFARX1 I_937 (I18813,I2859,I18524,I18830,);
not I_938 (I18516,I18830);
not I_939 (I18852,I18813);
nand I_940 (I18501,I18852,I18691);
nor I_941 (I18883,I222121,I222142);
not I_942 (I18900,I18883);
nor I_943 (I18917,I18852,I18900);
nor I_944 (I18934,I18558,I18917);
DFFARX1 I_945 (I18934,I2859,I18524,I18510,);
nor I_946 (I18965,I18618,I18900);
nor I_947 (I18498,I18813,I18965);
nor I_948 (I18507,I18748,I18883);
nor I_949 (I18495,I18618,I18883);
not I_950 (I19051,I2866);
DFFARX1 I_951 (I9030,I2859,I19051,I19077,);
not I_952 (I19085,I19077);
nand I_953 (I19102,I9018,I9024);
and I_954 (I19119,I19102,I9027);
DFFARX1 I_955 (I19119,I2859,I19051,I19145,);
DFFARX1 I_956 (I9009,I2859,I19051,I19162,);
and I_957 (I19170,I19162,I9015);
nor I_958 (I19187,I19145,I19170);
DFFARX1 I_959 (I19187,I2859,I19051,I19019,);
nand I_960 (I19218,I19162,I9015);
nand I_961 (I19235,I19085,I19218);
not I_962 (I19031,I19235);
DFFARX1 I_963 (I9009,I2859,I19051,I19275,);
DFFARX1 I_964 (I19275,I2859,I19051,I19040,);
nand I_965 (I19297,I9012,I9006);
and I_966 (I19314,I19297,I9021);
DFFARX1 I_967 (I19314,I2859,I19051,I19340,);
DFFARX1 I_968 (I19340,I2859,I19051,I19357,);
not I_969 (I19043,I19357);
not I_970 (I19379,I19340);
nand I_971 (I19028,I19379,I19218);
nor I_972 (I19410,I9006,I9006);
not I_973 (I19427,I19410);
nor I_974 (I19444,I19379,I19427);
nor I_975 (I19461,I19085,I19444);
DFFARX1 I_976 (I19461,I2859,I19051,I19037,);
nor I_977 (I19492,I19145,I19427);
nor I_978 (I19025,I19340,I19492);
nor I_979 (I19034,I19275,I19410);
nor I_980 (I19022,I19145,I19410);
not I_981 (I19578,I2866);
DFFARX1 I_982 (I328615,I2859,I19578,I19604,);
not I_983 (I19612,I19604);
nand I_984 (I19629,I328612,I328627);
and I_985 (I19646,I19629,I328609);
DFFARX1 I_986 (I19646,I2859,I19578,I19672,);
DFFARX1 I_987 (I328606,I2859,I19578,I19689,);
and I_988 (I19697,I19689,I328606);
nor I_989 (I19714,I19672,I19697);
DFFARX1 I_990 (I19714,I2859,I19578,I19546,);
nand I_991 (I19745,I19689,I328606);
nand I_992 (I19762,I19612,I19745);
not I_993 (I19558,I19762);
DFFARX1 I_994 (I328609,I2859,I19578,I19802,);
DFFARX1 I_995 (I19802,I2859,I19578,I19567,);
nand I_996 (I19824,I328621,I328612);
and I_997 (I19841,I19824,I328624);
DFFARX1 I_998 (I19841,I2859,I19578,I19867,);
DFFARX1 I_999 (I19867,I2859,I19578,I19884,);
not I_1000 (I19570,I19884);
not I_1001 (I19906,I19867);
nand I_1002 (I19555,I19906,I19745);
nor I_1003 (I19937,I328618,I328612);
not I_1004 (I19954,I19937);
nor I_1005 (I19971,I19906,I19954);
nor I_1006 (I19988,I19612,I19971);
DFFARX1 I_1007 (I19988,I2859,I19578,I19564,);
nor I_1008 (I20019,I19672,I19954);
nor I_1009 (I19552,I19867,I20019);
nor I_1010 (I19561,I19802,I19937);
nor I_1011 (I19549,I19672,I19937);
not I_1012 (I20105,I2866);
DFFARX1 I_1013 (I564782,I2859,I20105,I20131,);
not I_1014 (I20139,I20131);
nand I_1015 (I20156,I564776,I564797);
and I_1016 (I20173,I20156,I564773);
DFFARX1 I_1017 (I20173,I2859,I20105,I20199,);
DFFARX1 I_1018 (I564794,I2859,I20105,I20216,);
and I_1019 (I20224,I20216,I564791);
nor I_1020 (I20241,I20199,I20224);
DFFARX1 I_1021 (I20241,I2859,I20105,I20073,);
nand I_1022 (I20272,I20216,I564791);
nand I_1023 (I20289,I20139,I20272);
not I_1024 (I20085,I20289);
DFFARX1 I_1025 (I564779,I2859,I20105,I20329,);
DFFARX1 I_1026 (I20329,I2859,I20105,I20094,);
nand I_1027 (I20351,I564788,I564785);
and I_1028 (I20368,I20351,I564770);
DFFARX1 I_1029 (I20368,I2859,I20105,I20394,);
DFFARX1 I_1030 (I20394,I2859,I20105,I20411,);
not I_1031 (I20097,I20411);
not I_1032 (I20433,I20394);
nand I_1033 (I20082,I20433,I20272);
nor I_1034 (I20464,I564770,I564785);
not I_1035 (I20481,I20464);
nor I_1036 (I20498,I20433,I20481);
nor I_1037 (I20515,I20139,I20498);
DFFARX1 I_1038 (I20515,I2859,I20105,I20091,);
nor I_1039 (I20546,I20199,I20481);
nor I_1040 (I20079,I20394,I20546);
nor I_1041 (I20088,I20329,I20464);
nor I_1042 (I20076,I20199,I20464);
not I_1043 (I20632,I2866);
DFFARX1 I_1044 (I142517,I2859,I20632,I20658,);
not I_1045 (I20666,I20658);
nand I_1046 (I20683,I142499,I142514);
and I_1047 (I20700,I20683,I142490);
DFFARX1 I_1048 (I20700,I2859,I20632,I20726,);
DFFARX1 I_1049 (I142493,I2859,I20632,I20743,);
and I_1050 (I20751,I20743,I142508);
nor I_1051 (I20768,I20726,I20751);
DFFARX1 I_1052 (I20768,I2859,I20632,I20600,);
nand I_1053 (I20799,I20743,I142508);
nand I_1054 (I20816,I20666,I20799);
not I_1055 (I20612,I20816);
DFFARX1 I_1056 (I142511,I2859,I20632,I20856,);
DFFARX1 I_1057 (I20856,I2859,I20632,I20621,);
nand I_1058 (I20878,I142490,I142502);
and I_1059 (I20895,I20878,I142496);
DFFARX1 I_1060 (I20895,I2859,I20632,I20921,);
DFFARX1 I_1061 (I20921,I2859,I20632,I20938,);
not I_1062 (I20624,I20938);
not I_1063 (I20960,I20921);
nand I_1064 (I20609,I20960,I20799);
nor I_1065 (I20991,I142505,I142502);
not I_1066 (I21008,I20991);
nor I_1067 (I21025,I20960,I21008);
nor I_1068 (I21042,I20666,I21025);
DFFARX1 I_1069 (I21042,I2859,I20632,I20618,);
nor I_1070 (I21073,I20726,I21008);
nor I_1071 (I20606,I20921,I21073);
nor I_1072 (I20615,I20856,I20991);
nor I_1073 (I20603,I20726,I20991);
not I_1074 (I21159,I2866);
DFFARX1 I_1075 (I367630,I2859,I21159,I21185,);
not I_1076 (I21193,I21185);
nand I_1077 (I21210,I367648,I367642);
and I_1078 (I21227,I21210,I367621);
DFFARX1 I_1079 (I21227,I2859,I21159,I21253,);
DFFARX1 I_1080 (I367639,I2859,I21159,I21270,);
and I_1081 (I21278,I21270,I367624);
nor I_1082 (I21295,I21253,I21278);
DFFARX1 I_1083 (I21295,I2859,I21159,I21127,);
nand I_1084 (I21326,I21270,I367624);
nand I_1085 (I21343,I21193,I21326);
not I_1086 (I21139,I21343);
DFFARX1 I_1087 (I367636,I2859,I21159,I21383,);
DFFARX1 I_1088 (I21383,I2859,I21159,I21148,);
nand I_1089 (I21405,I367645,I367633);
and I_1090 (I21422,I21405,I367627);
DFFARX1 I_1091 (I21422,I2859,I21159,I21448,);
DFFARX1 I_1092 (I21448,I2859,I21159,I21465,);
not I_1093 (I21151,I21465);
not I_1094 (I21487,I21448);
nand I_1095 (I21136,I21487,I21326);
nor I_1096 (I21518,I367621,I367633);
not I_1097 (I21535,I21518);
nor I_1098 (I21552,I21487,I21535);
nor I_1099 (I21569,I21193,I21552);
DFFARX1 I_1100 (I21569,I2859,I21159,I21145,);
nor I_1101 (I21600,I21253,I21535);
nor I_1102 (I21133,I21448,I21600);
nor I_1103 (I21142,I21383,I21518);
nor I_1104 (I21130,I21253,I21518);
not I_1105 (I21686,I2866);
DFFARX1 I_1106 (I471854,I2859,I21686,I21712,);
not I_1107 (I21720,I21712);
nand I_1108 (I21737,I471869,I471848);
and I_1109 (I21754,I21737,I471851);
DFFARX1 I_1110 (I21754,I2859,I21686,I21780,);
DFFARX1 I_1111 (I471872,I2859,I21686,I21797,);
and I_1112 (I21805,I21797,I471851);
nor I_1113 (I21822,I21780,I21805);
DFFARX1 I_1114 (I21822,I2859,I21686,I21654,);
nand I_1115 (I21853,I21797,I471851);
nand I_1116 (I21870,I21720,I21853);
not I_1117 (I21666,I21870);
DFFARX1 I_1118 (I471848,I2859,I21686,I21910,);
DFFARX1 I_1119 (I21910,I2859,I21686,I21675,);
nand I_1120 (I21932,I471860,I471857);
and I_1121 (I21949,I21932,I471863);
DFFARX1 I_1122 (I21949,I2859,I21686,I21975,);
DFFARX1 I_1123 (I21975,I2859,I21686,I21992,);
not I_1124 (I21678,I21992);
not I_1125 (I22014,I21975);
nand I_1126 (I21663,I22014,I21853);
nor I_1127 (I22045,I471866,I471857);
not I_1128 (I22062,I22045);
nor I_1129 (I22079,I22014,I22062);
nor I_1130 (I22096,I21720,I22079);
DFFARX1 I_1131 (I22096,I2859,I21686,I21672,);
nor I_1132 (I22127,I21780,I22062);
nor I_1133 (I21660,I21975,I22127);
nor I_1134 (I21669,I21910,I22045);
nor I_1135 (I21657,I21780,I22045);
not I_1136 (I22213,I2866);
DFFARX1 I_1137 (I320183,I2859,I22213,I22239,);
not I_1138 (I22247,I22239);
nand I_1139 (I22264,I320180,I320195);
and I_1140 (I22281,I22264,I320177);
DFFARX1 I_1141 (I22281,I2859,I22213,I22307,);
DFFARX1 I_1142 (I320174,I2859,I22213,I22324,);
and I_1143 (I22332,I22324,I320174);
nor I_1144 (I22349,I22307,I22332);
DFFARX1 I_1145 (I22349,I2859,I22213,I22181,);
nand I_1146 (I22380,I22324,I320174);
nand I_1147 (I22397,I22247,I22380);
not I_1148 (I22193,I22397);
DFFARX1 I_1149 (I320177,I2859,I22213,I22437,);
DFFARX1 I_1150 (I22437,I2859,I22213,I22202,);
nand I_1151 (I22459,I320189,I320180);
and I_1152 (I22476,I22459,I320192);
DFFARX1 I_1153 (I22476,I2859,I22213,I22502,);
DFFARX1 I_1154 (I22502,I2859,I22213,I22519,);
not I_1155 (I22205,I22519);
not I_1156 (I22541,I22502);
nand I_1157 (I22190,I22541,I22380);
nor I_1158 (I22572,I320186,I320180);
not I_1159 (I22589,I22572);
nor I_1160 (I22606,I22541,I22589);
nor I_1161 (I22623,I22247,I22606);
DFFARX1 I_1162 (I22623,I2859,I22213,I22199,);
nor I_1163 (I22654,I22307,I22589);
nor I_1164 (I22187,I22502,I22654);
nor I_1165 (I22196,I22437,I22572);
nor I_1166 (I22184,I22307,I22572);
not I_1167 (I22740,I2866);
DFFARX1 I_1168 (I420392,I2859,I22740,I22766,);
not I_1169 (I22774,I22766);
nand I_1170 (I22791,I420389,I420395);
and I_1171 (I22808,I22791,I420392);
DFFARX1 I_1172 (I22808,I2859,I22740,I22834,);
DFFARX1 I_1173 (I420395,I2859,I22740,I22851,);
and I_1174 (I22859,I22851,I420389);
nor I_1175 (I22876,I22834,I22859);
DFFARX1 I_1176 (I22876,I2859,I22740,I22708,);
nand I_1177 (I22907,I22851,I420389);
nand I_1178 (I22924,I22774,I22907);
not I_1179 (I22720,I22924);
DFFARX1 I_1180 (I420398,I2859,I22740,I22964,);
DFFARX1 I_1181 (I22964,I2859,I22740,I22729,);
nand I_1182 (I22986,I420401,I420410);
and I_1183 (I23003,I22986,I420404);
DFFARX1 I_1184 (I23003,I2859,I22740,I23029,);
DFFARX1 I_1185 (I23029,I2859,I22740,I23046,);
not I_1186 (I22732,I23046);
not I_1187 (I23068,I23029);
nand I_1188 (I22717,I23068,I22907);
nor I_1189 (I23099,I420407,I420410);
not I_1190 (I23116,I23099);
nor I_1191 (I23133,I23068,I23116);
nor I_1192 (I23150,I22774,I23133);
DFFARX1 I_1193 (I23150,I2859,I22740,I22726,);
nor I_1194 (I23181,I22834,I23116);
nor I_1195 (I22714,I23029,I23181);
nor I_1196 (I22723,I22964,I23099);
nor I_1197 (I22711,I22834,I23099);
not I_1198 (I23267,I2866);
DFFARX1 I_1199 (I139882,I2859,I23267,I23293,);
not I_1200 (I23301,I23293);
nand I_1201 (I23318,I139864,I139879);
and I_1202 (I23335,I23318,I139855);
DFFARX1 I_1203 (I23335,I2859,I23267,I23361,);
DFFARX1 I_1204 (I139858,I2859,I23267,I23378,);
and I_1205 (I23386,I23378,I139873);
nor I_1206 (I23403,I23361,I23386);
DFFARX1 I_1207 (I23403,I2859,I23267,I23235,);
nand I_1208 (I23434,I23378,I139873);
nand I_1209 (I23451,I23301,I23434);
not I_1210 (I23247,I23451);
DFFARX1 I_1211 (I139876,I2859,I23267,I23491,);
DFFARX1 I_1212 (I23491,I2859,I23267,I23256,);
nand I_1213 (I23513,I139855,I139867);
and I_1214 (I23530,I23513,I139861);
DFFARX1 I_1215 (I23530,I2859,I23267,I23556,);
DFFARX1 I_1216 (I23556,I2859,I23267,I23573,);
not I_1217 (I23259,I23573);
not I_1218 (I23595,I23556);
nand I_1219 (I23244,I23595,I23434);
nor I_1220 (I23626,I139870,I139867);
not I_1221 (I23643,I23626);
nor I_1222 (I23660,I23595,I23643);
nor I_1223 (I23677,I23301,I23660);
DFFARX1 I_1224 (I23677,I2859,I23267,I23253,);
nor I_1225 (I23708,I23361,I23643);
nor I_1226 (I23241,I23556,I23708);
nor I_1227 (I23250,I23491,I23626);
nor I_1228 (I23238,I23361,I23626);
not I_1229 (I23794,I2866);
DFFARX1 I_1230 (I245825,I2859,I23794,I23820,);
not I_1231 (I23828,I23820);
nand I_1232 (I23845,I245837,I245822);
and I_1233 (I23862,I23845,I245816);
DFFARX1 I_1234 (I23862,I2859,I23794,I23888,);
DFFARX1 I_1235 (I245831,I2859,I23794,I23905,);
and I_1236 (I23913,I23905,I245819);
nor I_1237 (I23930,I23888,I23913);
DFFARX1 I_1238 (I23930,I2859,I23794,I23762,);
nand I_1239 (I23961,I23905,I245819);
nand I_1240 (I23978,I23828,I23961);
not I_1241 (I23774,I23978);
DFFARX1 I_1242 (I245828,I2859,I23794,I24018,);
DFFARX1 I_1243 (I24018,I2859,I23794,I23783,);
nand I_1244 (I24040,I245834,I245840);
and I_1245 (I24057,I24040,I245816);
DFFARX1 I_1246 (I24057,I2859,I23794,I24083,);
DFFARX1 I_1247 (I24083,I2859,I23794,I24100,);
not I_1248 (I23786,I24100);
not I_1249 (I24122,I24083);
nand I_1250 (I23771,I24122,I23961);
nor I_1251 (I24153,I245819,I245840);
not I_1252 (I24170,I24153);
nor I_1253 (I24187,I24122,I24170);
nor I_1254 (I24204,I23828,I24187);
DFFARX1 I_1255 (I24204,I2859,I23794,I23780,);
nor I_1256 (I24235,I23888,I24170);
nor I_1257 (I23768,I24083,I24235);
nor I_1258 (I23777,I24018,I24153);
nor I_1259 (I23765,I23888,I24153);
not I_1260 (I24321,I2866);
DFFARX1 I_1261 (I476478,I2859,I24321,I24347,);
not I_1262 (I24355,I24347);
nand I_1263 (I24372,I476493,I476472);
and I_1264 (I24389,I24372,I476475);
DFFARX1 I_1265 (I24389,I2859,I24321,I24415,);
DFFARX1 I_1266 (I476496,I2859,I24321,I24432,);
and I_1267 (I24440,I24432,I476475);
nor I_1268 (I24457,I24415,I24440);
DFFARX1 I_1269 (I24457,I2859,I24321,I24289,);
nand I_1270 (I24488,I24432,I476475);
nand I_1271 (I24505,I24355,I24488);
not I_1272 (I24301,I24505);
DFFARX1 I_1273 (I476472,I2859,I24321,I24545,);
DFFARX1 I_1274 (I24545,I2859,I24321,I24310,);
nand I_1275 (I24567,I476484,I476481);
and I_1276 (I24584,I24567,I476487);
DFFARX1 I_1277 (I24584,I2859,I24321,I24610,);
DFFARX1 I_1278 (I24610,I2859,I24321,I24627,);
not I_1279 (I24313,I24627);
not I_1280 (I24649,I24610);
nand I_1281 (I24298,I24649,I24488);
nor I_1282 (I24680,I476490,I476481);
not I_1283 (I24697,I24680);
nor I_1284 (I24714,I24649,I24697);
nor I_1285 (I24731,I24355,I24714);
DFFARX1 I_1286 (I24731,I2859,I24321,I24307,);
nor I_1287 (I24762,I24415,I24697);
nor I_1288 (I24295,I24610,I24762);
nor I_1289 (I24304,I24545,I24680);
nor I_1290 (I24292,I24415,I24680);
not I_1291 (I24848,I2866);
DFFARX1 I_1292 (I460294,I2859,I24848,I24874,);
not I_1293 (I24882,I24874);
nand I_1294 (I24899,I460309,I460288);
and I_1295 (I24916,I24899,I460291);
DFFARX1 I_1296 (I24916,I2859,I24848,I24942,);
DFFARX1 I_1297 (I460312,I2859,I24848,I24959,);
and I_1298 (I24967,I24959,I460291);
nor I_1299 (I24984,I24942,I24967);
DFFARX1 I_1300 (I24984,I2859,I24848,I24816,);
nand I_1301 (I25015,I24959,I460291);
nand I_1302 (I25032,I24882,I25015);
not I_1303 (I24828,I25032);
DFFARX1 I_1304 (I460288,I2859,I24848,I25072,);
DFFARX1 I_1305 (I25072,I2859,I24848,I24837,);
nand I_1306 (I25094,I460300,I460297);
and I_1307 (I25111,I25094,I460303);
DFFARX1 I_1308 (I25111,I2859,I24848,I25137,);
DFFARX1 I_1309 (I25137,I2859,I24848,I25154,);
not I_1310 (I24840,I25154);
not I_1311 (I25176,I25137);
nand I_1312 (I24825,I25176,I25015);
nor I_1313 (I25207,I460306,I460297);
not I_1314 (I25224,I25207);
nor I_1315 (I25241,I25176,I25224);
nor I_1316 (I25258,I24882,I25241);
DFFARX1 I_1317 (I25258,I2859,I24848,I24834,);
nor I_1318 (I25289,I24942,I25224);
nor I_1319 (I24822,I25137,I25289);
nor I_1320 (I24831,I25072,I25207);
nor I_1321 (I24819,I24942,I25207);
not I_1322 (I25375,I2866);
DFFARX1 I_1323 (I333358,I2859,I25375,I25401,);
not I_1324 (I25409,I25401);
nand I_1325 (I25426,I333355,I333370);
and I_1326 (I25443,I25426,I333352);
DFFARX1 I_1327 (I25443,I2859,I25375,I25469,);
DFFARX1 I_1328 (I333349,I2859,I25375,I25486,);
and I_1329 (I25494,I25486,I333349);
nor I_1330 (I25511,I25469,I25494);
DFFARX1 I_1331 (I25511,I2859,I25375,I25343,);
nand I_1332 (I25542,I25486,I333349);
nand I_1333 (I25559,I25409,I25542);
not I_1334 (I25355,I25559);
DFFARX1 I_1335 (I333352,I2859,I25375,I25599,);
DFFARX1 I_1336 (I25599,I2859,I25375,I25364,);
nand I_1337 (I25621,I333364,I333355);
and I_1338 (I25638,I25621,I333367);
DFFARX1 I_1339 (I25638,I2859,I25375,I25664,);
DFFARX1 I_1340 (I25664,I2859,I25375,I25681,);
not I_1341 (I25367,I25681);
not I_1342 (I25703,I25664);
nand I_1343 (I25352,I25703,I25542);
nor I_1344 (I25734,I333361,I333355);
not I_1345 (I25751,I25734);
nor I_1346 (I25768,I25703,I25751);
nor I_1347 (I25785,I25409,I25768);
DFFARX1 I_1348 (I25785,I2859,I25375,I25361,);
nor I_1349 (I25816,I25469,I25751);
nor I_1350 (I25349,I25664,I25816);
nor I_1351 (I25358,I25599,I25734);
nor I_1352 (I25346,I25469,I25734);
not I_1353 (I25902,I2866);
DFFARX1 I_1354 (I374736,I2859,I25902,I25928,);
not I_1355 (I25936,I25928);
nand I_1356 (I25953,I374754,I374748);
and I_1357 (I25970,I25953,I374727);
DFFARX1 I_1358 (I25970,I2859,I25902,I25996,);
DFFARX1 I_1359 (I374745,I2859,I25902,I26013,);
and I_1360 (I26021,I26013,I374730);
nor I_1361 (I26038,I25996,I26021);
DFFARX1 I_1362 (I26038,I2859,I25902,I25870,);
nand I_1363 (I26069,I26013,I374730);
nand I_1364 (I26086,I25936,I26069);
not I_1365 (I25882,I26086);
DFFARX1 I_1366 (I374742,I2859,I25902,I26126,);
DFFARX1 I_1367 (I26126,I2859,I25902,I25891,);
nand I_1368 (I26148,I374751,I374739);
and I_1369 (I26165,I26148,I374733);
DFFARX1 I_1370 (I26165,I2859,I25902,I26191,);
DFFARX1 I_1371 (I26191,I2859,I25902,I26208,);
not I_1372 (I25894,I26208);
not I_1373 (I26230,I26191);
nand I_1374 (I25879,I26230,I26069);
nor I_1375 (I26261,I374727,I374739);
not I_1376 (I26278,I26261);
nor I_1377 (I26295,I26230,I26278);
nor I_1378 (I26312,I25936,I26295);
DFFARX1 I_1379 (I26312,I2859,I25902,I25888,);
nor I_1380 (I26343,I25996,I26278);
nor I_1381 (I25876,I26191,I26343);
nor I_1382 (I25885,I26126,I26261);
nor I_1383 (I25873,I25996,I26261);
not I_1384 (I26429,I2866);
DFFARX1 I_1385 (I391532,I2859,I26429,I26455,);
not I_1386 (I26463,I26455);
nand I_1387 (I26480,I391550,I391544);
and I_1388 (I26497,I26480,I391523);
DFFARX1 I_1389 (I26497,I2859,I26429,I26523,);
DFFARX1 I_1390 (I391541,I2859,I26429,I26540,);
and I_1391 (I26548,I26540,I391526);
nor I_1392 (I26565,I26523,I26548);
DFFARX1 I_1393 (I26565,I2859,I26429,I26397,);
nand I_1394 (I26596,I26540,I391526);
nand I_1395 (I26613,I26463,I26596);
not I_1396 (I26409,I26613);
DFFARX1 I_1397 (I391538,I2859,I26429,I26653,);
DFFARX1 I_1398 (I26653,I2859,I26429,I26418,);
nand I_1399 (I26675,I391547,I391535);
and I_1400 (I26692,I26675,I391529);
DFFARX1 I_1401 (I26692,I2859,I26429,I26718,);
DFFARX1 I_1402 (I26718,I2859,I26429,I26735,);
not I_1403 (I26421,I26735);
not I_1404 (I26757,I26718);
nand I_1405 (I26406,I26757,I26596);
nor I_1406 (I26788,I391523,I391535);
not I_1407 (I26805,I26788);
nor I_1408 (I26822,I26757,I26805);
nor I_1409 (I26839,I26463,I26822);
DFFARX1 I_1410 (I26839,I2859,I26429,I26415,);
nor I_1411 (I26870,I26523,I26805);
nor I_1412 (I26403,I26718,I26870);
nor I_1413 (I26412,I26653,I26788);
nor I_1414 (I26400,I26523,I26788);
not I_1415 (I26956,I2866);
DFFARX1 I_1416 (I505208,I2859,I26956,I26982,);
not I_1417 (I26990,I26982);
nand I_1418 (I27007,I505202,I505223);
and I_1419 (I27024,I27007,I505214);
DFFARX1 I_1420 (I27024,I2859,I26956,I27050,);
DFFARX1 I_1421 (I505205,I2859,I26956,I27067,);
and I_1422 (I27075,I27067,I505217);
nor I_1423 (I27092,I27050,I27075);
DFFARX1 I_1424 (I27092,I2859,I26956,I26924,);
nand I_1425 (I27123,I27067,I505217);
nand I_1426 (I27140,I26990,I27123);
not I_1427 (I26936,I27140);
DFFARX1 I_1428 (I505205,I2859,I26956,I27180,);
DFFARX1 I_1429 (I27180,I2859,I26956,I26945,);
nand I_1430 (I27202,I505226,I505211);
and I_1431 (I27219,I27202,I505202);
DFFARX1 I_1432 (I27219,I2859,I26956,I27245,);
DFFARX1 I_1433 (I27245,I2859,I26956,I27262,);
not I_1434 (I26948,I27262);
not I_1435 (I27284,I27245);
nand I_1436 (I26933,I27284,I27123);
nor I_1437 (I27315,I505220,I505211);
not I_1438 (I27332,I27315);
nor I_1439 (I27349,I27284,I27332);
nor I_1440 (I27366,I26990,I27349);
DFFARX1 I_1441 (I27366,I2859,I26956,I26942,);
nor I_1442 (I27397,I27050,I27332);
nor I_1443 (I26930,I27245,I27397);
nor I_1444 (I26939,I27180,I27315);
nor I_1445 (I26927,I27050,I27315);
not I_1446 (I27483,I2866);
DFFARX1 I_1447 (I120910,I2859,I27483,I27509,);
not I_1448 (I27517,I27509);
nand I_1449 (I27534,I120892,I120907);
and I_1450 (I27551,I27534,I120883);
DFFARX1 I_1451 (I27551,I2859,I27483,I27577,);
DFFARX1 I_1452 (I120886,I2859,I27483,I27594,);
and I_1453 (I27602,I27594,I120901);
nor I_1454 (I27619,I27577,I27602);
DFFARX1 I_1455 (I27619,I2859,I27483,I27451,);
nand I_1456 (I27650,I27594,I120901);
nand I_1457 (I27667,I27517,I27650);
not I_1458 (I27463,I27667);
DFFARX1 I_1459 (I120904,I2859,I27483,I27707,);
DFFARX1 I_1460 (I27707,I2859,I27483,I27472,);
nand I_1461 (I27729,I120883,I120895);
and I_1462 (I27746,I27729,I120889);
DFFARX1 I_1463 (I27746,I2859,I27483,I27772,);
DFFARX1 I_1464 (I27772,I2859,I27483,I27789,);
not I_1465 (I27475,I27789);
not I_1466 (I27811,I27772);
nand I_1467 (I27460,I27811,I27650);
nor I_1468 (I27842,I120898,I120895);
not I_1469 (I27859,I27842);
nor I_1470 (I27876,I27811,I27859);
nor I_1471 (I27893,I27517,I27876);
DFFARX1 I_1472 (I27893,I2859,I27483,I27469,);
nor I_1473 (I27924,I27577,I27859);
nor I_1474 (I27457,I27772,I27924);
nor I_1475 (I27466,I27707,I27842);
nor I_1476 (I27454,I27577,I27842);
not I_1477 (I28010,I2866);
DFFARX1 I_1478 (I403160,I2859,I28010,I28036,);
not I_1479 (I28044,I28036);
nand I_1480 (I28061,I403178,I403172);
and I_1481 (I28078,I28061,I403151);
DFFARX1 I_1482 (I28078,I2859,I28010,I28104,);
DFFARX1 I_1483 (I403169,I2859,I28010,I28121,);
and I_1484 (I28129,I28121,I403154);
nor I_1485 (I28146,I28104,I28129);
DFFARX1 I_1486 (I28146,I2859,I28010,I27978,);
nand I_1487 (I28177,I28121,I403154);
nand I_1488 (I28194,I28044,I28177);
not I_1489 (I27990,I28194);
DFFARX1 I_1490 (I403166,I2859,I28010,I28234,);
DFFARX1 I_1491 (I28234,I2859,I28010,I27999,);
nand I_1492 (I28256,I403175,I403163);
and I_1493 (I28273,I28256,I403157);
DFFARX1 I_1494 (I28273,I2859,I28010,I28299,);
DFFARX1 I_1495 (I28299,I2859,I28010,I28316,);
not I_1496 (I28002,I28316);
not I_1497 (I28338,I28299);
nand I_1498 (I27987,I28338,I28177);
nor I_1499 (I28369,I403151,I403163);
not I_1500 (I28386,I28369);
nor I_1501 (I28403,I28338,I28386);
nor I_1502 (I28420,I28044,I28403);
DFFARX1 I_1503 (I28420,I2859,I28010,I27996,);
nor I_1504 (I28451,I28104,I28386);
nor I_1505 (I27984,I28299,I28451);
nor I_1506 (I27993,I28234,I28369);
nor I_1507 (I27981,I28104,I28369);
not I_1508 (I28537,I2866);
DFFARX1 I_1509 (I255651,I2859,I28537,I28563,);
not I_1510 (I28571,I28563);
nand I_1511 (I28588,I255663,I255648);
and I_1512 (I28605,I28588,I255642);
DFFARX1 I_1513 (I28605,I2859,I28537,I28631,);
DFFARX1 I_1514 (I255657,I2859,I28537,I28648,);
and I_1515 (I28656,I28648,I255645);
nor I_1516 (I28673,I28631,I28656);
DFFARX1 I_1517 (I28673,I2859,I28537,I28505,);
nand I_1518 (I28704,I28648,I255645);
nand I_1519 (I28721,I28571,I28704);
not I_1520 (I28517,I28721);
DFFARX1 I_1521 (I255654,I2859,I28537,I28761,);
DFFARX1 I_1522 (I28761,I2859,I28537,I28526,);
nand I_1523 (I28783,I255660,I255666);
and I_1524 (I28800,I28783,I255642);
DFFARX1 I_1525 (I28800,I2859,I28537,I28826,);
DFFARX1 I_1526 (I28826,I2859,I28537,I28843,);
not I_1527 (I28529,I28843);
not I_1528 (I28865,I28826);
nand I_1529 (I28514,I28865,I28704);
nor I_1530 (I28896,I255645,I255666);
not I_1531 (I28913,I28896);
nor I_1532 (I28930,I28865,I28913);
nor I_1533 (I28947,I28571,I28930);
DFFARX1 I_1534 (I28947,I2859,I28537,I28523,);
nor I_1535 (I28978,I28631,I28913);
nor I_1536 (I28511,I28826,I28978);
nor I_1537 (I28520,I28761,I28896);
nor I_1538 (I28508,I28631,I28896);
not I_1539 (I29064,I2866);
DFFARX1 I_1540 (I171306,I2859,I29064,I29090,);
not I_1541 (I29098,I29090);
nand I_1542 (I29115,I171300,I171291);
and I_1543 (I29132,I29115,I171312);
DFFARX1 I_1544 (I29132,I2859,I29064,I29158,);
DFFARX1 I_1545 (I171294,I2859,I29064,I29175,);
and I_1546 (I29183,I29175,I171288);
nor I_1547 (I29200,I29158,I29183);
DFFARX1 I_1548 (I29200,I2859,I29064,I29032,);
nand I_1549 (I29231,I29175,I171288);
nand I_1550 (I29248,I29098,I29231);
not I_1551 (I29044,I29248);
DFFARX1 I_1552 (I171288,I2859,I29064,I29288,);
DFFARX1 I_1553 (I29288,I2859,I29064,I29053,);
nand I_1554 (I29310,I171315,I171297);
and I_1555 (I29327,I29310,I171303);
DFFARX1 I_1556 (I29327,I2859,I29064,I29353,);
DFFARX1 I_1557 (I29353,I2859,I29064,I29370,);
not I_1558 (I29056,I29370);
not I_1559 (I29392,I29353);
nand I_1560 (I29041,I29392,I29231);
nor I_1561 (I29423,I171309,I171297);
not I_1562 (I29440,I29423);
nor I_1563 (I29457,I29392,I29440);
nor I_1564 (I29474,I29098,I29457);
DFFARX1 I_1565 (I29474,I2859,I29064,I29050,);
nor I_1566 (I29505,I29158,I29440);
nor I_1567 (I29038,I29353,I29505);
nor I_1568 (I29047,I29288,I29423);
nor I_1569 (I29035,I29158,I29423);
not I_1570 (I29591,I2866);
DFFARX1 I_1571 (I59644,I2859,I29591,I29617,);
not I_1572 (I29625,I29617);
nand I_1573 (I29642,I59638,I59632);
and I_1574 (I29659,I29642,I59653);
DFFARX1 I_1575 (I29659,I2859,I29591,I29685,);
DFFARX1 I_1576 (I59650,I2859,I29591,I29702,);
and I_1577 (I29710,I29702,I59647);
nor I_1578 (I29727,I29685,I29710);
DFFARX1 I_1579 (I29727,I2859,I29591,I29559,);
nand I_1580 (I29758,I29702,I59647);
nand I_1581 (I29775,I29625,I29758);
not I_1582 (I29571,I29775);
DFFARX1 I_1583 (I59632,I2859,I29591,I29815,);
DFFARX1 I_1584 (I29815,I2859,I29591,I29580,);
nand I_1585 (I29837,I59635,I59635);
and I_1586 (I29854,I29837,I59656);
DFFARX1 I_1587 (I29854,I2859,I29591,I29880,);
DFFARX1 I_1588 (I29880,I2859,I29591,I29897,);
not I_1589 (I29583,I29897);
not I_1590 (I29919,I29880);
nand I_1591 (I29568,I29919,I29758);
nor I_1592 (I29950,I59641,I59635);
not I_1593 (I29967,I29950);
nor I_1594 (I29984,I29919,I29967);
nor I_1595 (I30001,I29625,I29984);
DFFARX1 I_1596 (I30001,I2859,I29591,I29577,);
nor I_1597 (I30032,I29685,I29967);
nor I_1598 (I29565,I29880,I30032);
nor I_1599 (I29574,I29815,I29950);
nor I_1600 (I29562,I29685,I29950);
not I_1601 (I30118,I2866);
DFFARX1 I_1602 (I94154,I2859,I30118,I30144,);
not I_1603 (I30152,I30144);
nand I_1604 (I30169,I94148,I94142);
and I_1605 (I30186,I30169,I94163);
DFFARX1 I_1606 (I30186,I2859,I30118,I30212,);
DFFARX1 I_1607 (I94160,I2859,I30118,I30229,);
and I_1608 (I30237,I30229,I94157);
nor I_1609 (I30254,I30212,I30237);
DFFARX1 I_1610 (I30254,I2859,I30118,I30086,);
nand I_1611 (I30285,I30229,I94157);
nand I_1612 (I30302,I30152,I30285);
not I_1613 (I30098,I30302);
DFFARX1 I_1614 (I94142,I2859,I30118,I30342,);
DFFARX1 I_1615 (I30342,I2859,I30118,I30107,);
nand I_1616 (I30364,I94145,I94145);
and I_1617 (I30381,I30364,I94166);
DFFARX1 I_1618 (I30381,I2859,I30118,I30407,);
DFFARX1 I_1619 (I30407,I2859,I30118,I30424,);
not I_1620 (I30110,I30424);
not I_1621 (I30446,I30407);
nand I_1622 (I30095,I30446,I30285);
nor I_1623 (I30477,I94151,I94145);
not I_1624 (I30494,I30477);
nor I_1625 (I30511,I30446,I30494);
nor I_1626 (I30528,I30152,I30511);
DFFARX1 I_1627 (I30528,I2859,I30118,I30104,);
nor I_1628 (I30559,I30212,I30494);
nor I_1629 (I30092,I30407,I30559);
nor I_1630 (I30101,I30342,I30477);
nor I_1631 (I30089,I30212,I30477);
not I_1632 (I30645,I2866);
DFFARX1 I_1633 (I67974,I2859,I30645,I30671,);
not I_1634 (I30679,I30671);
nand I_1635 (I30696,I67968,I67962);
and I_1636 (I30713,I30696,I67983);
DFFARX1 I_1637 (I30713,I2859,I30645,I30739,);
DFFARX1 I_1638 (I67980,I2859,I30645,I30756,);
and I_1639 (I30764,I30756,I67977);
nor I_1640 (I30781,I30739,I30764);
DFFARX1 I_1641 (I30781,I2859,I30645,I30613,);
nand I_1642 (I30812,I30756,I67977);
nand I_1643 (I30829,I30679,I30812);
not I_1644 (I30625,I30829);
DFFARX1 I_1645 (I67962,I2859,I30645,I30869,);
DFFARX1 I_1646 (I30869,I2859,I30645,I30634,);
nand I_1647 (I30891,I67965,I67965);
and I_1648 (I30908,I30891,I67986);
DFFARX1 I_1649 (I30908,I2859,I30645,I30934,);
DFFARX1 I_1650 (I30934,I2859,I30645,I30951,);
not I_1651 (I30637,I30951);
not I_1652 (I30973,I30934);
nand I_1653 (I30622,I30973,I30812);
nor I_1654 (I31004,I67971,I67965);
not I_1655 (I31021,I31004);
nor I_1656 (I31038,I30973,I31021);
nor I_1657 (I31055,I30679,I31038);
DFFARX1 I_1658 (I31055,I2859,I30645,I30631,);
nor I_1659 (I31086,I30739,I31021);
nor I_1660 (I30619,I30934,I31086);
nor I_1661 (I30628,I30869,I31004);
nor I_1662 (I30616,I30739,I31004);
not I_1663 (I31172,I2866);
DFFARX1 I_1664 (I145679,I2859,I31172,I31198,);
not I_1665 (I31206,I31198);
nand I_1666 (I31223,I145661,I145676);
and I_1667 (I31240,I31223,I145652);
DFFARX1 I_1668 (I31240,I2859,I31172,I31266,);
DFFARX1 I_1669 (I145655,I2859,I31172,I31283,);
and I_1670 (I31291,I31283,I145670);
nor I_1671 (I31308,I31266,I31291);
DFFARX1 I_1672 (I31308,I2859,I31172,I31140,);
nand I_1673 (I31339,I31283,I145670);
nand I_1674 (I31356,I31206,I31339);
not I_1675 (I31152,I31356);
DFFARX1 I_1676 (I145673,I2859,I31172,I31396,);
DFFARX1 I_1677 (I31396,I2859,I31172,I31161,);
nand I_1678 (I31418,I145652,I145664);
and I_1679 (I31435,I31418,I145658);
DFFARX1 I_1680 (I31435,I2859,I31172,I31461,);
DFFARX1 I_1681 (I31461,I2859,I31172,I31478,);
not I_1682 (I31164,I31478);
not I_1683 (I31500,I31461);
nand I_1684 (I31149,I31500,I31339);
nor I_1685 (I31531,I145667,I145664);
not I_1686 (I31548,I31531);
nor I_1687 (I31565,I31500,I31548);
nor I_1688 (I31582,I31206,I31565);
DFFARX1 I_1689 (I31582,I2859,I31172,I31158,);
nor I_1690 (I31613,I31266,I31548);
nor I_1691 (I31146,I31461,I31613);
nor I_1692 (I31155,I31396,I31531);
nor I_1693 (I31143,I31266,I31531);
not I_1694 (I31699,I2866);
DFFARX1 I_1695 (I335466,I2859,I31699,I31725,);
not I_1696 (I31733,I31725);
nand I_1697 (I31750,I335463,I335478);
and I_1698 (I31767,I31750,I335460);
DFFARX1 I_1699 (I31767,I2859,I31699,I31793,);
DFFARX1 I_1700 (I335457,I2859,I31699,I31810,);
and I_1701 (I31818,I31810,I335457);
nor I_1702 (I31835,I31793,I31818);
DFFARX1 I_1703 (I31835,I2859,I31699,I31667,);
nand I_1704 (I31866,I31810,I335457);
nand I_1705 (I31883,I31733,I31866);
not I_1706 (I31679,I31883);
DFFARX1 I_1707 (I335460,I2859,I31699,I31923,);
DFFARX1 I_1708 (I31923,I2859,I31699,I31688,);
nand I_1709 (I31945,I335472,I335463);
and I_1710 (I31962,I31945,I335475);
DFFARX1 I_1711 (I31962,I2859,I31699,I31988,);
DFFARX1 I_1712 (I31988,I2859,I31699,I32005,);
not I_1713 (I31691,I32005);
not I_1714 (I32027,I31988);
nand I_1715 (I31676,I32027,I31866);
nor I_1716 (I32058,I335469,I335463);
not I_1717 (I32075,I32058);
nor I_1718 (I32092,I32027,I32075);
nor I_1719 (I32109,I31733,I32092);
DFFARX1 I_1720 (I32109,I2859,I31699,I31685,);
nor I_1721 (I32140,I31793,I32075);
nor I_1722 (I31673,I31988,I32140);
nor I_1723 (I31682,I31923,I32058);
nor I_1724 (I31670,I31793,I32058);
not I_1725 (I32226,I2866);
DFFARX1 I_1726 (I166410,I2859,I32226,I32252,);
not I_1727 (I32260,I32252);
nand I_1728 (I32277,I166404,I166395);
and I_1729 (I32294,I32277,I166416);
DFFARX1 I_1730 (I32294,I2859,I32226,I32320,);
DFFARX1 I_1731 (I166398,I2859,I32226,I32337,);
and I_1732 (I32345,I32337,I166392);
nor I_1733 (I32362,I32320,I32345);
DFFARX1 I_1734 (I32362,I2859,I32226,I32194,);
nand I_1735 (I32393,I32337,I166392);
nand I_1736 (I32410,I32260,I32393);
not I_1737 (I32206,I32410);
DFFARX1 I_1738 (I166392,I2859,I32226,I32450,);
DFFARX1 I_1739 (I32450,I2859,I32226,I32215,);
nand I_1740 (I32472,I166419,I166401);
and I_1741 (I32489,I32472,I166407);
DFFARX1 I_1742 (I32489,I2859,I32226,I32515,);
DFFARX1 I_1743 (I32515,I2859,I32226,I32532,);
not I_1744 (I32218,I32532);
not I_1745 (I32554,I32515);
nand I_1746 (I32203,I32554,I32393);
nor I_1747 (I32585,I166413,I166401);
not I_1748 (I32602,I32585);
nor I_1749 (I32619,I32554,I32602);
nor I_1750 (I32636,I32260,I32619);
DFFARX1 I_1751 (I32636,I2859,I32226,I32212,);
nor I_1752 (I32667,I32320,I32602);
nor I_1753 (I32200,I32515,I32667);
nor I_1754 (I32209,I32450,I32585);
nor I_1755 (I32197,I32320,I32585);
not I_1756 (I32753,I2866);
DFFARX1 I_1757 (I563592,I2859,I32753,I32779,);
not I_1758 (I32787,I32779);
nand I_1759 (I32804,I563586,I563607);
and I_1760 (I32821,I32804,I563583);
DFFARX1 I_1761 (I32821,I2859,I32753,I32847,);
DFFARX1 I_1762 (I563604,I2859,I32753,I32864,);
and I_1763 (I32872,I32864,I563601);
nor I_1764 (I32889,I32847,I32872);
DFFARX1 I_1765 (I32889,I2859,I32753,I32721,);
nand I_1766 (I32920,I32864,I563601);
nand I_1767 (I32937,I32787,I32920);
not I_1768 (I32733,I32937);
DFFARX1 I_1769 (I563589,I2859,I32753,I32977,);
DFFARX1 I_1770 (I32977,I2859,I32753,I32742,);
nand I_1771 (I32999,I563598,I563595);
and I_1772 (I33016,I32999,I563580);
DFFARX1 I_1773 (I33016,I2859,I32753,I33042,);
DFFARX1 I_1774 (I33042,I2859,I32753,I33059,);
not I_1775 (I32745,I33059);
not I_1776 (I33081,I33042);
nand I_1777 (I32730,I33081,I32920);
nor I_1778 (I33112,I563580,I563595);
not I_1779 (I33129,I33112);
nor I_1780 (I33146,I33081,I33129);
nor I_1781 (I33163,I32787,I33146);
DFFARX1 I_1782 (I33163,I2859,I32753,I32739,);
nor I_1783 (I33194,I32847,I33129);
nor I_1784 (I32727,I33042,I33194);
nor I_1785 (I32736,I32977,I33112);
nor I_1786 (I32724,I32847,I33112);
not I_1787 (I33280,I2866);
DFFARX1 I_1788 (I445266,I2859,I33280,I33306,);
not I_1789 (I33314,I33306);
nand I_1790 (I33331,I445281,I445260);
and I_1791 (I33348,I33331,I445263);
DFFARX1 I_1792 (I33348,I2859,I33280,I33374,);
DFFARX1 I_1793 (I445284,I2859,I33280,I33391,);
and I_1794 (I33399,I33391,I445263);
nor I_1795 (I33416,I33374,I33399);
DFFARX1 I_1796 (I33416,I2859,I33280,I33248,);
nand I_1797 (I33447,I33391,I445263);
nand I_1798 (I33464,I33314,I33447);
not I_1799 (I33260,I33464);
DFFARX1 I_1800 (I445260,I2859,I33280,I33504,);
DFFARX1 I_1801 (I33504,I2859,I33280,I33269,);
nand I_1802 (I33526,I445272,I445269);
and I_1803 (I33543,I33526,I445275);
DFFARX1 I_1804 (I33543,I2859,I33280,I33569,);
DFFARX1 I_1805 (I33569,I2859,I33280,I33586,);
not I_1806 (I33272,I33586);
not I_1807 (I33608,I33569);
nand I_1808 (I33257,I33608,I33447);
nor I_1809 (I33639,I445278,I445269);
not I_1810 (I33656,I33639);
nor I_1811 (I33673,I33608,I33656);
nor I_1812 (I33690,I33314,I33673);
DFFARX1 I_1813 (I33690,I2859,I33280,I33266,);
nor I_1814 (I33721,I33374,I33656);
nor I_1815 (I33254,I33569,I33721);
nor I_1816 (I33263,I33504,I33639);
nor I_1817 (I33251,I33374,I33639);
not I_1818 (I33807,I2866);
DFFARX1 I_1819 (I564187,I2859,I33807,I33833,);
not I_1820 (I33841,I33833);
nand I_1821 (I33858,I564181,I564202);
and I_1822 (I33875,I33858,I564178);
DFFARX1 I_1823 (I33875,I2859,I33807,I33901,);
DFFARX1 I_1824 (I564199,I2859,I33807,I33918,);
and I_1825 (I33926,I33918,I564196);
nor I_1826 (I33943,I33901,I33926);
DFFARX1 I_1827 (I33943,I2859,I33807,I33775,);
nand I_1828 (I33974,I33918,I564196);
nand I_1829 (I33991,I33841,I33974);
not I_1830 (I33787,I33991);
DFFARX1 I_1831 (I564184,I2859,I33807,I34031,);
DFFARX1 I_1832 (I34031,I2859,I33807,I33796,);
nand I_1833 (I34053,I564193,I564190);
and I_1834 (I34070,I34053,I564175);
DFFARX1 I_1835 (I34070,I2859,I33807,I34096,);
DFFARX1 I_1836 (I34096,I2859,I33807,I34113,);
not I_1837 (I33799,I34113);
not I_1838 (I34135,I34096);
nand I_1839 (I33784,I34135,I33974);
nor I_1840 (I34166,I564175,I564190);
not I_1841 (I34183,I34166);
nor I_1842 (I34200,I34135,I34183);
nor I_1843 (I34217,I33841,I34200);
DFFARX1 I_1844 (I34217,I2859,I33807,I33793,);
nor I_1845 (I34248,I33901,I34183);
nor I_1846 (I33781,I34096,I34248);
nor I_1847 (I33790,I34031,I34166);
nor I_1848 (I33778,I33901,I34166);
not I_1849 (I34334,I2866);
DFFARX1 I_1850 (I306518,I2859,I34334,I34360,);
not I_1851 (I34368,I34360);
nand I_1852 (I34385,I306509,I306527);
and I_1853 (I34402,I34385,I306506);
DFFARX1 I_1854 (I34402,I2859,I34334,I34428,);
DFFARX1 I_1855 (I306509,I2859,I34334,I34445,);
and I_1856 (I34453,I34445,I306512);
nor I_1857 (I34470,I34428,I34453);
DFFARX1 I_1858 (I34470,I2859,I34334,I34302,);
nand I_1859 (I34501,I34445,I306512);
nand I_1860 (I34518,I34368,I34501);
not I_1861 (I34314,I34518);
DFFARX1 I_1862 (I306506,I2859,I34334,I34558,);
DFFARX1 I_1863 (I34558,I2859,I34334,I34323,);
nand I_1864 (I34580,I306524,I306515);
and I_1865 (I34597,I34580,I306530);
DFFARX1 I_1866 (I34597,I2859,I34334,I34623,);
DFFARX1 I_1867 (I34623,I2859,I34334,I34640,);
not I_1868 (I34326,I34640);
not I_1869 (I34662,I34623);
nand I_1870 (I34311,I34662,I34501);
nor I_1871 (I34693,I306521,I306515);
not I_1872 (I34710,I34693);
nor I_1873 (I34727,I34662,I34710);
nor I_1874 (I34744,I34368,I34727);
DFFARX1 I_1875 (I34744,I2859,I34334,I34320,);
nor I_1876 (I34775,I34428,I34710);
nor I_1877 (I34308,I34623,I34775);
nor I_1878 (I34317,I34558,I34693);
nor I_1879 (I34305,I34428,I34693);
not I_1880 (I34861,I2866);
DFFARX1 I_1881 (I535032,I2859,I34861,I34887,);
not I_1882 (I34895,I34887);
nand I_1883 (I34912,I535026,I535047);
and I_1884 (I34929,I34912,I535023);
DFFARX1 I_1885 (I34929,I2859,I34861,I34955,);
DFFARX1 I_1886 (I535044,I2859,I34861,I34972,);
and I_1887 (I34980,I34972,I535041);
nor I_1888 (I34997,I34955,I34980);
DFFARX1 I_1889 (I34997,I2859,I34861,I34829,);
nand I_1890 (I35028,I34972,I535041);
nand I_1891 (I35045,I34895,I35028);
not I_1892 (I34841,I35045);
DFFARX1 I_1893 (I535029,I2859,I34861,I35085,);
DFFARX1 I_1894 (I35085,I2859,I34861,I34850,);
nand I_1895 (I35107,I535038,I535035);
and I_1896 (I35124,I35107,I535020);
DFFARX1 I_1897 (I35124,I2859,I34861,I35150,);
DFFARX1 I_1898 (I35150,I2859,I34861,I35167,);
not I_1899 (I34853,I35167);
not I_1900 (I35189,I35150);
nand I_1901 (I34838,I35189,I35028);
nor I_1902 (I35220,I535020,I535035);
not I_1903 (I35237,I35220);
nor I_1904 (I35254,I35189,I35237);
nor I_1905 (I35271,I34895,I35254);
DFFARX1 I_1906 (I35271,I2859,I34861,I34847,);
nor I_1907 (I35302,I34955,I35237);
nor I_1908 (I34835,I35150,I35302);
nor I_1909 (I34844,I35085,I35220);
nor I_1910 (I34832,I34955,I35220);
not I_1911 (I35388,I2866);
DFFARX1 I_1912 (I451046,I2859,I35388,I35414,);
not I_1913 (I35422,I35414);
nand I_1914 (I35439,I451061,I451040);
and I_1915 (I35456,I35439,I451043);
DFFARX1 I_1916 (I35456,I2859,I35388,I35482,);
DFFARX1 I_1917 (I451064,I2859,I35388,I35499,);
and I_1918 (I35507,I35499,I451043);
nor I_1919 (I35524,I35482,I35507);
DFFARX1 I_1920 (I35524,I2859,I35388,I35356,);
nand I_1921 (I35555,I35499,I451043);
nand I_1922 (I35572,I35422,I35555);
not I_1923 (I35368,I35572);
DFFARX1 I_1924 (I451040,I2859,I35388,I35612,);
DFFARX1 I_1925 (I35612,I2859,I35388,I35377,);
nand I_1926 (I35634,I451052,I451049);
and I_1927 (I35651,I35634,I451055);
DFFARX1 I_1928 (I35651,I2859,I35388,I35677,);
DFFARX1 I_1929 (I35677,I2859,I35388,I35694,);
not I_1930 (I35380,I35694);
not I_1931 (I35716,I35677);
nand I_1932 (I35365,I35716,I35555);
nor I_1933 (I35747,I451058,I451049);
not I_1934 (I35764,I35747);
nor I_1935 (I35781,I35716,I35764);
nor I_1936 (I35798,I35422,I35781);
DFFARX1 I_1937 (I35798,I2859,I35388,I35374,);
nor I_1938 (I35829,I35482,I35764);
nor I_1939 (I35362,I35677,I35829);
nor I_1940 (I35371,I35612,I35747);
nor I_1941 (I35359,I35482,I35747);
not I_1942 (I35915,I2866);
DFFARX1 I_1943 (I109029,I2859,I35915,I35941,);
not I_1944 (I35949,I35941);
nand I_1945 (I35966,I109023,I109017);
and I_1946 (I35983,I35966,I109038);
DFFARX1 I_1947 (I35983,I2859,I35915,I36009,);
DFFARX1 I_1948 (I109035,I2859,I35915,I36026,);
and I_1949 (I36034,I36026,I109032);
nor I_1950 (I36051,I36009,I36034);
DFFARX1 I_1951 (I36051,I2859,I35915,I35883,);
nand I_1952 (I36082,I36026,I109032);
nand I_1953 (I36099,I35949,I36082);
not I_1954 (I35895,I36099);
DFFARX1 I_1955 (I109017,I2859,I35915,I36139,);
DFFARX1 I_1956 (I36139,I2859,I35915,I35904,);
nand I_1957 (I36161,I109020,I109020);
and I_1958 (I36178,I36161,I109041);
DFFARX1 I_1959 (I36178,I2859,I35915,I36204,);
DFFARX1 I_1960 (I36204,I2859,I35915,I36221,);
not I_1961 (I35907,I36221);
not I_1962 (I36243,I36204);
nand I_1963 (I35892,I36243,I36082);
nor I_1964 (I36274,I109026,I109020);
not I_1965 (I36291,I36274);
nor I_1966 (I36308,I36243,I36291);
nor I_1967 (I36325,I35949,I36308);
DFFARX1 I_1968 (I36325,I2859,I35915,I35901,);
nor I_1969 (I36356,I36009,I36291);
nor I_1970 (I35889,I36204,I36356);
nor I_1971 (I35898,I36139,I36274);
nor I_1972 (I35886,I36009,I36274);
not I_1973 (I36442,I2866);
DFFARX1 I_1974 (I155165,I2859,I36442,I36468,);
not I_1975 (I36476,I36468);
nand I_1976 (I36493,I155147,I155162);
and I_1977 (I36510,I36493,I155138);
DFFARX1 I_1978 (I36510,I2859,I36442,I36536,);
DFFARX1 I_1979 (I155141,I2859,I36442,I36553,);
and I_1980 (I36561,I36553,I155156);
nor I_1981 (I36578,I36536,I36561);
DFFARX1 I_1982 (I36578,I2859,I36442,I36410,);
nand I_1983 (I36609,I36553,I155156);
nand I_1984 (I36626,I36476,I36609);
not I_1985 (I36422,I36626);
DFFARX1 I_1986 (I155159,I2859,I36442,I36666,);
DFFARX1 I_1987 (I36666,I2859,I36442,I36431,);
nand I_1988 (I36688,I155138,I155150);
and I_1989 (I36705,I36688,I155144);
DFFARX1 I_1990 (I36705,I2859,I36442,I36731,);
DFFARX1 I_1991 (I36731,I2859,I36442,I36748,);
not I_1992 (I36434,I36748);
not I_1993 (I36770,I36731);
nand I_1994 (I36419,I36770,I36609);
nor I_1995 (I36801,I155153,I155150);
not I_1996 (I36818,I36801);
nor I_1997 (I36835,I36770,I36818);
nor I_1998 (I36852,I36476,I36835);
DFFARX1 I_1999 (I36852,I2859,I36442,I36428,);
nor I_2000 (I36883,I36536,I36818);
nor I_2001 (I36416,I36731,I36883);
nor I_2002 (I36425,I36666,I36801);
nor I_2003 (I36413,I36536,I36801);
not I_2004 (I36969,I2866);
DFFARX1 I_2005 (I198506,I2859,I36969,I36995,);
not I_2006 (I37003,I36995);
nand I_2007 (I37020,I198500,I198491);
and I_2008 (I37037,I37020,I198512);
DFFARX1 I_2009 (I37037,I2859,I36969,I37063,);
DFFARX1 I_2010 (I198494,I2859,I36969,I37080,);
and I_2011 (I37088,I37080,I198488);
nor I_2012 (I37105,I37063,I37088);
DFFARX1 I_2013 (I37105,I2859,I36969,I36937,);
nand I_2014 (I37136,I37080,I198488);
nand I_2015 (I37153,I37003,I37136);
not I_2016 (I36949,I37153);
DFFARX1 I_2017 (I198488,I2859,I36969,I37193,);
DFFARX1 I_2018 (I37193,I2859,I36969,I36958,);
nand I_2019 (I37215,I198515,I198497);
and I_2020 (I37232,I37215,I198503);
DFFARX1 I_2021 (I37232,I2859,I36969,I37258,);
DFFARX1 I_2022 (I37258,I2859,I36969,I37275,);
not I_2023 (I36961,I37275);
not I_2024 (I37297,I37258);
nand I_2025 (I36946,I37297,I37136);
nor I_2026 (I37328,I198509,I198497);
not I_2027 (I37345,I37328);
nor I_2028 (I37362,I37297,I37345);
nor I_2029 (I37379,I37003,I37362);
DFFARX1 I_2030 (I37379,I2859,I36969,I36955,);
nor I_2031 (I37410,I37063,I37345);
nor I_2032 (I36943,I37258,I37410);
nor I_2033 (I36952,I37193,I37328);
nor I_2034 (I36940,I37063,I37328);
not I_2035 (I37496,I2866);
DFFARX1 I_2036 (I203693,I2859,I37496,I37522,);
not I_2037 (I37530,I37522);
nand I_2038 (I37547,I203714,I203708);
and I_2039 (I37564,I37547,I203690);
DFFARX1 I_2040 (I37564,I2859,I37496,I37590,);
DFFARX1 I_2041 (I203693,I2859,I37496,I37607,);
and I_2042 (I37615,I37607,I203702);
nor I_2043 (I37632,I37590,I37615);
DFFARX1 I_2044 (I37632,I2859,I37496,I37464,);
nand I_2045 (I37663,I37607,I203702);
nand I_2046 (I37680,I37530,I37663);
not I_2047 (I37476,I37680);
DFFARX1 I_2048 (I203699,I2859,I37496,I37720,);
DFFARX1 I_2049 (I37720,I2859,I37496,I37485,);
nand I_2050 (I37742,I203705,I203696);
and I_2051 (I37759,I37742,I203690);
DFFARX1 I_2052 (I37759,I2859,I37496,I37785,);
DFFARX1 I_2053 (I37785,I2859,I37496,I37802,);
not I_2054 (I37488,I37802);
not I_2055 (I37824,I37785);
nand I_2056 (I37473,I37824,I37663);
nor I_2057 (I37855,I203711,I203696);
not I_2058 (I37872,I37855);
nor I_2059 (I37889,I37824,I37872);
nor I_2060 (I37906,I37530,I37889);
DFFARX1 I_2061 (I37906,I2859,I37496,I37482,);
nor I_2062 (I37937,I37590,I37872);
nor I_2063 (I37470,I37785,I37937);
nor I_2064 (I37479,I37720,I37855);
nor I_2065 (I37467,I37590,I37855);
not I_2066 (I38023,I2866);
DFFARX1 I_2067 (I319129,I2859,I38023,I38049,);
not I_2068 (I38057,I38049);
nand I_2069 (I38074,I319126,I319141);
and I_2070 (I38091,I38074,I319123);
DFFARX1 I_2071 (I38091,I2859,I38023,I38117,);
DFFARX1 I_2072 (I319120,I2859,I38023,I38134,);
and I_2073 (I38142,I38134,I319120);
nor I_2074 (I38159,I38117,I38142);
DFFARX1 I_2075 (I38159,I2859,I38023,I37991,);
nand I_2076 (I38190,I38134,I319120);
nand I_2077 (I38207,I38057,I38190);
not I_2078 (I38003,I38207);
DFFARX1 I_2079 (I319123,I2859,I38023,I38247,);
DFFARX1 I_2080 (I38247,I2859,I38023,I38012,);
nand I_2081 (I38269,I319135,I319126);
and I_2082 (I38286,I38269,I319138);
DFFARX1 I_2083 (I38286,I2859,I38023,I38312,);
DFFARX1 I_2084 (I38312,I2859,I38023,I38329,);
not I_2085 (I38015,I38329);
not I_2086 (I38351,I38312);
nand I_2087 (I38000,I38351,I38190);
nor I_2088 (I38382,I319132,I319126);
not I_2089 (I38399,I38382);
nor I_2090 (I38416,I38351,I38399);
nor I_2091 (I38433,I38057,I38416);
DFFARX1 I_2092 (I38433,I2859,I38023,I38009,);
nor I_2093 (I38464,I38117,I38399);
nor I_2094 (I37997,I38312,I38464);
nor I_2095 (I38006,I38247,I38382);
nor I_2096 (I37994,I38117,I38382);
not I_2097 (I38550,I2866);
DFFARX1 I_2098 (I531620,I2859,I38550,I38576,);
not I_2099 (I38584,I38576);
nand I_2100 (I38601,I531626,I531644);
and I_2101 (I38618,I38601,I531641);
DFFARX1 I_2102 (I38618,I2859,I38550,I38644,);
DFFARX1 I_2103 (I531638,I2859,I38550,I38661,);
and I_2104 (I38669,I38661,I531632);
nor I_2105 (I38686,I38644,I38669);
DFFARX1 I_2106 (I38686,I2859,I38550,I38518,);
nand I_2107 (I38717,I38661,I531632);
nand I_2108 (I38734,I38584,I38717);
not I_2109 (I38530,I38734);
DFFARX1 I_2110 (I531620,I2859,I38550,I38774,);
DFFARX1 I_2111 (I38774,I2859,I38550,I38539,);
nand I_2112 (I38796,I531635,I531623);
and I_2113 (I38813,I38796,I531647);
DFFARX1 I_2114 (I38813,I2859,I38550,I38839,);
DFFARX1 I_2115 (I38839,I2859,I38550,I38856,);
not I_2116 (I38542,I38856);
not I_2117 (I38878,I38839);
nand I_2118 (I38527,I38878,I38717);
nor I_2119 (I38909,I531629,I531623);
not I_2120 (I38926,I38909);
nor I_2121 (I38943,I38878,I38926);
nor I_2122 (I38960,I38584,I38943);
DFFARX1 I_2123 (I38960,I2859,I38550,I38536,);
nor I_2124 (I38991,I38644,I38926);
nor I_2125 (I38524,I38839,I38991);
nor I_2126 (I38533,I38774,I38909);
nor I_2127 (I38521,I38644,I38909);
not I_2128 (I39077,I2866);
DFFARX1 I_2129 (I98319,I2859,I39077,I39103,);
not I_2130 (I39111,I39103);
nand I_2131 (I39128,I98313,I98307);
and I_2132 (I39145,I39128,I98328);
DFFARX1 I_2133 (I39145,I2859,I39077,I39171,);
DFFARX1 I_2134 (I98325,I2859,I39077,I39188,);
and I_2135 (I39196,I39188,I98322);
nor I_2136 (I39213,I39171,I39196);
DFFARX1 I_2137 (I39213,I2859,I39077,I39045,);
nand I_2138 (I39244,I39188,I98322);
nand I_2139 (I39261,I39111,I39244);
not I_2140 (I39057,I39261);
DFFARX1 I_2141 (I98307,I2859,I39077,I39301,);
DFFARX1 I_2142 (I39301,I2859,I39077,I39066,);
nand I_2143 (I39323,I98310,I98310);
and I_2144 (I39340,I39323,I98331);
DFFARX1 I_2145 (I39340,I2859,I39077,I39366,);
DFFARX1 I_2146 (I39366,I2859,I39077,I39383,);
not I_2147 (I39069,I39383);
not I_2148 (I39405,I39366);
nand I_2149 (I39054,I39405,I39244);
nor I_2150 (I39436,I98316,I98310);
not I_2151 (I39453,I39436);
nor I_2152 (I39470,I39405,I39453);
nor I_2153 (I39487,I39111,I39470);
DFFARX1 I_2154 (I39487,I2859,I39077,I39063,);
nor I_2155 (I39518,I39171,I39453);
nor I_2156 (I39051,I39366,I39518);
nor I_2157 (I39060,I39301,I39436);
nor I_2158 (I39048,I39171,I39436);
not I_2159 (I39604,I2866);
DFFARX1 I_2160 (I69164,I2859,I39604,I39630,);
not I_2161 (I39638,I39630);
nand I_2162 (I39655,I69158,I69152);
and I_2163 (I39672,I39655,I69173);
DFFARX1 I_2164 (I39672,I2859,I39604,I39698,);
DFFARX1 I_2165 (I69170,I2859,I39604,I39715,);
and I_2166 (I39723,I39715,I69167);
nor I_2167 (I39740,I39698,I39723);
DFFARX1 I_2168 (I39740,I2859,I39604,I39572,);
nand I_2169 (I39771,I39715,I69167);
nand I_2170 (I39788,I39638,I39771);
not I_2171 (I39584,I39788);
DFFARX1 I_2172 (I69152,I2859,I39604,I39828,);
DFFARX1 I_2173 (I39828,I2859,I39604,I39593,);
nand I_2174 (I39850,I69155,I69155);
and I_2175 (I39867,I39850,I69176);
DFFARX1 I_2176 (I39867,I2859,I39604,I39893,);
DFFARX1 I_2177 (I39893,I2859,I39604,I39910,);
not I_2178 (I39596,I39910);
not I_2179 (I39932,I39893);
nand I_2180 (I39581,I39932,I39771);
nor I_2181 (I39963,I69161,I69155);
not I_2182 (I39980,I39963);
nor I_2183 (I39997,I39932,I39980);
nor I_2184 (I40014,I39638,I39997);
DFFARX1 I_2185 (I40014,I2859,I39604,I39590,);
nor I_2186 (I40045,I39698,I39980);
nor I_2187 (I39578,I39893,I40045);
nor I_2188 (I39587,I39828,I39963);
nor I_2189 (I39575,I39698,I39963);
not I_2190 (I40131,I2866);
DFFARX1 I_2191 (I530485,I2859,I40131,I40157,);
not I_2192 (I40165,I40157);
nand I_2193 (I40182,I530488,I530482);
and I_2194 (I40199,I40182,I530479);
DFFARX1 I_2195 (I40199,I2859,I40131,I40225,);
DFFARX1 I_2196 (I530464,I2859,I40131,I40242,);
and I_2197 (I40250,I40242,I530473);
nor I_2198 (I40267,I40225,I40250);
DFFARX1 I_2199 (I40267,I2859,I40131,I40099,);
nand I_2200 (I40298,I40242,I530473);
nand I_2201 (I40315,I40165,I40298);
not I_2202 (I40111,I40315);
DFFARX1 I_2203 (I530464,I2859,I40131,I40355,);
DFFARX1 I_2204 (I40355,I2859,I40131,I40120,);
nand I_2205 (I40377,I530467,I530470);
and I_2206 (I40394,I40377,I530476);
DFFARX1 I_2207 (I40394,I2859,I40131,I40420,);
DFFARX1 I_2208 (I40420,I2859,I40131,I40437,);
not I_2209 (I40123,I40437);
not I_2210 (I40459,I40420);
nand I_2211 (I40108,I40459,I40298);
nor I_2212 (I40490,I530467,I530470);
not I_2213 (I40507,I40490);
nor I_2214 (I40524,I40459,I40507);
nor I_2215 (I40541,I40165,I40524);
DFFARX1 I_2216 (I40541,I2859,I40131,I40117,);
nor I_2217 (I40572,I40225,I40507);
nor I_2218 (I40105,I40420,I40572);
nor I_2219 (I40114,I40355,I40490);
nor I_2220 (I40102,I40225,I40490);
not I_2221 (I40658,I2866);
DFFARX1 I_2222 (I517769,I2859,I40658,I40684,);
not I_2223 (I40692,I40684);
nand I_2224 (I40709,I517772,I517766);
and I_2225 (I40726,I40709,I517763);
DFFARX1 I_2226 (I40726,I2859,I40658,I40752,);
DFFARX1 I_2227 (I517748,I2859,I40658,I40769,);
and I_2228 (I40777,I40769,I517757);
nor I_2229 (I40794,I40752,I40777);
DFFARX1 I_2230 (I40794,I2859,I40658,I40626,);
nand I_2231 (I40825,I40769,I517757);
nand I_2232 (I40842,I40692,I40825);
not I_2233 (I40638,I40842);
DFFARX1 I_2234 (I517748,I2859,I40658,I40882,);
DFFARX1 I_2235 (I40882,I2859,I40658,I40647,);
nand I_2236 (I40904,I517751,I517754);
and I_2237 (I40921,I40904,I517760);
DFFARX1 I_2238 (I40921,I2859,I40658,I40947,);
DFFARX1 I_2239 (I40947,I2859,I40658,I40964,);
not I_2240 (I40650,I40964);
not I_2241 (I40986,I40947);
nand I_2242 (I40635,I40986,I40825);
nor I_2243 (I41017,I517751,I517754);
not I_2244 (I41034,I41017);
nor I_2245 (I41051,I40986,I41034);
nor I_2246 (I41068,I40692,I41051);
DFFARX1 I_2247 (I41068,I2859,I40658,I40644,);
nor I_2248 (I41099,I40752,I41034);
nor I_2249 (I40632,I40947,I41099);
nor I_2250 (I40641,I40882,I41017);
nor I_2251 (I40629,I40752,I41017);
not I_2252 (I41185,I2866);
DFFARX1 I_2253 (I293224,I2859,I41185,I41211,);
not I_2254 (I41219,I41211);
nand I_2255 (I41236,I293215,I293233);
and I_2256 (I41253,I41236,I293212);
DFFARX1 I_2257 (I41253,I2859,I41185,I41279,);
DFFARX1 I_2258 (I293215,I2859,I41185,I41296,);
and I_2259 (I41304,I41296,I293218);
nor I_2260 (I41321,I41279,I41304);
DFFARX1 I_2261 (I41321,I2859,I41185,I41153,);
nand I_2262 (I41352,I41296,I293218);
nand I_2263 (I41369,I41219,I41352);
not I_2264 (I41165,I41369);
DFFARX1 I_2265 (I293212,I2859,I41185,I41409,);
DFFARX1 I_2266 (I41409,I2859,I41185,I41174,);
nand I_2267 (I41431,I293230,I293221);
and I_2268 (I41448,I41431,I293236);
DFFARX1 I_2269 (I41448,I2859,I41185,I41474,);
DFFARX1 I_2270 (I41474,I2859,I41185,I41491,);
not I_2271 (I41177,I41491);
not I_2272 (I41513,I41474);
nand I_2273 (I41162,I41513,I41352);
nor I_2274 (I41544,I293227,I293221);
not I_2275 (I41561,I41544);
nor I_2276 (I41578,I41513,I41561);
nor I_2277 (I41595,I41219,I41578);
DFFARX1 I_2278 (I41595,I2859,I41185,I41171,);
nor I_2279 (I41626,I41279,I41561);
nor I_2280 (I41159,I41474,I41626);
nor I_2281 (I41168,I41409,I41544);
nor I_2282 (I41156,I41279,I41544);
not I_2283 (I41712,I2866);
DFFARX1 I_2284 (I387656,I2859,I41712,I41738,);
not I_2285 (I41746,I41738);
nand I_2286 (I41763,I387674,I387668);
and I_2287 (I41780,I41763,I387647);
DFFARX1 I_2288 (I41780,I2859,I41712,I41806,);
DFFARX1 I_2289 (I387665,I2859,I41712,I41823,);
and I_2290 (I41831,I41823,I387650);
nor I_2291 (I41848,I41806,I41831);
DFFARX1 I_2292 (I41848,I2859,I41712,I41680,);
nand I_2293 (I41879,I41823,I387650);
nand I_2294 (I41896,I41746,I41879);
not I_2295 (I41692,I41896);
DFFARX1 I_2296 (I387662,I2859,I41712,I41936,);
DFFARX1 I_2297 (I41936,I2859,I41712,I41701,);
nand I_2298 (I41958,I387671,I387659);
and I_2299 (I41975,I41958,I387653);
DFFARX1 I_2300 (I41975,I2859,I41712,I42001,);
DFFARX1 I_2301 (I42001,I2859,I41712,I42018,);
not I_2302 (I41704,I42018);
not I_2303 (I42040,I42001);
nand I_2304 (I41689,I42040,I41879);
nor I_2305 (I42071,I387647,I387659);
not I_2306 (I42088,I42071);
nor I_2307 (I42105,I42040,I42088);
nor I_2308 (I42122,I41746,I42105);
DFFARX1 I_2309 (I42122,I2859,I41712,I41698,);
nor I_2310 (I42153,I41806,I42088);
nor I_2311 (I41686,I42001,I42153);
nor I_2312 (I41695,I41936,I42071);
nor I_2313 (I41683,I41806,I42071);
not I_2314 (I42239,I2866);
DFFARX1 I_2315 (I321237,I2859,I42239,I42265,);
not I_2316 (I42273,I42265);
nand I_2317 (I42290,I321234,I321249);
and I_2318 (I42307,I42290,I321231);
DFFARX1 I_2319 (I42307,I2859,I42239,I42333,);
DFFARX1 I_2320 (I321228,I2859,I42239,I42350,);
and I_2321 (I42358,I42350,I321228);
nor I_2322 (I42375,I42333,I42358);
DFFARX1 I_2323 (I42375,I2859,I42239,I42207,);
nand I_2324 (I42406,I42350,I321228);
nand I_2325 (I42423,I42273,I42406);
not I_2326 (I42219,I42423);
DFFARX1 I_2327 (I321231,I2859,I42239,I42463,);
DFFARX1 I_2328 (I42463,I2859,I42239,I42228,);
nand I_2329 (I42485,I321243,I321234);
and I_2330 (I42502,I42485,I321246);
DFFARX1 I_2331 (I42502,I2859,I42239,I42528,);
DFFARX1 I_2332 (I42528,I2859,I42239,I42545,);
not I_2333 (I42231,I42545);
not I_2334 (I42567,I42528);
nand I_2335 (I42216,I42567,I42406);
nor I_2336 (I42598,I321240,I321234);
not I_2337 (I42615,I42598);
nor I_2338 (I42632,I42567,I42615);
nor I_2339 (I42649,I42273,I42632);
DFFARX1 I_2340 (I42649,I2859,I42239,I42225,);
nor I_2341 (I42680,I42333,I42615);
nor I_2342 (I42213,I42528,I42680);
nor I_2343 (I42222,I42463,I42598);
nor I_2344 (I42210,I42333,I42598);
not I_2345 (I42766,I2866);
DFFARX1 I_2346 (I423758,I2859,I42766,I42792,);
not I_2347 (I42800,I42792);
nand I_2348 (I42817,I423755,I423761);
and I_2349 (I42834,I42817,I423758);
DFFARX1 I_2350 (I42834,I2859,I42766,I42860,);
DFFARX1 I_2351 (I423761,I2859,I42766,I42877,);
and I_2352 (I42885,I42877,I423755);
nor I_2353 (I42902,I42860,I42885);
DFFARX1 I_2354 (I42902,I2859,I42766,I42734,);
nand I_2355 (I42933,I42877,I423755);
nand I_2356 (I42950,I42800,I42933);
not I_2357 (I42746,I42950);
DFFARX1 I_2358 (I423764,I2859,I42766,I42990,);
DFFARX1 I_2359 (I42990,I2859,I42766,I42755,);
nand I_2360 (I43012,I423767,I423776);
and I_2361 (I43029,I43012,I423770);
DFFARX1 I_2362 (I43029,I2859,I42766,I43055,);
DFFARX1 I_2363 (I43055,I2859,I42766,I43072,);
not I_2364 (I42758,I43072);
not I_2365 (I43094,I43055);
nand I_2366 (I42743,I43094,I42933);
nor I_2367 (I43125,I423773,I423776);
not I_2368 (I43142,I43125);
nor I_2369 (I43159,I43094,I43142);
nor I_2370 (I43176,I42800,I43159);
DFFARX1 I_2371 (I43176,I2859,I42766,I42752,);
nor I_2372 (I43207,I42860,I43142);
nor I_2373 (I42740,I43055,I43207);
nor I_2374 (I42749,I42990,I43125);
nor I_2375 (I42737,I42860,I43125);
not I_2376 (I43293,I2866);
DFFARX1 I_2377 (I316922,I2859,I43293,I43319,);
not I_2378 (I43327,I43319);
nand I_2379 (I43344,I316913,I316931);
and I_2380 (I43361,I43344,I316910);
DFFARX1 I_2381 (I43361,I2859,I43293,I43387,);
DFFARX1 I_2382 (I316913,I2859,I43293,I43404,);
and I_2383 (I43412,I43404,I316916);
nor I_2384 (I43429,I43387,I43412);
DFFARX1 I_2385 (I43429,I2859,I43293,I43261,);
nand I_2386 (I43460,I43404,I316916);
nand I_2387 (I43477,I43327,I43460);
not I_2388 (I43273,I43477);
DFFARX1 I_2389 (I316910,I2859,I43293,I43517,);
DFFARX1 I_2390 (I43517,I2859,I43293,I43282,);
nand I_2391 (I43539,I316928,I316919);
and I_2392 (I43556,I43539,I316934);
DFFARX1 I_2393 (I43556,I2859,I43293,I43582,);
DFFARX1 I_2394 (I43582,I2859,I43293,I43599,);
not I_2395 (I43285,I43599);
not I_2396 (I43621,I43582);
nand I_2397 (I43270,I43621,I43460);
nor I_2398 (I43652,I316925,I316919);
not I_2399 (I43669,I43652);
nor I_2400 (I43686,I43621,I43669);
nor I_2401 (I43703,I43327,I43686);
DFFARX1 I_2402 (I43703,I2859,I43293,I43279,);
nor I_2403 (I43734,I43387,I43669);
nor I_2404 (I43267,I43582,I43734);
nor I_2405 (I43276,I43517,I43652);
nor I_2406 (I43264,I43387,I43652);
not I_2407 (I43820,I2866);
DFFARX1 I_2408 (I89394,I2859,I43820,I43846,);
not I_2409 (I43854,I43846);
nand I_2410 (I43871,I89388,I89382);
and I_2411 (I43888,I43871,I89403);
DFFARX1 I_2412 (I43888,I2859,I43820,I43914,);
DFFARX1 I_2413 (I89400,I2859,I43820,I43931,);
and I_2414 (I43939,I43931,I89397);
nor I_2415 (I43956,I43914,I43939);
DFFARX1 I_2416 (I43956,I2859,I43820,I43788,);
nand I_2417 (I43987,I43931,I89397);
nand I_2418 (I44004,I43854,I43987);
not I_2419 (I43800,I44004);
DFFARX1 I_2420 (I89382,I2859,I43820,I44044,);
DFFARX1 I_2421 (I44044,I2859,I43820,I43809,);
nand I_2422 (I44066,I89385,I89385);
and I_2423 (I44083,I44066,I89406);
DFFARX1 I_2424 (I44083,I2859,I43820,I44109,);
DFFARX1 I_2425 (I44109,I2859,I43820,I44126,);
not I_2426 (I43812,I44126);
not I_2427 (I44148,I44109);
nand I_2428 (I43797,I44148,I43987);
nor I_2429 (I44179,I89391,I89385);
not I_2430 (I44196,I44179);
nor I_2431 (I44213,I44148,I44196);
nor I_2432 (I44230,I43854,I44213);
DFFARX1 I_2433 (I44230,I2859,I43820,I43806,);
nor I_2434 (I44261,I43914,I44196);
nor I_2435 (I43794,I44109,I44261);
nor I_2436 (I43803,I44044,I44179);
nor I_2437 (I43791,I43914,I44179);
not I_2438 (I44347,I2866);
DFFARX1 I_2439 (I463184,I2859,I44347,I44373,);
not I_2440 (I44381,I44373);
nand I_2441 (I44398,I463199,I463178);
and I_2442 (I44415,I44398,I463181);
DFFARX1 I_2443 (I44415,I2859,I44347,I44441,);
DFFARX1 I_2444 (I463202,I2859,I44347,I44458,);
and I_2445 (I44466,I44458,I463181);
nor I_2446 (I44483,I44441,I44466);
DFFARX1 I_2447 (I44483,I2859,I44347,I44315,);
nand I_2448 (I44514,I44458,I463181);
nand I_2449 (I44531,I44381,I44514);
not I_2450 (I44327,I44531);
DFFARX1 I_2451 (I463178,I2859,I44347,I44571,);
DFFARX1 I_2452 (I44571,I2859,I44347,I44336,);
nand I_2453 (I44593,I463190,I463187);
and I_2454 (I44610,I44593,I463193);
DFFARX1 I_2455 (I44610,I2859,I44347,I44636,);
DFFARX1 I_2456 (I44636,I2859,I44347,I44653,);
not I_2457 (I44339,I44653);
not I_2458 (I44675,I44636);
nand I_2459 (I44324,I44675,I44514);
nor I_2460 (I44706,I463196,I463187);
not I_2461 (I44723,I44706);
nor I_2462 (I44740,I44675,I44723);
nor I_2463 (I44757,I44381,I44740);
DFFARX1 I_2464 (I44757,I2859,I44347,I44333,);
nor I_2465 (I44788,I44441,I44723);
nor I_2466 (I44321,I44636,I44788);
nor I_2467 (I44330,I44571,I44706);
nor I_2468 (I44318,I44441,I44706);
not I_2469 (I44874,I2866);
DFFARX1 I_2470 (I428807,I2859,I44874,I44900,);
not I_2471 (I44908,I44900);
nand I_2472 (I44925,I428804,I428810);
and I_2473 (I44942,I44925,I428807);
DFFARX1 I_2474 (I44942,I2859,I44874,I44968,);
DFFARX1 I_2475 (I428810,I2859,I44874,I44985,);
and I_2476 (I44993,I44985,I428804);
nor I_2477 (I45010,I44968,I44993);
DFFARX1 I_2478 (I45010,I2859,I44874,I44842,);
nand I_2479 (I45041,I44985,I428804);
nand I_2480 (I45058,I44908,I45041);
not I_2481 (I44854,I45058);
DFFARX1 I_2482 (I428813,I2859,I44874,I45098,);
DFFARX1 I_2483 (I45098,I2859,I44874,I44863,);
nand I_2484 (I45120,I428816,I428825);
and I_2485 (I45137,I45120,I428819);
DFFARX1 I_2486 (I45137,I2859,I44874,I45163,);
DFFARX1 I_2487 (I45163,I2859,I44874,I45180,);
not I_2488 (I44866,I45180);
not I_2489 (I45202,I45163);
nand I_2490 (I44851,I45202,I45041);
nor I_2491 (I45233,I428822,I428825);
not I_2492 (I45250,I45233);
nor I_2493 (I45267,I45202,I45250);
nor I_2494 (I45284,I44908,I45267);
DFFARX1 I_2495 (I45284,I2859,I44874,I44860,);
nor I_2496 (I45315,I44968,I45250);
nor I_2497 (I44848,I45163,I45315);
nor I_2498 (I44857,I45098,I45233);
nor I_2499 (I44845,I44968,I45233);
not I_2500 (I45401,I2866);
DFFARX1 I_2501 (I220948,I2859,I45401,I45427,);
not I_2502 (I45435,I45427);
nand I_2503 (I45452,I220969,I220963);
and I_2504 (I45469,I45452,I220945);
DFFARX1 I_2505 (I45469,I2859,I45401,I45495,);
DFFARX1 I_2506 (I220948,I2859,I45401,I45512,);
and I_2507 (I45520,I45512,I220957);
nor I_2508 (I45537,I45495,I45520);
DFFARX1 I_2509 (I45537,I2859,I45401,I45369,);
nand I_2510 (I45568,I45512,I220957);
nand I_2511 (I45585,I45435,I45568);
not I_2512 (I45381,I45585);
DFFARX1 I_2513 (I220954,I2859,I45401,I45625,);
DFFARX1 I_2514 (I45625,I2859,I45401,I45390,);
nand I_2515 (I45647,I220960,I220951);
and I_2516 (I45664,I45647,I220945);
DFFARX1 I_2517 (I45664,I2859,I45401,I45690,);
DFFARX1 I_2518 (I45690,I2859,I45401,I45707,);
not I_2519 (I45393,I45707);
not I_2520 (I45729,I45690);
nand I_2521 (I45378,I45729,I45568);
nor I_2522 (I45760,I220966,I220951);
not I_2523 (I45777,I45760);
nor I_2524 (I45794,I45729,I45777);
nor I_2525 (I45811,I45435,I45794);
DFFARX1 I_2526 (I45811,I2859,I45401,I45387,);
nor I_2527 (I45842,I45495,I45777);
nor I_2528 (I45375,I45690,I45842);
nor I_2529 (I45384,I45625,I45760);
nor I_2530 (I45372,I45495,I45760);
not I_2531 (I45928,I2866);
DFFARX1 I_2532 (I532742,I2859,I45928,I45954,);
not I_2533 (I45962,I45954);
nand I_2534 (I45979,I532748,I532766);
and I_2535 (I45996,I45979,I532763);
DFFARX1 I_2536 (I45996,I2859,I45928,I46022,);
DFFARX1 I_2537 (I532760,I2859,I45928,I46039,);
and I_2538 (I46047,I46039,I532754);
nor I_2539 (I46064,I46022,I46047);
DFFARX1 I_2540 (I46064,I2859,I45928,I45896,);
nand I_2541 (I46095,I46039,I532754);
nand I_2542 (I46112,I45962,I46095);
not I_2543 (I45908,I46112);
DFFARX1 I_2544 (I532742,I2859,I45928,I46152,);
DFFARX1 I_2545 (I46152,I2859,I45928,I45917,);
nand I_2546 (I46174,I532757,I532745);
and I_2547 (I46191,I46174,I532769);
DFFARX1 I_2548 (I46191,I2859,I45928,I46217,);
DFFARX1 I_2549 (I46217,I2859,I45928,I46234,);
not I_2550 (I45920,I46234);
not I_2551 (I46256,I46217);
nand I_2552 (I45905,I46256,I46095);
nor I_2553 (I46287,I532751,I532745);
not I_2554 (I46304,I46287);
nor I_2555 (I46321,I46256,I46304);
nor I_2556 (I46338,I45962,I46321);
DFFARX1 I_2557 (I46338,I2859,I45928,I45914,);
nor I_2558 (I46369,I46022,I46304);
nor I_2559 (I45902,I46217,I46369);
nor I_2560 (I45911,I46152,I46287);
nor I_2561 (I45899,I46022,I46287);
not I_2562 (I46455,I2866);
DFFARX1 I_2563 (I81659,I2859,I46455,I46481,);
not I_2564 (I46489,I46481);
nand I_2565 (I46506,I81653,I81647);
and I_2566 (I46523,I46506,I81668);
DFFARX1 I_2567 (I46523,I2859,I46455,I46549,);
DFFARX1 I_2568 (I81665,I2859,I46455,I46566,);
and I_2569 (I46574,I46566,I81662);
nor I_2570 (I46591,I46549,I46574);
DFFARX1 I_2571 (I46591,I2859,I46455,I46423,);
nand I_2572 (I46622,I46566,I81662);
nand I_2573 (I46639,I46489,I46622);
not I_2574 (I46435,I46639);
DFFARX1 I_2575 (I81647,I2859,I46455,I46679,);
DFFARX1 I_2576 (I46679,I2859,I46455,I46444,);
nand I_2577 (I46701,I81650,I81650);
and I_2578 (I46718,I46701,I81671);
DFFARX1 I_2579 (I46718,I2859,I46455,I46744,);
DFFARX1 I_2580 (I46744,I2859,I46455,I46761,);
not I_2581 (I46447,I46761);
not I_2582 (I46783,I46744);
nand I_2583 (I46432,I46783,I46622);
nor I_2584 (I46814,I81656,I81650);
not I_2585 (I46831,I46814);
nor I_2586 (I46848,I46783,I46831);
nor I_2587 (I46865,I46489,I46848);
DFFARX1 I_2588 (I46865,I2859,I46455,I46441,);
nor I_2589 (I46896,I46549,I46831);
nor I_2590 (I46429,I46744,I46896);
nor I_2591 (I46438,I46679,I46814);
nor I_2592 (I46426,I46549,I46814);
not I_2593 (I46982,I2866);
DFFARX1 I_2594 (I311720,I2859,I46982,I47008,);
not I_2595 (I47016,I47008);
nand I_2596 (I47033,I311711,I311729);
and I_2597 (I47050,I47033,I311708);
DFFARX1 I_2598 (I47050,I2859,I46982,I47076,);
DFFARX1 I_2599 (I311711,I2859,I46982,I47093,);
and I_2600 (I47101,I47093,I311714);
nor I_2601 (I47118,I47076,I47101);
DFFARX1 I_2602 (I47118,I2859,I46982,I46950,);
nand I_2603 (I47149,I47093,I311714);
nand I_2604 (I47166,I47016,I47149);
not I_2605 (I46962,I47166);
DFFARX1 I_2606 (I311708,I2859,I46982,I47206,);
DFFARX1 I_2607 (I47206,I2859,I46982,I46971,);
nand I_2608 (I47228,I311726,I311717);
and I_2609 (I47245,I47228,I311732);
DFFARX1 I_2610 (I47245,I2859,I46982,I47271,);
DFFARX1 I_2611 (I47271,I2859,I46982,I47288,);
not I_2612 (I46974,I47288);
not I_2613 (I47310,I47271);
nand I_2614 (I46959,I47310,I47149);
nor I_2615 (I47341,I311723,I311717);
not I_2616 (I47358,I47341);
nor I_2617 (I47375,I47310,I47358);
nor I_2618 (I47392,I47016,I47375);
DFFARX1 I_2619 (I47392,I2859,I46982,I46968,);
nor I_2620 (I47423,I47076,I47358);
nor I_2621 (I46956,I47271,I47423);
nor I_2622 (I46965,I47206,I47341);
nor I_2623 (I46953,I47076,I47341);
not I_2624 (I47509,I2866);
DFFARX1 I_2625 (I396700,I2859,I47509,I47535,);
not I_2626 (I47543,I47535);
nand I_2627 (I47560,I396718,I396712);
and I_2628 (I47577,I47560,I396691);
DFFARX1 I_2629 (I47577,I2859,I47509,I47603,);
DFFARX1 I_2630 (I396709,I2859,I47509,I47620,);
and I_2631 (I47628,I47620,I396694);
nor I_2632 (I47645,I47603,I47628);
DFFARX1 I_2633 (I47645,I2859,I47509,I47477,);
nand I_2634 (I47676,I47620,I396694);
nand I_2635 (I47693,I47543,I47676);
not I_2636 (I47489,I47693);
DFFARX1 I_2637 (I396706,I2859,I47509,I47733,);
DFFARX1 I_2638 (I47733,I2859,I47509,I47498,);
nand I_2639 (I47755,I396715,I396703);
and I_2640 (I47772,I47755,I396697);
DFFARX1 I_2641 (I47772,I2859,I47509,I47798,);
DFFARX1 I_2642 (I47798,I2859,I47509,I47815,);
not I_2643 (I47501,I47815);
not I_2644 (I47837,I47798);
nand I_2645 (I47486,I47837,I47676);
nor I_2646 (I47868,I396691,I396703);
not I_2647 (I47885,I47868);
nor I_2648 (I47902,I47837,I47885);
nor I_2649 (I47919,I47543,I47902);
DFFARX1 I_2650 (I47919,I2859,I47509,I47495,);
nor I_2651 (I47950,I47603,I47885);
nor I_2652 (I47483,I47798,I47950);
nor I_2653 (I47492,I47733,I47868);
nor I_2654 (I47480,I47603,I47868);
not I_2655 (I48036,I2866);
DFFARX1 I_2656 (I566567,I2859,I48036,I48062,);
not I_2657 (I48070,I48062);
nand I_2658 (I48087,I566561,I566582);
and I_2659 (I48104,I48087,I566558);
DFFARX1 I_2660 (I48104,I2859,I48036,I48130,);
DFFARX1 I_2661 (I566579,I2859,I48036,I48147,);
and I_2662 (I48155,I48147,I566576);
nor I_2663 (I48172,I48130,I48155);
DFFARX1 I_2664 (I48172,I2859,I48036,I48004,);
nand I_2665 (I48203,I48147,I566576);
nand I_2666 (I48220,I48070,I48203);
not I_2667 (I48016,I48220);
DFFARX1 I_2668 (I566564,I2859,I48036,I48260,);
DFFARX1 I_2669 (I48260,I2859,I48036,I48025,);
nand I_2670 (I48282,I566573,I566570);
and I_2671 (I48299,I48282,I566555);
DFFARX1 I_2672 (I48299,I2859,I48036,I48325,);
DFFARX1 I_2673 (I48325,I2859,I48036,I48342,);
not I_2674 (I48028,I48342);
not I_2675 (I48364,I48325);
nand I_2676 (I48013,I48364,I48203);
nor I_2677 (I48395,I566555,I566570);
not I_2678 (I48412,I48395);
nor I_2679 (I48429,I48364,I48412);
nor I_2680 (I48446,I48070,I48429);
DFFARX1 I_2681 (I48446,I2859,I48036,I48022,);
nor I_2682 (I48477,I48130,I48412);
nor I_2683 (I48010,I48325,I48477);
nor I_2684 (I48019,I48260,I48395);
nor I_2685 (I48007,I48130,I48395);
not I_2686 (I48563,I2866);
DFFARX1 I_2687 (I274150,I2859,I48563,I48589,);
not I_2688 (I48597,I48589);
nand I_2689 (I48614,I274141,I274159);
and I_2690 (I48631,I48614,I274138);
DFFARX1 I_2691 (I48631,I2859,I48563,I48657,);
DFFARX1 I_2692 (I274141,I2859,I48563,I48674,);
and I_2693 (I48682,I48674,I274144);
nor I_2694 (I48699,I48657,I48682);
DFFARX1 I_2695 (I48699,I2859,I48563,I48531,);
nand I_2696 (I48730,I48674,I274144);
nand I_2697 (I48747,I48597,I48730);
not I_2698 (I48543,I48747);
DFFARX1 I_2699 (I274138,I2859,I48563,I48787,);
DFFARX1 I_2700 (I48787,I2859,I48563,I48552,);
nand I_2701 (I48809,I274156,I274147);
and I_2702 (I48826,I48809,I274162);
DFFARX1 I_2703 (I48826,I2859,I48563,I48852,);
DFFARX1 I_2704 (I48852,I2859,I48563,I48869,);
not I_2705 (I48555,I48869);
not I_2706 (I48891,I48852);
nand I_2707 (I48540,I48891,I48730);
nor I_2708 (I48922,I274153,I274147);
not I_2709 (I48939,I48922);
nor I_2710 (I48956,I48891,I48939);
nor I_2711 (I48973,I48597,I48956);
DFFARX1 I_2712 (I48973,I2859,I48563,I48549,);
nor I_2713 (I49004,I48657,I48939);
nor I_2714 (I48537,I48852,I49004);
nor I_2715 (I48546,I48787,I48922);
nor I_2716 (I48534,I48657,I48922);
not I_2717 (I49090,I2866);
DFFARX1 I_2718 (I550502,I2859,I49090,I49116,);
not I_2719 (I49124,I49116);
nand I_2720 (I49141,I550496,I550517);
and I_2721 (I49158,I49141,I550493);
DFFARX1 I_2722 (I49158,I2859,I49090,I49184,);
DFFARX1 I_2723 (I550514,I2859,I49090,I49201,);
and I_2724 (I49209,I49201,I550511);
nor I_2725 (I49226,I49184,I49209);
DFFARX1 I_2726 (I49226,I2859,I49090,I49058,);
nand I_2727 (I49257,I49201,I550511);
nand I_2728 (I49274,I49124,I49257);
not I_2729 (I49070,I49274);
DFFARX1 I_2730 (I550499,I2859,I49090,I49314,);
DFFARX1 I_2731 (I49314,I2859,I49090,I49079,);
nand I_2732 (I49336,I550508,I550505);
and I_2733 (I49353,I49336,I550490);
DFFARX1 I_2734 (I49353,I2859,I49090,I49379,);
DFFARX1 I_2735 (I49379,I2859,I49090,I49396,);
not I_2736 (I49082,I49396);
not I_2737 (I49418,I49379);
nand I_2738 (I49067,I49418,I49257);
nor I_2739 (I49449,I550490,I550505);
not I_2740 (I49466,I49449);
nor I_2741 (I49483,I49418,I49466);
nor I_2742 (I49500,I49124,I49483);
DFFARX1 I_2743 (I49500,I2859,I49090,I49076,);
nor I_2744 (I49531,I49184,I49466);
nor I_2745 (I49064,I49379,I49531);
nor I_2746 (I49073,I49314,I49449);
nor I_2747 (I49061,I49184,I49449);
not I_2748 (I49617,I2866);
DFFARX1 I_2749 (I486882,I2859,I49617,I49643,);
not I_2750 (I49651,I49643);
nand I_2751 (I49668,I486897,I486876);
and I_2752 (I49685,I49668,I486879);
DFFARX1 I_2753 (I49685,I2859,I49617,I49711,);
DFFARX1 I_2754 (I486900,I2859,I49617,I49728,);
and I_2755 (I49736,I49728,I486879);
nor I_2756 (I49753,I49711,I49736);
DFFARX1 I_2757 (I49753,I2859,I49617,I49585,);
nand I_2758 (I49784,I49728,I486879);
nand I_2759 (I49801,I49651,I49784);
not I_2760 (I49597,I49801);
DFFARX1 I_2761 (I486876,I2859,I49617,I49841,);
DFFARX1 I_2762 (I49841,I2859,I49617,I49606,);
nand I_2763 (I49863,I486888,I486885);
and I_2764 (I49880,I49863,I486891);
DFFARX1 I_2765 (I49880,I2859,I49617,I49906,);
DFFARX1 I_2766 (I49906,I2859,I49617,I49923,);
not I_2767 (I49609,I49923);
not I_2768 (I49945,I49906);
nand I_2769 (I49594,I49945,I49784);
nor I_2770 (I49976,I486894,I486885);
not I_2771 (I49993,I49976);
nor I_2772 (I50010,I49945,I49993);
nor I_2773 (I50027,I49651,I50010);
DFFARX1 I_2774 (I50027,I2859,I49617,I49603,);
nor I_2775 (I50058,I49711,I49993);
nor I_2776 (I49591,I49906,I50058);
nor I_2777 (I49600,I49841,I49976);
nor I_2778 (I49588,I49711,I49976);
not I_2779 (I50147,I2866);
DFFARX1 I_2780 (I112460,I2859,I50147,I50173,);
not I_2781 (I50181,I50173);
DFFARX1 I_2782 (I112457,I2859,I50147,I50207,);
not I_2783 (I50215,I112454);
or I_2784 (I50232,I112466,I112454);
nor I_2785 (I50249,I50207,I112466);
nand I_2786 (I50124,I50215,I50249);
nor I_2787 (I50280,I112475,I112466);
nand I_2788 (I50118,I50280,I50215);
not I_2789 (I50311,I112472);
nand I_2790 (I50328,I50215,I50311);
nor I_2791 (I50345,I112451,I112451);
not I_2792 (I50362,I50345);
nor I_2793 (I50379,I50362,I50328);
nor I_2794 (I50396,I50280,I50379);
DFFARX1 I_2795 (I50396,I2859,I50147,I50133,);
nor I_2796 (I50130,I50345,I50232);
DFFARX1 I_2797 (I50345,I2859,I50147,I50136,);
nor I_2798 (I50455,I50311,I112451);
nor I_2799 (I50472,I50455,I112454);
nor I_2800 (I50489,I112463,I112478);
DFFARX1 I_2801 (I50489,I2859,I50147,I50515,);
nor I_2802 (I50115,I50515,I50472);
DFFARX1 I_2803 (I50515,I2859,I50147,I50546,);
nand I_2804 (I50554,I50546,I112469);
nor I_2805 (I50139,I50181,I50554);
not I_2806 (I50585,I50515);
nand I_2807 (I50602,I50585,I112469);
nor I_2808 (I50619,I50181,I50602);
nor I_2809 (I50121,I50207,I50619);
nor I_2810 (I50650,I112463,I112475);
nor I_2811 (I50667,I50207,I50650);
DFFARX1 I_2812 (I50667,I2859,I50147,I50112,);
and I_2813 (I50127,I50280,I112463);
not I_2814 (I50742,I2866);
DFFARX1 I_2815 (I216197,I2859,I50742,I50768,);
not I_2816 (I50776,I50768);
DFFARX1 I_2817 (I216203,I2859,I50742,I50802,);
not I_2818 (I50810,I216185);
or I_2819 (I50827,I216209,I216185);
nor I_2820 (I50844,I50802,I216209);
nand I_2821 (I50719,I50810,I50844);
nor I_2822 (I50875,I216200,I216209);
nand I_2823 (I50713,I50875,I50810);
not I_2824 (I50906,I216191);
nand I_2825 (I50923,I50810,I50906);
nor I_2826 (I50940,I216194,I216188);
not I_2827 (I50957,I50940);
nor I_2828 (I50974,I50957,I50923);
nor I_2829 (I50991,I50875,I50974);
DFFARX1 I_2830 (I50991,I2859,I50742,I50728,);
nor I_2831 (I50725,I50940,I50827);
DFFARX1 I_2832 (I50940,I2859,I50742,I50731,);
nor I_2833 (I51050,I50906,I216194);
nor I_2834 (I51067,I51050,I216185);
nor I_2835 (I51084,I216206,I216185);
DFFARX1 I_2836 (I51084,I2859,I50742,I51110,);
nor I_2837 (I50710,I51110,I51067);
DFFARX1 I_2838 (I51110,I2859,I50742,I51141,);
nand I_2839 (I51149,I51141,I216188);
nor I_2840 (I50734,I50776,I51149);
not I_2841 (I51180,I51110);
nand I_2842 (I51197,I51180,I216188);
nor I_2843 (I51214,I50776,I51197);
nor I_2844 (I50716,I50802,I51214);
nor I_2845 (I51245,I216206,I216200);
nor I_2846 (I51262,I50802,I51245);
DFFARX1 I_2847 (I51262,I2859,I50742,I50707,);
and I_2848 (I50722,I50875,I216206);
not I_2849 (I51337,I2866);
DFFARX1 I_2850 (I135121,I2859,I51337,I51363,);
not I_2851 (I51371,I51363);
DFFARX1 I_2852 (I135118,I2859,I51337,I51397,);
not I_2853 (I51405,I135115);
or I_2854 (I51422,I135127,I135115);
nor I_2855 (I51439,I51397,I135127);
nand I_2856 (I51314,I51405,I51439);
nor I_2857 (I51470,I135136,I135127);
nand I_2858 (I51308,I51470,I51405);
not I_2859 (I51501,I135133);
nand I_2860 (I51518,I51405,I51501);
nor I_2861 (I51535,I135112,I135112);
not I_2862 (I51552,I51535);
nor I_2863 (I51569,I51552,I51518);
nor I_2864 (I51586,I51470,I51569);
DFFARX1 I_2865 (I51586,I2859,I51337,I51323,);
nor I_2866 (I51320,I51535,I51422);
DFFARX1 I_2867 (I51535,I2859,I51337,I51326,);
nor I_2868 (I51645,I51501,I135112);
nor I_2869 (I51662,I51645,I135115);
nor I_2870 (I51679,I135124,I135139);
DFFARX1 I_2871 (I51679,I2859,I51337,I51705,);
nor I_2872 (I51305,I51705,I51662);
DFFARX1 I_2873 (I51705,I2859,I51337,I51736,);
nand I_2874 (I51744,I51736,I135130);
nor I_2875 (I51329,I51371,I51744);
not I_2876 (I51775,I51705);
nand I_2877 (I51792,I51775,I135130);
nor I_2878 (I51809,I51371,I51792);
nor I_2879 (I51311,I51397,I51809);
nor I_2880 (I51840,I135124,I135136);
nor I_2881 (I51857,I51397,I51840);
DFFARX1 I_2882 (I51857,I2859,I51337,I51302,);
and I_2883 (I51317,I51470,I135124);
not I_2884 (I51932,I2866);
DFFARX1 I_2885 (I377963,I2859,I51932,I51958,);
not I_2886 (I51966,I51958);
DFFARX1 I_2887 (I377984,I2859,I51932,I51992,);
not I_2888 (I52000,I377966);
or I_2889 (I52017,I377957,I377966);
nor I_2890 (I52034,I51992,I377957);
nand I_2891 (I51909,I52000,I52034);
nor I_2892 (I52065,I377969,I377957);
nand I_2893 (I51903,I52065,I52000);
not I_2894 (I52096,I377960);
nand I_2895 (I52113,I52000,I52096);
nor I_2896 (I52130,I377978,I377981);
not I_2897 (I52147,I52130);
nor I_2898 (I52164,I52147,I52113);
nor I_2899 (I52181,I52065,I52164);
DFFARX1 I_2900 (I52181,I2859,I51932,I51918,);
nor I_2901 (I51915,I52130,I52017);
DFFARX1 I_2902 (I52130,I2859,I51932,I51921,);
nor I_2903 (I52240,I52096,I377978);
nor I_2904 (I52257,I52240,I377966);
nor I_2905 (I52274,I377972,I377975);
DFFARX1 I_2906 (I52274,I2859,I51932,I52300,);
nor I_2907 (I51900,I52300,I52257);
DFFARX1 I_2908 (I52300,I2859,I51932,I52331,);
nand I_2909 (I52339,I52331,I377957);
nor I_2910 (I51924,I51966,I52339);
not I_2911 (I52370,I52300);
nand I_2912 (I52387,I52370,I377957);
nor I_2913 (I52404,I51966,I52387);
nor I_2914 (I51906,I51992,I52404);
nor I_2915 (I52435,I377972,I377969);
nor I_2916 (I52452,I51992,I52435);
DFFARX1 I_2917 (I52452,I2859,I51932,I51897,);
and I_2918 (I51912,I52065,I377972);
not I_2919 (I52527,I2866);
DFFARX1 I_2920 (I442373,I2859,I52527,I52553,);
not I_2921 (I52561,I52553);
DFFARX1 I_2922 (I442370,I2859,I52527,I52587,);
not I_2923 (I52595,I442379);
or I_2924 (I52612,I442370,I442379);
nor I_2925 (I52629,I52587,I442370);
nand I_2926 (I52504,I52595,I52629);
nor I_2927 (I52660,I442382,I442370);
nand I_2928 (I52498,I52660,I52595);
not I_2929 (I52691,I442376);
nand I_2930 (I52708,I52595,I52691);
nor I_2931 (I52725,I442373,I442391);
not I_2932 (I52742,I52725);
nor I_2933 (I52759,I52742,I52708);
nor I_2934 (I52776,I52660,I52759);
DFFARX1 I_2935 (I52776,I2859,I52527,I52513,);
nor I_2936 (I52510,I52725,I52612);
DFFARX1 I_2937 (I52725,I2859,I52527,I52516,);
nor I_2938 (I52835,I52691,I442373);
nor I_2939 (I52852,I52835,I442379);
nor I_2940 (I52869,I442394,I442388);
DFFARX1 I_2941 (I52869,I2859,I52527,I52895,);
nor I_2942 (I52495,I52895,I52852);
DFFARX1 I_2943 (I52895,I2859,I52527,I52926,);
nand I_2944 (I52934,I52926,I442385);
nor I_2945 (I52519,I52561,I52934);
not I_2946 (I52965,I52895);
nand I_2947 (I52982,I52965,I442385);
nor I_2948 (I52999,I52561,I52982);
nor I_2949 (I52501,I52587,I52999);
nor I_2950 (I53030,I442394,I442382);
nor I_2951 (I53047,I52587,I53030);
DFFARX1 I_2952 (I53047,I2859,I52527,I52492,);
and I_2953 (I52507,I52660,I442394);
not I_2954 (I53122,I2866);
DFFARX1 I_2955 (I40120,I2859,I53122,I53148,);
not I_2956 (I53156,I53148);
DFFARX1 I_2957 (I40114,I2859,I53122,I53182,);
not I_2958 (I53190,I40123);
or I_2959 (I53207,I40108,I40123);
nor I_2960 (I53224,I53182,I40108);
nand I_2961 (I53099,I53190,I53224);
nor I_2962 (I53255,I40099,I40108);
nand I_2963 (I53093,I53255,I53190);
not I_2964 (I53286,I40099);
nand I_2965 (I53303,I53190,I53286);
nor I_2966 (I53320,I40102,I40117);
not I_2967 (I53337,I53320);
nor I_2968 (I53354,I53337,I53303);
nor I_2969 (I53371,I53255,I53354);
DFFARX1 I_2970 (I53371,I2859,I53122,I53108,);
nor I_2971 (I53105,I53320,I53207);
DFFARX1 I_2972 (I53320,I2859,I53122,I53111,);
nor I_2973 (I53430,I53286,I40102);
nor I_2974 (I53447,I53430,I40123);
nor I_2975 (I53464,I40102,I40111);
DFFARX1 I_2976 (I53464,I2859,I53122,I53490,);
nor I_2977 (I53090,I53490,I53447);
DFFARX1 I_2978 (I53490,I2859,I53122,I53521,);
nand I_2979 (I53529,I53521,I40105);
nor I_2980 (I53114,I53156,I53529);
not I_2981 (I53560,I53490);
nand I_2982 (I53577,I53560,I40105);
nor I_2983 (I53594,I53156,I53577);
nor I_2984 (I53096,I53182,I53594);
nor I_2985 (I53625,I40102,I40099);
nor I_2986 (I53642,I53182,I53625);
DFFARX1 I_2987 (I53642,I2859,I53122,I53087,);
and I_2988 (I53102,I53255,I40102);
not I_2989 (I53717,I2866);
DFFARX1 I_2990 (I499595,I2859,I53717,I53743,);
not I_2991 (I53751,I53743);
DFFARX1 I_2992 (I499592,I2859,I53717,I53777,);
not I_2993 (I53785,I499601);
or I_2994 (I53802,I499592,I499601);
nor I_2995 (I53819,I53777,I499592);
nand I_2996 (I53694,I53785,I53819);
nor I_2997 (I53850,I499604,I499592);
nand I_2998 (I53688,I53850,I53785);
not I_2999 (I53881,I499598);
nand I_3000 (I53898,I53785,I53881);
nor I_3001 (I53915,I499595,I499613);
not I_3002 (I53932,I53915);
nor I_3003 (I53949,I53932,I53898);
nor I_3004 (I53966,I53850,I53949);
DFFARX1 I_3005 (I53966,I2859,I53717,I53703,);
nor I_3006 (I53700,I53915,I53802);
DFFARX1 I_3007 (I53915,I2859,I53717,I53706,);
nor I_3008 (I54025,I53881,I499595);
nor I_3009 (I54042,I54025,I499601);
nor I_3010 (I54059,I499616,I499610);
DFFARX1 I_3011 (I54059,I2859,I53717,I54085,);
nor I_3012 (I53685,I54085,I54042);
DFFARX1 I_3013 (I54085,I2859,I53717,I54116,);
nand I_3014 (I54124,I54116,I499607);
nor I_3015 (I53709,I53751,I54124);
not I_3016 (I54155,I54085);
nand I_3017 (I54172,I54155,I499607);
nor I_3018 (I54189,I53751,I54172);
nor I_3019 (I53691,I53777,I54189);
nor I_3020 (I54220,I499616,I499604);
nor I_3021 (I54237,I53777,I54220);
DFFARX1 I_3022 (I54237,I2859,I53717,I53682,);
and I_3023 (I53697,I53850,I499616);
not I_3024 (I54309,I2866);
DFFARX1 I_3025 (I320707,I2859,I54309,I54335,);
DFFARX1 I_3026 (I54335,I2859,I54309,I54352,);
not I_3027 (I54301,I54352);
not I_3028 (I54374,I54335);
DFFARX1 I_3029 (I320701,I2859,I54309,I54400,);
not I_3030 (I54408,I54400);
and I_3031 (I54425,I54374,I320719);
not I_3032 (I54442,I320707);
nand I_3033 (I54459,I54442,I320719);
not I_3034 (I54476,I320701);
nor I_3035 (I54493,I54476,I320713);
nand I_3036 (I54510,I54493,I320704);
nor I_3037 (I54527,I54510,I54459);
DFFARX1 I_3038 (I54527,I2859,I54309,I54277,);
not I_3039 (I54558,I54510);
not I_3040 (I54575,I320713);
nand I_3041 (I54592,I54575,I320719);
nor I_3042 (I54609,I320713,I320707);
nand I_3043 (I54289,I54425,I54609);
nand I_3044 (I54283,I54374,I320713);
nand I_3045 (I54654,I54476,I320716);
DFFARX1 I_3046 (I54654,I2859,I54309,I54298,);
DFFARX1 I_3047 (I54654,I2859,I54309,I54292,);
not I_3048 (I54699,I320716);
nor I_3049 (I54716,I54699,I320722);
and I_3050 (I54733,I54716,I320704);
or I_3051 (I54750,I54733,I320710);
DFFARX1 I_3052 (I54750,I2859,I54309,I54776,);
nand I_3053 (I54784,I54776,I54442);
nor I_3054 (I54286,I54784,I54592);
nor I_3055 (I54280,I54776,I54408);
DFFARX1 I_3056 (I54776,I2859,I54309,I54838,);
not I_3057 (I54846,I54838);
nor I_3058 (I54295,I54846,I54558);
not I_3059 (I54904,I2866);
DFFARX1 I_3060 (I384432,I2859,I54904,I54930,);
DFFARX1 I_3061 (I54930,I2859,I54904,I54947,);
not I_3062 (I54896,I54947);
not I_3063 (I54969,I54930);
DFFARX1 I_3064 (I384441,I2859,I54904,I54995,);
not I_3065 (I55003,I54995);
and I_3066 (I55020,I54969,I384429);
not I_3067 (I55037,I384420);
nand I_3068 (I55054,I55037,I384429);
not I_3069 (I55071,I384426);
nor I_3070 (I55088,I55071,I384444);
nand I_3071 (I55105,I55088,I384417);
nor I_3072 (I55122,I55105,I55054);
DFFARX1 I_3073 (I55122,I2859,I54904,I54872,);
not I_3074 (I55153,I55105);
not I_3075 (I55170,I384444);
nand I_3076 (I55187,I55170,I384429);
nor I_3077 (I55204,I384444,I384420);
nand I_3078 (I54884,I55020,I55204);
nand I_3079 (I54878,I54969,I384444);
nand I_3080 (I55249,I55071,I384423);
DFFARX1 I_3081 (I55249,I2859,I54904,I54893,);
DFFARX1 I_3082 (I55249,I2859,I54904,I54887,);
not I_3083 (I55294,I384423);
nor I_3084 (I55311,I55294,I384435);
and I_3085 (I55328,I55311,I384417);
or I_3086 (I55345,I55328,I384438);
DFFARX1 I_3087 (I55345,I2859,I54904,I55371,);
nand I_3088 (I55379,I55371,I55037);
nor I_3089 (I54881,I55379,I55187);
nor I_3090 (I54875,I55371,I55003);
DFFARX1 I_3091 (I55371,I2859,I54904,I55433,);
not I_3092 (I55441,I55433);
nor I_3093 (I54890,I55441,I55153);
not I_3094 (I55499,I2866);
DFFARX1 I_3095 (I492656,I2859,I55499,I55525,);
DFFARX1 I_3096 (I55525,I2859,I55499,I55542,);
not I_3097 (I55491,I55542);
not I_3098 (I55564,I55525);
DFFARX1 I_3099 (I492656,I2859,I55499,I55590,);
not I_3100 (I55598,I55590);
and I_3101 (I55615,I55564,I492659);
not I_3102 (I55632,I492671);
nand I_3103 (I55649,I55632,I492659);
not I_3104 (I55666,I492677);
nor I_3105 (I55683,I55666,I492668);
nand I_3106 (I55700,I55683,I492674);
nor I_3107 (I55717,I55700,I55649);
DFFARX1 I_3108 (I55717,I2859,I55499,I55467,);
not I_3109 (I55748,I55700);
not I_3110 (I55765,I492668);
nand I_3111 (I55782,I55765,I492659);
nor I_3112 (I55799,I492668,I492671);
nand I_3113 (I55479,I55615,I55799);
nand I_3114 (I55473,I55564,I492668);
nand I_3115 (I55844,I55666,I492665);
DFFARX1 I_3116 (I55844,I2859,I55499,I55488,);
DFFARX1 I_3117 (I55844,I2859,I55499,I55482,);
not I_3118 (I55889,I492665);
nor I_3119 (I55906,I55889,I492662);
and I_3120 (I55923,I55906,I492680);
or I_3121 (I55940,I55923,I492659);
DFFARX1 I_3122 (I55940,I2859,I55499,I55966,);
nand I_3123 (I55974,I55966,I55632);
nor I_3124 (I55476,I55974,I55782);
nor I_3125 (I55470,I55966,I55598);
DFFARX1 I_3126 (I55966,I2859,I55499,I56028,);
not I_3127 (I56036,I56028);
nor I_3128 (I55485,I56036,I55748);
not I_3129 (I56094,I2866);
DFFARX1 I_3130 (I540396,I2859,I56094,I56120,);
DFFARX1 I_3131 (I56120,I2859,I56094,I56137,);
not I_3132 (I56086,I56137);
not I_3133 (I56159,I56120);
DFFARX1 I_3134 (I540387,I2859,I56094,I56185,);
not I_3135 (I56193,I56185);
and I_3136 (I56210,I56159,I540381);
not I_3137 (I56227,I540375);
nand I_3138 (I56244,I56227,I540381);
not I_3139 (I56261,I540402);
nor I_3140 (I56278,I56261,I540375);
nand I_3141 (I56295,I56278,I540399);
nor I_3142 (I56312,I56295,I56244);
DFFARX1 I_3143 (I56312,I2859,I56094,I56062,);
not I_3144 (I56343,I56295);
not I_3145 (I56360,I540375);
nand I_3146 (I56377,I56360,I540381);
nor I_3147 (I56394,I540375,I540375);
nand I_3148 (I56074,I56210,I56394);
nand I_3149 (I56068,I56159,I540375);
nand I_3150 (I56439,I56261,I540384);
DFFARX1 I_3151 (I56439,I2859,I56094,I56083,);
DFFARX1 I_3152 (I56439,I2859,I56094,I56077,);
not I_3153 (I56484,I540384);
nor I_3154 (I56501,I56484,I540390);
and I_3155 (I56518,I56501,I540393);
or I_3156 (I56535,I56518,I540378);
DFFARX1 I_3157 (I56535,I2859,I56094,I56561,);
nand I_3158 (I56569,I56561,I56227);
nor I_3159 (I56071,I56569,I56377);
nor I_3160 (I56065,I56561,I56193);
DFFARX1 I_3161 (I56561,I2859,I56094,I56623,);
not I_3162 (I56631,I56623);
nor I_3163 (I56080,I56631,I56343);
not I_3164 (I56689,I2866);
DFFARX1 I_3165 (I549321,I2859,I56689,I56715,);
DFFARX1 I_3166 (I56715,I2859,I56689,I56732,);
not I_3167 (I56681,I56732);
not I_3168 (I56754,I56715);
DFFARX1 I_3169 (I549312,I2859,I56689,I56780,);
not I_3170 (I56788,I56780);
and I_3171 (I56805,I56754,I549306);
not I_3172 (I56822,I549300);
nand I_3173 (I56839,I56822,I549306);
not I_3174 (I56856,I549327);
nor I_3175 (I56873,I56856,I549300);
nand I_3176 (I56890,I56873,I549324);
nor I_3177 (I56907,I56890,I56839);
DFFARX1 I_3178 (I56907,I2859,I56689,I56657,);
not I_3179 (I56938,I56890);
not I_3180 (I56955,I549300);
nand I_3181 (I56972,I56955,I549306);
nor I_3182 (I56989,I549300,I549300);
nand I_3183 (I56669,I56805,I56989);
nand I_3184 (I56663,I56754,I549300);
nand I_3185 (I57034,I56856,I549309);
DFFARX1 I_3186 (I57034,I2859,I56689,I56678,);
DFFARX1 I_3187 (I57034,I2859,I56689,I56672,);
not I_3188 (I57079,I549309);
nor I_3189 (I57096,I57079,I549315);
and I_3190 (I57113,I57096,I549318);
or I_3191 (I57130,I57113,I549303);
DFFARX1 I_3192 (I57130,I2859,I56689,I57156,);
nand I_3193 (I57164,I57156,I56822);
nor I_3194 (I56666,I57164,I56972);
nor I_3195 (I56660,I57156,I56788);
DFFARX1 I_3196 (I57156,I2859,I56689,I57218,);
not I_3197 (I57226,I57218);
nor I_3198 (I56675,I57226,I56938);
not I_3199 (I57284,I2866);
DFFARX1 I_3200 (I31149,I2859,I57284,I57310,);
DFFARX1 I_3201 (I57310,I2859,I57284,I57327,);
not I_3202 (I57276,I57327);
not I_3203 (I57349,I57310);
DFFARX1 I_3204 (I31143,I2859,I57284,I57375,);
not I_3205 (I57383,I57375);
and I_3206 (I57400,I57349,I31140);
not I_3207 (I57417,I31161);
nand I_3208 (I57434,I57417,I31140);
not I_3209 (I57451,I31155);
nor I_3210 (I57468,I57451,I31146);
nand I_3211 (I57485,I57468,I31152);
nor I_3212 (I57502,I57485,I57434);
DFFARX1 I_3213 (I57502,I2859,I57284,I57252,);
not I_3214 (I57533,I57485);
not I_3215 (I57550,I31146);
nand I_3216 (I57567,I57550,I31140);
nor I_3217 (I57584,I31146,I31161);
nand I_3218 (I57264,I57400,I57584);
nand I_3219 (I57258,I57349,I31146);
nand I_3220 (I57629,I57451,I31140);
DFFARX1 I_3221 (I57629,I2859,I57284,I57273,);
DFFARX1 I_3222 (I57629,I2859,I57284,I57267,);
not I_3223 (I57674,I31140);
nor I_3224 (I57691,I57674,I31158);
and I_3225 (I57708,I57691,I31164);
or I_3226 (I57725,I57708,I31143);
DFFARX1 I_3227 (I57725,I2859,I57284,I57751,);
nand I_3228 (I57759,I57751,I57417);
nor I_3229 (I57261,I57759,I57567);
nor I_3230 (I57255,I57751,I57383);
DFFARX1 I_3231 (I57751,I2859,I57284,I57813,);
not I_3232 (I57821,I57813);
nor I_3233 (I57270,I57821,I57533);
not I_3234 (I57879,I2866);
DFFARX1 I_3235 (I36946,I2859,I57879,I57905,);
DFFARX1 I_3236 (I57905,I2859,I57879,I57922,);
not I_3237 (I57871,I57922);
not I_3238 (I57944,I57905);
DFFARX1 I_3239 (I36940,I2859,I57879,I57970,);
not I_3240 (I57978,I57970);
and I_3241 (I57995,I57944,I36937);
not I_3242 (I58012,I36958);
nand I_3243 (I58029,I58012,I36937);
not I_3244 (I58046,I36952);
nor I_3245 (I58063,I58046,I36943);
nand I_3246 (I58080,I58063,I36949);
nor I_3247 (I58097,I58080,I58029);
DFFARX1 I_3248 (I58097,I2859,I57879,I57847,);
not I_3249 (I58128,I58080);
not I_3250 (I58145,I36943);
nand I_3251 (I58162,I58145,I36937);
nor I_3252 (I58179,I36943,I36958);
nand I_3253 (I57859,I57995,I58179);
nand I_3254 (I57853,I57944,I36943);
nand I_3255 (I58224,I58046,I36937);
DFFARX1 I_3256 (I58224,I2859,I57879,I57868,);
DFFARX1 I_3257 (I58224,I2859,I57879,I57862,);
not I_3258 (I58269,I36937);
nor I_3259 (I58286,I58269,I36955);
and I_3260 (I58303,I58286,I36961);
or I_3261 (I58320,I58303,I36940);
DFFARX1 I_3262 (I58320,I2859,I57879,I58346,);
nand I_3263 (I58354,I58346,I58012);
nor I_3264 (I57856,I58354,I58162);
nor I_3265 (I57850,I58346,I57978);
DFFARX1 I_3266 (I58346,I2859,I57879,I58408,);
not I_3267 (I58416,I58408);
nor I_3268 (I57865,I58416,I58128);
not I_3269 (I58474,I2866);
DFFARX1 I_3270 (I188720,I2859,I58474,I58500,);
DFFARX1 I_3271 (I58500,I2859,I58474,I58517,);
not I_3272 (I58466,I58517);
not I_3273 (I58539,I58500);
DFFARX1 I_3274 (I188708,I2859,I58474,I58565,);
not I_3275 (I58573,I58565);
and I_3276 (I58590,I58539,I188717);
not I_3277 (I58607,I188714);
nand I_3278 (I58624,I58607,I188717);
not I_3279 (I58641,I188705);
nor I_3280 (I58658,I58641,I188711);
nand I_3281 (I58675,I58658,I188696);
nor I_3282 (I58692,I58675,I58624);
DFFARX1 I_3283 (I58692,I2859,I58474,I58442,);
not I_3284 (I58723,I58675);
not I_3285 (I58740,I188711);
nand I_3286 (I58757,I58740,I188717);
nor I_3287 (I58774,I188711,I188714);
nand I_3288 (I58454,I58590,I58774);
nand I_3289 (I58448,I58539,I188711);
nand I_3290 (I58819,I58641,I188696);
DFFARX1 I_3291 (I58819,I2859,I58474,I58463,);
DFFARX1 I_3292 (I58819,I2859,I58474,I58457,);
not I_3293 (I58864,I188696);
nor I_3294 (I58881,I58864,I188702);
and I_3295 (I58898,I58881,I188699);
or I_3296 (I58915,I58898,I188723);
DFFARX1 I_3297 (I58915,I2859,I58474,I58941,);
nand I_3298 (I58949,I58941,I58607);
nor I_3299 (I58451,I58949,I58757);
nor I_3300 (I58445,I58941,I58573);
DFFARX1 I_3301 (I58941,I2859,I58474,I59003,);
not I_3302 (I59011,I59003);
nor I_3303 (I58460,I59011,I58723);
not I_3304 (I59069,I2866);
DFFARX1 I_3305 (I439480,I2859,I59069,I59095,);
DFFARX1 I_3306 (I59095,I2859,I59069,I59112,);
not I_3307 (I59061,I59112);
not I_3308 (I59134,I59095);
DFFARX1 I_3309 (I439480,I2859,I59069,I59160,);
not I_3310 (I59168,I59160);
and I_3311 (I59185,I59134,I439483);
not I_3312 (I59202,I439495);
nand I_3313 (I59219,I59202,I439483);
not I_3314 (I59236,I439501);
nor I_3315 (I59253,I59236,I439492);
nand I_3316 (I59270,I59253,I439498);
nor I_3317 (I59287,I59270,I59219);
DFFARX1 I_3318 (I59287,I2859,I59069,I59037,);
not I_3319 (I59318,I59270);
not I_3320 (I59335,I439492);
nand I_3321 (I59352,I59335,I439483);
nor I_3322 (I59369,I439492,I439495);
nand I_3323 (I59049,I59185,I59369);
nand I_3324 (I59043,I59134,I439492);
nand I_3325 (I59414,I59236,I439489);
DFFARX1 I_3326 (I59414,I2859,I59069,I59058,);
DFFARX1 I_3327 (I59414,I2859,I59069,I59052,);
not I_3328 (I59459,I439489);
nor I_3329 (I59476,I59459,I439486);
and I_3330 (I59493,I59476,I439504);
or I_3331 (I59510,I59493,I439483);
DFFARX1 I_3332 (I59510,I2859,I59069,I59536,);
nand I_3333 (I59544,I59536,I59202);
nor I_3334 (I59046,I59544,I59352);
nor I_3335 (I59040,I59536,I59168);
DFFARX1 I_3336 (I59536,I2859,I59069,I59598,);
not I_3337 (I59606,I59598);
nor I_3338 (I59055,I59606,I59318);
not I_3339 (I59664,I2866);
DFFARX1 I_3340 (I478206,I2859,I59664,I59690,);
DFFARX1 I_3341 (I59690,I2859,I59664,I59707,);
not I_3342 (I59656,I59707);
not I_3343 (I59729,I59690);
DFFARX1 I_3344 (I478206,I2859,I59664,I59755,);
not I_3345 (I59763,I59755);
and I_3346 (I59780,I59729,I478209);
not I_3347 (I59797,I478221);
nand I_3348 (I59814,I59797,I478209);
not I_3349 (I59831,I478227);
nor I_3350 (I59848,I59831,I478218);
nand I_3351 (I59865,I59848,I478224);
nor I_3352 (I59882,I59865,I59814);
DFFARX1 I_3353 (I59882,I2859,I59664,I59632,);
not I_3354 (I59913,I59865);
not I_3355 (I59930,I478218);
nand I_3356 (I59947,I59930,I478209);
nor I_3357 (I59964,I478218,I478221);
nand I_3358 (I59644,I59780,I59964);
nand I_3359 (I59638,I59729,I478218);
nand I_3360 (I60009,I59831,I478215);
DFFARX1 I_3361 (I60009,I2859,I59664,I59653,);
DFFARX1 I_3362 (I60009,I2859,I59664,I59647,);
not I_3363 (I60054,I478215);
nor I_3364 (I60071,I60054,I478212);
and I_3365 (I60088,I60071,I478230);
or I_3366 (I60105,I60088,I478209);
DFFARX1 I_3367 (I60105,I2859,I59664,I60131,);
nand I_3368 (I60139,I60131,I59797);
nor I_3369 (I59641,I60139,I59947);
nor I_3370 (I59635,I60131,I59763);
DFFARX1 I_3371 (I60131,I2859,I59664,I60193,);
not I_3372 (I60201,I60193);
nor I_3373 (I59650,I60201,I59913);
not I_3374 (I60259,I2866);
DFFARX1 I_3375 (I392184,I2859,I60259,I60285,);
DFFARX1 I_3376 (I60285,I2859,I60259,I60302,);
not I_3377 (I60251,I60302);
not I_3378 (I60324,I60285);
DFFARX1 I_3379 (I392193,I2859,I60259,I60350,);
not I_3380 (I60358,I60350);
and I_3381 (I60375,I60324,I392181);
not I_3382 (I60392,I392172);
nand I_3383 (I60409,I60392,I392181);
not I_3384 (I60426,I392178);
nor I_3385 (I60443,I60426,I392196);
nand I_3386 (I60460,I60443,I392169);
nor I_3387 (I60477,I60460,I60409);
DFFARX1 I_3388 (I60477,I2859,I60259,I60227,);
not I_3389 (I60508,I60460);
not I_3390 (I60525,I392196);
nand I_3391 (I60542,I60525,I392181);
nor I_3392 (I60559,I392196,I392172);
nand I_3393 (I60239,I60375,I60559);
nand I_3394 (I60233,I60324,I392196);
nand I_3395 (I60604,I60426,I392175);
DFFARX1 I_3396 (I60604,I2859,I60259,I60248,);
DFFARX1 I_3397 (I60604,I2859,I60259,I60242,);
not I_3398 (I60649,I392175);
nor I_3399 (I60666,I60649,I392187);
and I_3400 (I60683,I60666,I392169);
or I_3401 (I60700,I60683,I392190);
DFFARX1 I_3402 (I60700,I2859,I60259,I60726,);
nand I_3403 (I60734,I60726,I60392);
nor I_3404 (I60236,I60734,I60542);
nor I_3405 (I60230,I60726,I60358);
DFFARX1 I_3406 (I60726,I2859,I60259,I60788,);
not I_3407 (I60796,I60788);
nor I_3408 (I60245,I60796,I60508);
not I_3409 (I60854,I2866);
DFFARX1 I_3410 (I15354,I2859,I60854,I60880,);
DFFARX1 I_3411 (I60880,I2859,I60854,I60897,);
not I_3412 (I60846,I60897);
not I_3413 (I60919,I60880);
DFFARX1 I_3414 (I15330,I2859,I60854,I60945,);
not I_3415 (I60953,I60945);
and I_3416 (I60970,I60919,I15345);
not I_3417 (I60987,I15333);
nand I_3418 (I61004,I60987,I15345);
not I_3419 (I61021,I15336);
nor I_3420 (I61038,I61021,I15348);
nand I_3421 (I61055,I61038,I15339);
nor I_3422 (I61072,I61055,I61004);
DFFARX1 I_3423 (I61072,I2859,I60854,I60822,);
not I_3424 (I61103,I61055);
not I_3425 (I61120,I15348);
nand I_3426 (I61137,I61120,I15345);
nor I_3427 (I61154,I15348,I15333);
nand I_3428 (I60834,I60970,I61154);
nand I_3429 (I60828,I60919,I15348);
nand I_3430 (I61199,I61021,I15342);
DFFARX1 I_3431 (I61199,I2859,I60854,I60843,);
DFFARX1 I_3432 (I61199,I2859,I60854,I60837,);
not I_3433 (I61244,I15342);
nor I_3434 (I61261,I61244,I15333);
and I_3435 (I61278,I61261,I15330);
or I_3436 (I61295,I61278,I15351);
DFFARX1 I_3437 (I61295,I2859,I60854,I61321,);
nand I_3438 (I61329,I61321,I60987);
nor I_3439 (I60831,I61329,I61137);
nor I_3440 (I60825,I61321,I60953);
DFFARX1 I_3441 (I61321,I2859,I60854,I61383,);
not I_3442 (I61391,I61383);
nor I_3443 (I60840,I61391,I61103);
not I_3444 (I61449,I2866);
DFFARX1 I_3445 (I210842,I2859,I61449,I61475,);
DFFARX1 I_3446 (I61475,I2859,I61449,I61492,);
not I_3447 (I61441,I61492);
not I_3448 (I61514,I61475);
DFFARX1 I_3449 (I210836,I2859,I61449,I61540,);
not I_3450 (I61548,I61540);
and I_3451 (I61565,I61514,I210851);
not I_3452 (I61582,I210848);
nand I_3453 (I61599,I61582,I210851);
not I_3454 (I61616,I210839);
nor I_3455 (I61633,I61616,I210830);
nand I_3456 (I61650,I61633,I210833);
nor I_3457 (I61667,I61650,I61599);
DFFARX1 I_3458 (I61667,I2859,I61449,I61417,);
not I_3459 (I61698,I61650);
not I_3460 (I61715,I210830);
nand I_3461 (I61732,I61715,I210851);
nor I_3462 (I61749,I210830,I210848);
nand I_3463 (I61429,I61565,I61749);
nand I_3464 (I61423,I61514,I210830);
nand I_3465 (I61794,I61616,I210854);
DFFARX1 I_3466 (I61794,I2859,I61449,I61438,);
DFFARX1 I_3467 (I61794,I2859,I61449,I61432,);
not I_3468 (I61839,I210854);
nor I_3469 (I61856,I61839,I210845);
and I_3470 (I61873,I61856,I210830);
or I_3471 (I61890,I61873,I210833);
DFFARX1 I_3472 (I61890,I2859,I61449,I61916,);
nand I_3473 (I61924,I61916,I61582);
nor I_3474 (I61426,I61924,I61732);
nor I_3475 (I61420,I61916,I61548);
DFFARX1 I_3476 (I61916,I2859,I61449,I61978,);
not I_3477 (I61986,I61978);
nor I_3478 (I61435,I61986,I61698);
not I_3479 (I62044,I2866);
DFFARX1 I_3480 (I522375,I2859,I62044,I62070,);
DFFARX1 I_3481 (I62070,I2859,I62044,I62087,);
not I_3482 (I62036,I62087);
not I_3483 (I62109,I62070);
DFFARX1 I_3484 (I522387,I2859,I62044,I62135,);
not I_3485 (I62143,I62135);
and I_3486 (I62160,I62109,I522381);
not I_3487 (I62177,I522393);
nand I_3488 (I62194,I62177,I522381);
not I_3489 (I62211,I522378);
nor I_3490 (I62228,I62211,I522390);
nand I_3491 (I62245,I62228,I522372);
nor I_3492 (I62262,I62245,I62194);
DFFARX1 I_3493 (I62262,I2859,I62044,I62012,);
not I_3494 (I62293,I62245);
not I_3495 (I62310,I522390);
nand I_3496 (I62327,I62310,I522381);
nor I_3497 (I62344,I522390,I522393);
nand I_3498 (I62024,I62160,I62344);
nand I_3499 (I62018,I62109,I522390);
nand I_3500 (I62389,I62211,I522384);
DFFARX1 I_3501 (I62389,I2859,I62044,I62033,);
DFFARX1 I_3502 (I62389,I2859,I62044,I62027,);
not I_3503 (I62434,I522384);
nor I_3504 (I62451,I62434,I522375);
and I_3505 (I62468,I62451,I522372);
or I_3506 (I62485,I62468,I522396);
DFFARX1 I_3507 (I62485,I2859,I62044,I62511,);
nand I_3508 (I62519,I62511,I62177);
nor I_3509 (I62021,I62519,I62327);
nor I_3510 (I62015,I62511,I62143);
DFFARX1 I_3511 (I62511,I2859,I62044,I62573,);
not I_3512 (I62581,I62573);
nor I_3513 (I62030,I62581,I62293);
not I_3514 (I62639,I2866);
DFFARX1 I_3515 (I168048,I2859,I62639,I62665,);
DFFARX1 I_3516 (I62665,I2859,I62639,I62682,);
not I_3517 (I62631,I62682);
not I_3518 (I62704,I62665);
DFFARX1 I_3519 (I168036,I2859,I62639,I62730,);
not I_3520 (I62738,I62730);
and I_3521 (I62755,I62704,I168045);
not I_3522 (I62772,I168042);
nand I_3523 (I62789,I62772,I168045);
not I_3524 (I62806,I168033);
nor I_3525 (I62823,I62806,I168039);
nand I_3526 (I62840,I62823,I168024);
nor I_3527 (I62857,I62840,I62789);
DFFARX1 I_3528 (I62857,I2859,I62639,I62607,);
not I_3529 (I62888,I62840);
not I_3530 (I62905,I168039);
nand I_3531 (I62922,I62905,I168045);
nor I_3532 (I62939,I168039,I168042);
nand I_3533 (I62619,I62755,I62939);
nand I_3534 (I62613,I62704,I168039);
nand I_3535 (I62984,I62806,I168024);
DFFARX1 I_3536 (I62984,I2859,I62639,I62628,);
DFFARX1 I_3537 (I62984,I2859,I62639,I62622,);
not I_3538 (I63029,I168024);
nor I_3539 (I63046,I63029,I168030);
and I_3540 (I63063,I63046,I168027);
or I_3541 (I63080,I63063,I168051);
DFFARX1 I_3542 (I63080,I2859,I62639,I63106,);
nand I_3543 (I63114,I63106,I62772);
nor I_3544 (I62616,I63114,I62922);
nor I_3545 (I62610,I63106,I62738);
DFFARX1 I_3546 (I63106,I2859,I62639,I63168,);
not I_3547 (I63176,I63168);
nor I_3548 (I62625,I63176,I62888);
not I_3549 (I63234,I2866);
DFFARX1 I_3550 (I512292,I2859,I63234,I63260,);
DFFARX1 I_3551 (I63260,I2859,I63234,I63277,);
not I_3552 (I63226,I63277);
not I_3553 (I63299,I63260);
DFFARX1 I_3554 (I512277,I2859,I63234,I63325,);
not I_3555 (I63333,I63325);
and I_3556 (I63350,I63299,I512295);
not I_3557 (I63367,I512277);
nand I_3558 (I63384,I63367,I512295);
not I_3559 (I63401,I512298);
nor I_3560 (I63418,I63401,I512289);
nand I_3561 (I63435,I63418,I512286);
nor I_3562 (I63452,I63435,I63384);
DFFARX1 I_3563 (I63452,I2859,I63234,I63202,);
not I_3564 (I63483,I63435);
not I_3565 (I63500,I512289);
nand I_3566 (I63517,I63500,I512295);
nor I_3567 (I63534,I512289,I512277);
nand I_3568 (I63214,I63350,I63534);
nand I_3569 (I63208,I63299,I512289);
nand I_3570 (I63579,I63401,I512283);
DFFARX1 I_3571 (I63579,I2859,I63234,I63223,);
DFFARX1 I_3572 (I63579,I2859,I63234,I63217,);
not I_3573 (I63624,I512283);
nor I_3574 (I63641,I63624,I512274);
and I_3575 (I63658,I63641,I512280);
or I_3576 (I63675,I63658,I512274);
DFFARX1 I_3577 (I63675,I2859,I63234,I63701,);
nand I_3578 (I63709,I63701,I63367);
nor I_3579 (I63211,I63709,I63517);
nor I_3580 (I63205,I63701,I63333);
DFFARX1 I_3581 (I63701,I2859,I63234,I63763,);
not I_3582 (I63771,I63763);
nor I_3583 (I63220,I63771,I63483);
not I_3584 (I63829,I2866);
DFFARX1 I_3585 (I218577,I2859,I63829,I63855,);
DFFARX1 I_3586 (I63855,I2859,I63829,I63872,);
not I_3587 (I63821,I63872);
not I_3588 (I63894,I63855);
DFFARX1 I_3589 (I218571,I2859,I63829,I63920,);
not I_3590 (I63928,I63920);
and I_3591 (I63945,I63894,I218586);
not I_3592 (I63962,I218583);
nand I_3593 (I63979,I63962,I218586);
not I_3594 (I63996,I218574);
nor I_3595 (I64013,I63996,I218565);
nand I_3596 (I64030,I64013,I218568);
nor I_3597 (I64047,I64030,I63979);
DFFARX1 I_3598 (I64047,I2859,I63829,I63797,);
not I_3599 (I64078,I64030);
not I_3600 (I64095,I218565);
nand I_3601 (I64112,I64095,I218586);
nor I_3602 (I64129,I218565,I218583);
nand I_3603 (I63809,I63945,I64129);
nand I_3604 (I63803,I63894,I218565);
nand I_3605 (I64174,I63996,I218589);
DFFARX1 I_3606 (I64174,I2859,I63829,I63818,);
DFFARX1 I_3607 (I64174,I2859,I63829,I63812,);
not I_3608 (I64219,I218589);
nor I_3609 (I64236,I64219,I218580);
and I_3610 (I64253,I64236,I218565);
or I_3611 (I64270,I64253,I218568);
DFFARX1 I_3612 (I64270,I2859,I63829,I64296,);
nand I_3613 (I64304,I64296,I63962);
nor I_3614 (I63806,I64304,I64112);
nor I_3615 (I63800,I64296,I63928);
DFFARX1 I_3616 (I64296,I2859,I63829,I64358,);
not I_3617 (I64366,I64358);
nor I_3618 (I63815,I64366,I64078);
not I_3619 (I64424,I2866);
DFFARX1 I_3620 (I146706,I2859,I64424,I64450,);
DFFARX1 I_3621 (I64450,I2859,I64424,I64467,);
not I_3622 (I64416,I64467);
not I_3623 (I64489,I64450);
DFFARX1 I_3624 (I146721,I2859,I64424,I64515,);
not I_3625 (I64523,I64515);
and I_3626 (I64540,I64489,I146718);
not I_3627 (I64557,I146706);
nand I_3628 (I64574,I64557,I146718);
not I_3629 (I64591,I146715);
nor I_3630 (I64608,I64591,I146730);
nand I_3631 (I64625,I64608,I146727);
nor I_3632 (I64642,I64625,I64574);
DFFARX1 I_3633 (I64642,I2859,I64424,I64392,);
not I_3634 (I64673,I64625);
not I_3635 (I64690,I146730);
nand I_3636 (I64707,I64690,I146718);
nor I_3637 (I64724,I146730,I146706);
nand I_3638 (I64404,I64540,I64724);
nand I_3639 (I64398,I64489,I146730);
nand I_3640 (I64769,I64591,I146724);
DFFARX1 I_3641 (I64769,I2859,I64424,I64413,);
DFFARX1 I_3642 (I64769,I2859,I64424,I64407,);
not I_3643 (I64814,I146724);
nor I_3644 (I64831,I64814,I146712);
and I_3645 (I64848,I64831,I146733);
or I_3646 (I64865,I64848,I146709);
DFFARX1 I_3647 (I64865,I2859,I64424,I64891,);
nand I_3648 (I64899,I64891,I64557);
nor I_3649 (I64401,I64899,I64707);
nor I_3650 (I64395,I64891,I64523);
DFFARX1 I_3651 (I64891,I2859,I64424,I64953,);
not I_3652 (I64961,I64953);
nor I_3653 (I64410,I64961,I64673);
not I_3654 (I65019,I2866);
DFFARX1 I_3655 (I372804,I2859,I65019,I65045,);
DFFARX1 I_3656 (I65045,I2859,I65019,I65062,);
not I_3657 (I65011,I65062);
not I_3658 (I65084,I65045);
DFFARX1 I_3659 (I372813,I2859,I65019,I65110,);
not I_3660 (I65118,I65110);
and I_3661 (I65135,I65084,I372801);
not I_3662 (I65152,I372792);
nand I_3663 (I65169,I65152,I372801);
not I_3664 (I65186,I372798);
nor I_3665 (I65203,I65186,I372816);
nand I_3666 (I65220,I65203,I372789);
nor I_3667 (I65237,I65220,I65169);
DFFARX1 I_3668 (I65237,I2859,I65019,I64987,);
not I_3669 (I65268,I65220);
not I_3670 (I65285,I372816);
nand I_3671 (I65302,I65285,I372801);
nor I_3672 (I65319,I372816,I372792);
nand I_3673 (I64999,I65135,I65319);
nand I_3674 (I64993,I65084,I372816);
nand I_3675 (I65364,I65186,I372795);
DFFARX1 I_3676 (I65364,I2859,I65019,I65008,);
DFFARX1 I_3677 (I65364,I2859,I65019,I65002,);
not I_3678 (I65409,I372795);
nor I_3679 (I65426,I65409,I372807);
and I_3680 (I65443,I65426,I372789);
or I_3681 (I65460,I65443,I372810);
DFFARX1 I_3682 (I65460,I2859,I65019,I65486,);
nand I_3683 (I65494,I65486,I65152);
nor I_3684 (I64996,I65494,I65302);
nor I_3685 (I64990,I65486,I65118);
DFFARX1 I_3686 (I65486,I2859,I65019,I65548,);
not I_3687 (I65556,I65548);
nor I_3688 (I65005,I65556,I65268);
not I_3689 (I65614,I2866);
DFFARX1 I_3690 (I461444,I2859,I65614,I65640,);
DFFARX1 I_3691 (I65640,I2859,I65614,I65657,);
not I_3692 (I65606,I65657);
not I_3693 (I65679,I65640);
DFFARX1 I_3694 (I461444,I2859,I65614,I65705,);
not I_3695 (I65713,I65705);
and I_3696 (I65730,I65679,I461447);
not I_3697 (I65747,I461459);
nand I_3698 (I65764,I65747,I461447);
not I_3699 (I65781,I461465);
nor I_3700 (I65798,I65781,I461456);
nand I_3701 (I65815,I65798,I461462);
nor I_3702 (I65832,I65815,I65764);
DFFARX1 I_3703 (I65832,I2859,I65614,I65582,);
not I_3704 (I65863,I65815);
not I_3705 (I65880,I461456);
nand I_3706 (I65897,I65880,I461447);
nor I_3707 (I65914,I461456,I461459);
nand I_3708 (I65594,I65730,I65914);
nand I_3709 (I65588,I65679,I461456);
nand I_3710 (I65959,I65781,I461453);
DFFARX1 I_3711 (I65959,I2859,I65614,I65603,);
DFFARX1 I_3712 (I65959,I2859,I65614,I65597,);
not I_3713 (I66004,I461453);
nor I_3714 (I66021,I66004,I461450);
and I_3715 (I66038,I66021,I461468);
or I_3716 (I66055,I66038,I461447);
DFFARX1 I_3717 (I66055,I2859,I65614,I66081,);
nand I_3718 (I66089,I66081,I65747);
nor I_3719 (I65591,I66089,I65897);
nor I_3720 (I65585,I66081,I65713);
DFFARX1 I_3721 (I66081,I2859,I65614,I66143,);
not I_3722 (I66151,I66143);
nor I_3723 (I65600,I66151,I65863);
not I_3724 (I66209,I2866);
DFFARX1 I_3725 (I1556,I2859,I66209,I66235,);
DFFARX1 I_3726 (I66235,I2859,I66209,I66252,);
not I_3727 (I66201,I66252);
not I_3728 (I66274,I66235);
DFFARX1 I_3729 (I2668,I2859,I66209,I66300,);
not I_3730 (I66308,I66300);
and I_3731 (I66325,I66274,I2804);
not I_3732 (I66342,I1876);
nand I_3733 (I66359,I66342,I2804);
not I_3734 (I66376,I2284);
nor I_3735 (I66393,I66376,I2340);
nand I_3736 (I66410,I66393,I1476);
nor I_3737 (I66427,I66410,I66359);
DFFARX1 I_3738 (I66427,I2859,I66209,I66177,);
not I_3739 (I66458,I66410);
not I_3740 (I66475,I2340);
nand I_3741 (I66492,I66475,I2804);
nor I_3742 (I66509,I2340,I1876);
nand I_3743 (I66189,I66325,I66509);
nand I_3744 (I66183,I66274,I2340);
nand I_3745 (I66554,I66376,I2772);
DFFARX1 I_3746 (I66554,I2859,I66209,I66198,);
DFFARX1 I_3747 (I66554,I2859,I66209,I66192,);
not I_3748 (I66599,I2772);
nor I_3749 (I66616,I66599,I1508);
and I_3750 (I66633,I66616,I2812);
or I_3751 (I66650,I66633,I2708);
DFFARX1 I_3752 (I66650,I2859,I66209,I66676,);
nand I_3753 (I66684,I66676,I66342);
nor I_3754 (I66186,I66684,I66492);
nor I_3755 (I66180,I66676,I66308);
DFFARX1 I_3756 (I66676,I2859,I66209,I66738,);
not I_3757 (I66746,I66738);
nor I_3758 (I66195,I66746,I66458);
not I_3759 (I66804,I2866);
DFFARX1 I_3760 (I22190,I2859,I66804,I66830,);
DFFARX1 I_3761 (I66830,I2859,I66804,I66847,);
not I_3762 (I66796,I66847);
not I_3763 (I66869,I66830);
DFFARX1 I_3764 (I22184,I2859,I66804,I66895,);
not I_3765 (I66903,I66895);
and I_3766 (I66920,I66869,I22181);
not I_3767 (I66937,I22202);
nand I_3768 (I66954,I66937,I22181);
not I_3769 (I66971,I22196);
nor I_3770 (I66988,I66971,I22187);
nand I_3771 (I67005,I66988,I22193);
nor I_3772 (I67022,I67005,I66954);
DFFARX1 I_3773 (I67022,I2859,I66804,I66772,);
not I_3774 (I67053,I67005);
not I_3775 (I67070,I22187);
nand I_3776 (I67087,I67070,I22181);
nor I_3777 (I67104,I22187,I22202);
nand I_3778 (I66784,I66920,I67104);
nand I_3779 (I66778,I66869,I22187);
nand I_3780 (I67149,I66971,I22181);
DFFARX1 I_3781 (I67149,I2859,I66804,I66793,);
DFFARX1 I_3782 (I67149,I2859,I66804,I66787,);
not I_3783 (I67194,I22181);
nor I_3784 (I67211,I67194,I22199);
and I_3785 (I67228,I67211,I22205);
or I_3786 (I67245,I67228,I22184);
DFFARX1 I_3787 (I67245,I2859,I66804,I67271,);
nand I_3788 (I67279,I67271,I66937);
nor I_3789 (I66781,I67279,I67087);
nor I_3790 (I66775,I67271,I66903);
DFFARX1 I_3791 (I67271,I2859,I66804,I67333,);
not I_3792 (I67341,I67333);
nor I_3793 (I66790,I67341,I67053);
not I_3794 (I67399,I2866);
DFFARX1 I_3795 (I565981,I2859,I67399,I67425,);
DFFARX1 I_3796 (I67425,I2859,I67399,I67442,);
not I_3797 (I67391,I67442);
not I_3798 (I67464,I67425);
DFFARX1 I_3799 (I565972,I2859,I67399,I67490,);
not I_3800 (I67498,I67490);
and I_3801 (I67515,I67464,I565966);
not I_3802 (I67532,I565960);
nand I_3803 (I67549,I67532,I565966);
not I_3804 (I67566,I565987);
nor I_3805 (I67583,I67566,I565960);
nand I_3806 (I67600,I67583,I565984);
nor I_3807 (I67617,I67600,I67549);
DFFARX1 I_3808 (I67617,I2859,I67399,I67367,);
not I_3809 (I67648,I67600);
not I_3810 (I67665,I565960);
nand I_3811 (I67682,I67665,I565966);
nor I_3812 (I67699,I565960,I565960);
nand I_3813 (I67379,I67515,I67699);
nand I_3814 (I67373,I67464,I565960);
nand I_3815 (I67744,I67566,I565969);
DFFARX1 I_3816 (I67744,I2859,I67399,I67388,);
DFFARX1 I_3817 (I67744,I2859,I67399,I67382,);
not I_3818 (I67789,I565969);
nor I_3819 (I67806,I67789,I565975);
and I_3820 (I67823,I67806,I565978);
or I_3821 (I67840,I67823,I565963);
DFFARX1 I_3822 (I67840,I2859,I67399,I67866,);
nand I_3823 (I67874,I67866,I67532);
nor I_3824 (I67376,I67874,I67682);
nor I_3825 (I67370,I67866,I67498);
DFFARX1 I_3826 (I67866,I2859,I67399,I67928,);
not I_3827 (I67936,I67928);
nor I_3828 (I67385,I67936,I67648);
not I_3829 (I67994,I2866);
DFFARX1 I_3830 (I180560,I2859,I67994,I68020,);
DFFARX1 I_3831 (I68020,I2859,I67994,I68037,);
not I_3832 (I67986,I68037);
not I_3833 (I68059,I68020);
DFFARX1 I_3834 (I180548,I2859,I67994,I68085,);
not I_3835 (I68093,I68085);
and I_3836 (I68110,I68059,I180557);
not I_3837 (I68127,I180554);
nand I_3838 (I68144,I68127,I180557);
not I_3839 (I68161,I180545);
nor I_3840 (I68178,I68161,I180551);
nand I_3841 (I68195,I68178,I180536);
nor I_3842 (I68212,I68195,I68144);
DFFARX1 I_3843 (I68212,I2859,I67994,I67962,);
not I_3844 (I68243,I68195);
not I_3845 (I68260,I180551);
nand I_3846 (I68277,I68260,I180557);
nor I_3847 (I68294,I180551,I180554);
nand I_3848 (I67974,I68110,I68294);
nand I_3849 (I67968,I68059,I180551);
nand I_3850 (I68339,I68161,I180536);
DFFARX1 I_3851 (I68339,I2859,I67994,I67983,);
DFFARX1 I_3852 (I68339,I2859,I67994,I67977,);
not I_3853 (I68384,I180536);
nor I_3854 (I68401,I68384,I180542);
and I_3855 (I68418,I68401,I180539);
or I_3856 (I68435,I68418,I180563);
DFFARX1 I_3857 (I68435,I2859,I67994,I68461,);
nand I_3858 (I68469,I68461,I68127);
nor I_3859 (I67971,I68469,I68277);
nor I_3860 (I67965,I68461,I68093);
DFFARX1 I_3861 (I68461,I2859,I67994,I68523,);
not I_3862 (I68531,I68523);
nor I_3863 (I67980,I68531,I68243);
not I_3864 (I68589,I2866);
DFFARX1 I_3865 (I537421,I2859,I68589,I68615,);
DFFARX1 I_3866 (I68615,I2859,I68589,I68632,);
not I_3867 (I68581,I68632);
not I_3868 (I68654,I68615);
DFFARX1 I_3869 (I537412,I2859,I68589,I68680,);
not I_3870 (I68688,I68680);
and I_3871 (I68705,I68654,I537406);
not I_3872 (I68722,I537400);
nand I_3873 (I68739,I68722,I537406);
not I_3874 (I68756,I537427);
nor I_3875 (I68773,I68756,I537400);
nand I_3876 (I68790,I68773,I537424);
nor I_3877 (I68807,I68790,I68739);
DFFARX1 I_3878 (I68807,I2859,I68589,I68557,);
not I_3879 (I68838,I68790);
not I_3880 (I68855,I537400);
nand I_3881 (I68872,I68855,I537406);
nor I_3882 (I68889,I537400,I537400);
nand I_3883 (I68569,I68705,I68889);
nand I_3884 (I68563,I68654,I537400);
nand I_3885 (I68934,I68756,I537409);
DFFARX1 I_3886 (I68934,I2859,I68589,I68578,);
DFFARX1 I_3887 (I68934,I2859,I68589,I68572,);
not I_3888 (I68979,I537409);
nor I_3889 (I68996,I68979,I537415);
and I_3890 (I69013,I68996,I537418);
or I_3891 (I69030,I69013,I537403);
DFFARX1 I_3892 (I69030,I2859,I68589,I69056,);
nand I_3893 (I69064,I69056,I68722);
nor I_3894 (I68566,I69064,I68872);
nor I_3895 (I68560,I69056,I68688);
DFFARX1 I_3896 (I69056,I2859,I68589,I69118,);
not I_3897 (I69126,I69118);
nor I_3898 (I68575,I69126,I68838);
not I_3899 (I69184,I2866);
DFFARX1 I_3900 (I429929,I2859,I69184,I69210,);
DFFARX1 I_3901 (I69210,I2859,I69184,I69227,);
not I_3902 (I69176,I69227);
not I_3903 (I69249,I69210);
DFFARX1 I_3904 (I429938,I2859,I69184,I69275,);
not I_3905 (I69283,I69275);
and I_3906 (I69300,I69249,I429932);
not I_3907 (I69317,I429926);
nand I_3908 (I69334,I69317,I429932);
not I_3909 (I69351,I429941);
nor I_3910 (I69368,I69351,I429929);
nand I_3911 (I69385,I69368,I429935);
nor I_3912 (I69402,I69385,I69334);
DFFARX1 I_3913 (I69402,I2859,I69184,I69152,);
not I_3914 (I69433,I69385);
not I_3915 (I69450,I429929);
nand I_3916 (I69467,I69450,I429932);
nor I_3917 (I69484,I429929,I429926);
nand I_3918 (I69164,I69300,I69484);
nand I_3919 (I69158,I69249,I429929);
nand I_3920 (I69529,I69351,I429932);
DFFARX1 I_3921 (I69529,I2859,I69184,I69173,);
DFFARX1 I_3922 (I69529,I2859,I69184,I69167,);
not I_3923 (I69574,I429932);
nor I_3924 (I69591,I69574,I429947);
and I_3925 (I69608,I69591,I429944);
or I_3926 (I69625,I69608,I429926);
DFFARX1 I_3927 (I69625,I2859,I69184,I69651,);
nand I_3928 (I69659,I69651,I69317);
nor I_3929 (I69161,I69659,I69467);
nor I_3930 (I69155,I69651,I69283);
DFFARX1 I_3931 (I69651,I2859,I69184,I69713,);
not I_3932 (I69721,I69713);
nor I_3933 (I69170,I69721,I69433);
not I_3934 (I69779,I2866);
DFFARX1 I_3935 (I153030,I2859,I69779,I69805,);
DFFARX1 I_3936 (I69805,I2859,I69779,I69822,);
not I_3937 (I69771,I69822);
not I_3938 (I69844,I69805);
DFFARX1 I_3939 (I153045,I2859,I69779,I69870,);
not I_3940 (I69878,I69870);
and I_3941 (I69895,I69844,I153042);
not I_3942 (I69912,I153030);
nand I_3943 (I69929,I69912,I153042);
not I_3944 (I69946,I153039);
nor I_3945 (I69963,I69946,I153054);
nand I_3946 (I69980,I69963,I153051);
nor I_3947 (I69997,I69980,I69929);
DFFARX1 I_3948 (I69997,I2859,I69779,I69747,);
not I_3949 (I70028,I69980);
not I_3950 (I70045,I153054);
nand I_3951 (I70062,I70045,I153042);
nor I_3952 (I70079,I153054,I153030);
nand I_3953 (I69759,I69895,I70079);
nand I_3954 (I69753,I69844,I153054);
nand I_3955 (I70124,I69946,I153048);
DFFARX1 I_3956 (I70124,I2859,I69779,I69768,);
DFFARX1 I_3957 (I70124,I2859,I69779,I69762,);
not I_3958 (I70169,I153048);
nor I_3959 (I70186,I70169,I153036);
and I_3960 (I70203,I70186,I153057);
or I_3961 (I70220,I70203,I153033);
DFFARX1 I_3962 (I70220,I2859,I69779,I70246,);
nand I_3963 (I70254,I70246,I69912);
nor I_3964 (I69756,I70254,I70062);
nor I_3965 (I69750,I70246,I69878);
DFFARX1 I_3966 (I70246,I2859,I69779,I70308,);
not I_3967 (I70316,I70308);
nor I_3968 (I69765,I70316,I70028);
not I_3969 (I70374,I2866);
DFFARX1 I_3970 (I373450,I2859,I70374,I70400,);
DFFARX1 I_3971 (I70400,I2859,I70374,I70417,);
not I_3972 (I70366,I70417);
not I_3973 (I70439,I70400);
DFFARX1 I_3974 (I373459,I2859,I70374,I70465,);
not I_3975 (I70473,I70465);
and I_3976 (I70490,I70439,I373447);
not I_3977 (I70507,I373438);
nand I_3978 (I70524,I70507,I373447);
not I_3979 (I70541,I373444);
nor I_3980 (I70558,I70541,I373462);
nand I_3981 (I70575,I70558,I373435);
nor I_3982 (I70592,I70575,I70524);
DFFARX1 I_3983 (I70592,I2859,I70374,I70342,);
not I_3984 (I70623,I70575);
not I_3985 (I70640,I373462);
nand I_3986 (I70657,I70640,I373447);
nor I_3987 (I70674,I373462,I373438);
nand I_3988 (I70354,I70490,I70674);
nand I_3989 (I70348,I70439,I373462);
nand I_3990 (I70719,I70541,I373441);
DFFARX1 I_3991 (I70719,I2859,I70374,I70363,);
DFFARX1 I_3992 (I70719,I2859,I70374,I70357,);
not I_3993 (I70764,I373441);
nor I_3994 (I70781,I70764,I373453);
and I_3995 (I70798,I70781,I373435);
or I_3996 (I70815,I70798,I373456);
DFFARX1 I_3997 (I70815,I2859,I70374,I70841,);
nand I_3998 (I70849,I70841,I70507);
nor I_3999 (I70351,I70849,I70657);
nor I_4000 (I70345,I70841,I70473);
DFFARX1 I_4001 (I70841,I2859,I70374,I70903,);
not I_4002 (I70911,I70903);
nor I_4003 (I70360,I70911,I70623);
not I_4004 (I70969,I2866);
DFFARX1 I_4005 (I40635,I2859,I70969,I70995,);
DFFARX1 I_4006 (I70995,I2859,I70969,I71012,);
not I_4007 (I70961,I71012);
not I_4008 (I71034,I70995);
DFFARX1 I_4009 (I40629,I2859,I70969,I71060,);
not I_4010 (I71068,I71060);
and I_4011 (I71085,I71034,I40626);
not I_4012 (I71102,I40647);
nand I_4013 (I71119,I71102,I40626);
not I_4014 (I71136,I40641);
nor I_4015 (I71153,I71136,I40632);
nand I_4016 (I71170,I71153,I40638);
nor I_4017 (I71187,I71170,I71119);
DFFARX1 I_4018 (I71187,I2859,I70969,I70937,);
not I_4019 (I71218,I71170);
not I_4020 (I71235,I40632);
nand I_4021 (I71252,I71235,I40626);
nor I_4022 (I71269,I40632,I40647);
nand I_4023 (I70949,I71085,I71269);
nand I_4024 (I70943,I71034,I40632);
nand I_4025 (I71314,I71136,I40626);
DFFARX1 I_4026 (I71314,I2859,I70969,I70958,);
DFFARX1 I_4027 (I71314,I2859,I70969,I70952,);
not I_4028 (I71359,I40626);
nor I_4029 (I71376,I71359,I40644);
and I_4030 (I71393,I71376,I40650);
or I_4031 (I71410,I71393,I40629);
DFFARX1 I_4032 (I71410,I2859,I70969,I71436,);
nand I_4033 (I71444,I71436,I71102);
nor I_4034 (I70946,I71444,I71252);
nor I_4035 (I70940,I71436,I71068);
DFFARX1 I_4036 (I71436,I2859,I70969,I71498,);
not I_4037 (I71506,I71498);
nor I_4038 (I70955,I71506,I71218);
not I_4039 (I71564,I2866);
DFFARX1 I_4040 (I1460,I2859,I71564,I71590,);
DFFARX1 I_4041 (I71590,I2859,I71564,I71607,);
not I_4042 (I71556,I71607);
not I_4043 (I71629,I71590);
DFFARX1 I_4044 (I2108,I2859,I71564,I71655,);
not I_4045 (I71663,I71655);
and I_4046 (I71680,I71629,I1396);
not I_4047 (I71697,I2652);
nand I_4048 (I71714,I71697,I1396);
not I_4049 (I71731,I2324);
nor I_4050 (I71748,I71731,I2780);
nand I_4051 (I71765,I71748,I1940);
nor I_4052 (I71782,I71765,I71714);
DFFARX1 I_4053 (I71782,I2859,I71564,I71532,);
not I_4054 (I71813,I71765);
not I_4055 (I71830,I2780);
nand I_4056 (I71847,I71830,I1396);
nor I_4057 (I71864,I2780,I2652);
nand I_4058 (I71544,I71680,I71864);
nand I_4059 (I71538,I71629,I2780);
nand I_4060 (I71909,I71731,I2836);
DFFARX1 I_4061 (I71909,I2859,I71564,I71553,);
DFFARX1 I_4062 (I71909,I2859,I71564,I71547,);
not I_4063 (I71954,I2836);
nor I_4064 (I71971,I71954,I2572);
and I_4065 (I71988,I71971,I1964);
or I_4066 (I72005,I71988,I2700);
DFFARX1 I_4067 (I72005,I2859,I71564,I72031,);
nand I_4068 (I72039,I72031,I71697);
nor I_4069 (I71541,I72039,I71847);
nor I_4070 (I71535,I72031,I71663);
DFFARX1 I_4071 (I72031,I2859,I71564,I72093,);
not I_4072 (I72101,I72093);
nor I_4073 (I71550,I72101,I71813);
not I_4074 (I72159,I2866);
DFFARX1 I_4075 (I500170,I2859,I72159,I72185,);
DFFARX1 I_4076 (I72185,I2859,I72159,I72202,);
not I_4077 (I72151,I72202);
not I_4078 (I72224,I72185);
DFFARX1 I_4079 (I500170,I2859,I72159,I72250,);
not I_4080 (I72258,I72250);
and I_4081 (I72275,I72224,I500173);
not I_4082 (I72292,I500185);
nand I_4083 (I72309,I72292,I500173);
not I_4084 (I72326,I500191);
nor I_4085 (I72343,I72326,I500182);
nand I_4086 (I72360,I72343,I500188);
nor I_4087 (I72377,I72360,I72309);
DFFARX1 I_4088 (I72377,I2859,I72159,I72127,);
not I_4089 (I72408,I72360);
not I_4090 (I72425,I500182);
nand I_4091 (I72442,I72425,I500173);
nor I_4092 (I72459,I500182,I500185);
nand I_4093 (I72139,I72275,I72459);
nand I_4094 (I72133,I72224,I500182);
nand I_4095 (I72504,I72326,I500179);
DFFARX1 I_4096 (I72504,I2859,I72159,I72148,);
DFFARX1 I_4097 (I72504,I2859,I72159,I72142,);
not I_4098 (I72549,I500179);
nor I_4099 (I72566,I72549,I500176);
and I_4100 (I72583,I72566,I500194);
or I_4101 (I72600,I72583,I500173);
DFFARX1 I_4102 (I72600,I2859,I72159,I72626,);
nand I_4103 (I72634,I72626,I72292);
nor I_4104 (I72136,I72634,I72442);
nor I_4105 (I72130,I72626,I72258);
DFFARX1 I_4106 (I72626,I2859,I72159,I72688,);
not I_4107 (I72696,I72688);
nor I_4108 (I72145,I72696,I72408);
not I_4109 (I72754,I2866);
DFFARX1 I_4110 (I383140,I2859,I72754,I72780,);
DFFARX1 I_4111 (I72780,I2859,I72754,I72797,);
not I_4112 (I72746,I72797);
not I_4113 (I72819,I72780);
DFFARX1 I_4114 (I383149,I2859,I72754,I72845,);
not I_4115 (I72853,I72845);
and I_4116 (I72870,I72819,I383137);
not I_4117 (I72887,I383128);
nand I_4118 (I72904,I72887,I383137);
not I_4119 (I72921,I383134);
nor I_4120 (I72938,I72921,I383152);
nand I_4121 (I72955,I72938,I383125);
nor I_4122 (I72972,I72955,I72904);
DFFARX1 I_4123 (I72972,I2859,I72754,I72722,);
not I_4124 (I73003,I72955);
not I_4125 (I73020,I383152);
nand I_4126 (I73037,I73020,I383137);
nor I_4127 (I73054,I383152,I383128);
nand I_4128 (I72734,I72870,I73054);
nand I_4129 (I72728,I72819,I383152);
nand I_4130 (I73099,I72921,I383131);
DFFARX1 I_4131 (I73099,I2859,I72754,I72743,);
DFFARX1 I_4132 (I73099,I2859,I72754,I72737,);
not I_4133 (I73144,I383131);
nor I_4134 (I73161,I73144,I383143);
and I_4135 (I73178,I73161,I383125);
or I_4136 (I73195,I73178,I383146);
DFFARX1 I_4137 (I73195,I2859,I72754,I73221,);
nand I_4138 (I73229,I73221,I72887);
nor I_4139 (I72731,I73229,I73037);
nor I_4140 (I72725,I73221,I72853);
DFFARX1 I_4141 (I73221,I2859,I72754,I73283,);
not I_4142 (I73291,I73283);
nor I_4143 (I72740,I73291,I73003);
not I_4144 (I73349,I2866);
DFFARX1 I_4145 (I567766,I2859,I73349,I73375,);
DFFARX1 I_4146 (I73375,I2859,I73349,I73392,);
not I_4147 (I73341,I73392);
not I_4148 (I73414,I73375);
DFFARX1 I_4149 (I567757,I2859,I73349,I73440,);
not I_4150 (I73448,I73440);
and I_4151 (I73465,I73414,I567751);
not I_4152 (I73482,I567745);
nand I_4153 (I73499,I73482,I567751);
not I_4154 (I73516,I567772);
nor I_4155 (I73533,I73516,I567745);
nand I_4156 (I73550,I73533,I567769);
nor I_4157 (I73567,I73550,I73499);
DFFARX1 I_4158 (I73567,I2859,I73349,I73317,);
not I_4159 (I73598,I73550);
not I_4160 (I73615,I567745);
nand I_4161 (I73632,I73615,I567751);
nor I_4162 (I73649,I567745,I567745);
nand I_4163 (I73329,I73465,I73649);
nand I_4164 (I73323,I73414,I567745);
nand I_4165 (I73694,I73516,I567754);
DFFARX1 I_4166 (I73694,I2859,I73349,I73338,);
DFFARX1 I_4167 (I73694,I2859,I73349,I73332,);
not I_4168 (I73739,I567754);
nor I_4169 (I73756,I73739,I567760);
and I_4170 (I73773,I73756,I567763);
or I_4171 (I73790,I73773,I567748);
DFFARX1 I_4172 (I73790,I2859,I73349,I73816,);
nand I_4173 (I73824,I73816,I73482);
nor I_4174 (I73326,I73824,I73632);
nor I_4175 (I73320,I73816,I73448);
DFFARX1 I_4176 (I73816,I2859,I73349,I73878,);
not I_4177 (I73886,I73878);
nor I_4178 (I73335,I73886,I73598);
not I_4179 (I73944,I2866);
DFFARX1 I_4180 (I444104,I2859,I73944,I73970,);
DFFARX1 I_4181 (I73970,I2859,I73944,I73987,);
not I_4182 (I73936,I73987);
not I_4183 (I74009,I73970);
DFFARX1 I_4184 (I444104,I2859,I73944,I74035,);
not I_4185 (I74043,I74035);
and I_4186 (I74060,I74009,I444107);
not I_4187 (I74077,I444119);
nand I_4188 (I74094,I74077,I444107);
not I_4189 (I74111,I444125);
nor I_4190 (I74128,I74111,I444116);
nand I_4191 (I74145,I74128,I444122);
nor I_4192 (I74162,I74145,I74094);
DFFARX1 I_4193 (I74162,I2859,I73944,I73912,);
not I_4194 (I74193,I74145);
not I_4195 (I74210,I444116);
nand I_4196 (I74227,I74210,I444107);
nor I_4197 (I74244,I444116,I444119);
nand I_4198 (I73924,I74060,I74244);
nand I_4199 (I73918,I74009,I444116);
nand I_4200 (I74289,I74111,I444113);
DFFARX1 I_4201 (I74289,I2859,I73944,I73933,);
DFFARX1 I_4202 (I74289,I2859,I73944,I73927,);
not I_4203 (I74334,I444113);
nor I_4204 (I74351,I74334,I444110);
and I_4205 (I74368,I74351,I444128);
or I_4206 (I74385,I74368,I444107);
DFFARX1 I_4207 (I74385,I2859,I73944,I74411,);
nand I_4208 (I74419,I74411,I74077);
nor I_4209 (I73921,I74419,I74227);
nor I_4210 (I73915,I74411,I74043);
DFFARX1 I_4211 (I74411,I2859,I73944,I74473,);
not I_4212 (I74481,I74473);
nor I_4213 (I73930,I74481,I74193);
not I_4214 (I74539,I2866);
DFFARX1 I_4215 (I155665,I2859,I74539,I74565,);
DFFARX1 I_4216 (I74565,I2859,I74539,I74582,);
not I_4217 (I74531,I74582);
not I_4218 (I74604,I74565);
DFFARX1 I_4219 (I155680,I2859,I74539,I74630,);
not I_4220 (I74638,I74630);
and I_4221 (I74655,I74604,I155677);
not I_4222 (I74672,I155665);
nand I_4223 (I74689,I74672,I155677);
not I_4224 (I74706,I155674);
nor I_4225 (I74723,I74706,I155689);
nand I_4226 (I74740,I74723,I155686);
nor I_4227 (I74757,I74740,I74689);
DFFARX1 I_4228 (I74757,I2859,I74539,I74507,);
not I_4229 (I74788,I74740);
not I_4230 (I74805,I155689);
nand I_4231 (I74822,I74805,I155677);
nor I_4232 (I74839,I155689,I155665);
nand I_4233 (I74519,I74655,I74839);
nand I_4234 (I74513,I74604,I155689);
nand I_4235 (I74884,I74706,I155683);
DFFARX1 I_4236 (I74884,I2859,I74539,I74528,);
DFFARX1 I_4237 (I74884,I2859,I74539,I74522,);
not I_4238 (I74929,I155683);
nor I_4239 (I74946,I74929,I155671);
and I_4240 (I74963,I74946,I155692);
or I_4241 (I74980,I74963,I155668);
DFFARX1 I_4242 (I74980,I2859,I74539,I75006,);
nand I_4243 (I75014,I75006,I74672);
nor I_4244 (I74516,I75014,I74822);
nor I_4245 (I74510,I75006,I74638);
DFFARX1 I_4246 (I75006,I2859,I74539,I75068,);
not I_4247 (I75076,I75068);
nor I_4248 (I74525,I75076,I74788);
not I_4249 (I75134,I2866);
DFFARX1 I_4250 (I211437,I2859,I75134,I75160,);
DFFARX1 I_4251 (I75160,I2859,I75134,I75177,);
not I_4252 (I75126,I75177);
not I_4253 (I75199,I75160);
DFFARX1 I_4254 (I211431,I2859,I75134,I75225,);
not I_4255 (I75233,I75225);
and I_4256 (I75250,I75199,I211446);
not I_4257 (I75267,I211443);
nand I_4258 (I75284,I75267,I211446);
not I_4259 (I75301,I211434);
nor I_4260 (I75318,I75301,I211425);
nand I_4261 (I75335,I75318,I211428);
nor I_4262 (I75352,I75335,I75284);
DFFARX1 I_4263 (I75352,I2859,I75134,I75102,);
not I_4264 (I75383,I75335);
not I_4265 (I75400,I211425);
nand I_4266 (I75417,I75400,I211446);
nor I_4267 (I75434,I211425,I211443);
nand I_4268 (I75114,I75250,I75434);
nand I_4269 (I75108,I75199,I211425);
nand I_4270 (I75479,I75301,I211449);
DFFARX1 I_4271 (I75479,I2859,I75134,I75123,);
DFFARX1 I_4272 (I75479,I2859,I75134,I75117,);
not I_4273 (I75524,I211449);
nor I_4274 (I75541,I75524,I211440);
and I_4275 (I75558,I75541,I211425);
or I_4276 (I75575,I75558,I211428);
DFFARX1 I_4277 (I75575,I2859,I75134,I75601,);
nand I_4278 (I75609,I75601,I75267);
nor I_4279 (I75111,I75609,I75417);
nor I_4280 (I75105,I75601,I75233);
DFFARX1 I_4281 (I75601,I2859,I75134,I75663,);
not I_4282 (I75671,I75663);
nor I_4283 (I75120,I75671,I75383);
not I_4284 (I75729,I2866);
DFFARX1 I_4285 (I231381,I2859,I75729,I75755,);
DFFARX1 I_4286 (I75755,I2859,I75729,I75772,);
not I_4287 (I75721,I75772);
not I_4288 (I75794,I75755);
DFFARX1 I_4289 (I231372,I2859,I75729,I75820,);
not I_4290 (I75828,I75820);
and I_4291 (I75845,I75794,I231390);
not I_4292 (I75862,I231387);
nand I_4293 (I75879,I75862,I231390);
not I_4294 (I75896,I231366);
nor I_4295 (I75913,I75896,I231369);
nand I_4296 (I75930,I75913,I231378);
nor I_4297 (I75947,I75930,I75879);
DFFARX1 I_4298 (I75947,I2859,I75729,I75697,);
not I_4299 (I75978,I75930);
not I_4300 (I75995,I231369);
nand I_4301 (I76012,I75995,I231390);
nor I_4302 (I76029,I231369,I231387);
nand I_4303 (I75709,I75845,I76029);
nand I_4304 (I75703,I75794,I231369);
nand I_4305 (I76074,I75896,I231384);
DFFARX1 I_4306 (I76074,I2859,I75729,I75718,);
DFFARX1 I_4307 (I76074,I2859,I75729,I75712,);
not I_4308 (I76119,I231384);
nor I_4309 (I76136,I76119,I231366);
and I_4310 (I76153,I76136,I231375);
or I_4311 (I76170,I76153,I231369);
DFFARX1 I_4312 (I76170,I2859,I75729,I76196,);
nand I_4313 (I76204,I76196,I75862);
nor I_4314 (I75706,I76204,I76012);
nor I_4315 (I75700,I76196,I75828);
DFFARX1 I_4316 (I76196,I2859,I75729,I76258,);
not I_4317 (I76266,I76258);
nor I_4318 (I75715,I76266,I75978);
not I_4319 (I76324,I2866);
DFFARX1 I_4320 (I202512,I2859,I76324,I76350,);
DFFARX1 I_4321 (I76350,I2859,I76324,I76367,);
not I_4322 (I76316,I76367);
not I_4323 (I76389,I76350);
DFFARX1 I_4324 (I202506,I2859,I76324,I76415,);
not I_4325 (I76423,I76415);
and I_4326 (I76440,I76389,I202521);
not I_4327 (I76457,I202518);
nand I_4328 (I76474,I76457,I202521);
not I_4329 (I76491,I202509);
nor I_4330 (I76508,I76491,I202500);
nand I_4331 (I76525,I76508,I202503);
nor I_4332 (I76542,I76525,I76474);
DFFARX1 I_4333 (I76542,I2859,I76324,I76292,);
not I_4334 (I76573,I76525);
not I_4335 (I76590,I202500);
nand I_4336 (I76607,I76590,I202521);
nor I_4337 (I76624,I202500,I202518);
nand I_4338 (I76304,I76440,I76624);
nand I_4339 (I76298,I76389,I202500);
nand I_4340 (I76669,I76491,I202524);
DFFARX1 I_4341 (I76669,I2859,I76324,I76313,);
DFFARX1 I_4342 (I76669,I2859,I76324,I76307,);
not I_4343 (I76714,I202524);
nor I_4344 (I76731,I76714,I202515);
and I_4345 (I76748,I76731,I202500);
or I_4346 (I76765,I76748,I202503);
DFFARX1 I_4347 (I76765,I2859,I76324,I76791,);
nand I_4348 (I76799,I76791,I76457);
nor I_4349 (I76301,I76799,I76607);
nor I_4350 (I76295,I76791,I76423);
DFFARX1 I_4351 (I76791,I2859,I76324,I76853,);
not I_4352 (I76861,I76853);
nor I_4353 (I76310,I76861,I76573);
not I_4354 (I76919,I2866);
DFFARX1 I_4355 (I181104,I2859,I76919,I76945,);
DFFARX1 I_4356 (I76945,I2859,I76919,I76962,);
not I_4357 (I76911,I76962);
not I_4358 (I76984,I76945);
DFFARX1 I_4359 (I181092,I2859,I76919,I77010,);
not I_4360 (I77018,I77010);
and I_4361 (I77035,I76984,I181101);
not I_4362 (I77052,I181098);
nand I_4363 (I77069,I77052,I181101);
not I_4364 (I77086,I181089);
nor I_4365 (I77103,I77086,I181095);
nand I_4366 (I77120,I77103,I181080);
nor I_4367 (I77137,I77120,I77069);
DFFARX1 I_4368 (I77137,I2859,I76919,I76887,);
not I_4369 (I77168,I77120);
not I_4370 (I77185,I181095);
nand I_4371 (I77202,I77185,I181101);
nor I_4372 (I77219,I181095,I181098);
nand I_4373 (I76899,I77035,I77219);
nand I_4374 (I76893,I76984,I181095);
nand I_4375 (I77264,I77086,I181080);
DFFARX1 I_4376 (I77264,I2859,I76919,I76908,);
DFFARX1 I_4377 (I77264,I2859,I76919,I76902,);
not I_4378 (I77309,I181080);
nor I_4379 (I77326,I77309,I181086);
and I_4380 (I77343,I77326,I181083);
or I_4381 (I77360,I77343,I181107);
DFFARX1 I_4382 (I77360,I2859,I76919,I77386,);
nand I_4383 (I77394,I77386,I77052);
nor I_4384 (I76896,I77394,I77202);
nor I_4385 (I76890,I77386,I77018);
DFFARX1 I_4386 (I77386,I2859,I76919,I77448,);
not I_4387 (I77456,I77448);
nor I_4388 (I76905,I77456,I77168);
not I_4389 (I77514,I2866);
DFFARX1 I_4390 (I502500,I2859,I77514,I77540,);
DFFARX1 I_4391 (I77540,I2859,I77514,I77557,);
not I_4392 (I77506,I77557);
not I_4393 (I77579,I77540);
DFFARX1 I_4394 (I502485,I2859,I77514,I77605,);
not I_4395 (I77613,I77605);
and I_4396 (I77630,I77579,I502503);
not I_4397 (I77647,I502485);
nand I_4398 (I77664,I77647,I502503);
not I_4399 (I77681,I502506);
nor I_4400 (I77698,I77681,I502497);
nand I_4401 (I77715,I77698,I502494);
nor I_4402 (I77732,I77715,I77664);
DFFARX1 I_4403 (I77732,I2859,I77514,I77482,);
not I_4404 (I77763,I77715);
not I_4405 (I77780,I502497);
nand I_4406 (I77797,I77780,I502503);
nor I_4407 (I77814,I502497,I502485);
nand I_4408 (I77494,I77630,I77814);
nand I_4409 (I77488,I77579,I502497);
nand I_4410 (I77859,I77681,I502491);
DFFARX1 I_4411 (I77859,I2859,I77514,I77503,);
DFFARX1 I_4412 (I77859,I2859,I77514,I77497,);
not I_4413 (I77904,I502491);
nor I_4414 (I77921,I77904,I502482);
and I_4415 (I77938,I77921,I502488);
or I_4416 (I77955,I77938,I502482);
DFFARX1 I_4417 (I77955,I2859,I77514,I77981,);
nand I_4418 (I77989,I77981,I77647);
nor I_4419 (I77491,I77989,I77797);
nor I_4420 (I77485,I77981,I77613);
DFFARX1 I_4421 (I77981,I2859,I77514,I78043,);
not I_4422 (I78051,I78043);
nor I_4423 (I77500,I78051,I77763);
not I_4424 (I78109,I2866);
DFFARX1 I_4425 (I37473,I2859,I78109,I78135,);
DFFARX1 I_4426 (I78135,I2859,I78109,I78152,);
not I_4427 (I78101,I78152);
not I_4428 (I78174,I78135);
DFFARX1 I_4429 (I37467,I2859,I78109,I78200,);
not I_4430 (I78208,I78200);
and I_4431 (I78225,I78174,I37464);
not I_4432 (I78242,I37485);
nand I_4433 (I78259,I78242,I37464);
not I_4434 (I78276,I37479);
nor I_4435 (I78293,I78276,I37470);
nand I_4436 (I78310,I78293,I37476);
nor I_4437 (I78327,I78310,I78259);
DFFARX1 I_4438 (I78327,I2859,I78109,I78077,);
not I_4439 (I78358,I78310);
not I_4440 (I78375,I37470);
nand I_4441 (I78392,I78375,I37464);
nor I_4442 (I78409,I37470,I37485);
nand I_4443 (I78089,I78225,I78409);
nand I_4444 (I78083,I78174,I37470);
nand I_4445 (I78454,I78276,I37464);
DFFARX1 I_4446 (I78454,I2859,I78109,I78098,);
DFFARX1 I_4447 (I78454,I2859,I78109,I78092,);
not I_4448 (I78499,I37464);
nor I_4449 (I78516,I78499,I37482);
and I_4450 (I78533,I78516,I37488);
or I_4451 (I78550,I78533,I37467);
DFFARX1 I_4452 (I78550,I2859,I78109,I78576,);
nand I_4453 (I78584,I78576,I78242);
nor I_4454 (I78086,I78584,I78392);
nor I_4455 (I78080,I78576,I78208);
DFFARX1 I_4456 (I78576,I2859,I78109,I78638,);
not I_4457 (I78646,I78638);
nor I_4458 (I78095,I78646,I78358);
not I_4459 (I78704,I2866);
DFFARX1 I_4460 (I127734,I2859,I78704,I78730,);
DFFARX1 I_4461 (I78730,I2859,I78704,I78747,);
not I_4462 (I78696,I78747);
not I_4463 (I78769,I78730);
DFFARX1 I_4464 (I127749,I2859,I78704,I78795,);
not I_4465 (I78803,I78795);
and I_4466 (I78820,I78769,I127746);
not I_4467 (I78837,I127734);
nand I_4468 (I78854,I78837,I127746);
not I_4469 (I78871,I127743);
nor I_4470 (I78888,I78871,I127758);
nand I_4471 (I78905,I78888,I127755);
nor I_4472 (I78922,I78905,I78854);
DFFARX1 I_4473 (I78922,I2859,I78704,I78672,);
not I_4474 (I78953,I78905);
not I_4475 (I78970,I127758);
nand I_4476 (I78987,I78970,I127746);
nor I_4477 (I79004,I127758,I127734);
nand I_4478 (I78684,I78820,I79004);
nand I_4479 (I78678,I78769,I127758);
nand I_4480 (I79049,I78871,I127752);
DFFARX1 I_4481 (I79049,I2859,I78704,I78693,);
DFFARX1 I_4482 (I79049,I2859,I78704,I78687,);
not I_4483 (I79094,I127752);
nor I_4484 (I79111,I79094,I127740);
and I_4485 (I79128,I79111,I127761);
or I_4486 (I79145,I79128,I127737);
DFFARX1 I_4487 (I79145,I2859,I78704,I79171,);
nand I_4488 (I79179,I79171,I78837);
nor I_4489 (I78681,I79179,I78987);
nor I_4490 (I78675,I79171,I78803);
DFFARX1 I_4491 (I79171,I2859,I78704,I79233,);
not I_4492 (I79241,I79233);
nor I_4493 (I78690,I79241,I78953);
not I_4494 (I79299,I2866);
DFFARX1 I_4495 (I369574,I2859,I79299,I79325,);
DFFARX1 I_4496 (I79325,I2859,I79299,I79342,);
not I_4497 (I79291,I79342);
not I_4498 (I79364,I79325);
DFFARX1 I_4499 (I369583,I2859,I79299,I79390,);
not I_4500 (I79398,I79390);
and I_4501 (I79415,I79364,I369571);
not I_4502 (I79432,I369562);
nand I_4503 (I79449,I79432,I369571);
not I_4504 (I79466,I369568);
nor I_4505 (I79483,I79466,I369586);
nand I_4506 (I79500,I79483,I369559);
nor I_4507 (I79517,I79500,I79449);
DFFARX1 I_4508 (I79517,I2859,I79299,I79267,);
not I_4509 (I79548,I79500);
not I_4510 (I79565,I369586);
nand I_4511 (I79582,I79565,I369571);
nor I_4512 (I79599,I369586,I369562);
nand I_4513 (I79279,I79415,I79599);
nand I_4514 (I79273,I79364,I369586);
nand I_4515 (I79644,I79466,I369565);
DFFARX1 I_4516 (I79644,I2859,I79299,I79288,);
DFFARX1 I_4517 (I79644,I2859,I79299,I79282,);
not I_4518 (I79689,I369565);
nor I_4519 (I79706,I79689,I369577);
and I_4520 (I79723,I79706,I369559);
or I_4521 (I79740,I79723,I369580);
DFFARX1 I_4522 (I79740,I2859,I79299,I79766,);
nand I_4523 (I79774,I79766,I79432);
nor I_4524 (I79276,I79774,I79582);
nor I_4525 (I79270,I79766,I79398);
DFFARX1 I_4526 (I79766,I2859,I79299,I79828,);
not I_4527 (I79836,I79828);
nor I_4528 (I79285,I79836,I79548);
not I_4529 (I79894,I2866);
DFFARX1 I_4530 (I358651,I2859,I79894,I79920,);
DFFARX1 I_4531 (I79920,I2859,I79894,I79937,);
not I_4532 (I79886,I79937);
not I_4533 (I79959,I79920);
DFFARX1 I_4534 (I358645,I2859,I79894,I79985,);
not I_4535 (I79993,I79985);
and I_4536 (I80010,I79959,I358663);
not I_4537 (I80027,I358651);
nand I_4538 (I80044,I80027,I358663);
not I_4539 (I80061,I358645);
nor I_4540 (I80078,I80061,I358657);
nand I_4541 (I80095,I80078,I358648);
nor I_4542 (I80112,I80095,I80044);
DFFARX1 I_4543 (I80112,I2859,I79894,I79862,);
not I_4544 (I80143,I80095);
not I_4545 (I80160,I358657);
nand I_4546 (I80177,I80160,I358663);
nor I_4547 (I80194,I358657,I358651);
nand I_4548 (I79874,I80010,I80194);
nand I_4549 (I79868,I79959,I358657);
nand I_4550 (I80239,I80061,I358660);
DFFARX1 I_4551 (I80239,I2859,I79894,I79883,);
DFFARX1 I_4552 (I80239,I2859,I79894,I79877,);
not I_4553 (I80284,I358660);
nor I_4554 (I80301,I80284,I358666);
and I_4555 (I80318,I80301,I358648);
or I_4556 (I80335,I80318,I358654);
DFFARX1 I_4557 (I80335,I2859,I79894,I80361,);
nand I_4558 (I80369,I80361,I80027);
nor I_4559 (I79871,I80369,I80177);
nor I_4560 (I79865,I80361,I79993);
DFFARX1 I_4561 (I80361,I2859,I79894,I80423,);
not I_4562 (I80431,I80423);
nor I_4563 (I79880,I80431,I80143);
not I_4564 (I80489,I2866);
DFFARX1 I_4565 (I219767,I2859,I80489,I80515,);
DFFARX1 I_4566 (I80515,I2859,I80489,I80532,);
not I_4567 (I80481,I80532);
not I_4568 (I80554,I80515);
DFFARX1 I_4569 (I219761,I2859,I80489,I80580,);
not I_4570 (I80588,I80580);
and I_4571 (I80605,I80554,I219776);
not I_4572 (I80622,I219773);
nand I_4573 (I80639,I80622,I219776);
not I_4574 (I80656,I219764);
nor I_4575 (I80673,I80656,I219755);
nand I_4576 (I80690,I80673,I219758);
nor I_4577 (I80707,I80690,I80639);
DFFARX1 I_4578 (I80707,I2859,I80489,I80457,);
not I_4579 (I80738,I80690);
not I_4580 (I80755,I219755);
nand I_4581 (I80772,I80755,I219776);
nor I_4582 (I80789,I219755,I219773);
nand I_4583 (I80469,I80605,I80789);
nand I_4584 (I80463,I80554,I219755);
nand I_4585 (I80834,I80656,I219779);
DFFARX1 I_4586 (I80834,I2859,I80489,I80478,);
DFFARX1 I_4587 (I80834,I2859,I80489,I80472,);
not I_4588 (I80879,I219779);
nor I_4589 (I80896,I80879,I219770);
and I_4590 (I80913,I80896,I219755);
or I_4591 (I80930,I80913,I219758);
DFFARX1 I_4592 (I80930,I2859,I80489,I80956,);
nand I_4593 (I80964,I80956,I80622);
nor I_4594 (I80466,I80964,I80772);
nor I_4595 (I80460,I80956,I80588);
DFFARX1 I_4596 (I80956,I2859,I80489,I81018,);
not I_4597 (I81026,I81018);
nor I_4598 (I80475,I81026,I80738);
not I_4599 (I81084,I2866);
DFFARX1 I_4600 (I304784,I2859,I81084,I81110,);
DFFARX1 I_4601 (I81110,I2859,I81084,I81127,);
not I_4602 (I81076,I81127);
not I_4603 (I81149,I81110);
DFFARX1 I_4604 (I304781,I2859,I81084,I81175,);
not I_4605 (I81183,I81175);
and I_4606 (I81200,I81149,I304787);
not I_4607 (I81217,I304772);
nand I_4608 (I81234,I81217,I304787);
not I_4609 (I81251,I304775);
nor I_4610 (I81268,I81251,I304796);
nand I_4611 (I81285,I81268,I304793);
nor I_4612 (I81302,I81285,I81234);
DFFARX1 I_4613 (I81302,I2859,I81084,I81052,);
not I_4614 (I81333,I81285);
not I_4615 (I81350,I304796);
nand I_4616 (I81367,I81350,I304787);
nor I_4617 (I81384,I304796,I304772);
nand I_4618 (I81064,I81200,I81384);
nand I_4619 (I81058,I81149,I304796);
nand I_4620 (I81429,I81251,I304772);
DFFARX1 I_4621 (I81429,I2859,I81084,I81073,);
DFFARX1 I_4622 (I81429,I2859,I81084,I81067,);
not I_4623 (I81474,I304772);
nor I_4624 (I81491,I81474,I304778);
and I_4625 (I81508,I81491,I304790);
or I_4626 (I81525,I81508,I304775);
DFFARX1 I_4627 (I81525,I2859,I81084,I81551,);
nand I_4628 (I81559,I81551,I81217);
nor I_4629 (I81061,I81559,I81367);
nor I_4630 (I81055,I81551,I81183);
DFFARX1 I_4631 (I81551,I2859,I81084,I81613,);
not I_4632 (I81621,I81613);
nor I_4633 (I81070,I81621,I81333);
not I_4634 (I81679,I2866);
DFFARX1 I_4635 (I377326,I2859,I81679,I81705,);
DFFARX1 I_4636 (I81705,I2859,I81679,I81722,);
not I_4637 (I81671,I81722);
not I_4638 (I81744,I81705);
DFFARX1 I_4639 (I377335,I2859,I81679,I81770,);
not I_4640 (I81778,I81770);
and I_4641 (I81795,I81744,I377323);
not I_4642 (I81812,I377314);
nand I_4643 (I81829,I81812,I377323);
not I_4644 (I81846,I377320);
nor I_4645 (I81863,I81846,I377338);
nand I_4646 (I81880,I81863,I377311);
nor I_4647 (I81897,I81880,I81829);
DFFARX1 I_4648 (I81897,I2859,I81679,I81647,);
not I_4649 (I81928,I81880);
not I_4650 (I81945,I377338);
nand I_4651 (I81962,I81945,I377323);
nor I_4652 (I81979,I377338,I377314);
nand I_4653 (I81659,I81795,I81979);
nand I_4654 (I81653,I81744,I377338);
nand I_4655 (I82024,I81846,I377317);
DFFARX1 I_4656 (I82024,I2859,I81679,I81668,);
DFFARX1 I_4657 (I82024,I2859,I81679,I81662,);
not I_4658 (I82069,I377317);
nor I_4659 (I82086,I82069,I377329);
and I_4660 (I82103,I82086,I377311);
or I_4661 (I82120,I82103,I377332);
DFFARX1 I_4662 (I82120,I2859,I81679,I82146,);
nand I_4663 (I82154,I82146,I81812);
nor I_4664 (I81656,I82154,I81962);
nor I_4665 (I81650,I82146,I81778);
DFFARX1 I_4666 (I82146,I2859,I81679,I82208,);
not I_4667 (I82216,I82208);
nor I_4668 (I81665,I82216,I81928);
not I_4669 (I82274,I2866);
DFFARX1 I_4670 (I187088,I2859,I82274,I82300,);
DFFARX1 I_4671 (I82300,I2859,I82274,I82317,);
not I_4672 (I82266,I82317);
not I_4673 (I82339,I82300);
DFFARX1 I_4674 (I187076,I2859,I82274,I82365,);
not I_4675 (I82373,I82365);
and I_4676 (I82390,I82339,I187085);
not I_4677 (I82407,I187082);
nand I_4678 (I82424,I82407,I187085);
not I_4679 (I82441,I187073);
nor I_4680 (I82458,I82441,I187079);
nand I_4681 (I82475,I82458,I187064);
nor I_4682 (I82492,I82475,I82424);
DFFARX1 I_4683 (I82492,I2859,I82274,I82242,);
not I_4684 (I82523,I82475);
not I_4685 (I82540,I187079);
nand I_4686 (I82557,I82540,I187085);
nor I_4687 (I82574,I187079,I187082);
nand I_4688 (I82254,I82390,I82574);
nand I_4689 (I82248,I82339,I187079);
nand I_4690 (I82619,I82441,I187064);
DFFARX1 I_4691 (I82619,I2859,I82274,I82263,);
DFFARX1 I_4692 (I82619,I2859,I82274,I82257,);
not I_4693 (I82664,I187064);
nor I_4694 (I82681,I82664,I187070);
and I_4695 (I82698,I82681,I187067);
or I_4696 (I82715,I82698,I187091);
DFFARX1 I_4697 (I82715,I2859,I82274,I82741,);
nand I_4698 (I82749,I82741,I82407);
nor I_4699 (I82251,I82749,I82557);
nor I_4700 (I82245,I82741,I82373);
DFFARX1 I_4701 (I82741,I2859,I82274,I82803,);
not I_4702 (I82811,I82803);
nor I_4703 (I82260,I82811,I82523);
not I_4704 (I82869,I2866);
DFFARX1 I_4705 (I448150,I2859,I82869,I82895,);
DFFARX1 I_4706 (I82895,I2859,I82869,I82912,);
not I_4707 (I82861,I82912);
not I_4708 (I82934,I82895);
DFFARX1 I_4709 (I448150,I2859,I82869,I82960,);
not I_4710 (I82968,I82960);
and I_4711 (I82985,I82934,I448153);
not I_4712 (I83002,I448165);
nand I_4713 (I83019,I83002,I448153);
not I_4714 (I83036,I448171);
nor I_4715 (I83053,I83036,I448162);
nand I_4716 (I83070,I83053,I448168);
nor I_4717 (I83087,I83070,I83019);
DFFARX1 I_4718 (I83087,I2859,I82869,I82837,);
not I_4719 (I83118,I83070);
not I_4720 (I83135,I448162);
nand I_4721 (I83152,I83135,I448153);
nor I_4722 (I83169,I448162,I448165);
nand I_4723 (I82849,I82985,I83169);
nand I_4724 (I82843,I82934,I448162);
nand I_4725 (I83214,I83036,I448159);
DFFARX1 I_4726 (I83214,I2859,I82869,I82858,);
DFFARX1 I_4727 (I83214,I2859,I82869,I82852,);
not I_4728 (I83259,I448159);
nor I_4729 (I83276,I83259,I448156);
and I_4730 (I83293,I83276,I448174);
or I_4731 (I83310,I83293,I448153);
DFFARX1 I_4732 (I83310,I2859,I82869,I83336,);
nand I_4733 (I83344,I83336,I83002);
nor I_4734 (I82846,I83344,I83152);
nor I_4735 (I82840,I83336,I82968);
DFFARX1 I_4736 (I83336,I2859,I82869,I83398,);
not I_4737 (I83406,I83398);
nor I_4738 (I82855,I83406,I83118);
not I_4739 (I83464,I2866);
DFFARX1 I_4740 (I233115,I2859,I83464,I83490,);
DFFARX1 I_4741 (I83490,I2859,I83464,I83507,);
not I_4742 (I83456,I83507);
not I_4743 (I83529,I83490);
DFFARX1 I_4744 (I233106,I2859,I83464,I83555,);
not I_4745 (I83563,I83555);
and I_4746 (I83580,I83529,I233124);
not I_4747 (I83597,I233121);
nand I_4748 (I83614,I83597,I233124);
not I_4749 (I83631,I233100);
nor I_4750 (I83648,I83631,I233103);
nand I_4751 (I83665,I83648,I233112);
nor I_4752 (I83682,I83665,I83614);
DFFARX1 I_4753 (I83682,I2859,I83464,I83432,);
not I_4754 (I83713,I83665);
not I_4755 (I83730,I233103);
nand I_4756 (I83747,I83730,I233124);
nor I_4757 (I83764,I233103,I233121);
nand I_4758 (I83444,I83580,I83764);
nand I_4759 (I83438,I83529,I233103);
nand I_4760 (I83809,I83631,I233118);
DFFARX1 I_4761 (I83809,I2859,I83464,I83453,);
DFFARX1 I_4762 (I83809,I2859,I83464,I83447,);
not I_4763 (I83854,I233118);
nor I_4764 (I83871,I83854,I233100);
and I_4765 (I83888,I83871,I233109);
or I_4766 (I83905,I83888,I233103);
DFFARX1 I_4767 (I83905,I2859,I83464,I83931,);
nand I_4768 (I83939,I83931,I83597);
nor I_4769 (I83441,I83939,I83747);
nor I_4770 (I83435,I83931,I83563);
DFFARX1 I_4771 (I83931,I2859,I83464,I83993,);
not I_4772 (I84001,I83993);
nor I_4773 (I83450,I84001,I83713);
not I_4774 (I84059,I2866);
DFFARX1 I_4775 (I243519,I2859,I84059,I84085,);
DFFARX1 I_4776 (I84085,I2859,I84059,I84102,);
not I_4777 (I84051,I84102);
not I_4778 (I84124,I84085);
DFFARX1 I_4779 (I243510,I2859,I84059,I84150,);
not I_4780 (I84158,I84150);
and I_4781 (I84175,I84124,I243528);
not I_4782 (I84192,I243525);
nand I_4783 (I84209,I84192,I243528);
not I_4784 (I84226,I243504);
nor I_4785 (I84243,I84226,I243507);
nand I_4786 (I84260,I84243,I243516);
nor I_4787 (I84277,I84260,I84209);
DFFARX1 I_4788 (I84277,I2859,I84059,I84027,);
not I_4789 (I84308,I84260);
not I_4790 (I84325,I243507);
nand I_4791 (I84342,I84325,I243528);
nor I_4792 (I84359,I243507,I243525);
nand I_4793 (I84039,I84175,I84359);
nand I_4794 (I84033,I84124,I243507);
nand I_4795 (I84404,I84226,I243522);
DFFARX1 I_4796 (I84404,I2859,I84059,I84048,);
DFFARX1 I_4797 (I84404,I2859,I84059,I84042,);
not I_4798 (I84449,I243522);
nor I_4799 (I84466,I84449,I243504);
and I_4800 (I84483,I84466,I243513);
or I_4801 (I84500,I84483,I243507);
DFFARX1 I_4802 (I84500,I2859,I84059,I84526,);
nand I_4803 (I84534,I84526,I84192);
nor I_4804 (I84036,I84534,I84342);
nor I_4805 (I84030,I84526,I84158);
DFFARX1 I_4806 (I84526,I2859,I84059,I84588,);
not I_4807 (I84596,I84588);
nor I_4808 (I84045,I84596,I84308);
not I_4809 (I84654,I2866);
DFFARX1 I_4810 (I532208,I2859,I84654,I84680,);
DFFARX1 I_4811 (I84680,I2859,I84654,I84697,);
not I_4812 (I84646,I84697);
not I_4813 (I84719,I84680);
DFFARX1 I_4814 (I532181,I2859,I84654,I84745,);
not I_4815 (I84753,I84745);
and I_4816 (I84770,I84719,I532205);
not I_4817 (I84787,I532202);
nand I_4818 (I84804,I84787,I532205);
not I_4819 (I84821,I532181);
nor I_4820 (I84838,I84821,I532199);
nand I_4821 (I84855,I84838,I532187);
nor I_4822 (I84872,I84855,I84804);
DFFARX1 I_4823 (I84872,I2859,I84654,I84622,);
not I_4824 (I84903,I84855);
not I_4825 (I84920,I532199);
nand I_4826 (I84937,I84920,I532205);
nor I_4827 (I84954,I532199,I532202);
nand I_4828 (I84634,I84770,I84954);
nand I_4829 (I84628,I84719,I532199);
nand I_4830 (I84999,I84821,I532193);
DFFARX1 I_4831 (I84999,I2859,I84654,I84643,);
DFFARX1 I_4832 (I84999,I2859,I84654,I84637,);
not I_4833 (I85044,I532193);
nor I_4834 (I85061,I85044,I532196);
and I_4835 (I85078,I85061,I532184);
or I_4836 (I85095,I85078,I532190);
DFFARX1 I_4837 (I85095,I2859,I84654,I85121,);
nand I_4838 (I85129,I85121,I84787);
nor I_4839 (I84631,I85129,I84937);
nor I_4840 (I84625,I85121,I84753);
DFFARX1 I_4841 (I85121,I2859,I84654,I85183,);
not I_4842 (I85191,I85183);
nor I_4843 (I84640,I85191,I84903);
not I_4844 (I85249,I2866);
DFFARX1 I_4845 (I468958,I2859,I85249,I85275,);
DFFARX1 I_4846 (I85275,I2859,I85249,I85292,);
not I_4847 (I85241,I85292);
not I_4848 (I85314,I85275);
DFFARX1 I_4849 (I468958,I2859,I85249,I85340,);
not I_4850 (I85348,I85340);
and I_4851 (I85365,I85314,I468961);
not I_4852 (I85382,I468973);
nand I_4853 (I85399,I85382,I468961);
not I_4854 (I85416,I468979);
nor I_4855 (I85433,I85416,I468970);
nand I_4856 (I85450,I85433,I468976);
nor I_4857 (I85467,I85450,I85399);
DFFARX1 I_4858 (I85467,I2859,I85249,I85217,);
not I_4859 (I85498,I85450);
not I_4860 (I85515,I468970);
nand I_4861 (I85532,I85515,I468961);
nor I_4862 (I85549,I468970,I468973);
nand I_4863 (I85229,I85365,I85549);
nand I_4864 (I85223,I85314,I468970);
nand I_4865 (I85594,I85416,I468967);
DFFARX1 I_4866 (I85594,I2859,I85249,I85238,);
DFFARX1 I_4867 (I85594,I2859,I85249,I85232,);
not I_4868 (I85639,I468967);
nor I_4869 (I85656,I85639,I468964);
and I_4870 (I85673,I85656,I468982);
or I_4871 (I85690,I85673,I468961);
DFFARX1 I_4872 (I85690,I2859,I85249,I85716,);
nand I_4873 (I85724,I85716,I85382);
nor I_4874 (I85226,I85724,I85532);
nor I_4875 (I85220,I85716,I85348);
DFFARX1 I_4876 (I85716,I2859,I85249,I85778,);
not I_4877 (I85786,I85778);
nor I_4878 (I85235,I85786,I85498);
not I_4879 (I85844,I2866);
DFFARX1 I_4880 (I514468,I2859,I85844,I85870,);
DFFARX1 I_4881 (I85870,I2859,I85844,I85887,);
not I_4882 (I85836,I85887);
not I_4883 (I85909,I85870);
DFFARX1 I_4884 (I514453,I2859,I85844,I85935,);
not I_4885 (I85943,I85935);
and I_4886 (I85960,I85909,I514471);
not I_4887 (I85977,I514453);
nand I_4888 (I85994,I85977,I514471);
not I_4889 (I86011,I514474);
nor I_4890 (I86028,I86011,I514465);
nand I_4891 (I86045,I86028,I514462);
nor I_4892 (I86062,I86045,I85994);
DFFARX1 I_4893 (I86062,I2859,I85844,I85812,);
not I_4894 (I86093,I86045);
not I_4895 (I86110,I514465);
nand I_4896 (I86127,I86110,I514471);
nor I_4897 (I86144,I514465,I514453);
nand I_4898 (I85824,I85960,I86144);
nand I_4899 (I85818,I85909,I514465);
nand I_4900 (I86189,I86011,I514459);
DFFARX1 I_4901 (I86189,I2859,I85844,I85833,);
DFFARX1 I_4902 (I86189,I2859,I85844,I85827,);
not I_4903 (I86234,I514459);
nor I_4904 (I86251,I86234,I514450);
and I_4905 (I86268,I86251,I514456);
or I_4906 (I86285,I86268,I514450);
DFFARX1 I_4907 (I86285,I2859,I85844,I86311,);
nand I_4908 (I86319,I86311,I85977);
nor I_4909 (I85821,I86319,I86127);
nor I_4910 (I85815,I86311,I85943);
DFFARX1 I_4911 (I86311,I2859,I85844,I86373,);
not I_4912 (I86381,I86373);
nor I_4913 (I85830,I86381,I86093);
not I_4914 (I86439,I2866);
DFFARX1 I_4915 (I150395,I2859,I86439,I86465,);
DFFARX1 I_4916 (I86465,I2859,I86439,I86482,);
not I_4917 (I86431,I86482);
not I_4918 (I86504,I86465);
DFFARX1 I_4919 (I150410,I2859,I86439,I86530,);
not I_4920 (I86538,I86530);
and I_4921 (I86555,I86504,I150407);
not I_4922 (I86572,I150395);
nand I_4923 (I86589,I86572,I150407);
not I_4924 (I86606,I150404);
nor I_4925 (I86623,I86606,I150419);
nand I_4926 (I86640,I86623,I150416);
nor I_4927 (I86657,I86640,I86589);
DFFARX1 I_4928 (I86657,I2859,I86439,I86407,);
not I_4929 (I86688,I86640);
not I_4930 (I86705,I150419);
nand I_4931 (I86722,I86705,I150407);
nor I_4932 (I86739,I150419,I150395);
nand I_4933 (I86419,I86555,I86739);
nand I_4934 (I86413,I86504,I150419);
nand I_4935 (I86784,I86606,I150413);
DFFARX1 I_4936 (I86784,I2859,I86439,I86428,);
DFFARX1 I_4937 (I86784,I2859,I86439,I86422,);
not I_4938 (I86829,I150413);
nor I_4939 (I86846,I86829,I150401);
and I_4940 (I86863,I86846,I150422);
or I_4941 (I86880,I86863,I150398);
DFFARX1 I_4942 (I86880,I2859,I86439,I86906,);
nand I_4943 (I86914,I86906,I86572);
nor I_4944 (I86416,I86914,I86722);
nor I_4945 (I86410,I86906,I86538);
DFFARX1 I_4946 (I86906,I2859,I86439,I86968,);
not I_4947 (I86976,I86968);
nor I_4948 (I86425,I86976,I86688);
not I_4949 (I87034,I2866);
DFFARX1 I_4950 (I206082,I2859,I87034,I87060,);
DFFARX1 I_4951 (I87060,I2859,I87034,I87077,);
not I_4952 (I87026,I87077);
not I_4953 (I87099,I87060);
DFFARX1 I_4954 (I206076,I2859,I87034,I87125,);
not I_4955 (I87133,I87125);
and I_4956 (I87150,I87099,I206091);
not I_4957 (I87167,I206088);
nand I_4958 (I87184,I87167,I206091);
not I_4959 (I87201,I206079);
nor I_4960 (I87218,I87201,I206070);
nand I_4961 (I87235,I87218,I206073);
nor I_4962 (I87252,I87235,I87184);
DFFARX1 I_4963 (I87252,I2859,I87034,I87002,);
not I_4964 (I87283,I87235);
not I_4965 (I87300,I206070);
nand I_4966 (I87317,I87300,I206091);
nor I_4967 (I87334,I206070,I206088);
nand I_4968 (I87014,I87150,I87334);
nand I_4969 (I87008,I87099,I206070);
nand I_4970 (I87379,I87201,I206094);
DFFARX1 I_4971 (I87379,I2859,I87034,I87023,);
DFFARX1 I_4972 (I87379,I2859,I87034,I87017,);
not I_4973 (I87424,I206094);
nor I_4974 (I87441,I87424,I206085);
and I_4975 (I87458,I87441,I206070);
or I_4976 (I87475,I87458,I206073);
DFFARX1 I_4977 (I87475,I2859,I87034,I87501,);
nand I_4978 (I87509,I87501,I87167);
nor I_4979 (I87011,I87509,I87317);
nor I_4980 (I87005,I87501,I87133);
DFFARX1 I_4981 (I87501,I2859,I87034,I87563,);
not I_4982 (I87571,I87563);
nor I_4983 (I87020,I87571,I87283);
not I_4984 (I87629,I2866);
DFFARX1 I_4985 (I15881,I2859,I87629,I87655,);
DFFARX1 I_4986 (I87655,I2859,I87629,I87672,);
not I_4987 (I87621,I87672);
not I_4988 (I87694,I87655);
DFFARX1 I_4989 (I15857,I2859,I87629,I87720,);
not I_4990 (I87728,I87720);
and I_4991 (I87745,I87694,I15872);
not I_4992 (I87762,I15860);
nand I_4993 (I87779,I87762,I15872);
not I_4994 (I87796,I15863);
nor I_4995 (I87813,I87796,I15875);
nand I_4996 (I87830,I87813,I15866);
nor I_4997 (I87847,I87830,I87779);
DFFARX1 I_4998 (I87847,I2859,I87629,I87597,);
not I_4999 (I87878,I87830);
not I_5000 (I87895,I15875);
nand I_5001 (I87912,I87895,I15872);
nor I_5002 (I87929,I15875,I15860);
nand I_5003 (I87609,I87745,I87929);
nand I_5004 (I87603,I87694,I15875);
nand I_5005 (I87974,I87796,I15869);
DFFARX1 I_5006 (I87974,I2859,I87629,I87618,);
DFFARX1 I_5007 (I87974,I2859,I87629,I87612,);
not I_5008 (I88019,I15869);
nor I_5009 (I88036,I88019,I15860);
and I_5010 (I88053,I88036,I15857);
or I_5011 (I88070,I88053,I15878);
DFFARX1 I_5012 (I88070,I2859,I87629,I88096,);
nand I_5013 (I88104,I88096,I87762);
nor I_5014 (I87606,I88104,I87912);
nor I_5015 (I87600,I88096,I87728);
DFFARX1 I_5016 (I88096,I2859,I87629,I88158,);
not I_5017 (I88166,I88158);
nor I_5018 (I87615,I88166,I87878);
not I_5019 (I88224,I2866);
DFFARX1 I_5020 (I395414,I2859,I88224,I88250,);
DFFARX1 I_5021 (I88250,I2859,I88224,I88267,);
not I_5022 (I88216,I88267);
not I_5023 (I88289,I88250);
DFFARX1 I_5024 (I395423,I2859,I88224,I88315,);
not I_5025 (I88323,I88315);
and I_5026 (I88340,I88289,I395411);
not I_5027 (I88357,I395402);
nand I_5028 (I88374,I88357,I395411);
not I_5029 (I88391,I395408);
nor I_5030 (I88408,I88391,I395426);
nand I_5031 (I88425,I88408,I395399);
nor I_5032 (I88442,I88425,I88374);
DFFARX1 I_5033 (I88442,I2859,I88224,I88192,);
not I_5034 (I88473,I88425);
not I_5035 (I88490,I395426);
nand I_5036 (I88507,I88490,I395411);
nor I_5037 (I88524,I395426,I395402);
nand I_5038 (I88204,I88340,I88524);
nand I_5039 (I88198,I88289,I395426);
nand I_5040 (I88569,I88391,I395405);
DFFARX1 I_5041 (I88569,I2859,I88224,I88213,);
DFFARX1 I_5042 (I88569,I2859,I88224,I88207,);
not I_5043 (I88614,I395405);
nor I_5044 (I88631,I88614,I395417);
and I_5045 (I88648,I88631,I395399);
or I_5046 (I88665,I88648,I395420);
DFFARX1 I_5047 (I88665,I2859,I88224,I88691,);
nand I_5048 (I88699,I88691,I88357);
nor I_5049 (I88201,I88699,I88507);
nor I_5050 (I88195,I88691,I88323);
DFFARX1 I_5051 (I88691,I2859,I88224,I88753,);
not I_5052 (I88761,I88753);
nor I_5053 (I88210,I88761,I88473);
not I_5054 (I88819,I2866);
DFFARX1 I_5055 (I288600,I2859,I88819,I88845,);
DFFARX1 I_5056 (I88845,I2859,I88819,I88862,);
not I_5057 (I88811,I88862);
not I_5058 (I88884,I88845);
DFFARX1 I_5059 (I288597,I2859,I88819,I88910,);
not I_5060 (I88918,I88910);
and I_5061 (I88935,I88884,I288603);
not I_5062 (I88952,I288588);
nand I_5063 (I88969,I88952,I288603);
not I_5064 (I88986,I288591);
nor I_5065 (I89003,I88986,I288612);
nand I_5066 (I89020,I89003,I288609);
nor I_5067 (I89037,I89020,I88969);
DFFARX1 I_5068 (I89037,I2859,I88819,I88787,);
not I_5069 (I89068,I89020);
not I_5070 (I89085,I288612);
nand I_5071 (I89102,I89085,I288603);
nor I_5072 (I89119,I288612,I288588);
nand I_5073 (I88799,I88935,I89119);
nand I_5074 (I88793,I88884,I288612);
nand I_5075 (I89164,I88986,I288588);
DFFARX1 I_5076 (I89164,I2859,I88819,I88808,);
DFFARX1 I_5077 (I89164,I2859,I88819,I88802,);
not I_5078 (I89209,I288588);
nor I_5079 (I89226,I89209,I288594);
and I_5080 (I89243,I89226,I288606);
or I_5081 (I89260,I89243,I288591);
DFFARX1 I_5082 (I89260,I2859,I88819,I89286,);
nand I_5083 (I89294,I89286,I88952);
nor I_5084 (I88796,I89294,I89102);
nor I_5085 (I88790,I89286,I88918);
DFFARX1 I_5086 (I89286,I2859,I88819,I89348,);
not I_5087 (I89356,I89348);
nor I_5088 (I88805,I89356,I89068);
not I_5089 (I89414,I2866);
DFFARX1 I_5090 (I170224,I2859,I89414,I89440,);
DFFARX1 I_5091 (I89440,I2859,I89414,I89457,);
not I_5092 (I89406,I89457);
not I_5093 (I89479,I89440);
DFFARX1 I_5094 (I170212,I2859,I89414,I89505,);
not I_5095 (I89513,I89505);
and I_5096 (I89530,I89479,I170221);
not I_5097 (I89547,I170218);
nand I_5098 (I89564,I89547,I170221);
not I_5099 (I89581,I170209);
nor I_5100 (I89598,I89581,I170215);
nand I_5101 (I89615,I89598,I170200);
nor I_5102 (I89632,I89615,I89564);
DFFARX1 I_5103 (I89632,I2859,I89414,I89382,);
not I_5104 (I89663,I89615);
not I_5105 (I89680,I170215);
nand I_5106 (I89697,I89680,I170221);
nor I_5107 (I89714,I170215,I170218);
nand I_5108 (I89394,I89530,I89714);
nand I_5109 (I89388,I89479,I170215);
nand I_5110 (I89759,I89581,I170200);
DFFARX1 I_5111 (I89759,I2859,I89414,I89403,);
DFFARX1 I_5112 (I89759,I2859,I89414,I89397,);
not I_5113 (I89804,I170200);
nor I_5114 (I89821,I89804,I170206);
and I_5115 (I89838,I89821,I170203);
or I_5116 (I89855,I89838,I170227);
DFFARX1 I_5117 (I89855,I2859,I89414,I89881,);
nand I_5118 (I89889,I89881,I89547);
nor I_5119 (I89391,I89889,I89697);
nor I_5120 (I89385,I89881,I89513);
DFFARX1 I_5121 (I89881,I2859,I89414,I89943,);
not I_5122 (I89951,I89943);
nor I_5123 (I89400,I89951,I89663);
not I_5124 (I90009,I2866);
DFFARX1 I_5125 (I442948,I2859,I90009,I90035,);
DFFARX1 I_5126 (I90035,I2859,I90009,I90052,);
not I_5127 (I90001,I90052);
not I_5128 (I90074,I90035);
DFFARX1 I_5129 (I442948,I2859,I90009,I90100,);
not I_5130 (I90108,I90100);
and I_5131 (I90125,I90074,I442951);
not I_5132 (I90142,I442963);
nand I_5133 (I90159,I90142,I442951);
not I_5134 (I90176,I442969);
nor I_5135 (I90193,I90176,I442960);
nand I_5136 (I90210,I90193,I442966);
nor I_5137 (I90227,I90210,I90159);
DFFARX1 I_5138 (I90227,I2859,I90009,I89977,);
not I_5139 (I90258,I90210);
not I_5140 (I90275,I442960);
nand I_5141 (I90292,I90275,I442951);
nor I_5142 (I90309,I442960,I442963);
nand I_5143 (I89989,I90125,I90309);
nand I_5144 (I89983,I90074,I442960);
nand I_5145 (I90354,I90176,I442957);
DFFARX1 I_5146 (I90354,I2859,I90009,I89998,);
DFFARX1 I_5147 (I90354,I2859,I90009,I89992,);
not I_5148 (I90399,I442957);
nor I_5149 (I90416,I90399,I442954);
and I_5150 (I90433,I90416,I442972);
or I_5151 (I90450,I90433,I442951);
DFFARX1 I_5152 (I90450,I2859,I90009,I90476,);
nand I_5153 (I90484,I90476,I90142);
nor I_5154 (I89986,I90484,I90292);
nor I_5155 (I89980,I90476,I90108);
DFFARX1 I_5156 (I90476,I2859,I90009,I90538,);
not I_5157 (I90546,I90538);
nor I_5158 (I89995,I90546,I90258);
not I_5159 (I90604,I2866);
DFFARX1 I_5160 (I33784,I2859,I90604,I90630,);
DFFARX1 I_5161 (I90630,I2859,I90604,I90647,);
not I_5162 (I90596,I90647);
not I_5163 (I90669,I90630);
DFFARX1 I_5164 (I33778,I2859,I90604,I90695,);
not I_5165 (I90703,I90695);
and I_5166 (I90720,I90669,I33775);
not I_5167 (I90737,I33796);
nand I_5168 (I90754,I90737,I33775);
not I_5169 (I90771,I33790);
nor I_5170 (I90788,I90771,I33781);
nand I_5171 (I90805,I90788,I33787);
nor I_5172 (I90822,I90805,I90754);
DFFARX1 I_5173 (I90822,I2859,I90604,I90572,);
not I_5174 (I90853,I90805);
not I_5175 (I90870,I33781);
nand I_5176 (I90887,I90870,I33775);
nor I_5177 (I90904,I33781,I33796);
nand I_5178 (I90584,I90720,I90904);
nand I_5179 (I90578,I90669,I33781);
nand I_5180 (I90949,I90771,I33775);
DFFARX1 I_5181 (I90949,I2859,I90604,I90593,);
DFFARX1 I_5182 (I90949,I2859,I90604,I90587,);
not I_5183 (I90994,I33775);
nor I_5184 (I91011,I90994,I33793);
and I_5185 (I91028,I91011,I33799);
or I_5186 (I91045,I91028,I33778);
DFFARX1 I_5187 (I91045,I2859,I90604,I91071,);
nand I_5188 (I91079,I91071,I90737);
nor I_5189 (I90581,I91079,I90887);
nor I_5190 (I90575,I91071,I90703);
DFFARX1 I_5191 (I91071,I2859,I90604,I91133,);
not I_5192 (I91141,I91133);
nor I_5193 (I90590,I91141,I90853);
not I_5194 (I91199,I2866);
DFFARX1 I_5195 (I330193,I2859,I91199,I91225,);
DFFARX1 I_5196 (I91225,I2859,I91199,I91242,);
not I_5197 (I91191,I91242);
not I_5198 (I91264,I91225);
DFFARX1 I_5199 (I330187,I2859,I91199,I91290,);
not I_5200 (I91298,I91290);
and I_5201 (I91315,I91264,I330205);
not I_5202 (I91332,I330193);
nand I_5203 (I91349,I91332,I330205);
not I_5204 (I91366,I330187);
nor I_5205 (I91383,I91366,I330199);
nand I_5206 (I91400,I91383,I330190);
nor I_5207 (I91417,I91400,I91349);
DFFARX1 I_5208 (I91417,I2859,I91199,I91167,);
not I_5209 (I91448,I91400);
not I_5210 (I91465,I330199);
nand I_5211 (I91482,I91465,I330205);
nor I_5212 (I91499,I330199,I330193);
nand I_5213 (I91179,I91315,I91499);
nand I_5214 (I91173,I91264,I330199);
nand I_5215 (I91544,I91366,I330202);
DFFARX1 I_5216 (I91544,I2859,I91199,I91188,);
DFFARX1 I_5217 (I91544,I2859,I91199,I91182,);
not I_5218 (I91589,I330202);
nor I_5219 (I91606,I91589,I330208);
and I_5220 (I91623,I91606,I330190);
or I_5221 (I91640,I91623,I330196);
DFFARX1 I_5222 (I91640,I2859,I91199,I91666,);
nand I_5223 (I91674,I91666,I91332);
nor I_5224 (I91176,I91674,I91482);
nor I_5225 (I91170,I91666,I91298);
DFFARX1 I_5226 (I91666,I2859,I91199,I91728,);
not I_5227 (I91736,I91728);
nor I_5228 (I91185,I91736,I91448);
not I_5229 (I91794,I2866);
DFFARX1 I_5230 (I27987,I2859,I91794,I91820,);
DFFARX1 I_5231 (I91820,I2859,I91794,I91837,);
not I_5232 (I91786,I91837);
not I_5233 (I91859,I91820);
DFFARX1 I_5234 (I27981,I2859,I91794,I91885,);
not I_5235 (I91893,I91885);
and I_5236 (I91910,I91859,I27978);
not I_5237 (I91927,I27999);
nand I_5238 (I91944,I91927,I27978);
not I_5239 (I91961,I27993);
nor I_5240 (I91978,I91961,I27984);
nand I_5241 (I91995,I91978,I27990);
nor I_5242 (I92012,I91995,I91944);
DFFARX1 I_5243 (I92012,I2859,I91794,I91762,);
not I_5244 (I92043,I91995);
not I_5245 (I92060,I27984);
nand I_5246 (I92077,I92060,I27978);
nor I_5247 (I92094,I27984,I27999);
nand I_5248 (I91774,I91910,I92094);
nand I_5249 (I91768,I91859,I27984);
nand I_5250 (I92139,I91961,I27978);
DFFARX1 I_5251 (I92139,I2859,I91794,I91783,);
DFFARX1 I_5252 (I92139,I2859,I91794,I91777,);
not I_5253 (I92184,I27978);
nor I_5254 (I92201,I92184,I27996);
and I_5255 (I92218,I92201,I28002);
or I_5256 (I92235,I92218,I27981);
DFFARX1 I_5257 (I92235,I2859,I91794,I92261,);
nand I_5258 (I92269,I92261,I91927);
nor I_5259 (I91771,I92269,I92077);
nor I_5260 (I91765,I92261,I91893);
DFFARX1 I_5261 (I92261,I2859,I91794,I92323,);
not I_5262 (I92331,I92323);
nor I_5263 (I91780,I92331,I92043);
not I_5264 (I92389,I2866);
DFFARX1 I_5265 (I323869,I2859,I92389,I92415,);
DFFARX1 I_5266 (I92415,I2859,I92389,I92432,);
not I_5267 (I92381,I92432);
not I_5268 (I92454,I92415);
DFFARX1 I_5269 (I323863,I2859,I92389,I92480,);
not I_5270 (I92488,I92480);
and I_5271 (I92505,I92454,I323881);
not I_5272 (I92522,I323869);
nand I_5273 (I92539,I92522,I323881);
not I_5274 (I92556,I323863);
nor I_5275 (I92573,I92556,I323875);
nand I_5276 (I92590,I92573,I323866);
nor I_5277 (I92607,I92590,I92539);
DFFARX1 I_5278 (I92607,I2859,I92389,I92357,);
not I_5279 (I92638,I92590);
not I_5280 (I92655,I323875);
nand I_5281 (I92672,I92655,I323881);
nor I_5282 (I92689,I323875,I323869);
nand I_5283 (I92369,I92505,I92689);
nand I_5284 (I92363,I92454,I323875);
nand I_5285 (I92734,I92556,I323878);
DFFARX1 I_5286 (I92734,I2859,I92389,I92378,);
DFFARX1 I_5287 (I92734,I2859,I92389,I92372,);
not I_5288 (I92779,I323878);
nor I_5289 (I92796,I92779,I323884);
and I_5290 (I92813,I92796,I323866);
or I_5291 (I92830,I92813,I323872);
DFFARX1 I_5292 (I92830,I2859,I92389,I92856,);
nand I_5293 (I92864,I92856,I92522);
nor I_5294 (I92366,I92864,I92672);
nor I_5295 (I92360,I92856,I92488);
DFFARX1 I_5296 (I92856,I2859,I92389,I92918,);
not I_5297 (I92926,I92918);
nor I_5298 (I92375,I92926,I92638);
not I_5299 (I92984,I2866);
DFFARX1 I_5300 (I366990,I2859,I92984,I93010,);
DFFARX1 I_5301 (I93010,I2859,I92984,I93027,);
not I_5302 (I92976,I93027);
not I_5303 (I93049,I93010);
DFFARX1 I_5304 (I366999,I2859,I92984,I93075,);
not I_5305 (I93083,I93075);
and I_5306 (I93100,I93049,I366987);
not I_5307 (I93117,I366978);
nand I_5308 (I93134,I93117,I366987);
not I_5309 (I93151,I366984);
nor I_5310 (I93168,I93151,I367002);
nand I_5311 (I93185,I93168,I366975);
nor I_5312 (I93202,I93185,I93134);
DFFARX1 I_5313 (I93202,I2859,I92984,I92952,);
not I_5314 (I93233,I93185);
not I_5315 (I93250,I367002);
nand I_5316 (I93267,I93250,I366987);
nor I_5317 (I93284,I367002,I366978);
nand I_5318 (I92964,I93100,I93284);
nand I_5319 (I92958,I93049,I367002);
nand I_5320 (I93329,I93151,I366981);
DFFARX1 I_5321 (I93329,I2859,I92984,I92973,);
DFFARX1 I_5322 (I93329,I2859,I92984,I92967,);
not I_5323 (I93374,I366981);
nor I_5324 (I93391,I93374,I366993);
and I_5325 (I93408,I93391,I366975);
or I_5326 (I93425,I93408,I366996);
DFFARX1 I_5327 (I93425,I2859,I92984,I93451,);
nand I_5328 (I93459,I93451,I93117);
nor I_5329 (I92961,I93459,I93267);
nor I_5330 (I92955,I93451,I93083);
DFFARX1 I_5331 (I93451,I2859,I92984,I93513,);
not I_5332 (I93521,I93513);
nor I_5333 (I92970,I93521,I93233);
not I_5334 (I93579,I2866);
DFFARX1 I_5335 (I475316,I2859,I93579,I93605,);
DFFARX1 I_5336 (I93605,I2859,I93579,I93622,);
not I_5337 (I93571,I93622);
not I_5338 (I93644,I93605);
DFFARX1 I_5339 (I475316,I2859,I93579,I93670,);
not I_5340 (I93678,I93670);
and I_5341 (I93695,I93644,I475319);
not I_5342 (I93712,I475331);
nand I_5343 (I93729,I93712,I475319);
not I_5344 (I93746,I475337);
nor I_5345 (I93763,I93746,I475328);
nand I_5346 (I93780,I93763,I475334);
nor I_5347 (I93797,I93780,I93729);
DFFARX1 I_5348 (I93797,I2859,I93579,I93547,);
not I_5349 (I93828,I93780);
not I_5350 (I93845,I475328);
nand I_5351 (I93862,I93845,I475319);
nor I_5352 (I93879,I475328,I475331);
nand I_5353 (I93559,I93695,I93879);
nand I_5354 (I93553,I93644,I475328);
nand I_5355 (I93924,I93746,I475325);
DFFARX1 I_5356 (I93924,I2859,I93579,I93568,);
DFFARX1 I_5357 (I93924,I2859,I93579,I93562,);
not I_5358 (I93969,I475325);
nor I_5359 (I93986,I93969,I475322);
and I_5360 (I94003,I93986,I475340);
or I_5361 (I94020,I94003,I475319);
DFFARX1 I_5362 (I94020,I2859,I93579,I94046,);
nand I_5363 (I94054,I94046,I93712);
nor I_5364 (I93556,I94054,I93862);
nor I_5365 (I93550,I94046,I93678);
DFFARX1 I_5366 (I94046,I2859,I93579,I94108,);
not I_5367 (I94116,I94108);
nor I_5368 (I93565,I94116,I93828);
not I_5369 (I94174,I2866);
DFFARX1 I_5370 (I418709,I2859,I94174,I94200,);
DFFARX1 I_5371 (I94200,I2859,I94174,I94217,);
not I_5372 (I94166,I94217);
not I_5373 (I94239,I94200);
DFFARX1 I_5374 (I418718,I2859,I94174,I94265,);
not I_5375 (I94273,I94265);
and I_5376 (I94290,I94239,I418712);
not I_5377 (I94307,I418706);
nand I_5378 (I94324,I94307,I418712);
not I_5379 (I94341,I418721);
nor I_5380 (I94358,I94341,I418709);
nand I_5381 (I94375,I94358,I418715);
nor I_5382 (I94392,I94375,I94324);
DFFARX1 I_5383 (I94392,I2859,I94174,I94142,);
not I_5384 (I94423,I94375);
not I_5385 (I94440,I418709);
nand I_5386 (I94457,I94440,I418712);
nor I_5387 (I94474,I418709,I418706);
nand I_5388 (I94154,I94290,I94474);
nand I_5389 (I94148,I94239,I418709);
nand I_5390 (I94519,I94341,I418712);
DFFARX1 I_5391 (I94519,I2859,I94174,I94163,);
DFFARX1 I_5392 (I94519,I2859,I94174,I94157,);
not I_5393 (I94564,I418712);
nor I_5394 (I94581,I94564,I418727);
and I_5395 (I94598,I94581,I418724);
or I_5396 (I94615,I94598,I418706);
DFFARX1 I_5397 (I94615,I2859,I94174,I94641,);
nand I_5398 (I94649,I94641,I94307);
nor I_5399 (I94151,I94649,I94457);
nor I_5400 (I94145,I94641,I94273);
DFFARX1 I_5401 (I94641,I2859,I94174,I94703,);
not I_5402 (I94711,I94703);
nor I_5403 (I94160,I94711,I94423);
not I_5404 (I94769,I2866);
DFFARX1 I_5405 (I131423,I2859,I94769,I94795,);
DFFARX1 I_5406 (I94795,I2859,I94769,I94812,);
not I_5407 (I94761,I94812);
not I_5408 (I94834,I94795);
DFFARX1 I_5409 (I131438,I2859,I94769,I94860,);
not I_5410 (I94868,I94860);
and I_5411 (I94885,I94834,I131435);
not I_5412 (I94902,I131423);
nand I_5413 (I94919,I94902,I131435);
not I_5414 (I94936,I131432);
nor I_5415 (I94953,I94936,I131447);
nand I_5416 (I94970,I94953,I131444);
nor I_5417 (I94987,I94970,I94919);
DFFARX1 I_5418 (I94987,I2859,I94769,I94737,);
not I_5419 (I95018,I94970);
not I_5420 (I95035,I131447);
nand I_5421 (I95052,I95035,I131435);
nor I_5422 (I95069,I131447,I131423);
nand I_5423 (I94749,I94885,I95069);
nand I_5424 (I94743,I94834,I131447);
nand I_5425 (I95114,I94936,I131441);
DFFARX1 I_5426 (I95114,I2859,I94769,I94758,);
DFFARX1 I_5427 (I95114,I2859,I94769,I94752,);
not I_5428 (I95159,I131441);
nor I_5429 (I95176,I95159,I131429);
and I_5430 (I95193,I95176,I131450);
or I_5431 (I95210,I95193,I131426);
DFFARX1 I_5432 (I95210,I2859,I94769,I95236,);
nand I_5433 (I95244,I95236,I94902);
nor I_5434 (I94746,I95244,I95052);
nor I_5435 (I94740,I95236,I94868);
DFFARX1 I_5436 (I95236,I2859,I94769,I95298,);
not I_5437 (I95306,I95298);
nor I_5438 (I94755,I95306,I95018);
not I_5439 (I95364,I2866);
DFFARX1 I_5440 (I321761,I2859,I95364,I95390,);
DFFARX1 I_5441 (I95390,I2859,I95364,I95407,);
not I_5442 (I95356,I95407);
not I_5443 (I95429,I95390);
DFFARX1 I_5444 (I321755,I2859,I95364,I95455,);
not I_5445 (I95463,I95455);
and I_5446 (I95480,I95429,I321773);
not I_5447 (I95497,I321761);
nand I_5448 (I95514,I95497,I321773);
not I_5449 (I95531,I321755);
nor I_5450 (I95548,I95531,I321767);
nand I_5451 (I95565,I95548,I321758);
nor I_5452 (I95582,I95565,I95514);
DFFARX1 I_5453 (I95582,I2859,I95364,I95332,);
not I_5454 (I95613,I95565);
not I_5455 (I95630,I321767);
nand I_5456 (I95647,I95630,I321773);
nor I_5457 (I95664,I321767,I321761);
nand I_5458 (I95344,I95480,I95664);
nand I_5459 (I95338,I95429,I321767);
nand I_5460 (I95709,I95531,I321770);
DFFARX1 I_5461 (I95709,I2859,I95364,I95353,);
DFFARX1 I_5462 (I95709,I2859,I95364,I95347,);
not I_5463 (I95754,I321770);
nor I_5464 (I95771,I95754,I321776);
and I_5465 (I95788,I95771,I321758);
or I_5466 (I95805,I95788,I321764);
DFFARX1 I_5467 (I95805,I2859,I95364,I95831,);
nand I_5468 (I95839,I95831,I95497);
nor I_5469 (I95341,I95839,I95647);
nor I_5470 (I95335,I95831,I95463);
DFFARX1 I_5471 (I95831,I2859,I95364,I95893,);
not I_5472 (I95901,I95893);
nor I_5473 (I95350,I95901,I95613);
not I_5474 (I95959,I2866);
DFFARX1 I_5475 (I213222,I2859,I95959,I95985,);
DFFARX1 I_5476 (I95985,I2859,I95959,I96002,);
not I_5477 (I95951,I96002);
not I_5478 (I96024,I95985);
DFFARX1 I_5479 (I213216,I2859,I95959,I96050,);
not I_5480 (I96058,I96050);
and I_5481 (I96075,I96024,I213231);
not I_5482 (I96092,I213228);
nand I_5483 (I96109,I96092,I213231);
not I_5484 (I96126,I213219);
nor I_5485 (I96143,I96126,I213210);
nand I_5486 (I96160,I96143,I213213);
nor I_5487 (I96177,I96160,I96109);
DFFARX1 I_5488 (I96177,I2859,I95959,I95927,);
not I_5489 (I96208,I96160);
not I_5490 (I96225,I213210);
nand I_5491 (I96242,I96225,I213231);
nor I_5492 (I96259,I213210,I213228);
nand I_5493 (I95939,I96075,I96259);
nand I_5494 (I95933,I96024,I213210);
nand I_5495 (I96304,I96126,I213234);
DFFARX1 I_5496 (I96304,I2859,I95959,I95948,);
DFFARX1 I_5497 (I96304,I2859,I95959,I95942,);
not I_5498 (I96349,I213234);
nor I_5499 (I96366,I96349,I213225);
and I_5500 (I96383,I96366,I213210);
or I_5501 (I96400,I96383,I213213);
DFFARX1 I_5502 (I96400,I2859,I95959,I96426,);
nand I_5503 (I96434,I96426,I96092);
nor I_5504 (I95936,I96434,I96242);
nor I_5505 (I95930,I96426,I96058);
DFFARX1 I_5506 (I96426,I2859,I95959,I96488,);
not I_5507 (I96496,I96488);
nor I_5508 (I95945,I96496,I96208);
not I_5509 (I96554,I2866);
DFFARX1 I_5510 (I10084,I2859,I96554,I96580,);
DFFARX1 I_5511 (I96580,I2859,I96554,I96597,);
not I_5512 (I96546,I96597);
not I_5513 (I96619,I96580);
DFFARX1 I_5514 (I10060,I2859,I96554,I96645,);
not I_5515 (I96653,I96645);
and I_5516 (I96670,I96619,I10075);
not I_5517 (I96687,I10063);
nand I_5518 (I96704,I96687,I10075);
not I_5519 (I96721,I10066);
nor I_5520 (I96738,I96721,I10078);
nand I_5521 (I96755,I96738,I10069);
nor I_5522 (I96772,I96755,I96704);
DFFARX1 I_5523 (I96772,I2859,I96554,I96522,);
not I_5524 (I96803,I96755);
not I_5525 (I96820,I10078);
nand I_5526 (I96837,I96820,I10075);
nor I_5527 (I96854,I10078,I10063);
nand I_5528 (I96534,I96670,I96854);
nand I_5529 (I96528,I96619,I10078);
nand I_5530 (I96899,I96721,I10072);
DFFARX1 I_5531 (I96899,I2859,I96554,I96543,);
DFFARX1 I_5532 (I96899,I2859,I96554,I96537,);
not I_5533 (I96944,I10072);
nor I_5534 (I96961,I96944,I10063);
and I_5535 (I96978,I96961,I10060);
or I_5536 (I96995,I96978,I10081);
DFFARX1 I_5537 (I96995,I2859,I96554,I97021,);
nand I_5538 (I97029,I97021,I96687);
nor I_5539 (I96531,I97029,I96837);
nor I_5540 (I96525,I97021,I96653);
DFFARX1 I_5541 (I97021,I2859,I96554,I97083,);
not I_5542 (I97091,I97083);
nor I_5543 (I96540,I97091,I96803);
not I_5544 (I97149,I2866);
DFFARX1 I_5545 (I486298,I2859,I97149,I97175,);
DFFARX1 I_5546 (I97175,I2859,I97149,I97192,);
not I_5547 (I97141,I97192);
not I_5548 (I97214,I97175);
DFFARX1 I_5549 (I486298,I2859,I97149,I97240,);
not I_5550 (I97248,I97240);
and I_5551 (I97265,I97214,I486301);
not I_5552 (I97282,I486313);
nand I_5553 (I97299,I97282,I486301);
not I_5554 (I97316,I486319);
nor I_5555 (I97333,I97316,I486310);
nand I_5556 (I97350,I97333,I486316);
nor I_5557 (I97367,I97350,I97299);
DFFARX1 I_5558 (I97367,I2859,I97149,I97117,);
not I_5559 (I97398,I97350);
not I_5560 (I97415,I486310);
nand I_5561 (I97432,I97415,I486301);
nor I_5562 (I97449,I486310,I486313);
nand I_5563 (I97129,I97265,I97449);
nand I_5564 (I97123,I97214,I486310);
nand I_5565 (I97494,I97316,I486307);
DFFARX1 I_5566 (I97494,I2859,I97149,I97138,);
DFFARX1 I_5567 (I97494,I2859,I97149,I97132,);
not I_5568 (I97539,I486307);
nor I_5569 (I97556,I97539,I486304);
and I_5570 (I97573,I97556,I486322);
or I_5571 (I97590,I97573,I486301);
DFFARX1 I_5572 (I97590,I2859,I97149,I97616,);
nand I_5573 (I97624,I97616,I97282);
nor I_5574 (I97126,I97624,I97432);
nor I_5575 (I97120,I97616,I97248);
DFFARX1 I_5576 (I97616,I2859,I97149,I97678,);
not I_5577 (I97686,I97678);
nor I_5578 (I97135,I97686,I97398);
not I_5579 (I97744,I2866);
DFFARX1 I_5580 (I174032,I2859,I97744,I97770,);
DFFARX1 I_5581 (I97770,I2859,I97744,I97787,);
not I_5582 (I97736,I97787);
not I_5583 (I97809,I97770);
DFFARX1 I_5584 (I174020,I2859,I97744,I97835,);
not I_5585 (I97843,I97835);
and I_5586 (I97860,I97809,I174029);
not I_5587 (I97877,I174026);
nand I_5588 (I97894,I97877,I174029);
not I_5589 (I97911,I174017);
nor I_5590 (I97928,I97911,I174023);
nand I_5591 (I97945,I97928,I174008);
nor I_5592 (I97962,I97945,I97894);
DFFARX1 I_5593 (I97962,I2859,I97744,I97712,);
not I_5594 (I97993,I97945);
not I_5595 (I98010,I174023);
nand I_5596 (I98027,I98010,I174029);
nor I_5597 (I98044,I174023,I174026);
nand I_5598 (I97724,I97860,I98044);
nand I_5599 (I97718,I97809,I174023);
nand I_5600 (I98089,I97911,I174008);
DFFARX1 I_5601 (I98089,I2859,I97744,I97733,);
DFFARX1 I_5602 (I98089,I2859,I97744,I97727,);
not I_5603 (I98134,I174008);
nor I_5604 (I98151,I98134,I174014);
and I_5605 (I98168,I98151,I174011);
or I_5606 (I98185,I98168,I174035);
DFFARX1 I_5607 (I98185,I2859,I97744,I98211,);
nand I_5608 (I98219,I98211,I97877);
nor I_5609 (I97721,I98219,I98027);
nor I_5610 (I97715,I98211,I97843);
DFFARX1 I_5611 (I98211,I2859,I97744,I98273,);
not I_5612 (I98281,I98273);
nor I_5613 (I97730,I98281,I97993);
not I_5614 (I98339,I2866);
DFFARX1 I_5615 (I41689,I2859,I98339,I98365,);
DFFARX1 I_5616 (I98365,I2859,I98339,I98382,);
not I_5617 (I98331,I98382);
not I_5618 (I98404,I98365);
DFFARX1 I_5619 (I41683,I2859,I98339,I98430,);
not I_5620 (I98438,I98430);
and I_5621 (I98455,I98404,I41680);
not I_5622 (I98472,I41701);
nand I_5623 (I98489,I98472,I41680);
not I_5624 (I98506,I41695);
nor I_5625 (I98523,I98506,I41686);
nand I_5626 (I98540,I98523,I41692);
nor I_5627 (I98557,I98540,I98489);
DFFARX1 I_5628 (I98557,I2859,I98339,I98307,);
not I_5629 (I98588,I98540);
not I_5630 (I98605,I41686);
nand I_5631 (I98622,I98605,I41680);
nor I_5632 (I98639,I41686,I41701);
nand I_5633 (I98319,I98455,I98639);
nand I_5634 (I98313,I98404,I41686);
nand I_5635 (I98684,I98506,I41680);
DFFARX1 I_5636 (I98684,I2859,I98339,I98328,);
DFFARX1 I_5637 (I98684,I2859,I98339,I98322,);
not I_5638 (I98729,I41680);
nor I_5639 (I98746,I98729,I41698);
and I_5640 (I98763,I98746,I41704);
or I_5641 (I98780,I98763,I41683);
DFFARX1 I_5642 (I98780,I2859,I98339,I98806,);
nand I_5643 (I98814,I98806,I98472);
nor I_5644 (I98316,I98814,I98622);
nor I_5645 (I98310,I98806,I98438);
DFFARX1 I_5646 (I98806,I2859,I98339,I98868,);
not I_5647 (I98876,I98868);
nor I_5648 (I98325,I98876,I98588);
not I_5649 (I98934,I2866);
DFFARX1 I_5650 (I43270,I2859,I98934,I98960,);
DFFARX1 I_5651 (I98960,I2859,I98934,I98977,);
not I_5652 (I98926,I98977);
not I_5653 (I98999,I98960);
DFFARX1 I_5654 (I43264,I2859,I98934,I99025,);
not I_5655 (I99033,I99025);
and I_5656 (I99050,I98999,I43261);
not I_5657 (I99067,I43282);
nand I_5658 (I99084,I99067,I43261);
not I_5659 (I99101,I43276);
nor I_5660 (I99118,I99101,I43267);
nand I_5661 (I99135,I99118,I43273);
nor I_5662 (I99152,I99135,I99084);
DFFARX1 I_5663 (I99152,I2859,I98934,I98902,);
not I_5664 (I99183,I99135);
not I_5665 (I99200,I43267);
nand I_5666 (I99217,I99200,I43261);
nor I_5667 (I99234,I43267,I43282);
nand I_5668 (I98914,I99050,I99234);
nand I_5669 (I98908,I98999,I43267);
nand I_5670 (I99279,I99101,I43261);
DFFARX1 I_5671 (I99279,I2859,I98934,I98923,);
DFFARX1 I_5672 (I99279,I2859,I98934,I98917,);
not I_5673 (I99324,I43261);
nor I_5674 (I99341,I99324,I43279);
and I_5675 (I99358,I99341,I43285);
or I_5676 (I99375,I99358,I43264);
DFFARX1 I_5677 (I99375,I2859,I98934,I99401,);
nand I_5678 (I99409,I99401,I99067);
nor I_5679 (I98911,I99409,I99217);
nor I_5680 (I98905,I99401,I99033);
DFFARX1 I_5681 (I99401,I2859,I98934,I99463,);
not I_5682 (I99471,I99463);
nor I_5683 (I98920,I99471,I99183);
not I_5684 (I99529,I2866);
DFFARX1 I_5685 (I513380,I2859,I99529,I99555,);
DFFARX1 I_5686 (I99555,I2859,I99529,I99572,);
not I_5687 (I99521,I99572);
not I_5688 (I99594,I99555);
DFFARX1 I_5689 (I513365,I2859,I99529,I99620,);
not I_5690 (I99628,I99620);
and I_5691 (I99645,I99594,I513383);
not I_5692 (I99662,I513365);
nand I_5693 (I99679,I99662,I513383);
not I_5694 (I99696,I513386);
nor I_5695 (I99713,I99696,I513377);
nand I_5696 (I99730,I99713,I513374);
nor I_5697 (I99747,I99730,I99679);
DFFARX1 I_5698 (I99747,I2859,I99529,I99497,);
not I_5699 (I99778,I99730);
not I_5700 (I99795,I513377);
nand I_5701 (I99812,I99795,I513383);
nor I_5702 (I99829,I513377,I513365);
nand I_5703 (I99509,I99645,I99829);
nand I_5704 (I99503,I99594,I513377);
nand I_5705 (I99874,I99696,I513371);
DFFARX1 I_5706 (I99874,I2859,I99529,I99518,);
DFFARX1 I_5707 (I99874,I2859,I99529,I99512,);
not I_5708 (I99919,I513371);
nor I_5709 (I99936,I99919,I513362);
and I_5710 (I99953,I99936,I513368);
or I_5711 (I99970,I99953,I513362);
DFFARX1 I_5712 (I99970,I2859,I99529,I99996,);
nand I_5713 (I100004,I99996,I99662);
nor I_5714 (I99506,I100004,I99812);
nor I_5715 (I99500,I99996,I99628);
DFFARX1 I_5716 (I99996,I2859,I99529,I100058,);
not I_5717 (I100066,I100058);
nor I_5718 (I99515,I100066,I99778);
not I_5719 (I100124,I2866);
DFFARX1 I_5720 (I111924,I2859,I100124,I100150,);
DFFARX1 I_5721 (I100150,I2859,I100124,I100167,);
not I_5722 (I100116,I100167);
not I_5723 (I100189,I100150);
DFFARX1 I_5724 (I111939,I2859,I100124,I100215,);
not I_5725 (I100223,I100215);
and I_5726 (I100240,I100189,I111936);
not I_5727 (I100257,I111924);
nand I_5728 (I100274,I100257,I111936);
not I_5729 (I100291,I111933);
nor I_5730 (I100308,I100291,I111948);
nand I_5731 (I100325,I100308,I111945);
nor I_5732 (I100342,I100325,I100274);
DFFARX1 I_5733 (I100342,I2859,I100124,I100092,);
not I_5734 (I100373,I100325);
not I_5735 (I100390,I111948);
nand I_5736 (I100407,I100390,I111936);
nor I_5737 (I100424,I111948,I111924);
nand I_5738 (I100104,I100240,I100424);
nand I_5739 (I100098,I100189,I111948);
nand I_5740 (I100469,I100291,I111942);
DFFARX1 I_5741 (I100469,I2859,I100124,I100113,);
DFFARX1 I_5742 (I100469,I2859,I100124,I100107,);
not I_5743 (I100514,I111942);
nor I_5744 (I100531,I100514,I111930);
and I_5745 (I100548,I100531,I111951);
or I_5746 (I100565,I100548,I111927);
DFFARX1 I_5747 (I100565,I2859,I100124,I100591,);
nand I_5748 (I100599,I100591,I100257);
nor I_5749 (I100101,I100599,I100407);
nor I_5750 (I100095,I100591,I100223);
DFFARX1 I_5751 (I100591,I2859,I100124,I100653,);
not I_5752 (I100661,I100653);
nor I_5753 (I100110,I100661,I100373);
not I_5754 (I100719,I2866);
DFFARX1 I_5755 (I2887,I2859,I100719,I100745,);
DFFARX1 I_5756 (I100745,I2859,I100719,I100762,);
not I_5757 (I100711,I100762);
not I_5758 (I100784,I100745);
DFFARX1 I_5759 (I2884,I2859,I100719,I100810,);
not I_5760 (I100818,I100810);
and I_5761 (I100835,I100784,I2875);
not I_5762 (I100852,I2872);
nand I_5763 (I100869,I100852,I2875);
not I_5764 (I100886,I2872);
nor I_5765 (I100903,I100886,I2869);
nand I_5766 (I100920,I100903,I2881);
nor I_5767 (I100937,I100920,I100869);
DFFARX1 I_5768 (I100937,I2859,I100719,I100687,);
not I_5769 (I100968,I100920);
not I_5770 (I100985,I2869);
nand I_5771 (I101002,I100985,I2875);
nor I_5772 (I101019,I2869,I2872);
nand I_5773 (I100699,I100835,I101019);
nand I_5774 (I100693,I100784,I2869);
nand I_5775 (I101064,I100886,I2878);
DFFARX1 I_5776 (I101064,I2859,I100719,I100708,);
DFFARX1 I_5777 (I101064,I2859,I100719,I100702,);
not I_5778 (I101109,I2878);
nor I_5779 (I101126,I101109,I2890);
and I_5780 (I101143,I101126,I2875);
or I_5781 (I101160,I101143,I2869);
DFFARX1 I_5782 (I101160,I2859,I100719,I101186,);
nand I_5783 (I101194,I101186,I100852);
nor I_5784 (I100696,I101194,I101002);
nor I_5785 (I100690,I101186,I100818);
DFFARX1 I_5786 (I101186,I2859,I100719,I101248,);
not I_5787 (I101256,I101248);
nor I_5788 (I100705,I101256,I100968);
not I_5789 (I101314,I2866);
DFFARX1 I_5790 (I134058,I2859,I101314,I101340,);
DFFARX1 I_5791 (I101340,I2859,I101314,I101357,);
not I_5792 (I101306,I101357);
not I_5793 (I101379,I101340);
DFFARX1 I_5794 (I134073,I2859,I101314,I101405,);
not I_5795 (I101413,I101405);
and I_5796 (I101430,I101379,I134070);
not I_5797 (I101447,I134058);
nand I_5798 (I101464,I101447,I134070);
not I_5799 (I101481,I134067);
nor I_5800 (I101498,I101481,I134082);
nand I_5801 (I101515,I101498,I134079);
nor I_5802 (I101532,I101515,I101464);
DFFARX1 I_5803 (I101532,I2859,I101314,I101282,);
not I_5804 (I101563,I101515);
not I_5805 (I101580,I134082);
nand I_5806 (I101597,I101580,I134070);
nor I_5807 (I101614,I134082,I134058);
nand I_5808 (I101294,I101430,I101614);
nand I_5809 (I101288,I101379,I134082);
nand I_5810 (I101659,I101481,I134076);
DFFARX1 I_5811 (I101659,I2859,I101314,I101303,);
DFFARX1 I_5812 (I101659,I2859,I101314,I101297,);
not I_5813 (I101704,I134076);
nor I_5814 (I101721,I101704,I134064);
and I_5815 (I101738,I101721,I134085);
or I_5816 (I101755,I101738,I134061);
DFFARX1 I_5817 (I101755,I2859,I101314,I101781,);
nand I_5818 (I101789,I101781,I101447);
nor I_5819 (I101291,I101789,I101597);
nor I_5820 (I101285,I101781,I101413);
DFFARX1 I_5821 (I101781,I2859,I101314,I101843,);
not I_5822 (I101851,I101843);
nor I_5823 (I101300,I101851,I101563);
not I_5824 (I101909,I2866);
DFFARX1 I_5825 (I493234,I2859,I101909,I101935,);
DFFARX1 I_5826 (I101935,I2859,I101909,I101952,);
not I_5827 (I101901,I101952);
not I_5828 (I101974,I101935);
DFFARX1 I_5829 (I493234,I2859,I101909,I102000,);
not I_5830 (I102008,I102000);
and I_5831 (I102025,I101974,I493237);
not I_5832 (I102042,I493249);
nand I_5833 (I102059,I102042,I493237);
not I_5834 (I102076,I493255);
nor I_5835 (I102093,I102076,I493246);
nand I_5836 (I102110,I102093,I493252);
nor I_5837 (I102127,I102110,I102059);
DFFARX1 I_5838 (I102127,I2859,I101909,I101877,);
not I_5839 (I102158,I102110);
not I_5840 (I102175,I493246);
nand I_5841 (I102192,I102175,I493237);
nor I_5842 (I102209,I493246,I493249);
nand I_5843 (I101889,I102025,I102209);
nand I_5844 (I101883,I101974,I493246);
nand I_5845 (I102254,I102076,I493243);
DFFARX1 I_5846 (I102254,I2859,I101909,I101898,);
DFFARX1 I_5847 (I102254,I2859,I101909,I101892,);
not I_5848 (I102299,I493243);
nor I_5849 (I102316,I102299,I493240);
and I_5850 (I102333,I102316,I493258);
or I_5851 (I102350,I102333,I493237);
DFFARX1 I_5852 (I102350,I2859,I101909,I102376,);
nand I_5853 (I102384,I102376,I102042);
nor I_5854 (I101886,I102384,I102192);
nor I_5855 (I101880,I102376,I102008);
DFFARX1 I_5856 (I102376,I2859,I101909,I102438,);
not I_5857 (I102446,I102438);
nor I_5858 (I101895,I102446,I102158);
not I_5859 (I102504,I2866);
DFFARX1 I_5860 (I494390,I2859,I102504,I102530,);
DFFARX1 I_5861 (I102530,I2859,I102504,I102547,);
not I_5862 (I102496,I102547);
not I_5863 (I102569,I102530);
DFFARX1 I_5864 (I494390,I2859,I102504,I102595,);
not I_5865 (I102603,I102595);
and I_5866 (I102620,I102569,I494393);
not I_5867 (I102637,I494405);
nand I_5868 (I102654,I102637,I494393);
not I_5869 (I102671,I494411);
nor I_5870 (I102688,I102671,I494402);
nand I_5871 (I102705,I102688,I494408);
nor I_5872 (I102722,I102705,I102654);
DFFARX1 I_5873 (I102722,I2859,I102504,I102472,);
not I_5874 (I102753,I102705);
not I_5875 (I102770,I494402);
nand I_5876 (I102787,I102770,I494393);
nor I_5877 (I102804,I494402,I494405);
nand I_5878 (I102484,I102620,I102804);
nand I_5879 (I102478,I102569,I494402);
nand I_5880 (I102849,I102671,I494399);
DFFARX1 I_5881 (I102849,I2859,I102504,I102493,);
DFFARX1 I_5882 (I102849,I2859,I102504,I102487,);
not I_5883 (I102894,I494399);
nor I_5884 (I102911,I102894,I494396);
and I_5885 (I102928,I102911,I494414);
or I_5886 (I102945,I102928,I494393);
DFFARX1 I_5887 (I102945,I2859,I102504,I102971,);
nand I_5888 (I102979,I102971,I102637);
nor I_5889 (I102481,I102979,I102787);
nor I_5890 (I102475,I102971,I102603);
DFFARX1 I_5891 (I102971,I2859,I102504,I103033,);
not I_5892 (I103041,I103033);
nor I_5893 (I102490,I103041,I102753);
not I_5894 (I103099,I2866);
DFFARX1 I_5895 (I516100,I2859,I103099,I103125,);
DFFARX1 I_5896 (I103125,I2859,I103099,I103142,);
not I_5897 (I103091,I103142);
not I_5898 (I103164,I103125);
DFFARX1 I_5899 (I516085,I2859,I103099,I103190,);
not I_5900 (I103198,I103190);
and I_5901 (I103215,I103164,I516103);
not I_5902 (I103232,I516085);
nand I_5903 (I103249,I103232,I516103);
not I_5904 (I103266,I516106);
nor I_5905 (I103283,I103266,I516097);
nand I_5906 (I103300,I103283,I516094);
nor I_5907 (I103317,I103300,I103249);
DFFARX1 I_5908 (I103317,I2859,I103099,I103067,);
not I_5909 (I103348,I103300);
not I_5910 (I103365,I516097);
nand I_5911 (I103382,I103365,I516103);
nor I_5912 (I103399,I516097,I516085);
nand I_5913 (I103079,I103215,I103399);
nand I_5914 (I103073,I103164,I516097);
nand I_5915 (I103444,I103266,I516091);
DFFARX1 I_5916 (I103444,I2859,I103099,I103088,);
DFFARX1 I_5917 (I103444,I2859,I103099,I103082,);
not I_5918 (I103489,I516091);
nor I_5919 (I103506,I103489,I516082);
and I_5920 (I103523,I103506,I516088);
or I_5921 (I103540,I103523,I516082);
DFFARX1 I_5922 (I103540,I2859,I103099,I103566,);
nand I_5923 (I103574,I103566,I103232);
nor I_5924 (I103076,I103574,I103382);
nor I_5925 (I103070,I103566,I103198);
DFFARX1 I_5926 (I103566,I2859,I103099,I103628,);
not I_5927 (I103636,I103628);
nor I_5928 (I103085,I103636,I103348);
not I_5929 (I103694,I2866);
DFFARX1 I_5930 (I407042,I2859,I103694,I103720,);
DFFARX1 I_5931 (I103720,I2859,I103694,I103737,);
not I_5932 (I103686,I103737);
not I_5933 (I103759,I103720);
DFFARX1 I_5934 (I407051,I2859,I103694,I103785,);
not I_5935 (I103793,I103785);
and I_5936 (I103810,I103759,I407039);
not I_5937 (I103827,I407030);
nand I_5938 (I103844,I103827,I407039);
not I_5939 (I103861,I407036);
nor I_5940 (I103878,I103861,I407054);
nand I_5941 (I103895,I103878,I407027);
nor I_5942 (I103912,I103895,I103844);
DFFARX1 I_5943 (I103912,I2859,I103694,I103662,);
not I_5944 (I103943,I103895);
not I_5945 (I103960,I407054);
nand I_5946 (I103977,I103960,I407039);
nor I_5947 (I103994,I407054,I407030);
nand I_5948 (I103674,I103810,I103994);
nand I_5949 (I103668,I103759,I407054);
nand I_5950 (I104039,I103861,I407033);
DFFARX1 I_5951 (I104039,I2859,I103694,I103683,);
DFFARX1 I_5952 (I104039,I2859,I103694,I103677,);
not I_5953 (I104084,I407033);
nor I_5954 (I104101,I104084,I407045);
and I_5955 (I104118,I104101,I407027);
or I_5956 (I104135,I104118,I407048);
DFFARX1 I_5957 (I104135,I2859,I103694,I104161,);
nand I_5958 (I104169,I104161,I103827);
nor I_5959 (I103671,I104169,I103977);
nor I_5960 (I103665,I104161,I103793);
DFFARX1 I_5961 (I104161,I2859,I103694,I104223,);
not I_5962 (I104231,I104223);
nor I_5963 (I103680,I104231,I103943);
not I_5964 (I104289,I2866);
DFFARX1 I_5965 (I167504,I2859,I104289,I104315,);
DFFARX1 I_5966 (I104315,I2859,I104289,I104332,);
not I_5967 (I104281,I104332);
not I_5968 (I104354,I104315);
DFFARX1 I_5969 (I167492,I2859,I104289,I104380,);
not I_5970 (I104388,I104380);
and I_5971 (I104405,I104354,I167501);
not I_5972 (I104422,I167498);
nand I_5973 (I104439,I104422,I167501);
not I_5974 (I104456,I167489);
nor I_5975 (I104473,I104456,I167495);
nand I_5976 (I104490,I104473,I167480);
nor I_5977 (I104507,I104490,I104439);
DFFARX1 I_5978 (I104507,I2859,I104289,I104257,);
not I_5979 (I104538,I104490);
not I_5980 (I104555,I167495);
nand I_5981 (I104572,I104555,I167501);
nor I_5982 (I104589,I167495,I167498);
nand I_5983 (I104269,I104405,I104589);
nand I_5984 (I104263,I104354,I167495);
nand I_5985 (I104634,I104456,I167480);
DFFARX1 I_5986 (I104634,I2859,I104289,I104278,);
DFFARX1 I_5987 (I104634,I2859,I104289,I104272,);
not I_5988 (I104679,I167480);
nor I_5989 (I104696,I104679,I167486);
and I_5990 (I104713,I104696,I167483);
or I_5991 (I104730,I104713,I167507);
DFFARX1 I_5992 (I104730,I2859,I104289,I104756,);
nand I_5993 (I104764,I104756,I104422);
nor I_5994 (I104266,I104764,I104572);
nor I_5995 (I104260,I104756,I104388);
DFFARX1 I_5996 (I104756,I2859,I104289,I104818,);
not I_5997 (I104826,I104818);
nor I_5998 (I104275,I104826,I104538);
not I_5999 (I104884,I2866);
DFFARX1 I_6000 (I448728,I2859,I104884,I104910,);
DFFARX1 I_6001 (I104910,I2859,I104884,I104927,);
not I_6002 (I104876,I104927);
not I_6003 (I104949,I104910);
DFFARX1 I_6004 (I448728,I2859,I104884,I104975,);
not I_6005 (I104983,I104975);
and I_6006 (I105000,I104949,I448731);
not I_6007 (I105017,I448743);
nand I_6008 (I105034,I105017,I448731);
not I_6009 (I105051,I448749);
nor I_6010 (I105068,I105051,I448740);
nand I_6011 (I105085,I105068,I448746);
nor I_6012 (I105102,I105085,I105034);
DFFARX1 I_6013 (I105102,I2859,I104884,I104852,);
not I_6014 (I105133,I105085);
not I_6015 (I105150,I448740);
nand I_6016 (I105167,I105150,I448731);
nor I_6017 (I105184,I448740,I448743);
nand I_6018 (I104864,I105000,I105184);
nand I_6019 (I104858,I104949,I448740);
nand I_6020 (I105229,I105051,I448737);
DFFARX1 I_6021 (I105229,I2859,I104884,I104873,);
DFFARX1 I_6022 (I105229,I2859,I104884,I104867,);
not I_6023 (I105274,I448737);
nor I_6024 (I105291,I105274,I448734);
and I_6025 (I105308,I105291,I448752);
or I_6026 (I105325,I105308,I448731);
DFFARX1 I_6027 (I105325,I2859,I104884,I105351,);
nand I_6028 (I105359,I105351,I105017);
nor I_6029 (I104861,I105359,I105167);
nor I_6030 (I104855,I105351,I104983);
DFFARX1 I_6031 (I105351,I2859,I104884,I105413,);
not I_6032 (I105421,I105413);
nor I_6033 (I104870,I105421,I105133);
not I_6034 (I105479,I2866);
DFFARX1 I_6035 (I339679,I2859,I105479,I105505,);
DFFARX1 I_6036 (I105505,I2859,I105479,I105522,);
not I_6037 (I105471,I105522);
not I_6038 (I105544,I105505);
DFFARX1 I_6039 (I339673,I2859,I105479,I105570,);
not I_6040 (I105578,I105570);
and I_6041 (I105595,I105544,I339691);
not I_6042 (I105612,I339679);
nand I_6043 (I105629,I105612,I339691);
not I_6044 (I105646,I339673);
nor I_6045 (I105663,I105646,I339685);
nand I_6046 (I105680,I105663,I339676);
nor I_6047 (I105697,I105680,I105629);
DFFARX1 I_6048 (I105697,I2859,I105479,I105447,);
not I_6049 (I105728,I105680);
not I_6050 (I105745,I339685);
nand I_6051 (I105762,I105745,I339691);
nor I_6052 (I105779,I339685,I339679);
nand I_6053 (I105459,I105595,I105779);
nand I_6054 (I105453,I105544,I339685);
nand I_6055 (I105824,I105646,I339688);
DFFARX1 I_6056 (I105824,I2859,I105479,I105468,);
DFFARX1 I_6057 (I105824,I2859,I105479,I105462,);
not I_6058 (I105869,I339688);
nor I_6059 (I105886,I105869,I339694);
and I_6060 (I105903,I105886,I339676);
or I_6061 (I105920,I105903,I339682);
DFFARX1 I_6062 (I105920,I2859,I105479,I105946,);
nand I_6063 (I105954,I105946,I105612);
nor I_6064 (I105456,I105954,I105762);
nor I_6065 (I105450,I105946,I105578);
DFFARX1 I_6066 (I105946,I2859,I105479,I106008,);
not I_6067 (I106016,I106008);
nor I_6068 (I105465,I106016,I105728);
not I_6069 (I106074,I2866);
DFFARX1 I_6070 (I282242,I2859,I106074,I106100,);
DFFARX1 I_6071 (I106100,I2859,I106074,I106117,);
not I_6072 (I106066,I106117);
not I_6073 (I106139,I106100);
DFFARX1 I_6074 (I282239,I2859,I106074,I106165,);
not I_6075 (I106173,I106165);
and I_6076 (I106190,I106139,I282245);
not I_6077 (I106207,I282230);
nand I_6078 (I106224,I106207,I282245);
not I_6079 (I106241,I282233);
nor I_6080 (I106258,I106241,I282254);
nand I_6081 (I106275,I106258,I282251);
nor I_6082 (I106292,I106275,I106224);
DFFARX1 I_6083 (I106292,I2859,I106074,I106042,);
not I_6084 (I106323,I106275);
not I_6085 (I106340,I282254);
nand I_6086 (I106357,I106340,I282245);
nor I_6087 (I106374,I282254,I282230);
nand I_6088 (I106054,I106190,I106374);
nand I_6089 (I106048,I106139,I282254);
nand I_6090 (I106419,I106241,I282230);
DFFARX1 I_6091 (I106419,I2859,I106074,I106063,);
DFFARX1 I_6092 (I106419,I2859,I106074,I106057,);
not I_6093 (I106464,I282230);
nor I_6094 (I106481,I106464,I282236);
and I_6095 (I106498,I106481,I282248);
or I_6096 (I106515,I106498,I282233);
DFFARX1 I_6097 (I106515,I2859,I106074,I106541,);
nand I_6098 (I106549,I106541,I106207);
nor I_6099 (I106051,I106549,I106357);
nor I_6100 (I106045,I106541,I106173);
DFFARX1 I_6101 (I106541,I2859,I106074,I106603,);
not I_6102 (I106611,I106603);
nor I_6103 (I106060,I106611,I106323);
not I_6104 (I106669,I2866);
DFFARX1 I_6105 (I315188,I2859,I106669,I106695,);
DFFARX1 I_6106 (I106695,I2859,I106669,I106712,);
not I_6107 (I106661,I106712);
not I_6108 (I106734,I106695);
DFFARX1 I_6109 (I315185,I2859,I106669,I106760,);
not I_6110 (I106768,I106760);
and I_6111 (I106785,I106734,I315191);
not I_6112 (I106802,I315176);
nand I_6113 (I106819,I106802,I315191);
not I_6114 (I106836,I315179);
nor I_6115 (I106853,I106836,I315200);
nand I_6116 (I106870,I106853,I315197);
nor I_6117 (I106887,I106870,I106819);
DFFARX1 I_6118 (I106887,I2859,I106669,I106637,);
not I_6119 (I106918,I106870);
not I_6120 (I106935,I315200);
nand I_6121 (I106952,I106935,I315191);
nor I_6122 (I106969,I315200,I315176);
nand I_6123 (I106649,I106785,I106969);
nand I_6124 (I106643,I106734,I315200);
nand I_6125 (I107014,I106836,I315176);
DFFARX1 I_6126 (I107014,I2859,I106669,I106658,);
DFFARX1 I_6127 (I107014,I2859,I106669,I106652,);
not I_6128 (I107059,I315176);
nor I_6129 (I107076,I107059,I315182);
and I_6130 (I107093,I107076,I315194);
or I_6131 (I107110,I107093,I315179);
DFFARX1 I_6132 (I107110,I2859,I106669,I107136,);
nand I_6133 (I107144,I107136,I106802);
nor I_6134 (I106646,I107144,I106952);
nor I_6135 (I106640,I107136,I106768);
DFFARX1 I_6136 (I107136,I2859,I106669,I107198,);
not I_6137 (I107206,I107198);
nor I_6138 (I106655,I107206,I106918);
not I_6139 (I107264,I2866);
DFFARX1 I_6140 (I279930,I2859,I107264,I107290,);
DFFARX1 I_6141 (I107290,I2859,I107264,I107307,);
not I_6142 (I107256,I107307);
not I_6143 (I107329,I107290);
DFFARX1 I_6144 (I279927,I2859,I107264,I107355,);
not I_6145 (I107363,I107355);
and I_6146 (I107380,I107329,I279933);
not I_6147 (I107397,I279918);
nand I_6148 (I107414,I107397,I279933);
not I_6149 (I107431,I279921);
nor I_6150 (I107448,I107431,I279942);
nand I_6151 (I107465,I107448,I279939);
nor I_6152 (I107482,I107465,I107414);
DFFARX1 I_6153 (I107482,I2859,I107264,I107232,);
not I_6154 (I107513,I107465);
not I_6155 (I107530,I279942);
nand I_6156 (I107547,I107530,I279933);
nor I_6157 (I107564,I279942,I279918);
nand I_6158 (I107244,I107380,I107564);
nand I_6159 (I107238,I107329,I279942);
nand I_6160 (I107609,I107431,I279918);
DFFARX1 I_6161 (I107609,I2859,I107264,I107253,);
DFFARX1 I_6162 (I107609,I2859,I107264,I107247,);
not I_6163 (I107654,I279918);
nor I_6164 (I107671,I107654,I279924);
and I_6165 (I107688,I107671,I279936);
or I_6166 (I107705,I107688,I279921);
DFFARX1 I_6167 (I107705,I2859,I107264,I107731,);
nand I_6168 (I107739,I107731,I107397);
nor I_6169 (I107241,I107739,I107547);
nor I_6170 (I107235,I107731,I107363);
DFFARX1 I_6171 (I107731,I2859,I107264,I107793,);
not I_6172 (I107801,I107793);
nor I_6173 (I107250,I107801,I107513);
not I_6174 (I107859,I2866);
DFFARX1 I_6175 (I173488,I2859,I107859,I107885,);
DFFARX1 I_6176 (I107885,I2859,I107859,I107902,);
not I_6177 (I107851,I107902);
not I_6178 (I107924,I107885);
DFFARX1 I_6179 (I173476,I2859,I107859,I107950,);
not I_6180 (I107958,I107950);
and I_6181 (I107975,I107924,I173485);
not I_6182 (I107992,I173482);
nand I_6183 (I108009,I107992,I173485);
not I_6184 (I108026,I173473);
nor I_6185 (I108043,I108026,I173479);
nand I_6186 (I108060,I108043,I173464);
nor I_6187 (I108077,I108060,I108009);
DFFARX1 I_6188 (I108077,I2859,I107859,I107827,);
not I_6189 (I108108,I108060);
not I_6190 (I108125,I173479);
nand I_6191 (I108142,I108125,I173485);
nor I_6192 (I108159,I173479,I173482);
nand I_6193 (I107839,I107975,I108159);
nand I_6194 (I107833,I107924,I173479);
nand I_6195 (I108204,I108026,I173464);
DFFARX1 I_6196 (I108204,I2859,I107859,I107848,);
DFFARX1 I_6197 (I108204,I2859,I107859,I107842,);
not I_6198 (I108249,I173464);
nor I_6199 (I108266,I108249,I173470);
and I_6200 (I108283,I108266,I173467);
or I_6201 (I108300,I108283,I173491);
DFFARX1 I_6202 (I108300,I2859,I107859,I108326,);
nand I_6203 (I108334,I108326,I107992);
nor I_6204 (I107836,I108334,I108142);
nor I_6205 (I107830,I108326,I107958);
DFFARX1 I_6206 (I108326,I2859,I107859,I108388,);
not I_6207 (I108396,I108388);
nor I_6208 (I107845,I108396,I108108);
not I_6209 (I108454,I2866);
DFFARX1 I_6210 (I432173,I2859,I108454,I108480,);
DFFARX1 I_6211 (I108480,I2859,I108454,I108497,);
not I_6212 (I108446,I108497);
not I_6213 (I108519,I108480);
DFFARX1 I_6214 (I432182,I2859,I108454,I108545,);
not I_6215 (I108553,I108545);
and I_6216 (I108570,I108519,I432176);
not I_6217 (I108587,I432170);
nand I_6218 (I108604,I108587,I432176);
not I_6219 (I108621,I432185);
nor I_6220 (I108638,I108621,I432173);
nand I_6221 (I108655,I108638,I432179);
nor I_6222 (I108672,I108655,I108604);
DFFARX1 I_6223 (I108672,I2859,I108454,I108422,);
not I_6224 (I108703,I108655);
not I_6225 (I108720,I432173);
nand I_6226 (I108737,I108720,I432176);
nor I_6227 (I108754,I432173,I432170);
nand I_6228 (I108434,I108570,I108754);
nand I_6229 (I108428,I108519,I432173);
nand I_6230 (I108799,I108621,I432176);
DFFARX1 I_6231 (I108799,I2859,I108454,I108443,);
DFFARX1 I_6232 (I108799,I2859,I108454,I108437,);
not I_6233 (I108844,I432176);
nor I_6234 (I108861,I108844,I432191);
and I_6235 (I108878,I108861,I432188);
or I_6236 (I108895,I108878,I432170);
DFFARX1 I_6237 (I108895,I2859,I108454,I108921,);
nand I_6238 (I108929,I108921,I108587);
nor I_6239 (I108431,I108929,I108737);
nor I_6240 (I108425,I108921,I108553);
DFFARX1 I_6241 (I108921,I2859,I108454,I108983,);
not I_6242 (I108991,I108983);
nor I_6243 (I108440,I108991,I108703);
not I_6244 (I109049,I2866);
DFFARX1 I_6245 (I548131,I2859,I109049,I109075,);
DFFARX1 I_6246 (I109075,I2859,I109049,I109092,);
not I_6247 (I109041,I109092);
not I_6248 (I109114,I109075);
DFFARX1 I_6249 (I548122,I2859,I109049,I109140,);
not I_6250 (I109148,I109140);
and I_6251 (I109165,I109114,I548116);
not I_6252 (I109182,I548110);
nand I_6253 (I109199,I109182,I548116);
not I_6254 (I109216,I548137);
nor I_6255 (I109233,I109216,I548110);
nand I_6256 (I109250,I109233,I548134);
nor I_6257 (I109267,I109250,I109199);
DFFARX1 I_6258 (I109267,I2859,I109049,I109017,);
not I_6259 (I109298,I109250);
not I_6260 (I109315,I548110);
nand I_6261 (I109332,I109315,I548116);
nor I_6262 (I109349,I548110,I548110);
nand I_6263 (I109029,I109165,I109349);
nand I_6264 (I109023,I109114,I548110);
nand I_6265 (I109394,I109216,I548119);
DFFARX1 I_6266 (I109394,I2859,I109049,I109038,);
DFFARX1 I_6267 (I109394,I2859,I109049,I109032,);
not I_6268 (I109439,I548119);
nor I_6269 (I109456,I109439,I548125);
and I_6270 (I109473,I109456,I548128);
or I_6271 (I109490,I109473,I548113);
DFFARX1 I_6272 (I109490,I2859,I109049,I109516,);
nand I_6273 (I109524,I109516,I109182);
nor I_6274 (I109026,I109524,I109332);
nor I_6275 (I109020,I109516,I109148);
DFFARX1 I_6276 (I109516,I2859,I109049,I109578,);
not I_6277 (I109586,I109578);
nor I_6278 (I109035,I109586,I109298);
not I_6279 (I109644,I2866);
DFFARX1 I_6280 (I398644,I2859,I109644,I109670,);
DFFARX1 I_6281 (I109670,I2859,I109644,I109687,);
not I_6282 (I109636,I109687);
not I_6283 (I109709,I109670);
DFFARX1 I_6284 (I398653,I2859,I109644,I109735,);
not I_6285 (I109743,I109735);
and I_6286 (I109760,I109709,I398641);
not I_6287 (I109777,I398632);
nand I_6288 (I109794,I109777,I398641);
not I_6289 (I109811,I398638);
nor I_6290 (I109828,I109811,I398656);
nand I_6291 (I109845,I109828,I398629);
nor I_6292 (I109862,I109845,I109794);
DFFARX1 I_6293 (I109862,I2859,I109644,I109612,);
not I_6294 (I109893,I109845);
not I_6295 (I109910,I398656);
nand I_6296 (I109927,I109910,I398641);
nor I_6297 (I109944,I398656,I398632);
nand I_6298 (I109624,I109760,I109944);
nand I_6299 (I109618,I109709,I398656);
nand I_6300 (I109989,I109811,I398635);
DFFARX1 I_6301 (I109989,I2859,I109644,I109633,);
DFFARX1 I_6302 (I109989,I2859,I109644,I109627,);
not I_6303 (I110034,I398635);
nor I_6304 (I110051,I110034,I398647);
and I_6305 (I110068,I110051,I398629);
or I_6306 (I110085,I110068,I398650);
DFFARX1 I_6307 (I110085,I2859,I109644,I110111,);
nand I_6308 (I110119,I110111,I109777);
nor I_6309 (I109621,I110119,I109927);
nor I_6310 (I109615,I110111,I109743);
DFFARX1 I_6311 (I110111,I2859,I109644,I110173,);
not I_6312 (I110181,I110173);
nor I_6313 (I109630,I110181,I109893);
not I_6314 (I110239,I2866);
DFFARX1 I_6315 (I234271,I2859,I110239,I110265,);
DFFARX1 I_6316 (I110265,I2859,I110239,I110282,);
not I_6317 (I110231,I110282);
not I_6318 (I110304,I110265);
DFFARX1 I_6319 (I234262,I2859,I110239,I110330,);
not I_6320 (I110338,I110330);
and I_6321 (I110355,I110304,I234280);
not I_6322 (I110372,I234277);
nand I_6323 (I110389,I110372,I234280);
not I_6324 (I110406,I234256);
nor I_6325 (I110423,I110406,I234259);
nand I_6326 (I110440,I110423,I234268);
nor I_6327 (I110457,I110440,I110389);
DFFARX1 I_6328 (I110457,I2859,I110239,I110207,);
not I_6329 (I110488,I110440);
not I_6330 (I110505,I234259);
nand I_6331 (I110522,I110505,I234280);
nor I_6332 (I110539,I234259,I234277);
nand I_6333 (I110219,I110355,I110539);
nand I_6334 (I110213,I110304,I234259);
nand I_6335 (I110584,I110406,I234274);
DFFARX1 I_6336 (I110584,I2859,I110239,I110228,);
DFFARX1 I_6337 (I110584,I2859,I110239,I110222,);
not I_6338 (I110629,I234274);
nor I_6339 (I110646,I110629,I234256);
and I_6340 (I110663,I110646,I234265);
or I_6341 (I110680,I110663,I234259);
DFFARX1 I_6342 (I110680,I2859,I110239,I110706,);
nand I_6343 (I110714,I110706,I110372);
nor I_6344 (I110216,I110714,I110522);
nor I_6345 (I110210,I110706,I110338);
DFFARX1 I_6346 (I110706,I2859,I110239,I110768,);
not I_6347 (I110776,I110768);
nor I_6348 (I110225,I110776,I110488);
not I_6349 (I110834,I2866);
DFFARX1 I_6350 (I168592,I2859,I110834,I110860,);
DFFARX1 I_6351 (I110860,I2859,I110834,I110877,);
not I_6352 (I110826,I110877);
not I_6353 (I110899,I110860);
DFFARX1 I_6354 (I168580,I2859,I110834,I110925,);
not I_6355 (I110933,I110925);
and I_6356 (I110950,I110899,I168589);
not I_6357 (I110967,I168586);
nand I_6358 (I110984,I110967,I168589);
not I_6359 (I111001,I168577);
nor I_6360 (I111018,I111001,I168583);
nand I_6361 (I111035,I111018,I168568);
nor I_6362 (I111052,I111035,I110984);
DFFARX1 I_6363 (I111052,I2859,I110834,I110802,);
not I_6364 (I111083,I111035);
not I_6365 (I111100,I168583);
nand I_6366 (I111117,I111100,I168589);
nor I_6367 (I111134,I168583,I168586);
nand I_6368 (I110814,I110950,I111134);
nand I_6369 (I110808,I110899,I168583);
nand I_6370 (I111179,I111001,I168568);
DFFARX1 I_6371 (I111179,I2859,I110834,I110823,);
DFFARX1 I_6372 (I111179,I2859,I110834,I110817,);
not I_6373 (I111224,I168568);
nor I_6374 (I111241,I111224,I168574);
and I_6375 (I111258,I111241,I168571);
or I_6376 (I111275,I111258,I168595);
DFFARX1 I_6377 (I111275,I2859,I110834,I111301,);
nand I_6378 (I111309,I111301,I110967);
nor I_6379 (I110811,I111309,I111117);
nor I_6380 (I110805,I111301,I110933);
DFFARX1 I_6381 (I111301,I2859,I110834,I111363,);
not I_6382 (I111371,I111363);
nor I_6383 (I110820,I111371,I111083);
not I_6384 (I111432,I2866);
DFFARX1 I_6385 (I265480,I2859,I111432,I111458,);
nand I_6386 (I111466,I265471,I265486);
and I_6387 (I111483,I111466,I265492);
DFFARX1 I_6388 (I111483,I2859,I111432,I111509,);
nor I_6389 (I111400,I111509,I111458);
not I_6390 (I111531,I111509);
DFFARX1 I_6391 (I265477,I2859,I111432,I111557,);
nand I_6392 (I111565,I111557,I265471);
not I_6393 (I111582,I111565);
DFFARX1 I_6394 (I111582,I2859,I111432,I111608,);
not I_6395 (I111424,I111608);
nor I_6396 (I111630,I111458,I111565);
nor I_6397 (I111406,I111509,I111630);
DFFARX1 I_6398 (I265474,I2859,I111432,I111670,);
DFFARX1 I_6399 (I111670,I2859,I111432,I111687,);
not I_6400 (I111695,I111687);
not I_6401 (I111712,I111670);
nand I_6402 (I111409,I111712,I111531);
nand I_6403 (I111743,I265468,I265483);
and I_6404 (I111760,I111743,I265468);
DFFARX1 I_6405 (I111760,I2859,I111432,I111786,);
nor I_6406 (I111794,I111786,I111458);
DFFARX1 I_6407 (I111794,I2859,I111432,I111397,);
DFFARX1 I_6408 (I111786,I2859,I111432,I111415,);
nor I_6409 (I111839,I265489,I265483);
not I_6410 (I111856,I111839);
nor I_6411 (I111418,I111695,I111856);
nand I_6412 (I111403,I111712,I111856);
nor I_6413 (I111412,I111458,I111839);
DFFARX1 I_6414 (I111839,I2859,I111432,I111421,);
not I_6415 (I111959,I2866);
DFFARX1 I_6416 (I217378,I2859,I111959,I111985,);
nand I_6417 (I111993,I217378,I217390);
and I_6418 (I112010,I111993,I217375);
DFFARX1 I_6419 (I112010,I2859,I111959,I112036,);
nor I_6420 (I111927,I112036,I111985);
not I_6421 (I112058,I112036);
DFFARX1 I_6422 (I217399,I2859,I111959,I112084,);
nand I_6423 (I112092,I112084,I217396);
not I_6424 (I112109,I112092);
DFFARX1 I_6425 (I112109,I2859,I111959,I112135,);
not I_6426 (I111951,I112135);
nor I_6427 (I112157,I111985,I112092);
nor I_6428 (I111933,I112036,I112157);
DFFARX1 I_6429 (I217387,I2859,I111959,I112197,);
DFFARX1 I_6430 (I112197,I2859,I111959,I112214,);
not I_6431 (I112222,I112214);
not I_6432 (I112239,I112197);
nand I_6433 (I111936,I112239,I112058);
nand I_6434 (I112270,I217375,I217384);
and I_6435 (I112287,I112270,I217393);
DFFARX1 I_6436 (I112287,I2859,I111959,I112313,);
nor I_6437 (I112321,I112313,I111985);
DFFARX1 I_6438 (I112321,I2859,I111959,I111924,);
DFFARX1 I_6439 (I112313,I2859,I111959,I111942,);
nor I_6440 (I112366,I217381,I217384);
not I_6441 (I112383,I112366);
nor I_6442 (I111945,I112222,I112383);
nand I_6443 (I111930,I112239,I112383);
nor I_6444 (I111939,I111985,I112366);
DFFARX1 I_6445 (I112366,I2859,I111959,I111948,);
not I_6446 (I112486,I2866);
DFFARX1 I_6447 (I426563,I2859,I112486,I112512,);
nand I_6448 (I112520,I426560,I426563);
and I_6449 (I112537,I112520,I426572);
DFFARX1 I_6450 (I112537,I2859,I112486,I112563,);
nor I_6451 (I112454,I112563,I112512);
not I_6452 (I112585,I112563);
DFFARX1 I_6453 (I426560,I2859,I112486,I112611,);
nand I_6454 (I112619,I112611,I426578);
not I_6455 (I112636,I112619);
DFFARX1 I_6456 (I112636,I2859,I112486,I112662,);
not I_6457 (I112478,I112662);
nor I_6458 (I112684,I112512,I112619);
nor I_6459 (I112460,I112563,I112684);
DFFARX1 I_6460 (I426566,I2859,I112486,I112724,);
DFFARX1 I_6461 (I112724,I2859,I112486,I112741,);
not I_6462 (I112749,I112741);
not I_6463 (I112766,I112724);
nand I_6464 (I112463,I112766,I112585);
nand I_6465 (I112797,I426575,I426581);
and I_6466 (I112814,I112797,I426566);
DFFARX1 I_6467 (I112814,I2859,I112486,I112840,);
nor I_6468 (I112848,I112840,I112512);
DFFARX1 I_6469 (I112848,I2859,I112486,I112451,);
DFFARX1 I_6470 (I112840,I2859,I112486,I112469,);
nor I_6471 (I112893,I426569,I426581);
not I_6472 (I112910,I112893);
nor I_6473 (I112472,I112749,I112910);
nand I_6474 (I112457,I112766,I112910);
nor I_6475 (I112466,I112512,I112893);
DFFARX1 I_6476 (I112893,I2859,I112486,I112475,);
not I_6477 (I113013,I2866);
DFFARX1 I_6478 (I21130,I2859,I113013,I113039,);
nand I_6479 (I113047,I21142,I21151);
and I_6480 (I113064,I113047,I21130);
DFFARX1 I_6481 (I113064,I2859,I113013,I113090,);
nor I_6482 (I112981,I113090,I113039);
not I_6483 (I113112,I113090);
DFFARX1 I_6484 (I21145,I2859,I113013,I113138,);
nand I_6485 (I113146,I113138,I21133);
not I_6486 (I113163,I113146);
DFFARX1 I_6487 (I113163,I2859,I113013,I113189,);
not I_6488 (I113005,I113189);
nor I_6489 (I113211,I113039,I113146);
nor I_6490 (I112987,I113090,I113211);
DFFARX1 I_6491 (I21136,I2859,I113013,I113251,);
DFFARX1 I_6492 (I113251,I2859,I113013,I113268,);
not I_6493 (I113276,I113268);
not I_6494 (I113293,I113251);
nand I_6495 (I112990,I113293,I113112);
nand I_6496 (I113324,I21127,I21127);
and I_6497 (I113341,I113324,I21139);
DFFARX1 I_6498 (I113341,I2859,I113013,I113367,);
nor I_6499 (I113375,I113367,I113039);
DFFARX1 I_6500 (I113375,I2859,I113013,I112978,);
DFFARX1 I_6501 (I113367,I2859,I113013,I112996,);
nor I_6502 (I113420,I21148,I21127);
not I_6503 (I113437,I113420);
nor I_6504 (I112999,I113276,I113437);
nand I_6505 (I112984,I113293,I113437);
nor I_6506 (I112993,I113039,I113420);
DFFARX1 I_6507 (I113420,I2859,I113013,I113002,);
not I_6508 (I113540,I2866);
DFFARX1 I_6509 (I162596,I2859,I113540,I113566,);
nand I_6510 (I113574,I162608,I162587);
and I_6511 (I113591,I113574,I162611);
DFFARX1 I_6512 (I113591,I2859,I113540,I113617,);
nor I_6513 (I113508,I113617,I113566);
not I_6514 (I113639,I113617);
DFFARX1 I_6515 (I162602,I2859,I113540,I113665,);
nand I_6516 (I113673,I113665,I162584);
not I_6517 (I113690,I113673);
DFFARX1 I_6518 (I113690,I2859,I113540,I113716,);
not I_6519 (I113532,I113716);
nor I_6520 (I113738,I113566,I113673);
nor I_6521 (I113514,I113617,I113738);
DFFARX1 I_6522 (I162599,I2859,I113540,I113778,);
DFFARX1 I_6523 (I113778,I2859,I113540,I113795,);
not I_6524 (I113803,I113795);
not I_6525 (I113820,I113778);
nand I_6526 (I113517,I113820,I113639);
nand I_6527 (I113851,I162584,I162590);
and I_6528 (I113868,I113851,I162593);
DFFARX1 I_6529 (I113868,I2859,I113540,I113894,);
nor I_6530 (I113902,I113894,I113566);
DFFARX1 I_6531 (I113902,I2859,I113540,I113505,);
DFFARX1 I_6532 (I113894,I2859,I113540,I113523,);
nor I_6533 (I113947,I162605,I162590);
not I_6534 (I113964,I113947);
nor I_6535 (I113526,I113803,I113964);
nand I_6536 (I113511,I113820,I113964);
nor I_6537 (I113520,I113566,I113947);
DFFARX1 I_6538 (I113947,I2859,I113540,I113529,);
not I_6539 (I114067,I2866);
DFFARX1 I_6540 (I342838,I2859,I114067,I114093,);
nand I_6541 (I114101,I342841,I342835);
and I_6542 (I114118,I114101,I342847);
DFFARX1 I_6543 (I114118,I2859,I114067,I114144,);
nor I_6544 (I114035,I114144,I114093);
not I_6545 (I114166,I114144);
DFFARX1 I_6546 (I342850,I2859,I114067,I114192,);
nand I_6547 (I114200,I114192,I342841);
not I_6548 (I114217,I114200);
DFFARX1 I_6549 (I114217,I2859,I114067,I114243,);
not I_6550 (I114059,I114243);
nor I_6551 (I114265,I114093,I114200);
nor I_6552 (I114041,I114144,I114265);
DFFARX1 I_6553 (I342853,I2859,I114067,I114305,);
DFFARX1 I_6554 (I114305,I2859,I114067,I114322,);
not I_6555 (I114330,I114322);
not I_6556 (I114347,I114305);
nand I_6557 (I114044,I114347,I114166);
nand I_6558 (I114378,I342835,I342844);
and I_6559 (I114395,I114378,I342838);
DFFARX1 I_6560 (I114395,I2859,I114067,I114421,);
nor I_6561 (I114429,I114421,I114093);
DFFARX1 I_6562 (I114429,I2859,I114067,I114032,);
DFFARX1 I_6563 (I114421,I2859,I114067,I114050,);
nor I_6564 (I114474,I342856,I342844);
not I_6565 (I114491,I114474);
nor I_6566 (I114053,I114330,I114491);
nand I_6567 (I114038,I114347,I114491);
nor I_6568 (I114047,I114093,I114474);
DFFARX1 I_6569 (I114474,I2859,I114067,I114056,);
not I_6570 (I114594,I2866);
DFFARX1 I_6571 (I317500,I2859,I114594,I114620,);
nand I_6572 (I114628,I317491,I317506);
and I_6573 (I114645,I114628,I317512);
DFFARX1 I_6574 (I114645,I2859,I114594,I114671,);
nor I_6575 (I114562,I114671,I114620);
not I_6576 (I114693,I114671);
DFFARX1 I_6577 (I317497,I2859,I114594,I114719,);
nand I_6578 (I114727,I114719,I317491);
not I_6579 (I114744,I114727);
DFFARX1 I_6580 (I114744,I2859,I114594,I114770,);
not I_6581 (I114586,I114770);
nor I_6582 (I114792,I114620,I114727);
nor I_6583 (I114568,I114671,I114792);
DFFARX1 I_6584 (I317494,I2859,I114594,I114832,);
DFFARX1 I_6585 (I114832,I2859,I114594,I114849,);
not I_6586 (I114857,I114849);
not I_6587 (I114874,I114832);
nand I_6588 (I114571,I114874,I114693);
nand I_6589 (I114905,I317488,I317503);
and I_6590 (I114922,I114905,I317488);
DFFARX1 I_6591 (I114922,I2859,I114594,I114948,);
nor I_6592 (I114956,I114948,I114620);
DFFARX1 I_6593 (I114956,I2859,I114594,I114559,);
DFFARX1 I_6594 (I114948,I2859,I114594,I114577,);
nor I_6595 (I115001,I317509,I317503);
not I_6596 (I115018,I115001);
nor I_6597 (I114580,I114857,I115018);
nand I_6598 (I114565,I114874,I115018);
nor I_6599 (I114574,I114620,I115001);
DFFARX1 I_6600 (I115001,I2859,I114594,I114583,);
not I_6601 (I115121,I2866);
DFFARX1 I_6602 (I415343,I2859,I115121,I115147,);
nand I_6603 (I115155,I415340,I415343);
and I_6604 (I115172,I115155,I415352);
DFFARX1 I_6605 (I115172,I2859,I115121,I115198,);
nor I_6606 (I115089,I115198,I115147);
not I_6607 (I115220,I115198);
DFFARX1 I_6608 (I415340,I2859,I115121,I115246,);
nand I_6609 (I115254,I115246,I415358);
not I_6610 (I115271,I115254);
DFFARX1 I_6611 (I115271,I2859,I115121,I115297,);
not I_6612 (I115113,I115297);
nor I_6613 (I115319,I115147,I115254);
nor I_6614 (I115095,I115198,I115319);
DFFARX1 I_6615 (I415346,I2859,I115121,I115359,);
DFFARX1 I_6616 (I115359,I2859,I115121,I115376,);
not I_6617 (I115384,I115376);
not I_6618 (I115401,I115359);
nand I_6619 (I115098,I115401,I115220);
nand I_6620 (I115432,I415355,I415361);
and I_6621 (I115449,I115432,I415346);
DFFARX1 I_6622 (I115449,I2859,I115121,I115475,);
nor I_6623 (I115483,I115475,I115147);
DFFARX1 I_6624 (I115483,I2859,I115121,I115086,);
DFFARX1 I_6625 (I115475,I2859,I115121,I115104,);
nor I_6626 (I115528,I415349,I415361);
not I_6627 (I115545,I115528);
nor I_6628 (I115107,I115384,I115545);
nand I_6629 (I115092,I115401,I115545);
nor I_6630 (I115101,I115147,I115528);
DFFARX1 I_6631 (I115528,I2859,I115121,I115110,);
not I_6632 (I115648,I2866);
DFFARX1 I_6633 (I251611,I2859,I115648,I115674,);
nand I_6634 (I115682,I251596,I251599);
and I_6635 (I115699,I115682,I251614);
DFFARX1 I_6636 (I115699,I2859,I115648,I115725,);
nor I_6637 (I115616,I115725,I115674);
not I_6638 (I115747,I115725);
DFFARX1 I_6639 (I251608,I2859,I115648,I115773,);
nand I_6640 (I115781,I115773,I251599);
not I_6641 (I115798,I115781);
DFFARX1 I_6642 (I115798,I2859,I115648,I115824,);
not I_6643 (I115640,I115824);
nor I_6644 (I115846,I115674,I115781);
nor I_6645 (I115622,I115725,I115846);
DFFARX1 I_6646 (I251605,I2859,I115648,I115886,);
DFFARX1 I_6647 (I115886,I2859,I115648,I115903,);
not I_6648 (I115911,I115903);
not I_6649 (I115928,I115886);
nand I_6650 (I115625,I115928,I115747);
nand I_6651 (I115959,I251620,I251596);
and I_6652 (I115976,I115959,I251617);
DFFARX1 I_6653 (I115976,I2859,I115648,I116002,);
nor I_6654 (I116010,I116002,I115674);
DFFARX1 I_6655 (I116010,I2859,I115648,I115613,);
DFFARX1 I_6656 (I116002,I2859,I115648,I115631,);
nor I_6657 (I116055,I251602,I251596);
not I_6658 (I116072,I116055);
nor I_6659 (I115634,I115911,I116072);
nand I_6660 (I115619,I115928,I116072);
nor I_6661 (I115628,I115674,I116055);
DFFARX1 I_6662 (I116055,I2859,I115648,I115637,);
not I_6663 (I116175,I2866);
DFFARX1 I_6664 (I412844,I2859,I116175,I116201,);
nand I_6665 (I116209,I412841,I412859);
and I_6666 (I116226,I116209,I412850);
DFFARX1 I_6667 (I116226,I2859,I116175,I116252,);
nor I_6668 (I116143,I116252,I116201);
not I_6669 (I116274,I116252);
DFFARX1 I_6670 (I412865,I2859,I116175,I116300,);
nand I_6671 (I116308,I116300,I412847);
not I_6672 (I116325,I116308);
DFFARX1 I_6673 (I116325,I2859,I116175,I116351,);
not I_6674 (I116167,I116351);
nor I_6675 (I116373,I116201,I116308);
nor I_6676 (I116149,I116252,I116373);
DFFARX1 I_6677 (I412853,I2859,I116175,I116413,);
DFFARX1 I_6678 (I116413,I2859,I116175,I116430,);
not I_6679 (I116438,I116430);
not I_6680 (I116455,I116413);
nand I_6681 (I116152,I116455,I116274);
nand I_6682 (I116486,I412841,I412868);
and I_6683 (I116503,I116486,I412856);
DFFARX1 I_6684 (I116503,I2859,I116175,I116529,);
nor I_6685 (I116537,I116529,I116201);
DFFARX1 I_6686 (I116537,I2859,I116175,I116140,);
DFFARX1 I_6687 (I116529,I2859,I116175,I116158,);
nor I_6688 (I116582,I412862,I412868);
not I_6689 (I116599,I116582);
nor I_6690 (I116161,I116438,I116599);
nand I_6691 (I116146,I116455,I116599);
nor I_6692 (I116155,I116201,I116582);
DFFARX1 I_6693 (I116582,I2859,I116175,I116164,);
not I_6694 (I116702,I2866);
DFFARX1 I_6695 (I239473,I2859,I116702,I116728,);
nand I_6696 (I116736,I239458,I239461);
and I_6697 (I116753,I116736,I239476);
DFFARX1 I_6698 (I116753,I2859,I116702,I116779,);
nor I_6699 (I116670,I116779,I116728);
not I_6700 (I116801,I116779);
DFFARX1 I_6701 (I239470,I2859,I116702,I116827,);
nand I_6702 (I116835,I116827,I239461);
not I_6703 (I116852,I116835);
DFFARX1 I_6704 (I116852,I2859,I116702,I116878,);
not I_6705 (I116694,I116878);
nor I_6706 (I116900,I116728,I116835);
nor I_6707 (I116676,I116779,I116900);
DFFARX1 I_6708 (I239467,I2859,I116702,I116940,);
DFFARX1 I_6709 (I116940,I2859,I116702,I116957,);
not I_6710 (I116965,I116957);
not I_6711 (I116982,I116940);
nand I_6712 (I116679,I116982,I116801);
nand I_6713 (I117013,I239482,I239458);
and I_6714 (I117030,I117013,I239479);
DFFARX1 I_6715 (I117030,I2859,I116702,I117056,);
nor I_6716 (I117064,I117056,I116728);
DFFARX1 I_6717 (I117064,I2859,I116702,I116667,);
DFFARX1 I_6718 (I117056,I2859,I116702,I116685,);
nor I_6719 (I117109,I239464,I239458);
not I_6720 (I117126,I117109);
nor I_6721 (I116688,I116965,I117126);
nand I_6722 (I116673,I116982,I117126);
nor I_6723 (I116682,I116728,I117109);
DFFARX1 I_6724 (I117109,I2859,I116702,I116691,);
not I_6725 (I117229,I2866);
DFFARX1 I_6726 (I394110,I2859,I117229,I117255,);
nand I_6727 (I117263,I394107,I394125);
and I_6728 (I117280,I117263,I394116);
DFFARX1 I_6729 (I117280,I2859,I117229,I117306,);
nor I_6730 (I117197,I117306,I117255);
not I_6731 (I117328,I117306);
DFFARX1 I_6732 (I394131,I2859,I117229,I117354,);
nand I_6733 (I117362,I117354,I394113);
not I_6734 (I117379,I117362);
DFFARX1 I_6735 (I117379,I2859,I117229,I117405,);
not I_6736 (I117221,I117405);
nor I_6737 (I117427,I117255,I117362);
nor I_6738 (I117203,I117306,I117427);
DFFARX1 I_6739 (I394119,I2859,I117229,I117467,);
DFFARX1 I_6740 (I117467,I2859,I117229,I117484,);
not I_6741 (I117492,I117484);
not I_6742 (I117509,I117467);
nand I_6743 (I117206,I117509,I117328);
nand I_6744 (I117540,I394107,I394134);
and I_6745 (I117557,I117540,I394122);
DFFARX1 I_6746 (I117557,I2859,I117229,I117583,);
nor I_6747 (I117591,I117583,I117255);
DFFARX1 I_6748 (I117591,I2859,I117229,I117194,);
DFFARX1 I_6749 (I117583,I2859,I117229,I117212,);
nor I_6750 (I117636,I394128,I394134);
not I_6751 (I117653,I117636);
nor I_6752 (I117215,I117492,I117653);
nand I_6753 (I117200,I117509,I117653);
nor I_6754 (I117209,I117255,I117636);
DFFARX1 I_6755 (I117636,I2859,I117229,I117218,);
not I_6756 (I117756,I2866);
DFFARX1 I_6757 (I567171,I2859,I117756,I117782,);
nand I_6758 (I117790,I567150,I567150);
and I_6759 (I117807,I117790,I567177);
DFFARX1 I_6760 (I117807,I2859,I117756,I117833,);
nor I_6761 (I117724,I117833,I117782);
not I_6762 (I117855,I117833);
DFFARX1 I_6763 (I567165,I2859,I117756,I117881,);
nand I_6764 (I117889,I117881,I567168);
not I_6765 (I117906,I117889);
DFFARX1 I_6766 (I117906,I2859,I117756,I117932,);
not I_6767 (I117748,I117932);
nor I_6768 (I117954,I117782,I117889);
nor I_6769 (I117730,I117833,I117954);
DFFARX1 I_6770 (I567159,I2859,I117756,I117994,);
DFFARX1 I_6771 (I117994,I2859,I117756,I118011,);
not I_6772 (I118019,I118011);
not I_6773 (I118036,I117994);
nand I_6774 (I117733,I118036,I117855);
nand I_6775 (I118067,I567156,I567153);
and I_6776 (I118084,I118067,I567174);
DFFARX1 I_6777 (I118084,I2859,I117756,I118110,);
nor I_6778 (I118118,I118110,I117782);
DFFARX1 I_6779 (I118118,I2859,I117756,I117721,);
DFFARX1 I_6780 (I118110,I2859,I117756,I117739,);
nor I_6781 (I118163,I567162,I567153);
not I_6782 (I118180,I118163);
nor I_6783 (I117742,I118019,I118180);
nand I_6784 (I117727,I118036,I118180);
nor I_6785 (I117736,I117782,I118163);
DFFARX1 I_6786 (I118163,I2859,I117756,I117745,);
not I_6787 (I118283,I2866);
DFFARX1 I_6788 (I541586,I2859,I118283,I118309,);
nand I_6789 (I118317,I541565,I541565);
and I_6790 (I118334,I118317,I541592);
DFFARX1 I_6791 (I118334,I2859,I118283,I118360,);
nor I_6792 (I118251,I118360,I118309);
not I_6793 (I118382,I118360);
DFFARX1 I_6794 (I541580,I2859,I118283,I118408,);
nand I_6795 (I118416,I118408,I541583);
not I_6796 (I118433,I118416);
DFFARX1 I_6797 (I118433,I2859,I118283,I118459,);
not I_6798 (I118275,I118459);
nor I_6799 (I118481,I118309,I118416);
nor I_6800 (I118257,I118360,I118481);
DFFARX1 I_6801 (I541574,I2859,I118283,I118521,);
DFFARX1 I_6802 (I118521,I2859,I118283,I118538,);
not I_6803 (I118546,I118538);
not I_6804 (I118563,I118521);
nand I_6805 (I118260,I118563,I118382);
nand I_6806 (I118594,I541571,I541568);
and I_6807 (I118611,I118594,I541589);
DFFARX1 I_6808 (I118611,I2859,I118283,I118637,);
nor I_6809 (I118645,I118637,I118309);
DFFARX1 I_6810 (I118645,I2859,I118283,I118248,);
DFFARX1 I_6811 (I118637,I2859,I118283,I118266,);
nor I_6812 (I118690,I541577,I541568);
not I_6813 (I118707,I118690);
nor I_6814 (I118269,I118546,I118707);
nand I_6815 (I118254,I118563,I118707);
nor I_6816 (I118263,I118309,I118690);
DFFARX1 I_6817 (I118690,I2859,I118283,I118272,);
not I_6818 (I118810,I2866);
DFFARX1 I_6819 (I182180,I2859,I118810,I118836,);
nand I_6820 (I118844,I182192,I182171);
and I_6821 (I118861,I118844,I182195);
DFFARX1 I_6822 (I118861,I2859,I118810,I118887,);
nor I_6823 (I118778,I118887,I118836);
not I_6824 (I118909,I118887);
DFFARX1 I_6825 (I182186,I2859,I118810,I118935,);
nand I_6826 (I118943,I118935,I182168);
not I_6827 (I118960,I118943);
DFFARX1 I_6828 (I118960,I2859,I118810,I118986,);
not I_6829 (I118802,I118986);
nor I_6830 (I119008,I118836,I118943);
nor I_6831 (I118784,I118887,I119008);
DFFARX1 I_6832 (I182183,I2859,I118810,I119048,);
DFFARX1 I_6833 (I119048,I2859,I118810,I119065,);
not I_6834 (I119073,I119065);
not I_6835 (I119090,I119048);
nand I_6836 (I118787,I119090,I118909);
nand I_6837 (I119121,I182168,I182174);
and I_6838 (I119138,I119121,I182177);
DFFARX1 I_6839 (I119138,I2859,I118810,I119164,);
nor I_6840 (I119172,I119164,I118836);
DFFARX1 I_6841 (I119172,I2859,I118810,I118775,);
DFFARX1 I_6842 (I119164,I2859,I118810,I118793,);
nor I_6843 (I119217,I182189,I182174);
not I_6844 (I119234,I119217);
nor I_6845 (I118796,I119073,I119234);
nand I_6846 (I118781,I119090,I119234);
nor I_6847 (I118790,I118836,I119217);
DFFARX1 I_6848 (I119217,I2859,I118810,I118799,);
not I_6849 (I119337,I2866);
DFFARX1 I_6850 (I63202,I2859,I119337,I119363,);
nand I_6851 (I119371,I63202,I63208);
and I_6852 (I119388,I119371,I63226);
DFFARX1 I_6853 (I119388,I2859,I119337,I119414,);
nor I_6854 (I119305,I119414,I119363);
not I_6855 (I119436,I119414);
DFFARX1 I_6856 (I63214,I2859,I119337,I119462,);
nand I_6857 (I119470,I119462,I63211);
not I_6858 (I119487,I119470);
DFFARX1 I_6859 (I119487,I2859,I119337,I119513,);
not I_6860 (I119329,I119513);
nor I_6861 (I119535,I119363,I119470);
nor I_6862 (I119311,I119414,I119535);
DFFARX1 I_6863 (I63220,I2859,I119337,I119575,);
DFFARX1 I_6864 (I119575,I2859,I119337,I119592,);
not I_6865 (I119600,I119592);
not I_6866 (I119617,I119575);
nand I_6867 (I119314,I119617,I119436);
nand I_6868 (I119648,I63205,I63205);
and I_6869 (I119665,I119648,I63217);
DFFARX1 I_6870 (I119665,I2859,I119337,I119691,);
nor I_6871 (I119699,I119691,I119363);
DFFARX1 I_6872 (I119699,I2859,I119337,I119302,);
DFFARX1 I_6873 (I119691,I2859,I119337,I119320,);
nor I_6874 (I119744,I63223,I63205);
not I_6875 (I119761,I119744);
nor I_6876 (I119323,I119600,I119761);
nand I_6877 (I119308,I119617,I119761);
nor I_6878 (I119317,I119363,I119744);
DFFARX1 I_6879 (I119744,I2859,I119337,I119326,);
not I_6880 (I119864,I2866);
DFFARX1 I_6881 (I249299,I2859,I119864,I119890,);
nand I_6882 (I119898,I249284,I249287);
and I_6883 (I119915,I119898,I249302);
DFFARX1 I_6884 (I119915,I2859,I119864,I119941,);
nor I_6885 (I119832,I119941,I119890);
not I_6886 (I119963,I119941);
DFFARX1 I_6887 (I249296,I2859,I119864,I119989,);
nand I_6888 (I119997,I119989,I249287);
not I_6889 (I120014,I119997);
DFFARX1 I_6890 (I120014,I2859,I119864,I120040,);
not I_6891 (I119856,I120040);
nor I_6892 (I120062,I119890,I119997);
nor I_6893 (I119838,I119941,I120062);
DFFARX1 I_6894 (I249293,I2859,I119864,I120102,);
DFFARX1 I_6895 (I120102,I2859,I119864,I120119,);
not I_6896 (I120127,I120119);
not I_6897 (I120144,I120102);
nand I_6898 (I119841,I120144,I119963);
nand I_6899 (I120175,I249308,I249284);
and I_6900 (I120192,I120175,I249305);
DFFARX1 I_6901 (I120192,I2859,I119864,I120218,);
nor I_6902 (I120226,I120218,I119890);
DFFARX1 I_6903 (I120226,I2859,I119864,I119829,);
DFFARX1 I_6904 (I120218,I2859,I119864,I119847,);
nor I_6905 (I120271,I249290,I249284);
not I_6906 (I120288,I120271);
nor I_6907 (I119850,I120127,I120288);
nand I_6908 (I119835,I120144,I120288);
nor I_6909 (I119844,I119890,I120271);
DFFARX1 I_6910 (I120271,I2859,I119864,I119853,);
not I_6911 (I120391,I2866);
DFFARX1 I_6912 (I333879,I2859,I120391,I120417,);
nand I_6913 (I120425,I333882,I333876);
and I_6914 (I120442,I120425,I333888);
DFFARX1 I_6915 (I120442,I2859,I120391,I120468,);
nor I_6916 (I120359,I120468,I120417);
not I_6917 (I120490,I120468);
DFFARX1 I_6918 (I333891,I2859,I120391,I120516,);
nand I_6919 (I120524,I120516,I333882);
not I_6920 (I120541,I120524);
DFFARX1 I_6921 (I120541,I2859,I120391,I120567,);
not I_6922 (I120383,I120567);
nor I_6923 (I120589,I120417,I120524);
nor I_6924 (I120365,I120468,I120589);
DFFARX1 I_6925 (I333894,I2859,I120391,I120629,);
DFFARX1 I_6926 (I120629,I2859,I120391,I120646,);
not I_6927 (I120654,I120646);
not I_6928 (I120671,I120629);
nand I_6929 (I120368,I120671,I120490);
nand I_6930 (I120702,I333876,I333885);
and I_6931 (I120719,I120702,I333879);
DFFARX1 I_6932 (I120719,I2859,I120391,I120745,);
nor I_6933 (I120753,I120745,I120417);
DFFARX1 I_6934 (I120753,I2859,I120391,I120356,);
DFFARX1 I_6935 (I120745,I2859,I120391,I120374,);
nor I_6936 (I120798,I333897,I333885);
not I_6937 (I120815,I120798);
nor I_6938 (I120377,I120654,I120815);
nand I_6939 (I120362,I120671,I120815);
nor I_6940 (I120371,I120417,I120798);
DFFARX1 I_6941 (I120798,I2859,I120391,I120380,);
not I_6942 (I120918,I2866);
DFFARX1 I_6943 (I522965,I2859,I120918,I120944,);
nand I_6944 (I120952,I522962,I522953);
and I_6945 (I120969,I120952,I522950);
DFFARX1 I_6946 (I120969,I2859,I120918,I120995,);
nor I_6947 (I120886,I120995,I120944);
not I_6948 (I121017,I120995);
DFFARX1 I_6949 (I522959,I2859,I120918,I121043,);
nand I_6950 (I121051,I121043,I522968);
not I_6951 (I121068,I121051);
DFFARX1 I_6952 (I121068,I2859,I120918,I121094,);
not I_6953 (I120910,I121094);
nor I_6954 (I121116,I120944,I121051);
nor I_6955 (I120892,I120995,I121116);
DFFARX1 I_6956 (I522971,I2859,I120918,I121156,);
DFFARX1 I_6957 (I121156,I2859,I120918,I121173,);
not I_6958 (I121181,I121173);
not I_6959 (I121198,I121156);
nand I_6960 (I120895,I121198,I121017);
nand I_6961 (I121229,I522950,I522956);
and I_6962 (I121246,I121229,I522974);
DFFARX1 I_6963 (I121246,I2859,I120918,I121272,);
nor I_6964 (I121280,I121272,I120944);
DFFARX1 I_6965 (I121280,I2859,I120918,I120883,);
DFFARX1 I_6966 (I121272,I2859,I120918,I120901,);
nor I_6967 (I121325,I522953,I522956);
not I_6968 (I121342,I121325);
nor I_6969 (I120904,I121181,I121342);
nand I_6970 (I120889,I121198,I121342);
nor I_6971 (I120898,I120944,I121325);
DFFARX1 I_6972 (I121325,I2859,I120918,I120907,);
not I_6973 (I121445,I2866);
DFFARX1 I_6974 (I79267,I2859,I121445,I121471,);
nand I_6975 (I121479,I79267,I79273);
and I_6976 (I121496,I121479,I79291);
DFFARX1 I_6977 (I121496,I2859,I121445,I121522,);
nor I_6978 (I121413,I121522,I121471);
not I_6979 (I121544,I121522);
DFFARX1 I_6980 (I79279,I2859,I121445,I121570,);
nand I_6981 (I121578,I121570,I79276);
not I_6982 (I121595,I121578);
DFFARX1 I_6983 (I121595,I2859,I121445,I121621,);
not I_6984 (I121437,I121621);
nor I_6985 (I121643,I121471,I121578);
nor I_6986 (I121419,I121522,I121643);
DFFARX1 I_6987 (I79285,I2859,I121445,I121683,);
DFFARX1 I_6988 (I121683,I2859,I121445,I121700,);
not I_6989 (I121708,I121700);
not I_6990 (I121725,I121683);
nand I_6991 (I121422,I121725,I121544);
nand I_6992 (I121756,I79270,I79270);
and I_6993 (I121773,I121756,I79282);
DFFARX1 I_6994 (I121773,I2859,I121445,I121799,);
nor I_6995 (I121807,I121799,I121471);
DFFARX1 I_6996 (I121807,I2859,I121445,I121410,);
DFFARX1 I_6997 (I121799,I2859,I121445,I121428,);
nor I_6998 (I121852,I79288,I79270);
not I_6999 (I121869,I121852);
nor I_7000 (I121431,I121708,I121869);
nand I_7001 (I121416,I121725,I121869);
nor I_7002 (I121425,I121471,I121852);
DFFARX1 I_7003 (I121852,I2859,I121445,I121434,);
not I_7004 (I121972,I2866);
DFFARX1 I_7005 (I481096,I2859,I121972,I121998,);
nand I_7006 (I122006,I481111,I481096);
and I_7007 (I122023,I122006,I481114);
DFFARX1 I_7008 (I122023,I2859,I121972,I122049,);
nor I_7009 (I121940,I122049,I121998);
not I_7010 (I122071,I122049);
DFFARX1 I_7011 (I481120,I2859,I121972,I122097,);
nand I_7012 (I122105,I122097,I481102);
not I_7013 (I122122,I122105);
DFFARX1 I_7014 (I122122,I2859,I121972,I122148,);
not I_7015 (I121964,I122148);
nor I_7016 (I122170,I121998,I122105);
nor I_7017 (I121946,I122049,I122170);
DFFARX1 I_7018 (I481099,I2859,I121972,I122210,);
DFFARX1 I_7019 (I122210,I2859,I121972,I122227,);
not I_7020 (I122235,I122227);
not I_7021 (I122252,I122210);
nand I_7022 (I121949,I122252,I122071);
nand I_7023 (I122283,I481099,I481105);
and I_7024 (I122300,I122283,I481117);
DFFARX1 I_7025 (I122300,I2859,I121972,I122326,);
nor I_7026 (I122334,I122326,I121998);
DFFARX1 I_7027 (I122334,I2859,I121972,I121937,);
DFFARX1 I_7028 (I122326,I2859,I121972,I121955,);
nor I_7029 (I122379,I481108,I481105);
not I_7030 (I122396,I122379);
nor I_7031 (I121958,I122235,I122396);
nand I_7032 (I121943,I122252,I122396);
nor I_7033 (I121952,I121998,I122379);
DFFARX1 I_7034 (I122379,I2859,I121972,I121961,);
not I_7035 (I122499,I2866);
DFFARX1 I_7036 (I350216,I2859,I122499,I122525,);
nand I_7037 (I122533,I350219,I350213);
and I_7038 (I122550,I122533,I350225);
DFFARX1 I_7039 (I122550,I2859,I122499,I122576,);
nor I_7040 (I122467,I122576,I122525);
not I_7041 (I122598,I122576);
DFFARX1 I_7042 (I350228,I2859,I122499,I122624,);
nand I_7043 (I122632,I122624,I350219);
not I_7044 (I122649,I122632);
DFFARX1 I_7045 (I122649,I2859,I122499,I122675,);
not I_7046 (I122491,I122675);
nor I_7047 (I122697,I122525,I122632);
nor I_7048 (I122473,I122576,I122697);
DFFARX1 I_7049 (I350231,I2859,I122499,I122737,);
DFFARX1 I_7050 (I122737,I2859,I122499,I122754,);
not I_7051 (I122762,I122754);
not I_7052 (I122779,I122737);
nand I_7053 (I122476,I122779,I122598);
nand I_7054 (I122810,I350213,I350222);
and I_7055 (I122827,I122810,I350216);
DFFARX1 I_7056 (I122827,I2859,I122499,I122853,);
nor I_7057 (I122861,I122853,I122525);
DFFARX1 I_7058 (I122861,I2859,I122499,I122464,);
DFFARX1 I_7059 (I122853,I2859,I122499,I122482,);
nor I_7060 (I122906,I350234,I350222);
not I_7061 (I122923,I122906);
nor I_7062 (I122485,I122762,I122923);
nand I_7063 (I122470,I122779,I122923);
nor I_7064 (I122479,I122525,I122906);
DFFARX1 I_7065 (I122906,I2859,I122499,I122488,);
not I_7066 (I123026,I2866);
DFFARX1 I_7067 (I204883,I2859,I123026,I123052,);
nand I_7068 (I123060,I204883,I204895);
and I_7069 (I123077,I123060,I204880);
DFFARX1 I_7070 (I123077,I2859,I123026,I123103,);
nor I_7071 (I122994,I123103,I123052);
not I_7072 (I123125,I123103);
DFFARX1 I_7073 (I204904,I2859,I123026,I123151,);
nand I_7074 (I123159,I123151,I204901);
not I_7075 (I123176,I123159);
DFFARX1 I_7076 (I123176,I2859,I123026,I123202,);
not I_7077 (I123018,I123202);
nor I_7078 (I123224,I123052,I123159);
nor I_7079 (I123000,I123103,I123224);
DFFARX1 I_7080 (I204892,I2859,I123026,I123264,);
DFFARX1 I_7081 (I123264,I2859,I123026,I123281,);
not I_7082 (I123289,I123281);
not I_7083 (I123306,I123264);
nand I_7084 (I123003,I123306,I123125);
nand I_7085 (I123337,I204880,I204889);
and I_7086 (I123354,I123337,I204898);
DFFARX1 I_7087 (I123354,I2859,I123026,I123380,);
nor I_7088 (I123388,I123380,I123052);
DFFARX1 I_7089 (I123388,I2859,I123026,I122991,);
DFFARX1 I_7090 (I123380,I2859,I123026,I123009,);
nor I_7091 (I123433,I204886,I204889);
not I_7092 (I123450,I123433);
nor I_7093 (I123012,I123289,I123450);
nand I_7094 (I122997,I123306,I123450);
nor I_7095 (I123006,I123052,I123433);
DFFARX1 I_7096 (I123433,I2859,I123026,I123015,);
not I_7097 (I123553,I2866);
DFFARX1 I_7098 (I510116,I2859,I123553,I123579,);
nand I_7099 (I123587,I510098,I510122);
and I_7100 (I123604,I123587,I510113);
DFFARX1 I_7101 (I123604,I2859,I123553,I123630,);
nor I_7102 (I123521,I123630,I123579);
not I_7103 (I123652,I123630);
DFFARX1 I_7104 (I510119,I2859,I123553,I123678,);
nand I_7105 (I123686,I123678,I510107);
not I_7106 (I123703,I123686);
DFFARX1 I_7107 (I123703,I2859,I123553,I123729,);
not I_7108 (I123545,I123729);
nor I_7109 (I123751,I123579,I123686);
nor I_7110 (I123527,I123630,I123751);
DFFARX1 I_7111 (I510098,I2859,I123553,I123791,);
DFFARX1 I_7112 (I123791,I2859,I123553,I123808,);
not I_7113 (I123816,I123808);
not I_7114 (I123833,I123791);
nand I_7115 (I123530,I123833,I123652);
nand I_7116 (I123864,I510104,I510101);
and I_7117 (I123881,I123864,I510110);
DFFARX1 I_7118 (I123881,I2859,I123553,I123907,);
nor I_7119 (I123915,I123907,I123579);
DFFARX1 I_7120 (I123915,I2859,I123553,I123518,);
DFFARX1 I_7121 (I123907,I2859,I123553,I123536,);
nor I_7122 (I123960,I510101,I510101);
not I_7123 (I123977,I123960);
nor I_7124 (I123539,I123816,I123977);
nand I_7125 (I123524,I123833,I123977);
nor I_7126 (I123533,I123579,I123960);
DFFARX1 I_7127 (I123960,I2859,I123553,I123542,);
not I_7128 (I124080,I2866);
DFFARX1 I_7129 (I325447,I2859,I124080,I124106,);
nand I_7130 (I124114,I325450,I325444);
and I_7131 (I124131,I124114,I325456);
DFFARX1 I_7132 (I124131,I2859,I124080,I124157,);
nor I_7133 (I124048,I124157,I124106);
not I_7134 (I124179,I124157);
DFFARX1 I_7135 (I325459,I2859,I124080,I124205,);
nand I_7136 (I124213,I124205,I325450);
not I_7137 (I124230,I124213);
DFFARX1 I_7138 (I124230,I2859,I124080,I124256,);
not I_7139 (I124072,I124256);
nor I_7140 (I124278,I124106,I124213);
nor I_7141 (I124054,I124157,I124278);
DFFARX1 I_7142 (I325462,I2859,I124080,I124318,);
DFFARX1 I_7143 (I124318,I2859,I124080,I124335,);
not I_7144 (I124343,I124335);
not I_7145 (I124360,I124318);
nand I_7146 (I124057,I124360,I124179);
nand I_7147 (I124391,I325444,I325453);
and I_7148 (I124408,I124391,I325447);
DFFARX1 I_7149 (I124408,I2859,I124080,I124434,);
nor I_7150 (I124442,I124434,I124106);
DFFARX1 I_7151 (I124442,I2859,I124080,I124045,);
DFFARX1 I_7152 (I124434,I2859,I124080,I124063,);
nor I_7153 (I124487,I325465,I325453);
not I_7154 (I124504,I124487);
nor I_7155 (I124066,I124343,I124504);
nand I_7156 (I124051,I124360,I124504);
nor I_7157 (I124060,I124106,I124487);
DFFARX1 I_7158 (I124487,I2859,I124080,I124069,);
not I_7159 (I124607,I2866);
DFFARX1 I_7160 (I343892,I2859,I124607,I124633,);
nand I_7161 (I124641,I343895,I343889);
and I_7162 (I124658,I124641,I343901);
DFFARX1 I_7163 (I124658,I2859,I124607,I124684,);
nor I_7164 (I124575,I124684,I124633);
not I_7165 (I124706,I124684);
DFFARX1 I_7166 (I343904,I2859,I124607,I124732,);
nand I_7167 (I124740,I124732,I343895);
not I_7168 (I124757,I124740);
DFFARX1 I_7169 (I124757,I2859,I124607,I124783,);
not I_7170 (I124599,I124783);
nor I_7171 (I124805,I124633,I124740);
nor I_7172 (I124581,I124684,I124805);
DFFARX1 I_7173 (I343907,I2859,I124607,I124845,);
DFFARX1 I_7174 (I124845,I2859,I124607,I124862,);
not I_7175 (I124870,I124862);
not I_7176 (I124887,I124845);
nand I_7177 (I124584,I124887,I124706);
nand I_7178 (I124918,I343889,I343898);
and I_7179 (I124935,I124918,I343892);
DFFARX1 I_7180 (I124935,I2859,I124607,I124961,);
nor I_7181 (I124969,I124961,I124633);
DFFARX1 I_7182 (I124969,I2859,I124607,I124572,);
DFFARX1 I_7183 (I124961,I2859,I124607,I124590,);
nor I_7184 (I125014,I343910,I343898);
not I_7185 (I125031,I125014);
nor I_7186 (I124593,I124870,I125031);
nand I_7187 (I124578,I124887,I125031);
nor I_7188 (I124587,I124633,I125014);
DFFARX1 I_7189 (I125014,I2859,I124607,I124596,);
not I_7190 (I125134,I2866);
DFFARX1 I_7191 (I529901,I2859,I125134,I125160,);
nand I_7192 (I125168,I529898,I529889);
and I_7193 (I125185,I125168,I529886);
DFFARX1 I_7194 (I125185,I2859,I125134,I125211,);
nor I_7195 (I125102,I125211,I125160);
not I_7196 (I125233,I125211);
DFFARX1 I_7197 (I529895,I2859,I125134,I125259,);
nand I_7198 (I125267,I125259,I529904);
not I_7199 (I125284,I125267);
DFFARX1 I_7200 (I125284,I2859,I125134,I125310,);
not I_7201 (I125126,I125310);
nor I_7202 (I125332,I125160,I125267);
nor I_7203 (I125108,I125211,I125332);
DFFARX1 I_7204 (I529907,I2859,I125134,I125372,);
DFFARX1 I_7205 (I125372,I2859,I125134,I125389,);
not I_7206 (I125397,I125389);
not I_7207 (I125414,I125372);
nand I_7208 (I125111,I125414,I125233);
nand I_7209 (I125445,I529886,I529892);
and I_7210 (I125462,I125445,I529910);
DFFARX1 I_7211 (I125462,I2859,I125134,I125488,);
nor I_7212 (I125496,I125488,I125160);
DFFARX1 I_7213 (I125496,I2859,I125134,I125099,);
DFFARX1 I_7214 (I125488,I2859,I125134,I125117,);
nor I_7215 (I125541,I529889,I529892);
not I_7216 (I125558,I125541);
nor I_7217 (I125120,I125397,I125558);
nand I_7218 (I125105,I125414,I125558);
nor I_7219 (I125114,I125160,I125541);
DFFARX1 I_7220 (I125541,I2859,I125134,I125123,);
not I_7221 (I125661,I2866);
DFFARX1 I_7222 (I328082,I2859,I125661,I125687,);
nand I_7223 (I125695,I328085,I328079);
and I_7224 (I125712,I125695,I328091);
DFFARX1 I_7225 (I125712,I2859,I125661,I125738,);
nor I_7226 (I125629,I125738,I125687);
not I_7227 (I125760,I125738);
DFFARX1 I_7228 (I328094,I2859,I125661,I125786,);
nand I_7229 (I125794,I125786,I328085);
not I_7230 (I125811,I125794);
DFFARX1 I_7231 (I125811,I2859,I125661,I125837,);
not I_7232 (I125653,I125837);
nor I_7233 (I125859,I125687,I125794);
nor I_7234 (I125635,I125738,I125859);
DFFARX1 I_7235 (I328097,I2859,I125661,I125899,);
DFFARX1 I_7236 (I125899,I2859,I125661,I125916,);
not I_7237 (I125924,I125916);
not I_7238 (I125941,I125899);
nand I_7239 (I125638,I125941,I125760);
nand I_7240 (I125972,I328079,I328088);
and I_7241 (I125989,I125972,I328082);
DFFARX1 I_7242 (I125989,I2859,I125661,I126015,);
nor I_7243 (I126023,I126015,I125687);
DFFARX1 I_7244 (I126023,I2859,I125661,I125626,);
DFFARX1 I_7245 (I126015,I2859,I125661,I125644,);
nor I_7246 (I126068,I328100,I328088);
not I_7247 (I126085,I126068);
nor I_7248 (I125647,I125924,I126085);
nand I_7249 (I125632,I125941,I126085);
nor I_7250 (I125641,I125687,I126068);
DFFARX1 I_7251 (I126068,I2859,I125661,I125650,);
not I_7252 (I126188,I2866);
DFFARX1 I_7253 (I551701,I2859,I126188,I126214,);
nand I_7254 (I126222,I551680,I551680);
and I_7255 (I126239,I126222,I551707);
DFFARX1 I_7256 (I126239,I2859,I126188,I126265,);
nor I_7257 (I126156,I126265,I126214);
not I_7258 (I126287,I126265);
DFFARX1 I_7259 (I551695,I2859,I126188,I126313,);
nand I_7260 (I126321,I126313,I551698);
not I_7261 (I126338,I126321);
DFFARX1 I_7262 (I126338,I2859,I126188,I126364,);
not I_7263 (I126180,I126364);
nor I_7264 (I126386,I126214,I126321);
nor I_7265 (I126162,I126265,I126386);
DFFARX1 I_7266 (I551689,I2859,I126188,I126426,);
DFFARX1 I_7267 (I126426,I2859,I126188,I126443,);
not I_7268 (I126451,I126443);
not I_7269 (I126468,I126426);
nand I_7270 (I126165,I126468,I126287);
nand I_7271 (I126499,I551686,I551683);
and I_7272 (I126516,I126499,I551704);
DFFARX1 I_7273 (I126516,I2859,I126188,I126542,);
nor I_7274 (I126550,I126542,I126214);
DFFARX1 I_7275 (I126550,I2859,I126188,I126153,);
DFFARX1 I_7276 (I126542,I2859,I126188,I126171,);
nor I_7277 (I126595,I551692,I551683);
not I_7278 (I126612,I126595);
nor I_7279 (I126174,I126451,I126612);
nand I_7280 (I126159,I126468,I126612);
nor I_7281 (I126168,I126214,I126595);
DFFARX1 I_7282 (I126595,I2859,I126188,I126177,);
not I_7283 (I126715,I2866);
DFFARX1 I_7284 (I161508,I2859,I126715,I126741,);
nand I_7285 (I126749,I161520,I161499);
and I_7286 (I126766,I126749,I161523);
DFFARX1 I_7287 (I126766,I2859,I126715,I126792,);
nor I_7288 (I126683,I126792,I126741);
not I_7289 (I126814,I126792);
DFFARX1 I_7290 (I161514,I2859,I126715,I126840,);
nand I_7291 (I126848,I126840,I161496);
not I_7292 (I126865,I126848);
DFFARX1 I_7293 (I126865,I2859,I126715,I126891,);
not I_7294 (I126707,I126891);
nor I_7295 (I126913,I126741,I126848);
nor I_7296 (I126689,I126792,I126913);
DFFARX1 I_7297 (I161511,I2859,I126715,I126953,);
DFFARX1 I_7298 (I126953,I2859,I126715,I126970,);
not I_7299 (I126978,I126970);
not I_7300 (I126995,I126953);
nand I_7301 (I126692,I126995,I126814);
nand I_7302 (I127026,I161496,I161502);
and I_7303 (I127043,I127026,I161505);
DFFARX1 I_7304 (I127043,I2859,I126715,I127069,);
nor I_7305 (I127077,I127069,I126741);
DFFARX1 I_7306 (I127077,I2859,I126715,I126680,);
DFFARX1 I_7307 (I127069,I2859,I126715,I126698,);
nor I_7308 (I127122,I161517,I161502);
not I_7309 (I127139,I127122);
nor I_7310 (I126701,I126978,I127139);
nand I_7311 (I126686,I126995,I127139);
nor I_7312 (I126695,I126741,I127122);
DFFARX1 I_7313 (I127122,I2859,I126715,I126704,);
not I_7314 (I127242,I2866);
DFFARX1 I_7315 (I205478,I2859,I127242,I127268,);
nand I_7316 (I127276,I205478,I205490);
and I_7317 (I127293,I127276,I205475);
DFFARX1 I_7318 (I127293,I2859,I127242,I127319,);
nor I_7319 (I127210,I127319,I127268);
not I_7320 (I127341,I127319);
DFFARX1 I_7321 (I205499,I2859,I127242,I127367,);
nand I_7322 (I127375,I127367,I205496);
not I_7323 (I127392,I127375);
DFFARX1 I_7324 (I127392,I2859,I127242,I127418,);
not I_7325 (I127234,I127418);
nor I_7326 (I127440,I127268,I127375);
nor I_7327 (I127216,I127319,I127440);
DFFARX1 I_7328 (I205487,I2859,I127242,I127480,);
DFFARX1 I_7329 (I127480,I2859,I127242,I127497,);
not I_7330 (I127505,I127497);
not I_7331 (I127522,I127480);
nand I_7332 (I127219,I127522,I127341);
nand I_7333 (I127553,I205475,I205484);
and I_7334 (I127570,I127553,I205493);
DFFARX1 I_7335 (I127570,I2859,I127242,I127596,);
nor I_7336 (I127604,I127596,I127268);
DFFARX1 I_7337 (I127604,I2859,I127242,I127207,);
DFFARX1 I_7338 (I127596,I2859,I127242,I127225,);
nor I_7339 (I127649,I205481,I205484);
not I_7340 (I127666,I127649);
nor I_7341 (I127228,I127505,I127666);
nand I_7342 (I127213,I127522,I127666);
nor I_7343 (I127222,I127268,I127649);
DFFARX1 I_7344 (I127649,I2859,I127242,I127231,);
not I_7345 (I127769,I2866);
DFFARX1 I_7346 (I84027,I2859,I127769,I127795,);
nand I_7347 (I127803,I84027,I84033);
and I_7348 (I127820,I127803,I84051);
DFFARX1 I_7349 (I127820,I2859,I127769,I127846,);
nor I_7350 (I127737,I127846,I127795);
not I_7351 (I127868,I127846);
DFFARX1 I_7352 (I84039,I2859,I127769,I127894,);
nand I_7353 (I127902,I127894,I84036);
not I_7354 (I127919,I127902);
DFFARX1 I_7355 (I127919,I2859,I127769,I127945,);
not I_7356 (I127761,I127945);
nor I_7357 (I127967,I127795,I127902);
nor I_7358 (I127743,I127846,I127967);
DFFARX1 I_7359 (I84045,I2859,I127769,I128007,);
DFFARX1 I_7360 (I128007,I2859,I127769,I128024,);
not I_7361 (I128032,I128024);
not I_7362 (I128049,I128007);
nand I_7363 (I127746,I128049,I127868);
nand I_7364 (I128080,I84030,I84030);
and I_7365 (I128097,I128080,I84042);
DFFARX1 I_7366 (I128097,I2859,I127769,I128123,);
nor I_7367 (I128131,I128123,I127795);
DFFARX1 I_7368 (I128131,I2859,I127769,I127734,);
DFFARX1 I_7369 (I128123,I2859,I127769,I127752,);
nor I_7370 (I128176,I84048,I84030);
not I_7371 (I128193,I128176);
nor I_7372 (I127755,I128032,I128193);
nand I_7373 (I127740,I128049,I128193);
nor I_7374 (I127749,I127795,I128176);
DFFARX1 I_7375 (I128176,I2859,I127769,I127758,);
not I_7376 (I128296,I2866);
DFFARX1 I_7377 (I177284,I2859,I128296,I128322,);
nand I_7378 (I128330,I177296,I177275);
and I_7379 (I128347,I128330,I177299);
DFFARX1 I_7380 (I128347,I2859,I128296,I128373,);
nor I_7381 (I128264,I128373,I128322);
not I_7382 (I128395,I128373);
DFFARX1 I_7383 (I177290,I2859,I128296,I128421,);
nand I_7384 (I128429,I128421,I177272);
not I_7385 (I128446,I128429);
DFFARX1 I_7386 (I128446,I2859,I128296,I128472,);
not I_7387 (I128288,I128472);
nor I_7388 (I128494,I128322,I128429);
nor I_7389 (I128270,I128373,I128494);
DFFARX1 I_7390 (I177287,I2859,I128296,I128534,);
DFFARX1 I_7391 (I128534,I2859,I128296,I128551,);
not I_7392 (I128559,I128551);
not I_7393 (I128576,I128534);
nand I_7394 (I128273,I128576,I128395);
nand I_7395 (I128607,I177272,I177278);
and I_7396 (I128624,I128607,I177281);
DFFARX1 I_7397 (I128624,I2859,I128296,I128650,);
nor I_7398 (I128658,I128650,I128322);
DFFARX1 I_7399 (I128658,I2859,I128296,I128261,);
DFFARX1 I_7400 (I128650,I2859,I128296,I128279,);
nor I_7401 (I128703,I177293,I177278);
not I_7402 (I128720,I128703);
nor I_7403 (I128282,I128559,I128720);
nand I_7404 (I128267,I128576,I128720);
nor I_7405 (I128276,I128322,I128703);
DFFARX1 I_7406 (I128703,I2859,I128296,I128285,);
not I_7407 (I128823,I2866);
DFFARX1 I_7408 (I356013,I2859,I128823,I128849,);
nand I_7409 (I128857,I356016,I356010);
and I_7410 (I128874,I128857,I356022);
DFFARX1 I_7411 (I128874,I2859,I128823,I128900,);
nor I_7412 (I128791,I128900,I128849);
not I_7413 (I128922,I128900);
DFFARX1 I_7414 (I356025,I2859,I128823,I128948,);
nand I_7415 (I128956,I128948,I356016);
not I_7416 (I128973,I128956);
DFFARX1 I_7417 (I128973,I2859,I128823,I128999,);
not I_7418 (I128815,I128999);
nor I_7419 (I129021,I128849,I128956);
nor I_7420 (I128797,I128900,I129021);
DFFARX1 I_7421 (I356028,I2859,I128823,I129061,);
DFFARX1 I_7422 (I129061,I2859,I128823,I129078,);
not I_7423 (I129086,I129078);
not I_7424 (I129103,I129061);
nand I_7425 (I128800,I129103,I128922);
nand I_7426 (I129134,I356010,I356019);
and I_7427 (I129151,I129134,I356013);
DFFARX1 I_7428 (I129151,I2859,I128823,I129177,);
nor I_7429 (I129185,I129177,I128849);
DFFARX1 I_7430 (I129185,I2859,I128823,I128788,);
DFFARX1 I_7431 (I129177,I2859,I128823,I128806,);
nor I_7432 (I129230,I356031,I356019);
not I_7433 (I129247,I129230);
nor I_7434 (I128809,I129086,I129247);
nand I_7435 (I128794,I129103,I129247);
nor I_7436 (I128803,I128849,I129230);
DFFARX1 I_7437 (I129230,I2859,I128823,I128812,);
not I_7438 (I129350,I2866);
DFFARX1 I_7439 (I17438,I2859,I129350,I129376,);
nand I_7440 (I129384,I17462,I17441);
and I_7441 (I129401,I129384,I17438);
DFFARX1 I_7442 (I129401,I2859,I129350,I129427,);
nor I_7443 (I129318,I129427,I129376);
not I_7444 (I129449,I129427);
DFFARX1 I_7445 (I17444,I2859,I129350,I129475,);
nand I_7446 (I129483,I129475,I17453);
not I_7447 (I129500,I129483);
DFFARX1 I_7448 (I129500,I2859,I129350,I129526,);
not I_7449 (I129342,I129526);
nor I_7450 (I129548,I129376,I129483);
nor I_7451 (I129324,I129427,I129548);
DFFARX1 I_7452 (I17447,I2859,I129350,I129588,);
DFFARX1 I_7453 (I129588,I2859,I129350,I129605,);
not I_7454 (I129613,I129605);
not I_7455 (I129630,I129588);
nand I_7456 (I129327,I129630,I129449);
nand I_7457 (I129661,I17459,I17441);
and I_7458 (I129678,I129661,I17450);
DFFARX1 I_7459 (I129678,I2859,I129350,I129704,);
nor I_7460 (I129712,I129704,I129376);
DFFARX1 I_7461 (I129712,I2859,I129350,I129315,);
DFFARX1 I_7462 (I129704,I2859,I129350,I129333,);
nor I_7463 (I129757,I17456,I17441);
not I_7464 (I129774,I129757);
nor I_7465 (I129336,I129613,I129774);
nand I_7466 (I129321,I129630,I129774);
nor I_7467 (I129330,I129376,I129757);
DFFARX1 I_7468 (I129757,I2859,I129350,I129339,);
not I_7469 (I129877,I2866);
DFFARX1 I_7470 (I63797,I2859,I129877,I129903,);
nand I_7471 (I129911,I63797,I63803);
and I_7472 (I129928,I129911,I63821);
DFFARX1 I_7473 (I129928,I2859,I129877,I129954,);
nor I_7474 (I129845,I129954,I129903);
not I_7475 (I129976,I129954);
DFFARX1 I_7476 (I63809,I2859,I129877,I130002,);
nand I_7477 (I130010,I130002,I63806);
not I_7478 (I130027,I130010);
DFFARX1 I_7479 (I130027,I2859,I129877,I130053,);
not I_7480 (I129869,I130053);
nor I_7481 (I130075,I129903,I130010);
nor I_7482 (I129851,I129954,I130075);
DFFARX1 I_7483 (I63815,I2859,I129877,I130115,);
DFFARX1 I_7484 (I130115,I2859,I129877,I130132,);
not I_7485 (I130140,I130132);
not I_7486 (I130157,I130115);
nand I_7487 (I129854,I130157,I129976);
nand I_7488 (I130188,I63800,I63800);
and I_7489 (I130205,I130188,I63812);
DFFARX1 I_7490 (I130205,I2859,I129877,I130231,);
nor I_7491 (I130239,I130231,I129903);
DFFARX1 I_7492 (I130239,I2859,I129877,I129842,);
DFFARX1 I_7493 (I130231,I2859,I129877,I129860,);
nor I_7494 (I130284,I63818,I63800);
not I_7495 (I130301,I130284);
nor I_7496 (I129863,I130140,I130301);
nand I_7497 (I129848,I130157,I130301);
nor I_7498 (I129857,I129903,I130284);
DFFARX1 I_7499 (I130284,I2859,I129877,I129866,);
not I_7500 (I130404,I2866);
DFFARX1 I_7501 (I433295,I2859,I130404,I130430,);
nand I_7502 (I130438,I433292,I433295);
and I_7503 (I130455,I130438,I433304);
DFFARX1 I_7504 (I130455,I2859,I130404,I130481,);
nor I_7505 (I130372,I130481,I130430);
not I_7506 (I130503,I130481);
DFFARX1 I_7507 (I433292,I2859,I130404,I130529,);
nand I_7508 (I130537,I130529,I433310);
not I_7509 (I130554,I130537);
DFFARX1 I_7510 (I130554,I2859,I130404,I130580,);
not I_7511 (I130396,I130580);
nor I_7512 (I130602,I130430,I130537);
nor I_7513 (I130378,I130481,I130602);
DFFARX1 I_7514 (I433298,I2859,I130404,I130642,);
DFFARX1 I_7515 (I130642,I2859,I130404,I130659,);
not I_7516 (I130667,I130659);
not I_7517 (I130684,I130642);
nand I_7518 (I130381,I130684,I130503);
nand I_7519 (I130715,I433307,I433313);
and I_7520 (I130732,I130715,I433298);
DFFARX1 I_7521 (I130732,I2859,I130404,I130758,);
nor I_7522 (I130766,I130758,I130430);
DFFARX1 I_7523 (I130766,I2859,I130404,I130369,);
DFFARX1 I_7524 (I130758,I2859,I130404,I130387,);
nor I_7525 (I130811,I433301,I433313);
not I_7526 (I130828,I130811);
nor I_7527 (I130390,I130667,I130828);
nand I_7528 (I130375,I130684,I130828);
nor I_7529 (I130384,I130430,I130811);
DFFARX1 I_7530 (I130811,I2859,I130404,I130393,);
not I_7531 (I130931,I2866);
DFFARX1 I_7532 (I341257,I2859,I130931,I130957,);
nand I_7533 (I130965,I341260,I341254);
and I_7534 (I130982,I130965,I341266);
DFFARX1 I_7535 (I130982,I2859,I130931,I131008,);
nor I_7536 (I130899,I131008,I130957);
not I_7537 (I131030,I131008);
DFFARX1 I_7538 (I341269,I2859,I130931,I131056,);
nand I_7539 (I131064,I131056,I341260);
not I_7540 (I131081,I131064);
DFFARX1 I_7541 (I131081,I2859,I130931,I131107,);
not I_7542 (I130923,I131107);
nor I_7543 (I131129,I130957,I131064);
nor I_7544 (I130905,I131008,I131129);
DFFARX1 I_7545 (I341272,I2859,I130931,I131169,);
DFFARX1 I_7546 (I131169,I2859,I130931,I131186,);
not I_7547 (I131194,I131186);
not I_7548 (I131211,I131169);
nand I_7549 (I130908,I131211,I131030);
nand I_7550 (I131242,I341254,I341263);
and I_7551 (I131259,I131242,I341257);
DFFARX1 I_7552 (I131259,I2859,I130931,I131285,);
nor I_7553 (I131293,I131285,I130957);
DFFARX1 I_7554 (I131293,I2859,I130931,I130896,);
DFFARX1 I_7555 (I131285,I2859,I130931,I130914,);
nor I_7556 (I131338,I341275,I341263);
not I_7557 (I131355,I131338);
nor I_7558 (I130917,I131194,I131355);
nand I_7559 (I130902,I131211,I131355);
nor I_7560 (I130911,I130957,I131338);
DFFARX1 I_7561 (I131338,I2859,I130931,I130920,);
not I_7562 (I131458,I2866);
DFFARX1 I_7563 (I362456,I2859,I131458,I131484,);
nand I_7564 (I131492,I362453,I362471);
and I_7565 (I131509,I131492,I362462);
DFFARX1 I_7566 (I131509,I2859,I131458,I131535,);
nor I_7567 (I131426,I131535,I131484);
not I_7568 (I131557,I131535);
DFFARX1 I_7569 (I362477,I2859,I131458,I131583,);
nand I_7570 (I131591,I131583,I362459);
not I_7571 (I131608,I131591);
DFFARX1 I_7572 (I131608,I2859,I131458,I131634,);
not I_7573 (I131450,I131634);
nor I_7574 (I131656,I131484,I131591);
nor I_7575 (I131432,I131535,I131656);
DFFARX1 I_7576 (I362465,I2859,I131458,I131696,);
DFFARX1 I_7577 (I131696,I2859,I131458,I131713,);
not I_7578 (I131721,I131713);
not I_7579 (I131738,I131696);
nand I_7580 (I131435,I131738,I131557);
nand I_7581 (I131769,I362453,I362480);
and I_7582 (I131786,I131769,I362468);
DFFARX1 I_7583 (I131786,I2859,I131458,I131812,);
nor I_7584 (I131820,I131812,I131484);
DFFARX1 I_7585 (I131820,I2859,I131458,I131423,);
DFFARX1 I_7586 (I131812,I2859,I131458,I131441,);
nor I_7587 (I131865,I362474,I362480);
not I_7588 (I131882,I131865);
nor I_7589 (I131444,I131721,I131882);
nand I_7590 (I131429,I131738,I131882);
nor I_7591 (I131438,I131484,I131865);
DFFARX1 I_7592 (I131865,I2859,I131458,I131447,);
not I_7593 (I131985,I2866);
DFFARX1 I_7594 (I381836,I2859,I131985,I132011,);
nand I_7595 (I132019,I381833,I381851);
and I_7596 (I132036,I132019,I381842);
DFFARX1 I_7597 (I132036,I2859,I131985,I132062,);
nor I_7598 (I131953,I132062,I132011);
not I_7599 (I132084,I132062);
DFFARX1 I_7600 (I381857,I2859,I131985,I132110,);
nand I_7601 (I132118,I132110,I381839);
not I_7602 (I132135,I132118);
DFFARX1 I_7603 (I132135,I2859,I131985,I132161,);
not I_7604 (I131977,I132161);
nor I_7605 (I132183,I132011,I132118);
nor I_7606 (I131959,I132062,I132183);
DFFARX1 I_7607 (I381845,I2859,I131985,I132223,);
DFFARX1 I_7608 (I132223,I2859,I131985,I132240,);
not I_7609 (I132248,I132240);
not I_7610 (I132265,I132223);
nand I_7611 (I131962,I132265,I132084);
nand I_7612 (I132296,I381833,I381860);
and I_7613 (I132313,I132296,I381848);
DFFARX1 I_7614 (I132313,I2859,I131985,I132339,);
nor I_7615 (I132347,I132339,I132011);
DFFARX1 I_7616 (I132347,I2859,I131985,I131950,);
DFFARX1 I_7617 (I132339,I2859,I131985,I131968,);
nor I_7618 (I132392,I381854,I381860);
not I_7619 (I132409,I132392);
nor I_7620 (I131971,I132248,I132409);
nand I_7621 (I131956,I132265,I132409);
nor I_7622 (I131965,I132011,I132392);
DFFARX1 I_7623 (I132392,I2859,I131985,I131974,);
not I_7624 (I132512,I2866);
DFFARX1 I_7625 (I551106,I2859,I132512,I132538,);
nand I_7626 (I132546,I551085,I551085);
and I_7627 (I132563,I132546,I551112);
DFFARX1 I_7628 (I132563,I2859,I132512,I132589,);
nor I_7629 (I132480,I132589,I132538);
not I_7630 (I132611,I132589);
DFFARX1 I_7631 (I551100,I2859,I132512,I132637,);
nand I_7632 (I132645,I132637,I551103);
not I_7633 (I132662,I132645);
DFFARX1 I_7634 (I132662,I2859,I132512,I132688,);
not I_7635 (I132504,I132688);
nor I_7636 (I132710,I132538,I132645);
nor I_7637 (I132486,I132589,I132710);
DFFARX1 I_7638 (I551094,I2859,I132512,I132750,);
DFFARX1 I_7639 (I132750,I2859,I132512,I132767,);
not I_7640 (I132775,I132767);
not I_7641 (I132792,I132750);
nand I_7642 (I132489,I132792,I132611);
nand I_7643 (I132823,I551091,I551088);
and I_7644 (I132840,I132823,I551109);
DFFARX1 I_7645 (I132840,I2859,I132512,I132866,);
nor I_7646 (I132874,I132866,I132538);
DFFARX1 I_7647 (I132874,I2859,I132512,I132477,);
DFFARX1 I_7648 (I132866,I2859,I132512,I132495,);
nor I_7649 (I132919,I551097,I551088);
not I_7650 (I132936,I132919);
nor I_7651 (I132498,I132775,I132936);
nand I_7652 (I132483,I132792,I132936);
nor I_7653 (I132492,I132538,I132919);
DFFARX1 I_7654 (I132919,I2859,I132512,I132501,);
not I_7655 (I133039,I2866);
DFFARX1 I_7656 (I452196,I2859,I133039,I133065,);
nand I_7657 (I133073,I452211,I452196);
and I_7658 (I133090,I133073,I452214);
DFFARX1 I_7659 (I133090,I2859,I133039,I133116,);
nor I_7660 (I133007,I133116,I133065);
not I_7661 (I133138,I133116);
DFFARX1 I_7662 (I452220,I2859,I133039,I133164,);
nand I_7663 (I133172,I133164,I452202);
not I_7664 (I133189,I133172);
DFFARX1 I_7665 (I133189,I2859,I133039,I133215,);
not I_7666 (I133031,I133215);
nor I_7667 (I133237,I133065,I133172);
nor I_7668 (I133013,I133116,I133237);
DFFARX1 I_7669 (I452199,I2859,I133039,I133277,);
DFFARX1 I_7670 (I133277,I2859,I133039,I133294,);
not I_7671 (I133302,I133294);
not I_7672 (I133319,I133277);
nand I_7673 (I133016,I133319,I133138);
nand I_7674 (I133350,I452199,I452205);
and I_7675 (I133367,I133350,I452217);
DFFARX1 I_7676 (I133367,I2859,I133039,I133393,);
nor I_7677 (I133401,I133393,I133065);
DFFARX1 I_7678 (I133401,I2859,I133039,I133004,);
DFFARX1 I_7679 (I133393,I2859,I133039,I133022,);
nor I_7680 (I133446,I452208,I452205);
not I_7681 (I133463,I133446);
nor I_7682 (I133025,I133302,I133463);
nand I_7683 (I133010,I133319,I133463);
nor I_7684 (I133019,I133065,I133446);
DFFARX1 I_7685 (I133446,I2859,I133039,I133028,);
not I_7686 (I133566,I2866);
DFFARX1 I_7687 (I10587,I2859,I133566,I133592,);
nand I_7688 (I133600,I10611,I10590);
and I_7689 (I133617,I133600,I10587);
DFFARX1 I_7690 (I133617,I2859,I133566,I133643,);
nor I_7691 (I133534,I133643,I133592);
not I_7692 (I133665,I133643);
DFFARX1 I_7693 (I10593,I2859,I133566,I133691,);
nand I_7694 (I133699,I133691,I10602);
not I_7695 (I133716,I133699);
DFFARX1 I_7696 (I133716,I2859,I133566,I133742,);
not I_7697 (I133558,I133742);
nor I_7698 (I133764,I133592,I133699);
nor I_7699 (I133540,I133643,I133764);
DFFARX1 I_7700 (I10596,I2859,I133566,I133804,);
DFFARX1 I_7701 (I133804,I2859,I133566,I133821,);
not I_7702 (I133829,I133821);
not I_7703 (I133846,I133804);
nand I_7704 (I133543,I133846,I133665);
nand I_7705 (I133877,I10608,I10590);
and I_7706 (I133894,I133877,I10599);
DFFARX1 I_7707 (I133894,I2859,I133566,I133920,);
nor I_7708 (I133928,I133920,I133592);
DFFARX1 I_7709 (I133928,I2859,I133566,I133531,);
DFFARX1 I_7710 (I133920,I2859,I133566,I133549,);
nor I_7711 (I133973,I10605,I10590);
not I_7712 (I133990,I133973);
nor I_7713 (I133552,I133829,I133990);
nand I_7714 (I133537,I133846,I133990);
nor I_7715 (I133546,I133592,I133973);
DFFARX1 I_7716 (I133973,I2859,I133566,I133555,);
not I_7717 (I134093,I2866);
DFFARX1 I_7718 (I214403,I2859,I134093,I134119,);
nand I_7719 (I134127,I214403,I214415);
and I_7720 (I134144,I134127,I214400);
DFFARX1 I_7721 (I134144,I2859,I134093,I134170,);
nor I_7722 (I134061,I134170,I134119);
not I_7723 (I134192,I134170);
DFFARX1 I_7724 (I214424,I2859,I134093,I134218,);
nand I_7725 (I134226,I134218,I214421);
not I_7726 (I134243,I134226);
DFFARX1 I_7727 (I134243,I2859,I134093,I134269,);
not I_7728 (I134085,I134269);
nor I_7729 (I134291,I134119,I134226);
nor I_7730 (I134067,I134170,I134291);
DFFARX1 I_7731 (I214412,I2859,I134093,I134331,);
DFFARX1 I_7732 (I134331,I2859,I134093,I134348,);
not I_7733 (I134356,I134348);
not I_7734 (I134373,I134331);
nand I_7735 (I134070,I134373,I134192);
nand I_7736 (I134404,I214400,I214409);
and I_7737 (I134421,I134404,I214418);
DFFARX1 I_7738 (I134421,I2859,I134093,I134447,);
nor I_7739 (I134455,I134447,I134119);
DFFARX1 I_7740 (I134455,I2859,I134093,I134058,);
DFFARX1 I_7741 (I134447,I2859,I134093,I134076,);
nor I_7742 (I134500,I214406,I214409);
not I_7743 (I134517,I134500);
nor I_7744 (I134079,I134356,I134517);
nand I_7745 (I134064,I134373,I134517);
nor I_7746 (I134073,I134119,I134500);
DFFARX1 I_7747 (I134500,I2859,I134093,I134082,);
not I_7748 (I134620,I2866);
DFFARX1 I_7749 (I190884,I2859,I134620,I134646,);
nand I_7750 (I134654,I190896,I190875);
and I_7751 (I134671,I134654,I190899);
DFFARX1 I_7752 (I134671,I2859,I134620,I134697,);
nor I_7753 (I134588,I134697,I134646);
not I_7754 (I134719,I134697);
DFFARX1 I_7755 (I190890,I2859,I134620,I134745,);
nand I_7756 (I134753,I134745,I190872);
not I_7757 (I134770,I134753);
DFFARX1 I_7758 (I134770,I2859,I134620,I134796,);
not I_7759 (I134612,I134796);
nor I_7760 (I134818,I134646,I134753);
nor I_7761 (I134594,I134697,I134818);
DFFARX1 I_7762 (I190887,I2859,I134620,I134858,);
DFFARX1 I_7763 (I134858,I2859,I134620,I134875,);
not I_7764 (I134883,I134875);
not I_7765 (I134900,I134858);
nand I_7766 (I134597,I134900,I134719);
nand I_7767 (I134931,I190872,I190878);
and I_7768 (I134948,I134931,I190881);
DFFARX1 I_7769 (I134948,I2859,I134620,I134974,);
nor I_7770 (I134982,I134974,I134646);
DFFARX1 I_7771 (I134982,I2859,I134620,I134585,);
DFFARX1 I_7772 (I134974,I2859,I134620,I134603,);
nor I_7773 (I135027,I190893,I190878);
not I_7774 (I135044,I135027);
nor I_7775 (I134606,I134883,I135044);
nand I_7776 (I134591,I134900,I135044);
nor I_7777 (I134600,I134646,I135027);
DFFARX1 I_7778 (I135027,I2859,I134620,I134609,);
not I_7779 (I135147,I2866);
DFFARX1 I_7780 (I462022,I2859,I135147,I135173,);
nand I_7781 (I135181,I462037,I462022);
and I_7782 (I135198,I135181,I462040);
DFFARX1 I_7783 (I135198,I2859,I135147,I135224,);
nor I_7784 (I135115,I135224,I135173);
not I_7785 (I135246,I135224);
DFFARX1 I_7786 (I462046,I2859,I135147,I135272,);
nand I_7787 (I135280,I135272,I462028);
not I_7788 (I135297,I135280);
DFFARX1 I_7789 (I135297,I2859,I135147,I135323,);
not I_7790 (I135139,I135323);
nor I_7791 (I135345,I135173,I135280);
nor I_7792 (I135121,I135224,I135345);
DFFARX1 I_7793 (I462025,I2859,I135147,I135385,);
DFFARX1 I_7794 (I135385,I2859,I135147,I135402,);
not I_7795 (I135410,I135402);
not I_7796 (I135427,I135385);
nand I_7797 (I135124,I135427,I135246);
nand I_7798 (I135458,I462025,I462031);
and I_7799 (I135475,I135458,I462043);
DFFARX1 I_7800 (I135475,I2859,I135147,I135501,);
nor I_7801 (I135509,I135501,I135173);
DFFARX1 I_7802 (I135509,I2859,I135147,I135112,);
DFFARX1 I_7803 (I135501,I2859,I135147,I135130,);
nor I_7804 (I135554,I462034,I462031);
not I_7805 (I135571,I135554);
nor I_7806 (I135133,I135410,I135571);
nand I_7807 (I135118,I135427,I135571);
nor I_7808 (I135127,I135173,I135554);
DFFARX1 I_7809 (I135554,I2859,I135147,I135136,);
not I_7810 (I135674,I2866);
DFFARX1 I_7811 (I77482,I2859,I135674,I135700,);
nand I_7812 (I135708,I77482,I77488);
and I_7813 (I135725,I135708,I77506);
DFFARX1 I_7814 (I135725,I2859,I135674,I135751,);
nor I_7815 (I135642,I135751,I135700);
not I_7816 (I135773,I135751);
DFFARX1 I_7817 (I77494,I2859,I135674,I135799,);
nand I_7818 (I135807,I135799,I77491);
not I_7819 (I135824,I135807);
DFFARX1 I_7820 (I135824,I2859,I135674,I135850,);
not I_7821 (I135666,I135850);
nor I_7822 (I135872,I135700,I135807);
nor I_7823 (I135648,I135751,I135872);
DFFARX1 I_7824 (I77500,I2859,I135674,I135912,);
DFFARX1 I_7825 (I135912,I2859,I135674,I135929,);
not I_7826 (I135937,I135929);
not I_7827 (I135954,I135912);
nand I_7828 (I135651,I135954,I135773);
nand I_7829 (I135985,I77485,I77485);
and I_7830 (I136002,I135985,I77497);
DFFARX1 I_7831 (I136002,I2859,I135674,I136028,);
nor I_7832 (I136036,I136028,I135700);
DFFARX1 I_7833 (I136036,I2859,I135674,I135639,);
DFFARX1 I_7834 (I136028,I2859,I135674,I135657,);
nor I_7835 (I136081,I77503,I77485);
not I_7836 (I136098,I136081);
nor I_7837 (I135660,I135937,I136098);
nand I_7838 (I135645,I135954,I136098);
nor I_7839 (I135654,I135700,I136081);
DFFARX1 I_7840 (I136081,I2859,I135674,I135663,);
not I_7841 (I136201,I2866);
DFFARX1 I_7842 (I376668,I2859,I136201,I136227,);
nand I_7843 (I136235,I376665,I376683);
and I_7844 (I136252,I136235,I376674);
DFFARX1 I_7845 (I136252,I2859,I136201,I136278,);
nor I_7846 (I136169,I136278,I136227);
not I_7847 (I136300,I136278);
DFFARX1 I_7848 (I376689,I2859,I136201,I136326,);
nand I_7849 (I136334,I136326,I376671);
not I_7850 (I136351,I136334);
DFFARX1 I_7851 (I136351,I2859,I136201,I136377,);
not I_7852 (I136193,I136377);
nor I_7853 (I136399,I136227,I136334);
nor I_7854 (I136175,I136278,I136399);
DFFARX1 I_7855 (I376677,I2859,I136201,I136439,);
DFFARX1 I_7856 (I136439,I2859,I136201,I136456,);
not I_7857 (I136464,I136456);
not I_7858 (I136481,I136439);
nand I_7859 (I136178,I136481,I136300);
nand I_7860 (I136512,I376665,I376692);
and I_7861 (I136529,I136512,I376680);
DFFARX1 I_7862 (I136529,I2859,I136201,I136555,);
nor I_7863 (I136563,I136555,I136227);
DFFARX1 I_7864 (I136563,I2859,I136201,I136166,);
DFFARX1 I_7865 (I136555,I2859,I136201,I136184,);
nor I_7866 (I136608,I376686,I376692);
not I_7867 (I136625,I136608);
nor I_7868 (I136187,I136464,I136625);
nand I_7869 (I136172,I136481,I136625);
nor I_7870 (I136181,I136227,I136608);
DFFARX1 I_7871 (I136608,I2859,I136201,I136190,);
not I_7872 (I136728,I2866);
DFFARX1 I_7873 (I241207,I2859,I136728,I136754,);
nand I_7874 (I136762,I241192,I241195);
and I_7875 (I136779,I136762,I241210);
DFFARX1 I_7876 (I136779,I2859,I136728,I136805,);
nor I_7877 (I136696,I136805,I136754);
not I_7878 (I136827,I136805);
DFFARX1 I_7879 (I241204,I2859,I136728,I136853,);
nand I_7880 (I136861,I136853,I241195);
not I_7881 (I136878,I136861);
DFFARX1 I_7882 (I136878,I2859,I136728,I136904,);
not I_7883 (I136720,I136904);
nor I_7884 (I136926,I136754,I136861);
nor I_7885 (I136702,I136805,I136926);
DFFARX1 I_7886 (I241201,I2859,I136728,I136966,);
DFFARX1 I_7887 (I136966,I2859,I136728,I136983,);
not I_7888 (I136991,I136983);
not I_7889 (I137008,I136966);
nand I_7890 (I136705,I137008,I136827);
nand I_7891 (I137039,I241216,I241192);
and I_7892 (I137056,I137039,I241213);
DFFARX1 I_7893 (I137056,I2859,I136728,I137082,);
nor I_7894 (I137090,I137082,I136754);
DFFARX1 I_7895 (I137090,I2859,I136728,I136693,);
DFFARX1 I_7896 (I137082,I2859,I136728,I136711,);
nor I_7897 (I137135,I241198,I241192);
not I_7898 (I137152,I137135);
nor I_7899 (I136714,I136991,I137152);
nand I_7900 (I136699,I137008,I137152);
nor I_7901 (I136708,I136754,I137135);
DFFARX1 I_7902 (I137135,I2859,I136728,I136717,);
not I_7903 (I137255,I2866);
DFFARX1 I_7904 (I34832,I2859,I137255,I137281,);
nand I_7905 (I137289,I34844,I34853);
and I_7906 (I137306,I137289,I34832);
DFFARX1 I_7907 (I137306,I2859,I137255,I137332,);
nor I_7908 (I137223,I137332,I137281);
not I_7909 (I137354,I137332);
DFFARX1 I_7910 (I34847,I2859,I137255,I137380,);
nand I_7911 (I137388,I137380,I34835);
not I_7912 (I137405,I137388);
DFFARX1 I_7913 (I137405,I2859,I137255,I137431,);
not I_7914 (I137247,I137431);
nor I_7915 (I137453,I137281,I137388);
nor I_7916 (I137229,I137332,I137453);
DFFARX1 I_7917 (I34838,I2859,I137255,I137493,);
DFFARX1 I_7918 (I137493,I2859,I137255,I137510,);
not I_7919 (I137518,I137510);
not I_7920 (I137535,I137493);
nand I_7921 (I137232,I137535,I137354);
nand I_7922 (I137566,I34829,I34829);
and I_7923 (I137583,I137566,I34841);
DFFARX1 I_7924 (I137583,I2859,I137255,I137609,);
nor I_7925 (I137617,I137609,I137281);
DFFARX1 I_7926 (I137617,I2859,I137255,I137220,);
DFFARX1 I_7927 (I137609,I2859,I137255,I137238,);
nor I_7928 (I137662,I34850,I34829);
not I_7929 (I137679,I137662);
nor I_7930 (I137241,I137518,I137679);
nand I_7931 (I137226,I137535,I137679);
nor I_7932 (I137235,I137281,I137662);
DFFARX1 I_7933 (I137662,I2859,I137255,I137244,);
not I_7934 (I137782,I2866);
DFFARX1 I_7935 (I39575,I2859,I137782,I137808,);
nand I_7936 (I137816,I39587,I39596);
and I_7937 (I137833,I137816,I39575);
DFFARX1 I_7938 (I137833,I2859,I137782,I137859,);
nor I_7939 (I137750,I137859,I137808);
not I_7940 (I137881,I137859);
DFFARX1 I_7941 (I39590,I2859,I137782,I137907,);
nand I_7942 (I137915,I137907,I39578);
not I_7943 (I137932,I137915);
DFFARX1 I_7944 (I137932,I2859,I137782,I137958,);
not I_7945 (I137774,I137958);
nor I_7946 (I137980,I137808,I137915);
nor I_7947 (I137756,I137859,I137980);
DFFARX1 I_7948 (I39581,I2859,I137782,I138020,);
DFFARX1 I_7949 (I138020,I2859,I137782,I138037,);
not I_7950 (I138045,I138037);
not I_7951 (I138062,I138020);
nand I_7952 (I137759,I138062,I137881);
nand I_7953 (I138093,I39572,I39572);
and I_7954 (I138110,I138093,I39584);
DFFARX1 I_7955 (I138110,I2859,I137782,I138136,);
nor I_7956 (I138144,I138136,I137808);
DFFARX1 I_7957 (I138144,I2859,I137782,I137747,);
DFFARX1 I_7958 (I138136,I2859,I137782,I137765,);
nor I_7959 (I138189,I39593,I39572);
not I_7960 (I138206,I138189);
nor I_7961 (I137768,I138045,I138206);
nand I_7962 (I137753,I138062,I138206);
nor I_7963 (I137762,I137808,I138189);
DFFARX1 I_7964 (I138189,I2859,I137782,I137771,);
not I_7965 (I138309,I2866);
DFFARX1 I_7966 (I249877,I2859,I138309,I138335,);
nand I_7967 (I138343,I249862,I249865);
and I_7968 (I138360,I138343,I249880);
DFFARX1 I_7969 (I138360,I2859,I138309,I138386,);
nor I_7970 (I138277,I138386,I138335);
not I_7971 (I138408,I138386);
DFFARX1 I_7972 (I249874,I2859,I138309,I138434,);
nand I_7973 (I138442,I138434,I249865);
not I_7974 (I138459,I138442);
DFFARX1 I_7975 (I138459,I2859,I138309,I138485,);
not I_7976 (I138301,I138485);
nor I_7977 (I138507,I138335,I138442);
nor I_7978 (I138283,I138386,I138507);
DFFARX1 I_7979 (I249871,I2859,I138309,I138547,);
DFFARX1 I_7980 (I138547,I2859,I138309,I138564,);
not I_7981 (I138572,I138564);
not I_7982 (I138589,I138547);
nand I_7983 (I138286,I138589,I138408);
nand I_7984 (I138620,I249886,I249862);
and I_7985 (I138637,I138620,I249883);
DFFARX1 I_7986 (I138637,I2859,I138309,I138663,);
nor I_7987 (I138671,I138663,I138335);
DFFARX1 I_7988 (I138671,I2859,I138309,I138274,);
DFFARX1 I_7989 (I138663,I2859,I138309,I138292,);
nor I_7990 (I138716,I249868,I249862);
not I_7991 (I138733,I138716);
nor I_7992 (I138295,I138572,I138733);
nand I_7993 (I138280,I138589,I138733);
nor I_7994 (I138289,I138335,I138716);
DFFARX1 I_7995 (I138716,I2859,I138309,I138298,);
not I_7996 (I138836,I2866);
DFFARX1 I_7997 (I108422,I2859,I138836,I138862,);
nand I_7998 (I138870,I108422,I108428);
and I_7999 (I138887,I138870,I108446);
DFFARX1 I_8000 (I138887,I2859,I138836,I138913,);
nor I_8001 (I138804,I138913,I138862);
not I_8002 (I138935,I138913);
DFFARX1 I_8003 (I108434,I2859,I138836,I138961,);
nand I_8004 (I138969,I138961,I108431);
not I_8005 (I138986,I138969);
DFFARX1 I_8006 (I138986,I2859,I138836,I139012,);
not I_8007 (I138828,I139012);
nor I_8008 (I139034,I138862,I138969);
nor I_8009 (I138810,I138913,I139034);
DFFARX1 I_8010 (I108440,I2859,I138836,I139074,);
DFFARX1 I_8011 (I139074,I2859,I138836,I139091,);
not I_8012 (I139099,I139091);
not I_8013 (I139116,I139074);
nand I_8014 (I138813,I139116,I138935);
nand I_8015 (I139147,I108425,I108425);
and I_8016 (I139164,I139147,I108437);
DFFARX1 I_8017 (I139164,I2859,I138836,I139190,);
nor I_8018 (I139198,I139190,I138862);
DFFARX1 I_8019 (I139198,I2859,I138836,I138801,);
DFFARX1 I_8020 (I139190,I2859,I138836,I138819,);
nor I_8021 (I139243,I108443,I108425);
not I_8022 (I139260,I139243);
nor I_8023 (I138822,I139099,I139260);
nand I_8024 (I138807,I139116,I139260);
nor I_8025 (I138816,I138862,I139243);
DFFARX1 I_8026 (I139243,I2859,I138836,I138825,);
not I_8027 (I139363,I2866);
DFFARX1 I_8028 (I256813,I2859,I139363,I139389,);
nand I_8029 (I139397,I256798,I256801);
and I_8030 (I139414,I139397,I256816);
DFFARX1 I_8031 (I139414,I2859,I139363,I139440,);
nor I_8032 (I139331,I139440,I139389);
not I_8033 (I139462,I139440);
DFFARX1 I_8034 (I256810,I2859,I139363,I139488,);
nand I_8035 (I139496,I139488,I256801);
not I_8036 (I139513,I139496);
DFFARX1 I_8037 (I139513,I2859,I139363,I139539,);
not I_8038 (I139355,I139539);
nor I_8039 (I139561,I139389,I139496);
nor I_8040 (I139337,I139440,I139561);
DFFARX1 I_8041 (I256807,I2859,I139363,I139601,);
DFFARX1 I_8042 (I139601,I2859,I139363,I139618,);
not I_8043 (I139626,I139618);
not I_8044 (I139643,I139601);
nand I_8045 (I139340,I139643,I139462);
nand I_8046 (I139674,I256822,I256798);
and I_8047 (I139691,I139674,I256819);
DFFARX1 I_8048 (I139691,I2859,I139363,I139717,);
nor I_8049 (I139725,I139717,I139389);
DFFARX1 I_8050 (I139725,I2859,I139363,I139328,);
DFFARX1 I_8051 (I139717,I2859,I139363,I139346,);
nor I_8052 (I139770,I256804,I256798);
not I_8053 (I139787,I139770);
nor I_8054 (I139349,I139626,I139787);
nand I_8055 (I139334,I139643,I139787);
nor I_8056 (I139343,I139389,I139770);
DFFARX1 I_8057 (I139770,I2859,I139363,I139352,);
not I_8058 (I139890,I2866);
DFFARX1 I_8059 (I494968,I2859,I139890,I139916,);
nand I_8060 (I139924,I494983,I494968);
and I_8061 (I139941,I139924,I494986);
DFFARX1 I_8062 (I139941,I2859,I139890,I139967,);
nor I_8063 (I139858,I139967,I139916);
not I_8064 (I139989,I139967);
DFFARX1 I_8065 (I494992,I2859,I139890,I140015,);
nand I_8066 (I140023,I140015,I494974);
not I_8067 (I140040,I140023);
DFFARX1 I_8068 (I140040,I2859,I139890,I140066,);
not I_8069 (I139882,I140066);
nor I_8070 (I140088,I139916,I140023);
nor I_8071 (I139864,I139967,I140088);
DFFARX1 I_8072 (I494971,I2859,I139890,I140128,);
DFFARX1 I_8073 (I140128,I2859,I139890,I140145,);
not I_8074 (I140153,I140145);
not I_8075 (I140170,I140128);
nand I_8076 (I139867,I140170,I139989);
nand I_8077 (I140201,I494971,I494977);
and I_8078 (I140218,I140201,I494989);
DFFARX1 I_8079 (I140218,I2859,I139890,I140244,);
nor I_8080 (I140252,I140244,I139916);
DFFARX1 I_8081 (I140252,I2859,I139890,I139855,);
DFFARX1 I_8082 (I140244,I2859,I139890,I139873,);
nor I_8083 (I140297,I494980,I494977);
not I_8084 (I140314,I140297);
nor I_8085 (I139876,I140153,I140314);
nand I_8086 (I139861,I140170,I140314);
nor I_8087 (I139870,I139916,I140297);
DFFARX1 I_8088 (I140297,I2859,I139890,I139879,);
not I_8089 (I140417,I2866);
DFFARX1 I_8090 (I260856,I2859,I140417,I140443,);
nand I_8091 (I140451,I260847,I260862);
and I_8092 (I140468,I140451,I260868);
DFFARX1 I_8093 (I140468,I2859,I140417,I140494,);
nor I_8094 (I140385,I140494,I140443);
not I_8095 (I140516,I140494);
DFFARX1 I_8096 (I260853,I2859,I140417,I140542,);
nand I_8097 (I140550,I140542,I260847);
not I_8098 (I140567,I140550);
DFFARX1 I_8099 (I140567,I2859,I140417,I140593,);
not I_8100 (I140409,I140593);
nor I_8101 (I140615,I140443,I140550);
nor I_8102 (I140391,I140494,I140615);
DFFARX1 I_8103 (I260850,I2859,I140417,I140655,);
DFFARX1 I_8104 (I140655,I2859,I140417,I140672,);
not I_8105 (I140680,I140672);
not I_8106 (I140697,I140655);
nand I_8107 (I140394,I140697,I140516);
nand I_8108 (I140728,I260844,I260859);
and I_8109 (I140745,I140728,I260844);
DFFARX1 I_8110 (I140745,I2859,I140417,I140771,);
nor I_8111 (I140779,I140771,I140443);
DFFARX1 I_8112 (I140779,I2859,I140417,I140382,);
DFFARX1 I_8113 (I140771,I2859,I140417,I140400,);
nor I_8114 (I140824,I260865,I260859);
not I_8115 (I140841,I140824);
nor I_8116 (I140403,I140680,I140841);
nand I_8117 (I140388,I140697,I140841);
nor I_8118 (I140397,I140443,I140824);
DFFARX1 I_8119 (I140824,I2859,I140417,I140406,);
not I_8120 (I140944,I2866);
DFFARX1 I_8121 (I432734,I2859,I140944,I140970,);
nand I_8122 (I140978,I432731,I432734);
and I_8123 (I140995,I140978,I432743);
DFFARX1 I_8124 (I140995,I2859,I140944,I141021,);
nor I_8125 (I140912,I141021,I140970);
not I_8126 (I141043,I141021);
DFFARX1 I_8127 (I432731,I2859,I140944,I141069,);
nand I_8128 (I141077,I141069,I432749);
not I_8129 (I141094,I141077);
DFFARX1 I_8130 (I141094,I2859,I140944,I141120,);
not I_8131 (I140936,I141120);
nor I_8132 (I141142,I140970,I141077);
nor I_8133 (I140918,I141021,I141142);
DFFARX1 I_8134 (I432737,I2859,I140944,I141182,);
DFFARX1 I_8135 (I141182,I2859,I140944,I141199,);
not I_8136 (I141207,I141199);
not I_8137 (I141224,I141182);
nand I_8138 (I140921,I141224,I141043);
nand I_8139 (I141255,I432746,I432752);
and I_8140 (I141272,I141255,I432737);
DFFARX1 I_8141 (I141272,I2859,I140944,I141298,);
nor I_8142 (I141306,I141298,I140970);
DFFARX1 I_8143 (I141306,I2859,I140944,I140909,);
DFFARX1 I_8144 (I141298,I2859,I140944,I140927,);
nor I_8145 (I141351,I432740,I432752);
not I_8146 (I141368,I141351);
nor I_8147 (I140930,I141207,I141368);
nand I_8148 (I140915,I141224,I141368);
nor I_8149 (I140924,I140970,I141351);
DFFARX1 I_8150 (I141351,I2859,I140944,I140933,);
not I_8151 (I141471,I2866);
DFFARX1 I_8152 (I363748,I2859,I141471,I141497,);
nand I_8153 (I141505,I363745,I363763);
and I_8154 (I141522,I141505,I363754);
DFFARX1 I_8155 (I141522,I2859,I141471,I141548,);
nor I_8156 (I141439,I141548,I141497);
not I_8157 (I141570,I141548);
DFFARX1 I_8158 (I363769,I2859,I141471,I141596,);
nand I_8159 (I141604,I141596,I363751);
not I_8160 (I141621,I141604);
DFFARX1 I_8161 (I141621,I2859,I141471,I141647,);
not I_8162 (I141463,I141647);
nor I_8163 (I141669,I141497,I141604);
nor I_8164 (I141445,I141548,I141669);
DFFARX1 I_8165 (I363757,I2859,I141471,I141709,);
DFFARX1 I_8166 (I141709,I2859,I141471,I141726,);
not I_8167 (I141734,I141726);
not I_8168 (I141751,I141709);
nand I_8169 (I141448,I141751,I141570);
nand I_8170 (I141782,I363745,I363772);
and I_8171 (I141799,I141782,I363760);
DFFARX1 I_8172 (I141799,I2859,I141471,I141825,);
nor I_8173 (I141833,I141825,I141497);
DFFARX1 I_8174 (I141833,I2859,I141471,I141436,);
DFFARX1 I_8175 (I141825,I2859,I141471,I141454,);
nor I_8176 (I141878,I363766,I363772);
not I_8177 (I141895,I141878);
nor I_8178 (I141457,I141734,I141895);
nand I_8179 (I141442,I141751,I141895);
nor I_8180 (I141451,I141497,I141878);
DFFARX1 I_8181 (I141878,I2859,I141471,I141460,);
not I_8182 (I141998,I2866);
DFFARX1 I_8183 (I60227,I2859,I141998,I142024,);
nand I_8184 (I142032,I60227,I60233);
and I_8185 (I142049,I142032,I60251);
DFFARX1 I_8186 (I142049,I2859,I141998,I142075,);
nor I_8187 (I141966,I142075,I142024);
not I_8188 (I142097,I142075);
DFFARX1 I_8189 (I60239,I2859,I141998,I142123,);
nand I_8190 (I142131,I142123,I60236);
not I_8191 (I142148,I142131);
DFFARX1 I_8192 (I142148,I2859,I141998,I142174,);
not I_8193 (I141990,I142174);
nor I_8194 (I142196,I142024,I142131);
nor I_8195 (I141972,I142075,I142196);
DFFARX1 I_8196 (I60245,I2859,I141998,I142236,);
DFFARX1 I_8197 (I142236,I2859,I141998,I142253,);
not I_8198 (I142261,I142253);
not I_8199 (I142278,I142236);
nand I_8200 (I141975,I142278,I142097);
nand I_8201 (I142309,I60230,I60230);
and I_8202 (I142326,I142309,I60242);
DFFARX1 I_8203 (I142326,I2859,I141998,I142352,);
nor I_8204 (I142360,I142352,I142024);
DFFARX1 I_8205 (I142360,I2859,I141998,I141963,);
DFFARX1 I_8206 (I142352,I2859,I141998,I141981,);
nor I_8207 (I142405,I60248,I60230);
not I_8208 (I142422,I142405);
nor I_8209 (I141984,I142261,I142422);
nand I_8210 (I141969,I142278,I142422);
nor I_8211 (I141978,I142024,I142405);
DFFARX1 I_8212 (I142405,I2859,I141998,I141987,);
not I_8213 (I142525,I2866);
DFFARX1 I_8214 (I56657,I2859,I142525,I142551,);
nand I_8215 (I142559,I56657,I56663);
and I_8216 (I142576,I142559,I56681);
DFFARX1 I_8217 (I142576,I2859,I142525,I142602,);
nor I_8218 (I142493,I142602,I142551);
not I_8219 (I142624,I142602);
DFFARX1 I_8220 (I56669,I2859,I142525,I142650,);
nand I_8221 (I142658,I142650,I56666);
not I_8222 (I142675,I142658);
DFFARX1 I_8223 (I142675,I2859,I142525,I142701,);
not I_8224 (I142517,I142701);
nor I_8225 (I142723,I142551,I142658);
nor I_8226 (I142499,I142602,I142723);
DFFARX1 I_8227 (I56675,I2859,I142525,I142763,);
DFFARX1 I_8228 (I142763,I2859,I142525,I142780,);
not I_8229 (I142788,I142780);
not I_8230 (I142805,I142763);
nand I_8231 (I142502,I142805,I142624);
nand I_8232 (I142836,I56660,I56660);
and I_8233 (I142853,I142836,I56672);
DFFARX1 I_8234 (I142853,I2859,I142525,I142879,);
nor I_8235 (I142887,I142879,I142551);
DFFARX1 I_8236 (I142887,I2859,I142525,I142490,);
DFFARX1 I_8237 (I142879,I2859,I142525,I142508,);
nor I_8238 (I142932,I56678,I56660);
not I_8239 (I142949,I142932);
nor I_8240 (I142511,I142788,I142949);
nand I_8241 (I142496,I142805,I142949);
nor I_8242 (I142505,I142551,I142932);
DFFARX1 I_8243 (I142932,I2859,I142525,I142514,);
not I_8244 (I143052,I2866);
DFFARX1 I_8245 (I379252,I2859,I143052,I143078,);
nand I_8246 (I143086,I379249,I379267);
and I_8247 (I143103,I143086,I379258);
DFFARX1 I_8248 (I143103,I2859,I143052,I143129,);
nor I_8249 (I143020,I143129,I143078);
not I_8250 (I143151,I143129);
DFFARX1 I_8251 (I379273,I2859,I143052,I143177,);
nand I_8252 (I143185,I143177,I379255);
not I_8253 (I143202,I143185);
DFFARX1 I_8254 (I143202,I2859,I143052,I143228,);
not I_8255 (I143044,I143228);
nor I_8256 (I143250,I143078,I143185);
nor I_8257 (I143026,I143129,I143250);
DFFARX1 I_8258 (I379261,I2859,I143052,I143290,);
DFFARX1 I_8259 (I143290,I2859,I143052,I143307,);
not I_8260 (I143315,I143307);
not I_8261 (I143332,I143290);
nand I_8262 (I143029,I143332,I143151);
nand I_8263 (I143363,I379249,I379276);
and I_8264 (I143380,I143363,I379264);
DFFARX1 I_8265 (I143380,I2859,I143052,I143406,);
nor I_8266 (I143414,I143406,I143078);
DFFARX1 I_8267 (I143414,I2859,I143052,I143017,);
DFFARX1 I_8268 (I143406,I2859,I143052,I143035,);
nor I_8269 (I143459,I379270,I379276);
not I_8270 (I143476,I143459);
nor I_8271 (I143038,I143315,I143476);
nand I_8272 (I143023,I143332,I143476);
nor I_8273 (I143032,I143078,I143459);
DFFARX1 I_8274 (I143459,I2859,I143052,I143041,);
not I_8275 (I143579,I2866);
DFFARX1 I_8276 (I509572,I2859,I143579,I143605,);
nand I_8277 (I143613,I509554,I509578);
and I_8278 (I143630,I143613,I509569);
DFFARX1 I_8279 (I143630,I2859,I143579,I143656,);
nor I_8280 (I143547,I143656,I143605);
not I_8281 (I143678,I143656);
DFFARX1 I_8282 (I509575,I2859,I143579,I143704,);
nand I_8283 (I143712,I143704,I509563);
not I_8284 (I143729,I143712);
DFFARX1 I_8285 (I143729,I2859,I143579,I143755,);
not I_8286 (I143571,I143755);
nor I_8287 (I143777,I143605,I143712);
nor I_8288 (I143553,I143656,I143777);
DFFARX1 I_8289 (I509554,I2859,I143579,I143817,);
DFFARX1 I_8290 (I143817,I2859,I143579,I143834,);
not I_8291 (I143842,I143834);
not I_8292 (I143859,I143817);
nand I_8293 (I143556,I143859,I143678);
nand I_8294 (I143890,I509560,I509557);
and I_8295 (I143907,I143890,I509566);
DFFARX1 I_8296 (I143907,I2859,I143579,I143933,);
nor I_8297 (I143941,I143933,I143605);
DFFARX1 I_8298 (I143941,I2859,I143579,I143544,);
DFFARX1 I_8299 (I143933,I2859,I143579,I143562,);
nor I_8300 (I143986,I509557,I509557);
not I_8301 (I144003,I143986);
nor I_8302 (I143565,I143842,I144003);
nand I_8303 (I143550,I143859,I144003);
nor I_8304 (I143559,I143605,I143986);
DFFARX1 I_8305 (I143986,I2859,I143579,I143568,);
not I_8306 (I144106,I2866);
DFFARX1 I_8307 (I312298,I2859,I144106,I144132,);
nand I_8308 (I144140,I312289,I312304);
and I_8309 (I144157,I144140,I312310);
DFFARX1 I_8310 (I144157,I2859,I144106,I144183,);
nor I_8311 (I144074,I144183,I144132);
not I_8312 (I144205,I144183);
DFFARX1 I_8313 (I312295,I2859,I144106,I144231,);
nand I_8314 (I144239,I144231,I312289);
not I_8315 (I144256,I144239);
DFFARX1 I_8316 (I144256,I2859,I144106,I144282,);
not I_8317 (I144098,I144282);
nor I_8318 (I144304,I144132,I144239);
nor I_8319 (I144080,I144183,I144304);
DFFARX1 I_8320 (I312292,I2859,I144106,I144344,);
DFFARX1 I_8321 (I144344,I2859,I144106,I144361,);
not I_8322 (I144369,I144361);
not I_8323 (I144386,I144344);
nand I_8324 (I144083,I144386,I144205);
nand I_8325 (I144417,I312286,I312301);
and I_8326 (I144434,I144417,I312286);
DFFARX1 I_8327 (I144434,I2859,I144106,I144460,);
nor I_8328 (I144468,I144460,I144132);
DFFARX1 I_8329 (I144468,I2859,I144106,I144071,);
DFFARX1 I_8330 (I144460,I2859,I144106,I144089,);
nor I_8331 (I144513,I312307,I312301);
not I_8332 (I144530,I144513);
nor I_8333 (I144092,I144369,I144530);
nand I_8334 (I144077,I144386,I144530);
nor I_8335 (I144086,I144132,I144513);
DFFARX1 I_8336 (I144513,I2859,I144106,I144095,);
not I_8337 (I144633,I2866);
DFFARX1 I_8338 (I332825,I2859,I144633,I144659,);
nand I_8339 (I144667,I332828,I332822);
and I_8340 (I144684,I144667,I332834);
DFFARX1 I_8341 (I144684,I2859,I144633,I144710,);
nor I_8342 (I144601,I144710,I144659);
not I_8343 (I144732,I144710);
DFFARX1 I_8344 (I332837,I2859,I144633,I144758,);
nand I_8345 (I144766,I144758,I332828);
not I_8346 (I144783,I144766);
DFFARX1 I_8347 (I144783,I2859,I144633,I144809,);
not I_8348 (I144625,I144809);
nor I_8349 (I144831,I144659,I144766);
nor I_8350 (I144607,I144710,I144831);
DFFARX1 I_8351 (I332840,I2859,I144633,I144871,);
DFFARX1 I_8352 (I144871,I2859,I144633,I144888,);
not I_8353 (I144896,I144888);
not I_8354 (I144913,I144871);
nand I_8355 (I144610,I144913,I144732);
nand I_8356 (I144944,I332822,I332831);
and I_8357 (I144961,I144944,I332825);
DFFARX1 I_8358 (I144961,I2859,I144633,I144987,);
nor I_8359 (I144995,I144987,I144659);
DFFARX1 I_8360 (I144995,I2859,I144633,I144598,);
DFFARX1 I_8361 (I144987,I2859,I144633,I144616,);
nor I_8362 (I145040,I332843,I332831);
not I_8363 (I145057,I145040);
nor I_8364 (I144619,I144896,I145057);
nand I_8365 (I144604,I144913,I145057);
nor I_8366 (I144613,I144659,I145040);
DFFARX1 I_8367 (I145040,I2859,I144633,I144622,);
not I_8368 (I145160,I2866);
DFFARX1 I_8369 (I209048,I2859,I145160,I145186,);
nand I_8370 (I145194,I209048,I209060);
and I_8371 (I145211,I145194,I209045);
DFFARX1 I_8372 (I145211,I2859,I145160,I145237,);
nor I_8373 (I145128,I145237,I145186);
not I_8374 (I145259,I145237);
DFFARX1 I_8375 (I209069,I2859,I145160,I145285,);
nand I_8376 (I145293,I145285,I209066);
not I_8377 (I145310,I145293);
DFFARX1 I_8378 (I145310,I2859,I145160,I145336,);
not I_8379 (I145152,I145336);
nor I_8380 (I145358,I145186,I145293);
nor I_8381 (I145134,I145237,I145358);
DFFARX1 I_8382 (I209057,I2859,I145160,I145398,);
DFFARX1 I_8383 (I145398,I2859,I145160,I145415,);
not I_8384 (I145423,I145415);
not I_8385 (I145440,I145398);
nand I_8386 (I145137,I145440,I145259);
nand I_8387 (I145471,I209045,I209054);
and I_8388 (I145488,I145471,I209063);
DFFARX1 I_8389 (I145488,I2859,I145160,I145514,);
nor I_8390 (I145522,I145514,I145186);
DFFARX1 I_8391 (I145522,I2859,I145160,I145125,);
DFFARX1 I_8392 (I145514,I2859,I145160,I145143,);
nor I_8393 (I145567,I209051,I209054);
not I_8394 (I145584,I145567);
nor I_8395 (I145146,I145423,I145584);
nand I_8396 (I145131,I145440,I145584);
nor I_8397 (I145140,I145186,I145567);
DFFARX1 I_8398 (I145567,I2859,I145160,I145149,);
not I_8399 (I145687,I2866);
DFFARX1 I_8400 (I308830,I2859,I145687,I145713,);
nand I_8401 (I145721,I308821,I308836);
and I_8402 (I145738,I145721,I308842);
DFFARX1 I_8403 (I145738,I2859,I145687,I145764,);
nor I_8404 (I145655,I145764,I145713);
not I_8405 (I145786,I145764);
DFFARX1 I_8406 (I308827,I2859,I145687,I145812,);
nand I_8407 (I145820,I145812,I308821);
not I_8408 (I145837,I145820);
DFFARX1 I_8409 (I145837,I2859,I145687,I145863,);
not I_8410 (I145679,I145863);
nor I_8411 (I145885,I145713,I145820);
nor I_8412 (I145661,I145764,I145885);
DFFARX1 I_8413 (I308824,I2859,I145687,I145925,);
DFFARX1 I_8414 (I145925,I2859,I145687,I145942,);
not I_8415 (I145950,I145942);
not I_8416 (I145967,I145925);
nand I_8417 (I145664,I145967,I145786);
nand I_8418 (I145998,I308818,I308833);
and I_8419 (I146015,I145998,I308818);
DFFARX1 I_8420 (I146015,I2859,I145687,I146041,);
nor I_8421 (I146049,I146041,I145713);
DFFARX1 I_8422 (I146049,I2859,I145687,I145652,);
DFFARX1 I_8423 (I146041,I2859,I145687,I145670,);
nor I_8424 (I146094,I308839,I308833);
not I_8425 (I146111,I146094);
nor I_8426 (I145673,I145950,I146111);
nand I_8427 (I145658,I145967,I146111);
nor I_8428 (I145667,I145713,I146094);
DFFARX1 I_8429 (I146094,I2859,I145687,I145676,);
not I_8430 (I146214,I2866);
DFFARX1 I_8431 (I53111,I2859,I146214,I146240,);
nand I_8432 (I146248,I53096,I53087);
and I_8433 (I146265,I146248,I53102);
DFFARX1 I_8434 (I146265,I2859,I146214,I146291,);
nor I_8435 (I146182,I146291,I146240);
not I_8436 (I146313,I146291);
DFFARX1 I_8437 (I53114,I2859,I146214,I146339,);
nand I_8438 (I146347,I146339,I53105);
not I_8439 (I146364,I146347);
DFFARX1 I_8440 (I146364,I2859,I146214,I146390,);
not I_8441 (I146206,I146390);
nor I_8442 (I146412,I146240,I146347);
nor I_8443 (I146188,I146291,I146412);
DFFARX1 I_8444 (I53093,I2859,I146214,I146452,);
DFFARX1 I_8445 (I146452,I2859,I146214,I146469,);
not I_8446 (I146477,I146469);
not I_8447 (I146494,I146452);
nand I_8448 (I146191,I146494,I146313);
nand I_8449 (I146525,I53099,I53090);
and I_8450 (I146542,I146525,I53087);
DFFARX1 I_8451 (I146542,I2859,I146214,I146568,);
nor I_8452 (I146576,I146568,I146240);
DFFARX1 I_8453 (I146576,I2859,I146214,I146179,);
DFFARX1 I_8454 (I146568,I2859,I146214,I146197,);
nor I_8455 (I146621,I53108,I53090);
not I_8456 (I146638,I146621);
nor I_8457 (I146200,I146477,I146638);
nand I_8458 (I146185,I146494,I146638);
nor I_8459 (I146194,I146240,I146621);
DFFARX1 I_8460 (I146621,I2859,I146214,I146203,);
not I_8461 (I146741,I2866);
DFFARX1 I_8462 (I556461,I2859,I146741,I146767,);
nand I_8463 (I146775,I556440,I556440);
and I_8464 (I146792,I146775,I556467);
DFFARX1 I_8465 (I146792,I2859,I146741,I146818,);
nor I_8466 (I146709,I146818,I146767);
not I_8467 (I146840,I146818);
DFFARX1 I_8468 (I556455,I2859,I146741,I146866,);
nand I_8469 (I146874,I146866,I556458);
not I_8470 (I146891,I146874);
DFFARX1 I_8471 (I146891,I2859,I146741,I146917,);
not I_8472 (I146733,I146917);
nor I_8473 (I146939,I146767,I146874);
nor I_8474 (I146715,I146818,I146939);
DFFARX1 I_8475 (I556449,I2859,I146741,I146979,);
DFFARX1 I_8476 (I146979,I2859,I146741,I146996,);
not I_8477 (I147004,I146996);
not I_8478 (I147021,I146979);
nand I_8479 (I146718,I147021,I146840);
nand I_8480 (I147052,I556446,I556443);
and I_8481 (I147069,I147052,I556464);
DFFARX1 I_8482 (I147069,I2859,I146741,I147095,);
nor I_8483 (I147103,I147095,I146767);
DFFARX1 I_8484 (I147103,I2859,I146741,I146706,);
DFFARX1 I_8485 (I147095,I2859,I146741,I146724,);
nor I_8486 (I147148,I556452,I556443);
not I_8487 (I147165,I147148);
nor I_8488 (I146727,I147004,I147165);
nand I_8489 (I146712,I147021,I147165);
nor I_8490 (I146721,I146767,I147148);
DFFARX1 I_8491 (I147148,I2859,I146741,I146730,);
not I_8492 (I147268,I2866);
DFFARX1 I_8493 (I254501,I2859,I147268,I147294,);
nand I_8494 (I147302,I254486,I254489);
and I_8495 (I147319,I147302,I254504);
DFFARX1 I_8496 (I147319,I2859,I147268,I147345,);
nor I_8497 (I147236,I147345,I147294);
not I_8498 (I147367,I147345);
DFFARX1 I_8499 (I254498,I2859,I147268,I147393,);
nand I_8500 (I147401,I147393,I254489);
not I_8501 (I147418,I147401);
DFFARX1 I_8502 (I147418,I2859,I147268,I147444,);
not I_8503 (I147260,I147444);
nor I_8504 (I147466,I147294,I147401);
nor I_8505 (I147242,I147345,I147466);
DFFARX1 I_8506 (I254495,I2859,I147268,I147506,);
DFFARX1 I_8507 (I147506,I2859,I147268,I147523,);
not I_8508 (I147531,I147523);
not I_8509 (I147548,I147506);
nand I_8510 (I147245,I147548,I147367);
nand I_8511 (I147579,I254510,I254486);
and I_8512 (I147596,I147579,I254507);
DFFARX1 I_8513 (I147596,I2859,I147268,I147622,);
nor I_8514 (I147630,I147622,I147294);
DFFARX1 I_8515 (I147630,I2859,I147268,I147233,);
DFFARX1 I_8516 (I147622,I2859,I147268,I147251,);
nor I_8517 (I147675,I254492,I254486);
not I_8518 (I147692,I147675);
nor I_8519 (I147254,I147531,I147692);
nand I_8520 (I147239,I147548,I147692);
nor I_8521 (I147248,I147294,I147675);
DFFARX1 I_8522 (I147675,I2859,I147268,I147257,);
not I_8523 (I147795,I2866);
DFFARX1 I_8524 (I270682,I2859,I147795,I147821,);
nand I_8525 (I147829,I270673,I270688);
and I_8526 (I147846,I147829,I270694);
DFFARX1 I_8527 (I147846,I2859,I147795,I147872,);
nor I_8528 (I147763,I147872,I147821);
not I_8529 (I147894,I147872);
DFFARX1 I_8530 (I270679,I2859,I147795,I147920,);
nand I_8531 (I147928,I147920,I270673);
not I_8532 (I147945,I147928);
DFFARX1 I_8533 (I147945,I2859,I147795,I147971,);
not I_8534 (I147787,I147971);
nor I_8535 (I147993,I147821,I147928);
nor I_8536 (I147769,I147872,I147993);
DFFARX1 I_8537 (I270676,I2859,I147795,I148033,);
DFFARX1 I_8538 (I148033,I2859,I147795,I148050,);
not I_8539 (I148058,I148050);
not I_8540 (I148075,I148033);
nand I_8541 (I147772,I148075,I147894);
nand I_8542 (I148106,I270670,I270685);
and I_8543 (I148123,I148106,I270670);
DFFARX1 I_8544 (I148123,I2859,I147795,I148149,);
nor I_8545 (I148157,I148149,I147821);
DFFARX1 I_8546 (I148157,I2859,I147795,I147760,);
DFFARX1 I_8547 (I148149,I2859,I147795,I147778,);
nor I_8548 (I148202,I270691,I270685);
not I_8549 (I148219,I148202);
nor I_8550 (I147781,I148058,I148219);
nand I_8551 (I147766,I148075,I148219);
nor I_8552 (I147775,I147821,I148202);
DFFARX1 I_8553 (I148202,I2859,I147795,I147784,);
not I_8554 (I148322,I2866);
DFFARX1 I_8555 (I76292,I2859,I148322,I148348,);
nand I_8556 (I148356,I76292,I76298);
and I_8557 (I148373,I148356,I76316);
DFFARX1 I_8558 (I148373,I2859,I148322,I148399,);
nor I_8559 (I148290,I148399,I148348);
not I_8560 (I148421,I148399);
DFFARX1 I_8561 (I76304,I2859,I148322,I148447,);
nand I_8562 (I148455,I148447,I76301);
not I_8563 (I148472,I148455);
DFFARX1 I_8564 (I148472,I2859,I148322,I148498,);
not I_8565 (I148314,I148498);
nor I_8566 (I148520,I148348,I148455);
nor I_8567 (I148296,I148399,I148520);
DFFARX1 I_8568 (I76310,I2859,I148322,I148560,);
DFFARX1 I_8569 (I148560,I2859,I148322,I148577,);
not I_8570 (I148585,I148577);
not I_8571 (I148602,I148560);
nand I_8572 (I148299,I148602,I148421);
nand I_8573 (I148633,I76295,I76295);
and I_8574 (I148650,I148633,I76307);
DFFARX1 I_8575 (I148650,I2859,I148322,I148676,);
nor I_8576 (I148684,I148676,I148348);
DFFARX1 I_8577 (I148684,I2859,I148322,I148287,);
DFFARX1 I_8578 (I148676,I2859,I148322,I148305,);
nor I_8579 (I148729,I76313,I76295);
not I_8580 (I148746,I148729);
nor I_8581 (I148308,I148585,I148746);
nand I_8582 (I148293,I148602,I148746);
nor I_8583 (I148302,I148348,I148729);
DFFARX1 I_8584 (I148729,I2859,I148322,I148311,);
not I_8585 (I148849,I2866);
DFFARX1 I_8586 (I24819,I2859,I148849,I148875,);
nand I_8587 (I148883,I24831,I24840);
and I_8588 (I148900,I148883,I24819);
DFFARX1 I_8589 (I148900,I2859,I148849,I148926,);
nor I_8590 (I148817,I148926,I148875);
not I_8591 (I148948,I148926);
DFFARX1 I_8592 (I24834,I2859,I148849,I148974,);
nand I_8593 (I148982,I148974,I24822);
not I_8594 (I148999,I148982);
DFFARX1 I_8595 (I148999,I2859,I148849,I149025,);
not I_8596 (I148841,I149025);
nor I_8597 (I149047,I148875,I148982);
nor I_8598 (I148823,I148926,I149047);
DFFARX1 I_8599 (I24825,I2859,I148849,I149087,);
DFFARX1 I_8600 (I149087,I2859,I148849,I149104,);
not I_8601 (I149112,I149104);
not I_8602 (I149129,I149087);
nand I_8603 (I148826,I149129,I148948);
nand I_8604 (I149160,I24816,I24816);
and I_8605 (I149177,I149160,I24828);
DFFARX1 I_8606 (I149177,I2859,I148849,I149203,);
nor I_8607 (I149211,I149203,I148875);
DFFARX1 I_8608 (I149211,I2859,I148849,I148814,);
DFFARX1 I_8609 (I149203,I2859,I148849,I148832,);
nor I_8610 (I149256,I24837,I24816);
not I_8611 (I149273,I149256);
nor I_8612 (I148835,I149112,I149273);
nand I_8613 (I148820,I149129,I149273);
nor I_8614 (I148829,I148875,I149256);
DFFARX1 I_8615 (I149256,I2859,I148849,I148838,);
not I_8616 (I149376,I2866);
DFFARX1 I_8617 (I324920,I2859,I149376,I149402,);
nand I_8618 (I149410,I324923,I324917);
and I_8619 (I149427,I149410,I324929);
DFFARX1 I_8620 (I149427,I2859,I149376,I149453,);
nor I_8621 (I149344,I149453,I149402);
not I_8622 (I149475,I149453);
DFFARX1 I_8623 (I324932,I2859,I149376,I149501,);
nand I_8624 (I149509,I149501,I324923);
not I_8625 (I149526,I149509);
DFFARX1 I_8626 (I149526,I2859,I149376,I149552,);
not I_8627 (I149368,I149552);
nor I_8628 (I149574,I149402,I149509);
nor I_8629 (I149350,I149453,I149574);
DFFARX1 I_8630 (I324935,I2859,I149376,I149614,);
DFFARX1 I_8631 (I149614,I2859,I149376,I149631,);
not I_8632 (I149639,I149631);
not I_8633 (I149656,I149614);
nand I_8634 (I149353,I149656,I149475);
nand I_8635 (I149687,I324917,I324926);
and I_8636 (I149704,I149687,I324920);
DFFARX1 I_8637 (I149704,I2859,I149376,I149730,);
nor I_8638 (I149738,I149730,I149402);
DFFARX1 I_8639 (I149738,I2859,I149376,I149341,);
DFFARX1 I_8640 (I149730,I2859,I149376,I149359,);
nor I_8641 (I149783,I324938,I324926);
not I_8642 (I149800,I149783);
nor I_8643 (I149362,I149639,I149800);
nand I_8644 (I149347,I149656,I149800);
nor I_8645 (I149356,I149402,I149783);
DFFARX1 I_8646 (I149783,I2859,I149376,I149365,);
not I_8647 (I149903,I2866);
DFFARX1 I_8648 (I374084,I2859,I149903,I149929,);
nand I_8649 (I149937,I374081,I374099);
and I_8650 (I149954,I149937,I374090);
DFFARX1 I_8651 (I149954,I2859,I149903,I149980,);
nor I_8652 (I149871,I149980,I149929);
not I_8653 (I150002,I149980);
DFFARX1 I_8654 (I374105,I2859,I149903,I150028,);
nand I_8655 (I150036,I150028,I374087);
not I_8656 (I150053,I150036);
DFFARX1 I_8657 (I150053,I2859,I149903,I150079,);
not I_8658 (I149895,I150079);
nor I_8659 (I150101,I149929,I150036);
nor I_8660 (I149877,I149980,I150101);
DFFARX1 I_8661 (I374093,I2859,I149903,I150141,);
DFFARX1 I_8662 (I150141,I2859,I149903,I150158,);
not I_8663 (I150166,I150158);
not I_8664 (I150183,I150141);
nand I_8665 (I149880,I150183,I150002);
nand I_8666 (I150214,I374081,I374108);
and I_8667 (I150231,I150214,I374096);
DFFARX1 I_8668 (I150231,I2859,I149903,I150257,);
nor I_8669 (I150265,I150257,I149929);
DFFARX1 I_8670 (I150265,I2859,I149903,I149868,);
DFFARX1 I_8671 (I150257,I2859,I149903,I149886,);
nor I_8672 (I150310,I374102,I374108);
not I_8673 (I150327,I150310);
nor I_8674 (I149889,I150166,I150327);
nand I_8675 (I149874,I150183,I150327);
nor I_8676 (I149883,I149929,I150310);
DFFARX1 I_8677 (I150310,I2859,I149903,I149892,);
not I_8678 (I150430,I2866);
DFFARX1 I_8679 (I353905,I2859,I150430,I150456,);
nand I_8680 (I150464,I353908,I353902);
and I_8681 (I150481,I150464,I353914);
DFFARX1 I_8682 (I150481,I2859,I150430,I150507,);
nor I_8683 (I150398,I150507,I150456);
not I_8684 (I150529,I150507);
DFFARX1 I_8685 (I353917,I2859,I150430,I150555,);
nand I_8686 (I150563,I150555,I353908);
not I_8687 (I150580,I150563);
DFFARX1 I_8688 (I150580,I2859,I150430,I150606,);
not I_8689 (I150422,I150606);
nor I_8690 (I150628,I150456,I150563);
nor I_8691 (I150404,I150507,I150628);
DFFARX1 I_8692 (I353920,I2859,I150430,I150668,);
DFFARX1 I_8693 (I150668,I2859,I150430,I150685,);
not I_8694 (I150693,I150685);
not I_8695 (I150710,I150668);
nand I_8696 (I150407,I150710,I150529);
nand I_8697 (I150741,I353902,I353911);
and I_8698 (I150758,I150741,I353905);
DFFARX1 I_8699 (I150758,I2859,I150430,I150784,);
nor I_8700 (I150792,I150784,I150456);
DFFARX1 I_8701 (I150792,I2859,I150430,I150395,);
DFFARX1 I_8702 (I150784,I2859,I150430,I150413,);
nor I_8703 (I150837,I353923,I353911);
not I_8704 (I150854,I150837);
nor I_8705 (I150416,I150693,I150854);
nand I_8706 (I150401,I150710,I150854);
nor I_8707 (I150410,I150456,I150837);
DFFARX1 I_8708 (I150837,I2859,I150430,I150419,);
not I_8709 (I150957,I2866);
DFFARX1 I_8710 (I478784,I2859,I150957,I150983,);
nand I_8711 (I150991,I478799,I478784);
and I_8712 (I151008,I150991,I478802);
DFFARX1 I_8713 (I151008,I2859,I150957,I151034,);
nor I_8714 (I150925,I151034,I150983);
not I_8715 (I151056,I151034);
DFFARX1 I_8716 (I478808,I2859,I150957,I151082,);
nand I_8717 (I151090,I151082,I478790);
not I_8718 (I151107,I151090);
DFFARX1 I_8719 (I151107,I2859,I150957,I151133,);
not I_8720 (I150949,I151133);
nor I_8721 (I151155,I150983,I151090);
nor I_8722 (I150931,I151034,I151155);
DFFARX1 I_8723 (I478787,I2859,I150957,I151195,);
DFFARX1 I_8724 (I151195,I2859,I150957,I151212,);
not I_8725 (I151220,I151212);
not I_8726 (I151237,I151195);
nand I_8727 (I150934,I151237,I151056);
nand I_8728 (I151268,I478787,I478793);
and I_8729 (I151285,I151268,I478805);
DFFARX1 I_8730 (I151285,I2859,I150957,I151311,);
nor I_8731 (I151319,I151311,I150983);
DFFARX1 I_8732 (I151319,I2859,I150957,I150922,);
DFFARX1 I_8733 (I151311,I2859,I150957,I150940,);
nor I_8734 (I151364,I478796,I478793);
not I_8735 (I151381,I151364);
nor I_8736 (I150943,I151220,I151381);
nand I_8737 (I150928,I151237,I151381);
nor I_8738 (I150937,I150983,I151364);
DFFARX1 I_8739 (I151364,I2859,I150957,I150946,);
not I_8740 (I151484,I2866);
DFFARX1 I_8741 (I264324,I2859,I151484,I151510,);
nand I_8742 (I151518,I264315,I264330);
and I_8743 (I151535,I151518,I264336);
DFFARX1 I_8744 (I151535,I2859,I151484,I151561,);
nor I_8745 (I151452,I151561,I151510);
not I_8746 (I151583,I151561);
DFFARX1 I_8747 (I264321,I2859,I151484,I151609,);
nand I_8748 (I151617,I151609,I264315);
not I_8749 (I151634,I151617);
DFFARX1 I_8750 (I151634,I2859,I151484,I151660,);
not I_8751 (I151476,I151660);
nor I_8752 (I151682,I151510,I151617);
nor I_8753 (I151458,I151561,I151682);
DFFARX1 I_8754 (I264318,I2859,I151484,I151722,);
DFFARX1 I_8755 (I151722,I2859,I151484,I151739,);
not I_8756 (I151747,I151739);
not I_8757 (I151764,I151722);
nand I_8758 (I151461,I151764,I151583);
nand I_8759 (I151795,I264312,I264327);
and I_8760 (I151812,I151795,I264312);
DFFARX1 I_8761 (I151812,I2859,I151484,I151838,);
nor I_8762 (I151846,I151838,I151510);
DFFARX1 I_8763 (I151846,I2859,I151484,I151449,);
DFFARX1 I_8764 (I151838,I2859,I151484,I151467,);
nor I_8765 (I151891,I264333,I264327);
not I_8766 (I151908,I151891);
nor I_8767 (I151470,I151747,I151908);
nand I_8768 (I151455,I151764,I151908);
nor I_8769 (I151464,I151510,I151891);
DFFARX1 I_8770 (I151891,I2859,I151484,I151473,);
not I_8771 (I152011,I2866);
DFFARX1 I_8772 (I169668,I2859,I152011,I152037,);
nand I_8773 (I152045,I169680,I169659);
and I_8774 (I152062,I152045,I169683);
DFFARX1 I_8775 (I152062,I2859,I152011,I152088,);
nor I_8776 (I151979,I152088,I152037);
not I_8777 (I152110,I152088);
DFFARX1 I_8778 (I169674,I2859,I152011,I152136,);
nand I_8779 (I152144,I152136,I169656);
not I_8780 (I152161,I152144);
DFFARX1 I_8781 (I152161,I2859,I152011,I152187,);
not I_8782 (I152003,I152187);
nor I_8783 (I152209,I152037,I152144);
nor I_8784 (I151985,I152088,I152209);
DFFARX1 I_8785 (I169671,I2859,I152011,I152249,);
DFFARX1 I_8786 (I152249,I2859,I152011,I152266,);
not I_8787 (I152274,I152266);
not I_8788 (I152291,I152249);
nand I_8789 (I151988,I152291,I152110);
nand I_8790 (I152322,I169656,I169662);
and I_8791 (I152339,I152322,I169665);
DFFARX1 I_8792 (I152339,I2859,I152011,I152365,);
nor I_8793 (I152373,I152365,I152037);
DFFARX1 I_8794 (I152373,I2859,I152011,I151976,);
DFFARX1 I_8795 (I152365,I2859,I152011,I151994,);
nor I_8796 (I152418,I169677,I169662);
not I_8797 (I152435,I152418);
nor I_8798 (I151997,I152274,I152435);
nand I_8799 (I151982,I152291,I152435);
nor I_8800 (I151991,I152037,I152418);
DFFARX1 I_8801 (I152418,I2859,I152011,I152000,);
not I_8802 (I152538,I2866);
DFFARX1 I_8803 (I229069,I2859,I152538,I152564,);
nand I_8804 (I152572,I229054,I229057);
and I_8805 (I152589,I152572,I229072);
DFFARX1 I_8806 (I152589,I2859,I152538,I152615,);
nor I_8807 (I152506,I152615,I152564);
not I_8808 (I152637,I152615);
DFFARX1 I_8809 (I229066,I2859,I152538,I152663,);
nand I_8810 (I152671,I152663,I229057);
not I_8811 (I152688,I152671);
DFFARX1 I_8812 (I152688,I2859,I152538,I152714,);
not I_8813 (I152530,I152714);
nor I_8814 (I152736,I152564,I152671);
nor I_8815 (I152512,I152615,I152736);
DFFARX1 I_8816 (I229063,I2859,I152538,I152776,);
DFFARX1 I_8817 (I152776,I2859,I152538,I152793,);
not I_8818 (I152801,I152793);
not I_8819 (I152818,I152776);
nand I_8820 (I152515,I152818,I152637);
nand I_8821 (I152849,I229078,I229054);
and I_8822 (I152866,I152849,I229075);
DFFARX1 I_8823 (I152866,I2859,I152538,I152892,);
nor I_8824 (I152900,I152892,I152564);
DFFARX1 I_8825 (I152900,I2859,I152538,I152503,);
DFFARX1 I_8826 (I152892,I2859,I152538,I152521,);
nor I_8827 (I152945,I229060,I229054);
not I_8828 (I152962,I152945);
nor I_8829 (I152524,I152801,I152962);
nand I_8830 (I152509,I152818,I152962);
nor I_8831 (I152518,I152564,I152945);
DFFARX1 I_8832 (I152945,I2859,I152538,I152527,);
not I_8833 (I153065,I2866);
DFFARX1 I_8834 (I74507,I2859,I153065,I153091,);
nand I_8835 (I153099,I74507,I74513);
and I_8836 (I153116,I153099,I74531);
DFFARX1 I_8837 (I153116,I2859,I153065,I153142,);
nor I_8838 (I153033,I153142,I153091);
not I_8839 (I153164,I153142);
DFFARX1 I_8840 (I74519,I2859,I153065,I153190,);
nand I_8841 (I153198,I153190,I74516);
not I_8842 (I153215,I153198);
DFFARX1 I_8843 (I153215,I2859,I153065,I153241,);
not I_8844 (I153057,I153241);
nor I_8845 (I153263,I153091,I153198);
nor I_8846 (I153039,I153142,I153263);
DFFARX1 I_8847 (I74525,I2859,I153065,I153303,);
DFFARX1 I_8848 (I153303,I2859,I153065,I153320,);
not I_8849 (I153328,I153320);
not I_8850 (I153345,I153303);
nand I_8851 (I153042,I153345,I153164);
nand I_8852 (I153376,I74510,I74510);
and I_8853 (I153393,I153376,I74522);
DFFARX1 I_8854 (I153393,I2859,I153065,I153419,);
nor I_8855 (I153427,I153419,I153091);
DFFARX1 I_8856 (I153427,I2859,I153065,I153030,);
DFFARX1 I_8857 (I153419,I2859,I153065,I153048,);
nor I_8858 (I153472,I74528,I74510);
not I_8859 (I153489,I153472);
nor I_8860 (I153051,I153328,I153489);
nand I_8861 (I153036,I153345,I153489);
nor I_8862 (I153045,I153091,I153472);
DFFARX1 I_8863 (I153472,I2859,I153065,I153054,);
not I_8864 (I153592,I2866);
DFFARX1 I_8865 (I465490,I2859,I153592,I153618,);
nand I_8866 (I153626,I465505,I465490);
and I_8867 (I153643,I153626,I465508);
DFFARX1 I_8868 (I153643,I2859,I153592,I153669,);
nor I_8869 (I153560,I153669,I153618);
not I_8870 (I153691,I153669);
DFFARX1 I_8871 (I465514,I2859,I153592,I153717,);
nand I_8872 (I153725,I153717,I465496);
not I_8873 (I153742,I153725);
DFFARX1 I_8874 (I153742,I2859,I153592,I153768,);
not I_8875 (I153584,I153768);
nor I_8876 (I153790,I153618,I153725);
nor I_8877 (I153566,I153669,I153790);
DFFARX1 I_8878 (I465493,I2859,I153592,I153830,);
DFFARX1 I_8879 (I153830,I2859,I153592,I153847,);
not I_8880 (I153855,I153847);
not I_8881 (I153872,I153830);
nand I_8882 (I153569,I153872,I153691);
nand I_8883 (I153903,I465493,I465499);
and I_8884 (I153920,I153903,I465511);
DFFARX1 I_8885 (I153920,I2859,I153592,I153946,);
nor I_8886 (I153954,I153946,I153618);
DFFARX1 I_8887 (I153954,I2859,I153592,I153557,);
DFFARX1 I_8888 (I153946,I2859,I153592,I153575,);
nor I_8889 (I153999,I465502,I465499);
not I_8890 (I154016,I153999);
nor I_8891 (I153578,I153855,I154016);
nand I_8892 (I153563,I153872,I154016);
nor I_8893 (I153572,I153618,I153999);
DFFARX1 I_8894 (I153999,I2859,I153592,I153581,);
not I_8895 (I154119,I2866);
DFFARX1 I_8896 (I449306,I2859,I154119,I154145,);
nand I_8897 (I154153,I449321,I449306);
and I_8898 (I154170,I154153,I449324);
DFFARX1 I_8899 (I154170,I2859,I154119,I154196,);
nor I_8900 (I154087,I154196,I154145);
not I_8901 (I154218,I154196);
DFFARX1 I_8902 (I449330,I2859,I154119,I154244,);
nand I_8903 (I154252,I154244,I449312);
not I_8904 (I154269,I154252);
DFFARX1 I_8905 (I154269,I2859,I154119,I154295,);
not I_8906 (I154111,I154295);
nor I_8907 (I154317,I154145,I154252);
nor I_8908 (I154093,I154196,I154317);
DFFARX1 I_8909 (I449309,I2859,I154119,I154357,);
DFFARX1 I_8910 (I154357,I2859,I154119,I154374,);
not I_8911 (I154382,I154374);
not I_8912 (I154399,I154357);
nand I_8913 (I154096,I154399,I154218);
nand I_8914 (I154430,I449309,I449315);
and I_8915 (I154447,I154430,I449327);
DFFARX1 I_8916 (I154447,I2859,I154119,I154473,);
nor I_8917 (I154481,I154473,I154145);
DFFARX1 I_8918 (I154481,I2859,I154119,I154084,);
DFFARX1 I_8919 (I154473,I2859,I154119,I154102,);
nor I_8920 (I154526,I449318,I449315);
not I_8921 (I154543,I154526);
nor I_8922 (I154105,I154382,I154543);
nand I_8923 (I154090,I154399,I154543);
nor I_8924 (I154099,I154145,I154526);
DFFARX1 I_8925 (I154526,I2859,I154119,I154108,);
not I_8926 (I154646,I2866);
DFFARX1 I_8927 (I338095,I2859,I154646,I154672,);
nand I_8928 (I154680,I338098,I338092);
and I_8929 (I154697,I154680,I338104);
DFFARX1 I_8930 (I154697,I2859,I154646,I154723,);
nor I_8931 (I154614,I154723,I154672);
not I_8932 (I154745,I154723);
DFFARX1 I_8933 (I338107,I2859,I154646,I154771,);
nand I_8934 (I154779,I154771,I338098);
not I_8935 (I154796,I154779);
DFFARX1 I_8936 (I154796,I2859,I154646,I154822,);
not I_8937 (I154638,I154822);
nor I_8938 (I154844,I154672,I154779);
nor I_8939 (I154620,I154723,I154844);
DFFARX1 I_8940 (I338110,I2859,I154646,I154884,);
DFFARX1 I_8941 (I154884,I2859,I154646,I154901,);
not I_8942 (I154909,I154901);
not I_8943 (I154926,I154884);
nand I_8944 (I154623,I154926,I154745);
nand I_8945 (I154957,I338092,I338101);
and I_8946 (I154974,I154957,I338095);
DFFARX1 I_8947 (I154974,I2859,I154646,I155000,);
nor I_8948 (I155008,I155000,I154672);
DFFARX1 I_8949 (I155008,I2859,I154646,I154611,);
DFFARX1 I_8950 (I155000,I2859,I154646,I154629,);
nor I_8951 (I155053,I338113,I338101);
not I_8952 (I155070,I155053);
nor I_8953 (I154632,I154909,I155070);
nand I_8954 (I154617,I154926,I155070);
nor I_8955 (I154626,I154672,I155053);
DFFARX1 I_8956 (I155053,I2859,I154646,I154635,);
not I_8957 (I155173,I2866);
DFFARX1 I_8958 (I12695,I2859,I155173,I155199,);
nand I_8959 (I155207,I12719,I12698);
and I_8960 (I155224,I155207,I12695);
DFFARX1 I_8961 (I155224,I2859,I155173,I155250,);
nor I_8962 (I155141,I155250,I155199);
not I_8963 (I155272,I155250);
DFFARX1 I_8964 (I12701,I2859,I155173,I155298,);
nand I_8965 (I155306,I155298,I12710);
not I_8966 (I155323,I155306);
DFFARX1 I_8967 (I155323,I2859,I155173,I155349,);
not I_8968 (I155165,I155349);
nor I_8969 (I155371,I155199,I155306);
nor I_8970 (I155147,I155250,I155371);
DFFARX1 I_8971 (I12704,I2859,I155173,I155411,);
DFFARX1 I_8972 (I155411,I2859,I155173,I155428,);
not I_8973 (I155436,I155428);
not I_8974 (I155453,I155411);
nand I_8975 (I155150,I155453,I155272);
nand I_8976 (I155484,I12716,I12698);
and I_8977 (I155501,I155484,I12707);
DFFARX1 I_8978 (I155501,I2859,I155173,I155527,);
nor I_8979 (I155535,I155527,I155199);
DFFARX1 I_8980 (I155535,I2859,I155173,I155138,);
DFFARX1 I_8981 (I155527,I2859,I155173,I155156,);
nor I_8982 (I155580,I12713,I12698);
not I_8983 (I155597,I155580);
nor I_8984 (I155159,I155436,I155597);
nand I_8985 (I155144,I155453,I155597);
nor I_8986 (I155153,I155199,I155580);
DFFARX1 I_8987 (I155580,I2859,I155173,I155162,);
not I_8988 (I155700,I2866);
DFFARX1 I_8989 (I467224,I2859,I155700,I155726,);
nand I_8990 (I155734,I467239,I467224);
and I_8991 (I155751,I155734,I467242);
DFFARX1 I_8992 (I155751,I2859,I155700,I155777,);
nor I_8993 (I155668,I155777,I155726);
not I_8994 (I155799,I155777);
DFFARX1 I_8995 (I467248,I2859,I155700,I155825,);
nand I_8996 (I155833,I155825,I467230);
not I_8997 (I155850,I155833);
DFFARX1 I_8998 (I155850,I2859,I155700,I155876,);
not I_8999 (I155692,I155876);
nor I_9000 (I155898,I155726,I155833);
nor I_9001 (I155674,I155777,I155898);
DFFARX1 I_9002 (I467227,I2859,I155700,I155938,);
DFFARX1 I_9003 (I155938,I2859,I155700,I155955,);
not I_9004 (I155963,I155955);
not I_9005 (I155980,I155938);
nand I_9006 (I155677,I155980,I155799);
nand I_9007 (I156011,I467227,I467233);
and I_9008 (I156028,I156011,I467245);
DFFARX1 I_9009 (I156028,I2859,I155700,I156054,);
nor I_9010 (I156062,I156054,I155726);
DFFARX1 I_9011 (I156062,I2859,I155700,I155665,);
DFFARX1 I_9012 (I156054,I2859,I155700,I155683,);
nor I_9013 (I156107,I467236,I467233);
not I_9014 (I156124,I156107);
nor I_9015 (I155686,I155963,I156124);
nand I_9016 (I155671,I155980,I156124);
nor I_9017 (I155680,I155726,I156107);
DFFARX1 I_9018 (I156107,I2859,I155700,I155689,);
not I_9019 (I156227,I2866);
DFFARX1 I_9020 (I441792,I2859,I156227,I156253,);
nand I_9021 (I156261,I441807,I441792);
and I_9022 (I156278,I156261,I441810);
DFFARX1 I_9023 (I156278,I2859,I156227,I156304,);
nor I_9024 (I156195,I156304,I156253);
not I_9025 (I156326,I156304);
DFFARX1 I_9026 (I441816,I2859,I156227,I156352,);
nand I_9027 (I156360,I156352,I441798);
not I_9028 (I156377,I156360);
DFFARX1 I_9029 (I156377,I2859,I156227,I156403,);
not I_9030 (I156219,I156403);
nor I_9031 (I156425,I156253,I156360);
nor I_9032 (I156201,I156304,I156425);
DFFARX1 I_9033 (I441795,I2859,I156227,I156465,);
DFFARX1 I_9034 (I156465,I2859,I156227,I156482,);
not I_9035 (I156490,I156482);
not I_9036 (I156507,I156465);
nand I_9037 (I156204,I156507,I156326);
nand I_9038 (I156538,I441795,I441801);
and I_9039 (I156555,I156538,I441813);
DFFARX1 I_9040 (I156555,I2859,I156227,I156581,);
nor I_9041 (I156589,I156581,I156253);
DFFARX1 I_9042 (I156589,I2859,I156227,I156192,);
DFFARX1 I_9043 (I156581,I2859,I156227,I156210,);
nor I_9044 (I156634,I441804,I441801);
not I_9045 (I156651,I156634);
nor I_9046 (I156213,I156490,I156651);
nand I_9047 (I156198,I156507,I156651);
nor I_9048 (I156207,I156253,I156634);
DFFARX1 I_9049 (I156634,I2859,I156227,I156216,);
not I_9050 (I156754,I2866);
DFFARX1 I_9051 (I38521,I2859,I156754,I156780,);
nand I_9052 (I156788,I38533,I38542);
and I_9053 (I156805,I156788,I38521);
DFFARX1 I_9054 (I156805,I2859,I156754,I156831,);
nor I_9055 (I156722,I156831,I156780);
not I_9056 (I156853,I156831);
DFFARX1 I_9057 (I38536,I2859,I156754,I156879,);
nand I_9058 (I156887,I156879,I38524);
not I_9059 (I156904,I156887);
DFFARX1 I_9060 (I156904,I2859,I156754,I156930,);
not I_9061 (I156746,I156930);
nor I_9062 (I156952,I156780,I156887);
nor I_9063 (I156728,I156831,I156952);
DFFARX1 I_9064 (I38527,I2859,I156754,I156992,);
DFFARX1 I_9065 (I156992,I2859,I156754,I157009,);
not I_9066 (I157017,I157009);
not I_9067 (I157034,I156992);
nand I_9068 (I156731,I157034,I156853);
nand I_9069 (I157065,I38518,I38518);
and I_9070 (I157082,I157065,I38530);
DFFARX1 I_9071 (I157082,I2859,I156754,I157108,);
nor I_9072 (I157116,I157108,I156780);
DFFARX1 I_9073 (I157116,I2859,I156754,I156719,);
DFFARX1 I_9074 (I157108,I2859,I156754,I156737,);
nor I_9075 (I157161,I38539,I38518);
not I_9076 (I157178,I157161);
nor I_9077 (I156740,I157017,I157178);
nand I_9078 (I156725,I157034,I157178);
nor I_9079 (I156734,I156780,I157161);
DFFARX1 I_9080 (I157161,I2859,I156754,I156743,);
not I_9081 (I157281,I2866);
DFFARX1 I_9082 (I310564,I2859,I157281,I157307,);
nand I_9083 (I157315,I310555,I310570);
and I_9084 (I157332,I157315,I310576);
DFFARX1 I_9085 (I157332,I2859,I157281,I157358,);
nor I_9086 (I157249,I157358,I157307);
not I_9087 (I157380,I157358);
DFFARX1 I_9088 (I310561,I2859,I157281,I157406,);
nand I_9089 (I157414,I157406,I310555);
not I_9090 (I157431,I157414);
DFFARX1 I_9091 (I157431,I2859,I157281,I157457,);
not I_9092 (I157273,I157457);
nor I_9093 (I157479,I157307,I157414);
nor I_9094 (I157255,I157358,I157479);
DFFARX1 I_9095 (I310558,I2859,I157281,I157519,);
DFFARX1 I_9096 (I157519,I2859,I157281,I157536,);
not I_9097 (I157544,I157536);
not I_9098 (I157561,I157519);
nand I_9099 (I157258,I157561,I157380);
nand I_9100 (I157592,I310552,I310567);
and I_9101 (I157609,I157592,I310552);
DFFARX1 I_9102 (I157609,I2859,I157281,I157635,);
nor I_9103 (I157643,I157635,I157307);
DFFARX1 I_9104 (I157643,I2859,I157281,I157246,);
DFFARX1 I_9105 (I157635,I2859,I157281,I157264,);
nor I_9106 (I157688,I310573,I310567);
not I_9107 (I157705,I157688);
nor I_9108 (I157267,I157544,I157705);
nand I_9109 (I157252,I157561,I157705);
nor I_9110 (I157261,I157307,I157688);
DFFARX1 I_9111 (I157688,I2859,I157281,I157270,);
not I_9112 (I157808,I2866);
DFFARX1 I_9113 (I458554,I2859,I157808,I157834,);
nand I_9114 (I157842,I458569,I458554);
and I_9115 (I157859,I157842,I458572);
DFFARX1 I_9116 (I157859,I2859,I157808,I157885,);
nor I_9117 (I157776,I157885,I157834);
not I_9118 (I157907,I157885);
DFFARX1 I_9119 (I458578,I2859,I157808,I157933,);
nand I_9120 (I157941,I157933,I458560);
not I_9121 (I157958,I157941);
DFFARX1 I_9122 (I157958,I2859,I157808,I157984,);
not I_9123 (I157800,I157984);
nor I_9124 (I158006,I157834,I157941);
nor I_9125 (I157782,I157885,I158006);
DFFARX1 I_9126 (I458557,I2859,I157808,I158046,);
DFFARX1 I_9127 (I158046,I2859,I157808,I158063,);
not I_9128 (I158071,I158063);
not I_9129 (I158088,I158046);
nand I_9130 (I157785,I158088,I157907);
nand I_9131 (I158119,I458557,I458563);
and I_9132 (I158136,I158119,I458575);
DFFARX1 I_9133 (I158136,I2859,I157808,I158162,);
nor I_9134 (I158170,I158162,I157834);
DFFARX1 I_9135 (I158170,I2859,I157808,I157773,);
DFFARX1 I_9136 (I158162,I2859,I157808,I157791,);
nor I_9137 (I158215,I458566,I458563);
not I_9138 (I158232,I158215);
nor I_9139 (I157794,I158071,I158232);
nand I_9140 (I157779,I158088,I158232);
nor I_9141 (I157788,I157834,I158215);
DFFARX1 I_9142 (I158215,I2859,I157808,I157797,);
not I_9143 (I158335,I2866);
DFFARX1 I_9144 (I257388,I2859,I158335,I158361,);
nand I_9145 (I158369,I257379,I257394);
and I_9146 (I158386,I158369,I257400);
DFFARX1 I_9147 (I158386,I2859,I158335,I158412,);
nor I_9148 (I158303,I158412,I158361);
not I_9149 (I158434,I158412);
DFFARX1 I_9150 (I257385,I2859,I158335,I158460,);
nand I_9151 (I158468,I158460,I257379);
not I_9152 (I158485,I158468);
DFFARX1 I_9153 (I158485,I2859,I158335,I158511,);
not I_9154 (I158327,I158511);
nor I_9155 (I158533,I158361,I158468);
nor I_9156 (I158309,I158412,I158533);
DFFARX1 I_9157 (I257382,I2859,I158335,I158573,);
DFFARX1 I_9158 (I158573,I2859,I158335,I158590,);
not I_9159 (I158598,I158590);
not I_9160 (I158615,I158573);
nand I_9161 (I158312,I158615,I158434);
nand I_9162 (I158646,I257376,I257391);
and I_9163 (I158663,I158646,I257376);
DFFARX1 I_9164 (I158663,I2859,I158335,I158689,);
nor I_9165 (I158697,I158689,I158361);
DFFARX1 I_9166 (I158697,I2859,I158335,I158300,);
DFFARX1 I_9167 (I158689,I2859,I158335,I158318,);
nor I_9168 (I158742,I257397,I257391);
not I_9169 (I158759,I158742);
nor I_9170 (I158321,I158598,I158759);
nand I_9171 (I158306,I158615,I158759);
nor I_9172 (I158315,I158361,I158742);
DFFARX1 I_9173 (I158742,I2859,I158335,I158324,);
not I_9174 (I158862,I2866);
DFFARX1 I_9175 (I434978,I2859,I158862,I158888,);
nand I_9176 (I158896,I434975,I434978);
and I_9177 (I158913,I158896,I434987);
DFFARX1 I_9178 (I158913,I2859,I158862,I158939,);
nor I_9179 (I158830,I158939,I158888);
not I_9180 (I158961,I158939);
DFFARX1 I_9181 (I434975,I2859,I158862,I158987,);
nand I_9182 (I158995,I158987,I434993);
not I_9183 (I159012,I158995);
DFFARX1 I_9184 (I159012,I2859,I158862,I159038,);
not I_9185 (I158854,I159038);
nor I_9186 (I159060,I158888,I158995);
nor I_9187 (I158836,I158939,I159060);
DFFARX1 I_9188 (I434981,I2859,I158862,I159100,);
DFFARX1 I_9189 (I159100,I2859,I158862,I159117,);
not I_9190 (I159125,I159117);
not I_9191 (I159142,I159100);
nand I_9192 (I158839,I159142,I158961);
nand I_9193 (I159173,I434990,I434996);
and I_9194 (I159190,I159173,I434981);
DFFARX1 I_9195 (I159190,I2859,I158862,I159216,);
nor I_9196 (I159224,I159216,I158888);
DFFARX1 I_9197 (I159224,I2859,I158862,I158827,);
DFFARX1 I_9198 (I159216,I2859,I158862,I158845,);
nor I_9199 (I159269,I434984,I434996);
not I_9200 (I159286,I159269);
nor I_9201 (I158848,I159125,I159286);
nand I_9202 (I158833,I159142,I159286);
nor I_9203 (I158842,I158888,I159269);
DFFARX1 I_9204 (I159269,I2859,I158862,I158851,);
not I_9205 (I159389,I2866);
DFFARX1 I_9206 (I253345,I2859,I159389,I159415,);
nand I_9207 (I159423,I253330,I253333);
and I_9208 (I159440,I159423,I253348);
DFFARX1 I_9209 (I159440,I2859,I159389,I159466,);
nor I_9210 (I159357,I159466,I159415);
not I_9211 (I159488,I159466);
DFFARX1 I_9212 (I253342,I2859,I159389,I159514,);
nand I_9213 (I159522,I159514,I253333);
not I_9214 (I159539,I159522);
DFFARX1 I_9215 (I159539,I2859,I159389,I159565,);
not I_9216 (I159381,I159565);
nor I_9217 (I159587,I159415,I159522);
nor I_9218 (I159363,I159466,I159587);
DFFARX1 I_9219 (I253339,I2859,I159389,I159627,);
DFFARX1 I_9220 (I159627,I2859,I159389,I159644,);
not I_9221 (I159652,I159644);
not I_9222 (I159669,I159627);
nand I_9223 (I159366,I159669,I159488);
nand I_9224 (I159700,I253354,I253330);
and I_9225 (I159717,I159700,I253351);
DFFARX1 I_9226 (I159717,I2859,I159389,I159743,);
nor I_9227 (I159751,I159743,I159415);
DFFARX1 I_9228 (I159751,I2859,I159389,I159354,);
DFFARX1 I_9229 (I159743,I2859,I159389,I159372,);
nor I_9230 (I159796,I253336,I253330);
not I_9231 (I159813,I159796);
nor I_9232 (I159375,I159652,I159813);
nand I_9233 (I159360,I159669,I159813);
nor I_9234 (I159369,I159415,I159796);
DFFARX1 I_9235 (I159796,I2859,I159389,I159378,);
not I_9236 (I159916,I2866);
DFFARX1 I_9237 (I160964,I2859,I159916,I159942,);
nand I_9238 (I159950,I160976,I160955);
and I_9239 (I159967,I159950,I160979);
DFFARX1 I_9240 (I159967,I2859,I159916,I159993,);
nor I_9241 (I159884,I159993,I159942);
not I_9242 (I160015,I159993);
DFFARX1 I_9243 (I160970,I2859,I159916,I160041,);
nand I_9244 (I160049,I160041,I160952);
not I_9245 (I160066,I160049);
DFFARX1 I_9246 (I160066,I2859,I159916,I160092,);
not I_9247 (I159908,I160092);
nor I_9248 (I160114,I159942,I160049);
nor I_9249 (I159890,I159993,I160114);
DFFARX1 I_9250 (I160967,I2859,I159916,I160154,);
DFFARX1 I_9251 (I160154,I2859,I159916,I160171,);
not I_9252 (I160179,I160171);
not I_9253 (I160196,I160154);
nand I_9254 (I159893,I160196,I160015);
nand I_9255 (I160227,I160952,I160958);
and I_9256 (I160244,I160227,I160961);
DFFARX1 I_9257 (I160244,I2859,I159916,I160270,);
nor I_9258 (I160278,I160270,I159942);
DFFARX1 I_9259 (I160278,I2859,I159916,I159881,);
DFFARX1 I_9260 (I160270,I2859,I159916,I159899,);
nor I_9261 (I160323,I160973,I160958);
not I_9262 (I160340,I160323);
nor I_9263 (I159902,I160179,I160340);
nand I_9264 (I159887,I160196,I160340);
nor I_9265 (I159896,I159942,I160323);
DFFARX1 I_9266 (I160323,I2859,I159916,I159905,);
not I_9267 (I160443,I2866);
DFFARX1 I_9268 (I501907,I2859,I160443,I160469,);
DFFARX1 I_9269 (I160469,I2859,I160443,I160486,);
not I_9270 (I160435,I160486);
not I_9271 (I160508,I160469);
nand I_9272 (I160525,I501919,I501907);
and I_9273 (I160542,I160525,I501910);
DFFARX1 I_9274 (I160542,I2859,I160443,I160568,);
not I_9275 (I160576,I160568);
DFFARX1 I_9276 (I501928,I2859,I160443,I160602,);
and I_9277 (I160610,I160602,I501904);
nand I_9278 (I160627,I160602,I501904);
nand I_9279 (I160414,I160576,I160627);
DFFARX1 I_9280 (I501922,I2859,I160443,I160667,);
nor I_9281 (I160675,I160667,I160610);
DFFARX1 I_9282 (I160675,I2859,I160443,I160408,);
nor I_9283 (I160423,I160667,I160568);
nand I_9284 (I160720,I501916,I501913);
and I_9285 (I160737,I160720,I501925);
DFFARX1 I_9286 (I160737,I2859,I160443,I160763,);
nor I_9287 (I160411,I160763,I160667);
not I_9288 (I160785,I160763);
nor I_9289 (I160802,I160785,I160576);
nor I_9290 (I160819,I160508,I160802);
DFFARX1 I_9291 (I160819,I2859,I160443,I160426,);
nor I_9292 (I160850,I160785,I160667);
nor I_9293 (I160867,I501904,I501913);
nor I_9294 (I160417,I160867,I160850);
not I_9295 (I160898,I160867);
nand I_9296 (I160420,I160627,I160898);
DFFARX1 I_9297 (I160867,I2859,I160443,I160432,);
DFFARX1 I_9298 (I160867,I2859,I160443,I160429,);
not I_9299 (I160987,I2866);
DFFARX1 I_9300 (I501329,I2859,I160987,I161013,);
DFFARX1 I_9301 (I161013,I2859,I160987,I161030,);
not I_9302 (I160979,I161030);
not I_9303 (I161052,I161013);
nand I_9304 (I161069,I501341,I501329);
and I_9305 (I161086,I161069,I501332);
DFFARX1 I_9306 (I161086,I2859,I160987,I161112,);
not I_9307 (I161120,I161112);
DFFARX1 I_9308 (I501350,I2859,I160987,I161146,);
and I_9309 (I161154,I161146,I501326);
nand I_9310 (I161171,I161146,I501326);
nand I_9311 (I160958,I161120,I161171);
DFFARX1 I_9312 (I501344,I2859,I160987,I161211,);
nor I_9313 (I161219,I161211,I161154);
DFFARX1 I_9314 (I161219,I2859,I160987,I160952,);
nor I_9315 (I160967,I161211,I161112);
nand I_9316 (I161264,I501338,I501335);
and I_9317 (I161281,I161264,I501347);
DFFARX1 I_9318 (I161281,I2859,I160987,I161307,);
nor I_9319 (I160955,I161307,I161211);
not I_9320 (I161329,I161307);
nor I_9321 (I161346,I161329,I161120);
nor I_9322 (I161363,I161052,I161346);
DFFARX1 I_9323 (I161363,I2859,I160987,I160970,);
nor I_9324 (I161394,I161329,I161211);
nor I_9325 (I161411,I501326,I501335);
nor I_9326 (I160961,I161411,I161394);
not I_9327 (I161442,I161411);
nand I_9328 (I160964,I161171,I161442);
DFFARX1 I_9329 (I161411,I2859,I160987,I160976,);
DFFARX1 I_9330 (I161411,I2859,I160987,I160973,);
not I_9331 (I161531,I2866);
DFFARX1 I_9332 (I294371,I2859,I161531,I161557,);
DFFARX1 I_9333 (I161557,I2859,I161531,I161574,);
not I_9334 (I161523,I161574);
not I_9335 (I161596,I161557);
nand I_9336 (I161613,I294392,I294383);
and I_9337 (I161630,I161613,I294371);
DFFARX1 I_9338 (I161630,I2859,I161531,I161656,);
not I_9339 (I161664,I161656);
DFFARX1 I_9340 (I294377,I2859,I161531,I161690,);
and I_9341 (I161698,I161690,I294374);
nand I_9342 (I161715,I161690,I294374);
nand I_9343 (I161502,I161664,I161715);
DFFARX1 I_9344 (I294368,I2859,I161531,I161755,);
nor I_9345 (I161763,I161755,I161698);
DFFARX1 I_9346 (I161763,I2859,I161531,I161496,);
nor I_9347 (I161511,I161755,I161656);
nand I_9348 (I161808,I294368,I294380);
and I_9349 (I161825,I161808,I294389);
DFFARX1 I_9350 (I161825,I2859,I161531,I161851,);
nor I_9351 (I161499,I161851,I161755);
not I_9352 (I161873,I161851);
nor I_9353 (I161890,I161873,I161664);
nor I_9354 (I161907,I161596,I161890);
DFFARX1 I_9355 (I161907,I2859,I161531,I161514,);
nor I_9356 (I161938,I161873,I161755);
nor I_9357 (I161955,I294386,I294380);
nor I_9358 (I161505,I161955,I161938);
not I_9359 (I161986,I161955);
nand I_9360 (I161508,I161715,I161986);
DFFARX1 I_9361 (I161955,I2859,I161531,I161520,);
DFFARX1 I_9362 (I161955,I2859,I161531,I161517,);
not I_9363 (I162075,I2866);
DFFARX1 I_9364 (I7437,I2859,I162075,I162101,);
DFFARX1 I_9365 (I162101,I2859,I162075,I162118,);
not I_9366 (I162067,I162118);
not I_9367 (I162140,I162101);
nand I_9368 (I162157,I7425,I7440);
and I_9369 (I162174,I162157,I7428);
DFFARX1 I_9370 (I162174,I2859,I162075,I162200,);
not I_9371 (I162208,I162200);
DFFARX1 I_9372 (I7449,I2859,I162075,I162234,);
and I_9373 (I162242,I162234,I7443);
nand I_9374 (I162259,I162234,I7443);
nand I_9375 (I162046,I162208,I162259);
DFFARX1 I_9376 (I7446,I2859,I162075,I162299,);
nor I_9377 (I162307,I162299,I162242);
DFFARX1 I_9378 (I162307,I2859,I162075,I162040,);
nor I_9379 (I162055,I162299,I162200);
nand I_9380 (I162352,I7425,I7428);
and I_9381 (I162369,I162352,I7431);
DFFARX1 I_9382 (I162369,I2859,I162075,I162395,);
nor I_9383 (I162043,I162395,I162299);
not I_9384 (I162417,I162395);
nor I_9385 (I162434,I162417,I162208);
nor I_9386 (I162451,I162140,I162434);
DFFARX1 I_9387 (I162451,I2859,I162075,I162058,);
nor I_9388 (I162482,I162417,I162299);
nor I_9389 (I162499,I7434,I7428);
nor I_9390 (I162049,I162499,I162482);
not I_9391 (I162530,I162499);
nand I_9392 (I162052,I162259,I162530);
DFFARX1 I_9393 (I162499,I2859,I162075,I162064,);
DFFARX1 I_9394 (I162499,I2859,I162075,I162061,);
not I_9395 (I162619,I2866);
DFFARX1 I_9396 (I19025,I2859,I162619,I162645,);
DFFARX1 I_9397 (I162645,I2859,I162619,I162662,);
not I_9398 (I162611,I162662);
not I_9399 (I162684,I162645);
nand I_9400 (I162701,I19040,I19019);
and I_9401 (I162718,I162701,I19022);
DFFARX1 I_9402 (I162718,I2859,I162619,I162744,);
not I_9403 (I162752,I162744);
DFFARX1 I_9404 (I19028,I2859,I162619,I162778,);
and I_9405 (I162786,I162778,I19022);
nand I_9406 (I162803,I162778,I19022);
nand I_9407 (I162590,I162752,I162803);
DFFARX1 I_9408 (I19037,I2859,I162619,I162843,);
nor I_9409 (I162851,I162843,I162786);
DFFARX1 I_9410 (I162851,I2859,I162619,I162584,);
nor I_9411 (I162599,I162843,I162744);
nand I_9412 (I162896,I19019,I19034);
and I_9413 (I162913,I162896,I19031);
DFFARX1 I_9414 (I162913,I2859,I162619,I162939,);
nor I_9415 (I162587,I162939,I162843);
not I_9416 (I162961,I162939);
nor I_9417 (I162978,I162961,I162752);
nor I_9418 (I162995,I162684,I162978);
DFFARX1 I_9419 (I162995,I2859,I162619,I162602,);
nor I_9420 (I163026,I162961,I162843);
nor I_9421 (I163043,I19043,I19034);
nor I_9422 (I162593,I163043,I163026);
not I_9423 (I163074,I163043);
nand I_9424 (I162596,I162803,I163074);
DFFARX1 I_9425 (I163043,I2859,I162619,I162608,);
DFFARX1 I_9426 (I163043,I2859,I162619,I162605,);
not I_9427 (I163163,I2866);
DFFARX1 I_9428 (I232525,I2859,I163163,I163189,);
DFFARX1 I_9429 (I163189,I2859,I163163,I163206,);
not I_9430 (I163155,I163206);
not I_9431 (I163228,I163189);
nand I_9432 (I163245,I232522,I232543);
and I_9433 (I163262,I163245,I232546);
DFFARX1 I_9434 (I163262,I2859,I163163,I163288,);
not I_9435 (I163296,I163288);
DFFARX1 I_9436 (I232531,I2859,I163163,I163322,);
and I_9437 (I163330,I163322,I232534);
nand I_9438 (I163347,I163322,I232534);
nand I_9439 (I163134,I163296,I163347);
DFFARX1 I_9440 (I232537,I2859,I163163,I163387,);
nor I_9441 (I163395,I163387,I163330);
DFFARX1 I_9442 (I163395,I2859,I163163,I163128,);
nor I_9443 (I163143,I163387,I163288);
nand I_9444 (I163440,I232522,I232528);
and I_9445 (I163457,I163440,I232540);
DFFARX1 I_9446 (I163457,I2859,I163163,I163483,);
nor I_9447 (I163131,I163483,I163387);
not I_9448 (I163505,I163483);
nor I_9449 (I163522,I163505,I163296);
nor I_9450 (I163539,I163228,I163522);
DFFARX1 I_9451 (I163539,I2859,I163163,I163146,);
nor I_9452 (I163570,I163505,I163387);
nor I_9453 (I163587,I232525,I232528);
nor I_9454 (I163137,I163587,I163570);
not I_9455 (I163618,I163587);
nand I_9456 (I163140,I163347,I163618);
DFFARX1 I_9457 (I163587,I2859,I163163,I163152,);
DFFARX1 I_9458 (I163587,I2859,I163163,I163149,);
not I_9459 (I163707,I2866);
DFFARX1 I_9460 (I49064,I2859,I163707,I163733,);
DFFARX1 I_9461 (I163733,I2859,I163707,I163750,);
not I_9462 (I163699,I163750);
not I_9463 (I163772,I163733);
nand I_9464 (I163789,I49079,I49058);
and I_9465 (I163806,I163789,I49061);
DFFARX1 I_9466 (I163806,I2859,I163707,I163832,);
not I_9467 (I163840,I163832);
DFFARX1 I_9468 (I49067,I2859,I163707,I163866,);
and I_9469 (I163874,I163866,I49061);
nand I_9470 (I163891,I163866,I49061);
nand I_9471 (I163678,I163840,I163891);
DFFARX1 I_9472 (I49076,I2859,I163707,I163931,);
nor I_9473 (I163939,I163931,I163874);
DFFARX1 I_9474 (I163939,I2859,I163707,I163672,);
nor I_9475 (I163687,I163931,I163832);
nand I_9476 (I163984,I49058,I49073);
and I_9477 (I164001,I163984,I49070);
DFFARX1 I_9478 (I164001,I2859,I163707,I164027,);
nor I_9479 (I163675,I164027,I163931);
not I_9480 (I164049,I164027);
nor I_9481 (I164066,I164049,I163840);
nor I_9482 (I164083,I163772,I164066);
DFFARX1 I_9483 (I164083,I2859,I163707,I163690,);
nor I_9484 (I164114,I164049,I163931);
nor I_9485 (I164131,I49082,I49073);
nor I_9486 (I163681,I164131,I164114);
not I_9487 (I164162,I164131);
nand I_9488 (I163684,I163891,I164162);
DFFARX1 I_9489 (I164131,I2859,I163707,I163696,);
DFFARX1 I_9490 (I164131,I2859,I163707,I163693,);
not I_9491 (I164251,I2866);
DFFARX1 I_9492 (I368273,I2859,I164251,I164277,);
DFFARX1 I_9493 (I164277,I2859,I164251,I164294,);
not I_9494 (I164243,I164294);
not I_9495 (I164316,I164277);
nand I_9496 (I164333,I368288,I368276);
and I_9497 (I164350,I164333,I368267);
DFFARX1 I_9498 (I164350,I2859,I164251,I164376,);
not I_9499 (I164384,I164376);
DFFARX1 I_9500 (I368279,I2859,I164251,I164410,);
and I_9501 (I164418,I164410,I368270);
nand I_9502 (I164435,I164410,I368270);
nand I_9503 (I164222,I164384,I164435);
DFFARX1 I_9504 (I368285,I2859,I164251,I164475,);
nor I_9505 (I164483,I164475,I164418);
DFFARX1 I_9506 (I164483,I2859,I164251,I164216,);
nor I_9507 (I164231,I164475,I164376);
nand I_9508 (I164528,I368294,I368282);
and I_9509 (I164545,I164528,I368291);
DFFARX1 I_9510 (I164545,I2859,I164251,I164571,);
nor I_9511 (I164219,I164571,I164475);
not I_9512 (I164593,I164571);
nor I_9513 (I164610,I164593,I164384);
nor I_9514 (I164627,I164316,I164610);
DFFARX1 I_9515 (I164627,I2859,I164251,I164234,);
nor I_9516 (I164658,I164593,I164475);
nor I_9517 (I164675,I368267,I368282);
nor I_9518 (I164225,I164675,I164658);
not I_9519 (I164706,I164675);
nand I_9520 (I164228,I164435,I164706);
DFFARX1 I_9521 (I164675,I2859,I164251,I164240,);
DFFARX1 I_9522 (I164675,I2859,I164251,I164237,);
not I_9523 (I164795,I2866);
DFFARX1 I_9524 (I157794,I2859,I164795,I164821,);
DFFARX1 I_9525 (I164821,I2859,I164795,I164838,);
not I_9526 (I164787,I164838);
not I_9527 (I164860,I164821);
nand I_9528 (I164877,I157773,I157797);
and I_9529 (I164894,I164877,I157800);
DFFARX1 I_9530 (I164894,I2859,I164795,I164920,);
not I_9531 (I164928,I164920);
DFFARX1 I_9532 (I157782,I2859,I164795,I164954,);
and I_9533 (I164962,I164954,I157788);
nand I_9534 (I164979,I164954,I157788);
nand I_9535 (I164766,I164928,I164979);
DFFARX1 I_9536 (I157776,I2859,I164795,I165019,);
nor I_9537 (I165027,I165019,I164962);
DFFARX1 I_9538 (I165027,I2859,I164795,I164760,);
nor I_9539 (I164775,I165019,I164920);
nand I_9540 (I165072,I157785,I157773);
and I_9541 (I165089,I165072,I157779);
DFFARX1 I_9542 (I165089,I2859,I164795,I165115,);
nor I_9543 (I164763,I165115,I165019);
not I_9544 (I165137,I165115);
nor I_9545 (I165154,I165137,I164928);
nor I_9546 (I165171,I164860,I165154);
DFFARX1 I_9547 (I165171,I2859,I164795,I164778,);
nor I_9548 (I165202,I165137,I165019);
nor I_9549 (I165219,I157791,I157773);
nor I_9550 (I164769,I165219,I165202);
not I_9551 (I165250,I165219);
nand I_9552 (I164772,I164979,I165250);
DFFARX1 I_9553 (I165219,I2859,I164795,I164784,);
DFFARX1 I_9554 (I165219,I2859,I164795,I164781,);
not I_9555 (I165339,I2866);
DFFARX1 I_9556 (I352860,I2859,I165339,I165365,);
DFFARX1 I_9557 (I165365,I2859,I165339,I165382,);
not I_9558 (I165331,I165382);
not I_9559 (I165404,I165365);
nand I_9560 (I165421,I352854,I352851);
and I_9561 (I165438,I165421,I352866);
DFFARX1 I_9562 (I165438,I2859,I165339,I165464,);
not I_9563 (I165472,I165464);
DFFARX1 I_9564 (I352854,I2859,I165339,I165498,);
and I_9565 (I165506,I165498,I352848);
nand I_9566 (I165523,I165498,I352848);
nand I_9567 (I165310,I165472,I165523);
DFFARX1 I_9568 (I352848,I2859,I165339,I165563,);
nor I_9569 (I165571,I165563,I165506);
DFFARX1 I_9570 (I165571,I2859,I165339,I165304,);
nor I_9571 (I165319,I165563,I165464);
nand I_9572 (I165616,I352863,I352857);
and I_9573 (I165633,I165616,I352851);
DFFARX1 I_9574 (I165633,I2859,I165339,I165659,);
nor I_9575 (I165307,I165659,I165563);
not I_9576 (I165681,I165659);
nor I_9577 (I165698,I165681,I165472);
nor I_9578 (I165715,I165404,I165698);
DFFARX1 I_9579 (I165715,I2859,I165339,I165322,);
nor I_9580 (I165746,I165681,I165563);
nor I_9581 (I165763,I352869,I352857);
nor I_9582 (I165313,I165763,I165746);
not I_9583 (I165794,I165763);
nand I_9584 (I165316,I165523,I165794);
DFFARX1 I_9585 (I165763,I2859,I165339,I165328,);
DFFARX1 I_9586 (I165763,I2859,I165339,I165325,);
not I_9587 (I165883,I2866);
DFFARX1 I_9588 (I425438,I2859,I165883,I165909,);
DFFARX1 I_9589 (I165909,I2859,I165883,I165926,);
not I_9590 (I165875,I165926);
not I_9591 (I165948,I165909);
nand I_9592 (I165965,I425438,I425456);
and I_9593 (I165982,I165965,I425450);
DFFARX1 I_9594 (I165982,I2859,I165883,I166008,);
not I_9595 (I166016,I166008);
DFFARX1 I_9596 (I425444,I2859,I165883,I166042,);
and I_9597 (I166050,I166042,I425453);
nand I_9598 (I166067,I166042,I425453);
nand I_9599 (I165854,I166016,I166067);
DFFARX1 I_9600 (I425441,I2859,I165883,I166107,);
nor I_9601 (I166115,I166107,I166050);
DFFARX1 I_9602 (I166115,I2859,I165883,I165848,);
nor I_9603 (I165863,I166107,I166008);
nand I_9604 (I166160,I425441,I425459);
and I_9605 (I166177,I166160,I425444);
DFFARX1 I_9606 (I166177,I2859,I165883,I166203,);
nor I_9607 (I165851,I166203,I166107);
not I_9608 (I166225,I166203);
nor I_9609 (I166242,I166225,I166016);
nor I_9610 (I166259,I165948,I166242);
DFFARX1 I_9611 (I166259,I2859,I165883,I165866,);
nor I_9612 (I166290,I166225,I166107);
nor I_9613 (I166307,I425447,I425459);
nor I_9614 (I165857,I166307,I166290);
not I_9615 (I166338,I166307);
nand I_9616 (I165860,I166067,I166338);
DFFARX1 I_9617 (I166307,I2859,I165883,I165872,);
DFFARX1 I_9618 (I166307,I2859,I165883,I165869,);
not I_9619 (I166427,I2866);
DFFARX1 I_9620 (I368919,I2859,I166427,I166453,);
DFFARX1 I_9621 (I166453,I2859,I166427,I166470,);
not I_9622 (I166419,I166470);
not I_9623 (I166492,I166453);
nand I_9624 (I166509,I368934,I368922);
and I_9625 (I166526,I166509,I368913);
DFFARX1 I_9626 (I166526,I2859,I166427,I166552,);
not I_9627 (I166560,I166552);
DFFARX1 I_9628 (I368925,I2859,I166427,I166586,);
and I_9629 (I166594,I166586,I368916);
nand I_9630 (I166611,I166586,I368916);
nand I_9631 (I166398,I166560,I166611);
DFFARX1 I_9632 (I368931,I2859,I166427,I166651,);
nor I_9633 (I166659,I166651,I166594);
DFFARX1 I_9634 (I166659,I2859,I166427,I166392,);
nor I_9635 (I166407,I166651,I166552);
nand I_9636 (I166704,I368940,I368928);
and I_9637 (I166721,I166704,I368937);
DFFARX1 I_9638 (I166721,I2859,I166427,I166747,);
nor I_9639 (I166395,I166747,I166651);
not I_9640 (I166769,I166747);
nor I_9641 (I166786,I166769,I166560);
nor I_9642 (I166803,I166492,I166786);
DFFARX1 I_9643 (I166803,I2859,I166427,I166410,);
nor I_9644 (I166834,I166769,I166651);
nor I_9645 (I166851,I368913,I368928);
nor I_9646 (I166401,I166851,I166834);
not I_9647 (I166882,I166851);
nand I_9648 (I166404,I166611,I166882);
DFFARX1 I_9649 (I166851,I2859,I166427,I166416,);
DFFARX1 I_9650 (I166851,I2859,I166427,I166413,);
not I_9651 (I166971,I2866);
DFFARX1 I_9652 (I109621,I2859,I166971,I166997,);
DFFARX1 I_9653 (I166997,I2859,I166971,I167014,);
not I_9654 (I166963,I167014);
not I_9655 (I167036,I166997);
nand I_9656 (I167053,I109633,I109612);
and I_9657 (I167070,I167053,I109615);
DFFARX1 I_9658 (I167070,I2859,I166971,I167096,);
not I_9659 (I167104,I167096);
DFFARX1 I_9660 (I109624,I2859,I166971,I167130,);
and I_9661 (I167138,I167130,I109636);
nand I_9662 (I167155,I167130,I109636);
nand I_9663 (I166942,I167104,I167155);
DFFARX1 I_9664 (I109630,I2859,I166971,I167195,);
nor I_9665 (I167203,I167195,I167138);
DFFARX1 I_9666 (I167203,I2859,I166971,I166936,);
nor I_9667 (I166951,I167195,I167096);
nand I_9668 (I167248,I109618,I109615);
and I_9669 (I167265,I167248,I109627);
DFFARX1 I_9670 (I167265,I2859,I166971,I167291,);
nor I_9671 (I166939,I167291,I167195);
not I_9672 (I167313,I167291);
nor I_9673 (I167330,I167313,I167104);
nor I_9674 (I167347,I167036,I167330);
DFFARX1 I_9675 (I167347,I2859,I166971,I166954,);
nor I_9676 (I167378,I167313,I167195);
nor I_9677 (I167395,I109612,I109615);
nor I_9678 (I166945,I167395,I167378);
not I_9679 (I167426,I167395);
nand I_9680 (I166948,I167155,I167426);
DFFARX1 I_9681 (I167395,I2859,I166971,I166960,);
DFFARX1 I_9682 (I167395,I2859,I166971,I166957,);
not I_9683 (I167515,I2866);
DFFARX1 I_9684 (I351806,I2859,I167515,I167541,);
DFFARX1 I_9685 (I167541,I2859,I167515,I167558,);
not I_9686 (I167507,I167558);
not I_9687 (I167580,I167541);
nand I_9688 (I167597,I351800,I351797);
and I_9689 (I167614,I167597,I351812);
DFFARX1 I_9690 (I167614,I2859,I167515,I167640,);
not I_9691 (I167648,I167640);
DFFARX1 I_9692 (I351800,I2859,I167515,I167674,);
and I_9693 (I167682,I167674,I351794);
nand I_9694 (I167699,I167674,I351794);
nand I_9695 (I167486,I167648,I167699);
DFFARX1 I_9696 (I351794,I2859,I167515,I167739,);
nor I_9697 (I167747,I167739,I167682);
DFFARX1 I_9698 (I167747,I2859,I167515,I167480,);
nor I_9699 (I167495,I167739,I167640);
nand I_9700 (I167792,I351809,I351803);
and I_9701 (I167809,I167792,I351797);
DFFARX1 I_9702 (I167809,I2859,I167515,I167835,);
nor I_9703 (I167483,I167835,I167739);
not I_9704 (I167857,I167835);
nor I_9705 (I167874,I167857,I167648);
nor I_9706 (I167891,I167580,I167874);
DFFARX1 I_9707 (I167891,I2859,I167515,I167498,);
nor I_9708 (I167922,I167857,I167739);
nor I_9709 (I167939,I351815,I351803);
nor I_9710 (I167489,I167939,I167922);
not I_9711 (I167970,I167939);
nand I_9712 (I167492,I167699,I167970);
DFFARX1 I_9713 (I167939,I2859,I167515,I167504,);
DFFARX1 I_9714 (I167939,I2859,I167515,I167501,);
not I_9715 (I168059,I2866);
DFFARX1 I_9716 (I298995,I2859,I168059,I168085,);
DFFARX1 I_9717 (I168085,I2859,I168059,I168102,);
not I_9718 (I168051,I168102);
not I_9719 (I168124,I168085);
nand I_9720 (I168141,I299016,I299007);
and I_9721 (I168158,I168141,I298995);
DFFARX1 I_9722 (I168158,I2859,I168059,I168184,);
not I_9723 (I168192,I168184);
DFFARX1 I_9724 (I299001,I2859,I168059,I168218,);
and I_9725 (I168226,I168218,I298998);
nand I_9726 (I168243,I168218,I298998);
nand I_9727 (I168030,I168192,I168243);
DFFARX1 I_9728 (I298992,I2859,I168059,I168283,);
nor I_9729 (I168291,I168283,I168226);
DFFARX1 I_9730 (I168291,I2859,I168059,I168024,);
nor I_9731 (I168039,I168283,I168184);
nand I_9732 (I168336,I298992,I299004);
and I_9733 (I168353,I168336,I299013);
DFFARX1 I_9734 (I168353,I2859,I168059,I168379,);
nor I_9735 (I168027,I168379,I168283);
not I_9736 (I168401,I168379);
nor I_9737 (I168418,I168401,I168192);
nor I_9738 (I168435,I168124,I168418);
DFFARX1 I_9739 (I168435,I2859,I168059,I168042,);
nor I_9740 (I168466,I168401,I168283);
nor I_9741 (I168483,I299010,I299004);
nor I_9742 (I168033,I168483,I168466);
not I_9743 (I168514,I168483);
nand I_9744 (I168036,I168243,I168514);
DFFARX1 I_9745 (I168483,I2859,I168059,I168048,);
DFFARX1 I_9746 (I168483,I2859,I168059,I168045,);
not I_9747 (I168603,I2866);
DFFARX1 I_9748 (I444685,I2859,I168603,I168629,);
DFFARX1 I_9749 (I168629,I2859,I168603,I168646,);
not I_9750 (I168595,I168646);
not I_9751 (I168668,I168629);
nand I_9752 (I168685,I444697,I444685);
and I_9753 (I168702,I168685,I444688);
DFFARX1 I_9754 (I168702,I2859,I168603,I168728,);
not I_9755 (I168736,I168728);
DFFARX1 I_9756 (I444706,I2859,I168603,I168762,);
and I_9757 (I168770,I168762,I444682);
nand I_9758 (I168787,I168762,I444682);
nand I_9759 (I168574,I168736,I168787);
DFFARX1 I_9760 (I444700,I2859,I168603,I168827,);
nor I_9761 (I168835,I168827,I168770);
DFFARX1 I_9762 (I168835,I2859,I168603,I168568,);
nor I_9763 (I168583,I168827,I168728);
nand I_9764 (I168880,I444694,I444691);
and I_9765 (I168897,I168880,I444703);
DFFARX1 I_9766 (I168897,I2859,I168603,I168923,);
nor I_9767 (I168571,I168923,I168827);
not I_9768 (I168945,I168923);
nor I_9769 (I168962,I168945,I168736);
nor I_9770 (I168979,I168668,I168962);
DFFARX1 I_9771 (I168979,I2859,I168603,I168586,);
nor I_9772 (I169010,I168945,I168827);
nor I_9773 (I169027,I444682,I444691);
nor I_9774 (I168577,I169027,I169010);
not I_9775 (I169058,I169027);
nand I_9776 (I168580,I168787,I169058);
DFFARX1 I_9777 (I169027,I2859,I168603,I168592,);
DFFARX1 I_9778 (I169027,I2859,I168603,I168589,);
not I_9779 (I169147,I2866);
DFFARX1 I_9780 (I511733,I2859,I169147,I169173,);
DFFARX1 I_9781 (I169173,I2859,I169147,I169190,);
not I_9782 (I169139,I169190);
not I_9783 (I169212,I169173);
nand I_9784 (I169229,I511745,I511748);
and I_9785 (I169246,I169229,I511751);
DFFARX1 I_9786 (I169246,I2859,I169147,I169272,);
not I_9787 (I169280,I169272);
DFFARX1 I_9788 (I511736,I2859,I169147,I169306,);
and I_9789 (I169314,I169306,I511742);
nand I_9790 (I169331,I169306,I511742);
nand I_9791 (I169118,I169280,I169331);
DFFARX1 I_9792 (I511730,I2859,I169147,I169371,);
nor I_9793 (I169379,I169371,I169314);
DFFARX1 I_9794 (I169379,I2859,I169147,I169112,);
nor I_9795 (I169127,I169371,I169272);
nand I_9796 (I169424,I511733,I511754);
and I_9797 (I169441,I169424,I511739);
DFFARX1 I_9798 (I169441,I2859,I169147,I169467,);
nor I_9799 (I169115,I169467,I169371);
not I_9800 (I169489,I169467);
nor I_9801 (I169506,I169489,I169280);
nor I_9802 (I169523,I169212,I169506);
DFFARX1 I_9803 (I169523,I2859,I169147,I169130,);
nor I_9804 (I169554,I169489,I169371);
nor I_9805 (I169571,I511730,I511754);
nor I_9806 (I169121,I169571,I169554);
not I_9807 (I169602,I169571);
nand I_9808 (I169124,I169331,I169602);
DFFARX1 I_9809 (I169571,I2859,I169147,I169136,);
DFFARX1 I_9810 (I169571,I2859,I169147,I169133,);
not I_9811 (I169691,I2866);
DFFARX1 I_9812 (I481677,I2859,I169691,I169717,);
DFFARX1 I_9813 (I169717,I2859,I169691,I169734,);
not I_9814 (I169683,I169734);
not I_9815 (I169756,I169717);
nand I_9816 (I169773,I481689,I481677);
and I_9817 (I169790,I169773,I481680);
DFFARX1 I_9818 (I169790,I2859,I169691,I169816,);
not I_9819 (I169824,I169816);
DFFARX1 I_9820 (I481698,I2859,I169691,I169850,);
and I_9821 (I169858,I169850,I481674);
nand I_9822 (I169875,I169850,I481674);
nand I_9823 (I169662,I169824,I169875);
DFFARX1 I_9824 (I481692,I2859,I169691,I169915,);
nor I_9825 (I169923,I169915,I169858);
DFFARX1 I_9826 (I169923,I2859,I169691,I169656,);
nor I_9827 (I169671,I169915,I169816);
nand I_9828 (I169968,I481686,I481683);
and I_9829 (I169985,I169968,I481695);
DFFARX1 I_9830 (I169985,I2859,I169691,I170011,);
nor I_9831 (I169659,I170011,I169915);
not I_9832 (I170033,I170011);
nor I_9833 (I170050,I170033,I169824);
nor I_9834 (I170067,I169756,I170050);
DFFARX1 I_9835 (I170067,I2859,I169691,I169674,);
nor I_9836 (I170098,I170033,I169915);
nor I_9837 (I170115,I481674,I481683);
nor I_9838 (I169665,I170115,I170098);
not I_9839 (I170146,I170115);
nand I_9840 (I169668,I169875,I170146);
DFFARX1 I_9841 (I170115,I2859,I169691,I169680,);
DFFARX1 I_9842 (I170115,I2859,I169691,I169677,);
not I_9843 (I170235,I2866);
DFFARX1 I_9844 (I539807,I2859,I170235,I170261,);
DFFARX1 I_9845 (I170261,I2859,I170235,I170278,);
not I_9846 (I170227,I170278);
not I_9847 (I170300,I170261);
nand I_9848 (I170317,I539783,I539804);
and I_9849 (I170334,I170317,I539801);
DFFARX1 I_9850 (I170334,I2859,I170235,I170360,);
not I_9851 (I170368,I170360);
DFFARX1 I_9852 (I539780,I2859,I170235,I170394,);
and I_9853 (I170402,I170394,I539792);
nand I_9854 (I170419,I170394,I539792);
nand I_9855 (I170206,I170368,I170419);
DFFARX1 I_9856 (I539795,I2859,I170235,I170459,);
nor I_9857 (I170467,I170459,I170402);
DFFARX1 I_9858 (I170467,I2859,I170235,I170200,);
nor I_9859 (I170215,I170459,I170360);
nand I_9860 (I170512,I539798,I539786);
and I_9861 (I170529,I170512,I539789);
DFFARX1 I_9862 (I170529,I2859,I170235,I170555,);
nor I_9863 (I170203,I170555,I170459);
not I_9864 (I170577,I170555);
nor I_9865 (I170594,I170577,I170368);
nor I_9866 (I170611,I170300,I170594);
DFFARX1 I_9867 (I170611,I2859,I170235,I170218,);
nor I_9868 (I170642,I170577,I170459);
nor I_9869 (I170659,I539780,I539786);
nor I_9870 (I170209,I170659,I170642);
not I_9871 (I170690,I170659);
nand I_9872 (I170212,I170419,I170690);
DFFARX1 I_9873 (I170659,I2859,I170235,I170224,);
DFFARX1 I_9874 (I170659,I2859,I170235,I170221,);
not I_9875 (I170779,I2866);
DFFARX1 I_9876 (I412201,I2859,I170779,I170805,);
DFFARX1 I_9877 (I170805,I2859,I170779,I170822,);
not I_9878 (I170771,I170822);
not I_9879 (I170844,I170805);
nand I_9880 (I170861,I412216,I412204);
and I_9881 (I170878,I170861,I412195);
DFFARX1 I_9882 (I170878,I2859,I170779,I170904,);
not I_9883 (I170912,I170904);
DFFARX1 I_9884 (I412207,I2859,I170779,I170938,);
and I_9885 (I170946,I170938,I412198);
nand I_9886 (I170963,I170938,I412198);
nand I_9887 (I170750,I170912,I170963);
DFFARX1 I_9888 (I412213,I2859,I170779,I171003,);
nor I_9889 (I171011,I171003,I170946);
DFFARX1 I_9890 (I171011,I2859,I170779,I170744,);
nor I_9891 (I170759,I171003,I170904);
nand I_9892 (I171056,I412222,I412210);
and I_9893 (I171073,I171056,I412219);
DFFARX1 I_9894 (I171073,I2859,I170779,I171099,);
nor I_9895 (I170747,I171099,I171003);
not I_9896 (I171121,I171099);
nor I_9897 (I171138,I171121,I170912);
nor I_9898 (I171155,I170844,I171138);
DFFARX1 I_9899 (I171155,I2859,I170779,I170762,);
nor I_9900 (I171186,I171121,I171003);
nor I_9901 (I171203,I412195,I412210);
nor I_9902 (I170753,I171203,I171186);
not I_9903 (I171234,I171203);
nand I_9904 (I170756,I170963,I171234);
DFFARX1 I_9905 (I171203,I2859,I170779,I170768,);
DFFARX1 I_9906 (I171203,I2859,I170779,I170765,);
not I_9907 (I171323,I2866);
DFFARX1 I_9908 (I406387,I2859,I171323,I171349,);
DFFARX1 I_9909 (I171349,I2859,I171323,I171366,);
not I_9910 (I171315,I171366);
not I_9911 (I171388,I171349);
nand I_9912 (I171405,I406402,I406390);
and I_9913 (I171422,I171405,I406381);
DFFARX1 I_9914 (I171422,I2859,I171323,I171448,);
not I_9915 (I171456,I171448);
DFFARX1 I_9916 (I406393,I2859,I171323,I171482,);
and I_9917 (I171490,I171482,I406384);
nand I_9918 (I171507,I171482,I406384);
nand I_9919 (I171294,I171456,I171507);
DFFARX1 I_9920 (I406399,I2859,I171323,I171547,);
nor I_9921 (I171555,I171547,I171490);
DFFARX1 I_9922 (I171555,I2859,I171323,I171288,);
nor I_9923 (I171303,I171547,I171448);
nand I_9924 (I171600,I406408,I406396);
and I_9925 (I171617,I171600,I406405);
DFFARX1 I_9926 (I171617,I2859,I171323,I171643,);
nor I_9927 (I171291,I171643,I171547);
not I_9928 (I171665,I171643);
nor I_9929 (I171682,I171665,I171456);
nor I_9930 (I171699,I171388,I171682);
DFFARX1 I_9931 (I171699,I2859,I171323,I171306,);
nor I_9932 (I171730,I171665,I171547);
nor I_9933 (I171747,I406381,I406396);
nor I_9934 (I171297,I171747,I171730);
not I_9935 (I171778,I171747);
nand I_9936 (I171300,I171507,I171778);
DFFARX1 I_9937 (I171747,I2859,I171323,I171312,);
DFFARX1 I_9938 (I171747,I2859,I171323,I171309,);
not I_9939 (I171867,I2866);
DFFARX1 I_9940 (I414779,I2859,I171867,I171893,);
DFFARX1 I_9941 (I171893,I2859,I171867,I171910,);
not I_9942 (I171859,I171910);
not I_9943 (I171932,I171893);
nand I_9944 (I171949,I414779,I414797);
and I_9945 (I171966,I171949,I414791);
DFFARX1 I_9946 (I171966,I2859,I171867,I171992,);
not I_9947 (I172000,I171992);
DFFARX1 I_9948 (I414785,I2859,I171867,I172026,);
and I_9949 (I172034,I172026,I414794);
nand I_9950 (I172051,I172026,I414794);
nand I_9951 (I171838,I172000,I172051);
DFFARX1 I_9952 (I414782,I2859,I171867,I172091,);
nor I_9953 (I172099,I172091,I172034);
DFFARX1 I_9954 (I172099,I2859,I171867,I171832,);
nor I_9955 (I171847,I172091,I171992);
nand I_9956 (I172144,I414782,I414800);
and I_9957 (I172161,I172144,I414785);
DFFARX1 I_9958 (I172161,I2859,I171867,I172187,);
nor I_9959 (I171835,I172187,I172091);
not I_9960 (I172209,I172187);
nor I_9961 (I172226,I172209,I172000);
nor I_9962 (I172243,I171932,I172226);
DFFARX1 I_9963 (I172243,I2859,I171867,I171850,);
nor I_9964 (I172274,I172209,I172091);
nor I_9965 (I172291,I414788,I414800);
nor I_9966 (I171841,I172291,I172274);
not I_9967 (I172322,I172291);
nand I_9968 (I171844,I172051,I172322);
DFFARX1 I_9969 (I172291,I2859,I171867,I171856,);
DFFARX1 I_9970 (I172291,I2859,I171867,I171853,);
not I_9971 (I172411,I2866);
DFFARX1 I_9972 (I146200,I2859,I172411,I172437,);
DFFARX1 I_9973 (I172437,I2859,I172411,I172454,);
not I_9974 (I172403,I172454);
not I_9975 (I172476,I172437);
nand I_9976 (I172493,I146179,I146203);
and I_9977 (I172510,I172493,I146206);
DFFARX1 I_9978 (I172510,I2859,I172411,I172536,);
not I_9979 (I172544,I172536);
DFFARX1 I_9980 (I146188,I2859,I172411,I172570,);
and I_9981 (I172578,I172570,I146194);
nand I_9982 (I172595,I172570,I146194);
nand I_9983 (I172382,I172544,I172595);
DFFARX1 I_9984 (I146182,I2859,I172411,I172635,);
nor I_9985 (I172643,I172635,I172578);
DFFARX1 I_9986 (I172643,I2859,I172411,I172376,);
nor I_9987 (I172391,I172635,I172536);
nand I_9988 (I172688,I146191,I146179);
and I_9989 (I172705,I172688,I146185);
DFFARX1 I_9990 (I172705,I2859,I172411,I172731,);
nor I_9991 (I172379,I172731,I172635);
not I_9992 (I172753,I172731);
nor I_9993 (I172770,I172753,I172544);
nor I_9994 (I172787,I172476,I172770);
DFFARX1 I_9995 (I172787,I2859,I172411,I172394,);
nor I_9996 (I172818,I172753,I172635);
nor I_9997 (I172835,I146197,I146179);
nor I_9998 (I172385,I172835,I172818);
not I_9999 (I172866,I172835);
nand I_10000 (I172388,I172595,I172866);
DFFARX1 I_10001 (I172835,I2859,I172411,I172400,);
DFFARX1 I_10002 (I172835,I2859,I172411,I172397,);
not I_10003 (I172955,I2866);
DFFARX1 I_10004 (I382485,I2859,I172955,I172981,);
DFFARX1 I_10005 (I172981,I2859,I172955,I172998,);
not I_10006 (I172947,I172998);
not I_10007 (I173020,I172981);
nand I_10008 (I173037,I382500,I382488);
and I_10009 (I173054,I173037,I382479);
DFFARX1 I_10010 (I173054,I2859,I172955,I173080,);
not I_10011 (I173088,I173080);
DFFARX1 I_10012 (I382491,I2859,I172955,I173114,);
and I_10013 (I173122,I173114,I382482);
nand I_10014 (I173139,I173114,I382482);
nand I_10015 (I172926,I173088,I173139);
DFFARX1 I_10016 (I382497,I2859,I172955,I173179,);
nor I_10017 (I173187,I173179,I173122);
DFFARX1 I_10018 (I173187,I2859,I172955,I172920,);
nor I_10019 (I172935,I173179,I173080);
nand I_10020 (I173232,I382506,I382494);
and I_10021 (I173249,I173232,I382503);
DFFARX1 I_10022 (I173249,I2859,I172955,I173275,);
nor I_10023 (I172923,I173275,I173179);
not I_10024 (I173297,I173275);
nor I_10025 (I173314,I173297,I173088);
nor I_10026 (I173331,I173020,I173314);
DFFARX1 I_10027 (I173331,I2859,I172955,I172938,);
nor I_10028 (I173362,I173297,I173179);
nor I_10029 (I173379,I382479,I382494);
nor I_10030 (I172929,I173379,I173362);
not I_10031 (I173410,I173379);
nand I_10032 (I172932,I173139,I173410);
DFFARX1 I_10033 (I173379,I2859,I172955,I172944,);
DFFARX1 I_10034 (I173379,I2859,I172955,I172941,);
not I_10035 (I173499,I2866);
DFFARX1 I_10036 (I159902,I2859,I173499,I173525,);
DFFARX1 I_10037 (I173525,I2859,I173499,I173542,);
not I_10038 (I173491,I173542);
not I_10039 (I173564,I173525);
nand I_10040 (I173581,I159881,I159905);
and I_10041 (I173598,I173581,I159908);
DFFARX1 I_10042 (I173598,I2859,I173499,I173624,);
not I_10043 (I173632,I173624);
DFFARX1 I_10044 (I159890,I2859,I173499,I173658,);
and I_10045 (I173666,I173658,I159896);
nand I_10046 (I173683,I173658,I159896);
nand I_10047 (I173470,I173632,I173683);
DFFARX1 I_10048 (I159884,I2859,I173499,I173723,);
nor I_10049 (I173731,I173723,I173666);
DFFARX1 I_10050 (I173731,I2859,I173499,I173464,);
nor I_10051 (I173479,I173723,I173624);
nand I_10052 (I173776,I159893,I159881);
and I_10053 (I173793,I173776,I159887);
DFFARX1 I_10054 (I173793,I2859,I173499,I173819,);
nor I_10055 (I173467,I173819,I173723);
not I_10056 (I173841,I173819);
nor I_10057 (I173858,I173841,I173632);
nor I_10058 (I173875,I173564,I173858);
DFFARX1 I_10059 (I173875,I2859,I173499,I173482,);
nor I_10060 (I173906,I173841,I173723);
nor I_10061 (I173923,I159899,I159881);
nor I_10062 (I173473,I173923,I173906);
not I_10063 (I173954,I173923);
nand I_10064 (I173476,I173683,I173954);
DFFARX1 I_10065 (I173923,I2859,I173499,I173488,);
DFFARX1 I_10066 (I173923,I2859,I173499,I173485,);
not I_10067 (I174043,I2866);
DFFARX1 I_10068 (I348644,I2859,I174043,I174069,);
DFFARX1 I_10069 (I174069,I2859,I174043,I174086,);
not I_10070 (I174035,I174086);
not I_10071 (I174108,I174069);
nand I_10072 (I174125,I348638,I348635);
and I_10073 (I174142,I174125,I348650);
DFFARX1 I_10074 (I174142,I2859,I174043,I174168,);
not I_10075 (I174176,I174168);
DFFARX1 I_10076 (I348638,I2859,I174043,I174202,);
and I_10077 (I174210,I174202,I348632);
nand I_10078 (I174227,I174202,I348632);
nand I_10079 (I174014,I174176,I174227);
DFFARX1 I_10080 (I348632,I2859,I174043,I174267,);
nor I_10081 (I174275,I174267,I174210);
DFFARX1 I_10082 (I174275,I2859,I174043,I174008,);
nor I_10083 (I174023,I174267,I174168);
nand I_10084 (I174320,I348647,I348641);
and I_10085 (I174337,I174320,I348635);
DFFARX1 I_10086 (I174337,I2859,I174043,I174363,);
nor I_10087 (I174011,I174363,I174267);
not I_10088 (I174385,I174363);
nor I_10089 (I174402,I174385,I174176);
nor I_10090 (I174419,I174108,I174402);
DFFARX1 I_10091 (I174419,I2859,I174043,I174026,);
nor I_10092 (I174450,I174385,I174267);
nor I_10093 (I174467,I348653,I348641);
nor I_10094 (I174017,I174467,I174450);
not I_10095 (I174498,I174467);
nand I_10096 (I174020,I174227,I174498);
DFFARX1 I_10097 (I174467,I2859,I174043,I174032,);
DFFARX1 I_10098 (I174467,I2859,I174043,I174029,);
not I_10099 (I174587,I2866);
DFFARX1 I_10100 (I500751,I2859,I174587,I174613,);
DFFARX1 I_10101 (I174613,I2859,I174587,I174630,);
not I_10102 (I174579,I174630);
not I_10103 (I174652,I174613);
nand I_10104 (I174669,I500763,I500751);
and I_10105 (I174686,I174669,I500754);
DFFARX1 I_10106 (I174686,I2859,I174587,I174712,);
not I_10107 (I174720,I174712);
DFFARX1 I_10108 (I500772,I2859,I174587,I174746,);
and I_10109 (I174754,I174746,I500748);
nand I_10110 (I174771,I174746,I500748);
nand I_10111 (I174558,I174720,I174771);
DFFARX1 I_10112 (I500766,I2859,I174587,I174811,);
nor I_10113 (I174819,I174811,I174754);
DFFARX1 I_10114 (I174819,I2859,I174587,I174552,);
nor I_10115 (I174567,I174811,I174712);
nand I_10116 (I174864,I500760,I500757);
and I_10117 (I174881,I174864,I500769);
DFFARX1 I_10118 (I174881,I2859,I174587,I174907,);
nor I_10119 (I174555,I174907,I174811);
not I_10120 (I174929,I174907);
nor I_10121 (I174946,I174929,I174720);
nor I_10122 (I174963,I174652,I174946);
DFFARX1 I_10123 (I174963,I2859,I174587,I174570,);
nor I_10124 (I174994,I174929,I174811);
nor I_10125 (I175011,I500748,I500757);
nor I_10126 (I174561,I175011,I174994);
not I_10127 (I175042,I175011);
nand I_10128 (I174564,I174771,I175042);
DFFARX1 I_10129 (I175011,I2859,I174587,I174576,);
DFFARX1 I_10130 (I175011,I2859,I174587,I174573,);
not I_10131 (I175131,I2866);
DFFARX1 I_10132 (I85821,I2859,I175131,I175157,);
DFFARX1 I_10133 (I175157,I2859,I175131,I175174,);
not I_10134 (I175123,I175174);
not I_10135 (I175196,I175157);
nand I_10136 (I175213,I85833,I85812);
and I_10137 (I175230,I175213,I85815);
DFFARX1 I_10138 (I175230,I2859,I175131,I175256,);
not I_10139 (I175264,I175256);
DFFARX1 I_10140 (I85824,I2859,I175131,I175290,);
and I_10141 (I175298,I175290,I85836);
nand I_10142 (I175315,I175290,I85836);
nand I_10143 (I175102,I175264,I175315);
DFFARX1 I_10144 (I85830,I2859,I175131,I175355,);
nor I_10145 (I175363,I175355,I175298);
DFFARX1 I_10146 (I175363,I2859,I175131,I175096,);
nor I_10147 (I175111,I175355,I175256);
nand I_10148 (I175408,I85818,I85815);
and I_10149 (I175425,I175408,I85827);
DFFARX1 I_10150 (I175425,I2859,I175131,I175451,);
nor I_10151 (I175099,I175451,I175355);
not I_10152 (I175473,I175451);
nor I_10153 (I175490,I175473,I175264);
nor I_10154 (I175507,I175196,I175490);
DFFARX1 I_10155 (I175507,I2859,I175131,I175114,);
nor I_10156 (I175538,I175473,I175355);
nor I_10157 (I175555,I85812,I85815);
nor I_10158 (I175105,I175555,I175538);
not I_10159 (I175586,I175555);
nand I_10160 (I175108,I175315,I175586);
DFFARX1 I_10161 (I175555,I2859,I175131,I175120,);
DFFARX1 I_10162 (I175555,I2859,I175131,I175117,);
not I_10163 (I175675,I2866);
DFFARX1 I_10164 (I446997,I2859,I175675,I175701,);
DFFARX1 I_10165 (I175701,I2859,I175675,I175718,);
not I_10166 (I175667,I175718);
not I_10167 (I175740,I175701);
nand I_10168 (I175757,I447009,I446997);
and I_10169 (I175774,I175757,I447000);
DFFARX1 I_10170 (I175774,I2859,I175675,I175800,);
not I_10171 (I175808,I175800);
DFFARX1 I_10172 (I447018,I2859,I175675,I175834,);
and I_10173 (I175842,I175834,I446994);
nand I_10174 (I175859,I175834,I446994);
nand I_10175 (I175646,I175808,I175859);
DFFARX1 I_10176 (I447012,I2859,I175675,I175899,);
nor I_10177 (I175907,I175899,I175842);
DFFARX1 I_10178 (I175907,I2859,I175675,I175640,);
nor I_10179 (I175655,I175899,I175800);
nand I_10180 (I175952,I447006,I447003);
and I_10181 (I175969,I175952,I447015);
DFFARX1 I_10182 (I175969,I2859,I175675,I175995,);
nor I_10183 (I175643,I175995,I175899);
not I_10184 (I176017,I175995);
nor I_10185 (I176034,I176017,I175808);
nor I_10186 (I176051,I175740,I176034);
DFFARX1 I_10187 (I176051,I2859,I175675,I175658,);
nor I_10188 (I176082,I176017,I175899);
nor I_10189 (I176099,I446994,I447003);
nor I_10190 (I175649,I176099,I176082);
not I_10191 (I176130,I176099);
nand I_10192 (I175652,I175859,I176130);
DFFARX1 I_10193 (I176099,I2859,I175675,I175664,);
DFFARX1 I_10194 (I176099,I2859,I175675,I175661,);
not I_10195 (I176219,I2866);
DFFARX1 I_10196 (I545162,I2859,I176219,I176245,);
DFFARX1 I_10197 (I176245,I2859,I176219,I176262,);
not I_10198 (I176211,I176262);
not I_10199 (I176284,I176245);
nand I_10200 (I176301,I545138,I545159);
and I_10201 (I176318,I176301,I545156);
DFFARX1 I_10202 (I176318,I2859,I176219,I176344,);
not I_10203 (I176352,I176344);
DFFARX1 I_10204 (I545135,I2859,I176219,I176378,);
and I_10205 (I176386,I176378,I545147);
nand I_10206 (I176403,I176378,I545147);
nand I_10207 (I176190,I176352,I176403);
DFFARX1 I_10208 (I545150,I2859,I176219,I176443,);
nor I_10209 (I176451,I176443,I176386);
DFFARX1 I_10210 (I176451,I2859,I176219,I176184,);
nor I_10211 (I176199,I176443,I176344);
nand I_10212 (I176496,I545153,I545141);
and I_10213 (I176513,I176496,I545144);
DFFARX1 I_10214 (I176513,I2859,I176219,I176539,);
nor I_10215 (I176187,I176539,I176443);
not I_10216 (I176561,I176539);
nor I_10217 (I176578,I176561,I176352);
nor I_10218 (I176595,I176284,I176578);
DFFARX1 I_10219 (I176595,I2859,I176219,I176202,);
nor I_10220 (I176626,I176561,I176443);
nor I_10221 (I176643,I545135,I545141);
nor I_10222 (I176193,I176643,I176626);
not I_10223 (I176674,I176643);
nand I_10224 (I176196,I176403,I176674);
DFFARX1 I_10225 (I176643,I2859,I176219,I176208,);
DFFARX1 I_10226 (I176643,I2859,I176219,I176205,);
not I_10227 (I176763,I2866);
DFFARX1 I_10228 (I37997,I2859,I176763,I176789,);
DFFARX1 I_10229 (I176789,I2859,I176763,I176806,);
not I_10230 (I176755,I176806);
not I_10231 (I176828,I176789);
nand I_10232 (I176845,I38012,I37991);
and I_10233 (I176862,I176845,I37994);
DFFARX1 I_10234 (I176862,I2859,I176763,I176888,);
not I_10235 (I176896,I176888);
DFFARX1 I_10236 (I38000,I2859,I176763,I176922,);
and I_10237 (I176930,I176922,I37994);
nand I_10238 (I176947,I176922,I37994);
nand I_10239 (I176734,I176896,I176947);
DFFARX1 I_10240 (I38009,I2859,I176763,I176987,);
nor I_10241 (I176995,I176987,I176930);
DFFARX1 I_10242 (I176995,I2859,I176763,I176728,);
nor I_10243 (I176743,I176987,I176888);
nand I_10244 (I177040,I37991,I38006);
and I_10245 (I177057,I177040,I38003);
DFFARX1 I_10246 (I177057,I2859,I176763,I177083,);
nor I_10247 (I176731,I177083,I176987);
not I_10248 (I177105,I177083);
nor I_10249 (I177122,I177105,I176896);
nor I_10250 (I177139,I176828,I177122);
DFFARX1 I_10251 (I177139,I2859,I176763,I176746,);
nor I_10252 (I177170,I177105,I176987);
nor I_10253 (I177187,I38015,I38006);
nor I_10254 (I176737,I177187,I177170);
not I_10255 (I177218,I177187);
nand I_10256 (I176740,I176947,I177218);
DFFARX1 I_10257 (I177187,I2859,I176763,I176752,);
DFFARX1 I_10258 (I177187,I2859,I176763,I176749,);
not I_10259 (I177307,I2866);
DFFARX1 I_10260 (I158848,I2859,I177307,I177333,);
DFFARX1 I_10261 (I177333,I2859,I177307,I177350,);
not I_10262 (I177299,I177350);
not I_10263 (I177372,I177333);
nand I_10264 (I177389,I158827,I158851);
and I_10265 (I177406,I177389,I158854);
DFFARX1 I_10266 (I177406,I2859,I177307,I177432,);
not I_10267 (I177440,I177432);
DFFARX1 I_10268 (I158836,I2859,I177307,I177466,);
and I_10269 (I177474,I177466,I158842);
nand I_10270 (I177491,I177466,I158842);
nand I_10271 (I177278,I177440,I177491);
DFFARX1 I_10272 (I158830,I2859,I177307,I177531,);
nor I_10273 (I177539,I177531,I177474);
DFFARX1 I_10274 (I177539,I2859,I177307,I177272,);
nor I_10275 (I177287,I177531,I177432);
nand I_10276 (I177584,I158839,I158827);
and I_10277 (I177601,I177584,I158833);
DFFARX1 I_10278 (I177601,I2859,I177307,I177627,);
nor I_10279 (I177275,I177627,I177531);
not I_10280 (I177649,I177627);
nor I_10281 (I177666,I177649,I177440);
nor I_10282 (I177683,I177372,I177666);
DFFARX1 I_10283 (I177683,I2859,I177307,I177290,);
nor I_10284 (I177714,I177649,I177531);
nor I_10285 (I177731,I158845,I158827);
nor I_10286 (I177281,I177731,I177714);
not I_10287 (I177762,I177731);
nand I_10288 (I177284,I177491,I177762);
DFFARX1 I_10289 (I177731,I2859,I177307,I177296,);
DFFARX1 I_10290 (I177731,I2859,I177307,I177293,);
not I_10291 (I177851,I2866);
DFFARX1 I_10292 (I296683,I2859,I177851,I177877,);
DFFARX1 I_10293 (I177877,I2859,I177851,I177894,);
not I_10294 (I177843,I177894);
not I_10295 (I177916,I177877);
nand I_10296 (I177933,I296704,I296695);
and I_10297 (I177950,I177933,I296683);
DFFARX1 I_10298 (I177950,I2859,I177851,I177976,);
not I_10299 (I177984,I177976);
DFFARX1 I_10300 (I296689,I2859,I177851,I178010,);
and I_10301 (I178018,I178010,I296686);
nand I_10302 (I178035,I178010,I296686);
nand I_10303 (I177822,I177984,I178035);
DFFARX1 I_10304 (I296680,I2859,I177851,I178075,);
nor I_10305 (I178083,I178075,I178018);
DFFARX1 I_10306 (I178083,I2859,I177851,I177816,);
nor I_10307 (I177831,I178075,I177976);
nand I_10308 (I178128,I296680,I296692);
and I_10309 (I178145,I178128,I296701);
DFFARX1 I_10310 (I178145,I2859,I177851,I178171,);
nor I_10311 (I177819,I178171,I178075);
not I_10312 (I178193,I178171);
nor I_10313 (I178210,I178193,I177984);
nor I_10314 (I178227,I177916,I178210);
DFFARX1 I_10315 (I178227,I2859,I177851,I177834,);
nor I_10316 (I178258,I178193,I178075);
nor I_10317 (I178275,I296698,I296692);
nor I_10318 (I177825,I178275,I178258);
not I_10319 (I178306,I178275);
nand I_10320 (I177828,I178035,I178306);
DFFARX1 I_10321 (I178275,I2859,I177851,I177840,);
DFFARX1 I_10322 (I178275,I2859,I177851,I177837,);
not I_10323 (I178395,I2866);
DFFARX1 I_10324 (I115107,I2859,I178395,I178421,);
DFFARX1 I_10325 (I178421,I2859,I178395,I178438,);
not I_10326 (I178387,I178438);
not I_10327 (I178460,I178421);
nand I_10328 (I178477,I115086,I115110);
and I_10329 (I178494,I178477,I115113);
DFFARX1 I_10330 (I178494,I2859,I178395,I178520,);
not I_10331 (I178528,I178520);
DFFARX1 I_10332 (I115095,I2859,I178395,I178554,);
and I_10333 (I178562,I178554,I115101);
nand I_10334 (I178579,I178554,I115101);
nand I_10335 (I178366,I178528,I178579);
DFFARX1 I_10336 (I115089,I2859,I178395,I178619,);
nor I_10337 (I178627,I178619,I178562);
DFFARX1 I_10338 (I178627,I2859,I178395,I178360,);
nor I_10339 (I178375,I178619,I178520);
nand I_10340 (I178672,I115098,I115086);
and I_10341 (I178689,I178672,I115092);
DFFARX1 I_10342 (I178689,I2859,I178395,I178715,);
nor I_10343 (I178363,I178715,I178619);
not I_10344 (I178737,I178715);
nor I_10345 (I178754,I178737,I178528);
nor I_10346 (I178771,I178460,I178754);
DFFARX1 I_10347 (I178771,I2859,I178395,I178378,);
nor I_10348 (I178802,I178737,I178619);
nor I_10349 (I178819,I115104,I115086);
nor I_10350 (I178369,I178819,I178802);
not I_10351 (I178850,I178819);
nand I_10352 (I178372,I178579,I178850);
DFFARX1 I_10353 (I178819,I2859,I178395,I178384,);
DFFARX1 I_10354 (I178819,I2859,I178395,I178381,);
not I_10355 (I178939,I2866);
DFFARX1 I_10356 (I290325,I2859,I178939,I178965,);
DFFARX1 I_10357 (I178965,I2859,I178939,I178982,);
not I_10358 (I178931,I178982);
not I_10359 (I179004,I178965);
nand I_10360 (I179021,I290346,I290337);
and I_10361 (I179038,I179021,I290325);
DFFARX1 I_10362 (I179038,I2859,I178939,I179064,);
not I_10363 (I179072,I179064);
DFFARX1 I_10364 (I290331,I2859,I178939,I179098,);
and I_10365 (I179106,I179098,I290328);
nand I_10366 (I179123,I179098,I290328);
nand I_10367 (I178910,I179072,I179123);
DFFARX1 I_10368 (I290322,I2859,I178939,I179163,);
nor I_10369 (I179171,I179163,I179106);
DFFARX1 I_10370 (I179171,I2859,I178939,I178904,);
nor I_10371 (I178919,I179163,I179064);
nand I_10372 (I179216,I290322,I290334);
and I_10373 (I179233,I179216,I290343);
DFFARX1 I_10374 (I179233,I2859,I178939,I179259,);
nor I_10375 (I178907,I179259,I179163);
not I_10376 (I179281,I179259);
nor I_10377 (I179298,I179281,I179072);
nor I_10378 (I179315,I179004,I179298);
DFFARX1 I_10379 (I179315,I2859,I178939,I178922,);
nor I_10380 (I179346,I179281,I179163);
nor I_10381 (I179363,I290340,I290334);
nor I_10382 (I178913,I179363,I179346);
not I_10383 (I179394,I179363);
nand I_10384 (I178916,I179123,I179394);
DFFARX1 I_10385 (I179363,I2859,I178939,I178928,);
DFFARX1 I_10386 (I179363,I2859,I178939,I178925,);
not I_10387 (I179483,I2866);
DFFARX1 I_10388 (I82846,I2859,I179483,I179509,);
DFFARX1 I_10389 (I179509,I2859,I179483,I179526,);
not I_10390 (I179475,I179526);
not I_10391 (I179548,I179509);
nand I_10392 (I179565,I82858,I82837);
and I_10393 (I179582,I179565,I82840);
DFFARX1 I_10394 (I179582,I2859,I179483,I179608,);
not I_10395 (I179616,I179608);
DFFARX1 I_10396 (I82849,I2859,I179483,I179642,);
and I_10397 (I179650,I179642,I82861);
nand I_10398 (I179667,I179642,I82861);
nand I_10399 (I179454,I179616,I179667);
DFFARX1 I_10400 (I82855,I2859,I179483,I179707,);
nor I_10401 (I179715,I179707,I179650);
DFFARX1 I_10402 (I179715,I2859,I179483,I179448,);
nor I_10403 (I179463,I179707,I179608);
nand I_10404 (I179760,I82843,I82840);
and I_10405 (I179777,I179760,I82852);
DFFARX1 I_10406 (I179777,I2859,I179483,I179803,);
nor I_10407 (I179451,I179803,I179707);
not I_10408 (I179825,I179803);
nor I_10409 (I179842,I179825,I179616);
nor I_10410 (I179859,I179548,I179842);
DFFARX1 I_10411 (I179859,I2859,I179483,I179466,);
nor I_10412 (I179890,I179825,I179707);
nor I_10413 (I179907,I82837,I82840);
nor I_10414 (I179457,I179907,I179890);
not I_10415 (I179938,I179907);
nand I_10416 (I179460,I179667,I179938);
DFFARX1 I_10417 (I179907,I2859,I179483,I179472,);
DFFARX1 I_10418 (I179907,I2859,I179483,I179469,);
not I_10419 (I180027,I2866);
DFFARX1 I_10420 (I542782,I2859,I180027,I180053,);
DFFARX1 I_10421 (I180053,I2859,I180027,I180070,);
not I_10422 (I180019,I180070);
not I_10423 (I180092,I180053);
nand I_10424 (I180109,I542758,I542779);
and I_10425 (I180126,I180109,I542776);
DFFARX1 I_10426 (I180126,I2859,I180027,I180152,);
not I_10427 (I180160,I180152);
DFFARX1 I_10428 (I542755,I2859,I180027,I180186,);
and I_10429 (I180194,I180186,I542767);
nand I_10430 (I180211,I180186,I542767);
nand I_10431 (I179998,I180160,I180211);
DFFARX1 I_10432 (I542770,I2859,I180027,I180251,);
nor I_10433 (I180259,I180251,I180194);
DFFARX1 I_10434 (I180259,I2859,I180027,I179992,);
nor I_10435 (I180007,I180251,I180152);
nand I_10436 (I180304,I542773,I542761);
and I_10437 (I180321,I180304,I542764);
DFFARX1 I_10438 (I180321,I2859,I180027,I180347,);
nor I_10439 (I179995,I180347,I180251);
not I_10440 (I180369,I180347);
nor I_10441 (I180386,I180369,I180160);
nor I_10442 (I180403,I180092,I180386);
DFFARX1 I_10443 (I180403,I2859,I180027,I180010,);
nor I_10444 (I180434,I180369,I180251);
nor I_10445 (I180451,I542755,I542761);
nor I_10446 (I180001,I180451,I180434);
not I_10447 (I180482,I180451);
nand I_10448 (I180004,I180211,I180482);
DFFARX1 I_10449 (I180451,I2859,I180027,I180016,);
DFFARX1 I_10450 (I180451,I2859,I180027,I180013,);
not I_10451 (I180571,I2866);
DFFARX1 I_10452 (I360238,I2859,I180571,I180597,);
DFFARX1 I_10453 (I180597,I2859,I180571,I180614,);
not I_10454 (I180563,I180614);
not I_10455 (I180636,I180597);
nand I_10456 (I180653,I360232,I360229);
and I_10457 (I180670,I180653,I360244);
DFFARX1 I_10458 (I180670,I2859,I180571,I180696,);
not I_10459 (I180704,I180696);
DFFARX1 I_10460 (I360232,I2859,I180571,I180730,);
and I_10461 (I180738,I180730,I360226);
nand I_10462 (I180755,I180730,I360226);
nand I_10463 (I180542,I180704,I180755);
DFFARX1 I_10464 (I360226,I2859,I180571,I180795,);
nor I_10465 (I180803,I180795,I180738);
DFFARX1 I_10466 (I180803,I2859,I180571,I180536,);
nor I_10467 (I180551,I180795,I180696);
nand I_10468 (I180848,I360241,I360235);
and I_10469 (I180865,I180848,I360229);
DFFARX1 I_10470 (I180865,I2859,I180571,I180891,);
nor I_10471 (I180539,I180891,I180795);
not I_10472 (I180913,I180891);
nor I_10473 (I180930,I180913,I180704);
nor I_10474 (I180947,I180636,I180930);
DFFARX1 I_10475 (I180947,I2859,I180571,I180554,);
nor I_10476 (I180978,I180913,I180795);
nor I_10477 (I180995,I360247,I360235);
nor I_10478 (I180545,I180995,I180978);
not I_10479 (I181026,I180995);
nand I_10480 (I180548,I180755,I181026);
DFFARX1 I_10481 (I180995,I2859,I180571,I180560,);
DFFARX1 I_10482 (I180995,I2859,I180571,I180557,);
not I_10483 (I181115,I2866);
DFFARX1 I_10484 (I116161,I2859,I181115,I181141,);
DFFARX1 I_10485 (I181141,I2859,I181115,I181158,);
not I_10486 (I181107,I181158);
not I_10487 (I181180,I181141);
nand I_10488 (I181197,I116140,I116164);
and I_10489 (I181214,I181197,I116167);
DFFARX1 I_10490 (I181214,I2859,I181115,I181240,);
not I_10491 (I181248,I181240);
DFFARX1 I_10492 (I116149,I2859,I181115,I181274,);
and I_10493 (I181282,I181274,I116155);
nand I_10494 (I181299,I181274,I116155);
nand I_10495 (I181086,I181248,I181299);
DFFARX1 I_10496 (I116143,I2859,I181115,I181339,);
nor I_10497 (I181347,I181339,I181282);
DFFARX1 I_10498 (I181347,I2859,I181115,I181080,);
nor I_10499 (I181095,I181339,I181240);
nand I_10500 (I181392,I116152,I116140);
and I_10501 (I181409,I181392,I116146);
DFFARX1 I_10502 (I181409,I2859,I181115,I181435,);
nor I_10503 (I181083,I181435,I181339);
not I_10504 (I181457,I181435);
nor I_10505 (I181474,I181457,I181248);
nor I_10506 (I181491,I181180,I181474);
DFFARX1 I_10507 (I181491,I2859,I181115,I181098,);
nor I_10508 (I181522,I181457,I181339);
nor I_10509 (I181539,I116158,I116140);
nor I_10510 (I181089,I181539,I181522);
not I_10511 (I181570,I181539);
nand I_10512 (I181092,I181299,I181570);
DFFARX1 I_10513 (I181539,I2859,I181115,I181104,);
DFFARX1 I_10514 (I181539,I2859,I181115,I181101,);
not I_10515 (I181659,I2866);
DFFARX1 I_10516 (I446419,I2859,I181659,I181685,);
DFFARX1 I_10517 (I181685,I2859,I181659,I181702,);
not I_10518 (I181651,I181702);
not I_10519 (I181724,I181685);
nand I_10520 (I181741,I446431,I446419);
and I_10521 (I181758,I181741,I446422);
DFFARX1 I_10522 (I181758,I2859,I181659,I181784,);
not I_10523 (I181792,I181784);
DFFARX1 I_10524 (I446440,I2859,I181659,I181818,);
and I_10525 (I181826,I181818,I446416);
nand I_10526 (I181843,I181818,I446416);
nand I_10527 (I181630,I181792,I181843);
DFFARX1 I_10528 (I446434,I2859,I181659,I181883,);
nor I_10529 (I181891,I181883,I181826);
DFFARX1 I_10530 (I181891,I2859,I181659,I181624,);
nor I_10531 (I181639,I181883,I181784);
nand I_10532 (I181936,I446428,I446425);
and I_10533 (I181953,I181936,I446437);
DFFARX1 I_10534 (I181953,I2859,I181659,I181979,);
nor I_10535 (I181627,I181979,I181883);
not I_10536 (I182001,I181979);
nor I_10537 (I182018,I182001,I181792);
nor I_10538 (I182035,I181724,I182018);
DFFARX1 I_10539 (I182035,I2859,I181659,I181642,);
nor I_10540 (I182066,I182001,I181883);
nor I_10541 (I182083,I446416,I446425);
nor I_10542 (I181633,I182083,I182066);
not I_10543 (I182114,I182083);
nand I_10544 (I181636,I181843,I182114);
DFFARX1 I_10545 (I182083,I2859,I181659,I181648,);
DFFARX1 I_10546 (I182083,I2859,I181659,I181645,);
not I_10547 (I182203,I2866);
DFFARX1 I_10548 (I364397,I2859,I182203,I182229,);
DFFARX1 I_10549 (I182229,I2859,I182203,I182246,);
not I_10550 (I182195,I182246);
not I_10551 (I182268,I182229);
nand I_10552 (I182285,I364412,I364400);
and I_10553 (I182302,I182285,I364391);
DFFARX1 I_10554 (I182302,I2859,I182203,I182328,);
not I_10555 (I182336,I182328);
DFFARX1 I_10556 (I364403,I2859,I182203,I182362,);
and I_10557 (I182370,I182362,I364394);
nand I_10558 (I182387,I182362,I364394);
nand I_10559 (I182174,I182336,I182387);
DFFARX1 I_10560 (I364409,I2859,I182203,I182427,);
nor I_10561 (I182435,I182427,I182370);
DFFARX1 I_10562 (I182435,I2859,I182203,I182168,);
nor I_10563 (I182183,I182427,I182328);
nand I_10564 (I182480,I364418,I364406);
and I_10565 (I182497,I182480,I364415);
DFFARX1 I_10566 (I182497,I2859,I182203,I182523,);
nor I_10567 (I182171,I182523,I182427);
not I_10568 (I182545,I182523);
nor I_10569 (I182562,I182545,I182336);
nor I_10570 (I182579,I182268,I182562);
DFFARX1 I_10571 (I182579,I2859,I182203,I182186,);
nor I_10572 (I182610,I182545,I182427);
nor I_10573 (I182627,I364391,I364406);
nor I_10574 (I182177,I182627,I182610);
not I_10575 (I182658,I182627);
nand I_10576 (I182180,I182387,I182658);
DFFARX1 I_10577 (I182627,I2859,I182203,I182192,);
DFFARX1 I_10578 (I182627,I2859,I182203,I182189,);
not I_10579 (I182747,I2866);
DFFARX1 I_10580 (I497861,I2859,I182747,I182773,);
DFFARX1 I_10581 (I182773,I2859,I182747,I182790,);
not I_10582 (I182739,I182790);
not I_10583 (I182812,I182773);
nand I_10584 (I182829,I497873,I497861);
and I_10585 (I182846,I182829,I497864);
DFFARX1 I_10586 (I182846,I2859,I182747,I182872,);
not I_10587 (I182880,I182872);
DFFARX1 I_10588 (I497882,I2859,I182747,I182906,);
and I_10589 (I182914,I182906,I497858);
nand I_10590 (I182931,I182906,I497858);
nand I_10591 (I182718,I182880,I182931);
DFFARX1 I_10592 (I497876,I2859,I182747,I182971,);
nor I_10593 (I182979,I182971,I182914);
DFFARX1 I_10594 (I182979,I2859,I182747,I182712,);
nor I_10595 (I182727,I182971,I182872);
nand I_10596 (I183024,I497870,I497867);
and I_10597 (I183041,I183024,I497879);
DFFARX1 I_10598 (I183041,I2859,I182747,I183067,);
nor I_10599 (I182715,I183067,I182971);
not I_10600 (I183089,I183067);
nor I_10601 (I183106,I183089,I182880);
nor I_10602 (I183123,I182812,I183106);
DFFARX1 I_10603 (I183123,I2859,I182747,I182730,);
nor I_10604 (I183154,I183089,I182971);
nor I_10605 (I183171,I497858,I497867);
nor I_10606 (I182721,I183171,I183154);
not I_10607 (I183202,I183171);
nand I_10608 (I182724,I182931,I183202);
DFFARX1 I_10609 (I183171,I2859,I182747,I182736,);
DFFARX1 I_10610 (I183171,I2859,I182747,I182733,);
not I_10611 (I183291,I2866);
DFFARX1 I_10612 (I492081,I2859,I183291,I183317,);
DFFARX1 I_10613 (I183317,I2859,I183291,I183334,);
not I_10614 (I183283,I183334);
not I_10615 (I183356,I183317);
nand I_10616 (I183373,I492093,I492081);
and I_10617 (I183390,I183373,I492084);
DFFARX1 I_10618 (I183390,I2859,I183291,I183416,);
not I_10619 (I183424,I183416);
DFFARX1 I_10620 (I492102,I2859,I183291,I183450,);
and I_10621 (I183458,I183450,I492078);
nand I_10622 (I183475,I183450,I492078);
nand I_10623 (I183262,I183424,I183475);
DFFARX1 I_10624 (I492096,I2859,I183291,I183515,);
nor I_10625 (I183523,I183515,I183458);
DFFARX1 I_10626 (I183523,I2859,I183291,I183256,);
nor I_10627 (I183271,I183515,I183416);
nand I_10628 (I183568,I492090,I492087);
and I_10629 (I183585,I183568,I492099);
DFFARX1 I_10630 (I183585,I2859,I183291,I183611,);
nor I_10631 (I183259,I183611,I183515);
not I_10632 (I183633,I183611);
nor I_10633 (I183650,I183633,I183424);
nor I_10634 (I183667,I183356,I183650);
DFFARX1 I_10635 (I183667,I2859,I183291,I183274,);
nor I_10636 (I183698,I183633,I183515);
nor I_10637 (I183715,I492078,I492087);
nor I_10638 (I183265,I183715,I183698);
not I_10639 (I183746,I183715);
nand I_10640 (I183268,I183475,I183746);
DFFARX1 I_10641 (I183715,I2859,I183291,I183280,);
DFFARX1 I_10642 (I183715,I2859,I183291,I183277,);
not I_10643 (I183835,I2866);
DFFARX1 I_10644 (I488035,I2859,I183835,I183861,);
DFFARX1 I_10645 (I183861,I2859,I183835,I183878,);
not I_10646 (I183827,I183878);
not I_10647 (I183900,I183861);
nand I_10648 (I183917,I488047,I488035);
and I_10649 (I183934,I183917,I488038);
DFFARX1 I_10650 (I183934,I2859,I183835,I183960,);
not I_10651 (I183968,I183960);
DFFARX1 I_10652 (I488056,I2859,I183835,I183994,);
and I_10653 (I184002,I183994,I488032);
nand I_10654 (I184019,I183994,I488032);
nand I_10655 (I183806,I183968,I184019);
DFFARX1 I_10656 (I488050,I2859,I183835,I184059,);
nor I_10657 (I184067,I184059,I184002);
DFFARX1 I_10658 (I184067,I2859,I183835,I183800,);
nor I_10659 (I183815,I184059,I183960);
nand I_10660 (I184112,I488044,I488041);
and I_10661 (I184129,I184112,I488053);
DFFARX1 I_10662 (I184129,I2859,I183835,I184155,);
nor I_10663 (I183803,I184155,I184059);
not I_10664 (I184177,I184155);
nor I_10665 (I184194,I184177,I183968);
nor I_10666 (I184211,I183900,I184194);
DFFARX1 I_10667 (I184211,I2859,I183835,I183818,);
nor I_10668 (I184242,I184177,I184059);
nor I_10669 (I184259,I488032,I488041);
nor I_10670 (I183809,I184259,I184242);
not I_10671 (I184290,I184259);
nand I_10672 (I183812,I184019,I184290);
DFFARX1 I_10673 (I184259,I2859,I183835,I183824,);
DFFARX1 I_10674 (I184259,I2859,I183835,I183821,);
not I_10675 (I184379,I2866);
DFFARX1 I_10676 (I569557,I2859,I184379,I184405,);
DFFARX1 I_10677 (I184405,I2859,I184379,I184422,);
not I_10678 (I184371,I184422);
not I_10679 (I184444,I184405);
nand I_10680 (I184461,I569533,I569554);
and I_10681 (I184478,I184461,I569551);
DFFARX1 I_10682 (I184478,I2859,I184379,I184504,);
not I_10683 (I184512,I184504);
DFFARX1 I_10684 (I569530,I2859,I184379,I184538,);
and I_10685 (I184546,I184538,I569542);
nand I_10686 (I184563,I184538,I569542);
nand I_10687 (I184350,I184512,I184563);
DFFARX1 I_10688 (I569545,I2859,I184379,I184603,);
nor I_10689 (I184611,I184603,I184546);
DFFARX1 I_10690 (I184611,I2859,I184379,I184344,);
nor I_10691 (I184359,I184603,I184504);
nand I_10692 (I184656,I569548,I569536);
and I_10693 (I184673,I184656,I569539);
DFFARX1 I_10694 (I184673,I2859,I184379,I184699,);
nor I_10695 (I184347,I184699,I184603);
not I_10696 (I184721,I184699);
nor I_10697 (I184738,I184721,I184512);
nor I_10698 (I184755,I184444,I184738);
DFFARX1 I_10699 (I184755,I2859,I184379,I184362,);
nor I_10700 (I184786,I184721,I184603);
nor I_10701 (I184803,I569530,I569536);
nor I_10702 (I184353,I184803,I184786);
not I_10703 (I184834,I184803);
nand I_10704 (I184356,I184563,I184834);
DFFARX1 I_10705 (I184803,I2859,I184379,I184368,);
DFFARX1 I_10706 (I184803,I2859,I184379,I184365,);
not I_10707 (I184923,I2866);
DFFARX1 I_10708 (I1860,I2859,I184923,I184949,);
DFFARX1 I_10709 (I184949,I2859,I184923,I184966,);
not I_10710 (I184915,I184966);
not I_10711 (I184988,I184949);
nand I_10712 (I185005,I2348,I1972);
and I_10713 (I185022,I185005,I2540);
DFFARX1 I_10714 (I185022,I2859,I184923,I185048,);
not I_10715 (I185056,I185048);
DFFARX1 I_10716 (I1540,I2859,I184923,I185082,);
and I_10717 (I185090,I185082,I2212);
nand I_10718 (I185107,I185082,I2212);
nand I_10719 (I184894,I185056,I185107);
DFFARX1 I_10720 (I2036,I2859,I184923,I185147,);
nor I_10721 (I185155,I185147,I185090);
DFFARX1 I_10722 (I185155,I2859,I184923,I184888,);
nor I_10723 (I184903,I185147,I185048);
nand I_10724 (I185200,I2004,I2636);
and I_10725 (I185217,I185200,I2148);
DFFARX1 I_10726 (I185217,I2859,I184923,I185243,);
nor I_10727 (I184891,I185243,I185147);
not I_10728 (I185265,I185243);
nor I_10729 (I185282,I185265,I185056);
nor I_10730 (I185299,I184988,I185282);
DFFARX1 I_10731 (I185299,I2859,I184923,I184906,);
nor I_10732 (I185330,I185265,I185147);
nor I_10733 (I185347,I2404,I2636);
nor I_10734 (I184897,I185347,I185330);
not I_10735 (I185378,I185347);
nand I_10736 (I184900,I185107,I185378);
DFFARX1 I_10737 (I185347,I2859,I184923,I184912,);
DFFARX1 I_10738 (I185347,I2859,I184923,I184909,);
not I_10739 (I185467,I2866);
DFFARX1 I_10740 (I248131,I2859,I185467,I185493,);
DFFARX1 I_10741 (I185493,I2859,I185467,I185510,);
not I_10742 (I185459,I185510);
not I_10743 (I185532,I185493);
nand I_10744 (I185549,I248128,I248149);
and I_10745 (I185566,I185549,I248152);
DFFARX1 I_10746 (I185566,I2859,I185467,I185592,);
not I_10747 (I185600,I185592);
DFFARX1 I_10748 (I248137,I2859,I185467,I185626,);
and I_10749 (I185634,I185626,I248140);
nand I_10750 (I185651,I185626,I248140);
nand I_10751 (I185438,I185600,I185651);
DFFARX1 I_10752 (I248143,I2859,I185467,I185691,);
nor I_10753 (I185699,I185691,I185634);
DFFARX1 I_10754 (I185699,I2859,I185467,I185432,);
nor I_10755 (I185447,I185691,I185592);
nand I_10756 (I185744,I248128,I248134);
and I_10757 (I185761,I185744,I248146);
DFFARX1 I_10758 (I185761,I2859,I185467,I185787,);
nor I_10759 (I185435,I185787,I185691);
not I_10760 (I185809,I185787);
nor I_10761 (I185826,I185809,I185600);
nor I_10762 (I185843,I185532,I185826);
DFFARX1 I_10763 (I185843,I2859,I185467,I185450,);
nor I_10764 (I185874,I185809,I185691);
nor I_10765 (I185891,I248131,I248134);
nor I_10766 (I185441,I185891,I185874);
not I_10767 (I185922,I185891);
nand I_10768 (I185444,I185651,I185922);
DFFARX1 I_10769 (I185891,I2859,I185467,I185456,);
DFFARX1 I_10770 (I185891,I2859,I185467,I185453,);
not I_10771 (I186011,I2866);
DFFARX1 I_10772 (I130390,I2859,I186011,I186037,);
DFFARX1 I_10773 (I186037,I2859,I186011,I186054,);
not I_10774 (I186003,I186054);
not I_10775 (I186076,I186037);
nand I_10776 (I186093,I130369,I130393);
and I_10777 (I186110,I186093,I130396);
DFFARX1 I_10778 (I186110,I2859,I186011,I186136,);
not I_10779 (I186144,I186136);
DFFARX1 I_10780 (I130378,I2859,I186011,I186170,);
and I_10781 (I186178,I186170,I130384);
nand I_10782 (I186195,I186170,I130384);
nand I_10783 (I185982,I186144,I186195);
DFFARX1 I_10784 (I130372,I2859,I186011,I186235,);
nor I_10785 (I186243,I186235,I186178);
DFFARX1 I_10786 (I186243,I2859,I186011,I185976,);
nor I_10787 (I185991,I186235,I186136);
nand I_10788 (I186288,I130381,I130369);
and I_10789 (I186305,I186288,I130375);
DFFARX1 I_10790 (I186305,I2859,I186011,I186331,);
nor I_10791 (I185979,I186331,I186235);
not I_10792 (I186353,I186331);
nor I_10793 (I186370,I186353,I186144);
nor I_10794 (I186387,I186076,I186370);
DFFARX1 I_10795 (I186387,I2859,I186011,I185994,);
nor I_10796 (I186418,I186353,I186235);
nor I_10797 (I186435,I130387,I130369);
nor I_10798 (I185985,I186435,I186418);
not I_10799 (I186466,I186435);
nand I_10800 (I185988,I186195,I186466);
DFFARX1 I_10801 (I186435,I2859,I186011,I186000,);
DFFARX1 I_10802 (I186435,I2859,I186011,I185997,);
not I_10803 (I186555,I2866);
DFFARX1 I_10804 (I111418,I2859,I186555,I186581,);
DFFARX1 I_10805 (I186581,I2859,I186555,I186598,);
not I_10806 (I186547,I186598);
not I_10807 (I186620,I186581);
nand I_10808 (I186637,I111397,I111421);
and I_10809 (I186654,I186637,I111424);
DFFARX1 I_10810 (I186654,I2859,I186555,I186680,);
not I_10811 (I186688,I186680);
DFFARX1 I_10812 (I111406,I2859,I186555,I186714,);
and I_10813 (I186722,I186714,I111412);
nand I_10814 (I186739,I186714,I111412);
nand I_10815 (I186526,I186688,I186739);
DFFARX1 I_10816 (I111400,I2859,I186555,I186779,);
nor I_10817 (I186787,I186779,I186722);
DFFARX1 I_10818 (I186787,I2859,I186555,I186520,);
nor I_10819 (I186535,I186779,I186680);
nand I_10820 (I186832,I111409,I111397);
and I_10821 (I186849,I186832,I111403);
DFFARX1 I_10822 (I186849,I2859,I186555,I186875,);
nor I_10823 (I186523,I186875,I186779);
not I_10824 (I186897,I186875);
nor I_10825 (I186914,I186897,I186688);
nor I_10826 (I186931,I186620,I186914);
DFFARX1 I_10827 (I186931,I2859,I186555,I186538,);
nor I_10828 (I186962,I186897,I186779);
nor I_10829 (I186979,I111415,I111397);
nor I_10830 (I186529,I186979,I186962);
not I_10831 (I187010,I186979);
nand I_10832 (I186532,I186739,I187010);
DFFARX1 I_10833 (I186979,I2859,I186555,I186544,);
DFFARX1 I_10834 (I186979,I2859,I186555,I186541,);
not I_10835 (I187099,I2866);
DFFARX1 I_10836 (I238883,I2859,I187099,I187125,);
DFFARX1 I_10837 (I187125,I2859,I187099,I187142,);
not I_10838 (I187091,I187142);
not I_10839 (I187164,I187125);
nand I_10840 (I187181,I238880,I238901);
and I_10841 (I187198,I187181,I238904);
DFFARX1 I_10842 (I187198,I2859,I187099,I187224,);
not I_10843 (I187232,I187224);
DFFARX1 I_10844 (I238889,I2859,I187099,I187258,);
and I_10845 (I187266,I187258,I238892);
nand I_10846 (I187283,I187258,I238892);
nand I_10847 (I187070,I187232,I187283);
DFFARX1 I_10848 (I238895,I2859,I187099,I187323,);
nor I_10849 (I187331,I187323,I187266);
DFFARX1 I_10850 (I187331,I2859,I187099,I187064,);
nor I_10851 (I187079,I187323,I187224);
nand I_10852 (I187376,I238880,I238886);
and I_10853 (I187393,I187376,I238898);
DFFARX1 I_10854 (I187393,I2859,I187099,I187419,);
nor I_10855 (I187067,I187419,I187323);
not I_10856 (I187441,I187419);
nor I_10857 (I187458,I187441,I187232);
nor I_10858 (I187475,I187164,I187458);
DFFARX1 I_10859 (I187475,I2859,I187099,I187082,);
nor I_10860 (I187506,I187441,I187323);
nor I_10861 (I187523,I238883,I238886);
nor I_10862 (I187073,I187523,I187506);
not I_10863 (I187554,I187523);
nand I_10864 (I187076,I187283,I187554);
DFFARX1 I_10865 (I187523,I2859,I187099,I187088,);
DFFARX1 I_10866 (I187523,I2859,I187099,I187085,);
not I_10867 (I187643,I2866);
DFFARX1 I_10868 (I507381,I2859,I187643,I187669,);
DFFARX1 I_10869 (I187669,I2859,I187643,I187686,);
not I_10870 (I187635,I187686);
not I_10871 (I187708,I187669);
nand I_10872 (I187725,I507393,I507396);
and I_10873 (I187742,I187725,I507399);
DFFARX1 I_10874 (I187742,I2859,I187643,I187768,);
not I_10875 (I187776,I187768);
DFFARX1 I_10876 (I507384,I2859,I187643,I187802,);
and I_10877 (I187810,I187802,I507390);
nand I_10878 (I187827,I187802,I507390);
nand I_10879 (I187614,I187776,I187827);
DFFARX1 I_10880 (I507378,I2859,I187643,I187867,);
nor I_10881 (I187875,I187867,I187810);
DFFARX1 I_10882 (I187875,I2859,I187643,I187608,);
nor I_10883 (I187623,I187867,I187768);
nand I_10884 (I187920,I507381,I507402);
and I_10885 (I187937,I187920,I507387);
DFFARX1 I_10886 (I187937,I2859,I187643,I187963,);
nor I_10887 (I187611,I187963,I187867);
not I_10888 (I187985,I187963);
nor I_10889 (I188002,I187985,I187776);
nor I_10890 (I188019,I187708,I188002);
DFFARX1 I_10891 (I188019,I2859,I187643,I187626,);
nor I_10892 (I188050,I187985,I187867);
nor I_10893 (I188067,I507378,I507402);
nor I_10894 (I187617,I188067,I188050);
not I_10895 (I188098,I188067);
nand I_10896 (I187620,I187827,I188098);
DFFARX1 I_10897 (I188067,I2859,I187643,I187632,);
DFFARX1 I_10898 (I188067,I2859,I187643,I187629,);
not I_10899 (I188187,I2866);
DFFARX1 I_10900 (I413493,I2859,I188187,I188213,);
DFFARX1 I_10901 (I188213,I2859,I188187,I188230,);
not I_10902 (I188179,I188230);
not I_10903 (I188252,I188213);
nand I_10904 (I188269,I413508,I413496);
and I_10905 (I188286,I188269,I413487);
DFFARX1 I_10906 (I188286,I2859,I188187,I188312,);
not I_10907 (I188320,I188312);
DFFARX1 I_10908 (I413499,I2859,I188187,I188346,);
and I_10909 (I188354,I188346,I413490);
nand I_10910 (I188371,I188346,I413490);
nand I_10911 (I188158,I188320,I188371);
DFFARX1 I_10912 (I413505,I2859,I188187,I188411,);
nor I_10913 (I188419,I188411,I188354);
DFFARX1 I_10914 (I188419,I2859,I188187,I188152,);
nor I_10915 (I188167,I188411,I188312);
nand I_10916 (I188464,I413514,I413502);
and I_10917 (I188481,I188464,I413511);
DFFARX1 I_10918 (I188481,I2859,I188187,I188507,);
nor I_10919 (I188155,I188507,I188411);
not I_10920 (I188529,I188507);
nor I_10921 (I188546,I188529,I188320);
nor I_10922 (I188563,I188252,I188546);
DFFARX1 I_10923 (I188563,I2859,I188187,I188170,);
nor I_10924 (I188594,I188529,I188411);
nor I_10925 (I188611,I413487,I413502);
nor I_10926 (I188161,I188611,I188594);
not I_10927 (I188642,I188611);
nand I_10928 (I188164,I188371,I188642);
DFFARX1 I_10929 (I188611,I2859,I188187,I188176,);
DFFARX1 I_10930 (I188611,I2859,I188187,I188173,);
not I_10931 (I188731,I2866);
DFFARX1 I_10932 (I390883,I2859,I188731,I188757,);
DFFARX1 I_10933 (I188757,I2859,I188731,I188774,);
not I_10934 (I188723,I188774);
not I_10935 (I188796,I188757);
nand I_10936 (I188813,I390898,I390886);
and I_10937 (I188830,I188813,I390877);
DFFARX1 I_10938 (I188830,I2859,I188731,I188856,);
not I_10939 (I188864,I188856);
DFFARX1 I_10940 (I390889,I2859,I188731,I188890,);
and I_10941 (I188898,I188890,I390880);
nand I_10942 (I188915,I188890,I390880);
nand I_10943 (I188702,I188864,I188915);
DFFARX1 I_10944 (I390895,I2859,I188731,I188955,);
nor I_10945 (I188963,I188955,I188898);
DFFARX1 I_10946 (I188963,I2859,I188731,I188696,);
nor I_10947 (I188711,I188955,I188856);
nand I_10948 (I189008,I390904,I390892);
and I_10949 (I189025,I189008,I390901);
DFFARX1 I_10950 (I189025,I2859,I188731,I189051,);
nor I_10951 (I188699,I189051,I188955);
not I_10952 (I189073,I189051);
nor I_10953 (I189090,I189073,I188864);
nor I_10954 (I189107,I188796,I189090);
DFFARX1 I_10955 (I189107,I2859,I188731,I188714,);
nor I_10956 (I189138,I189073,I188955);
nor I_10957 (I189155,I390877,I390892);
nor I_10958 (I188705,I189155,I189138);
not I_10959 (I189186,I189155);
nand I_10960 (I188708,I188915,I189186);
DFFARX1 I_10961 (I189155,I2859,I188731,I188720,);
DFFARX1 I_10962 (I189155,I2859,I188731,I188717,);
not I_10963 (I189275,I2866);
DFFARX1 I_10964 (I91771,I2859,I189275,I189301,);
DFFARX1 I_10965 (I189301,I2859,I189275,I189318,);
not I_10966 (I189267,I189318);
not I_10967 (I189340,I189301);
nand I_10968 (I189357,I91783,I91762);
and I_10969 (I189374,I189357,I91765);
DFFARX1 I_10970 (I189374,I2859,I189275,I189400,);
not I_10971 (I189408,I189400);
DFFARX1 I_10972 (I91774,I2859,I189275,I189434,);
and I_10973 (I189442,I189434,I91786);
nand I_10974 (I189459,I189434,I91786);
nand I_10975 (I189246,I189408,I189459);
DFFARX1 I_10976 (I91780,I2859,I189275,I189499,);
nor I_10977 (I189507,I189499,I189442);
DFFARX1 I_10978 (I189507,I2859,I189275,I189240,);
nor I_10979 (I189255,I189499,I189400);
nand I_10980 (I189552,I91768,I91765);
and I_10981 (I189569,I189552,I91777);
DFFARX1 I_10982 (I189569,I2859,I189275,I189595,);
nor I_10983 (I189243,I189595,I189499);
not I_10984 (I189617,I189595);
nor I_10985 (I189634,I189617,I189408);
nor I_10986 (I189651,I189340,I189634);
DFFARX1 I_10987 (I189651,I2859,I189275,I189258,);
nor I_10988 (I189682,I189617,I189499);
nor I_10989 (I189699,I91762,I91765);
nor I_10990 (I189249,I189699,I189682);
not I_10991 (I189730,I189699);
nand I_10992 (I189252,I189459,I189730);
DFFARX1 I_10993 (I189699,I2859,I189275,I189264,);
DFFARX1 I_10994 (I189699,I2859,I189275,I189261,);
not I_10995 (I189819,I2866);
DFFARX1 I_10996 (I528170,I2859,I189819,I189845,);
DFFARX1 I_10997 (I189845,I2859,I189819,I189862,);
not I_10998 (I189811,I189862);
not I_10999 (I189884,I189845);
nand I_11000 (I189901,I528167,I528164);
and I_11001 (I189918,I189901,I528152);
DFFARX1 I_11002 (I189918,I2859,I189819,I189944,);
not I_11003 (I189952,I189944);
DFFARX1 I_11004 (I528176,I2859,I189819,I189978,);
and I_11005 (I189986,I189978,I528161);
nand I_11006 (I190003,I189978,I528161);
nand I_11007 (I189790,I189952,I190003);
DFFARX1 I_11008 (I528155,I2859,I189819,I190043,);
nor I_11009 (I190051,I190043,I189986);
DFFARX1 I_11010 (I190051,I2859,I189819,I189784,);
nor I_11011 (I189799,I190043,I189944);
nand I_11012 (I190096,I528152,I528158);
and I_11013 (I190113,I190096,I528173);
DFFARX1 I_11014 (I190113,I2859,I189819,I190139,);
nor I_11015 (I189787,I190139,I190043);
not I_11016 (I190161,I190139);
nor I_11017 (I190178,I190161,I189952);
nor I_11018 (I190195,I189884,I190178);
DFFARX1 I_11019 (I190195,I2859,I189819,I189802,);
nor I_11020 (I190226,I190161,I190043);
nor I_11021 (I190243,I528155,I528158);
nor I_11022 (I189793,I190243,I190226);
not I_11023 (I190274,I190243);
nand I_11024 (I189796,I190003,I190274);
DFFARX1 I_11025 (I190243,I2859,I189819,I189808,);
DFFARX1 I_11026 (I190243,I2859,I189819,I189805,);
not I_11027 (I190363,I2866);
DFFARX1 I_11028 (I312867,I2859,I190363,I190389,);
DFFARX1 I_11029 (I190389,I2859,I190363,I190406,);
not I_11030 (I190355,I190406);
not I_11031 (I190428,I190389);
nand I_11032 (I190445,I312888,I312879);
and I_11033 (I190462,I190445,I312867);
DFFARX1 I_11034 (I190462,I2859,I190363,I190488,);
not I_11035 (I190496,I190488);
DFFARX1 I_11036 (I312873,I2859,I190363,I190522,);
and I_11037 (I190530,I190522,I312870);
nand I_11038 (I190547,I190522,I312870);
nand I_11039 (I190334,I190496,I190547);
DFFARX1 I_11040 (I312864,I2859,I190363,I190587,);
nor I_11041 (I190595,I190587,I190530);
DFFARX1 I_11042 (I190595,I2859,I190363,I190328,);
nor I_11043 (I190343,I190587,I190488);
nand I_11044 (I190640,I312864,I312876);
and I_11045 (I190657,I190640,I312885);
DFFARX1 I_11046 (I190657,I2859,I190363,I190683,);
nor I_11047 (I190331,I190683,I190587);
not I_11048 (I190705,I190683);
nor I_11049 (I190722,I190705,I190496);
nor I_11050 (I190739,I190428,I190722);
DFFARX1 I_11051 (I190739,I2859,I190363,I190346,);
nor I_11052 (I190770,I190705,I190587);
nor I_11053 (I190787,I312882,I312876);
nor I_11054 (I190337,I190787,I190770);
not I_11055 (I190818,I190787);
nand I_11056 (I190340,I190547,I190818);
DFFARX1 I_11057 (I190787,I2859,I190363,I190352,);
DFFARX1 I_11058 (I190787,I2859,I190363,I190349,);
not I_11059 (I190907,I2866);
DFFARX1 I_11060 (I571342,I2859,I190907,I190933,);
DFFARX1 I_11061 (I190933,I2859,I190907,I190950,);
not I_11062 (I190899,I190950);
not I_11063 (I190972,I190933);
nand I_11064 (I190989,I571318,I571339);
and I_11065 (I191006,I190989,I571336);
DFFARX1 I_11066 (I191006,I2859,I190907,I191032,);
not I_11067 (I191040,I191032);
DFFARX1 I_11068 (I571315,I2859,I190907,I191066,);
and I_11069 (I191074,I191066,I571327);
nand I_11070 (I191091,I191066,I571327);
nand I_11071 (I190878,I191040,I191091);
DFFARX1 I_11072 (I571330,I2859,I190907,I191131,);
nor I_11073 (I191139,I191131,I191074);
DFFARX1 I_11074 (I191139,I2859,I190907,I190872,);
nor I_11075 (I190887,I191131,I191032);
nand I_11076 (I191184,I571333,I571321);
and I_11077 (I191201,I191184,I571324);
DFFARX1 I_11078 (I191201,I2859,I190907,I191227,);
nor I_11079 (I190875,I191227,I191131);
not I_11080 (I191249,I191227);
nor I_11081 (I191266,I191249,I191040);
nor I_11082 (I191283,I190972,I191266);
DFFARX1 I_11083 (I191283,I2859,I190907,I190890,);
nor I_11084 (I191314,I191249,I191131);
nor I_11085 (I191331,I571315,I571321);
nor I_11086 (I190881,I191331,I191314);
not I_11087 (I191362,I191331);
nand I_11088 (I190884,I191091,I191362);
DFFARX1 I_11089 (I191331,I2859,I190907,I190896,);
DFFARX1 I_11090 (I191331,I2859,I190907,I190893,);
not I_11091 (I191451,I2866);
DFFARX1 I_11092 (I139349,I2859,I191451,I191477,);
DFFARX1 I_11093 (I191477,I2859,I191451,I191494,);
not I_11094 (I191443,I191494);
not I_11095 (I191516,I191477);
nand I_11096 (I191533,I139328,I139352);
and I_11097 (I191550,I191533,I139355);
DFFARX1 I_11098 (I191550,I2859,I191451,I191576,);
not I_11099 (I191584,I191576);
DFFARX1 I_11100 (I139337,I2859,I191451,I191610,);
and I_11101 (I191618,I191610,I139343);
nand I_11102 (I191635,I191610,I139343);
nand I_11103 (I191422,I191584,I191635);
DFFARX1 I_11104 (I139331,I2859,I191451,I191675,);
nor I_11105 (I191683,I191675,I191618);
DFFARX1 I_11106 (I191683,I2859,I191451,I191416,);
nor I_11107 (I191431,I191675,I191576);
nand I_11108 (I191728,I139340,I139328);
and I_11109 (I191745,I191728,I139334);
DFFARX1 I_11110 (I191745,I2859,I191451,I191771,);
nor I_11111 (I191419,I191771,I191675);
not I_11112 (I191793,I191771);
nor I_11113 (I191810,I191793,I191584);
nor I_11114 (I191827,I191516,I191810);
DFFARX1 I_11115 (I191827,I2859,I191451,I191434,);
nor I_11116 (I191858,I191793,I191675);
nor I_11117 (I191875,I139346,I139328);
nor I_11118 (I191425,I191875,I191858);
not I_11119 (I191906,I191875);
nand I_11120 (I191428,I191635,I191906);
DFFARX1 I_11121 (I191875,I2859,I191451,I191440,);
DFFARX1 I_11122 (I191875,I2859,I191451,I191437,);
not I_11123 (I191995,I2866);
DFFARX1 I_11124 (I79871,I2859,I191995,I192021,);
DFFARX1 I_11125 (I192021,I2859,I191995,I192038,);
not I_11126 (I191987,I192038);
not I_11127 (I192060,I192021);
nand I_11128 (I192077,I79883,I79862);
and I_11129 (I192094,I192077,I79865);
DFFARX1 I_11130 (I192094,I2859,I191995,I192120,);
not I_11131 (I192128,I192120);
DFFARX1 I_11132 (I79874,I2859,I191995,I192154,);
and I_11133 (I192162,I192154,I79886);
nand I_11134 (I192179,I192154,I79886);
nand I_11135 (I191966,I192128,I192179);
DFFARX1 I_11136 (I79880,I2859,I191995,I192219,);
nor I_11137 (I192227,I192219,I192162);
DFFARX1 I_11138 (I192227,I2859,I191995,I191960,);
nor I_11139 (I191975,I192219,I192120);
nand I_11140 (I192272,I79868,I79865);
and I_11141 (I192289,I192272,I79877);
DFFARX1 I_11142 (I192289,I2859,I191995,I192315,);
nor I_11143 (I191963,I192315,I192219);
not I_11144 (I192337,I192315);
nor I_11145 (I192354,I192337,I192128);
nor I_11146 (I192371,I192060,I192354);
DFFARX1 I_11147 (I192371,I2859,I191995,I191978,);
nor I_11148 (I192402,I192337,I192219);
nor I_11149 (I192419,I79862,I79865);
nor I_11150 (I191969,I192419,I192402);
not I_11151 (I192450,I192419);
nand I_11152 (I191972,I192179,I192450);
DFFARX1 I_11153 (I192419,I2859,I191995,I191984,);
DFFARX1 I_11154 (I192419,I2859,I191995,I191981,);
not I_11155 (I192539,I2866);
DFFARX1 I_11156 (I479365,I2859,I192539,I192565,);
DFFARX1 I_11157 (I192565,I2859,I192539,I192582,);
not I_11158 (I192531,I192582);
not I_11159 (I192604,I192565);
nand I_11160 (I192621,I479377,I479365);
and I_11161 (I192638,I192621,I479368);
DFFARX1 I_11162 (I192638,I2859,I192539,I192664,);
not I_11163 (I192672,I192664);
DFFARX1 I_11164 (I479386,I2859,I192539,I192698,);
and I_11165 (I192706,I192698,I479362);
nand I_11166 (I192723,I192698,I479362);
nand I_11167 (I192510,I192672,I192723);
DFFARX1 I_11168 (I479380,I2859,I192539,I192763,);
nor I_11169 (I192771,I192763,I192706);
DFFARX1 I_11170 (I192771,I2859,I192539,I192504,);
nor I_11171 (I192519,I192763,I192664);
nand I_11172 (I192816,I479374,I479371);
and I_11173 (I192833,I192816,I479383);
DFFARX1 I_11174 (I192833,I2859,I192539,I192859,);
nor I_11175 (I192507,I192859,I192763);
not I_11176 (I192881,I192859);
nor I_11177 (I192898,I192881,I192672);
nor I_11178 (I192915,I192604,I192898);
DFFARX1 I_11179 (I192915,I2859,I192539,I192522,);
nor I_11180 (I192946,I192881,I192763);
nor I_11181 (I192963,I479362,I479371);
nor I_11182 (I192513,I192963,I192946);
not I_11183 (I192994,I192963);
nand I_11184 (I192516,I192723,I192994);
DFFARX1 I_11185 (I192963,I2859,I192539,I192528,);
DFFARX1 I_11186 (I192963,I2859,I192539,I192525,);
not I_11187 (I193083,I2866);
DFFARX1 I_11188 (I305353,I2859,I193083,I193109,);
DFFARX1 I_11189 (I193109,I2859,I193083,I193126,);
not I_11190 (I193075,I193126);
not I_11191 (I193148,I193109);
nand I_11192 (I193165,I305374,I305365);
and I_11193 (I193182,I193165,I305353);
DFFARX1 I_11194 (I193182,I2859,I193083,I193208,);
not I_11195 (I193216,I193208);
DFFARX1 I_11196 (I305359,I2859,I193083,I193242,);
and I_11197 (I193250,I193242,I305356);
nand I_11198 (I193267,I193242,I305356);
nand I_11199 (I193054,I193216,I193267);
DFFARX1 I_11200 (I305350,I2859,I193083,I193307,);
nor I_11201 (I193315,I193307,I193250);
DFFARX1 I_11202 (I193315,I2859,I193083,I193048,);
nor I_11203 (I193063,I193307,I193208);
nand I_11204 (I193360,I305350,I305362);
and I_11205 (I193377,I193360,I305371);
DFFARX1 I_11206 (I193377,I2859,I193083,I193403,);
nor I_11207 (I193051,I193403,I193307);
not I_11208 (I193425,I193403);
nor I_11209 (I193442,I193425,I193216);
nor I_11210 (I193459,I193148,I193442);
DFFARX1 I_11211 (I193459,I2859,I193083,I193066,);
nor I_11212 (I193490,I193425,I193307);
nor I_11213 (I193507,I305368,I305362);
nor I_11214 (I193057,I193507,I193490);
not I_11215 (I193538,I193507);
nand I_11216 (I193060,I193267,I193538);
DFFARX1 I_11217 (I193507,I2859,I193083,I193072,);
DFFARX1 I_11218 (I193507,I2859,I193083,I193069,);
not I_11219 (I193627,I2866);
DFFARX1 I_11220 (I11126,I2859,I193627,I193653,);
DFFARX1 I_11221 (I193653,I2859,I193627,I193670,);
not I_11222 (I193619,I193670);
not I_11223 (I193692,I193653);
nand I_11224 (I193709,I11114,I11129);
and I_11225 (I193726,I193709,I11117);
DFFARX1 I_11226 (I193726,I2859,I193627,I193752,);
not I_11227 (I193760,I193752);
DFFARX1 I_11228 (I11138,I2859,I193627,I193786,);
and I_11229 (I193794,I193786,I11132);
nand I_11230 (I193811,I193786,I11132);
nand I_11231 (I193598,I193760,I193811);
DFFARX1 I_11232 (I11135,I2859,I193627,I193851,);
nor I_11233 (I193859,I193851,I193794);
DFFARX1 I_11234 (I193859,I2859,I193627,I193592,);
nor I_11235 (I193607,I193851,I193752);
nand I_11236 (I193904,I11114,I11117);
and I_11237 (I193921,I193904,I11120);
DFFARX1 I_11238 (I193921,I2859,I193627,I193947,);
nor I_11239 (I193595,I193947,I193851);
not I_11240 (I193969,I193947);
nor I_11241 (I193986,I193969,I193760);
nor I_11242 (I194003,I193692,I193986);
DFFARX1 I_11243 (I194003,I2859,I193627,I193610,);
nor I_11244 (I194034,I193969,I193851);
nor I_11245 (I194051,I11123,I11117);
nor I_11246 (I193601,I194051,I194034);
not I_11247 (I194082,I194051);
nand I_11248 (I193604,I193811,I194082);
DFFARX1 I_11249 (I194051,I2859,I193627,I193616,);
DFFARX1 I_11250 (I194051,I2859,I193627,I193613,);
not I_11251 (I194171,I2866);
DFFARX1 I_11252 (I148308,I2859,I194171,I194197,);
DFFARX1 I_11253 (I194197,I2859,I194171,I194214,);
not I_11254 (I194163,I194214);
not I_11255 (I194236,I194197);
nand I_11256 (I194253,I148287,I148311);
and I_11257 (I194270,I194253,I148314);
DFFARX1 I_11258 (I194270,I2859,I194171,I194296,);
not I_11259 (I194304,I194296);
DFFARX1 I_11260 (I148296,I2859,I194171,I194330,);
and I_11261 (I194338,I194330,I148302);
nand I_11262 (I194355,I194330,I148302);
nand I_11263 (I194142,I194304,I194355);
DFFARX1 I_11264 (I148290,I2859,I194171,I194395,);
nor I_11265 (I194403,I194395,I194338);
DFFARX1 I_11266 (I194403,I2859,I194171,I194136,);
nor I_11267 (I194151,I194395,I194296);
nand I_11268 (I194448,I148299,I148287);
and I_11269 (I194465,I194448,I148293);
DFFARX1 I_11270 (I194465,I2859,I194171,I194491,);
nor I_11271 (I194139,I194491,I194395);
not I_11272 (I194513,I194491);
nor I_11273 (I194530,I194513,I194304);
nor I_11274 (I194547,I194236,I194530);
DFFARX1 I_11275 (I194547,I2859,I194171,I194154,);
nor I_11276 (I194578,I194513,I194395);
nor I_11277 (I194595,I148305,I148287);
nor I_11278 (I194145,I194595,I194578);
not I_11279 (I194626,I194595);
nand I_11280 (I194148,I194355,I194626);
DFFARX1 I_11281 (I194595,I2859,I194171,I194160,);
DFFARX1 I_11282 (I194595,I2859,I194171,I194157,);
not I_11283 (I194715,I2866);
DFFARX1 I_11284 (I360765,I2859,I194715,I194741,);
DFFARX1 I_11285 (I194741,I2859,I194715,I194758,);
not I_11286 (I194707,I194758);
not I_11287 (I194780,I194741);
nand I_11288 (I194797,I360759,I360756);
and I_11289 (I194814,I194797,I360771);
DFFARX1 I_11290 (I194814,I2859,I194715,I194840,);
not I_11291 (I194848,I194840);
DFFARX1 I_11292 (I360759,I2859,I194715,I194874,);
and I_11293 (I194882,I194874,I360753);
nand I_11294 (I194899,I194874,I360753);
nand I_11295 (I194686,I194848,I194899);
DFFARX1 I_11296 (I360753,I2859,I194715,I194939,);
nor I_11297 (I194947,I194939,I194882);
DFFARX1 I_11298 (I194947,I2859,I194715,I194680,);
nor I_11299 (I194695,I194939,I194840);
nand I_11300 (I194992,I360768,I360762);
and I_11301 (I195009,I194992,I360756);
DFFARX1 I_11302 (I195009,I2859,I194715,I195035,);
nor I_11303 (I194683,I195035,I194939);
not I_11304 (I195057,I195035);
nor I_11305 (I195074,I195057,I194848);
nor I_11306 (I195091,I194780,I195074);
DFFARX1 I_11307 (I195091,I2859,I194715,I194698,);
nor I_11308 (I195122,I195057,I194939);
nor I_11309 (I195139,I360774,I360762);
nor I_11310 (I194689,I195139,I195122);
not I_11311 (I195170,I195139);
nand I_11312 (I194692,I194899,I195170);
DFFARX1 I_11313 (I195139,I2859,I194715,I194704,);
DFFARX1 I_11314 (I195139,I2859,I194715,I194701,);
not I_11315 (I195259,I2866);
DFFARX1 I_11316 (I348117,I2859,I195259,I195285,);
DFFARX1 I_11317 (I195285,I2859,I195259,I195302,);
not I_11318 (I195251,I195302);
not I_11319 (I195324,I195285);
nand I_11320 (I195341,I348111,I348108);
and I_11321 (I195358,I195341,I348123);
DFFARX1 I_11322 (I195358,I2859,I195259,I195384,);
not I_11323 (I195392,I195384);
DFFARX1 I_11324 (I348111,I2859,I195259,I195418,);
and I_11325 (I195426,I195418,I348105);
nand I_11326 (I195443,I195418,I348105);
nand I_11327 (I195230,I195392,I195443);
DFFARX1 I_11328 (I348105,I2859,I195259,I195483,);
nor I_11329 (I195491,I195483,I195426);
DFFARX1 I_11330 (I195491,I2859,I195259,I195224,);
nor I_11331 (I195239,I195483,I195384);
nand I_11332 (I195536,I348120,I348114);
and I_11333 (I195553,I195536,I348108);
DFFARX1 I_11334 (I195553,I2859,I195259,I195579,);
nor I_11335 (I195227,I195579,I195483);
not I_11336 (I195601,I195579);
nor I_11337 (I195618,I195601,I195392);
nor I_11338 (I195635,I195324,I195618);
DFFARX1 I_11339 (I195635,I2859,I195259,I195242,);
nor I_11340 (I195666,I195601,I195483);
nor I_11341 (I195683,I348126,I348114);
nor I_11342 (I195233,I195683,I195666);
not I_11343 (I195714,I195683);
nand I_11344 (I195236,I195443,I195714);
DFFARX1 I_11345 (I195683,I2859,I195259,I195248,);
DFFARX1 I_11346 (I195683,I2859,I195259,I195245,);
not I_11347 (I195803,I2866);
DFFARX1 I_11348 (I294949,I2859,I195803,I195829,);
DFFARX1 I_11349 (I195829,I2859,I195803,I195846,);
not I_11350 (I195795,I195846);
not I_11351 (I195868,I195829);
nand I_11352 (I195885,I294970,I294961);
and I_11353 (I195902,I195885,I294949);
DFFARX1 I_11354 (I195902,I2859,I195803,I195928,);
not I_11355 (I195936,I195928);
DFFARX1 I_11356 (I294955,I2859,I195803,I195962,);
and I_11357 (I195970,I195962,I294952);
nand I_11358 (I195987,I195962,I294952);
nand I_11359 (I195774,I195936,I195987);
DFFARX1 I_11360 (I294946,I2859,I195803,I196027,);
nor I_11361 (I196035,I196027,I195970);
DFFARX1 I_11362 (I196035,I2859,I195803,I195768,);
nor I_11363 (I195783,I196027,I195928);
nand I_11364 (I196080,I294946,I294958);
and I_11365 (I196097,I196080,I294967);
DFFARX1 I_11366 (I196097,I2859,I195803,I196123,);
nor I_11367 (I195771,I196123,I196027);
not I_11368 (I196145,I196123);
nor I_11369 (I196162,I196145,I195936);
nor I_11370 (I196179,I195868,I196162);
DFFARX1 I_11371 (I196179,I2859,I195803,I195786,);
nor I_11372 (I196210,I196145,I196027);
nor I_11373 (I196227,I294964,I294958);
nor I_11374 (I195777,I196227,I196210);
not I_11375 (I196258,I196227);
nand I_11376 (I195780,I195987,I196258);
DFFARX1 I_11377 (I196227,I2859,I195803,I195792,);
DFFARX1 I_11378 (I196227,I2859,I195803,I195789,);
not I_11379 (I196347,I2866);
DFFARX1 I_11380 (I493815,I2859,I196347,I196373,);
DFFARX1 I_11381 (I196373,I2859,I196347,I196390,);
not I_11382 (I196339,I196390);
not I_11383 (I196412,I196373);
nand I_11384 (I196429,I493827,I493815);
and I_11385 (I196446,I196429,I493818);
DFFARX1 I_11386 (I196446,I2859,I196347,I196472,);
not I_11387 (I196480,I196472);
DFFARX1 I_11388 (I493836,I2859,I196347,I196506,);
and I_11389 (I196514,I196506,I493812);
nand I_11390 (I196531,I196506,I493812);
nand I_11391 (I196318,I196480,I196531);
DFFARX1 I_11392 (I493830,I2859,I196347,I196571,);
nor I_11393 (I196579,I196571,I196514);
DFFARX1 I_11394 (I196579,I2859,I196347,I196312,);
nor I_11395 (I196327,I196571,I196472);
nand I_11396 (I196624,I493824,I493821);
and I_11397 (I196641,I196624,I493833);
DFFARX1 I_11398 (I196641,I2859,I196347,I196667,);
nor I_11399 (I196315,I196667,I196571);
not I_11400 (I196689,I196667);
nor I_11401 (I196706,I196689,I196480);
nor I_11402 (I196723,I196412,I196706);
DFFARX1 I_11403 (I196723,I2859,I196347,I196330,);
nor I_11404 (I196754,I196689,I196571);
nor I_11405 (I196771,I493812,I493821);
nor I_11406 (I196321,I196771,I196754);
not I_11407 (I196802,I196771);
nand I_11408 (I196324,I196531,I196802);
DFFARX1 I_11409 (I196771,I2859,I196347,I196336,);
DFFARX1 I_11410 (I196771,I2859,I196347,I196333,);
not I_11411 (I196891,I2866);
DFFARX1 I_11412 (I47483,I2859,I196891,I196917,);
DFFARX1 I_11413 (I196917,I2859,I196891,I196934,);
not I_11414 (I196883,I196934);
not I_11415 (I196956,I196917);
nand I_11416 (I196973,I47498,I47477);
and I_11417 (I196990,I196973,I47480);
DFFARX1 I_11418 (I196990,I2859,I196891,I197016,);
not I_11419 (I197024,I197016);
DFFARX1 I_11420 (I47486,I2859,I196891,I197050,);
and I_11421 (I197058,I197050,I47480);
nand I_11422 (I197075,I197050,I47480);
nand I_11423 (I196862,I197024,I197075);
DFFARX1 I_11424 (I47495,I2859,I196891,I197115,);
nor I_11425 (I197123,I197115,I197058);
DFFARX1 I_11426 (I197123,I2859,I196891,I196856,);
nor I_11427 (I196871,I197115,I197016);
nand I_11428 (I197168,I47477,I47492);
and I_11429 (I197185,I197168,I47489);
DFFARX1 I_11430 (I197185,I2859,I196891,I197211,);
nor I_11431 (I196859,I197211,I197115);
not I_11432 (I197233,I197211);
nor I_11433 (I197250,I197233,I197024);
nor I_11434 (I197267,I196956,I197250);
DFFARX1 I_11435 (I197267,I2859,I196891,I196874,);
nor I_11436 (I197298,I197233,I197115);
nor I_11437 (I197315,I47501,I47492);
nor I_11438 (I196865,I197315,I197298);
not I_11439 (I197346,I197315);
nand I_11440 (I196868,I197075,I197346);
DFFARX1 I_11441 (I197315,I2859,I196891,I196880,);
DFFARX1 I_11442 (I197315,I2859,I196891,I196877,);
not I_11443 (I197435,I2866);
DFFARX1 I_11444 (I237149,I2859,I197435,I197461,);
DFFARX1 I_11445 (I197461,I2859,I197435,I197478,);
not I_11446 (I197427,I197478);
not I_11447 (I197500,I197461);
nand I_11448 (I197517,I237146,I237167);
and I_11449 (I197534,I197517,I237170);
DFFARX1 I_11450 (I197534,I2859,I197435,I197560,);
not I_11451 (I197568,I197560);
DFFARX1 I_11452 (I237155,I2859,I197435,I197594,);
and I_11453 (I197602,I197594,I237158);
nand I_11454 (I197619,I197594,I237158);
nand I_11455 (I197406,I197568,I197619);
DFFARX1 I_11456 (I237161,I2859,I197435,I197659,);
nor I_11457 (I197667,I197659,I197602);
DFFARX1 I_11458 (I197667,I2859,I197435,I197400,);
nor I_11459 (I197415,I197659,I197560);
nand I_11460 (I197712,I237146,I237152);
and I_11461 (I197729,I197712,I237164);
DFFARX1 I_11462 (I197729,I2859,I197435,I197755,);
nor I_11463 (I197403,I197755,I197659);
not I_11464 (I197777,I197755);
nor I_11465 (I197794,I197777,I197568);
nor I_11466 (I197811,I197500,I197794);
DFFARX1 I_11467 (I197811,I2859,I197435,I197418,);
nor I_11468 (I197842,I197777,I197659);
nor I_11469 (I197859,I237149,I237152);
nor I_11470 (I197409,I197859,I197842);
not I_11471 (I197890,I197859);
nand I_11472 (I197412,I197619,I197890);
DFFARX1 I_11473 (I197859,I2859,I197435,I197424,);
DFFARX1 I_11474 (I197859,I2859,I197435,I197421,);
not I_11475 (I197979,I2866);
DFFARX1 I_11476 (I61426,I2859,I197979,I198005,);
DFFARX1 I_11477 (I198005,I2859,I197979,I198022,);
not I_11478 (I197971,I198022);
not I_11479 (I198044,I198005);
nand I_11480 (I198061,I61438,I61417);
and I_11481 (I198078,I198061,I61420);
DFFARX1 I_11482 (I198078,I2859,I197979,I198104,);
not I_11483 (I198112,I198104);
DFFARX1 I_11484 (I61429,I2859,I197979,I198138,);
and I_11485 (I198146,I198138,I61441);
nand I_11486 (I198163,I198138,I61441);
nand I_11487 (I197950,I198112,I198163);
DFFARX1 I_11488 (I61435,I2859,I197979,I198203,);
nor I_11489 (I198211,I198203,I198146);
DFFARX1 I_11490 (I198211,I2859,I197979,I197944,);
nor I_11491 (I197959,I198203,I198104);
nand I_11492 (I198256,I61423,I61420);
and I_11493 (I198273,I198256,I61432);
DFFARX1 I_11494 (I198273,I2859,I197979,I198299,);
nor I_11495 (I197947,I198299,I198203);
not I_11496 (I198321,I198299);
nor I_11497 (I198338,I198321,I198112);
nor I_11498 (I198355,I198044,I198338);
DFFARX1 I_11499 (I198355,I2859,I197979,I197962,);
nor I_11500 (I198386,I198321,I198203);
nor I_11501 (I198403,I61417,I61420);
nor I_11502 (I197953,I198403,I198386);
not I_11503 (I198434,I198403);
nand I_11504 (I197956,I198163,I198434);
DFFARX1 I_11505 (I198403,I2859,I197979,I197968,);
DFFARX1 I_11506 (I198403,I2859,I197979,I197965,);
not I_11507 (I198523,I2866);
DFFARX1 I_11508 (I495549,I2859,I198523,I198549,);
DFFARX1 I_11509 (I198549,I2859,I198523,I198566,);
not I_11510 (I198515,I198566);
not I_11511 (I198588,I198549);
nand I_11512 (I198605,I495561,I495549);
and I_11513 (I198622,I198605,I495552);
DFFARX1 I_11514 (I198622,I2859,I198523,I198648,);
not I_11515 (I198656,I198648);
DFFARX1 I_11516 (I495570,I2859,I198523,I198682,);
and I_11517 (I198690,I198682,I495546);
nand I_11518 (I198707,I198682,I495546);
nand I_11519 (I198494,I198656,I198707);
DFFARX1 I_11520 (I495564,I2859,I198523,I198747,);
nor I_11521 (I198755,I198747,I198690);
DFFARX1 I_11522 (I198755,I2859,I198523,I198488,);
nor I_11523 (I198503,I198747,I198648);
nand I_11524 (I198800,I495558,I495555);
and I_11525 (I198817,I198800,I495567);
DFFARX1 I_11526 (I198817,I2859,I198523,I198843,);
nor I_11527 (I198491,I198843,I198747);
not I_11528 (I198865,I198843);
nor I_11529 (I198882,I198865,I198656);
nor I_11530 (I198899,I198588,I198882);
DFFARX1 I_11531 (I198899,I2859,I198523,I198506,);
nor I_11532 (I198930,I198865,I198747);
nor I_11533 (I198947,I495546,I495555);
nor I_11534 (I198497,I198947,I198930);
not I_11535 (I198978,I198947);
nand I_11536 (I198500,I198707,I198978);
DFFARX1 I_11537 (I198947,I2859,I198523,I198512,);
DFFARX1 I_11538 (I198947,I2859,I198523,I198509,);
not I_11539 (I199067,I2866);
DFFARX1 I_11540 (I100696,I2859,I199067,I199093,);
DFFARX1 I_11541 (I199093,I2859,I199067,I199110,);
not I_11542 (I199059,I199110);
not I_11543 (I199132,I199093);
nand I_11544 (I199149,I100708,I100687);
and I_11545 (I199166,I199149,I100690);
DFFARX1 I_11546 (I199166,I2859,I199067,I199192,);
not I_11547 (I199200,I199192);
DFFARX1 I_11548 (I100699,I2859,I199067,I199226,);
and I_11549 (I199234,I199226,I100711);
nand I_11550 (I199251,I199226,I100711);
nand I_11551 (I199038,I199200,I199251);
DFFARX1 I_11552 (I100705,I2859,I199067,I199291,);
nor I_11553 (I199299,I199291,I199234);
DFFARX1 I_11554 (I199299,I2859,I199067,I199032,);
nor I_11555 (I199047,I199291,I199192);
nand I_11556 (I199344,I100693,I100690);
and I_11557 (I199361,I199344,I100702);
DFFARX1 I_11558 (I199361,I2859,I199067,I199387,);
nor I_11559 (I199035,I199387,I199291);
not I_11560 (I199409,I199387);
nor I_11561 (I199426,I199409,I199200);
nor I_11562 (I199443,I199132,I199426);
DFFARX1 I_11563 (I199443,I2859,I199067,I199050,);
nor I_11564 (I199474,I199409,I199291);
nor I_11565 (I199491,I100687,I100690);
nor I_11566 (I199041,I199491,I199474);
not I_11567 (I199522,I199491);
nand I_11568 (I199044,I199251,I199522);
DFFARX1 I_11569 (I199491,I2859,I199067,I199056,);
DFFARX1 I_11570 (I199491,I2859,I199067,I199053,);
not I_11571 (I199611,I2866);
DFFARX1 I_11572 (I29565,I2859,I199611,I199637,);
DFFARX1 I_11573 (I199637,I2859,I199611,I199654,);
not I_11574 (I199603,I199654);
not I_11575 (I199676,I199637);
nand I_11576 (I199693,I29580,I29559);
and I_11577 (I199710,I199693,I29562);
DFFARX1 I_11578 (I199710,I2859,I199611,I199736,);
not I_11579 (I199744,I199736);
DFFARX1 I_11580 (I29568,I2859,I199611,I199770,);
and I_11581 (I199778,I199770,I29562);
nand I_11582 (I199795,I199770,I29562);
nand I_11583 (I199582,I199744,I199795);
DFFARX1 I_11584 (I29577,I2859,I199611,I199835,);
nor I_11585 (I199843,I199835,I199778);
DFFARX1 I_11586 (I199843,I2859,I199611,I199576,);
nor I_11587 (I199591,I199835,I199736);
nand I_11588 (I199888,I29559,I29574);
and I_11589 (I199905,I199888,I29571);
DFFARX1 I_11590 (I199905,I2859,I199611,I199931,);
nor I_11591 (I199579,I199931,I199835);
not I_11592 (I199953,I199931);
nor I_11593 (I199970,I199953,I199744);
nor I_11594 (I199987,I199676,I199970);
DFFARX1 I_11595 (I199987,I2859,I199611,I199594,);
nor I_11596 (I200018,I199953,I199835);
nor I_11597 (I200035,I29583,I29574);
nor I_11598 (I199585,I200035,I200018);
not I_11599 (I200066,I200035);
nand I_11600 (I199588,I199795,I200066);
DFFARX1 I_11601 (I200035,I2859,I199611,I199600,);
DFFARX1 I_11602 (I200035,I2859,I199611,I199597,);
not I_11603 (I200152,I2866);
DFFARX1 I_11604 (I51915,I2859,I200152,I200178,);
DFFARX1 I_11605 (I200178,I2859,I200152,I200195,);
not I_11606 (I200144,I200195);
DFFARX1 I_11607 (I51903,I2859,I200152,I200226,);
not I_11608 (I200234,I51909);
nor I_11609 (I200251,I200178,I200234);
not I_11610 (I200268,I51900);
not I_11611 (I200285,I51918);
nand I_11612 (I200302,I200285,I51900);
nor I_11613 (I200319,I200234,I200302);
nor I_11614 (I200336,I200226,I200319);
DFFARX1 I_11615 (I200285,I2859,I200152,I200141,);
nor I_11616 (I200367,I51918,I51897);
nand I_11617 (I200384,I200367,I51924);
nor I_11618 (I200401,I200384,I200268);
nand I_11619 (I200126,I200401,I51909);
DFFARX1 I_11620 (I200384,I2859,I200152,I200138,);
nand I_11621 (I200446,I200268,I51918);
nor I_11622 (I200463,I200268,I51918);
nand I_11623 (I200132,I200251,I200463);
not I_11624 (I200494,I51912);
nor I_11625 (I200511,I200494,I200446);
DFFARX1 I_11626 (I200511,I2859,I200152,I200120,);
nor I_11627 (I200542,I200494,I51897);
and I_11628 (I200559,I200542,I51921);
or I_11629 (I200576,I200559,I51906);
DFFARX1 I_11630 (I200576,I2859,I200152,I200602,);
nor I_11631 (I200610,I200602,I200226);
nor I_11632 (I200129,I200178,I200610);
not I_11633 (I200641,I200602);
nor I_11634 (I200658,I200641,I200336);
DFFARX1 I_11635 (I200658,I2859,I200152,I200135,);
nand I_11636 (I200689,I200641,I200268);
nor I_11637 (I200123,I200494,I200689);
not I_11638 (I200747,I2866);
DFFARX1 I_11639 (I126168,I2859,I200747,I200773,);
DFFARX1 I_11640 (I200773,I2859,I200747,I200790,);
not I_11641 (I200739,I200790);
DFFARX1 I_11642 (I126156,I2859,I200747,I200821,);
not I_11643 (I200829,I126159);
nor I_11644 (I200846,I200773,I200829);
not I_11645 (I200863,I126162);
not I_11646 (I200880,I126174);
nand I_11647 (I200897,I200880,I126162);
nor I_11648 (I200914,I200829,I200897);
nor I_11649 (I200931,I200821,I200914);
DFFARX1 I_11650 (I200880,I2859,I200747,I200736,);
nor I_11651 (I200962,I126174,I126165);
nand I_11652 (I200979,I200962,I126153);
nor I_11653 (I200996,I200979,I200863);
nand I_11654 (I200721,I200996,I126159);
DFFARX1 I_11655 (I200979,I2859,I200747,I200733,);
nand I_11656 (I201041,I200863,I126174);
nor I_11657 (I201058,I200863,I126174);
nand I_11658 (I200727,I200846,I201058);
not I_11659 (I201089,I126171);
nor I_11660 (I201106,I201089,I201041);
DFFARX1 I_11661 (I201106,I2859,I200747,I200715,);
nor I_11662 (I201137,I201089,I126177);
and I_11663 (I201154,I201137,I126180);
or I_11664 (I201171,I201154,I126153);
DFFARX1 I_11665 (I201171,I2859,I200747,I201197,);
nor I_11666 (I201205,I201197,I200821);
nor I_11667 (I200724,I200773,I201205);
not I_11668 (I201236,I201197);
nor I_11669 (I201253,I201236,I200931);
DFFARX1 I_11670 (I201253,I2859,I200747,I200730,);
nand I_11671 (I201284,I201236,I200863);
nor I_11672 (I200718,I201089,I201284);
not I_11673 (I201342,I2866);
DFFARX1 I_11674 (I42743,I2859,I201342,I201368,);
DFFARX1 I_11675 (I201368,I2859,I201342,I201385,);
not I_11676 (I201334,I201385);
DFFARX1 I_11677 (I42755,I2859,I201342,I201416,);
not I_11678 (I201424,I42746);
nor I_11679 (I201441,I201368,I201424);
not I_11680 (I201458,I42737);
not I_11681 (I201475,I42734);
nand I_11682 (I201492,I201475,I42737);
nor I_11683 (I201509,I201424,I201492);
nor I_11684 (I201526,I201416,I201509);
DFFARX1 I_11685 (I201475,I2859,I201342,I201331,);
nor I_11686 (I201557,I42734,I42734);
nand I_11687 (I201574,I201557,I42752);
nor I_11688 (I201591,I201574,I201458);
nand I_11689 (I201316,I201591,I42746);
DFFARX1 I_11690 (I201574,I2859,I201342,I201328,);
nand I_11691 (I201636,I201458,I42734);
nor I_11692 (I201653,I201458,I42734);
nand I_11693 (I201322,I201441,I201653);
not I_11694 (I201684,I42758);
nor I_11695 (I201701,I201684,I201636);
DFFARX1 I_11696 (I201701,I2859,I201342,I201310,);
nor I_11697 (I201732,I201684,I42737);
and I_11698 (I201749,I201732,I42740);
or I_11699 (I201766,I201749,I42749);
DFFARX1 I_11700 (I201766,I2859,I201342,I201792,);
nor I_11701 (I201800,I201792,I201416);
nor I_11702 (I201319,I201368,I201800);
not I_11703 (I201831,I201792);
nor I_11704 (I201848,I201831,I201526);
DFFARX1 I_11705 (I201848,I2859,I201342,I201325,);
nand I_11706 (I201879,I201831,I201458);
nor I_11707 (I201313,I201684,I201879);
not I_11708 (I201937,I2866);
DFFARX1 I_11709 (I174552,I2859,I201937,I201963,);
DFFARX1 I_11710 (I201963,I2859,I201937,I201980,);
not I_11711 (I201929,I201980);
DFFARX1 I_11712 (I174576,I2859,I201937,I202011,);
not I_11713 (I202019,I174555);
nor I_11714 (I202036,I201963,I202019);
not I_11715 (I202053,I174561);
not I_11716 (I202070,I174567);
nand I_11717 (I202087,I202070,I174561);
nor I_11718 (I202104,I202019,I202087);
nor I_11719 (I202121,I202011,I202104);
DFFARX1 I_11720 (I202070,I2859,I201937,I201926,);
nor I_11721 (I202152,I174567,I174579);
nand I_11722 (I202169,I202152,I174573);
nor I_11723 (I202186,I202169,I202053);
nand I_11724 (I201911,I202186,I174555);
DFFARX1 I_11725 (I202169,I2859,I201937,I201923,);
nand I_11726 (I202231,I202053,I174567);
nor I_11727 (I202248,I202053,I174567);
nand I_11728 (I201917,I202036,I202248);
not I_11729 (I202279,I174558);
nor I_11730 (I202296,I202279,I202231);
DFFARX1 I_11731 (I202296,I2859,I201937,I201905,);
nor I_11732 (I202327,I202279,I174552);
and I_11733 (I202344,I202327,I174570);
or I_11734 (I202361,I202344,I174564);
DFFARX1 I_11735 (I202361,I2859,I201937,I202387,);
nor I_11736 (I202395,I202387,I202011);
nor I_11737 (I201914,I201963,I202395);
not I_11738 (I202426,I202387);
nor I_11739 (I202443,I202426,I202121);
DFFARX1 I_11740 (I202443,I2859,I201937,I201920,);
nand I_11741 (I202474,I202426,I202053);
nor I_11742 (I201908,I202279,I202474);
not I_11743 (I202532,I2866);
DFFARX1 I_11744 (I423194,I2859,I202532,I202558,);
DFFARX1 I_11745 (I202558,I2859,I202532,I202575,);
not I_11746 (I202524,I202575);
DFFARX1 I_11747 (I423197,I2859,I202532,I202606,);
not I_11748 (I202614,I423200);
nor I_11749 (I202631,I202558,I202614);
not I_11750 (I202648,I423212);
not I_11751 (I202665,I423203);
nand I_11752 (I202682,I202665,I423212);
nor I_11753 (I202699,I202614,I202682);
nor I_11754 (I202716,I202606,I202699);
DFFARX1 I_11755 (I202665,I2859,I202532,I202521,);
nor I_11756 (I202747,I423203,I423209);
nand I_11757 (I202764,I202747,I423197);
nor I_11758 (I202781,I202764,I202648);
nand I_11759 (I202506,I202781,I423200);
DFFARX1 I_11760 (I202764,I2859,I202532,I202518,);
nand I_11761 (I202826,I202648,I423203);
nor I_11762 (I202843,I202648,I423203);
nand I_11763 (I202512,I202631,I202843);
not I_11764 (I202874,I423200);
nor I_11765 (I202891,I202874,I202826);
DFFARX1 I_11766 (I202891,I2859,I202532,I202500,);
nor I_11767 (I202922,I202874,I423206);
and I_11768 (I202939,I202922,I423194);
or I_11769 (I202956,I202939,I423215);
DFFARX1 I_11770 (I202956,I2859,I202532,I202982,);
nor I_11771 (I202990,I202982,I202606);
nor I_11772 (I202509,I202558,I202990);
not I_11773 (I203021,I202982);
nor I_11774 (I203038,I203021,I202716);
DFFARX1 I_11775 (I203038,I2859,I202532,I202515,);
nand I_11776 (I203069,I203021,I202648);
nor I_11777 (I202503,I202874,I203069);
not I_11778 (I203127,I2866);
DFFARX1 I_11779 (I454526,I2859,I203127,I203153,);
DFFARX1 I_11780 (I203153,I2859,I203127,I203170,);
not I_11781 (I203119,I203170);
DFFARX1 I_11782 (I454508,I2859,I203127,I203201,);
not I_11783 (I203209,I454514);
nor I_11784 (I203226,I203153,I203209);
not I_11785 (I203243,I454529);
not I_11786 (I203260,I454520);
nand I_11787 (I203277,I203260,I454529);
nor I_11788 (I203294,I203209,I203277);
nor I_11789 (I203311,I203201,I203294);
DFFARX1 I_11790 (I203260,I2859,I203127,I203116,);
nor I_11791 (I203342,I454520,I454532);
nand I_11792 (I203359,I203342,I454511);
nor I_11793 (I203376,I203359,I203243);
nand I_11794 (I203101,I203376,I454514);
DFFARX1 I_11795 (I203359,I2859,I203127,I203113,);
nand I_11796 (I203421,I203243,I454520);
nor I_11797 (I203438,I203243,I454520);
nand I_11798 (I203107,I203226,I203438);
not I_11799 (I203469,I454517);
nor I_11800 (I203486,I203469,I203421);
DFFARX1 I_11801 (I203486,I2859,I203127,I203095,);
nor I_11802 (I203517,I203469,I454523);
and I_11803 (I203534,I203517,I454508);
or I_11804 (I203551,I203534,I454511);
DFFARX1 I_11805 (I203551,I2859,I203127,I203577,);
nor I_11806 (I203585,I203577,I203201);
nor I_11807 (I203104,I203153,I203585);
not I_11808 (I203616,I203577);
nor I_11809 (I203633,I203616,I203311);
DFFARX1 I_11810 (I203633,I2859,I203127,I203110,);
nand I_11811 (I203664,I203616,I203243);
nor I_11812 (I203098,I203469,I203664);
not I_11813 (I203722,I2866);
DFFARX1 I_11814 (I357600,I2859,I203722,I203748,);
DFFARX1 I_11815 (I203748,I2859,I203722,I203765,);
not I_11816 (I203714,I203765);
DFFARX1 I_11817 (I357597,I2859,I203722,I203796,);
not I_11818 (I203804,I357597);
nor I_11819 (I203821,I203748,I203804);
not I_11820 (I203838,I357594);
not I_11821 (I203855,I357609);
nand I_11822 (I203872,I203855,I357594);
nor I_11823 (I203889,I203804,I203872);
nor I_11824 (I203906,I203796,I203889);
DFFARX1 I_11825 (I203855,I2859,I203722,I203711,);
nor I_11826 (I203937,I357609,I357603);
nand I_11827 (I203954,I203937,I357591);
nor I_11828 (I203971,I203954,I203838);
nand I_11829 (I203696,I203971,I357597);
DFFARX1 I_11830 (I203954,I2859,I203722,I203708,);
nand I_11831 (I204016,I203838,I357609);
nor I_11832 (I204033,I203838,I357609);
nand I_11833 (I203702,I203821,I204033);
not I_11834 (I204064,I357612);
nor I_11835 (I204081,I204064,I204016);
DFFARX1 I_11836 (I204081,I2859,I203722,I203690,);
nor I_11837 (I204112,I204064,I357591);
and I_11838 (I204129,I204112,I357606);
or I_11839 (I204146,I204129,I357594);
DFFARX1 I_11840 (I204146,I2859,I203722,I204172,);
nor I_11841 (I204180,I204172,I203796);
nor I_11842 (I203699,I203748,I204180);
not I_11843 (I204211,I204172);
nor I_11844 (I204228,I204211,I203906);
DFFARX1 I_11845 (I204228,I2859,I203722,I203705,);
nand I_11846 (I204259,I204211,I203838);
nor I_11847 (I203693,I204064,I204259);
not I_11848 (I204317,I2866);
DFFARX1 I_11849 (I525271,I2859,I204317,I204343,);
DFFARX1 I_11850 (I204343,I2859,I204317,I204360,);
not I_11851 (I204309,I204360);
DFFARX1 I_11852 (I525277,I2859,I204317,I204391,);
not I_11853 (I204399,I525265);
nor I_11854 (I204416,I204343,I204399);
not I_11855 (I204433,I525268);
not I_11856 (I204450,I525274);
nand I_11857 (I204467,I204450,I525268);
nor I_11858 (I204484,I204399,I204467);
nor I_11859 (I204501,I204391,I204484);
DFFARX1 I_11860 (I204450,I2859,I204317,I204306,);
nor I_11861 (I204532,I525274,I525265);
nand I_11862 (I204549,I204532,I525283);
nor I_11863 (I204566,I204549,I204433);
nand I_11864 (I204291,I204566,I525265);
DFFARX1 I_11865 (I204549,I2859,I204317,I204303,);
nand I_11866 (I204611,I204433,I525274);
nor I_11867 (I204628,I204433,I525274);
nand I_11868 (I204297,I204416,I204628);
not I_11869 (I204659,I525262);
nor I_11870 (I204676,I204659,I204611);
DFFARX1 I_11871 (I204676,I2859,I204317,I204285,);
nor I_11872 (I204707,I204659,I525286);
and I_11873 (I204724,I204707,I525262);
or I_11874 (I204741,I204724,I525280);
DFFARX1 I_11875 (I204741,I2859,I204317,I204767,);
nor I_11876 (I204775,I204767,I204391);
nor I_11877 (I204294,I204343,I204775);
not I_11878 (I204806,I204767);
nor I_11879 (I204823,I204806,I204501);
DFFARX1 I_11880 (I204823,I2859,I204317,I204300,);
nand I_11881 (I204854,I204806,I204433);
nor I_11882 (I204288,I204659,I204854);
not I_11883 (I204912,I2866);
DFFARX1 I_11884 (I33257,I2859,I204912,I204938,);
DFFARX1 I_11885 (I204938,I2859,I204912,I204955,);
not I_11886 (I204904,I204955);
DFFARX1 I_11887 (I33269,I2859,I204912,I204986,);
not I_11888 (I204994,I33260);
nor I_11889 (I205011,I204938,I204994);
not I_11890 (I205028,I33251);
not I_11891 (I205045,I33248);
nand I_11892 (I205062,I205045,I33251);
nor I_11893 (I205079,I204994,I205062);
nor I_11894 (I205096,I204986,I205079);
DFFARX1 I_11895 (I205045,I2859,I204912,I204901,);
nor I_11896 (I205127,I33248,I33248);
nand I_11897 (I205144,I205127,I33266);
nor I_11898 (I205161,I205144,I205028);
nand I_11899 (I204886,I205161,I33260);
DFFARX1 I_11900 (I205144,I2859,I204912,I204898,);
nand I_11901 (I205206,I205028,I33248);
nor I_11902 (I205223,I205028,I33248);
nand I_11903 (I204892,I205011,I205223);
not I_11904 (I205254,I33272);
nor I_11905 (I205271,I205254,I205206);
DFFARX1 I_11906 (I205271,I2859,I204912,I204880,);
nor I_11907 (I205302,I205254,I33251);
and I_11908 (I205319,I205302,I33254);
or I_11909 (I205336,I205319,I33263);
DFFARX1 I_11910 (I205336,I2859,I204912,I205362,);
nor I_11911 (I205370,I205362,I204986);
nor I_11912 (I204889,I204938,I205370);
not I_11913 (I205401,I205362);
nor I_11914 (I205418,I205401,I205096);
DFFARX1 I_11915 (I205418,I2859,I204912,I204895,);
nand I_11916 (I205449,I205401,I205028);
nor I_11917 (I204883,I205254,I205449);
not I_11918 (I205507,I2866);
DFFARX1 I_11919 (I506290,I2859,I205507,I205533,);
DFFARX1 I_11920 (I205533,I2859,I205507,I205550,);
not I_11921 (I205499,I205550);
DFFARX1 I_11922 (I506305,I2859,I205507,I205581,);
not I_11923 (I205589,I506314);
nor I_11924 (I205606,I205533,I205589);
not I_11925 (I205623,I506293);
not I_11926 (I205640,I506299);
nand I_11927 (I205657,I205640,I506293);
nor I_11928 (I205674,I205589,I205657);
nor I_11929 (I205691,I205581,I205674);
DFFARX1 I_11930 (I205640,I2859,I205507,I205496,);
nor I_11931 (I205722,I506299,I506311);
nand I_11932 (I205739,I205722,I506308);
nor I_11933 (I205756,I205739,I205623);
nand I_11934 (I205481,I205756,I506314);
DFFARX1 I_11935 (I205739,I2859,I205507,I205493,);
nand I_11936 (I205801,I205623,I506299);
nor I_11937 (I205818,I205623,I506299);
nand I_11938 (I205487,I205606,I205818);
not I_11939 (I205849,I506290);
nor I_11940 (I205866,I205849,I205801);
DFFARX1 I_11941 (I205866,I2859,I205507,I205475,);
nor I_11942 (I205897,I205849,I506302);
and I_11943 (I205914,I205897,I506296);
or I_11944 (I205931,I205914,I506293);
DFFARX1 I_11945 (I205931,I2859,I205507,I205957,);
nor I_11946 (I205965,I205957,I205581);
nor I_11947 (I205484,I205533,I205965);
not I_11948 (I205996,I205957);
nor I_11949 (I206013,I205996,I205691);
DFFARX1 I_11950 (I206013,I2859,I205507,I205490,);
nand I_11951 (I206044,I205996,I205623);
nor I_11952 (I205478,I205849,I206044);
not I_11953 (I206102,I2866);
DFFARX1 I_11954 (I196312,I2859,I206102,I206128,);
DFFARX1 I_11955 (I206128,I2859,I206102,I206145,);
not I_11956 (I206094,I206145);
DFFARX1 I_11957 (I196336,I2859,I206102,I206176,);
not I_11958 (I206184,I196315);
nor I_11959 (I206201,I206128,I206184);
not I_11960 (I206218,I196321);
not I_11961 (I206235,I196327);
nand I_11962 (I206252,I206235,I196321);
nor I_11963 (I206269,I206184,I206252);
nor I_11964 (I206286,I206176,I206269);
DFFARX1 I_11965 (I206235,I2859,I206102,I206091,);
nor I_11966 (I206317,I196327,I196339);
nand I_11967 (I206334,I206317,I196333);
nor I_11968 (I206351,I206334,I206218);
nand I_11969 (I206076,I206351,I196315);
DFFARX1 I_11970 (I206334,I2859,I206102,I206088,);
nand I_11971 (I206396,I206218,I196327);
nor I_11972 (I206413,I206218,I196327);
nand I_11973 (I206082,I206201,I206413);
not I_11974 (I206444,I196318);
nor I_11975 (I206461,I206444,I206396);
DFFARX1 I_11976 (I206461,I2859,I206102,I206070,);
nor I_11977 (I206492,I206444,I196312);
and I_11978 (I206509,I206492,I196330);
or I_11979 (I206526,I206509,I196324);
DFFARX1 I_11980 (I206526,I2859,I206102,I206552,);
nor I_11981 (I206560,I206552,I206176);
nor I_11982 (I206079,I206128,I206560);
not I_11983 (I206591,I206552);
nor I_11984 (I206608,I206591,I206286);
DFFARX1 I_11985 (I206608,I2859,I206102,I206085,);
nand I_11986 (I206639,I206591,I206218);
nor I_11987 (I206073,I206444,I206639);
not I_11988 (I206697,I2866);
DFFARX1 I_11989 (I148829,I2859,I206697,I206723,);
DFFARX1 I_11990 (I206723,I2859,I206697,I206740,);
not I_11991 (I206689,I206740);
DFFARX1 I_11992 (I148817,I2859,I206697,I206771,);
not I_11993 (I206779,I148820);
nor I_11994 (I206796,I206723,I206779);
not I_11995 (I206813,I148823);
not I_11996 (I206830,I148835);
nand I_11997 (I206847,I206830,I148823);
nor I_11998 (I206864,I206779,I206847);
nor I_11999 (I206881,I206771,I206864);
DFFARX1 I_12000 (I206830,I2859,I206697,I206686,);
nor I_12001 (I206912,I148835,I148826);
nand I_12002 (I206929,I206912,I148814);
nor I_12003 (I206946,I206929,I206813);
nand I_12004 (I206671,I206946,I148820);
DFFARX1 I_12005 (I206929,I2859,I206697,I206683,);
nand I_12006 (I206991,I206813,I148835);
nor I_12007 (I207008,I206813,I148835);
nand I_12008 (I206677,I206796,I207008);
not I_12009 (I207039,I148832);
nor I_12010 (I207056,I207039,I206991);
DFFARX1 I_12011 (I207056,I2859,I206697,I206665,);
nor I_12012 (I207087,I207039,I148838);
and I_12013 (I207104,I207087,I148841);
or I_12014 (I207121,I207104,I148814);
DFFARX1 I_12015 (I207121,I2859,I206697,I207147,);
nor I_12016 (I207155,I207147,I206771);
nor I_12017 (I206674,I206723,I207155);
not I_12018 (I207186,I207147);
nor I_12019 (I207203,I207186,I206881);
DFFARX1 I_12020 (I207203,I2859,I206697,I206680,);
nand I_12021 (I207234,I207186,I206813);
nor I_12022 (I206668,I207039,I207234);
not I_12023 (I207292,I2866);
DFFARX1 I_12024 (I54872,I2859,I207292,I207318,);
DFFARX1 I_12025 (I207318,I2859,I207292,I207335,);
not I_12026 (I207284,I207335);
DFFARX1 I_12027 (I54896,I2859,I207292,I207366,);
not I_12028 (I207374,I54890);
nor I_12029 (I207391,I207318,I207374);
not I_12030 (I207408,I54884);
not I_12031 (I207425,I54881);
nand I_12032 (I207442,I207425,I54884);
nor I_12033 (I207459,I207374,I207442);
nor I_12034 (I207476,I207366,I207459);
DFFARX1 I_12035 (I207425,I2859,I207292,I207281,);
nor I_12036 (I207507,I54881,I54875);
nand I_12037 (I207524,I207507,I54893);
nor I_12038 (I207541,I207524,I207408);
nand I_12039 (I207266,I207541,I54890);
DFFARX1 I_12040 (I207524,I2859,I207292,I207278,);
nand I_12041 (I207586,I207408,I54881);
nor I_12042 (I207603,I207408,I54881);
nand I_12043 (I207272,I207391,I207603);
not I_12044 (I207634,I54887);
nor I_12045 (I207651,I207634,I207586);
DFFARX1 I_12046 (I207651,I2859,I207292,I207260,);
nor I_12047 (I207682,I207634,I54872);
and I_12048 (I207699,I207682,I54878);
or I_12049 (I207716,I207699,I54875);
DFFARX1 I_12050 (I207716,I2859,I207292,I207742,);
nor I_12051 (I207750,I207742,I207366);
nor I_12052 (I207269,I207318,I207750);
not I_12053 (I207781,I207742);
nor I_12054 (I207798,I207781,I207476);
DFFARX1 I_12055 (I207798,I2859,I207292,I207275,);
nand I_12056 (I207829,I207781,I207408);
nor I_12057 (I207263,I207634,I207829);
not I_12058 (I207887,I2866);
DFFARX1 I_12059 (I104852,I2859,I207887,I207913,);
DFFARX1 I_12060 (I207913,I2859,I207887,I207930,);
not I_12061 (I207879,I207930);
DFFARX1 I_12062 (I104876,I2859,I207887,I207961,);
not I_12063 (I207969,I104870);
nor I_12064 (I207986,I207913,I207969);
not I_12065 (I208003,I104864);
not I_12066 (I208020,I104861);
nand I_12067 (I208037,I208020,I104864);
nor I_12068 (I208054,I207969,I208037);
nor I_12069 (I208071,I207961,I208054);
DFFARX1 I_12070 (I208020,I2859,I207887,I207876,);
nor I_12071 (I208102,I104861,I104855);
nand I_12072 (I208119,I208102,I104873);
nor I_12073 (I208136,I208119,I208003);
nand I_12074 (I207861,I208136,I104870);
DFFARX1 I_12075 (I208119,I2859,I207887,I207873,);
nand I_12076 (I208181,I208003,I104861);
nor I_12077 (I208198,I208003,I104861);
nand I_12078 (I207867,I207986,I208198);
not I_12079 (I208229,I104867);
nor I_12080 (I208246,I208229,I208181);
DFFARX1 I_12081 (I208246,I2859,I207887,I207855,);
nor I_12082 (I208277,I208229,I104852);
and I_12083 (I208294,I208277,I104858);
or I_12084 (I208311,I208294,I104855);
DFFARX1 I_12085 (I208311,I2859,I207887,I208337,);
nor I_12086 (I208345,I208337,I207961);
nor I_12087 (I207864,I207913,I208345);
not I_12088 (I208376,I208337);
nor I_12089 (I208393,I208376,I208071);
DFFARX1 I_12090 (I208393,I2859,I207887,I207870,);
nand I_12091 (I208424,I208376,I208003);
nor I_12092 (I207858,I208229,I208424);
not I_12093 (I208482,I2866);
DFFARX1 I_12094 (I554655,I2859,I208482,I208508,);
DFFARX1 I_12095 (I208508,I2859,I208482,I208525,);
not I_12096 (I208474,I208525);
DFFARX1 I_12097 (I554661,I2859,I208482,I208556,);
not I_12098 (I208564,I554676);
nor I_12099 (I208581,I208508,I208564);
not I_12100 (I208598,I554667);
not I_12101 (I208615,I554664);
nand I_12102 (I208632,I208615,I554667);
nor I_12103 (I208649,I208564,I208632);
nor I_12104 (I208666,I208556,I208649);
DFFARX1 I_12105 (I208615,I2859,I208482,I208471,);
nor I_12106 (I208697,I554664,I554655);
nand I_12107 (I208714,I208697,I554679);
nor I_12108 (I208731,I208714,I208598);
nand I_12109 (I208456,I208731,I554676);
DFFARX1 I_12110 (I208714,I2859,I208482,I208468,);
nand I_12111 (I208776,I208598,I554664);
nor I_12112 (I208793,I208598,I554664);
nand I_12113 (I208462,I208581,I208793);
not I_12114 (I208824,I554673);
nor I_12115 (I208841,I208824,I208776);
DFFARX1 I_12116 (I208841,I2859,I208482,I208450,);
nor I_12117 (I208872,I208824,I554658);
and I_12118 (I208889,I208872,I554670);
or I_12119 (I208906,I208889,I554682);
DFFARX1 I_12120 (I208906,I2859,I208482,I208932,);
nor I_12121 (I208940,I208932,I208556);
nor I_12122 (I208459,I208508,I208940);
not I_12123 (I208971,I208932);
nor I_12124 (I208988,I208971,I208666);
DFFARX1 I_12125 (I208988,I2859,I208482,I208465,);
nand I_12126 (I209019,I208971,I208598);
nor I_12127 (I208453,I208824,I209019);
not I_12128 (I209077,I2866);
DFFARX1 I_12129 (I359181,I2859,I209077,I209103,);
DFFARX1 I_12130 (I209103,I2859,I209077,I209120,);
not I_12131 (I209069,I209120);
DFFARX1 I_12132 (I359178,I2859,I209077,I209151,);
not I_12133 (I209159,I359178);
nor I_12134 (I209176,I209103,I209159);
not I_12135 (I209193,I359175);
not I_12136 (I209210,I359190);
nand I_12137 (I209227,I209210,I359175);
nor I_12138 (I209244,I209159,I209227);
nor I_12139 (I209261,I209151,I209244);
DFFARX1 I_12140 (I209210,I2859,I209077,I209066,);
nor I_12141 (I209292,I359190,I359184);
nand I_12142 (I209309,I209292,I359172);
nor I_12143 (I209326,I209309,I209193);
nand I_12144 (I209051,I209326,I359178);
DFFARX1 I_12145 (I209309,I2859,I209077,I209063,);
nand I_12146 (I209371,I209193,I359190);
nor I_12147 (I209388,I209193,I359190);
nand I_12148 (I209057,I209176,I209388);
not I_12149 (I209419,I359193);
nor I_12150 (I209436,I209419,I209371);
DFFARX1 I_12151 (I209436,I2859,I209077,I209045,);
nor I_12152 (I209467,I209419,I359172);
and I_12153 (I209484,I209467,I359187);
or I_12154 (I209501,I209484,I359175);
DFFARX1 I_12155 (I209501,I2859,I209077,I209527,);
nor I_12156 (I209535,I209527,I209151);
nor I_12157 (I209054,I209103,I209535);
not I_12158 (I209566,I209527);
nor I_12159 (I209583,I209566,I209261);
DFFARX1 I_12160 (I209583,I2859,I209077,I209060,);
nand I_12161 (I209614,I209566,I209193);
nor I_12162 (I209048,I209419,I209614);
not I_12163 (I209672,I2866);
DFFARX1 I_12164 (I242351,I2859,I209672,I209698,);
DFFARX1 I_12165 (I209698,I2859,I209672,I209715,);
not I_12166 (I209664,I209715);
DFFARX1 I_12167 (I242363,I2859,I209672,I209746,);
not I_12168 (I209754,I242348);
nor I_12169 (I209771,I209698,I209754);
not I_12170 (I209788,I242366);
not I_12171 (I209805,I242357);
nand I_12172 (I209822,I209805,I242366);
nor I_12173 (I209839,I209754,I209822);
nor I_12174 (I209856,I209746,I209839);
DFFARX1 I_12175 (I209805,I2859,I209672,I209661,);
nor I_12176 (I209887,I242357,I242369);
nand I_12177 (I209904,I209887,I242372);
nor I_12178 (I209921,I209904,I209788);
nand I_12179 (I209646,I209921,I242348);
DFFARX1 I_12180 (I209904,I2859,I209672,I209658,);
nand I_12181 (I209966,I209788,I242357);
nor I_12182 (I209983,I209788,I242357);
nand I_12183 (I209652,I209771,I209983);
not I_12184 (I210014,I242348);
nor I_12185 (I210031,I210014,I209966);
DFFARX1 I_12186 (I210031,I2859,I209672,I209640,);
nor I_12187 (I210062,I210014,I242360);
and I_12188 (I210079,I210062,I242354);
or I_12189 (I210096,I210079,I242351);
DFFARX1 I_12190 (I210096,I2859,I209672,I210122,);
nor I_12191 (I210130,I210122,I209746);
nor I_12192 (I209649,I209698,I210130);
not I_12193 (I210161,I210122);
nor I_12194 (I210178,I210161,I209856);
DFFARX1 I_12195 (I210178,I2859,I209672,I209655,);
nand I_12196 (I210209,I210161,I209788);
nor I_12197 (I209643,I210014,I210209);
not I_12198 (I210267,I2866);
DFFARX1 I_12199 (I78077,I2859,I210267,I210293,);
DFFARX1 I_12200 (I210293,I2859,I210267,I210310,);
not I_12201 (I210259,I210310);
DFFARX1 I_12202 (I78101,I2859,I210267,I210341,);
not I_12203 (I210349,I78095);
nor I_12204 (I210366,I210293,I210349);
not I_12205 (I210383,I78089);
not I_12206 (I210400,I78086);
nand I_12207 (I210417,I210400,I78089);
nor I_12208 (I210434,I210349,I210417);
nor I_12209 (I210451,I210341,I210434);
DFFARX1 I_12210 (I210400,I2859,I210267,I210256,);
nor I_12211 (I210482,I78086,I78080);
nand I_12212 (I210499,I210482,I78098);
nor I_12213 (I210516,I210499,I210383);
nand I_12214 (I210241,I210516,I78095);
DFFARX1 I_12215 (I210499,I2859,I210267,I210253,);
nand I_12216 (I210561,I210383,I78086);
nor I_12217 (I210578,I210383,I78086);
nand I_12218 (I210247,I210366,I210578);
not I_12219 (I210609,I78092);
nor I_12220 (I210626,I210609,I210561);
DFFARX1 I_12221 (I210626,I2859,I210267,I210235,);
nor I_12222 (I210657,I210609,I78077);
and I_12223 (I210674,I210657,I78083);
or I_12224 (I210691,I210674,I78080);
DFFARX1 I_12225 (I210691,I2859,I210267,I210717,);
nor I_12226 (I210725,I210717,I210341);
nor I_12227 (I210244,I210293,I210725);
not I_12228 (I210756,I210717);
nor I_12229 (I210773,I210756,I210451);
DFFARX1 I_12230 (I210773,I2859,I210267,I210250,);
nand I_12231 (I210804,I210756,I210383);
nor I_12232 (I210238,I210609,I210804);
not I_12233 (I210862,I2866);
DFFARX1 I_12234 (I469554,I2859,I210862,I210888,);
DFFARX1 I_12235 (I210888,I2859,I210862,I210905,);
not I_12236 (I210854,I210905);
DFFARX1 I_12237 (I469536,I2859,I210862,I210936,);
not I_12238 (I210944,I469542);
nor I_12239 (I210961,I210888,I210944);
not I_12240 (I210978,I469557);
not I_12241 (I210995,I469548);
nand I_12242 (I211012,I210995,I469557);
nor I_12243 (I211029,I210944,I211012);
nor I_12244 (I211046,I210936,I211029);
DFFARX1 I_12245 (I210995,I2859,I210862,I210851,);
nor I_12246 (I211077,I469548,I469560);
nand I_12247 (I211094,I211077,I469539);
nor I_12248 (I211111,I211094,I210978);
nand I_12249 (I210836,I211111,I469542);
DFFARX1 I_12250 (I211094,I2859,I210862,I210848,);
nand I_12251 (I211156,I210978,I469548);
nor I_12252 (I211173,I210978,I469548);
nand I_12253 (I210842,I210961,I211173);
not I_12254 (I211204,I469545);
nor I_12255 (I211221,I211204,I211156);
DFFARX1 I_12256 (I211221,I2859,I210862,I210830,);
nor I_12257 (I211252,I211204,I469551);
and I_12258 (I211269,I211252,I469536);
or I_12259 (I211286,I211269,I469539);
DFFARX1 I_12260 (I211286,I2859,I210862,I211312,);
nor I_12261 (I211320,I211312,I210936);
nor I_12262 (I210839,I210888,I211320);
not I_12263 (I211351,I211312);
nor I_12264 (I211368,I211351,I211046);
DFFARX1 I_12265 (I211368,I2859,I210862,I210845,);
nand I_12266 (I211399,I211351,I210978);
nor I_12267 (I210833,I211204,I211399);
not I_12268 (I211457,I2866);
DFFARX1 I_12269 (I479958,I2859,I211457,I211483,);
DFFARX1 I_12270 (I211483,I2859,I211457,I211500,);
not I_12271 (I211449,I211500);
DFFARX1 I_12272 (I479940,I2859,I211457,I211531,);
not I_12273 (I211539,I479946);
nor I_12274 (I211556,I211483,I211539);
not I_12275 (I211573,I479961);
not I_12276 (I211590,I479952);
nand I_12277 (I211607,I211590,I479961);
nor I_12278 (I211624,I211539,I211607);
nor I_12279 (I211641,I211531,I211624);
DFFARX1 I_12280 (I211590,I2859,I211457,I211446,);
nor I_12281 (I211672,I479952,I479964);
nand I_12282 (I211689,I211672,I479943);
nor I_12283 (I211706,I211689,I211573);
nand I_12284 (I211431,I211706,I479946);
DFFARX1 I_12285 (I211689,I2859,I211457,I211443,);
nand I_12286 (I211751,I211573,I479952);
nor I_12287 (I211768,I211573,I479952);
nand I_12288 (I211437,I211556,I211768);
not I_12289 (I211799,I479949);
nor I_12290 (I211816,I211799,I211751);
DFFARX1 I_12291 (I211816,I2859,I211457,I211425,);
nor I_12292 (I211847,I211799,I479955);
and I_12293 (I211864,I211847,I479940);
or I_12294 (I211881,I211864,I479943);
DFFARX1 I_12295 (I211881,I2859,I211457,I211907,);
nor I_12296 (I211915,I211907,I211531);
nor I_12297 (I211434,I211483,I211915);
not I_12298 (I211946,I211907);
nor I_12299 (I211963,I211946,I211641);
DFFARX1 I_12300 (I211963,I2859,I211457,I211440,);
nand I_12301 (I211994,I211946,I211573);
nor I_12302 (I211428,I211799,I211994);
not I_12303 (I212052,I2866);
DFFARX1 I_12304 (I267789,I2859,I212052,I212078,);
DFFARX1 I_12305 (I212078,I2859,I212052,I212095,);
not I_12306 (I212044,I212095);
DFFARX1 I_12307 (I267783,I2859,I212052,I212126,);
not I_12308 (I212134,I267780);
nor I_12309 (I212151,I212078,I212134);
not I_12310 (I212168,I267792);
not I_12311 (I212185,I267795);
nand I_12312 (I212202,I212185,I267792);
nor I_12313 (I212219,I212134,I212202);
nor I_12314 (I212236,I212126,I212219);
DFFARX1 I_12315 (I212185,I2859,I212052,I212041,);
nor I_12316 (I212267,I267795,I267804);
nand I_12317 (I212284,I212267,I267798);
nor I_12318 (I212301,I212284,I212168);
nand I_12319 (I212026,I212301,I267780);
DFFARX1 I_12320 (I212284,I2859,I212052,I212038,);
nand I_12321 (I212346,I212168,I267795);
nor I_12322 (I212363,I212168,I267795);
nand I_12323 (I212032,I212151,I212363);
not I_12324 (I212394,I267786);
nor I_12325 (I212411,I212394,I212346);
DFFARX1 I_12326 (I212411,I2859,I212052,I212020,);
nor I_12327 (I212442,I212394,I267801);
and I_12328 (I212459,I212442,I267780);
or I_12329 (I212476,I212459,I267783);
DFFARX1 I_12330 (I212476,I2859,I212052,I212502,);
nor I_12331 (I212510,I212502,I212126);
nor I_12332 (I212029,I212078,I212510);
not I_12333 (I212541,I212502);
nor I_12334 (I212558,I212541,I212236);
DFFARX1 I_12335 (I212558,I2859,I212052,I212035,);
nand I_12336 (I212589,I212541,I212168);
nor I_12337 (I212023,I212394,I212589);
not I_12338 (I212647,I2866);
DFFARX1 I_12339 (I97712,I2859,I212647,I212673,);
DFFARX1 I_12340 (I212673,I2859,I212647,I212690,);
not I_12341 (I212639,I212690);
DFFARX1 I_12342 (I97736,I2859,I212647,I212721,);
not I_12343 (I212729,I97730);
nor I_12344 (I212746,I212673,I212729);
not I_12345 (I212763,I97724);
not I_12346 (I212780,I97721);
nand I_12347 (I212797,I212780,I97724);
nor I_12348 (I212814,I212729,I212797);
nor I_12349 (I212831,I212721,I212814);
DFFARX1 I_12350 (I212780,I2859,I212647,I212636,);
nor I_12351 (I212862,I97721,I97715);
nand I_12352 (I212879,I212862,I97733);
nor I_12353 (I212896,I212879,I212763);
nand I_12354 (I212621,I212896,I97730);
DFFARX1 I_12355 (I212879,I2859,I212647,I212633,);
nand I_12356 (I212941,I212763,I97721);
nor I_12357 (I212958,I212763,I97721);
nand I_12358 (I212627,I212746,I212958);
not I_12359 (I212989,I97727);
nor I_12360 (I213006,I212989,I212941);
DFFARX1 I_12361 (I213006,I2859,I212647,I212615,);
nor I_12362 (I213037,I212989,I97712);
and I_12363 (I213054,I213037,I97718);
or I_12364 (I213071,I213054,I97715);
DFFARX1 I_12365 (I213071,I2859,I212647,I213097,);
nor I_12366 (I213105,I213097,I212721);
nor I_12367 (I212624,I212673,I213105);
not I_12368 (I213136,I213097);
nor I_12369 (I213153,I213136,I212831);
DFFARX1 I_12370 (I213153,I2859,I212647,I212630,);
nand I_12371 (I213184,I213136,I212763);
nor I_12372 (I212618,I212989,I213184);
not I_12373 (I213242,I2866);
DFFARX1 I_12374 (I351276,I2859,I213242,I213268,);
DFFARX1 I_12375 (I213268,I2859,I213242,I213285,);
not I_12376 (I213234,I213285);
DFFARX1 I_12377 (I351273,I2859,I213242,I213316,);
not I_12378 (I213324,I351273);
nor I_12379 (I213341,I213268,I213324);
not I_12380 (I213358,I351270);
not I_12381 (I213375,I351285);
nand I_12382 (I213392,I213375,I351270);
nor I_12383 (I213409,I213324,I213392);
nor I_12384 (I213426,I213316,I213409);
DFFARX1 I_12385 (I213375,I2859,I213242,I213231,);
nor I_12386 (I213457,I351285,I351279);
nand I_12387 (I213474,I213457,I351267);
nor I_12388 (I213491,I213474,I213358);
nand I_12389 (I213216,I213491,I351273);
DFFARX1 I_12390 (I213474,I2859,I213242,I213228,);
nand I_12391 (I213536,I213358,I351285);
nor I_12392 (I213553,I213358,I351285);
nand I_12393 (I213222,I213341,I213553);
not I_12394 (I213584,I351288);
nor I_12395 (I213601,I213584,I213536);
DFFARX1 I_12396 (I213601,I2859,I213242,I213210,);
nor I_12397 (I213632,I213584,I351267);
and I_12398 (I213649,I213632,I351282);
or I_12399 (I213666,I213649,I351270);
DFFARX1 I_12400 (I213666,I2859,I213242,I213692,);
nor I_12401 (I213700,I213692,I213316);
nor I_12402 (I213219,I213268,I213700);
not I_12403 (I213731,I213692);
nor I_12404 (I213748,I213731,I213426);
DFFARX1 I_12405 (I213748,I2859,I213242,I213225,);
nand I_12406 (I213779,I213731,I213358);
nor I_12407 (I213213,I213584,I213779);
not I_12408 (I213837,I2866);
DFFARX1 I_12409 (I420950,I2859,I213837,I213863,);
DFFARX1 I_12410 (I213863,I2859,I213837,I213880,);
not I_12411 (I213829,I213880);
DFFARX1 I_12412 (I420953,I2859,I213837,I213911,);
not I_12413 (I213919,I420956);
nor I_12414 (I213936,I213863,I213919);
not I_12415 (I213953,I420968);
not I_12416 (I213970,I420959);
nand I_12417 (I213987,I213970,I420968);
nor I_12418 (I214004,I213919,I213987);
nor I_12419 (I214021,I213911,I214004);
DFFARX1 I_12420 (I213970,I2859,I213837,I213826,);
nor I_12421 (I214052,I420959,I420965);
nand I_12422 (I214069,I214052,I420953);
nor I_12423 (I214086,I214069,I213953);
nand I_12424 (I213811,I214086,I420956);
DFFARX1 I_12425 (I214069,I2859,I213837,I213823,);
nand I_12426 (I214131,I213953,I420959);
nor I_12427 (I214148,I213953,I420959);
nand I_12428 (I213817,I213936,I214148);
not I_12429 (I214179,I420956);
nor I_12430 (I214196,I214179,I214131);
DFFARX1 I_12431 (I214196,I2859,I213837,I213805,);
nor I_12432 (I214227,I214179,I420962);
and I_12433 (I214244,I214227,I420950);
or I_12434 (I214261,I214244,I420971);
DFFARX1 I_12435 (I214261,I2859,I213837,I214287,);
nor I_12436 (I214295,I214287,I213911);
nor I_12437 (I213814,I213863,I214295);
not I_12438 (I214326,I214287);
nor I_12439 (I214343,I214326,I214021);
DFFARX1 I_12440 (I214343,I2859,I213837,I213820,);
nand I_12441 (I214374,I214326,I213953);
nor I_12442 (I213808,I214179,I214374);
not I_12443 (I214432,I2866);
DFFARX1 I_12444 (I514994,I2859,I214432,I214458,);
DFFARX1 I_12445 (I214458,I2859,I214432,I214475,);
not I_12446 (I214424,I214475);
DFFARX1 I_12447 (I515009,I2859,I214432,I214506,);
not I_12448 (I214514,I515018);
nor I_12449 (I214531,I214458,I214514);
not I_12450 (I214548,I514997);
not I_12451 (I214565,I515003);
nand I_12452 (I214582,I214565,I514997);
nor I_12453 (I214599,I214514,I214582);
nor I_12454 (I214616,I214506,I214599);
DFFARX1 I_12455 (I214565,I2859,I214432,I214421,);
nor I_12456 (I214647,I515003,I515015);
nand I_12457 (I214664,I214647,I515012);
nor I_12458 (I214681,I214664,I214548);
nand I_12459 (I214406,I214681,I515018);
DFFARX1 I_12460 (I214664,I2859,I214432,I214418,);
nand I_12461 (I214726,I214548,I515003);
nor I_12462 (I214743,I214548,I515003);
nand I_12463 (I214412,I214531,I214743);
not I_12464 (I214774,I514994);
nor I_12465 (I214791,I214774,I214726);
DFFARX1 I_12466 (I214791,I2859,I214432,I214400,);
nor I_12467 (I214822,I214774,I515006);
and I_12468 (I214839,I214822,I515000);
or I_12469 (I214856,I214839,I514997);
DFFARX1 I_12470 (I214856,I2859,I214432,I214882,);
nor I_12471 (I214890,I214882,I214506);
nor I_12472 (I214409,I214458,I214890);
not I_12473 (I214921,I214882);
nor I_12474 (I214938,I214921,I214616);
DFFARX1 I_12475 (I214938,I2859,I214432,I214415,);
nand I_12476 (I214969,I214921,I214548);
nor I_12477 (I214403,I214774,I214969);
not I_12478 (I215027,I2866);
DFFARX1 I_12479 (I536805,I2859,I215027,I215053,);
DFFARX1 I_12480 (I215053,I2859,I215027,I215070,);
not I_12481 (I215019,I215070);
DFFARX1 I_12482 (I536811,I2859,I215027,I215101,);
not I_12483 (I215109,I536826);
nor I_12484 (I215126,I215053,I215109);
not I_12485 (I215143,I536817);
not I_12486 (I215160,I536814);
nand I_12487 (I215177,I215160,I536817);
nor I_12488 (I215194,I215109,I215177);
nor I_12489 (I215211,I215101,I215194);
DFFARX1 I_12490 (I215160,I2859,I215027,I215016,);
nor I_12491 (I215242,I536814,I536805);
nand I_12492 (I215259,I215242,I536829);
nor I_12493 (I215276,I215259,I215143);
nand I_12494 (I215001,I215276,I536826);
DFFARX1 I_12495 (I215259,I2859,I215027,I215013,);
nand I_12496 (I215321,I215143,I536814);
nor I_12497 (I215338,I215143,I536814);
nand I_12498 (I215007,I215126,I215338);
not I_12499 (I215369,I536823);
nor I_12500 (I215386,I215369,I215321);
DFFARX1 I_12501 (I215386,I2859,I215027,I214995,);
nor I_12502 (I215417,I215369,I536808);
and I_12503 (I215434,I215417,I536820);
or I_12504 (I215451,I215434,I536832);
DFFARX1 I_12505 (I215451,I2859,I215027,I215477,);
nor I_12506 (I215485,I215477,I215101);
nor I_12507 (I215004,I215053,I215485);
not I_12508 (I215516,I215477);
nor I_12509 (I215533,I215516,I215211);
DFFARX1 I_12510 (I215533,I2859,I215027,I215010,);
nand I_12511 (I215564,I215516,I215143);
nor I_12512 (I214998,I215369,I215564);
not I_12513 (I215622,I2866);
DFFARX1 I_12514 (I99497,I2859,I215622,I215648,);
DFFARX1 I_12515 (I215648,I2859,I215622,I215665,);
not I_12516 (I215614,I215665);
DFFARX1 I_12517 (I99521,I2859,I215622,I215696,);
not I_12518 (I215704,I99515);
nor I_12519 (I215721,I215648,I215704);
not I_12520 (I215738,I99509);
not I_12521 (I215755,I99506);
nand I_12522 (I215772,I215755,I99509);
nor I_12523 (I215789,I215704,I215772);
nor I_12524 (I215806,I215696,I215789);
DFFARX1 I_12525 (I215755,I2859,I215622,I215611,);
nor I_12526 (I215837,I99506,I99500);
nand I_12527 (I215854,I215837,I99518);
nor I_12528 (I215871,I215854,I215738);
nand I_12529 (I215596,I215871,I99515);
DFFARX1 I_12530 (I215854,I2859,I215622,I215608,);
nand I_12531 (I215916,I215738,I99506);
nor I_12532 (I215933,I215738,I99506);
nand I_12533 (I215602,I215721,I215933);
not I_12534 (I215964,I99512);
nor I_12535 (I215981,I215964,I215916);
DFFARX1 I_12536 (I215981,I2859,I215622,I215590,);
nor I_12537 (I216012,I215964,I99497);
and I_12538 (I216029,I216012,I99503);
or I_12539 (I216046,I216029,I99500);
DFFARX1 I_12540 (I216046,I2859,I215622,I216072,);
nor I_12541 (I216080,I216072,I215696);
nor I_12542 (I215599,I215648,I216080);
not I_12543 (I216111,I216072);
nor I_12544 (I216128,I216111,I215806);
DFFARX1 I_12545 (I216128,I2859,I215622,I215605,);
nand I_12546 (I216159,I216111,I215738);
nor I_12547 (I215593,I215964,I216159);
not I_12548 (I216217,I2866);
DFFARX1 I_12549 (I468398,I2859,I216217,I216243,);
DFFARX1 I_12550 (I216243,I2859,I216217,I216260,);
not I_12551 (I216209,I216260);
DFFARX1 I_12552 (I468380,I2859,I216217,I216291,);
not I_12553 (I216299,I468386);
nor I_12554 (I216316,I216243,I216299);
not I_12555 (I216333,I468401);
not I_12556 (I216350,I468392);
nand I_12557 (I216367,I216350,I468401);
nor I_12558 (I216384,I216299,I216367);
nor I_12559 (I216401,I216291,I216384);
DFFARX1 I_12560 (I216350,I2859,I216217,I216206,);
nor I_12561 (I216432,I468392,I468404);
nand I_12562 (I216449,I216432,I468383);
nor I_12563 (I216466,I216449,I216333);
nand I_12564 (I216191,I216466,I468386);
DFFARX1 I_12565 (I216449,I2859,I216217,I216203,);
nand I_12566 (I216511,I216333,I468392);
nor I_12567 (I216528,I216333,I468392);
nand I_12568 (I216197,I216316,I216528);
not I_12569 (I216559,I468389);
nor I_12570 (I216576,I216559,I216511);
DFFARX1 I_12571 (I216576,I2859,I216217,I216185,);
nor I_12572 (I216607,I216559,I468395);
and I_12573 (I216624,I216607,I468380);
or I_12574 (I216641,I216624,I468383);
DFFARX1 I_12575 (I216641,I2859,I216217,I216667,);
nor I_12576 (I216675,I216667,I216291);
nor I_12577 (I216194,I216243,I216675);
not I_12578 (I216706,I216667);
nor I_12579 (I216723,I216706,I216401);
DFFARX1 I_12580 (I216723,I2859,I216217,I216200,);
nand I_12581 (I216754,I216706,I216333);
nor I_12582 (I216188,I216559,I216754);
not I_12583 (I216812,I2866);
DFFARX1 I_12584 (I322818,I2859,I216812,I216838,);
DFFARX1 I_12585 (I216838,I2859,I216812,I216855,);
not I_12586 (I216804,I216855);
DFFARX1 I_12587 (I322815,I2859,I216812,I216886,);
not I_12588 (I216894,I322815);
nor I_12589 (I216911,I216838,I216894);
not I_12590 (I216928,I322812);
not I_12591 (I216945,I322827);
nand I_12592 (I216962,I216945,I322812);
nor I_12593 (I216979,I216894,I216962);
nor I_12594 (I216996,I216886,I216979);
DFFARX1 I_12595 (I216945,I2859,I216812,I216801,);
nor I_12596 (I217027,I322827,I322821);
nand I_12597 (I217044,I217027,I322809);
nor I_12598 (I217061,I217044,I216928);
nand I_12599 (I216786,I217061,I322815);
DFFARX1 I_12600 (I217044,I2859,I216812,I216798,);
nand I_12601 (I217106,I216928,I322827);
nor I_12602 (I217123,I216928,I322827);
nand I_12603 (I216792,I216911,I217123);
not I_12604 (I217154,I322830);
nor I_12605 (I217171,I217154,I217106);
DFFARX1 I_12606 (I217171,I2859,I216812,I216780,);
nor I_12607 (I217202,I217154,I322809);
and I_12608 (I217219,I217202,I322824);
or I_12609 (I217236,I217219,I322812);
DFFARX1 I_12610 (I217236,I2859,I216812,I217262,);
nor I_12611 (I217270,I217262,I216886);
nor I_12612 (I216789,I216838,I217270);
not I_12613 (I217301,I217262);
nor I_12614 (I217318,I217301,I216996);
DFFARX1 I_12615 (I217318,I2859,I216812,I216795,);
nand I_12616 (I217349,I217301,I216928);
nor I_12617 (I216783,I217154,I217349);
not I_12618 (I217407,I2866);
DFFARX1 I_12619 (I175640,I2859,I217407,I217433,);
DFFARX1 I_12620 (I217433,I2859,I217407,I217450,);
not I_12621 (I217399,I217450);
DFFARX1 I_12622 (I175664,I2859,I217407,I217481,);
not I_12623 (I217489,I175643);
nor I_12624 (I217506,I217433,I217489);
not I_12625 (I217523,I175649);
not I_12626 (I217540,I175655);
nand I_12627 (I217557,I217540,I175649);
nor I_12628 (I217574,I217489,I217557);
nor I_12629 (I217591,I217481,I217574);
DFFARX1 I_12630 (I217540,I2859,I217407,I217396,);
nor I_12631 (I217622,I175655,I175667);
nand I_12632 (I217639,I217622,I175661);
nor I_12633 (I217656,I217639,I217523);
nand I_12634 (I217381,I217656,I175643);
DFFARX1 I_12635 (I217639,I2859,I217407,I217393,);
nand I_12636 (I217701,I217523,I175655);
nor I_12637 (I217718,I217523,I175655);
nand I_12638 (I217387,I217506,I217718);
not I_12639 (I217749,I175646);
nor I_12640 (I217766,I217749,I217701);
DFFARX1 I_12641 (I217766,I2859,I217407,I217375,);
nor I_12642 (I217797,I217749,I175640);
and I_12643 (I217814,I217797,I175658);
or I_12644 (I217831,I217814,I175652);
DFFARX1 I_12645 (I217831,I2859,I217407,I217857,);
nor I_12646 (I217865,I217857,I217481);
nor I_12647 (I217384,I217433,I217865);
not I_12648 (I217896,I217857);
nor I_12649 (I217913,I217896,I217591);
DFFARX1 I_12650 (I217913,I2859,I217407,I217390,);
nand I_12651 (I217944,I217896,I217523);
nor I_12652 (I217378,I217749,I217944);
not I_12653 (I218002,I2866);
DFFARX1 I_12654 (I132492,I2859,I218002,I218028,);
DFFARX1 I_12655 (I218028,I2859,I218002,I218045,);
not I_12656 (I217994,I218045);
DFFARX1 I_12657 (I132480,I2859,I218002,I218076,);
not I_12658 (I218084,I132483);
nor I_12659 (I218101,I218028,I218084);
not I_12660 (I218118,I132486);
not I_12661 (I218135,I132498);
nand I_12662 (I218152,I218135,I132486);
nor I_12663 (I218169,I218084,I218152);
nor I_12664 (I218186,I218076,I218169);
DFFARX1 I_12665 (I218135,I2859,I218002,I217991,);
nor I_12666 (I218217,I132498,I132489);
nand I_12667 (I218234,I218217,I132477);
nor I_12668 (I218251,I218234,I218118);
nand I_12669 (I217976,I218251,I132483);
DFFARX1 I_12670 (I218234,I2859,I218002,I217988,);
nand I_12671 (I218296,I218118,I132498);
nor I_12672 (I218313,I218118,I132498);
nand I_12673 (I217982,I218101,I218313);
not I_12674 (I218344,I132495);
nor I_12675 (I218361,I218344,I218296);
DFFARX1 I_12676 (I218361,I2859,I218002,I217970,);
nor I_12677 (I218392,I218344,I132501);
and I_12678 (I218409,I218392,I132504);
or I_12679 (I218426,I218409,I132477);
DFFARX1 I_12680 (I218426,I2859,I218002,I218452,);
nor I_12681 (I218460,I218452,I218076);
nor I_12682 (I217979,I218028,I218460);
not I_12683 (I218491,I218452);
nor I_12684 (I218508,I218491,I218186);
DFFARX1 I_12685 (I218508,I2859,I218002,I217985,);
nand I_12686 (I218539,I218491,I218118);
nor I_12687 (I217973,I218344,I218539);
not I_12688 (I218597,I2866);
DFFARX1 I_12689 (I434414,I2859,I218597,I218623,);
DFFARX1 I_12690 (I218623,I2859,I218597,I218640,);
not I_12691 (I218589,I218640);
DFFARX1 I_12692 (I434417,I2859,I218597,I218671,);
not I_12693 (I218679,I434420);
nor I_12694 (I218696,I218623,I218679);
not I_12695 (I218713,I434432);
not I_12696 (I218730,I434423);
nand I_12697 (I218747,I218730,I434432);
nor I_12698 (I218764,I218679,I218747);
nor I_12699 (I218781,I218671,I218764);
DFFARX1 I_12700 (I218730,I2859,I218597,I218586,);
nor I_12701 (I218812,I434423,I434429);
nand I_12702 (I218829,I218812,I434417);
nor I_12703 (I218846,I218829,I218713);
nand I_12704 (I218571,I218846,I434420);
DFFARX1 I_12705 (I218829,I2859,I218597,I218583,);
nand I_12706 (I218891,I218713,I434423);
nor I_12707 (I218908,I218713,I434423);
nand I_12708 (I218577,I218696,I218908);
not I_12709 (I218939,I434420);
nor I_12710 (I218956,I218939,I218891);
DFFARX1 I_12711 (I218956,I2859,I218597,I218565,);
nor I_12712 (I218987,I218939,I434426);
and I_12713 (I219004,I218987,I434414);
or I_12714 (I219021,I219004,I434435);
DFFARX1 I_12715 (I219021,I2859,I218597,I219047,);
nor I_12716 (I219055,I219047,I218671);
nor I_12717 (I218574,I218623,I219055);
not I_12718 (I219086,I219047);
nor I_12719 (I219103,I219086,I218781);
DFFARX1 I_12720 (I219103,I2859,I218597,I218580,);
nand I_12721 (I219134,I219086,I218713);
nor I_12722 (I218568,I218939,I219134);
not I_12723 (I219192,I2866);
DFFARX1 I_12724 (I354438,I2859,I219192,I219218,);
DFFARX1 I_12725 (I219218,I2859,I219192,I219235,);
not I_12726 (I219184,I219235);
DFFARX1 I_12727 (I354435,I2859,I219192,I219266,);
not I_12728 (I219274,I354435);
nor I_12729 (I219291,I219218,I219274);
not I_12730 (I219308,I354432);
not I_12731 (I219325,I354447);
nand I_12732 (I219342,I219325,I354432);
nor I_12733 (I219359,I219274,I219342);
nor I_12734 (I219376,I219266,I219359);
DFFARX1 I_12735 (I219325,I2859,I219192,I219181,);
nor I_12736 (I219407,I354447,I354441);
nand I_12737 (I219424,I219407,I354429);
nor I_12738 (I219441,I219424,I219308);
nand I_12739 (I219166,I219441,I354435);
DFFARX1 I_12740 (I219424,I2859,I219192,I219178,);
nand I_12741 (I219486,I219308,I354447);
nor I_12742 (I219503,I219308,I354447);
nand I_12743 (I219172,I219291,I219503);
not I_12744 (I219534,I354450);
nor I_12745 (I219551,I219534,I219486);
DFFARX1 I_12746 (I219551,I2859,I219192,I219160,);
nor I_12747 (I219582,I219534,I354429);
and I_12748 (I219599,I219582,I354444);
or I_12749 (I219616,I219599,I354432);
DFFARX1 I_12750 (I219616,I2859,I219192,I219642,);
nor I_12751 (I219650,I219642,I219266);
nor I_12752 (I219169,I219218,I219650);
not I_12753 (I219681,I219642);
nor I_12754 (I219698,I219681,I219376);
DFFARX1 I_12755 (I219698,I2859,I219192,I219175,);
nand I_12756 (I219729,I219681,I219308);
nor I_12757 (I219163,I219534,I219729);
not I_12758 (I219787,I2866);
DFFARX1 I_12759 (I568340,I2859,I219787,I219813,);
DFFARX1 I_12760 (I219813,I2859,I219787,I219830,);
not I_12761 (I219779,I219830);
DFFARX1 I_12762 (I568346,I2859,I219787,I219861,);
not I_12763 (I219869,I568361);
nor I_12764 (I219886,I219813,I219869);
not I_12765 (I219903,I568352);
not I_12766 (I219920,I568349);
nand I_12767 (I219937,I219920,I568352);
nor I_12768 (I219954,I219869,I219937);
nor I_12769 (I219971,I219861,I219954);
DFFARX1 I_12770 (I219920,I2859,I219787,I219776,);
nor I_12771 (I220002,I568349,I568340);
nand I_12772 (I220019,I220002,I568364);
nor I_12773 (I220036,I220019,I219903);
nand I_12774 (I219761,I220036,I568361);
DFFARX1 I_12775 (I220019,I2859,I219787,I219773,);
nand I_12776 (I220081,I219903,I568349);
nor I_12777 (I220098,I219903,I568349);
nand I_12778 (I219767,I219886,I220098);
not I_12779 (I220129,I568358);
nor I_12780 (I220146,I220129,I220081);
DFFARX1 I_12781 (I220146,I2859,I219787,I219755,);
nor I_12782 (I220177,I220129,I568343);
and I_12783 (I220194,I220177,I568355);
or I_12784 (I220211,I220194,I568367);
DFFARX1 I_12785 (I220211,I2859,I219787,I220237,);
nor I_12786 (I220245,I220237,I219861);
nor I_12787 (I219764,I219813,I220245);
not I_12788 (I220276,I220237);
nor I_12789 (I220293,I220276,I219971);
DFFARX1 I_12790 (I220293,I2859,I219787,I219770,);
nand I_12791 (I220324,I220276,I219903);
nor I_12792 (I219758,I220129,I220324);
not I_12793 (I220382,I2866);
DFFARX1 I_12794 (I470710,I2859,I220382,I220408,);
DFFARX1 I_12795 (I220408,I2859,I220382,I220425,);
not I_12796 (I220374,I220425);
DFFARX1 I_12797 (I470692,I2859,I220382,I220456,);
not I_12798 (I220464,I470698);
nor I_12799 (I220481,I220408,I220464);
not I_12800 (I220498,I470713);
not I_12801 (I220515,I470704);
nand I_12802 (I220532,I220515,I470713);
nor I_12803 (I220549,I220464,I220532);
nor I_12804 (I220566,I220456,I220549);
DFFARX1 I_12805 (I220515,I2859,I220382,I220371,);
nor I_12806 (I220597,I470704,I470716);
nand I_12807 (I220614,I220597,I470695);
nor I_12808 (I220631,I220614,I220498);
nand I_12809 (I220356,I220631,I470698);
DFFARX1 I_12810 (I220614,I2859,I220382,I220368,);
nand I_12811 (I220676,I220498,I470704);
nor I_12812 (I220693,I220498,I470704);
nand I_12813 (I220362,I220481,I220693);
not I_12814 (I220724,I470701);
nor I_12815 (I220741,I220724,I220676);
DFFARX1 I_12816 (I220741,I2859,I220382,I220350,);
nor I_12817 (I220772,I220724,I470707);
and I_12818 (I220789,I220772,I470692);
or I_12819 (I220806,I220789,I470695);
DFFARX1 I_12820 (I220806,I2859,I220382,I220832,);
nor I_12821 (I220840,I220832,I220456);
nor I_12822 (I220359,I220408,I220840);
not I_12823 (I220871,I220832);
nor I_12824 (I220888,I220871,I220566);
DFFARX1 I_12825 (I220888,I2859,I220382,I220365,);
nand I_12826 (I220919,I220871,I220498);
nor I_12827 (I220353,I220724,I220919);
not I_12828 (I220977,I2866);
DFFARX1 I_12829 (I199032,I2859,I220977,I221003,);
DFFARX1 I_12830 (I221003,I2859,I220977,I221020,);
not I_12831 (I220969,I221020);
DFFARX1 I_12832 (I199056,I2859,I220977,I221051,);
not I_12833 (I221059,I199035);
nor I_12834 (I221076,I221003,I221059);
not I_12835 (I221093,I199041);
not I_12836 (I221110,I199047);
nand I_12837 (I221127,I221110,I199041);
nor I_12838 (I221144,I221059,I221127);
nor I_12839 (I221161,I221051,I221144);
DFFARX1 I_12840 (I221110,I2859,I220977,I220966,);
nor I_12841 (I221192,I199047,I199059);
nand I_12842 (I221209,I221192,I199053);
nor I_12843 (I221226,I221209,I221093);
nand I_12844 (I220951,I221226,I199035);
DFFARX1 I_12845 (I221209,I2859,I220977,I220963,);
nand I_12846 (I221271,I221093,I199047);
nor I_12847 (I221288,I221093,I199047);
nand I_12848 (I220957,I221076,I221288);
not I_12849 (I221319,I199038);
nor I_12850 (I221336,I221319,I221271);
DFFARX1 I_12851 (I221336,I2859,I220977,I220945,);
nor I_12852 (I221367,I221319,I199032);
and I_12853 (I221384,I221367,I199050);
or I_12854 (I221401,I221384,I199044);
DFFARX1 I_12855 (I221401,I2859,I220977,I221427,);
nor I_12856 (I221435,I221427,I221051);
nor I_12857 (I220954,I221003,I221435);
not I_12858 (I221466,I221427);
nor I_12859 (I221483,I221466,I221161);
DFFARX1 I_12860 (I221483,I2859,I220977,I220960,);
nand I_12861 (I221514,I221466,I221093);
nor I_12862 (I220948,I221319,I221514);
not I_12863 (I221572,I2866);
DFFARX1 I_12864 (I276450,I2859,I221572,I221598,);
not I_12865 (I221606,I221598);
DFFARX1 I_12866 (I276462,I2859,I221572,I221632,);
not I_12867 (I221640,I276453);
nand I_12868 (I221657,I221640,I276456);
not I_12869 (I221674,I221657);
nor I_12870 (I221691,I221674,I276459);
nor I_12871 (I221708,I221606,I221691);
DFFARX1 I_12872 (I221708,I2859,I221572,I221558,);
not I_12873 (I221739,I276459);
nand I_12874 (I221756,I221739,I221674);
and I_12875 (I221773,I221739,I276453);
nand I_12876 (I221790,I221773,I276465);
nor I_12877 (I221555,I221790,I221739);
and I_12878 (I221546,I221632,I221790);
not I_12879 (I221835,I221790);
nand I_12880 (I221549,I221632,I221835);
nor I_12881 (I221543,I221598,I221790);
not I_12882 (I221880,I276471);
nor I_12883 (I221897,I221880,I276453);
nand I_12884 (I221914,I221897,I221739);
nor I_12885 (I221552,I221657,I221914);
nor I_12886 (I221945,I221880,I276450);
and I_12887 (I221962,I221945,I276468);
or I_12888 (I221979,I221962,I276474);
DFFARX1 I_12889 (I221979,I2859,I221572,I222005,);
nor I_12890 (I222013,I222005,I221756);
DFFARX1 I_12891 (I222013,I2859,I221572,I221540,);
DFFARX1 I_12892 (I222005,I2859,I221572,I221564,);
not I_12893 (I222058,I222005);
nor I_12894 (I222075,I222058,I221632);
nor I_12895 (I222092,I221897,I222075);
DFFARX1 I_12896 (I222092,I2859,I221572,I221561,);
not I_12897 (I222150,I2866);
DFFARX1 I_12898 (I415922,I2859,I222150,I222176,);
not I_12899 (I222184,I222176);
DFFARX1 I_12900 (I415913,I2859,I222150,I222210,);
not I_12901 (I222218,I415907);
nand I_12902 (I222235,I222218,I415919);
not I_12903 (I222252,I222235);
nor I_12904 (I222269,I222252,I415910);
nor I_12905 (I222286,I222184,I222269);
DFFARX1 I_12906 (I222286,I2859,I222150,I222136,);
not I_12907 (I222317,I415910);
nand I_12908 (I222334,I222317,I222252);
and I_12909 (I222351,I222317,I415916);
nand I_12910 (I222368,I222351,I415901);
nor I_12911 (I222133,I222368,I222317);
and I_12912 (I222124,I222210,I222368);
not I_12913 (I222413,I222368);
nand I_12914 (I222127,I222210,I222413);
nor I_12915 (I222121,I222176,I222368);
not I_12916 (I222458,I415901);
nor I_12917 (I222475,I222458,I415916);
nand I_12918 (I222492,I222475,I222317);
nor I_12919 (I222130,I222235,I222492);
nor I_12920 (I222523,I222458,I415904);
and I_12921 (I222540,I222523,I415907);
or I_12922 (I222557,I222540,I415904);
DFFARX1 I_12923 (I222557,I2859,I222150,I222583,);
nor I_12924 (I222591,I222583,I222334);
DFFARX1 I_12925 (I222591,I2859,I222150,I222118,);
DFFARX1 I_12926 (I222583,I2859,I222150,I222142,);
not I_12927 (I222636,I222583);
nor I_12928 (I222653,I222636,I222210);
nor I_12929 (I222670,I222475,I222653);
DFFARX1 I_12930 (I222670,I2859,I222150,I222139,);
not I_12931 (I222728,I2866);
DFFARX1 I_12932 (I136699,I2859,I222728,I222754,);
not I_12933 (I222762,I222754);
DFFARX1 I_12934 (I136714,I2859,I222728,I222788,);
not I_12935 (I222796,I136717);
nand I_12936 (I222813,I222796,I136696);
not I_12937 (I222830,I222813);
nor I_12938 (I222847,I222830,I136720);
nor I_12939 (I222864,I222762,I222847);
DFFARX1 I_12940 (I222864,I2859,I222728,I222714,);
not I_12941 (I222895,I136720);
nand I_12942 (I222912,I222895,I222830);
and I_12943 (I222929,I222895,I136702);
nand I_12944 (I222946,I222929,I136693);
nor I_12945 (I222711,I222946,I222895);
and I_12946 (I222702,I222788,I222946);
not I_12947 (I222991,I222946);
nand I_12948 (I222705,I222788,I222991);
nor I_12949 (I222699,I222754,I222946);
not I_12950 (I223036,I136693);
nor I_12951 (I223053,I223036,I136702);
nand I_12952 (I223070,I223053,I222895);
nor I_12953 (I222708,I222813,I223070);
nor I_12954 (I223101,I223036,I136708);
and I_12955 (I223118,I223101,I136711);
or I_12956 (I223135,I223118,I136705);
DFFARX1 I_12957 (I223135,I2859,I222728,I223161,);
nor I_12958 (I223169,I223161,I222912);
DFFARX1 I_12959 (I223169,I2859,I222728,I222696,);
DFFARX1 I_12960 (I223161,I2859,I222728,I222720,);
not I_12961 (I223214,I223161);
nor I_12962 (I223231,I223214,I222788);
nor I_12963 (I223248,I223053,I223231);
DFFARX1 I_12964 (I223248,I2859,I222728,I222717,);
not I_12965 (I223306,I2866);
DFFARX1 I_12966 (I527008,I2859,I223306,I223332,);
not I_12967 (I223340,I223332);
DFFARX1 I_12968 (I527020,I2859,I223306,I223366,);
not I_12969 (I223374,I527011);
nand I_12970 (I223391,I223374,I526999);
not I_12971 (I223408,I223391);
nor I_12972 (I223425,I223408,I526996);
nor I_12973 (I223442,I223340,I223425);
DFFARX1 I_12974 (I223442,I2859,I223306,I223292,);
not I_12975 (I223473,I526996);
nand I_12976 (I223490,I223473,I223408);
and I_12977 (I223507,I223473,I527002);
nand I_12978 (I223524,I223507,I526999);
nor I_12979 (I223289,I223524,I223473);
and I_12980 (I223280,I223366,I223524);
not I_12981 (I223569,I223524);
nand I_12982 (I223283,I223366,I223569);
nor I_12983 (I223277,I223332,I223524);
not I_12984 (I223614,I527017);
nor I_12985 (I223631,I223614,I527002);
nand I_12986 (I223648,I223631,I223473);
nor I_12987 (I223286,I223391,I223648);
nor I_12988 (I223679,I223614,I527005);
and I_12989 (I223696,I223679,I526996);
or I_12990 (I223713,I223696,I527014);
DFFARX1 I_12991 (I223713,I2859,I223306,I223739,);
nor I_12992 (I223747,I223739,I223490);
DFFARX1 I_12993 (I223747,I2859,I223306,I223274,);
DFFARX1 I_12994 (I223739,I2859,I223306,I223298,);
not I_12995 (I223792,I223739);
nor I_12996 (I223809,I223792,I223366);
nor I_12997 (I223826,I223631,I223809);
DFFARX1 I_12998 (I223826,I2859,I223306,I223295,);
not I_12999 (I223884,I2866);
DFFARX1 I_13000 (I387007,I2859,I223884,I223910,);
not I_13001 (I223918,I223910);
DFFARX1 I_13002 (I387004,I2859,I223884,I223944,);
not I_13003 (I223952,I387001);
nand I_13004 (I223969,I223952,I387028);
not I_13005 (I223986,I223969);
nor I_13006 (I224003,I223986,I387016);
nor I_13007 (I224020,I223918,I224003);
DFFARX1 I_13008 (I224020,I2859,I223884,I223870,);
not I_13009 (I224051,I387016);
nand I_13010 (I224068,I224051,I223986);
and I_13011 (I224085,I224051,I387022);
nand I_13012 (I224102,I224085,I387013);
nor I_13013 (I223867,I224102,I224051);
and I_13014 (I223858,I223944,I224102);
not I_13015 (I224147,I224102);
nand I_13016 (I223861,I223944,I224147);
nor I_13017 (I223855,I223910,I224102);
not I_13018 (I224192,I387010);
nor I_13019 (I224209,I224192,I387022);
nand I_13020 (I224226,I224209,I224051);
nor I_13021 (I223864,I223969,I224226);
nor I_13022 (I224257,I224192,I387025);
and I_13023 (I224274,I224257,I387019);
or I_13024 (I224291,I224274,I387001);
DFFARX1 I_13025 (I224291,I2859,I223884,I224317,);
nor I_13026 (I224325,I224317,I224068);
DFFARX1 I_13027 (I224325,I2859,I223884,I223852,);
DFFARX1 I_13028 (I224317,I2859,I223884,I223876,);
not I_13029 (I224370,I224317);
nor I_13030 (I224387,I224370,I223944);
nor I_13031 (I224404,I224209,I224387);
DFFARX1 I_13032 (I224404,I2859,I223884,I223873,);
not I_13033 (I224462,I2866);
DFFARX1 I_13034 (I64407,I2859,I224462,I224488,);
not I_13035 (I224496,I224488);
DFFARX1 I_13036 (I64392,I2859,I224462,I224522,);
not I_13037 (I224530,I64410);
nand I_13038 (I224547,I224530,I64395);
not I_13039 (I224564,I224547);
nor I_13040 (I224581,I224564,I64392);
nor I_13041 (I224598,I224496,I224581);
DFFARX1 I_13042 (I224598,I2859,I224462,I224448,);
not I_13043 (I224629,I64392);
nand I_13044 (I224646,I224629,I224564);
and I_13045 (I224663,I224629,I64395);
nand I_13046 (I224680,I224663,I64416);
nor I_13047 (I224445,I224680,I224629);
and I_13048 (I224436,I224522,I224680);
not I_13049 (I224725,I224680);
nand I_13050 (I224439,I224522,I224725);
nor I_13051 (I224433,I224488,I224680);
not I_13052 (I224770,I64404);
nor I_13053 (I224787,I224770,I64395);
nand I_13054 (I224804,I224787,I224629);
nor I_13055 (I224442,I224547,I224804);
nor I_13056 (I224835,I224770,I64398);
and I_13057 (I224852,I224835,I64413);
or I_13058 (I224869,I224852,I64401);
DFFARX1 I_13059 (I224869,I2859,I224462,I224895,);
nor I_13060 (I224903,I224895,I224646);
DFFARX1 I_13061 (I224903,I2859,I224462,I224430,);
DFFARX1 I_13062 (I224895,I2859,I224462,I224454,);
not I_13063 (I224948,I224895);
nor I_13064 (I224965,I224948,I224522);
nor I_13065 (I224982,I224787,I224965);
DFFARX1 I_13066 (I224982,I2859,I224462,I224451,);
not I_13067 (I225040,I2866);
DFFARX1 I_13068 (I277028,I2859,I225040,I225066,);
not I_13069 (I225074,I225066);
DFFARX1 I_13070 (I277040,I2859,I225040,I225100,);
not I_13071 (I225108,I277031);
nand I_13072 (I225125,I225108,I277034);
not I_13073 (I225142,I225125);
nor I_13074 (I225159,I225142,I277037);
nor I_13075 (I225176,I225074,I225159);
DFFARX1 I_13076 (I225176,I2859,I225040,I225026,);
not I_13077 (I225207,I277037);
nand I_13078 (I225224,I225207,I225142);
and I_13079 (I225241,I225207,I277031);
nand I_13080 (I225258,I225241,I277043);
nor I_13081 (I225023,I225258,I225207);
and I_13082 (I225014,I225100,I225258);
not I_13083 (I225303,I225258);
nand I_13084 (I225017,I225100,I225303);
nor I_13085 (I225011,I225066,I225258);
not I_13086 (I225348,I277049);
nor I_13087 (I225365,I225348,I277031);
nand I_13088 (I225382,I225365,I225207);
nor I_13089 (I225020,I225125,I225382);
nor I_13090 (I225413,I225348,I277028);
and I_13091 (I225430,I225413,I277046);
or I_13092 (I225447,I225430,I277052);
DFFARX1 I_13093 (I225447,I2859,I225040,I225473,);
nor I_13094 (I225481,I225473,I225224);
DFFARX1 I_13095 (I225481,I2859,I225040,I225008,);
DFFARX1 I_13096 (I225473,I2859,I225040,I225032,);
not I_13097 (I225526,I225473);
nor I_13098 (I225543,I225526,I225100);
nor I_13099 (I225560,I225365,I225543);
DFFARX1 I_13100 (I225560,I2859,I225040,I225029,);
not I_13101 (I225618,I2866);
DFFARX1 I_13102 (I325977,I2859,I225618,I225644,);
not I_13103 (I225652,I225644);
DFFARX1 I_13104 (I325977,I2859,I225618,I225678,);
not I_13105 (I225686,I325974);
nand I_13106 (I225703,I225686,I325989);
not I_13107 (I225720,I225703);
nor I_13108 (I225737,I225720,I325983);
nor I_13109 (I225754,I225652,I225737);
DFFARX1 I_13110 (I225754,I2859,I225618,I225604,);
not I_13111 (I225785,I325983);
nand I_13112 (I225802,I225785,I225720);
and I_13113 (I225819,I225785,I325980);
nand I_13114 (I225836,I225819,I325971);
nor I_13115 (I225601,I225836,I225785);
and I_13116 (I225592,I225678,I225836);
not I_13117 (I225881,I225836);
nand I_13118 (I225595,I225678,I225881);
nor I_13119 (I225589,I225644,I225836);
not I_13120 (I225926,I325992);
nor I_13121 (I225943,I225926,I325980);
nand I_13122 (I225960,I225943,I225785);
nor I_13123 (I225598,I225703,I225960);
nor I_13124 (I225991,I225926,I325971);
and I_13125 (I226008,I225991,I325974);
or I_13126 (I226025,I226008,I325986);
DFFARX1 I_13127 (I226025,I2859,I225618,I226051,);
nor I_13128 (I226059,I226051,I225802);
DFFARX1 I_13129 (I226059,I2859,I225618,I225586,);
DFFARX1 I_13130 (I226051,I2859,I225618,I225610,);
not I_13131 (I226104,I226051);
nor I_13132 (I226121,I226104,I225678);
nor I_13133 (I226138,I225943,I226121);
DFFARX1 I_13134 (I226138,I2859,I225618,I225607,);
not I_13135 (I226196,I2866);
DFFARX1 I_13136 (I336517,I2859,I226196,I226222,);
not I_13137 (I226230,I226222);
DFFARX1 I_13138 (I336517,I2859,I226196,I226256,);
not I_13139 (I226264,I336514);
nand I_13140 (I226281,I226264,I336529);
not I_13141 (I226298,I226281);
nor I_13142 (I226315,I226298,I336523);
nor I_13143 (I226332,I226230,I226315);
DFFARX1 I_13144 (I226332,I2859,I226196,I226182,);
not I_13145 (I226363,I336523);
nand I_13146 (I226380,I226363,I226298);
and I_13147 (I226397,I226363,I336520);
nand I_13148 (I226414,I226397,I336511);
nor I_13149 (I226179,I226414,I226363);
and I_13150 (I226170,I226256,I226414);
not I_13151 (I226459,I226414);
nand I_13152 (I226173,I226256,I226459);
nor I_13153 (I226167,I226222,I226414);
not I_13154 (I226504,I336532);
nor I_13155 (I226521,I226504,I336520);
nand I_13156 (I226538,I226521,I226363);
nor I_13157 (I226176,I226281,I226538);
nor I_13158 (I226569,I226504,I336511);
and I_13159 (I226586,I226569,I336514);
or I_13160 (I226603,I226586,I336526);
DFFARX1 I_13161 (I226603,I2859,I226196,I226629,);
nor I_13162 (I226637,I226629,I226380);
DFFARX1 I_13163 (I226637,I2859,I226196,I226164,);
DFFARX1 I_13164 (I226629,I2859,I226196,I226188,);
not I_13165 (I226682,I226629);
nor I_13166 (I226699,I226682,I226256);
nor I_13167 (I226716,I226521,I226699);
DFFARX1 I_13168 (I226716,I2859,I226196,I226185,);
not I_13169 (I226774,I2866);
DFFARX1 I_13170 (I441214,I2859,I226774,I226800,);
not I_13171 (I226808,I226800);
DFFARX1 I_13172 (I441220,I2859,I226774,I226834,);
not I_13173 (I226842,I441214);
nand I_13174 (I226859,I226842,I441217);
not I_13175 (I226876,I226859);
nor I_13176 (I226893,I226876,I441235);
nor I_13177 (I226910,I226808,I226893);
DFFARX1 I_13178 (I226910,I2859,I226774,I226760,);
not I_13179 (I226941,I441235);
nand I_13180 (I226958,I226941,I226876);
and I_13181 (I226975,I226941,I441238);
nand I_13182 (I226992,I226975,I441217);
nor I_13183 (I226757,I226992,I226941);
and I_13184 (I226748,I226834,I226992);
not I_13185 (I227037,I226992);
nand I_13186 (I226751,I226834,I227037);
nor I_13187 (I226745,I226800,I226992);
not I_13188 (I227082,I441223);
nor I_13189 (I227099,I227082,I441238);
nand I_13190 (I227116,I227099,I226941);
nor I_13191 (I226754,I226859,I227116);
nor I_13192 (I227147,I227082,I441229);
and I_13193 (I227164,I227147,I441226);
or I_13194 (I227181,I227164,I441232);
DFFARX1 I_13195 (I227181,I2859,I226774,I227207,);
nor I_13196 (I227215,I227207,I226958);
DFFARX1 I_13197 (I227215,I2859,I226774,I226742,);
DFFARX1 I_13198 (I227207,I2859,I226774,I226766,);
not I_13199 (I227260,I227207);
nor I_13200 (I227277,I227260,I226834);
nor I_13201 (I227294,I227099,I227277);
DFFARX1 I_13202 (I227294,I2859,I226774,I226763,);
not I_13203 (I227352,I2866);
DFFARX1 I_13204 (I296102,I2859,I227352,I227378,);
not I_13205 (I227386,I227378);
DFFARX1 I_13206 (I296114,I2859,I227352,I227412,);
not I_13207 (I227420,I296105);
nand I_13208 (I227437,I227420,I296108);
not I_13209 (I227454,I227437);
nor I_13210 (I227471,I227454,I296111);
nor I_13211 (I227488,I227386,I227471);
DFFARX1 I_13212 (I227488,I2859,I227352,I227338,);
not I_13213 (I227519,I296111);
nand I_13214 (I227536,I227519,I227454);
and I_13215 (I227553,I227519,I296105);
nand I_13216 (I227570,I227553,I296117);
nor I_13217 (I227335,I227570,I227519);
and I_13218 (I227326,I227412,I227570);
not I_13219 (I227615,I227570);
nand I_13220 (I227329,I227412,I227615);
nor I_13221 (I227323,I227378,I227570);
not I_13222 (I227660,I296123);
nor I_13223 (I227677,I227660,I296105);
nand I_13224 (I227694,I227677,I227519);
nor I_13225 (I227332,I227437,I227694);
nor I_13226 (I227725,I227660,I296102);
and I_13227 (I227742,I227725,I296120);
or I_13228 (I227759,I227742,I296126);
DFFARX1 I_13229 (I227759,I2859,I227352,I227785,);
nor I_13230 (I227793,I227785,I227536);
DFFARX1 I_13231 (I227793,I2859,I227352,I227320,);
DFFARX1 I_13232 (I227785,I2859,I227352,I227344,);
not I_13233 (I227838,I227785);
nor I_13234 (I227855,I227838,I227412);
nor I_13235 (I227872,I227677,I227855);
DFFARX1 I_13236 (I227872,I2859,I227352,I227341,);
not I_13237 (I227930,I2866);
DFFARX1 I_13238 (I112984,I2859,I227930,I227956,);
not I_13239 (I227964,I227956);
DFFARX1 I_13240 (I112999,I2859,I227930,I227990,);
not I_13241 (I227998,I113002);
nand I_13242 (I228015,I227998,I112981);
not I_13243 (I228032,I228015);
nor I_13244 (I228049,I228032,I113005);
nor I_13245 (I228066,I227964,I228049);
DFFARX1 I_13246 (I228066,I2859,I227930,I227916,);
not I_13247 (I228097,I113005);
nand I_13248 (I228114,I228097,I228032);
and I_13249 (I228131,I228097,I112987);
nand I_13250 (I228148,I228131,I112978);
nor I_13251 (I227913,I228148,I228097);
and I_13252 (I227904,I227990,I228148);
not I_13253 (I228193,I228148);
nand I_13254 (I227907,I227990,I228193);
nor I_13255 (I227901,I227956,I228148);
not I_13256 (I228238,I112978);
nor I_13257 (I228255,I228238,I112987);
nand I_13258 (I228272,I228255,I228097);
nor I_13259 (I227910,I228015,I228272);
nor I_13260 (I228303,I228238,I112993);
and I_13261 (I228320,I228303,I112996);
or I_13262 (I228337,I228320,I112990);
DFFARX1 I_13263 (I228337,I2859,I227930,I228363,);
nor I_13264 (I228371,I228363,I228114);
DFFARX1 I_13265 (I228371,I2859,I227930,I227898,);
DFFARX1 I_13266 (I228363,I2859,I227930,I227922,);
not I_13267 (I228416,I228363);
nor I_13268 (I228433,I228416,I227990);
nor I_13269 (I228450,I228255,I228433);
DFFARX1 I_13270 (I228450,I2859,I227930,I227919,);
not I_13271 (I228508,I2866);
DFFARX1 I_13272 (I307084,I2859,I228508,I228534,);
not I_13273 (I228542,I228534);
DFFARX1 I_13274 (I307096,I2859,I228508,I228568,);
not I_13275 (I228576,I307087);
nand I_13276 (I228593,I228576,I307090);
not I_13277 (I228610,I228593);
nor I_13278 (I228627,I228610,I307093);
nor I_13279 (I228644,I228542,I228627);
DFFARX1 I_13280 (I228644,I2859,I228508,I228494,);
not I_13281 (I228675,I307093);
nand I_13282 (I228692,I228675,I228610);
and I_13283 (I228709,I228675,I307087);
nand I_13284 (I228726,I228709,I307099);
nor I_13285 (I228491,I228726,I228675);
and I_13286 (I228482,I228568,I228726);
not I_13287 (I228771,I228726);
nand I_13288 (I228485,I228568,I228771);
nor I_13289 (I228479,I228534,I228726);
not I_13290 (I228816,I307105);
nor I_13291 (I228833,I228816,I307087);
nand I_13292 (I228850,I228833,I228675);
nor I_13293 (I228488,I228593,I228850);
nor I_13294 (I228881,I228816,I307084);
and I_13295 (I228898,I228881,I307102);
or I_13296 (I228915,I228898,I307108);
DFFARX1 I_13297 (I228915,I2859,I228508,I228941,);
nor I_13298 (I228949,I228941,I228692);
DFFARX1 I_13299 (I228949,I2859,I228508,I228476,);
DFFARX1 I_13300 (I228941,I2859,I228508,I228500,);
not I_13301 (I228994,I228941);
nor I_13302 (I229011,I228994,I228568);
nor I_13303 (I229028,I228833,I229011);
DFFARX1 I_13304 (I229028,I2859,I228508,I228497,);
not I_13305 (I229086,I2866);
DFFARX1 I_13306 (I309396,I2859,I229086,I229112,);
not I_13307 (I229120,I229112);
DFFARX1 I_13308 (I309408,I2859,I229086,I229146,);
not I_13309 (I229154,I309399);
nand I_13310 (I229171,I229154,I309402);
not I_13311 (I229188,I229171);
nor I_13312 (I229205,I229188,I309405);
nor I_13313 (I229222,I229120,I229205);
DFFARX1 I_13314 (I229222,I2859,I229086,I229072,);
not I_13315 (I229253,I309405);
nand I_13316 (I229270,I229253,I229188);
and I_13317 (I229287,I229253,I309399);
nand I_13318 (I229304,I229287,I309411);
nor I_13319 (I229069,I229304,I229253);
and I_13320 (I229060,I229146,I229304);
not I_13321 (I229349,I229304);
nand I_13322 (I229063,I229146,I229349);
nor I_13323 (I229057,I229112,I229304);
not I_13324 (I229394,I309417);
nor I_13325 (I229411,I229394,I309399);
nand I_13326 (I229428,I229411,I229253);
nor I_13327 (I229066,I229171,I229428);
nor I_13328 (I229459,I229394,I309396);
and I_13329 (I229476,I229459,I309414);
or I_13330 (I229493,I229476,I309420);
DFFARX1 I_13331 (I229493,I2859,I229086,I229519,);
nor I_13332 (I229527,I229519,I229270);
DFFARX1 I_13333 (I229527,I2859,I229086,I229054,);
DFFARX1 I_13334 (I229519,I2859,I229086,I229078,);
not I_13335 (I229572,I229519);
nor I_13336 (I229589,I229572,I229146);
nor I_13337 (I229606,I229411,I229589);
DFFARX1 I_13338 (I229606,I2859,I229086,I229075,);
not I_13339 (I229664,I2866);
DFFARX1 I_13340 (I327558,I2859,I229664,I229690,);
not I_13341 (I229698,I229690);
DFFARX1 I_13342 (I327558,I2859,I229664,I229724,);
not I_13343 (I229732,I327555);
nand I_13344 (I229749,I229732,I327570);
not I_13345 (I229766,I229749);
nor I_13346 (I229783,I229766,I327564);
nor I_13347 (I229800,I229698,I229783);
DFFARX1 I_13348 (I229800,I2859,I229664,I229650,);
not I_13349 (I229831,I327564);
nand I_13350 (I229848,I229831,I229766);
and I_13351 (I229865,I229831,I327561);
nand I_13352 (I229882,I229865,I327552);
nor I_13353 (I229647,I229882,I229831);
and I_13354 (I229638,I229724,I229882);
not I_13355 (I229927,I229882);
nand I_13356 (I229641,I229724,I229927);
nor I_13357 (I229635,I229690,I229882);
not I_13358 (I229972,I327573);
nor I_13359 (I229989,I229972,I327561);
nand I_13360 (I230006,I229989,I229831);
nor I_13361 (I229644,I229749,I230006);
nor I_13362 (I230037,I229972,I327552);
and I_13363 (I230054,I230037,I327555);
or I_13364 (I230071,I230054,I327567);
DFFARX1 I_13365 (I230071,I2859,I229664,I230097,);
nor I_13366 (I230105,I230097,I229848);
DFFARX1 I_13367 (I230105,I2859,I229664,I229632,);
DFFARX1 I_13368 (I230097,I2859,I229664,I229656,);
not I_13369 (I230150,I230097);
nor I_13370 (I230167,I230150,I229724);
nor I_13371 (I230184,I229989,I230167);
DFFARX1 I_13372 (I230184,I2859,I229664,I229653,);
not I_13373 (I230242,I2866);
DFFARX1 I_13374 (I459710,I2859,I230242,I230268,);
not I_13375 (I230276,I230268);
DFFARX1 I_13376 (I459716,I2859,I230242,I230302,);
not I_13377 (I230310,I459710);
nand I_13378 (I230327,I230310,I459713);
not I_13379 (I230344,I230327);
nor I_13380 (I230361,I230344,I459731);
nor I_13381 (I230378,I230276,I230361);
DFFARX1 I_13382 (I230378,I2859,I230242,I230228,);
not I_13383 (I230409,I459731);
nand I_13384 (I230426,I230409,I230344);
and I_13385 (I230443,I230409,I459734);
nand I_13386 (I230460,I230443,I459713);
nor I_13387 (I230225,I230460,I230409);
and I_13388 (I230216,I230302,I230460);
not I_13389 (I230505,I230460);
nand I_13390 (I230219,I230302,I230505);
nor I_13391 (I230213,I230268,I230460);
not I_13392 (I230550,I459719);
nor I_13393 (I230567,I230550,I459734);
nand I_13394 (I230584,I230567,I230409);
nor I_13395 (I230222,I230327,I230584);
nor I_13396 (I230615,I230550,I459725);
and I_13397 (I230632,I230615,I459722);
or I_13398 (I230649,I230632,I459728);
DFFARX1 I_13399 (I230649,I2859,I230242,I230675,);
nor I_13400 (I230683,I230675,I230426);
DFFARX1 I_13401 (I230683,I2859,I230242,I230210,);
DFFARX1 I_13402 (I230675,I2859,I230242,I230234,);
not I_13403 (I230728,I230675);
nor I_13404 (I230745,I230728,I230302);
nor I_13405 (I230762,I230567,I230745);
DFFARX1 I_13406 (I230762,I2859,I230242,I230231,);
not I_13407 (I230820,I2866);
DFFARX1 I_13408 (I116673,I2859,I230820,I230846,);
not I_13409 (I230854,I230846);
DFFARX1 I_13410 (I116688,I2859,I230820,I230880,);
not I_13411 (I230888,I116691);
nand I_13412 (I230905,I230888,I116670);
not I_13413 (I230922,I230905);
nor I_13414 (I230939,I230922,I116694);
nor I_13415 (I230956,I230854,I230939);
DFFARX1 I_13416 (I230956,I2859,I230820,I230806,);
not I_13417 (I230987,I116694);
nand I_13418 (I231004,I230987,I230922);
and I_13419 (I231021,I230987,I116676);
nand I_13420 (I231038,I231021,I116667);
nor I_13421 (I230803,I231038,I230987);
and I_13422 (I230794,I230880,I231038);
not I_13423 (I231083,I231038);
nand I_13424 (I230797,I230880,I231083);
nor I_13425 (I230791,I230846,I231038);
not I_13426 (I231128,I116667);
nor I_13427 (I231145,I231128,I116676);
nand I_13428 (I231162,I231145,I230987);
nor I_13429 (I230800,I230905,I231162);
nor I_13430 (I231193,I231128,I116682);
and I_13431 (I231210,I231193,I116685);
or I_13432 (I231227,I231210,I116679);
DFFARX1 I_13433 (I231227,I2859,I230820,I231253,);
nor I_13434 (I231261,I231253,I231004);
DFFARX1 I_13435 (I231261,I2859,I230820,I230788,);
DFFARX1 I_13436 (I231253,I2859,I230820,I230812,);
not I_13437 (I231306,I231253);
nor I_13438 (I231323,I231306,I230880);
nor I_13439 (I231340,I231145,I231323);
DFFARX1 I_13440 (I231340,I2859,I230820,I230809,);
not I_13441 (I231398,I2866);
DFFARX1 I_13442 (I19570,I2859,I231398,I231424,);
not I_13443 (I231432,I231424);
DFFARX1 I_13444 (I19549,I2859,I231398,I231458,);
not I_13445 (I231466,I19546);
nand I_13446 (I231483,I231466,I19561);
not I_13447 (I231500,I231483);
nor I_13448 (I231517,I231500,I19549);
nor I_13449 (I231534,I231432,I231517);
DFFARX1 I_13450 (I231534,I2859,I231398,I231384,);
not I_13451 (I231565,I19549);
nand I_13452 (I231582,I231565,I231500);
and I_13453 (I231599,I231565,I19552);
nand I_13454 (I231616,I231599,I19567);
nor I_13455 (I231381,I231616,I231565);
and I_13456 (I231372,I231458,I231616);
not I_13457 (I231661,I231616);
nand I_13458 (I231375,I231458,I231661);
nor I_13459 (I231369,I231424,I231616);
not I_13460 (I231706,I19558);
nor I_13461 (I231723,I231706,I19552);
nand I_13462 (I231740,I231723,I231565);
nor I_13463 (I231378,I231483,I231740);
nor I_13464 (I231771,I231706,I19546);
and I_13465 (I231788,I231771,I19555);
or I_13466 (I231805,I231788,I19564);
DFFARX1 I_13467 (I231805,I2859,I231398,I231831,);
nor I_13468 (I231839,I231831,I231582);
DFFARX1 I_13469 (I231839,I2859,I231398,I231366,);
DFFARX1 I_13470 (I231831,I2859,I231398,I231390,);
not I_13471 (I231884,I231831);
nor I_13472 (I231901,I231884,I231458);
nor I_13473 (I231918,I231723,I231901);
DFFARX1 I_13474 (I231918,I2859,I231398,I231387,);
not I_13475 (I231976,I2866);
DFFARX1 I_13476 (I438362,I2859,I231976,I232002,);
not I_13477 (I232010,I232002);
DFFARX1 I_13478 (I438353,I2859,I231976,I232036,);
not I_13479 (I232044,I438347);
nand I_13480 (I232061,I232044,I438359);
not I_13481 (I232078,I232061);
nor I_13482 (I232095,I232078,I438350);
nor I_13483 (I232112,I232010,I232095);
DFFARX1 I_13484 (I232112,I2859,I231976,I231962,);
not I_13485 (I232143,I438350);
nand I_13486 (I232160,I232143,I232078);
and I_13487 (I232177,I232143,I438356);
nand I_13488 (I232194,I232177,I438341);
nor I_13489 (I231959,I232194,I232143);
and I_13490 (I231950,I232036,I232194);
not I_13491 (I232239,I232194);
nand I_13492 (I231953,I232036,I232239);
nor I_13493 (I231947,I232002,I232194);
not I_13494 (I232284,I438341);
nor I_13495 (I232301,I232284,I438356);
nand I_13496 (I232318,I232301,I232143);
nor I_13497 (I231956,I232061,I232318);
nor I_13498 (I232349,I232284,I438344);
and I_13499 (I232366,I232349,I438347);
or I_13500 (I232383,I232366,I438344);
DFFARX1 I_13501 (I232383,I2859,I231976,I232409,);
nor I_13502 (I232417,I232409,I232160);
DFFARX1 I_13503 (I232417,I2859,I231976,I231944,);
DFFARX1 I_13504 (I232409,I2859,I231976,I231968,);
not I_13505 (I232462,I232409);
nor I_13506 (I232479,I232462,I232036);
nor I_13507 (I232496,I232301,I232479);
DFFARX1 I_13508 (I232496,I2859,I231976,I231965,);
not I_13509 (I232554,I2866);
DFFARX1 I_13510 (I311130,I2859,I232554,I232580,);
not I_13511 (I232588,I232580);
DFFARX1 I_13512 (I311142,I2859,I232554,I232614,);
not I_13513 (I232622,I311133);
nand I_13514 (I232639,I232622,I311136);
not I_13515 (I232656,I232639);
nor I_13516 (I232673,I232656,I311139);
nor I_13517 (I232690,I232588,I232673);
DFFARX1 I_13518 (I232690,I2859,I232554,I232540,);
not I_13519 (I232721,I311139);
nand I_13520 (I232738,I232721,I232656);
and I_13521 (I232755,I232721,I311133);
nand I_13522 (I232772,I232755,I311145);
nor I_13523 (I232537,I232772,I232721);
and I_13524 (I232528,I232614,I232772);
not I_13525 (I232817,I232772);
nand I_13526 (I232531,I232614,I232817);
nor I_13527 (I232525,I232580,I232772);
not I_13528 (I232862,I311151);
nor I_13529 (I232879,I232862,I311133);
nand I_13530 (I232896,I232879,I232721);
nor I_13531 (I232534,I232639,I232896);
nor I_13532 (I232927,I232862,I311130);
and I_13533 (I232944,I232927,I311148);
or I_13534 (I232961,I232944,I311154);
DFFARX1 I_13535 (I232961,I2859,I232554,I232987,);
nor I_13536 (I232995,I232987,I232738);
DFFARX1 I_13537 (I232995,I2859,I232554,I232522,);
DFFARX1 I_13538 (I232987,I2859,I232554,I232546,);
not I_13539 (I233040,I232987);
nor I_13540 (I233057,I233040,I232614);
nor I_13541 (I233074,I232879,I233057);
DFFARX1 I_13542 (I233074,I2859,I232554,I232543,);
not I_13543 (I233132,I2866);
DFFARX1 I_13544 (I46447,I2859,I233132,I233158,);
not I_13545 (I233166,I233158);
DFFARX1 I_13546 (I46426,I2859,I233132,I233192,);
not I_13547 (I233200,I46423);
nand I_13548 (I233217,I233200,I46438);
not I_13549 (I233234,I233217);
nor I_13550 (I233251,I233234,I46426);
nor I_13551 (I233268,I233166,I233251);
DFFARX1 I_13552 (I233268,I2859,I233132,I233118,);
not I_13553 (I233299,I46426);
nand I_13554 (I233316,I233299,I233234);
and I_13555 (I233333,I233299,I46429);
nand I_13556 (I233350,I233333,I46444);
nor I_13557 (I233115,I233350,I233299);
and I_13558 (I233106,I233192,I233350);
not I_13559 (I233395,I233350);
nand I_13560 (I233109,I233192,I233395);
nor I_13561 (I233103,I233158,I233350);
not I_13562 (I233440,I46435);
nor I_13563 (I233457,I233440,I46429);
nand I_13564 (I233474,I233457,I233299);
nor I_13565 (I233112,I233217,I233474);
nor I_13566 (I233505,I233440,I46423);
and I_13567 (I233522,I233505,I46432);
or I_13568 (I233539,I233522,I46441);
DFFARX1 I_13569 (I233539,I2859,I233132,I233565,);
nor I_13570 (I233573,I233565,I233316);
DFFARX1 I_13571 (I233573,I2859,I233132,I233100,);
DFFARX1 I_13572 (I233565,I2859,I233132,I233124,);
not I_13573 (I233618,I233565);
nor I_13574 (I233635,I233618,I233192);
nor I_13575 (I233652,I233457,I233635);
DFFARX1 I_13576 (I233652,I2859,I233132,I233121,);
not I_13577 (I233710,I2866);
DFFARX1 I_13578 (I114038,I2859,I233710,I233736,);
not I_13579 (I233744,I233736);
DFFARX1 I_13580 (I114053,I2859,I233710,I233770,);
not I_13581 (I233778,I114056);
nand I_13582 (I233795,I233778,I114035);
not I_13583 (I233812,I233795);
nor I_13584 (I233829,I233812,I114059);
nor I_13585 (I233846,I233744,I233829);
DFFARX1 I_13586 (I233846,I2859,I233710,I233696,);
not I_13587 (I233877,I114059);
nand I_13588 (I233894,I233877,I233812);
and I_13589 (I233911,I233877,I114041);
nand I_13590 (I233928,I233911,I114032);
nor I_13591 (I233693,I233928,I233877);
and I_13592 (I233684,I233770,I233928);
not I_13593 (I233973,I233928);
nand I_13594 (I233687,I233770,I233973);
nor I_13595 (I233681,I233736,I233928);
not I_13596 (I234018,I114032);
nor I_13597 (I234035,I234018,I114041);
nand I_13598 (I234052,I234035,I233877);
nor I_13599 (I233690,I233795,I234052);
nor I_13600 (I234083,I234018,I114047);
and I_13601 (I234100,I234083,I114050);
or I_13602 (I234117,I234100,I114044);
DFFARX1 I_13603 (I234117,I2859,I233710,I234143,);
nor I_13604 (I234151,I234143,I233894);
DFFARX1 I_13605 (I234151,I2859,I233710,I233678,);
DFFARX1 I_13606 (I234143,I2859,I233710,I233702,);
not I_13607 (I234196,I234143);
nor I_13608 (I234213,I234196,I233770);
nor I_13609 (I234230,I234035,I234213);
DFFARX1 I_13610 (I234230,I2859,I233710,I233699,);
not I_13611 (I234288,I2866);
DFFARX1 I_13612 (I51323,I2859,I234288,I234314,);
not I_13613 (I234322,I234314);
DFFARX1 I_13614 (I51302,I2859,I234288,I234348,);
not I_13615 (I234356,I51302);
nand I_13616 (I234373,I234356,I51329);
not I_13617 (I234390,I234373);
nor I_13618 (I234407,I234390,I51305);
nor I_13619 (I234424,I234322,I234407);
DFFARX1 I_13620 (I234424,I2859,I234288,I234274,);
not I_13621 (I234455,I51305);
nand I_13622 (I234472,I234455,I234390);
and I_13623 (I234489,I234455,I51326);
nand I_13624 (I234506,I234489,I51308);
nor I_13625 (I234271,I234506,I234455);
and I_13626 (I234262,I234348,I234506);
not I_13627 (I234551,I234506);
nand I_13628 (I234265,I234348,I234551);
nor I_13629 (I234259,I234314,I234506);
not I_13630 (I234596,I51311);
nor I_13631 (I234613,I234596,I51326);
nand I_13632 (I234630,I234613,I234455);
nor I_13633 (I234268,I234373,I234630);
nor I_13634 (I234661,I234596,I51317);
and I_13635 (I234678,I234661,I51314);
or I_13636 (I234695,I234678,I51320);
DFFARX1 I_13637 (I234695,I2859,I234288,I234721,);
nor I_13638 (I234729,I234721,I234472);
DFFARX1 I_13639 (I234729,I2859,I234288,I234256,);
DFFARX1 I_13640 (I234721,I2859,I234288,I234280,);
not I_13641 (I234774,I234721);
nor I_13642 (I234791,I234774,I234348);
nor I_13643 (I234808,I234613,I234791);
DFFARX1 I_13644 (I234808,I2859,I234288,I234277,);
not I_13645 (I234866,I2866);
DFFARX1 I_13646 (I71547,I2859,I234866,I234892,);
not I_13647 (I234900,I234892);
DFFARX1 I_13648 (I71532,I2859,I234866,I234926,);
not I_13649 (I234934,I71550);
nand I_13650 (I234951,I234934,I71535);
not I_13651 (I234968,I234951);
nor I_13652 (I234985,I234968,I71532);
nor I_13653 (I235002,I234900,I234985);
DFFARX1 I_13654 (I235002,I2859,I234866,I234852,);
not I_13655 (I235033,I71532);
nand I_13656 (I235050,I235033,I234968);
and I_13657 (I235067,I235033,I71535);
nand I_13658 (I235084,I235067,I71556);
nor I_13659 (I234849,I235084,I235033);
and I_13660 (I234840,I234926,I235084);
not I_13661 (I235129,I235084);
nand I_13662 (I234843,I234926,I235129);
nor I_13663 (I234837,I234892,I235084);
not I_13664 (I235174,I71544);
nor I_13665 (I235191,I235174,I71535);
nand I_13666 (I235208,I235191,I235033);
nor I_13667 (I234846,I234951,I235208);
nor I_13668 (I235239,I235174,I71538);
and I_13669 (I235256,I235239,I71553);
or I_13670 (I235273,I235256,I71541);
DFFARX1 I_13671 (I235273,I2859,I234866,I235299,);
nor I_13672 (I235307,I235299,I235050);
DFFARX1 I_13673 (I235307,I2859,I234866,I234834,);
DFFARX1 I_13674 (I235299,I2859,I234866,I234858,);
not I_13675 (I235352,I235299);
nor I_13676 (I235369,I235352,I234926);
nor I_13677 (I235386,I235191,I235369);
DFFARX1 I_13678 (I235386,I2859,I234866,I234855,);
not I_13679 (I235444,I2866);
DFFARX1 I_13680 (I45920,I2859,I235444,I235470,);
not I_13681 (I235478,I235470);
DFFARX1 I_13682 (I45899,I2859,I235444,I235504,);
not I_13683 (I235512,I45896);
nand I_13684 (I235529,I235512,I45911);
not I_13685 (I235546,I235529);
nor I_13686 (I235563,I235546,I45899);
nor I_13687 (I235580,I235478,I235563);
DFFARX1 I_13688 (I235580,I2859,I235444,I235430,);
not I_13689 (I235611,I45899);
nand I_13690 (I235628,I235611,I235546);
and I_13691 (I235645,I235611,I45902);
nand I_13692 (I235662,I235645,I45917);
nor I_13693 (I235427,I235662,I235611);
and I_13694 (I235418,I235504,I235662);
not I_13695 (I235707,I235662);
nand I_13696 (I235421,I235504,I235707);
nor I_13697 (I235415,I235470,I235662);
not I_13698 (I235752,I45908);
nor I_13699 (I235769,I235752,I45902);
nand I_13700 (I235786,I235769,I235611);
nor I_13701 (I235424,I235529,I235786);
nor I_13702 (I235817,I235752,I45896);
and I_13703 (I235834,I235817,I45905);
or I_13704 (I235851,I235834,I45914);
DFFARX1 I_13705 (I235851,I2859,I235444,I235877,);
nor I_13706 (I235885,I235877,I235628);
DFFARX1 I_13707 (I235885,I2859,I235444,I235412,);
DFFARX1 I_13708 (I235877,I2859,I235444,I235436,);
not I_13709 (I235930,I235877);
nor I_13710 (I235947,I235930,I235504);
nor I_13711 (I235964,I235769,I235947);
DFFARX1 I_13712 (I235964,I2859,I235444,I235433,);
not I_13713 (I236022,I2866);
DFFARX1 I_13714 (I474738,I2859,I236022,I236048,);
not I_13715 (I236056,I236048);
DFFARX1 I_13716 (I474744,I2859,I236022,I236082,);
not I_13717 (I236090,I474738);
nand I_13718 (I236107,I236090,I474741);
not I_13719 (I236124,I236107);
nor I_13720 (I236141,I236124,I474759);
nor I_13721 (I236158,I236056,I236141);
DFFARX1 I_13722 (I236158,I2859,I236022,I236008,);
not I_13723 (I236189,I474759);
nand I_13724 (I236206,I236189,I236124);
and I_13725 (I236223,I236189,I474762);
nand I_13726 (I236240,I236223,I474741);
nor I_13727 (I236005,I236240,I236189);
and I_13728 (I235996,I236082,I236240);
not I_13729 (I236285,I236240);
nand I_13730 (I235999,I236082,I236285);
nor I_13731 (I235993,I236048,I236240);
not I_13732 (I236330,I474747);
nor I_13733 (I236347,I236330,I474762);
nand I_13734 (I236364,I236347,I236189);
nor I_13735 (I236002,I236107,I236364);
nor I_13736 (I236395,I236330,I474753);
and I_13737 (I236412,I236395,I474750);
or I_13738 (I236429,I236412,I474756);
DFFARX1 I_13739 (I236429,I2859,I236022,I236455,);
nor I_13740 (I236463,I236455,I236206);
DFFARX1 I_13741 (I236463,I2859,I236022,I235990,);
DFFARX1 I_13742 (I236455,I2859,I236022,I236014,);
not I_13743 (I236508,I236455);
nor I_13744 (I236525,I236508,I236082);
nor I_13745 (I236542,I236347,I236525);
DFFARX1 I_13746 (I236542,I2859,I236022,I236011,);
not I_13747 (I236600,I2866);
DFFARX1 I_13748 (I511204,I2859,I236600,I236626,);
not I_13749 (I236634,I236626);
DFFARX1 I_13750 (I511198,I2859,I236600,I236660,);
not I_13751 (I236668,I511207);
nand I_13752 (I236685,I236668,I511186);
not I_13753 (I236702,I236685);
nor I_13754 (I236719,I236702,I511195);
nor I_13755 (I236736,I236634,I236719);
DFFARX1 I_13756 (I236736,I2859,I236600,I236586,);
not I_13757 (I236767,I511195);
nand I_13758 (I236784,I236767,I236702);
and I_13759 (I236801,I236767,I511210);
nand I_13760 (I236818,I236801,I511189);
nor I_13761 (I236583,I236818,I236767);
and I_13762 (I236574,I236660,I236818);
not I_13763 (I236863,I236818);
nand I_13764 (I236577,I236660,I236863);
nor I_13765 (I236571,I236626,I236818);
not I_13766 (I236908,I511192);
nor I_13767 (I236925,I236908,I511210);
nand I_13768 (I236942,I236925,I236767);
nor I_13769 (I236580,I236685,I236942);
nor I_13770 (I236973,I236908,I511201);
and I_13771 (I236990,I236973,I511189);
or I_13772 (I237007,I236990,I511186);
DFFARX1 I_13773 (I237007,I2859,I236600,I237033,);
nor I_13774 (I237041,I237033,I236784);
DFFARX1 I_13775 (I237041,I2859,I236600,I236568,);
DFFARX1 I_13776 (I237033,I2859,I236600,I236592,);
not I_13777 (I237086,I237033);
nor I_13778 (I237103,I237086,I236660);
nor I_13779 (I237120,I236925,I237103);
DFFARX1 I_13780 (I237120,I2859,I236600,I236589,);
not I_13781 (I237178,I2866);
DFFARX1 I_13782 (I16387,I2859,I237178,I237204,);
not I_13783 (I237212,I237204);
DFFARX1 I_13784 (I16390,I2859,I237178,I237238,);
not I_13785 (I237246,I16384);
nand I_13786 (I237263,I237246,I16408);
not I_13787 (I237280,I237263);
nor I_13788 (I237297,I237280,I16387);
nor I_13789 (I237314,I237212,I237297);
DFFARX1 I_13790 (I237314,I2859,I237178,I237164,);
not I_13791 (I237345,I16387);
nand I_13792 (I237362,I237345,I237280);
and I_13793 (I237379,I237345,I16402);
nand I_13794 (I237396,I237379,I16396);
nor I_13795 (I237161,I237396,I237345);
and I_13796 (I237152,I237238,I237396);
not I_13797 (I237441,I237396);
nand I_13798 (I237155,I237238,I237441);
nor I_13799 (I237149,I237204,I237396);
not I_13800 (I237486,I16405);
nor I_13801 (I237503,I237486,I16402);
nand I_13802 (I237520,I237503,I237345);
nor I_13803 (I237158,I237263,I237520);
nor I_13804 (I237551,I237486,I16384);
and I_13805 (I237568,I237551,I16393);
or I_13806 (I237585,I237568,I16399);
DFFARX1 I_13807 (I237585,I2859,I237178,I237611,);
nor I_13808 (I237619,I237611,I237362);
DFFARX1 I_13809 (I237619,I2859,I237178,I237146,);
DFFARX1 I_13810 (I237611,I2859,I237178,I237170,);
not I_13811 (I237664,I237611);
nor I_13812 (I237681,I237664,I237238);
nor I_13813 (I237698,I237503,I237681);
DFFARX1 I_13814 (I237698,I2859,I237178,I237167,);
not I_13815 (I237756,I2866);
DFFARX1 I_13816 (I528742,I2859,I237756,I237782,);
not I_13817 (I237790,I237782);
DFFARX1 I_13818 (I528754,I2859,I237756,I237816,);
not I_13819 (I237824,I528745);
nand I_13820 (I237841,I237824,I528733);
not I_13821 (I237858,I237841);
nor I_13822 (I237875,I237858,I528730);
nor I_13823 (I237892,I237790,I237875);
DFFARX1 I_13824 (I237892,I2859,I237756,I237742,);
not I_13825 (I237923,I528730);
nand I_13826 (I237940,I237923,I237858);
and I_13827 (I237957,I237923,I528736);
nand I_13828 (I237974,I237957,I528733);
nor I_13829 (I237739,I237974,I237923);
and I_13830 (I237730,I237816,I237974);
not I_13831 (I238019,I237974);
nand I_13832 (I237733,I237816,I238019);
nor I_13833 (I237727,I237782,I237974);
not I_13834 (I238064,I528751);
nor I_13835 (I238081,I238064,I528736);
nand I_13836 (I238098,I238081,I237923);
nor I_13837 (I237736,I237841,I238098);
nor I_13838 (I238129,I238064,I528739);
and I_13839 (I238146,I238129,I528730);
or I_13840 (I238163,I238146,I528748);
DFFARX1 I_13841 (I238163,I2859,I237756,I238189,);
nor I_13842 (I238197,I238189,I237940);
DFFARX1 I_13843 (I238197,I2859,I237756,I237724,);
DFFARX1 I_13844 (I238189,I2859,I237756,I237748,);
not I_13845 (I238242,I238189);
nor I_13846 (I238259,I238242,I237816);
nor I_13847 (I238276,I238081,I238259);
DFFARX1 I_13848 (I238276,I2859,I237756,I237745,);
not I_13849 (I238334,I2866);
DFFARX1 I_13850 (I315754,I2859,I238334,I238360,);
not I_13851 (I238368,I238360);
DFFARX1 I_13852 (I315766,I2859,I238334,I238394,);
not I_13853 (I238402,I315757);
nand I_13854 (I238419,I238402,I315760);
not I_13855 (I238436,I238419);
nor I_13856 (I238453,I238436,I315763);
nor I_13857 (I238470,I238368,I238453);
DFFARX1 I_13858 (I238470,I2859,I238334,I238320,);
not I_13859 (I238501,I315763);
nand I_13860 (I238518,I238501,I238436);
and I_13861 (I238535,I238501,I315757);
nand I_13862 (I238552,I238535,I315769);
nor I_13863 (I238317,I238552,I238501);
and I_13864 (I238308,I238394,I238552);
not I_13865 (I238597,I238552);
nand I_13866 (I238311,I238394,I238597);
nor I_13867 (I238305,I238360,I238552);
not I_13868 (I238642,I315775);
nor I_13869 (I238659,I238642,I315757);
nand I_13870 (I238676,I238659,I238501);
nor I_13871 (I238314,I238419,I238676);
nor I_13872 (I238707,I238642,I315754);
and I_13873 (I238724,I238707,I315772);
or I_13874 (I238741,I238724,I315778);
DFFARX1 I_13875 (I238741,I2859,I238334,I238767,);
nor I_13876 (I238775,I238767,I238518);
DFFARX1 I_13877 (I238775,I2859,I238334,I238302,);
DFFARX1 I_13878 (I238767,I2859,I238334,I238326,);
not I_13879 (I238820,I238767);
nor I_13880 (I238837,I238820,I238394);
nor I_13881 (I238854,I238659,I238837);
DFFARX1 I_13882 (I238854,I2859,I238334,I238323,);
not I_13883 (I238912,I2866);
DFFARX1 I_13884 (I75712,I2859,I238912,I238938,);
not I_13885 (I238946,I238938);
DFFARX1 I_13886 (I75697,I2859,I238912,I238972,);
not I_13887 (I238980,I75715);
nand I_13888 (I238997,I238980,I75700);
not I_13889 (I239014,I238997);
nor I_13890 (I239031,I239014,I75697);
nor I_13891 (I239048,I238946,I239031);
DFFARX1 I_13892 (I239048,I2859,I238912,I238898,);
not I_13893 (I239079,I75697);
nand I_13894 (I239096,I239079,I239014);
and I_13895 (I239113,I239079,I75700);
nand I_13896 (I239130,I239113,I75721);
nor I_13897 (I238895,I239130,I239079);
and I_13898 (I238886,I238972,I239130);
not I_13899 (I239175,I239130);
nand I_13900 (I238889,I238972,I239175);
nor I_13901 (I238883,I238938,I239130);
not I_13902 (I239220,I75709);
nor I_13903 (I239237,I239220,I75700);
nand I_13904 (I239254,I239237,I239079);
nor I_13905 (I238892,I238997,I239254);
nor I_13906 (I239285,I239220,I75703);
and I_13907 (I239302,I239285,I75718);
or I_13908 (I239319,I239302,I75706);
DFFARX1 I_13909 (I239319,I2859,I238912,I239345,);
nor I_13910 (I239353,I239345,I239096);
DFFARX1 I_13911 (I239353,I2859,I238912,I238880,);
DFFARX1 I_13912 (I239345,I2859,I238912,I238904,);
not I_13913 (I239398,I239345);
nor I_13914 (I239415,I239398,I238972);
nor I_13915 (I239432,I239237,I239415);
DFFARX1 I_13916 (I239432,I2859,I238912,I238901,);
not I_13917 (I239490,I2866);
DFFARX1 I_13918 (I164228,I2859,I239490,I239516,);
not I_13919 (I239524,I239516);
DFFARX1 I_13920 (I164240,I2859,I239490,I239550,);
not I_13921 (I239558,I164216);
nand I_13922 (I239575,I239558,I164243);
not I_13923 (I239592,I239575);
nor I_13924 (I239609,I239592,I164231);
nor I_13925 (I239626,I239524,I239609);
DFFARX1 I_13926 (I239626,I2859,I239490,I239476,);
not I_13927 (I239657,I164231);
nand I_13928 (I239674,I239657,I239592);
and I_13929 (I239691,I239657,I164216);
nand I_13930 (I239708,I239691,I164219);
nor I_13931 (I239473,I239708,I239657);
and I_13932 (I239464,I239550,I239708);
not I_13933 (I239753,I239708);
nand I_13934 (I239467,I239550,I239753);
nor I_13935 (I239461,I239516,I239708);
not I_13936 (I239798,I164225);
nor I_13937 (I239815,I239798,I164216);
nand I_13938 (I239832,I239815,I239657);
nor I_13939 (I239470,I239575,I239832);
nor I_13940 (I239863,I239798,I164234);
and I_13941 (I239880,I239863,I164222);
or I_13942 (I239897,I239880,I164237);
DFFARX1 I_13943 (I239897,I2859,I239490,I239923,);
nor I_13944 (I239931,I239923,I239674);
DFFARX1 I_13945 (I239931,I2859,I239490,I239458,);
DFFARX1 I_13946 (I239923,I2859,I239490,I239482,);
not I_13947 (I239976,I239923);
nor I_13948 (I239993,I239976,I239550);
nor I_13949 (I240010,I239815,I239993);
DFFARX1 I_13950 (I240010,I2859,I239490,I239479,);
not I_13951 (I240068,I2866);
DFFARX1 I_13952 (I262578,I2859,I240068,I240094,);
not I_13953 (I240102,I240094);
DFFARX1 I_13954 (I262590,I2859,I240068,I240128,);
not I_13955 (I240136,I262581);
nand I_13956 (I240153,I240136,I262584);
not I_13957 (I240170,I240153);
nor I_13958 (I240187,I240170,I262587);
nor I_13959 (I240204,I240102,I240187);
DFFARX1 I_13960 (I240204,I2859,I240068,I240054,);
not I_13961 (I240235,I262587);
nand I_13962 (I240252,I240235,I240170);
and I_13963 (I240269,I240235,I262581);
nand I_13964 (I240286,I240269,I262593);
nor I_13965 (I240051,I240286,I240235);
and I_13966 (I240042,I240128,I240286);
not I_13967 (I240331,I240286);
nand I_13968 (I240045,I240128,I240331);
nor I_13969 (I240039,I240094,I240286);
not I_13970 (I240376,I262599);
nor I_13971 (I240393,I240376,I262581);
nand I_13972 (I240410,I240393,I240235);
nor I_13973 (I240048,I240153,I240410);
nor I_13974 (I240441,I240376,I262578);
and I_13975 (I240458,I240441,I262596);
or I_13976 (I240475,I240458,I262602);
DFFARX1 I_13977 (I240475,I2859,I240068,I240501,);
nor I_13978 (I240509,I240501,I240252);
DFFARX1 I_13979 (I240509,I2859,I240068,I240036,);
DFFARX1 I_13980 (I240501,I2859,I240068,I240060,);
not I_13981 (I240554,I240501);
nor I_13982 (I240571,I240554,I240128);
nor I_13983 (I240588,I240393,I240571);
DFFARX1 I_13984 (I240588,I2859,I240068,I240057,);
not I_13985 (I240646,I2866);
DFFARX1 I_13986 (I183812,I2859,I240646,I240672,);
not I_13987 (I240680,I240672);
DFFARX1 I_13988 (I183824,I2859,I240646,I240706,);
not I_13989 (I240714,I183800);
nand I_13990 (I240731,I240714,I183827);
not I_13991 (I240748,I240731);
nor I_13992 (I240765,I240748,I183815);
nor I_13993 (I240782,I240680,I240765);
DFFARX1 I_13994 (I240782,I2859,I240646,I240632,);
not I_13995 (I240813,I183815);
nand I_13996 (I240830,I240813,I240748);
and I_13997 (I240847,I240813,I183800);
nand I_13998 (I240864,I240847,I183803);
nor I_13999 (I240629,I240864,I240813);
and I_14000 (I240620,I240706,I240864);
not I_14001 (I240909,I240864);
nand I_14002 (I240623,I240706,I240909);
nor I_14003 (I240617,I240672,I240864);
not I_14004 (I240954,I183809);
nor I_14005 (I240971,I240954,I183800);
nand I_14006 (I240988,I240971,I240813);
nor I_14007 (I240626,I240731,I240988);
nor I_14008 (I241019,I240954,I183818);
and I_14009 (I241036,I241019,I183806);
or I_14010 (I241053,I241036,I183821);
DFFARX1 I_14011 (I241053,I2859,I240646,I241079,);
nor I_14012 (I241087,I241079,I240830);
DFFARX1 I_14013 (I241087,I2859,I240646,I240614,);
DFFARX1 I_14014 (I241079,I2859,I240646,I240638,);
not I_14015 (I241132,I241079);
nor I_14016 (I241149,I241132,I240706);
nor I_14017 (I241166,I240971,I241149);
DFFARX1 I_14018 (I241166,I2859,I240646,I240635,);
not I_14019 (I241224,I2866);
DFFARX1 I_14020 (I291478,I2859,I241224,I241250,);
not I_14021 (I241258,I241250);
DFFARX1 I_14022 (I291490,I2859,I241224,I241284,);
not I_14023 (I241292,I291481);
nand I_14024 (I241309,I241292,I291484);
not I_14025 (I241326,I241309);
nor I_14026 (I241343,I241326,I291487);
nor I_14027 (I241360,I241258,I241343);
DFFARX1 I_14028 (I241360,I2859,I241224,I241210,);
not I_14029 (I241391,I291487);
nand I_14030 (I241408,I241391,I241326);
and I_14031 (I241425,I241391,I291481);
nand I_14032 (I241442,I241425,I291493);
nor I_14033 (I241207,I241442,I241391);
and I_14034 (I241198,I241284,I241442);
not I_14035 (I241487,I241442);
nand I_14036 (I241201,I241284,I241487);
nor I_14037 (I241195,I241250,I241442);
not I_14038 (I241532,I291499);
nor I_14039 (I241549,I241532,I291481);
nand I_14040 (I241566,I241549,I241391);
nor I_14041 (I241204,I241309,I241566);
nor I_14042 (I241597,I241532,I291478);
and I_14043 (I241614,I241597,I291496);
or I_14044 (I241631,I241614,I291502);
DFFARX1 I_14045 (I241631,I2859,I241224,I241657,);
nor I_14046 (I241665,I241657,I241408);
DFFARX1 I_14047 (I241665,I2859,I241224,I241192,);
DFFARX1 I_14048 (I241657,I2859,I241224,I241216,);
not I_14049 (I241710,I241657);
nor I_14050 (I241727,I241710,I241284);
nor I_14051 (I241744,I241549,I241727);
DFFARX1 I_14052 (I241744,I2859,I241224,I241213,);
not I_14053 (I241802,I2866);
DFFARX1 I_14054 (I487454,I2859,I241802,I241828,);
not I_14055 (I241836,I241828);
DFFARX1 I_14056 (I487460,I2859,I241802,I241862,);
not I_14057 (I241870,I487454);
nand I_14058 (I241887,I241870,I487457);
not I_14059 (I241904,I241887);
nor I_14060 (I241921,I241904,I487475);
nor I_14061 (I241938,I241836,I241921);
DFFARX1 I_14062 (I241938,I2859,I241802,I241788,);
not I_14063 (I241969,I487475);
nand I_14064 (I241986,I241969,I241904);
and I_14065 (I242003,I241969,I487478);
nand I_14066 (I242020,I242003,I487457);
nor I_14067 (I241785,I242020,I241969);
and I_14068 (I241776,I241862,I242020);
not I_14069 (I242065,I242020);
nand I_14070 (I241779,I241862,I242065);
nor I_14071 (I241773,I241828,I242020);
not I_14072 (I242110,I487463);
nor I_14073 (I242127,I242110,I487478);
nand I_14074 (I242144,I242127,I241969);
nor I_14075 (I241782,I241887,I242144);
nor I_14076 (I242175,I242110,I487469);
and I_14077 (I242192,I242175,I487466);
or I_14078 (I242209,I242192,I487472);
DFFARX1 I_14079 (I242209,I2859,I241802,I242235,);
nor I_14080 (I242243,I242235,I241986);
DFFARX1 I_14081 (I242243,I2859,I241802,I241770,);
DFFARX1 I_14082 (I242235,I2859,I241802,I241794,);
not I_14083 (I242288,I242235);
nor I_14084 (I242305,I242288,I241862);
nor I_14085 (I242322,I242127,I242305);
DFFARX1 I_14086 (I242322,I2859,I241802,I241791,);
not I_14087 (I242380,I2866);
DFFARX1 I_14088 (I447572,I2859,I242380,I242406,);
not I_14089 (I242414,I242406);
DFFARX1 I_14090 (I447578,I2859,I242380,I242440,);
not I_14091 (I242448,I447572);
nand I_14092 (I242465,I242448,I447575);
not I_14093 (I242482,I242465);
nor I_14094 (I242499,I242482,I447593);
nor I_14095 (I242516,I242414,I242499);
DFFARX1 I_14096 (I242516,I2859,I242380,I242366,);
not I_14097 (I242547,I447593);
nand I_14098 (I242564,I242547,I242482);
and I_14099 (I242581,I242547,I447596);
nand I_14100 (I242598,I242581,I447575);
nor I_14101 (I242363,I242598,I242547);
and I_14102 (I242354,I242440,I242598);
not I_14103 (I242643,I242598);
nand I_14104 (I242357,I242440,I242643);
nor I_14105 (I242351,I242406,I242598);
not I_14106 (I242688,I447581);
nor I_14107 (I242705,I242688,I447596);
nand I_14108 (I242722,I242705,I242547);
nor I_14109 (I242360,I242465,I242722);
nor I_14110 (I242753,I242688,I447587);
and I_14111 (I242770,I242753,I447584);
or I_14112 (I242787,I242770,I447590);
DFFARX1 I_14113 (I242787,I2859,I242380,I242813,);
nor I_14114 (I242821,I242813,I242564);
DFFARX1 I_14115 (I242821,I2859,I242380,I242348,);
DFFARX1 I_14116 (I242813,I2859,I242380,I242372,);
not I_14117 (I242866,I242813);
nor I_14118 (I242883,I242866,I242440);
nor I_14119 (I242900,I242705,I242883);
DFFARX1 I_14120 (I242900,I2859,I242380,I242369,);
not I_14121 (I242958,I2866);
DFFARX1 I_14122 (I349692,I2859,I242958,I242984,);
not I_14123 (I242992,I242984);
DFFARX1 I_14124 (I349692,I2859,I242958,I243018,);
not I_14125 (I243026,I349689);
nand I_14126 (I243043,I243026,I349704);
not I_14127 (I243060,I243043);
nor I_14128 (I243077,I243060,I349698);
nor I_14129 (I243094,I242992,I243077);
DFFARX1 I_14130 (I243094,I2859,I242958,I242944,);
not I_14131 (I243125,I349698);
nand I_14132 (I243142,I243125,I243060);
and I_14133 (I243159,I243125,I349695);
nand I_14134 (I243176,I243159,I349686);
nor I_14135 (I242941,I243176,I243125);
and I_14136 (I242932,I243018,I243176);
not I_14137 (I243221,I243176);
nand I_14138 (I242935,I243018,I243221);
nor I_14139 (I242929,I242984,I243176);
not I_14140 (I243266,I349707);
nor I_14141 (I243283,I243266,I349695);
nand I_14142 (I243300,I243283,I243125);
nor I_14143 (I242938,I243043,I243300);
nor I_14144 (I243331,I243266,I349686);
and I_14145 (I243348,I243331,I349689);
or I_14146 (I243365,I243348,I349701);
DFFARX1 I_14147 (I243365,I2859,I242958,I243391,);
nor I_14148 (I243399,I243391,I243142);
DFFARX1 I_14149 (I243399,I2859,I242958,I242926,);
DFFARX1 I_14150 (I243391,I2859,I242958,I242950,);
not I_14151 (I243444,I243391);
nor I_14152 (I243461,I243444,I243018);
nor I_14153 (I243478,I243283,I243461);
DFFARX1 I_14154 (I243478,I2859,I242958,I242947,);
not I_14155 (I243536,I2866);
DFFARX1 I_14156 (I103677,I2859,I243536,I243562,);
not I_14157 (I243570,I243562);
DFFARX1 I_14158 (I103662,I2859,I243536,I243596,);
not I_14159 (I243604,I103680);
nand I_14160 (I243621,I243604,I103665);
not I_14161 (I243638,I243621);
nor I_14162 (I243655,I243638,I103662);
nor I_14163 (I243672,I243570,I243655);
DFFARX1 I_14164 (I243672,I2859,I243536,I243522,);
not I_14165 (I243703,I103662);
nand I_14166 (I243720,I243703,I243638);
and I_14167 (I243737,I243703,I103665);
nand I_14168 (I243754,I243737,I103686);
nor I_14169 (I243519,I243754,I243703);
and I_14170 (I243510,I243596,I243754);
not I_14171 (I243799,I243754);
nand I_14172 (I243513,I243596,I243799);
nor I_14173 (I243507,I243562,I243754);
not I_14174 (I243844,I103674);
nor I_14175 (I243861,I243844,I103665);
nand I_14176 (I243878,I243861,I243703);
nor I_14177 (I243516,I243621,I243878);
nor I_14178 (I243909,I243844,I103668);
and I_14179 (I243926,I243909,I103683);
or I_14180 (I243943,I243926,I103671);
DFFARX1 I_14181 (I243943,I2859,I243536,I243969,);
nor I_14182 (I243977,I243969,I243720);
DFFARX1 I_14183 (I243977,I2859,I243536,I243504,);
DFFARX1 I_14184 (I243969,I2859,I243536,I243528,);
not I_14185 (I244022,I243969);
nor I_14186 (I244039,I244022,I243596);
nor I_14187 (I244056,I243861,I244039);
DFFARX1 I_14188 (I244056,I2859,I243536,I243525,);
not I_14189 (I244114,I2866);
DFFARX1 I_14190 (I34326,I2859,I244114,I244140,);
not I_14191 (I244148,I244140);
DFFARX1 I_14192 (I34305,I2859,I244114,I244174,);
not I_14193 (I244182,I34302);
nand I_14194 (I244199,I244182,I34317);
not I_14195 (I244216,I244199);
nor I_14196 (I244233,I244216,I34305);
nor I_14197 (I244250,I244148,I244233);
DFFARX1 I_14198 (I244250,I2859,I244114,I244100,);
not I_14199 (I244281,I34305);
nand I_14200 (I244298,I244281,I244216);
and I_14201 (I244315,I244281,I34308);
nand I_14202 (I244332,I244315,I34323);
nor I_14203 (I244097,I244332,I244281);
and I_14204 (I244088,I244174,I244332);
not I_14205 (I244377,I244332);
nand I_14206 (I244091,I244174,I244377);
nor I_14207 (I244085,I244140,I244332);
not I_14208 (I244422,I34314);
nor I_14209 (I244439,I244422,I34308);
nand I_14210 (I244456,I244439,I244281);
nor I_14211 (I244094,I244199,I244456);
nor I_14212 (I244487,I244422,I34302);
and I_14213 (I244504,I244487,I34311);
or I_14214 (I244521,I244504,I34320);
DFFARX1 I_14215 (I244521,I2859,I244114,I244547,);
nor I_14216 (I244555,I244547,I244298);
DFFARX1 I_14217 (I244555,I2859,I244114,I244082,);
DFFARX1 I_14218 (I244547,I2859,I244114,I244106,);
not I_14219 (I244600,I244547);
nor I_14220 (I244617,I244600,I244174);
nor I_14221 (I244634,I244439,I244617);
DFFARX1 I_14222 (I244634,I2859,I244114,I244103,);
not I_14223 (I244692,I2866);
DFFARX1 I_14224 (I568935,I2859,I244692,I244718,);
not I_14225 (I244726,I244718);
DFFARX1 I_14226 (I568935,I2859,I244692,I244752,);
not I_14227 (I244760,I568959);
nand I_14228 (I244777,I244760,I568941);
not I_14229 (I244794,I244777);
nor I_14230 (I244811,I244794,I568956);
nor I_14231 (I244828,I244726,I244811);
DFFARX1 I_14232 (I244828,I2859,I244692,I244678,);
not I_14233 (I244859,I568956);
nand I_14234 (I244876,I244859,I244794);
and I_14235 (I244893,I244859,I568938);
nand I_14236 (I244910,I244893,I568947);
nor I_14237 (I244675,I244910,I244859);
and I_14238 (I244666,I244752,I244910);
not I_14239 (I244955,I244910);
nand I_14240 (I244669,I244752,I244955);
nor I_14241 (I244663,I244718,I244910);
not I_14242 (I245000,I568944);
nor I_14243 (I245017,I245000,I568938);
nand I_14244 (I245034,I245017,I244859);
nor I_14245 (I244672,I244777,I245034);
nor I_14246 (I245065,I245000,I568953);
and I_14247 (I245082,I245065,I568962);
or I_14248 (I245099,I245082,I568950);
DFFARX1 I_14249 (I245099,I2859,I244692,I245125,);
nor I_14250 (I245133,I245125,I244876);
DFFARX1 I_14251 (I245133,I2859,I244692,I244660,);
DFFARX1 I_14252 (I245125,I2859,I244692,I244684,);
not I_14253 (I245178,I245125);
nor I_14254 (I245195,I245178,I244752);
nor I_14255 (I245212,I245017,I245195);
DFFARX1 I_14256 (I245212,I2859,I244692,I244681,);
not I_14257 (I245270,I2866);
DFFARX1 I_14258 (I191972,I2859,I245270,I245296,);
not I_14259 (I245304,I245296);
DFFARX1 I_14260 (I191984,I2859,I245270,I245330,);
not I_14261 (I245338,I191960);
nand I_14262 (I245355,I245338,I191987);
not I_14263 (I245372,I245355);
nor I_14264 (I245389,I245372,I191975);
nor I_14265 (I245406,I245304,I245389);
DFFARX1 I_14266 (I245406,I2859,I245270,I245256,);
not I_14267 (I245437,I191975);
nand I_14268 (I245454,I245437,I245372);
and I_14269 (I245471,I245437,I191960);
nand I_14270 (I245488,I245471,I191963);
nor I_14271 (I245253,I245488,I245437);
and I_14272 (I245244,I245330,I245488);
not I_14273 (I245533,I245488);
nand I_14274 (I245247,I245330,I245533);
nor I_14275 (I245241,I245296,I245488);
not I_14276 (I245578,I191969);
nor I_14277 (I245595,I245578,I191960);
nand I_14278 (I245612,I245595,I245437);
nor I_14279 (I245250,I245355,I245612);
nor I_14280 (I245643,I245578,I191978);
and I_14281 (I245660,I245643,I191966);
or I_14282 (I245677,I245660,I191981);
DFFARX1 I_14283 (I245677,I2859,I245270,I245703,);
nor I_14284 (I245711,I245703,I245454);
DFFARX1 I_14285 (I245711,I2859,I245270,I245238,);
DFFARX1 I_14286 (I245703,I2859,I245270,I245262,);
not I_14287 (I245756,I245703);
nor I_14288 (I245773,I245756,I245330);
nor I_14289 (I245790,I245595,I245773);
DFFARX1 I_14290 (I245790,I2859,I245270,I245259,);
not I_14291 (I245848,I2866);
DFFARX1 I_14292 (I308240,I2859,I245848,I245874,);
not I_14293 (I245882,I245874);
DFFARX1 I_14294 (I308252,I2859,I245848,I245908,);
not I_14295 (I245916,I308243);
nand I_14296 (I245933,I245916,I308246);
not I_14297 (I245950,I245933);
nor I_14298 (I245967,I245950,I308249);
nor I_14299 (I245984,I245882,I245967);
DFFARX1 I_14300 (I245984,I2859,I245848,I245834,);
not I_14301 (I246015,I308249);
nand I_14302 (I246032,I246015,I245950);
and I_14303 (I246049,I246015,I308243);
nand I_14304 (I246066,I246049,I308255);
nor I_14305 (I245831,I246066,I246015);
and I_14306 (I245822,I245908,I246066);
not I_14307 (I246111,I246066);
nand I_14308 (I245825,I245908,I246111);
nor I_14309 (I245819,I245874,I246066);
not I_14310 (I246156,I308261);
nor I_14311 (I246173,I246156,I308243);
nand I_14312 (I246190,I246173,I246015);
nor I_14313 (I245828,I245933,I246190);
nor I_14314 (I246221,I246156,I308240);
and I_14315 (I246238,I246221,I308258);
or I_14316 (I246255,I246238,I308264);
DFFARX1 I_14317 (I246255,I2859,I245848,I246281,);
nor I_14318 (I246289,I246281,I246032);
DFFARX1 I_14319 (I246289,I2859,I245848,I245816,);
DFFARX1 I_14320 (I246281,I2859,I245848,I245840,);
not I_14321 (I246334,I246281);
nor I_14322 (I246351,I246334,I245908);
nor I_14323 (I246368,I246173,I246351);
DFFARX1 I_14324 (I246368,I2859,I245848,I245837,);
not I_14325 (I246426,I2866);
DFFARX1 I_14326 (I513924,I2859,I246426,I246452,);
not I_14327 (I246460,I246452);
DFFARX1 I_14328 (I513918,I2859,I246426,I246486,);
not I_14329 (I246494,I513927);
nand I_14330 (I246511,I246494,I513906);
not I_14331 (I246528,I246511);
nor I_14332 (I246545,I246528,I513915);
nor I_14333 (I246562,I246460,I246545);
DFFARX1 I_14334 (I246562,I2859,I246426,I246412,);
not I_14335 (I246593,I513915);
nand I_14336 (I246610,I246593,I246528);
and I_14337 (I246627,I246593,I513930);
nand I_14338 (I246644,I246627,I513909);
nor I_14339 (I246409,I246644,I246593);
and I_14340 (I246400,I246486,I246644);
not I_14341 (I246689,I246644);
nand I_14342 (I246403,I246486,I246689);
nor I_14343 (I246397,I246452,I246644);
not I_14344 (I246734,I513912);
nor I_14345 (I246751,I246734,I513930);
nand I_14346 (I246768,I246751,I246593);
nor I_14347 (I246406,I246511,I246768);
nor I_14348 (I246799,I246734,I513921);
and I_14349 (I246816,I246799,I513909);
or I_14350 (I246833,I246816,I513906);
DFFARX1 I_14351 (I246833,I2859,I246426,I246859,);
nor I_14352 (I246867,I246859,I246610);
DFFARX1 I_14353 (I246867,I2859,I246426,I246394,);
DFFARX1 I_14354 (I246859,I2859,I246426,I246418,);
not I_14355 (I246912,I246859);
nor I_14356 (I246929,I246912,I246486);
nor I_14357 (I246946,I246751,I246929);
DFFARX1 I_14358 (I246946,I2859,I246426,I246415,);
not I_14359 (I247004,I2866);
DFFARX1 I_14360 (I264890,I2859,I247004,I247030,);
not I_14361 (I247038,I247030);
DFFARX1 I_14362 (I264902,I2859,I247004,I247064,);
not I_14363 (I247072,I264893);
nand I_14364 (I247089,I247072,I264896);
not I_14365 (I247106,I247089);
nor I_14366 (I247123,I247106,I264899);
nor I_14367 (I247140,I247038,I247123);
DFFARX1 I_14368 (I247140,I2859,I247004,I246990,);
not I_14369 (I247171,I264899);
nand I_14370 (I247188,I247171,I247106);
and I_14371 (I247205,I247171,I264893);
nand I_14372 (I247222,I247205,I264905);
nor I_14373 (I246987,I247222,I247171);
and I_14374 (I246978,I247064,I247222);
not I_14375 (I247267,I247222);
nand I_14376 (I246981,I247064,I247267);
nor I_14377 (I246975,I247030,I247222);
not I_14378 (I247312,I264911);
nor I_14379 (I247329,I247312,I264893);
nand I_14380 (I247346,I247329,I247171);
nor I_14381 (I246984,I247089,I247346);
nor I_14382 (I247377,I247312,I264890);
and I_14383 (I247394,I247377,I264908);
or I_14384 (I247411,I247394,I264914);
DFFARX1 I_14385 (I247411,I2859,I247004,I247437,);
nor I_14386 (I247445,I247437,I247188);
DFFARX1 I_14387 (I247445,I2859,I247004,I246972,);
DFFARX1 I_14388 (I247437,I2859,I247004,I246996,);
not I_14389 (I247490,I247437);
nor I_14390 (I247507,I247490,I247064);
nor I_14391 (I247524,I247329,I247507);
DFFARX1 I_14392 (I247524,I2859,I247004,I246993,);
not I_14393 (I247582,I2866);
DFFARX1 I_14394 (I277606,I2859,I247582,I247608,);
not I_14395 (I247616,I247608);
DFFARX1 I_14396 (I277618,I2859,I247582,I247642,);
not I_14397 (I247650,I277609);
nand I_14398 (I247667,I247650,I277612);
not I_14399 (I247684,I247667);
nor I_14400 (I247701,I247684,I277615);
nor I_14401 (I247718,I247616,I247701);
DFFARX1 I_14402 (I247718,I2859,I247582,I247568,);
not I_14403 (I247749,I277615);
nand I_14404 (I247766,I247749,I247684);
and I_14405 (I247783,I247749,I277609);
nand I_14406 (I247800,I247783,I277621);
nor I_14407 (I247565,I247800,I247749);
and I_14408 (I247556,I247642,I247800);
not I_14409 (I247845,I247800);
nand I_14410 (I247559,I247642,I247845);
nor I_14411 (I247553,I247608,I247800);
not I_14412 (I247890,I277627);
nor I_14413 (I247907,I247890,I277609);
nand I_14414 (I247924,I247907,I247749);
nor I_14415 (I247562,I247667,I247924);
nor I_14416 (I247955,I247890,I277606);
and I_14417 (I247972,I247955,I277624);
or I_14418 (I247989,I247972,I277630);
DFFARX1 I_14419 (I247989,I2859,I247582,I248015,);
nor I_14420 (I248023,I248015,I247766);
DFFARX1 I_14421 (I248023,I2859,I247582,I247550,);
DFFARX1 I_14422 (I248015,I2859,I247582,I247574,);
not I_14423 (I248068,I248015);
nor I_14424 (I248085,I248068,I247642);
nor I_14425 (I248102,I247907,I248085);
DFFARX1 I_14426 (I248102,I2859,I247582,I247571,);
not I_14427 (I248160,I2866);
DFFARX1 I_14428 (I508484,I2859,I248160,I248186,);
not I_14429 (I248194,I248186);
DFFARX1 I_14430 (I508478,I2859,I248160,I248220,);
not I_14431 (I248228,I508487);
nand I_14432 (I248245,I248228,I508466);
not I_14433 (I248262,I248245);
nor I_14434 (I248279,I248262,I508475);
nor I_14435 (I248296,I248194,I248279);
DFFARX1 I_14436 (I248296,I2859,I248160,I248146,);
not I_14437 (I248327,I508475);
nand I_14438 (I248344,I248327,I248262);
and I_14439 (I248361,I248327,I508490);
nand I_14440 (I248378,I248361,I508469);
nor I_14441 (I248143,I248378,I248327);
and I_14442 (I248134,I248220,I248378);
not I_14443 (I248423,I248378);
nand I_14444 (I248137,I248220,I248423);
nor I_14445 (I248131,I248186,I248378);
not I_14446 (I248468,I508472);
nor I_14447 (I248485,I248468,I508490);
nand I_14448 (I248502,I248485,I248327);
nor I_14449 (I248140,I248245,I248502);
nor I_14450 (I248533,I248468,I508481);
and I_14451 (I248550,I248533,I508469);
or I_14452 (I248567,I248550,I508466);
DFFARX1 I_14453 (I248567,I2859,I248160,I248593,);
nor I_14454 (I248601,I248593,I248344);
DFFARX1 I_14455 (I248601,I2859,I248160,I248128,);
DFFARX1 I_14456 (I248593,I2859,I248160,I248152,);
not I_14457 (I248646,I248593);
nor I_14458 (I248663,I248646,I248220);
nor I_14459 (I248680,I248485,I248663);
DFFARX1 I_14460 (I248680,I2859,I248160,I248149,);
not I_14461 (I248738,I2866);
DFFARX1 I_14462 (I499014,I2859,I248738,I248764,);
not I_14463 (I248772,I248764);
DFFARX1 I_14464 (I499020,I2859,I248738,I248798,);
not I_14465 (I248806,I499014);
nand I_14466 (I248823,I248806,I499017);
not I_14467 (I248840,I248823);
nor I_14468 (I248857,I248840,I499035);
nor I_14469 (I248874,I248772,I248857);
DFFARX1 I_14470 (I248874,I2859,I248738,I248724,);
not I_14471 (I248905,I499035);
nand I_14472 (I248922,I248905,I248840);
and I_14473 (I248939,I248905,I499038);
nand I_14474 (I248956,I248939,I499017);
nor I_14475 (I248721,I248956,I248905);
and I_14476 (I248712,I248798,I248956);
not I_14477 (I249001,I248956);
nand I_14478 (I248715,I248798,I249001);
nor I_14479 (I248709,I248764,I248956);
not I_14480 (I249046,I499023);
nor I_14481 (I249063,I249046,I499038);
nand I_14482 (I249080,I249063,I248905);
nor I_14483 (I248718,I248823,I249080);
nor I_14484 (I249111,I249046,I499029);
and I_14485 (I249128,I249111,I499026);
or I_14486 (I249145,I249128,I499032);
DFFARX1 I_14487 (I249145,I2859,I248738,I249171,);
nor I_14488 (I249179,I249171,I248922);
DFFARX1 I_14489 (I249179,I2859,I248738,I248706,);
DFFARX1 I_14490 (I249171,I2859,I248738,I248730,);
not I_14491 (I249224,I249171);
nor I_14492 (I249241,I249224,I248798);
nor I_14493 (I249258,I249063,I249241);
DFFARX1 I_14494 (I249258,I2859,I248738,I248727,);
not I_14495 (I249316,I2866);
DFFARX1 I_14496 (I185988,I2859,I249316,I249342,);
not I_14497 (I249350,I249342);
DFFARX1 I_14498 (I186000,I2859,I249316,I249376,);
not I_14499 (I249384,I185976);
nand I_14500 (I249401,I249384,I186003);
not I_14501 (I249418,I249401);
nor I_14502 (I249435,I249418,I185991);
nor I_14503 (I249452,I249350,I249435);
DFFARX1 I_14504 (I249452,I2859,I249316,I249302,);
not I_14505 (I249483,I185991);
nand I_14506 (I249500,I249483,I249418);
and I_14507 (I249517,I249483,I185976);
nand I_14508 (I249534,I249517,I185979);
nor I_14509 (I249299,I249534,I249483);
and I_14510 (I249290,I249376,I249534);
not I_14511 (I249579,I249534);
nand I_14512 (I249293,I249376,I249579);
nor I_14513 (I249287,I249342,I249534);
not I_14514 (I249624,I185985);
nor I_14515 (I249641,I249624,I185976);
nand I_14516 (I249658,I249641,I249483);
nor I_14517 (I249296,I249401,I249658);
nor I_14518 (I249689,I249624,I185994);
and I_14519 (I249706,I249689,I185982);
or I_14520 (I249723,I249706,I185997);
DFFARX1 I_14521 (I249723,I2859,I249316,I249749,);
nor I_14522 (I249757,I249749,I249500);
DFFARX1 I_14523 (I249757,I2859,I249316,I249284,);
DFFARX1 I_14524 (I249749,I2859,I249316,I249308,);
not I_14525 (I249802,I249749);
nor I_14526 (I249819,I249802,I249376);
nor I_14527 (I249836,I249641,I249819);
DFFARX1 I_14528 (I249836,I2859,I249316,I249305,);
not I_14529 (I249894,I2866);
DFFARX1 I_14530 (I62622,I2859,I249894,I249920,);
not I_14531 (I249928,I249920);
DFFARX1 I_14532 (I62607,I2859,I249894,I249954,);
not I_14533 (I249962,I62625);
nand I_14534 (I249979,I249962,I62610);
not I_14535 (I249996,I249979);
nor I_14536 (I250013,I249996,I62607);
nor I_14537 (I250030,I249928,I250013);
DFFARX1 I_14538 (I250030,I2859,I249894,I249880,);
not I_14539 (I250061,I62607);
nand I_14540 (I250078,I250061,I249996);
and I_14541 (I250095,I250061,I62610);
nand I_14542 (I250112,I250095,I62631);
nor I_14543 (I249877,I250112,I250061);
and I_14544 (I249868,I249954,I250112);
not I_14545 (I250157,I250112);
nand I_14546 (I249871,I249954,I250157);
nor I_14547 (I249865,I249920,I250112);
not I_14548 (I250202,I62619);
nor I_14549 (I250219,I250202,I62610);
nand I_14550 (I250236,I250219,I250061);
nor I_14551 (I249874,I249979,I250236);
nor I_14552 (I250267,I250202,I62613);
and I_14553 (I250284,I250267,I62628);
or I_14554 (I250301,I250284,I62616);
DFFARX1 I_14555 (I250301,I2859,I249894,I250327,);
nor I_14556 (I250335,I250327,I250078);
DFFARX1 I_14557 (I250335,I2859,I249894,I249862,);
DFFARX1 I_14558 (I250327,I2859,I249894,I249886,);
not I_14559 (I250380,I250327);
nor I_14560 (I250397,I250380,I249954);
nor I_14561 (I250414,I250219,I250397);
DFFARX1 I_14562 (I250414,I2859,I249894,I249883,);
not I_14563 (I250472,I2866);
DFFARX1 I_14564 (I533864,I2859,I250472,I250498,);
not I_14565 (I250506,I250498);
DFFARX1 I_14566 (I533882,I2859,I250472,I250532,);
not I_14567 (I250540,I533879);
nand I_14568 (I250557,I250540,I533870);
not I_14569 (I250574,I250557);
nor I_14570 (I250591,I250574,I533867);
nor I_14571 (I250608,I250506,I250591);
DFFARX1 I_14572 (I250608,I2859,I250472,I250458,);
not I_14573 (I250639,I533867);
nand I_14574 (I250656,I250639,I250574);
and I_14575 (I250673,I250639,I533873);
nand I_14576 (I250690,I250673,I533888);
nor I_14577 (I250455,I250690,I250639);
and I_14578 (I250446,I250532,I250690);
not I_14579 (I250735,I250690);
nand I_14580 (I250449,I250532,I250735);
nor I_14581 (I250443,I250498,I250690);
not I_14582 (I250780,I533864);
nor I_14583 (I250797,I250780,I533873);
nand I_14584 (I250814,I250797,I250639);
nor I_14585 (I250452,I250557,I250814);
nor I_14586 (I250845,I250780,I533885);
and I_14587 (I250862,I250845,I533876);
or I_14588 (I250879,I250862,I533891);
DFFARX1 I_14589 (I250879,I2859,I250472,I250905,);
nor I_14590 (I250913,I250905,I250656);
DFFARX1 I_14591 (I250913,I2859,I250472,I250440,);
DFFARX1 I_14592 (I250905,I2859,I250472,I250464,);
not I_14593 (I250958,I250905);
nor I_14594 (I250975,I250958,I250532);
nor I_14595 (I250992,I250797,I250975);
DFFARX1 I_14596 (I250992,I2859,I250472,I250461,);
not I_14597 (I251050,I2866);
DFFARX1 I_14598 (I128267,I2859,I251050,I251076,);
not I_14599 (I251084,I251076);
DFFARX1 I_14600 (I128282,I2859,I251050,I251110,);
not I_14601 (I251118,I128285);
nand I_14602 (I251135,I251118,I128264);
not I_14603 (I251152,I251135);
nor I_14604 (I251169,I251152,I128288);
nor I_14605 (I251186,I251084,I251169);
DFFARX1 I_14606 (I251186,I2859,I251050,I251036,);
not I_14607 (I251217,I128288);
nand I_14608 (I251234,I251217,I251152);
and I_14609 (I251251,I251217,I128270);
nand I_14610 (I251268,I251251,I128261);
nor I_14611 (I251033,I251268,I251217);
and I_14612 (I251024,I251110,I251268);
not I_14613 (I251313,I251268);
nand I_14614 (I251027,I251110,I251313);
nor I_14615 (I251021,I251076,I251268);
not I_14616 (I251358,I128261);
nor I_14617 (I251375,I251358,I128270);
nand I_14618 (I251392,I251375,I251217);
nor I_14619 (I251030,I251135,I251392);
nor I_14620 (I251423,I251358,I128276);
and I_14621 (I251440,I251423,I128279);
or I_14622 (I251457,I251440,I128273);
DFFARX1 I_14623 (I251457,I2859,I251050,I251483,);
nor I_14624 (I251491,I251483,I251234);
DFFARX1 I_14625 (I251491,I2859,I251050,I251018,);
DFFARX1 I_14626 (I251483,I2859,I251050,I251042,);
not I_14627 (I251536,I251483);
nor I_14628 (I251553,I251536,I251110);
nor I_14629 (I251570,I251375,I251553);
DFFARX1 I_14630 (I251570,I2859,I251050,I251039,);
not I_14631 (I251628,I2866);
DFFARX1 I_14632 (I302460,I2859,I251628,I251654,);
not I_14633 (I251662,I251654);
DFFARX1 I_14634 (I302472,I2859,I251628,I251688,);
not I_14635 (I251696,I302463);
nand I_14636 (I251713,I251696,I302466);
not I_14637 (I251730,I251713);
nor I_14638 (I251747,I251730,I302469);
nor I_14639 (I251764,I251662,I251747);
DFFARX1 I_14640 (I251764,I2859,I251628,I251614,);
not I_14641 (I251795,I302469);
nand I_14642 (I251812,I251795,I251730);
and I_14643 (I251829,I251795,I302463);
nand I_14644 (I251846,I251829,I302475);
nor I_14645 (I251611,I251846,I251795);
and I_14646 (I251602,I251688,I251846);
not I_14647 (I251891,I251846);
nand I_14648 (I251605,I251688,I251891);
nor I_14649 (I251599,I251654,I251846);
not I_14650 (I251936,I302481);
nor I_14651 (I251953,I251936,I302463);
nand I_14652 (I251970,I251953,I251795);
nor I_14653 (I251608,I251713,I251970);
nor I_14654 (I252001,I251936,I302460);
and I_14655 (I252018,I252001,I302478);
or I_14656 (I252035,I252018,I302484);
DFFARX1 I_14657 (I252035,I2859,I251628,I252061,);
nor I_14658 (I252069,I252061,I251812);
DFFARX1 I_14659 (I252069,I2859,I251628,I251596,);
DFFARX1 I_14660 (I252061,I2859,I251628,I251620,);
not I_14661 (I252114,I252061);
nor I_14662 (I252131,I252114,I251688);
nor I_14663 (I252148,I251953,I252131);
DFFARX1 I_14664 (I252148,I2859,I251628,I251617,);
not I_14665 (I252206,I2866);
DFFARX1 I_14666 (I552870,I2859,I252206,I252232,);
not I_14667 (I252240,I252232);
DFFARX1 I_14668 (I552870,I2859,I252206,I252266,);
not I_14669 (I252274,I552894);
nand I_14670 (I252291,I252274,I552876);
not I_14671 (I252308,I252291);
nor I_14672 (I252325,I252308,I552891);
nor I_14673 (I252342,I252240,I252325);
DFFARX1 I_14674 (I252342,I2859,I252206,I252192,);
not I_14675 (I252373,I552891);
nand I_14676 (I252390,I252373,I252308);
and I_14677 (I252407,I252373,I552873);
nand I_14678 (I252424,I252407,I552882);
nor I_14679 (I252189,I252424,I252373);
and I_14680 (I252180,I252266,I252424);
not I_14681 (I252469,I252424);
nand I_14682 (I252183,I252266,I252469);
nor I_14683 (I252177,I252232,I252424);
not I_14684 (I252514,I552879);
nor I_14685 (I252531,I252514,I552873);
nand I_14686 (I252548,I252531,I252373);
nor I_14687 (I252186,I252291,I252548);
nor I_14688 (I252579,I252514,I552888);
and I_14689 (I252596,I252579,I552897);
or I_14690 (I252613,I252596,I552885);
DFFARX1 I_14691 (I252613,I2859,I252206,I252639,);
nor I_14692 (I252647,I252639,I252390);
DFFARX1 I_14693 (I252647,I2859,I252206,I252174,);
DFFARX1 I_14694 (I252639,I2859,I252206,I252198,);
not I_14695 (I252692,I252639);
nor I_14696 (I252709,I252692,I252266);
nor I_14697 (I252726,I252531,I252709);
DFFARX1 I_14698 (I252726,I2859,I252206,I252195,);
not I_14699 (I252784,I2866);
DFFARX1 I_14700 (I431630,I2859,I252784,I252810,);
not I_14701 (I252818,I252810);
DFFARX1 I_14702 (I431621,I2859,I252784,I252844,);
not I_14703 (I252852,I431615);
nand I_14704 (I252869,I252852,I431627);
not I_14705 (I252886,I252869);
nor I_14706 (I252903,I252886,I431618);
nor I_14707 (I252920,I252818,I252903);
DFFARX1 I_14708 (I252920,I2859,I252784,I252770,);
not I_14709 (I252951,I431618);
nand I_14710 (I252968,I252951,I252886);
and I_14711 (I252985,I252951,I431624);
nand I_14712 (I253002,I252985,I431609);
nor I_14713 (I252767,I253002,I252951);
and I_14714 (I252758,I252844,I253002);
not I_14715 (I253047,I253002);
nand I_14716 (I252761,I252844,I253047);
nor I_14717 (I252755,I252810,I253002);
not I_14718 (I253092,I431609);
nor I_14719 (I253109,I253092,I431624);
nand I_14720 (I253126,I253109,I252951);
nor I_14721 (I252764,I252869,I253126);
nor I_14722 (I253157,I253092,I431612);
and I_14723 (I253174,I253157,I431615);
or I_14724 (I253191,I253174,I431612);
DFFARX1 I_14725 (I253191,I2859,I252784,I253217,);
nor I_14726 (I253225,I253217,I252968);
DFFARX1 I_14727 (I253225,I2859,I252784,I252752,);
DFFARX1 I_14728 (I253217,I2859,I252784,I252776,);
not I_14729 (I253270,I253217);
nor I_14730 (I253287,I253270,I252844);
nor I_14731 (I253304,I253109,I253287);
DFFARX1 I_14732 (I253304,I2859,I252784,I252773,);
not I_14733 (I253362,I2866);
DFFARX1 I_14734 (I1668,I2859,I253362,I253388,);
not I_14735 (I253396,I253388);
DFFARX1 I_14736 (I1748,I2859,I253362,I253422,);
not I_14737 (I253430,I1628);
nand I_14738 (I253447,I253430,I1420);
not I_14739 (I253464,I253447);
nor I_14740 (I253481,I253464,I2044);
nor I_14741 (I253498,I253396,I253481);
DFFARX1 I_14742 (I253498,I2859,I253362,I253348,);
not I_14743 (I253529,I2044);
nand I_14744 (I253546,I253529,I253464);
and I_14745 (I253563,I253529,I2020);
nand I_14746 (I253580,I253563,I1692);
nor I_14747 (I253345,I253580,I253529);
and I_14748 (I253336,I253422,I253580);
not I_14749 (I253625,I253580);
nand I_14750 (I253339,I253422,I253625);
nor I_14751 (I253333,I253388,I253580);
not I_14752 (I253670,I2588);
nor I_14753 (I253687,I253670,I2020);
nand I_14754 (I253704,I253687,I253529);
nor I_14755 (I253342,I253447,I253704);
nor I_14756 (I253735,I253670,I1804);
and I_14757 (I253752,I253735,I1724);
or I_14758 (I253769,I253752,I1564);
DFFARX1 I_14759 (I253769,I2859,I253362,I253795,);
nor I_14760 (I253803,I253795,I253546);
DFFARX1 I_14761 (I253803,I2859,I253362,I253330,);
DFFARX1 I_14762 (I253795,I2859,I253362,I253354,);
not I_14763 (I253848,I253795);
nor I_14764 (I253865,I253848,I253422);
nor I_14765 (I253882,I253687,I253865);
DFFARX1 I_14766 (I253882,I2859,I253362,I253351,);
not I_14767 (I253940,I2866);
DFFARX1 I_14768 (I267202,I2859,I253940,I253966,);
not I_14769 (I253974,I253966);
DFFARX1 I_14770 (I267214,I2859,I253940,I254000,);
not I_14771 (I254008,I267205);
nand I_14772 (I254025,I254008,I267208);
not I_14773 (I254042,I254025);
nor I_14774 (I254059,I254042,I267211);
nor I_14775 (I254076,I253974,I254059);
DFFARX1 I_14776 (I254076,I2859,I253940,I253926,);
not I_14777 (I254107,I267211);
nand I_14778 (I254124,I254107,I254042);
and I_14779 (I254141,I254107,I267205);
nand I_14780 (I254158,I254141,I267217);
nor I_14781 (I253923,I254158,I254107);
and I_14782 (I253914,I254000,I254158);
not I_14783 (I254203,I254158);
nand I_14784 (I253917,I254000,I254203);
nor I_14785 (I253911,I253966,I254158);
not I_14786 (I254248,I267223);
nor I_14787 (I254265,I254248,I267205);
nand I_14788 (I254282,I254265,I254107);
nor I_14789 (I253920,I254025,I254282);
nor I_14790 (I254313,I254248,I267202);
and I_14791 (I254330,I254313,I267220);
or I_14792 (I254347,I254330,I267226);
DFFARX1 I_14793 (I254347,I2859,I253940,I254373,);
nor I_14794 (I254381,I254373,I254124);
DFFARX1 I_14795 (I254381,I2859,I253940,I253908,);
DFFARX1 I_14796 (I254373,I2859,I253940,I253932,);
not I_14797 (I254426,I254373);
nor I_14798 (I254443,I254426,I254000);
nor I_14799 (I254460,I254265,I254443);
DFFARX1 I_14800 (I254460,I2859,I253940,I253929,);
not I_14801 (I254518,I2866);
DFFARX1 I_14802 (I405095,I2859,I254518,I254544,);
not I_14803 (I254552,I254544);
DFFARX1 I_14804 (I405092,I2859,I254518,I254578,);
not I_14805 (I254586,I405089);
nand I_14806 (I254603,I254586,I405116);
not I_14807 (I254620,I254603);
nor I_14808 (I254637,I254620,I405104);
nor I_14809 (I254654,I254552,I254637);
DFFARX1 I_14810 (I254654,I2859,I254518,I254504,);
not I_14811 (I254685,I405104);
nand I_14812 (I254702,I254685,I254620);
and I_14813 (I254719,I254685,I405110);
nand I_14814 (I254736,I254719,I405101);
nor I_14815 (I254501,I254736,I254685);
and I_14816 (I254492,I254578,I254736);
not I_14817 (I254781,I254736);
nand I_14818 (I254495,I254578,I254781);
nor I_14819 (I254489,I254544,I254736);
not I_14820 (I254826,I405098);
nor I_14821 (I254843,I254826,I405110);
nand I_14822 (I254860,I254843,I254685);
nor I_14823 (I254498,I254603,I254860);
nor I_14824 (I254891,I254826,I405113);
and I_14825 (I254908,I254891,I405107);
or I_14826 (I254925,I254908,I405089);
DFFARX1 I_14827 (I254925,I2859,I254518,I254951,);
nor I_14828 (I254959,I254951,I254702);
DFFARX1 I_14829 (I254959,I2859,I254518,I254486,);
DFFARX1 I_14830 (I254951,I2859,I254518,I254510,);
not I_14831 (I255004,I254951);
nor I_14832 (I255021,I255004,I254578);
nor I_14833 (I255038,I254843,I255021);
DFFARX1 I_14834 (I255038,I2859,I254518,I254507,);
not I_14835 (I255096,I2866);
DFFARX1 I_14836 (I427142,I2859,I255096,I255122,);
not I_14837 (I255130,I255122);
DFFARX1 I_14838 (I427133,I2859,I255096,I255156,);
not I_14839 (I255164,I427127);
nand I_14840 (I255181,I255164,I427139);
not I_14841 (I255198,I255181);
nor I_14842 (I255215,I255198,I427130);
nor I_14843 (I255232,I255130,I255215);
DFFARX1 I_14844 (I255232,I2859,I255096,I255082,);
not I_14845 (I255263,I427130);
nand I_14846 (I255280,I255263,I255198);
and I_14847 (I255297,I255263,I427136);
nand I_14848 (I255314,I255297,I427121);
nor I_14849 (I255079,I255314,I255263);
and I_14850 (I255070,I255156,I255314);
not I_14851 (I255359,I255314);
nand I_14852 (I255073,I255156,I255359);
nor I_14853 (I255067,I255122,I255314);
not I_14854 (I255404,I427121);
nor I_14855 (I255421,I255404,I427136);
nand I_14856 (I255438,I255421,I255263);
nor I_14857 (I255076,I255181,I255438);
nor I_14858 (I255469,I255404,I427124);
and I_14859 (I255486,I255469,I427127);
or I_14860 (I255503,I255486,I427124);
DFFARX1 I_14861 (I255503,I2859,I255096,I255529,);
nor I_14862 (I255537,I255529,I255280);
DFFARX1 I_14863 (I255537,I2859,I255096,I255064,);
DFFARX1 I_14864 (I255529,I2859,I255096,I255088,);
not I_14865 (I255582,I255529);
nor I_14866 (I255599,I255582,I255156);
nor I_14867 (I255616,I255421,I255599);
DFFARX1 I_14868 (I255616,I2859,I255096,I255085,);
not I_14869 (I255674,I2866);
DFFARX1 I_14870 (I279340,I2859,I255674,I255700,);
not I_14871 (I255708,I255700);
DFFARX1 I_14872 (I279352,I2859,I255674,I255734,);
not I_14873 (I255742,I279343);
nand I_14874 (I255759,I255742,I279346);
not I_14875 (I255776,I255759);
nor I_14876 (I255793,I255776,I279349);
nor I_14877 (I255810,I255708,I255793);
DFFARX1 I_14878 (I255810,I2859,I255674,I255660,);
not I_14879 (I255841,I279349);
nand I_14880 (I255858,I255841,I255776);
and I_14881 (I255875,I255841,I279343);
nand I_14882 (I255892,I255875,I279355);
nor I_14883 (I255657,I255892,I255841);
and I_14884 (I255648,I255734,I255892);
not I_14885 (I255937,I255892);
nand I_14886 (I255651,I255734,I255937);
nor I_14887 (I255645,I255700,I255892);
not I_14888 (I255982,I279361);
nor I_14889 (I255999,I255982,I279343);
nand I_14890 (I256016,I255999,I255841);
nor I_14891 (I255654,I255759,I256016);
nor I_14892 (I256047,I255982,I279340);
and I_14893 (I256064,I256047,I279358);
or I_14894 (I256081,I256064,I279364);
DFFARX1 I_14895 (I256081,I2859,I255674,I256107,);
nor I_14896 (I256115,I256107,I255858);
DFFARX1 I_14897 (I256115,I2859,I255674,I255642,);
DFFARX1 I_14898 (I256107,I2859,I255674,I255666,);
not I_14899 (I256160,I256107);
nor I_14900 (I256177,I256160,I255734);
nor I_14901 (I256194,I255999,I256177);
DFFARX1 I_14902 (I256194,I2859,I255674,I255663,);
not I_14903 (I256252,I2866);
DFFARX1 I_14904 (I95942,I2859,I256252,I256278,);
not I_14905 (I256286,I256278);
DFFARX1 I_14906 (I95927,I2859,I256252,I256312,);
not I_14907 (I256320,I95945);
nand I_14908 (I256337,I256320,I95930);
not I_14909 (I256354,I256337);
nor I_14910 (I256371,I256354,I95927);
nor I_14911 (I256388,I256286,I256371);
DFFARX1 I_14912 (I256388,I2859,I256252,I256238,);
not I_14913 (I256419,I95927);
nand I_14914 (I256436,I256419,I256354);
and I_14915 (I256453,I256419,I95930);
nand I_14916 (I256470,I256453,I95951);
nor I_14917 (I256235,I256470,I256419);
and I_14918 (I256226,I256312,I256470);
not I_14919 (I256515,I256470);
nand I_14920 (I256229,I256312,I256515);
nor I_14921 (I256223,I256278,I256470);
not I_14922 (I256560,I95939);
nor I_14923 (I256577,I256560,I95930);
nand I_14924 (I256594,I256577,I256419);
nor I_14925 (I256232,I256337,I256594);
nor I_14926 (I256625,I256560,I95933);
and I_14927 (I256642,I256625,I95948);
or I_14928 (I256659,I256642,I95936);
DFFARX1 I_14929 (I256659,I2859,I256252,I256685,);
nor I_14930 (I256693,I256685,I256436);
DFFARX1 I_14931 (I256693,I2859,I256252,I256220,);
DFFARX1 I_14932 (I256685,I2859,I256252,I256244,);
not I_14933 (I256738,I256685);
nor I_14934 (I256755,I256738,I256312);
nor I_14935 (I256772,I256577,I256755);
DFFARX1 I_14936 (I256772,I2859,I256252,I256241,);
not I_14937 (I256830,I2866);
DFFARX1 I_14938 (I410909,I2859,I256830,I256856,);
not I_14939 (I256864,I256856);
DFFARX1 I_14940 (I410906,I2859,I256830,I256890,);
not I_14941 (I256898,I410903);
nand I_14942 (I256915,I256898,I410930);
not I_14943 (I256932,I256915);
nor I_14944 (I256949,I256932,I410918);
nor I_14945 (I256966,I256864,I256949);
DFFARX1 I_14946 (I256966,I2859,I256830,I256816,);
not I_14947 (I256997,I410918);
nand I_14948 (I257014,I256997,I256932);
and I_14949 (I257031,I256997,I410924);
nand I_14950 (I257048,I257031,I410915);
nor I_14951 (I256813,I257048,I256997);
and I_14952 (I256804,I256890,I257048);
not I_14953 (I257093,I257048);
nand I_14954 (I256807,I256890,I257093);
nor I_14955 (I256801,I256856,I257048);
not I_14956 (I257138,I410912);
nor I_14957 (I257155,I257138,I410924);
nand I_14958 (I257172,I257155,I256997);
nor I_14959 (I256810,I256915,I257172);
nor I_14960 (I257203,I257138,I410927);
and I_14961 (I257220,I257203,I410921);
or I_14962 (I257237,I257220,I410903);
DFFARX1 I_14963 (I257237,I2859,I256830,I257263,);
nor I_14964 (I257271,I257263,I257014);
DFFARX1 I_14965 (I257271,I2859,I256830,I256798,);
DFFARX1 I_14966 (I257263,I2859,I256830,I256822,);
not I_14967 (I257316,I257263);
nor I_14968 (I257333,I257316,I256890);
nor I_14969 (I257350,I257155,I257333);
DFFARX1 I_14970 (I257350,I2859,I256830,I256819,);
not I_14971 (I257408,I2866);
DFFARX1 I_14972 (I518904,I2859,I257408,I257434,);
not I_14973 (I257442,I257434);
nand I_14974 (I257459,I518928,I518910);
and I_14975 (I257476,I257459,I518916);
DFFARX1 I_14976 (I257476,I2859,I257408,I257502,);
not I_14977 (I257510,I518922);
DFFARX1 I_14978 (I518907,I2859,I257408,I257536,);
not I_14979 (I257544,I257536);
nor I_14980 (I257561,I257544,I257442);
and I_14981 (I257578,I257561,I518922);
nor I_14982 (I257595,I257544,I257510);
nor I_14983 (I257391,I257502,I257595);
DFFARX1 I_14984 (I518919,I2859,I257408,I257635,);
nor I_14985 (I257643,I257635,I257502);
not I_14986 (I257660,I257643);
not I_14987 (I257677,I257635);
nor I_14988 (I257694,I257677,I257578);
DFFARX1 I_14989 (I257694,I2859,I257408,I257394,);
nand I_14990 (I257725,I518925,I518913);
and I_14991 (I257742,I257725,I518907);
DFFARX1 I_14992 (I257742,I2859,I257408,I257768,);
nor I_14993 (I257776,I257768,I257635);
DFFARX1 I_14994 (I257776,I2859,I257408,I257376,);
nand I_14995 (I257807,I257768,I257677);
nand I_14996 (I257385,I257660,I257807);
not I_14997 (I257838,I257768);
nor I_14998 (I257855,I257838,I257578);
DFFARX1 I_14999 (I257855,I2859,I257408,I257397,);
nor I_15000 (I257886,I518904,I518913);
or I_15001 (I257388,I257635,I257886);
nor I_15002 (I257379,I257768,I257886);
or I_15003 (I257382,I257502,I257886);
DFFARX1 I_15004 (I257886,I2859,I257408,I257400,);
not I_15005 (I257986,I2866);
DFFARX1 I_15006 (I543972,I2859,I257986,I258012,);
not I_15007 (I258020,I258012);
nand I_15008 (I258037,I543957,I543945);
and I_15009 (I258054,I258037,I543960);
DFFARX1 I_15010 (I258054,I2859,I257986,I258080,);
not I_15011 (I258088,I543945);
DFFARX1 I_15012 (I543963,I2859,I257986,I258114,);
not I_15013 (I258122,I258114);
nor I_15014 (I258139,I258122,I258020);
and I_15015 (I258156,I258139,I543945);
nor I_15016 (I258173,I258122,I258088);
nor I_15017 (I257969,I258080,I258173);
DFFARX1 I_15018 (I543951,I2859,I257986,I258213,);
nor I_15019 (I258221,I258213,I258080);
not I_15020 (I258238,I258221);
not I_15021 (I258255,I258213);
nor I_15022 (I258272,I258255,I258156);
DFFARX1 I_15023 (I258272,I2859,I257986,I257972,);
nand I_15024 (I258303,I543948,I543954);
and I_15025 (I258320,I258303,I543969);
DFFARX1 I_15026 (I258320,I2859,I257986,I258346,);
nor I_15027 (I258354,I258346,I258213);
DFFARX1 I_15028 (I258354,I2859,I257986,I257954,);
nand I_15029 (I258385,I258346,I258255);
nand I_15030 (I257963,I258238,I258385);
not I_15031 (I258416,I258346);
nor I_15032 (I258433,I258416,I258156);
DFFARX1 I_15033 (I258433,I2859,I257986,I257975,);
nor I_15034 (I258464,I543966,I543954);
or I_15035 (I257966,I258213,I258464);
nor I_15036 (I257957,I258346,I258464);
or I_15037 (I257960,I258080,I258464);
DFFARX1 I_15038 (I258464,I2859,I257986,I257978,);
not I_15039 (I258564,I2866);
DFFARX1 I_15040 (I105447,I2859,I258564,I258590,);
not I_15041 (I258598,I258590);
nand I_15042 (I258615,I105450,I105471);
and I_15043 (I258632,I258615,I105459);
DFFARX1 I_15044 (I258632,I2859,I258564,I258658,);
not I_15045 (I258666,I105456);
DFFARX1 I_15046 (I105447,I2859,I258564,I258692,);
not I_15047 (I258700,I258692);
nor I_15048 (I258717,I258700,I258598);
and I_15049 (I258734,I258717,I105456);
nor I_15050 (I258751,I258700,I258666);
nor I_15051 (I258547,I258658,I258751);
DFFARX1 I_15052 (I105465,I2859,I258564,I258791,);
nor I_15053 (I258799,I258791,I258658);
not I_15054 (I258816,I258799);
not I_15055 (I258833,I258791);
nor I_15056 (I258850,I258833,I258734);
DFFARX1 I_15057 (I258850,I2859,I258564,I258550,);
nand I_15058 (I258881,I105450,I105453);
and I_15059 (I258898,I258881,I105462);
DFFARX1 I_15060 (I258898,I2859,I258564,I258924,);
nor I_15061 (I258932,I258924,I258791);
DFFARX1 I_15062 (I258932,I2859,I258564,I258532,);
nand I_15063 (I258963,I258924,I258833);
nand I_15064 (I258541,I258816,I258963);
not I_15065 (I258994,I258924);
nor I_15066 (I259011,I258994,I258734);
DFFARX1 I_15067 (I259011,I2859,I258564,I258553,);
nor I_15068 (I259042,I105468,I105453);
or I_15069 (I258544,I258791,I259042);
nor I_15070 (I258535,I258924,I259042);
or I_15071 (I258538,I258658,I259042);
DFFARX1 I_15072 (I259042,I2859,I258564,I258556,);
not I_15073 (I259142,I2866);
DFFARX1 I_15074 (I410281,I2859,I259142,I259168,);
not I_15075 (I259176,I259168);
nand I_15076 (I259193,I410257,I410272);
and I_15077 (I259210,I259193,I410284);
DFFARX1 I_15078 (I259210,I2859,I259142,I259236,);
not I_15079 (I259244,I410269);
DFFARX1 I_15080 (I410260,I2859,I259142,I259270,);
not I_15081 (I259278,I259270);
nor I_15082 (I259295,I259278,I259176);
and I_15083 (I259312,I259295,I410269);
nor I_15084 (I259329,I259278,I259244);
nor I_15085 (I259125,I259236,I259329);
DFFARX1 I_15086 (I410257,I2859,I259142,I259369,);
nor I_15087 (I259377,I259369,I259236);
not I_15088 (I259394,I259377);
not I_15089 (I259411,I259369);
nor I_15090 (I259428,I259411,I259312);
DFFARX1 I_15091 (I259428,I2859,I259142,I259128,);
nand I_15092 (I259459,I410275,I410266);
and I_15093 (I259476,I259459,I410278);
DFFARX1 I_15094 (I259476,I2859,I259142,I259502,);
nor I_15095 (I259510,I259502,I259369);
DFFARX1 I_15096 (I259510,I2859,I259142,I259110,);
nand I_15097 (I259541,I259502,I259411);
nand I_15098 (I259119,I259394,I259541);
not I_15099 (I259572,I259502);
nor I_15100 (I259589,I259572,I259312);
DFFARX1 I_15101 (I259589,I2859,I259142,I259131,);
nor I_15102 (I259620,I410263,I410266);
or I_15103 (I259122,I259369,I259620);
nor I_15104 (I259113,I259502,I259620);
or I_15105 (I259116,I259236,I259620);
DFFARX1 I_15106 (I259620,I2859,I259142,I259134,);
not I_15107 (I259720,I2866);
DFFARX1 I_15108 (I431054,I2859,I259720,I259746,);
not I_15109 (I259754,I259746);
nand I_15110 (I259771,I431051,I431069);
and I_15111 (I259788,I259771,I431066);
DFFARX1 I_15112 (I259788,I2859,I259720,I259814,);
not I_15113 (I259822,I431048);
DFFARX1 I_15114 (I431051,I2859,I259720,I259848,);
not I_15115 (I259856,I259848);
nor I_15116 (I259873,I259856,I259754);
and I_15117 (I259890,I259873,I431048);
nor I_15118 (I259907,I259856,I259822);
nor I_15119 (I259703,I259814,I259907);
DFFARX1 I_15120 (I431060,I2859,I259720,I259947,);
nor I_15121 (I259955,I259947,I259814);
not I_15122 (I259972,I259955);
not I_15123 (I259989,I259947);
nor I_15124 (I260006,I259989,I259890);
DFFARX1 I_15125 (I260006,I2859,I259720,I259706,);
nand I_15126 (I260037,I431063,I431048);
and I_15127 (I260054,I260037,I431054);
DFFARX1 I_15128 (I260054,I2859,I259720,I260080,);
nor I_15129 (I260088,I260080,I259947);
DFFARX1 I_15130 (I260088,I2859,I259720,I259688,);
nand I_15131 (I260119,I260080,I259989);
nand I_15132 (I259697,I259972,I260119);
not I_15133 (I260150,I260080);
nor I_15134 (I260167,I260150,I259890);
DFFARX1 I_15135 (I260167,I2859,I259720,I259709,);
nor I_15136 (I260198,I431057,I431048);
or I_15137 (I259700,I259947,I260198);
nor I_15138 (I259691,I260080,I260198);
or I_15139 (I259694,I259814,I260198);
DFFARX1 I_15140 (I260198,I2859,I259720,I259712,);
not I_15141 (I260298,I2866);
DFFARX1 I_15142 (I115637,I2859,I260298,I260324,);
not I_15143 (I260332,I260324);
nand I_15144 (I260349,I115640,I115616);
and I_15145 (I260366,I260349,I115613);
DFFARX1 I_15146 (I260366,I2859,I260298,I260392,);
not I_15147 (I260400,I115619);
DFFARX1 I_15148 (I115613,I2859,I260298,I260426,);
not I_15149 (I260434,I260426);
nor I_15150 (I260451,I260434,I260332);
and I_15151 (I260468,I260451,I115619);
nor I_15152 (I260485,I260434,I260400);
nor I_15153 (I260281,I260392,I260485);
DFFARX1 I_15154 (I115622,I2859,I260298,I260525,);
nor I_15155 (I260533,I260525,I260392);
not I_15156 (I260550,I260533);
not I_15157 (I260567,I260525);
nor I_15158 (I260584,I260567,I260468);
DFFARX1 I_15159 (I260584,I2859,I260298,I260284,);
nand I_15160 (I260615,I115625,I115634);
and I_15161 (I260632,I260615,I115631);
DFFARX1 I_15162 (I260632,I2859,I260298,I260658,);
nor I_15163 (I260666,I260658,I260525);
DFFARX1 I_15164 (I260666,I2859,I260298,I260266,);
nand I_15165 (I260697,I260658,I260567);
nand I_15166 (I260275,I260550,I260697);
not I_15167 (I260728,I260658);
nor I_15168 (I260745,I260728,I260468);
DFFARX1 I_15169 (I260745,I2859,I260298,I260287,);
nor I_15170 (I260776,I115628,I115634);
or I_15171 (I260278,I260525,I260776);
nor I_15172 (I260269,I260658,I260776);
or I_15173 (I260272,I260392,I260776);
DFFARX1 I_15174 (I260776,I2859,I260298,I260290,);
not I_15175 (I260876,I2866);
DFFARX1 I_15176 (I199585,I2859,I260876,I260902,);
not I_15177 (I260910,I260902);
nand I_15178 (I260927,I199576,I199594);
and I_15179 (I260944,I260927,I199597);
DFFARX1 I_15180 (I260944,I2859,I260876,I260970,);
not I_15181 (I260978,I199591);
DFFARX1 I_15182 (I199579,I2859,I260876,I261004,);
not I_15183 (I261012,I261004);
nor I_15184 (I261029,I261012,I260910);
and I_15185 (I261046,I261029,I199591);
nor I_15186 (I261063,I261012,I260978);
nor I_15187 (I260859,I260970,I261063);
DFFARX1 I_15188 (I199588,I2859,I260876,I261103,);
nor I_15189 (I261111,I261103,I260970);
not I_15190 (I261128,I261111);
not I_15191 (I261145,I261103);
nor I_15192 (I261162,I261145,I261046);
DFFARX1 I_15193 (I261162,I2859,I260876,I260862,);
nand I_15194 (I261193,I199603,I199600);
and I_15195 (I261210,I261193,I199582);
DFFARX1 I_15196 (I261210,I2859,I260876,I261236,);
nor I_15197 (I261244,I261236,I261103);
DFFARX1 I_15198 (I261244,I2859,I260876,I260844,);
nand I_15199 (I261275,I261236,I261145);
nand I_15200 (I260853,I261128,I261275);
not I_15201 (I261306,I261236);
nor I_15202 (I261323,I261306,I261046);
DFFARX1 I_15203 (I261323,I2859,I260876,I260865,);
nor I_15204 (I261354,I199576,I199600);
or I_15205 (I260856,I261103,I261354);
nor I_15206 (I260847,I261236,I261354);
or I_15207 (I260850,I260970,I261354);
DFFARX1 I_15208 (I261354,I2859,I260876,I260868,);
not I_15209 (I261454,I2866);
DFFARX1 I_15210 (I66772,I2859,I261454,I261480,);
not I_15211 (I261488,I261480);
nand I_15212 (I261505,I66775,I66796);
and I_15213 (I261522,I261505,I66784);
DFFARX1 I_15214 (I261522,I2859,I261454,I261548,);
not I_15215 (I261556,I66781);
DFFARX1 I_15216 (I66772,I2859,I261454,I261582,);
not I_15217 (I261590,I261582);
nor I_15218 (I261607,I261590,I261488);
and I_15219 (I261624,I261607,I66781);
nor I_15220 (I261641,I261590,I261556);
nor I_15221 (I261437,I261548,I261641);
DFFARX1 I_15222 (I66790,I2859,I261454,I261681,);
nor I_15223 (I261689,I261681,I261548);
not I_15224 (I261706,I261689);
not I_15225 (I261723,I261681);
nor I_15226 (I261740,I261723,I261624);
DFFARX1 I_15227 (I261740,I2859,I261454,I261440,);
nand I_15228 (I261771,I66775,I66778);
and I_15229 (I261788,I261771,I66787);
DFFARX1 I_15230 (I261788,I2859,I261454,I261814,);
nor I_15231 (I261822,I261814,I261681);
DFFARX1 I_15232 (I261822,I2859,I261454,I261422,);
nand I_15233 (I261853,I261814,I261723);
nand I_15234 (I261431,I261706,I261853);
not I_15235 (I261884,I261814);
nor I_15236 (I261901,I261884,I261624);
DFFARX1 I_15237 (I261901,I2859,I261454,I261443,);
nor I_15238 (I261932,I66793,I66778);
or I_15239 (I261434,I261681,I261932);
nor I_15240 (I261425,I261814,I261932);
or I_15241 (I261428,I261548,I261932);
DFFARX1 I_15242 (I261932,I2859,I261454,I261446,);
not I_15243 (I262032,I2866);
DFFARX1 I_15244 (I72722,I2859,I262032,I262058,);
not I_15245 (I262066,I262058);
nand I_15246 (I262083,I72725,I72746);
and I_15247 (I262100,I262083,I72734);
DFFARX1 I_15248 (I262100,I2859,I262032,I262126,);
not I_15249 (I262134,I72731);
DFFARX1 I_15250 (I72722,I2859,I262032,I262160,);
not I_15251 (I262168,I262160);
nor I_15252 (I262185,I262168,I262066);
and I_15253 (I262202,I262185,I72731);
nor I_15254 (I262219,I262168,I262134);
nor I_15255 (I262015,I262126,I262219);
DFFARX1 I_15256 (I72740,I2859,I262032,I262259,);
nor I_15257 (I262267,I262259,I262126);
not I_15258 (I262284,I262267);
not I_15259 (I262301,I262259);
nor I_15260 (I262318,I262301,I262202);
DFFARX1 I_15261 (I262318,I2859,I262032,I262018,);
nand I_15262 (I262349,I72725,I72728);
and I_15263 (I262366,I262349,I72737);
DFFARX1 I_15264 (I262366,I2859,I262032,I262392,);
nor I_15265 (I262400,I262392,I262259);
DFFARX1 I_15266 (I262400,I2859,I262032,I262000,);
nand I_15267 (I262431,I262392,I262301);
nand I_15268 (I262009,I262284,I262431);
not I_15269 (I262462,I262392);
nor I_15270 (I262479,I262462,I262202);
DFFARX1 I_15271 (I262479,I2859,I262032,I262021,);
nor I_15272 (I262510,I72743,I72728);
or I_15273 (I262012,I262259,I262510);
nor I_15274 (I262003,I262392,I262510);
or I_15275 (I262006,I262126,I262510);
DFFARX1 I_15276 (I262510,I2859,I262032,I262024,);
not I_15277 (I262610,I2866);
DFFARX1 I_15278 (I125123,I2859,I262610,I262636,);
not I_15279 (I262644,I262636);
nand I_15280 (I262661,I125126,I125102);
and I_15281 (I262678,I262661,I125099);
DFFARX1 I_15282 (I262678,I2859,I262610,I262704,);
not I_15283 (I262712,I125105);
DFFARX1 I_15284 (I125099,I2859,I262610,I262738,);
not I_15285 (I262746,I262738);
nor I_15286 (I262763,I262746,I262644);
and I_15287 (I262780,I262763,I125105);
nor I_15288 (I262797,I262746,I262712);
nor I_15289 (I262593,I262704,I262797);
DFFARX1 I_15290 (I125108,I2859,I262610,I262837,);
nor I_15291 (I262845,I262837,I262704);
not I_15292 (I262862,I262845);
not I_15293 (I262879,I262837);
nor I_15294 (I262896,I262879,I262780);
DFFARX1 I_15295 (I262896,I2859,I262610,I262596,);
nand I_15296 (I262927,I125111,I125120);
and I_15297 (I262944,I262927,I125117);
DFFARX1 I_15298 (I262944,I2859,I262610,I262970,);
nor I_15299 (I262978,I262970,I262837);
DFFARX1 I_15300 (I262978,I2859,I262610,I262578,);
nand I_15301 (I263009,I262970,I262879);
nand I_15302 (I262587,I262862,I263009);
not I_15303 (I263040,I262970);
nor I_15304 (I263057,I263040,I262780);
DFFARX1 I_15305 (I263057,I2859,I262610,I262599,);
nor I_15306 (I263088,I125114,I125120);
or I_15307 (I262590,I262837,I263088);
nor I_15308 (I262581,I262970,I263088);
or I_15309 (I262584,I262704,I263088);
DFFARX1 I_15310 (I263088,I2859,I262610,I262602,);
not I_15311 (I263188,I2866);
DFFARX1 I_15312 (I365061,I2859,I263188,I263214,);
not I_15313 (I263222,I263214);
nand I_15314 (I263239,I365037,I365052);
and I_15315 (I263256,I263239,I365064);
DFFARX1 I_15316 (I263256,I2859,I263188,I263282,);
not I_15317 (I263290,I365049);
DFFARX1 I_15318 (I365040,I2859,I263188,I263316,);
not I_15319 (I263324,I263316);
nor I_15320 (I263341,I263324,I263222);
and I_15321 (I263358,I263341,I365049);
nor I_15322 (I263375,I263324,I263290);
nor I_15323 (I263171,I263282,I263375);
DFFARX1 I_15324 (I365037,I2859,I263188,I263415,);
nor I_15325 (I263423,I263415,I263282);
not I_15326 (I263440,I263423);
not I_15327 (I263457,I263415);
nor I_15328 (I263474,I263457,I263358);
DFFARX1 I_15329 (I263474,I2859,I263188,I263174,);
nand I_15330 (I263505,I365055,I365046);
and I_15331 (I263522,I263505,I365058);
DFFARX1 I_15332 (I263522,I2859,I263188,I263548,);
nor I_15333 (I263556,I263548,I263415);
DFFARX1 I_15334 (I263556,I2859,I263188,I263156,);
nand I_15335 (I263587,I263548,I263457);
nand I_15336 (I263165,I263440,I263587);
not I_15337 (I263618,I263548);
nor I_15338 (I263635,I263618,I263358);
DFFARX1 I_15339 (I263635,I2859,I263188,I263177,);
nor I_15340 (I263666,I365043,I365046);
or I_15341 (I263168,I263415,I263666);
nor I_15342 (I263159,I263548,I263666);
or I_15343 (I263162,I263282,I263666);
DFFARX1 I_15344 (I263666,I2859,I263188,I263180,);
not I_15345 (I263766,I2866);
DFFARX1 I_15346 (I453370,I2859,I263766,I263792,);
not I_15347 (I263800,I263792);
nand I_15348 (I263817,I453352,I453364);
and I_15349 (I263834,I263817,I453367);
DFFARX1 I_15350 (I263834,I2859,I263766,I263860,);
not I_15351 (I263868,I453361);
DFFARX1 I_15352 (I453358,I2859,I263766,I263894,);
not I_15353 (I263902,I263894);
nor I_15354 (I263919,I263902,I263800);
and I_15355 (I263936,I263919,I453361);
nor I_15356 (I263953,I263902,I263868);
nor I_15357 (I263749,I263860,I263953);
DFFARX1 I_15358 (I453376,I2859,I263766,I263993,);
nor I_15359 (I264001,I263993,I263860);
not I_15360 (I264018,I264001);
not I_15361 (I264035,I263993);
nor I_15362 (I264052,I264035,I263936);
DFFARX1 I_15363 (I264052,I2859,I263766,I263752,);
nand I_15364 (I264083,I453355,I453355);
and I_15365 (I264100,I264083,I453352);
DFFARX1 I_15366 (I264100,I2859,I263766,I264126,);
nor I_15367 (I264134,I264126,I263993);
DFFARX1 I_15368 (I264134,I2859,I263766,I263734,);
nand I_15369 (I264165,I264126,I264035);
nand I_15370 (I263743,I264018,I264165);
not I_15371 (I264196,I264126);
nor I_15372 (I264213,I264196,I263936);
DFFARX1 I_15373 (I264213,I2859,I263766,I263755,);
nor I_15374 (I264244,I453373,I453355);
or I_15375 (I263746,I263993,I264244);
nor I_15376 (I263737,I264126,I264244);
or I_15377 (I263740,I263860,I264244);
DFFARX1 I_15378 (I264244,I2859,I263766,I263758,);
not I_15379 (I264344,I2866);
DFFARX1 I_15380 (I46953,I2859,I264344,I264370,);
not I_15381 (I264378,I264370);
nand I_15382 (I264395,I46962,I46971);
and I_15383 (I264412,I264395,I46950);
DFFARX1 I_15384 (I264412,I2859,I264344,I264438,);
not I_15385 (I264446,I46953);
DFFARX1 I_15386 (I46968,I2859,I264344,I264472,);
not I_15387 (I264480,I264472);
nor I_15388 (I264497,I264480,I264378);
and I_15389 (I264514,I264497,I46953);
nor I_15390 (I264531,I264480,I264446);
nor I_15391 (I264327,I264438,I264531);
DFFARX1 I_15392 (I46959,I2859,I264344,I264571,);
nor I_15393 (I264579,I264571,I264438);
not I_15394 (I264596,I264579);
not I_15395 (I264613,I264571);
nor I_15396 (I264630,I264613,I264514);
DFFARX1 I_15397 (I264630,I2859,I264344,I264330,);
nand I_15398 (I264661,I46974,I46950);
and I_15399 (I264678,I264661,I46956);
DFFARX1 I_15400 (I264678,I2859,I264344,I264704,);
nor I_15401 (I264712,I264704,I264571);
DFFARX1 I_15402 (I264712,I2859,I264344,I264312,);
nand I_15403 (I264743,I264704,I264613);
nand I_15404 (I264321,I264596,I264743);
not I_15405 (I264774,I264704);
nor I_15406 (I264791,I264774,I264514);
DFFARX1 I_15407 (I264791,I2859,I264344,I264333,);
nor I_15408 (I264822,I46965,I46950);
or I_15409 (I264324,I264571,I264822);
nor I_15410 (I264315,I264704,I264822);
or I_15411 (I264318,I264438,I264822);
DFFARX1 I_15412 (I264822,I2859,I264344,I264336,);
not I_15413 (I264922,I2866);
DFFARX1 I_15414 (I450480,I2859,I264922,I264948,);
not I_15415 (I264956,I264948);
nand I_15416 (I264973,I450462,I450474);
and I_15417 (I264990,I264973,I450477);
DFFARX1 I_15418 (I264990,I2859,I264922,I265016,);
not I_15419 (I265024,I450471);
DFFARX1 I_15420 (I450468,I2859,I264922,I265050,);
not I_15421 (I265058,I265050);
nor I_15422 (I265075,I265058,I264956);
and I_15423 (I265092,I265075,I450471);
nor I_15424 (I265109,I265058,I265024);
nor I_15425 (I264905,I265016,I265109);
DFFARX1 I_15426 (I450486,I2859,I264922,I265149,);
nor I_15427 (I265157,I265149,I265016);
not I_15428 (I265174,I265157);
not I_15429 (I265191,I265149);
nor I_15430 (I265208,I265191,I265092);
DFFARX1 I_15431 (I265208,I2859,I264922,I264908,);
nand I_15432 (I265239,I450465,I450465);
and I_15433 (I265256,I265239,I450462);
DFFARX1 I_15434 (I265256,I2859,I264922,I265282,);
nor I_15435 (I265290,I265282,I265149);
DFFARX1 I_15436 (I265290,I2859,I264922,I264890,);
nand I_15437 (I265321,I265282,I265191);
nand I_15438 (I264899,I265174,I265321);
not I_15439 (I265352,I265282);
nor I_15440 (I265369,I265352,I265092);
DFFARX1 I_15441 (I265369,I2859,I264922,I264911,);
nor I_15442 (I265400,I450483,I450465);
or I_15443 (I264902,I265149,I265400);
nor I_15444 (I264893,I265282,I265400);
or I_15445 (I264896,I265016,I265400);
DFFARX1 I_15446 (I265400,I2859,I264922,I264914,);
not I_15447 (I265500,I2866);
DFFARX1 I_15448 (I9545,I2859,I265500,I265526,);
not I_15449 (I265534,I265526);
nand I_15450 (I265551,I9542,I9533);
and I_15451 (I265568,I265551,I9533);
DFFARX1 I_15452 (I265568,I2859,I265500,I265594,);
not I_15453 (I265602,I9536);
DFFARX1 I_15454 (I9551,I2859,I265500,I265628,);
not I_15455 (I265636,I265628);
nor I_15456 (I265653,I265636,I265534);
and I_15457 (I265670,I265653,I9536);
nor I_15458 (I265687,I265636,I265602);
nor I_15459 (I265483,I265594,I265687);
DFFARX1 I_15460 (I9536,I2859,I265500,I265727,);
nor I_15461 (I265735,I265727,I265594);
not I_15462 (I265752,I265735);
not I_15463 (I265769,I265727);
nor I_15464 (I265786,I265769,I265670);
DFFARX1 I_15465 (I265786,I2859,I265500,I265486,);
nand I_15466 (I265817,I9554,I9539);
and I_15467 (I265834,I265817,I9557);
DFFARX1 I_15468 (I265834,I2859,I265500,I265860,);
nor I_15469 (I265868,I265860,I265727);
DFFARX1 I_15470 (I265868,I2859,I265500,I265468,);
nand I_15471 (I265899,I265860,I265769);
nand I_15472 (I265477,I265752,I265899);
not I_15473 (I265930,I265860);
nor I_15474 (I265947,I265930,I265670);
DFFARX1 I_15475 (I265947,I2859,I265500,I265489,);
nor I_15476 (I265978,I9548,I9539);
or I_15477 (I265480,I265727,I265978);
nor I_15478 (I265471,I265860,I265978);
or I_15479 (I265474,I265594,I265978);
DFFARX1 I_15480 (I265978,I2859,I265500,I265492,);
not I_15481 (I266078,I2866);
DFFARX1 I_15482 (I101282,I2859,I266078,I266104,);
not I_15483 (I266112,I266104);
nand I_15484 (I266129,I101285,I101306);
and I_15485 (I266146,I266129,I101294);
DFFARX1 I_15486 (I266146,I2859,I266078,I266172,);
not I_15487 (I266180,I101291);
DFFARX1 I_15488 (I101282,I2859,I266078,I266206,);
not I_15489 (I266214,I266206);
nor I_15490 (I266231,I266214,I266112);
and I_15491 (I266248,I266231,I101291);
nor I_15492 (I266265,I266214,I266180);
nor I_15493 (I266061,I266172,I266265);
DFFARX1 I_15494 (I101300,I2859,I266078,I266305,);
nor I_15495 (I266313,I266305,I266172);
not I_15496 (I266330,I266313);
not I_15497 (I266347,I266305);
nor I_15498 (I266364,I266347,I266248);
DFFARX1 I_15499 (I266364,I2859,I266078,I266064,);
nand I_15500 (I266395,I101285,I101288);
and I_15501 (I266412,I266395,I101297);
DFFARX1 I_15502 (I266412,I2859,I266078,I266438,);
nor I_15503 (I266446,I266438,I266305);
DFFARX1 I_15504 (I266446,I2859,I266078,I266046,);
nand I_15505 (I266477,I266438,I266347);
nand I_15506 (I266055,I266330,I266477);
not I_15507 (I266508,I266438);
nor I_15508 (I266525,I266508,I266248);
DFFARX1 I_15509 (I266525,I2859,I266078,I266067,);
nor I_15510 (I266556,I101303,I101288);
or I_15511 (I266058,I266305,I266556);
nor I_15512 (I266049,I266438,I266556);
or I_15513 (I266052,I266172,I266556);
DFFARX1 I_15514 (I266556,I2859,I266078,I266070,);
not I_15515 (I266656,I2866);
DFFARX1 I_15516 (I89977,I2859,I266656,I266682,);
not I_15517 (I266690,I266682);
nand I_15518 (I266707,I89980,I90001);
and I_15519 (I266724,I266707,I89989);
DFFARX1 I_15520 (I266724,I2859,I266656,I266750,);
not I_15521 (I266758,I89986);
DFFARX1 I_15522 (I89977,I2859,I266656,I266784,);
not I_15523 (I266792,I266784);
nor I_15524 (I266809,I266792,I266690);
and I_15525 (I266826,I266809,I89986);
nor I_15526 (I266843,I266792,I266758);
nor I_15527 (I266639,I266750,I266843);
DFFARX1 I_15528 (I89995,I2859,I266656,I266883,);
nor I_15529 (I266891,I266883,I266750);
not I_15530 (I266908,I266891);
not I_15531 (I266925,I266883);
nor I_15532 (I266942,I266925,I266826);
DFFARX1 I_15533 (I266942,I2859,I266656,I266642,);
nand I_15534 (I266973,I89980,I89983);
and I_15535 (I266990,I266973,I89992);
DFFARX1 I_15536 (I266990,I2859,I266656,I267016,);
nor I_15537 (I267024,I267016,I266883);
DFFARX1 I_15538 (I267024,I2859,I266656,I266624,);
nand I_15539 (I267055,I267016,I266925);
nand I_15540 (I266633,I266908,I267055);
not I_15541 (I267086,I267016);
nor I_15542 (I267103,I267086,I266826);
DFFARX1 I_15543 (I267103,I2859,I266656,I266645,);
nor I_15544 (I267134,I89998,I89983);
or I_15545 (I266636,I266883,I267134);
nor I_15546 (I266627,I267016,I267134);
or I_15547 (I266630,I266750,I267134);
DFFARX1 I_15548 (I267134,I2859,I266656,I266648,);
not I_15549 (I267234,I2866);
DFFARX1 I_15550 (I388963,I2859,I267234,I267260,);
not I_15551 (I267268,I267260);
nand I_15552 (I267285,I388939,I388954);
and I_15553 (I267302,I267285,I388966);
DFFARX1 I_15554 (I267302,I2859,I267234,I267328,);
not I_15555 (I267336,I388951);
DFFARX1 I_15556 (I388942,I2859,I267234,I267362,);
not I_15557 (I267370,I267362);
nor I_15558 (I267387,I267370,I267268);
and I_15559 (I267404,I267387,I388951);
nor I_15560 (I267421,I267370,I267336);
nor I_15561 (I267217,I267328,I267421);
DFFARX1 I_15562 (I388939,I2859,I267234,I267461,);
nor I_15563 (I267469,I267461,I267328);
not I_15564 (I267486,I267469);
not I_15565 (I267503,I267461);
nor I_15566 (I267520,I267503,I267404);
DFFARX1 I_15567 (I267520,I2859,I267234,I267220,);
nand I_15568 (I267551,I388957,I388948);
and I_15569 (I267568,I267551,I388960);
DFFARX1 I_15570 (I267568,I2859,I267234,I267594,);
nor I_15571 (I267602,I267594,I267461);
DFFARX1 I_15572 (I267602,I2859,I267234,I267202,);
nand I_15573 (I267633,I267594,I267503);
nand I_15574 (I267211,I267486,I267633);
not I_15575 (I267664,I267594);
nor I_15576 (I267681,I267664,I267404);
DFFARX1 I_15577 (I267681,I2859,I267234,I267223,);
nor I_15578 (I267712,I388945,I388948);
or I_15579 (I267214,I267461,I267712);
nor I_15580 (I267205,I267594,I267712);
or I_15581 (I267208,I267328,I267712);
DFFARX1 I_15582 (I267712,I2859,I267234,I267226,);
not I_15583 (I267812,I2866);
DFFARX1 I_15584 (I443544,I2859,I267812,I267838,);
not I_15585 (I267846,I267838);
nand I_15586 (I267863,I443526,I443538);
and I_15587 (I267880,I267863,I443541);
DFFARX1 I_15588 (I267880,I2859,I267812,I267906,);
not I_15589 (I267914,I443535);
DFFARX1 I_15590 (I443532,I2859,I267812,I267940,);
not I_15591 (I267948,I267940);
nor I_15592 (I267965,I267948,I267846);
and I_15593 (I267982,I267965,I443535);
nor I_15594 (I267999,I267948,I267914);
nor I_15595 (I267795,I267906,I267999);
DFFARX1 I_15596 (I443550,I2859,I267812,I268039,);
nor I_15597 (I268047,I268039,I267906);
not I_15598 (I268064,I268047);
not I_15599 (I268081,I268039);
nor I_15600 (I268098,I268081,I267982);
DFFARX1 I_15601 (I268098,I2859,I267812,I267798,);
nand I_15602 (I268129,I443529,I443529);
and I_15603 (I268146,I268129,I443526);
DFFARX1 I_15604 (I268146,I2859,I267812,I268172,);
nor I_15605 (I268180,I268172,I268039);
DFFARX1 I_15606 (I268180,I2859,I267812,I267780,);
nand I_15607 (I268211,I268172,I268081);
nand I_15608 (I267789,I268064,I268211);
not I_15609 (I268242,I268172);
nor I_15610 (I268259,I268242,I267982);
DFFARX1 I_15611 (I268259,I2859,I267812,I267801,);
nor I_15612 (I268290,I443547,I443529);
or I_15613 (I267792,I268039,I268290);
nor I_15614 (I267783,I268172,I268290);
or I_15615 (I267786,I267906,I268290);
DFFARX1 I_15616 (I268290,I2859,I267812,I267804,);
not I_15617 (I268390,I2866);
DFFARX1 I_15618 (I14815,I2859,I268390,I268416,);
not I_15619 (I268424,I268416);
nand I_15620 (I268441,I14812,I14803);
and I_15621 (I268458,I268441,I14803);
DFFARX1 I_15622 (I268458,I2859,I268390,I268484,);
not I_15623 (I268492,I14806);
DFFARX1 I_15624 (I14821,I2859,I268390,I268518,);
not I_15625 (I268526,I268518);
nor I_15626 (I268543,I268526,I268424);
and I_15627 (I268560,I268543,I14806);
nor I_15628 (I268577,I268526,I268492);
nor I_15629 (I268373,I268484,I268577);
DFFARX1 I_15630 (I14806,I2859,I268390,I268617,);
nor I_15631 (I268625,I268617,I268484);
not I_15632 (I268642,I268625);
not I_15633 (I268659,I268617);
nor I_15634 (I268676,I268659,I268560);
DFFARX1 I_15635 (I268676,I2859,I268390,I268376,);
nand I_15636 (I268707,I14824,I14809);
and I_15637 (I268724,I268707,I14827);
DFFARX1 I_15638 (I268724,I2859,I268390,I268750,);
nor I_15639 (I268758,I268750,I268617);
DFFARX1 I_15640 (I268758,I2859,I268390,I268358,);
nand I_15641 (I268789,I268750,I268659);
nand I_15642 (I268367,I268642,I268789);
not I_15643 (I268820,I268750);
nor I_15644 (I268837,I268820,I268560);
DFFARX1 I_15645 (I268837,I2859,I268390,I268379,);
nor I_15646 (I268868,I14818,I14809);
or I_15647 (I268370,I268617,I268868);
nor I_15648 (I268361,I268750,I268868);
or I_15649 (I268364,I268484,I268868);
DFFARX1 I_15650 (I268868,I2859,I268390,I268382,);
not I_15651 (I268968,I2866);
DFFARX1 I_15652 (I548732,I2859,I268968,I268994,);
not I_15653 (I269002,I268994);
nand I_15654 (I269019,I548717,I548705);
and I_15655 (I269036,I269019,I548720);
DFFARX1 I_15656 (I269036,I2859,I268968,I269062,);
not I_15657 (I269070,I548705);
DFFARX1 I_15658 (I548723,I2859,I268968,I269096,);
not I_15659 (I269104,I269096);
nor I_15660 (I269121,I269104,I269002);
and I_15661 (I269138,I269121,I548705);
nor I_15662 (I269155,I269104,I269070);
nor I_15663 (I268951,I269062,I269155);
DFFARX1 I_15664 (I548711,I2859,I268968,I269195,);
nor I_15665 (I269203,I269195,I269062);
not I_15666 (I269220,I269203);
not I_15667 (I269237,I269195);
nor I_15668 (I269254,I269237,I269138);
DFFARX1 I_15669 (I269254,I2859,I268968,I268954,);
nand I_15670 (I269285,I548708,I548714);
and I_15671 (I269302,I269285,I548729);
DFFARX1 I_15672 (I269302,I2859,I268968,I269328,);
nor I_15673 (I269336,I269328,I269195);
DFFARX1 I_15674 (I269336,I2859,I268968,I268936,);
nand I_15675 (I269367,I269328,I269237);
nand I_15676 (I268945,I269220,I269367);
not I_15677 (I269398,I269328);
nor I_15678 (I269415,I269398,I269138);
DFFARX1 I_15679 (I269415,I2859,I268968,I268957,);
nor I_15680 (I269446,I548726,I548714);
or I_15681 (I268948,I269195,I269446);
nor I_15682 (I268939,I269328,I269446);
or I_15683 (I268942,I269062,I269446);
DFFARX1 I_15684 (I269446,I2859,I268968,I268960,);
not I_15685 (I269546,I2866);
DFFARX1 I_15686 (I426005,I2859,I269546,I269572,);
not I_15687 (I269580,I269572);
nand I_15688 (I269597,I426002,I426020);
and I_15689 (I269614,I269597,I426017);
DFFARX1 I_15690 (I269614,I2859,I269546,I269640,);
not I_15691 (I269648,I425999);
DFFARX1 I_15692 (I426002,I2859,I269546,I269674,);
not I_15693 (I269682,I269674);
nor I_15694 (I269699,I269682,I269580);
and I_15695 (I269716,I269699,I425999);
nor I_15696 (I269733,I269682,I269648);
nor I_15697 (I269529,I269640,I269733);
DFFARX1 I_15698 (I426011,I2859,I269546,I269773,);
nor I_15699 (I269781,I269773,I269640);
not I_15700 (I269798,I269781);
not I_15701 (I269815,I269773);
nor I_15702 (I269832,I269815,I269716);
DFFARX1 I_15703 (I269832,I2859,I269546,I269532,);
nand I_15704 (I269863,I426014,I425999);
and I_15705 (I269880,I269863,I426005);
DFFARX1 I_15706 (I269880,I2859,I269546,I269906,);
nor I_15707 (I269914,I269906,I269773);
DFFARX1 I_15708 (I269914,I2859,I269546,I269514,);
nand I_15709 (I269945,I269906,I269815);
nand I_15710 (I269523,I269798,I269945);
not I_15711 (I269976,I269906);
nor I_15712 (I269993,I269976,I269716);
DFFARX1 I_15713 (I269993,I2859,I269546,I269535,);
nor I_15714 (I270024,I426008,I425999);
or I_15715 (I269526,I269773,I270024);
nor I_15716 (I269517,I269906,I270024);
or I_15717 (I269520,I269640,I270024);
DFFARX1 I_15718 (I270024,I2859,I269546,I269538,);
not I_15719 (I270124,I2866);
DFFARX1 I_15720 (I140933,I2859,I270124,I270150,);
not I_15721 (I270158,I270150);
nand I_15722 (I270175,I140936,I140912);
and I_15723 (I270192,I270175,I140909);
DFFARX1 I_15724 (I270192,I2859,I270124,I270218,);
not I_15725 (I270226,I140915);
DFFARX1 I_15726 (I140909,I2859,I270124,I270252,);
not I_15727 (I270260,I270252);
nor I_15728 (I270277,I270260,I270158);
and I_15729 (I270294,I270277,I140915);
nor I_15730 (I270311,I270260,I270226);
nor I_15731 (I270107,I270218,I270311);
DFFARX1 I_15732 (I140918,I2859,I270124,I270351,);
nor I_15733 (I270359,I270351,I270218);
not I_15734 (I270376,I270359);
not I_15735 (I270393,I270351);
nor I_15736 (I270410,I270393,I270294);
DFFARX1 I_15737 (I270410,I2859,I270124,I270110,);
nand I_15738 (I270441,I140921,I140930);
and I_15739 (I270458,I270441,I140927);
DFFARX1 I_15740 (I270458,I2859,I270124,I270484,);
nor I_15741 (I270492,I270484,I270351);
DFFARX1 I_15742 (I270492,I2859,I270124,I270092,);
nand I_15743 (I270523,I270484,I270393);
nand I_15744 (I270101,I270376,I270523);
not I_15745 (I270554,I270484);
nor I_15746 (I270571,I270554,I270294);
DFFARX1 I_15747 (I270571,I2859,I270124,I270113,);
nor I_15748 (I270602,I140924,I140930);
or I_15749 (I270104,I270351,I270602);
nor I_15750 (I270095,I270484,I270602);
or I_15751 (I270098,I270218,I270602);
DFFARX1 I_15752 (I270602,I2859,I270124,I270116,);
not I_15753 (I270702,I2866);
DFFARX1 I_15754 (I546947,I2859,I270702,I270728,);
not I_15755 (I270736,I270728);
nand I_15756 (I270753,I546932,I546920);
and I_15757 (I270770,I270753,I546935);
DFFARX1 I_15758 (I270770,I2859,I270702,I270796,);
not I_15759 (I270804,I546920);
DFFARX1 I_15760 (I546938,I2859,I270702,I270830,);
not I_15761 (I270838,I270830);
nor I_15762 (I270855,I270838,I270736);
and I_15763 (I270872,I270855,I546920);
nor I_15764 (I270889,I270838,I270804);
nor I_15765 (I270685,I270796,I270889);
DFFARX1 I_15766 (I546926,I2859,I270702,I270929,);
nor I_15767 (I270937,I270929,I270796);
not I_15768 (I270954,I270937);
not I_15769 (I270971,I270929);
nor I_15770 (I270988,I270971,I270872);
DFFARX1 I_15771 (I270988,I2859,I270702,I270688,);
nand I_15772 (I271019,I546923,I546929);
and I_15773 (I271036,I271019,I546944);
DFFARX1 I_15774 (I271036,I2859,I270702,I271062,);
nor I_15775 (I271070,I271062,I270929);
DFFARX1 I_15776 (I271070,I2859,I270702,I270670,);
nand I_15777 (I271101,I271062,I270971);
nand I_15778 (I270679,I270954,I271101);
not I_15779 (I271132,I271062);
nor I_15780 (I271149,I271132,I270872);
DFFARX1 I_15781 (I271149,I2859,I270702,I270691,);
nor I_15782 (I271180,I546941,I546929);
or I_15783 (I270682,I270929,I271180);
nor I_15784 (I270673,I271062,I271180);
or I_15785 (I270676,I270796,I271180);
DFFARX1 I_15786 (I271180,I2859,I270702,I270694,);
not I_15787 (I271280,I2866);
DFFARX1 I_15788 (I363123,I2859,I271280,I271306,);
not I_15789 (I271314,I271306);
nand I_15790 (I271331,I363099,I363114);
and I_15791 (I271348,I271331,I363126);
DFFARX1 I_15792 (I271348,I2859,I271280,I271374,);
not I_15793 (I271382,I363111);
DFFARX1 I_15794 (I363102,I2859,I271280,I271408,);
not I_15795 (I271416,I271408);
nor I_15796 (I271433,I271416,I271314);
and I_15797 (I271450,I271433,I363111);
nor I_15798 (I271467,I271416,I271382);
nor I_15799 (I271263,I271374,I271467);
DFFARX1 I_15800 (I363099,I2859,I271280,I271507,);
nor I_15801 (I271515,I271507,I271374);
not I_15802 (I271532,I271515);
not I_15803 (I271549,I271507);
nor I_15804 (I271566,I271549,I271450);
DFFARX1 I_15805 (I271566,I2859,I271280,I271266,);
nand I_15806 (I271597,I363117,I363108);
and I_15807 (I271614,I271597,I363120);
DFFARX1 I_15808 (I271614,I2859,I271280,I271640,);
nor I_15809 (I271648,I271640,I271507);
DFFARX1 I_15810 (I271648,I2859,I271280,I271248,);
nand I_15811 (I271679,I271640,I271549);
nand I_15812 (I271257,I271532,I271679);
not I_15813 (I271710,I271640);
nor I_15814 (I271727,I271710,I271450);
DFFARX1 I_15815 (I271727,I2859,I271280,I271269,);
nor I_15816 (I271758,I363105,I363108);
or I_15817 (I271260,I271507,I271758);
nor I_15818 (I271251,I271640,I271758);
or I_15819 (I271254,I271374,I271758);
DFFARX1 I_15820 (I271758,I2859,I271280,I271272,);
not I_15821 (I271858,I2866);
DFFARX1 I_15822 (I2244,I2859,I271858,I271884,);
not I_15823 (I271892,I271884);
nand I_15824 (I271909,I2460,I2740);
and I_15825 (I271926,I271909,I2252);
DFFARX1 I_15826 (I271926,I2859,I271858,I271952,);
not I_15827 (I271960,I2620);
DFFARX1 I_15828 (I2468,I2859,I271858,I271986,);
not I_15829 (I271994,I271986);
nor I_15830 (I272011,I271994,I271892);
and I_15831 (I272028,I272011,I2620);
nor I_15832 (I272045,I271994,I271960);
nor I_15833 (I271841,I271952,I272045);
DFFARX1 I_15834 (I1892,I2859,I271858,I272085,);
nor I_15835 (I272093,I272085,I271952);
not I_15836 (I272110,I272093);
not I_15837 (I272127,I272085);
nor I_15838 (I272144,I272127,I272028);
DFFARX1 I_15839 (I272144,I2859,I271858,I271844,);
nand I_15840 (I272175,I1716,I1772);
and I_15841 (I272192,I272175,I1492);
DFFARX1 I_15842 (I272192,I2859,I271858,I272218,);
nor I_15843 (I272226,I272218,I272085);
DFFARX1 I_15844 (I272226,I2859,I271858,I271826,);
nand I_15845 (I272257,I272218,I272127);
nand I_15846 (I271835,I272110,I272257);
not I_15847 (I272288,I272218);
nor I_15848 (I272305,I272288,I272028);
DFFARX1 I_15849 (I272305,I2859,I271858,I271847,);
nor I_15850 (I272336,I1660,I1772);
or I_15851 (I271838,I272085,I272336);
nor I_15852 (I271829,I272218,I272336);
or I_15853 (I271832,I271952,I272336);
DFFARX1 I_15854 (I272336,I2859,I271858,I271850,);
not I_15855 (I272436,I2866);
DFFARX1 I_15856 (I30089,I2859,I272436,I272462,);
not I_15857 (I272470,I272462);
nand I_15858 (I272487,I30098,I30107);
and I_15859 (I272504,I272487,I30086);
DFFARX1 I_15860 (I272504,I2859,I272436,I272530,);
not I_15861 (I272538,I30089);
DFFARX1 I_15862 (I30104,I2859,I272436,I272564,);
not I_15863 (I272572,I272564);
nor I_15864 (I272589,I272572,I272470);
and I_15865 (I272606,I272589,I30089);
nor I_15866 (I272623,I272572,I272538);
nor I_15867 (I272419,I272530,I272623);
DFFARX1 I_15868 (I30095,I2859,I272436,I272663,);
nor I_15869 (I272671,I272663,I272530);
not I_15870 (I272688,I272671);
not I_15871 (I272705,I272663);
nor I_15872 (I272722,I272705,I272606);
DFFARX1 I_15873 (I272722,I2859,I272436,I272422,);
nand I_15874 (I272753,I30110,I30086);
and I_15875 (I272770,I272753,I30092);
DFFARX1 I_15876 (I272770,I2859,I272436,I272796,);
nor I_15877 (I272804,I272796,I272663);
DFFARX1 I_15878 (I272804,I2859,I272436,I272404,);
nand I_15879 (I272835,I272796,I272705);
nand I_15880 (I272413,I272688,I272835);
not I_15881 (I272866,I272796);
nor I_15882 (I272883,I272866,I272606);
DFFARX1 I_15883 (I272883,I2859,I272436,I272425,);
nor I_15884 (I272914,I30101,I30086);
or I_15885 (I272416,I272663,I272914);
nor I_15886 (I272407,I272796,I272914);
or I_15887 (I272410,I272530,I272914);
DFFARX1 I_15888 (I272914,I2859,I272436,I272428,);
not I_15889 (I273014,I2866);
DFFARX1 I_15890 (I390255,I2859,I273014,I273040,);
not I_15891 (I273048,I273040);
nand I_15892 (I273065,I390231,I390246);
and I_15893 (I273082,I273065,I390258);
DFFARX1 I_15894 (I273082,I2859,I273014,I273108,);
not I_15895 (I273116,I390243);
DFFARX1 I_15896 (I390234,I2859,I273014,I273142,);
not I_15897 (I273150,I273142);
nor I_15898 (I273167,I273150,I273048);
and I_15899 (I273184,I273167,I390243);
nor I_15900 (I273201,I273150,I273116);
nor I_15901 (I272997,I273108,I273201);
DFFARX1 I_15902 (I390231,I2859,I273014,I273241,);
nor I_15903 (I273249,I273241,I273108);
not I_15904 (I273266,I273249);
not I_15905 (I273283,I273241);
nor I_15906 (I273300,I273283,I273184);
DFFARX1 I_15907 (I273300,I2859,I273014,I273000,);
nand I_15908 (I273331,I390249,I390240);
and I_15909 (I273348,I273331,I390252);
DFFARX1 I_15910 (I273348,I2859,I273014,I273374,);
nor I_15911 (I273382,I273374,I273241);
DFFARX1 I_15912 (I273382,I2859,I273014,I272982,);
nand I_15913 (I273413,I273374,I273283);
nand I_15914 (I272991,I273266,I273413);
not I_15915 (I273444,I273374);
nor I_15916 (I273461,I273444,I273184);
DFFARX1 I_15917 (I273461,I2859,I273014,I273003,);
nor I_15918 (I273492,I390237,I390240);
or I_15919 (I272994,I273241,I273492);
nor I_15920 (I272985,I273374,I273492);
or I_15921 (I272988,I273108,I273492);
DFFARX1 I_15922 (I273492,I2859,I273014,I273006,);
not I_15923 (I273592,I2866);
DFFARX1 I_15924 (I366353,I2859,I273592,I273618,);
not I_15925 (I273626,I273618);
nand I_15926 (I273643,I366329,I366344);
and I_15927 (I273660,I273643,I366356);
DFFARX1 I_15928 (I273660,I2859,I273592,I273686,);
not I_15929 (I273694,I366341);
DFFARX1 I_15930 (I366332,I2859,I273592,I273720,);
not I_15931 (I273728,I273720);
nor I_15932 (I273745,I273728,I273626);
and I_15933 (I273762,I273745,I366341);
nor I_15934 (I273779,I273728,I273694);
nor I_15935 (I273575,I273686,I273779);
DFFARX1 I_15936 (I366329,I2859,I273592,I273819,);
nor I_15937 (I273827,I273819,I273686);
not I_15938 (I273844,I273827);
not I_15939 (I273861,I273819);
nor I_15940 (I273878,I273861,I273762);
DFFARX1 I_15941 (I273878,I2859,I273592,I273578,);
nand I_15942 (I273909,I366347,I366338);
and I_15943 (I273926,I273909,I366350);
DFFARX1 I_15944 (I273926,I2859,I273592,I273952,);
nor I_15945 (I273960,I273952,I273819);
DFFARX1 I_15946 (I273960,I2859,I273592,I273560,);
nand I_15947 (I273991,I273952,I273861);
nand I_15948 (I273569,I273844,I273991);
not I_15949 (I274022,I273952);
nor I_15950 (I274039,I274022,I273762);
DFFARX1 I_15951 (I274039,I2859,I273592,I273581,);
nor I_15952 (I274070,I366335,I366338);
or I_15953 (I273572,I273819,I274070);
nor I_15954 (I273563,I273952,I274070);
or I_15955 (I273566,I273686,I274070);
DFFARX1 I_15956 (I274070,I2859,I273592,I273584,);
not I_15957 (I274170,I2866);
DFFARX1 I_15958 (I517170,I2859,I274170,I274196,);
not I_15959 (I274204,I274196);
nand I_15960 (I274221,I517194,I517176);
and I_15961 (I274238,I274221,I517182);
DFFARX1 I_15962 (I274238,I2859,I274170,I274264,);
not I_15963 (I274272,I517188);
DFFARX1 I_15964 (I517173,I2859,I274170,I274298,);
not I_15965 (I274306,I274298);
nor I_15966 (I274323,I274306,I274204);
and I_15967 (I274340,I274323,I517188);
nor I_15968 (I274357,I274306,I274272);
nor I_15969 (I274153,I274264,I274357);
DFFARX1 I_15970 (I517185,I2859,I274170,I274397,);
nor I_15971 (I274405,I274397,I274264);
not I_15972 (I274422,I274405);
not I_15973 (I274439,I274397);
nor I_15974 (I274456,I274439,I274340);
DFFARX1 I_15975 (I274456,I2859,I274170,I274156,);
nand I_15976 (I274487,I517191,I517179);
and I_15977 (I274504,I274487,I517173);
DFFARX1 I_15978 (I274504,I2859,I274170,I274530,);
nor I_15979 (I274538,I274530,I274397);
DFFARX1 I_15980 (I274538,I2859,I274170,I274138,);
nand I_15981 (I274569,I274530,I274439);
nand I_15982 (I274147,I274422,I274569);
not I_15983 (I274600,I274530);
nor I_15984 (I274617,I274600,I274340);
DFFARX1 I_15985 (I274617,I2859,I274170,I274159,);
nor I_15986 (I274648,I517170,I517179);
or I_15987 (I274150,I274397,I274648);
nor I_15988 (I274141,I274530,I274648);
or I_15989 (I274144,I274264,I274648);
DFFARX1 I_15990 (I274648,I2859,I274170,I274162,);
not I_15991 (I274748,I2866);
DFFARX1 I_15992 (I466664,I2859,I274748,I274774,);
not I_15993 (I274782,I274774);
nand I_15994 (I274799,I466646,I466658);
and I_15995 (I274816,I274799,I466661);
DFFARX1 I_15996 (I274816,I2859,I274748,I274842,);
not I_15997 (I274850,I466655);
DFFARX1 I_15998 (I466652,I2859,I274748,I274876,);
not I_15999 (I274884,I274876);
nor I_16000 (I274901,I274884,I274782);
and I_16001 (I274918,I274901,I466655);
nor I_16002 (I274935,I274884,I274850);
nor I_16003 (I274731,I274842,I274935);
DFFARX1 I_16004 (I466670,I2859,I274748,I274975,);
nor I_16005 (I274983,I274975,I274842);
not I_16006 (I275000,I274983);
not I_16007 (I275017,I274975);
nor I_16008 (I275034,I275017,I274918);
DFFARX1 I_16009 (I275034,I2859,I274748,I274734,);
nand I_16010 (I275065,I466649,I466649);
and I_16011 (I275082,I275065,I466646);
DFFARX1 I_16012 (I275082,I2859,I274748,I275108,);
nor I_16013 (I275116,I275108,I274975);
DFFARX1 I_16014 (I275116,I2859,I274748,I274716,);
nand I_16015 (I275147,I275108,I275017);
nand I_16016 (I274725,I275000,I275147);
not I_16017 (I275178,I275108);
nor I_16018 (I275195,I275178,I274918);
DFFARX1 I_16019 (I275195,I2859,I274748,I274737,);
nor I_16020 (I275226,I466667,I466649);
or I_16021 (I274728,I274975,I275226);
nor I_16022 (I274719,I275108,I275226);
or I_16023 (I274722,I274842,I275226);
DFFARX1 I_16024 (I275226,I2859,I274748,I274740,);
not I_16025 (I275326,I2866);
DFFARX1 I_16026 (I389609,I2859,I275326,I275352,);
not I_16027 (I275360,I275352);
nand I_16028 (I275377,I389585,I389600);
and I_16029 (I275394,I275377,I389612);
DFFARX1 I_16030 (I275394,I2859,I275326,I275420,);
not I_16031 (I275428,I389597);
DFFARX1 I_16032 (I389588,I2859,I275326,I275454,);
not I_16033 (I275462,I275454);
nor I_16034 (I275479,I275462,I275360);
and I_16035 (I275496,I275479,I389597);
nor I_16036 (I275513,I275462,I275428);
nor I_16037 (I275309,I275420,I275513);
DFFARX1 I_16038 (I389585,I2859,I275326,I275553,);
nor I_16039 (I275561,I275553,I275420);
not I_16040 (I275578,I275561);
not I_16041 (I275595,I275553);
nor I_16042 (I275612,I275595,I275496);
DFFARX1 I_16043 (I275612,I2859,I275326,I275312,);
nand I_16044 (I275643,I389603,I389594);
and I_16045 (I275660,I275643,I389606);
DFFARX1 I_16046 (I275660,I2859,I275326,I275686,);
nor I_16047 (I275694,I275686,I275553);
DFFARX1 I_16048 (I275694,I2859,I275326,I275294,);
nand I_16049 (I275725,I275686,I275595);
nand I_16050 (I275303,I275578,I275725);
not I_16051 (I275756,I275686);
nor I_16052 (I275773,I275756,I275496);
DFFARX1 I_16053 (I275773,I2859,I275326,I275315,);
nor I_16054 (I275804,I389591,I389594);
or I_16055 (I275306,I275553,I275804);
nor I_16056 (I275297,I275686,I275804);
or I_16057 (I275300,I275420,I275804);
DFFARX1 I_16058 (I275804,I2859,I275326,I275318,);
not I_16059 (I275904,I2866);
DFFARX1 I_16060 (I240036,I2859,I275904,I275930,);
not I_16061 (I275938,I275930);
nand I_16062 (I275955,I240045,I240054);
and I_16063 (I275972,I275955,I240060);
DFFARX1 I_16064 (I275972,I2859,I275904,I275998,);
not I_16065 (I276006,I240057);
DFFARX1 I_16066 (I240042,I2859,I275904,I276032,);
not I_16067 (I276040,I276032);
nor I_16068 (I276057,I276040,I275938);
and I_16069 (I276074,I276057,I240057);
nor I_16070 (I276091,I276040,I276006);
nor I_16071 (I275887,I275998,I276091);
DFFARX1 I_16072 (I240051,I2859,I275904,I276131,);
nor I_16073 (I276139,I276131,I275998);
not I_16074 (I276156,I276139);
not I_16075 (I276173,I276131);
nor I_16076 (I276190,I276173,I276074);
DFFARX1 I_16077 (I276190,I2859,I275904,I275890,);
nand I_16078 (I276221,I240048,I240039);
and I_16079 (I276238,I276221,I240036);
DFFARX1 I_16080 (I276238,I2859,I275904,I276264,);
nor I_16081 (I276272,I276264,I276131);
DFFARX1 I_16082 (I276272,I2859,I275904,I275872,);
nand I_16083 (I276303,I276264,I276173);
nand I_16084 (I275881,I276156,I276303);
not I_16085 (I276334,I276264);
nor I_16086 (I276351,I276334,I276074);
DFFARX1 I_16087 (I276351,I2859,I275904,I275893,);
nor I_16088 (I276382,I240039,I240039);
or I_16089 (I275884,I276131,I276382);
nor I_16090 (I275875,I276264,I276382);
or I_16091 (I275878,I275998,I276382);
DFFARX1 I_16092 (I276382,I2859,I275904,I275896,);
not I_16093 (I276482,I2866);
DFFARX1 I_16094 (I215590,I2859,I276482,I276508,);
not I_16095 (I276516,I276508);
nand I_16096 (I276533,I215605,I215590);
and I_16097 (I276550,I276533,I215593);
DFFARX1 I_16098 (I276550,I2859,I276482,I276576,);
not I_16099 (I276584,I215593);
DFFARX1 I_16100 (I215602,I2859,I276482,I276610,);
not I_16101 (I276618,I276610);
nor I_16102 (I276635,I276618,I276516);
and I_16103 (I276652,I276635,I215593);
nor I_16104 (I276669,I276618,I276584);
nor I_16105 (I276465,I276576,I276669);
DFFARX1 I_16106 (I215596,I2859,I276482,I276709,);
nor I_16107 (I276717,I276709,I276576);
not I_16108 (I276734,I276717);
not I_16109 (I276751,I276709);
nor I_16110 (I276768,I276751,I276652);
DFFARX1 I_16111 (I276768,I2859,I276482,I276468,);
nand I_16112 (I276799,I215599,I215608);
and I_16113 (I276816,I276799,I215614);
DFFARX1 I_16114 (I276816,I2859,I276482,I276842,);
nor I_16115 (I276850,I276842,I276709);
DFFARX1 I_16116 (I276850,I2859,I276482,I276450,);
nand I_16117 (I276881,I276842,I276751);
nand I_16118 (I276459,I276734,I276881);
not I_16119 (I276912,I276842);
nor I_16120 (I276929,I276912,I276652);
DFFARX1 I_16121 (I276929,I2859,I276482,I276471,);
nor I_16122 (I276960,I215611,I215608);
or I_16123 (I276462,I276709,I276960);
nor I_16124 (I276453,I276842,I276960);
or I_16125 (I276456,I276576,I276960);
DFFARX1 I_16126 (I276960,I2859,I276482,I276474,);
not I_16127 (I277060,I2866);
DFFARX1 I_16128 (I323351,I2859,I277060,I277086,);
not I_16129 (I277094,I277086);
nand I_16130 (I277111,I323339,I323357);
and I_16131 (I277128,I277111,I323354);
DFFARX1 I_16132 (I277128,I2859,I277060,I277154,);
not I_16133 (I277162,I323345);
DFFARX1 I_16134 (I323342,I2859,I277060,I277188,);
not I_16135 (I277196,I277188);
nor I_16136 (I277213,I277196,I277094);
and I_16137 (I277230,I277213,I323345);
nor I_16138 (I277247,I277196,I277162);
nor I_16139 (I277043,I277154,I277247);
DFFARX1 I_16140 (I323336,I2859,I277060,I277287,);
nor I_16141 (I277295,I277287,I277154);
not I_16142 (I277312,I277295);
not I_16143 (I277329,I277287);
nor I_16144 (I277346,I277329,I277230);
DFFARX1 I_16145 (I277346,I2859,I277060,I277046,);
nand I_16146 (I277377,I323336,I323339);
and I_16147 (I277394,I277377,I323342);
DFFARX1 I_16148 (I277394,I2859,I277060,I277420,);
nor I_16149 (I277428,I277420,I277287);
DFFARX1 I_16150 (I277428,I2859,I277060,I277028,);
nand I_16151 (I277459,I277420,I277329);
nand I_16152 (I277037,I277312,I277459);
not I_16153 (I277490,I277420);
nor I_16154 (I277507,I277490,I277230);
DFFARX1 I_16155 (I277507,I2859,I277060,I277049,);
nor I_16156 (I277538,I323348,I323339);
or I_16157 (I277040,I277287,I277538);
nor I_16158 (I277031,I277420,I277538);
or I_16159 (I277034,I277154,I277538);
DFFARX1 I_16160 (I277538,I2859,I277060,I277052,);
not I_16161 (I277638,I2866);
DFFARX1 I_16162 (I129866,I2859,I277638,I277664,);
not I_16163 (I277672,I277664);
nand I_16164 (I277689,I129869,I129845);
and I_16165 (I277706,I277689,I129842);
DFFARX1 I_16166 (I277706,I2859,I277638,I277732,);
not I_16167 (I277740,I129848);
DFFARX1 I_16168 (I129842,I2859,I277638,I277766,);
not I_16169 (I277774,I277766);
nor I_16170 (I277791,I277774,I277672);
and I_16171 (I277808,I277791,I129848);
nor I_16172 (I277825,I277774,I277740);
nor I_16173 (I277621,I277732,I277825);
DFFARX1 I_16174 (I129851,I2859,I277638,I277865,);
nor I_16175 (I277873,I277865,I277732);
not I_16176 (I277890,I277873);
not I_16177 (I277907,I277865);
nor I_16178 (I277924,I277907,I277808);
DFFARX1 I_16179 (I277924,I2859,I277638,I277624,);
nand I_16180 (I277955,I129854,I129863);
and I_16181 (I277972,I277955,I129860);
DFFARX1 I_16182 (I277972,I2859,I277638,I277998,);
nor I_16183 (I278006,I277998,I277865);
DFFARX1 I_16184 (I278006,I2859,I277638,I277606,);
nand I_16185 (I278037,I277998,I277907);
nand I_16186 (I277615,I277890,I278037);
not I_16187 (I278068,I277998);
nor I_16188 (I278085,I278068,I277808);
DFFARX1 I_16189 (I278085,I2859,I277638,I277627,);
nor I_16190 (I278116,I129857,I129863);
or I_16191 (I277618,I277865,I278116);
nor I_16192 (I277609,I277998,I278116);
or I_16193 (I277612,I277732,I278116);
DFFARX1 I_16194 (I278116,I2859,I277638,I277630,);
not I_16195 (I278216,I2866);
DFFARX1 I_16196 (I357079,I2859,I278216,I278242,);
not I_16197 (I278250,I278242);
nand I_16198 (I278267,I357067,I357085);
and I_16199 (I278284,I278267,I357082);
DFFARX1 I_16200 (I278284,I2859,I278216,I278310,);
not I_16201 (I278318,I357073);
DFFARX1 I_16202 (I357070,I2859,I278216,I278344,);
not I_16203 (I278352,I278344);
nor I_16204 (I278369,I278352,I278250);
and I_16205 (I278386,I278369,I357073);
nor I_16206 (I278403,I278352,I278318);
nor I_16207 (I278199,I278310,I278403);
DFFARX1 I_16208 (I357064,I2859,I278216,I278443,);
nor I_16209 (I278451,I278443,I278310);
not I_16210 (I278468,I278451);
not I_16211 (I278485,I278443);
nor I_16212 (I278502,I278485,I278386);
DFFARX1 I_16213 (I278502,I2859,I278216,I278202,);
nand I_16214 (I278533,I357064,I357067);
and I_16215 (I278550,I278533,I357070);
DFFARX1 I_16216 (I278550,I2859,I278216,I278576,);
nor I_16217 (I278584,I278576,I278443);
DFFARX1 I_16218 (I278584,I2859,I278216,I278184,);
nand I_16219 (I278615,I278576,I278485);
nand I_16220 (I278193,I278468,I278615);
not I_16221 (I278646,I278576);
nor I_16222 (I278663,I278646,I278386);
DFFARX1 I_16223 (I278663,I2859,I278216,I278205,);
nor I_16224 (I278694,I357076,I357067);
or I_16225 (I278196,I278443,I278694);
nor I_16226 (I278187,I278576,I278694);
or I_16227 (I278190,I278310,I278694);
DFFARX1 I_16228 (I278694,I2859,I278216,I278208,);
not I_16229 (I278794,I2866);
DFFARX1 I_16230 (I519482,I2859,I278794,I278820,);
not I_16231 (I278828,I278820);
nand I_16232 (I278845,I519506,I519488);
and I_16233 (I278862,I278845,I519494);
DFFARX1 I_16234 (I278862,I2859,I278794,I278888,);
not I_16235 (I278896,I519500);
DFFARX1 I_16236 (I519485,I2859,I278794,I278922,);
not I_16237 (I278930,I278922);
nor I_16238 (I278947,I278930,I278828);
and I_16239 (I278964,I278947,I519500);
nor I_16240 (I278981,I278930,I278896);
nor I_16241 (I278777,I278888,I278981);
DFFARX1 I_16242 (I519497,I2859,I278794,I279021,);
nor I_16243 (I279029,I279021,I278888);
not I_16244 (I279046,I279029);
not I_16245 (I279063,I279021);
nor I_16246 (I279080,I279063,I278964);
DFFARX1 I_16247 (I279080,I2859,I278794,I278780,);
nand I_16248 (I279111,I519503,I519491);
and I_16249 (I279128,I279111,I519485);
DFFARX1 I_16250 (I279128,I2859,I278794,I279154,);
nor I_16251 (I279162,I279154,I279021);
DFFARX1 I_16252 (I279162,I2859,I278794,I278762,);
nand I_16253 (I279193,I279154,I279063);
nand I_16254 (I278771,I279046,I279193);
not I_16255 (I279224,I279154);
nor I_16256 (I279241,I279224,I278964);
DFFARX1 I_16257 (I279241,I2859,I278794,I278783,);
nor I_16258 (I279272,I519482,I519491);
or I_16259 (I278774,I279021,I279272);
nor I_16260 (I278765,I279154,I279272);
or I_16261 (I278768,I278888,I279272);
DFFARX1 I_16262 (I279272,I2859,I278794,I278786,);
not I_16263 (I279372,I2866);
DFFARX1 I_16264 (I527574,I2859,I279372,I279398,);
not I_16265 (I279406,I279398);
nand I_16266 (I279423,I527598,I527580);
and I_16267 (I279440,I279423,I527586);
DFFARX1 I_16268 (I279440,I2859,I279372,I279466,);
not I_16269 (I279474,I527592);
DFFARX1 I_16270 (I527577,I2859,I279372,I279500,);
not I_16271 (I279508,I279500);
nor I_16272 (I279525,I279508,I279406);
and I_16273 (I279542,I279525,I527592);
nor I_16274 (I279559,I279508,I279474);
nor I_16275 (I279355,I279466,I279559);
DFFARX1 I_16276 (I527589,I2859,I279372,I279599,);
nor I_16277 (I279607,I279599,I279466);
not I_16278 (I279624,I279607);
not I_16279 (I279641,I279599);
nor I_16280 (I279658,I279641,I279542);
DFFARX1 I_16281 (I279658,I2859,I279372,I279358,);
nand I_16282 (I279689,I527595,I527583);
and I_16283 (I279706,I279689,I527577);
DFFARX1 I_16284 (I279706,I2859,I279372,I279732,);
nor I_16285 (I279740,I279732,I279599);
DFFARX1 I_16286 (I279740,I2859,I279372,I279340,);
nand I_16287 (I279771,I279732,I279641);
nand I_16288 (I279349,I279624,I279771);
not I_16289 (I279802,I279732);
nor I_16290 (I279819,I279802,I279542);
DFFARX1 I_16291 (I279819,I2859,I279372,I279361,);
nor I_16292 (I279850,I527574,I527583);
or I_16293 (I279352,I279599,I279850);
nor I_16294 (I279343,I279732,I279850);
or I_16295 (I279346,I279466,I279850);
DFFARX1 I_16296 (I279850,I2859,I279372,I279364,);
not I_16297 (I279950,I2866);
DFFARX1 I_16298 (I346539,I2859,I279950,I279976,);
not I_16299 (I279984,I279976);
nand I_16300 (I280001,I346527,I346545);
and I_16301 (I280018,I280001,I346542);
DFFARX1 I_16302 (I280018,I2859,I279950,I280044,);
not I_16303 (I280052,I346533);
DFFARX1 I_16304 (I346530,I2859,I279950,I280078,);
not I_16305 (I280086,I280078);
nor I_16306 (I280103,I280086,I279984);
and I_16307 (I280120,I280103,I346533);
nor I_16308 (I280137,I280086,I280052);
nor I_16309 (I279933,I280044,I280137);
DFFARX1 I_16310 (I346524,I2859,I279950,I280177,);
nor I_16311 (I280185,I280177,I280044);
not I_16312 (I280202,I280185);
not I_16313 (I280219,I280177);
nor I_16314 (I280236,I280219,I280120);
DFFARX1 I_16315 (I280236,I2859,I279950,I279936,);
nand I_16316 (I280267,I346524,I346527);
and I_16317 (I280284,I280267,I346530);
DFFARX1 I_16318 (I280284,I2859,I279950,I280310,);
nor I_16319 (I280318,I280310,I280177);
DFFARX1 I_16320 (I280318,I2859,I279950,I279918,);
nand I_16321 (I280349,I280310,I280219);
nand I_16322 (I279927,I280202,I280349);
not I_16323 (I280380,I280310);
nor I_16324 (I280397,I280380,I280120);
DFFARX1 I_16325 (I280397,I2859,I279950,I279939,);
nor I_16326 (I280428,I346536,I346527);
or I_16327 (I279930,I280177,I280428);
nor I_16328 (I279921,I280310,I280428);
or I_16329 (I279924,I280044,I280428);
DFFARX1 I_16330 (I280428,I2859,I279950,I279942,);
not I_16331 (I280528,I2866);
DFFARX1 I_16332 (I5856,I2859,I280528,I280554,);
not I_16333 (I280562,I280554);
nand I_16334 (I280579,I5853,I5844);
and I_16335 (I280596,I280579,I5844);
DFFARX1 I_16336 (I280596,I2859,I280528,I280622,);
not I_16337 (I280630,I5847);
DFFARX1 I_16338 (I5862,I2859,I280528,I280656,);
not I_16339 (I280664,I280656);
nor I_16340 (I280681,I280664,I280562);
and I_16341 (I280698,I280681,I5847);
nor I_16342 (I280715,I280664,I280630);
nor I_16343 (I280511,I280622,I280715);
DFFARX1 I_16344 (I5847,I2859,I280528,I280755,);
nor I_16345 (I280763,I280755,I280622);
not I_16346 (I280780,I280763);
not I_16347 (I280797,I280755);
nor I_16348 (I280814,I280797,I280698);
DFFARX1 I_16349 (I280814,I2859,I280528,I280514,);
nand I_16350 (I280845,I5865,I5850);
and I_16351 (I280862,I280845,I5868);
DFFARX1 I_16352 (I280862,I2859,I280528,I280888,);
nor I_16353 (I280896,I280888,I280755);
DFFARX1 I_16354 (I280896,I2859,I280528,I280496,);
nand I_16355 (I280927,I280888,I280797);
nand I_16356 (I280505,I280780,I280927);
not I_16357 (I280958,I280888);
nor I_16358 (I280975,I280958,I280698);
DFFARX1 I_16359 (I280975,I2859,I280528,I280517,);
nor I_16360 (I281006,I5859,I5850);
or I_16361 (I280508,I280755,I281006);
nor I_16362 (I280499,I280888,I281006);
or I_16363 (I280502,I280622,I281006);
DFFARX1 I_16364 (I281006,I2859,I280528,I280520,);
not I_16365 (I281106,I2866);
DFFARX1 I_16366 (I408343,I2859,I281106,I281132,);
not I_16367 (I281140,I281132);
nand I_16368 (I281157,I408319,I408334);
and I_16369 (I281174,I281157,I408346);
DFFARX1 I_16370 (I281174,I2859,I281106,I281200,);
not I_16371 (I281208,I408331);
DFFARX1 I_16372 (I408322,I2859,I281106,I281234,);
not I_16373 (I281242,I281234);
nor I_16374 (I281259,I281242,I281140);
and I_16375 (I281276,I281259,I408331);
nor I_16376 (I281293,I281242,I281208);
nor I_16377 (I281089,I281200,I281293);
DFFARX1 I_16378 (I408319,I2859,I281106,I281333,);
nor I_16379 (I281341,I281333,I281200);
not I_16380 (I281358,I281341);
not I_16381 (I281375,I281333);
nor I_16382 (I281392,I281375,I281276);
DFFARX1 I_16383 (I281392,I2859,I281106,I281092,);
nand I_16384 (I281423,I408337,I408328);
and I_16385 (I281440,I281423,I408340);
DFFARX1 I_16386 (I281440,I2859,I281106,I281466,);
nor I_16387 (I281474,I281466,I281333);
DFFARX1 I_16388 (I281474,I2859,I281106,I281074,);
nand I_16389 (I281505,I281466,I281375);
nand I_16390 (I281083,I281358,I281505);
not I_16391 (I281536,I281466);
nor I_16392 (I281553,I281536,I281276);
DFFARX1 I_16393 (I281553,I2859,I281106,I281095,);
nor I_16394 (I281584,I408325,I408328);
or I_16395 (I281086,I281333,I281584);
nor I_16396 (I281077,I281466,I281584);
or I_16397 (I281080,I281200,I281584);
DFFARX1 I_16398 (I281584,I2859,I281106,I281098,);
not I_16399 (I281684,I2866);
DFFARX1 I_16400 (I119326,I2859,I281684,I281710,);
not I_16401 (I281718,I281710);
nand I_16402 (I281735,I119329,I119305);
and I_16403 (I281752,I281735,I119302);
DFFARX1 I_16404 (I281752,I2859,I281684,I281778,);
not I_16405 (I281786,I119308);
DFFARX1 I_16406 (I119302,I2859,I281684,I281812,);
not I_16407 (I281820,I281812);
nor I_16408 (I281837,I281820,I281718);
and I_16409 (I281854,I281837,I119308);
nor I_16410 (I281871,I281820,I281786);
nor I_16411 (I281667,I281778,I281871);
DFFARX1 I_16412 (I119311,I2859,I281684,I281911,);
nor I_16413 (I281919,I281911,I281778);
not I_16414 (I281936,I281919);
not I_16415 (I281953,I281911);
nor I_16416 (I281970,I281953,I281854);
DFFARX1 I_16417 (I281970,I2859,I281684,I281670,);
nand I_16418 (I282001,I119314,I119323);
and I_16419 (I282018,I282001,I119320);
DFFARX1 I_16420 (I282018,I2859,I281684,I282044,);
nor I_16421 (I282052,I282044,I281911);
DFFARX1 I_16422 (I282052,I2859,I281684,I281652,);
nand I_16423 (I282083,I282044,I281953);
nand I_16424 (I281661,I281936,I282083);
not I_16425 (I282114,I282044);
nor I_16426 (I282131,I282114,I281854);
DFFARX1 I_16427 (I282131,I2859,I281684,I281673,);
nor I_16428 (I282162,I119317,I119323);
or I_16429 (I281664,I281911,I282162);
nor I_16430 (I281655,I282044,I282162);
or I_16431 (I281658,I281778,I282162);
DFFARX1 I_16432 (I282162,I2859,I281684,I281676,);
not I_16433 (I282262,I2866);
DFFARX1 I_16434 (I485738,I2859,I282262,I282288,);
not I_16435 (I282296,I282288);
nand I_16436 (I282313,I485720,I485732);
and I_16437 (I282330,I282313,I485735);
DFFARX1 I_16438 (I282330,I2859,I282262,I282356,);
not I_16439 (I282364,I485729);
DFFARX1 I_16440 (I485726,I2859,I282262,I282390,);
not I_16441 (I282398,I282390);
nor I_16442 (I282415,I282398,I282296);
and I_16443 (I282432,I282415,I485729);
nor I_16444 (I282449,I282398,I282364);
nor I_16445 (I282245,I282356,I282449);
DFFARX1 I_16446 (I485744,I2859,I282262,I282489,);
nor I_16447 (I282497,I282489,I282356);
not I_16448 (I282514,I282497);
not I_16449 (I282531,I282489);
nor I_16450 (I282548,I282531,I282432);
DFFARX1 I_16451 (I282548,I2859,I282262,I282248,);
nand I_16452 (I282579,I485723,I485723);
and I_16453 (I282596,I282579,I485720);
DFFARX1 I_16454 (I282596,I2859,I282262,I282622,);
nor I_16455 (I282630,I282622,I282489);
DFFARX1 I_16456 (I282630,I2859,I282262,I282230,);
nand I_16457 (I282661,I282622,I282531);
nand I_16458 (I282239,I282514,I282661);
not I_16459 (I282692,I282622);
nor I_16460 (I282709,I282692,I282432);
DFFARX1 I_16461 (I282709,I2859,I282262,I282251,);
nor I_16462 (I282740,I485741,I485723);
or I_16463 (I282242,I282489,I282740);
nor I_16464 (I282233,I282622,I282740);
or I_16465 (I282236,I282356,I282740);
DFFARX1 I_16466 (I282740,I2859,I282262,I282254,);
not I_16467 (I282840,I2866);
DFFARX1 I_16468 (I78672,I2859,I282840,I282866,);
not I_16469 (I282874,I282866);
nand I_16470 (I282891,I78675,I78696);
and I_16471 (I282908,I282891,I78684);
DFFARX1 I_16472 (I282908,I2859,I282840,I282934,);
not I_16473 (I282942,I78681);
DFFARX1 I_16474 (I78672,I2859,I282840,I282968,);
not I_16475 (I282976,I282968);
nor I_16476 (I282993,I282976,I282874);
and I_16477 (I283010,I282993,I78681);
nor I_16478 (I283027,I282976,I282942);
nor I_16479 (I282823,I282934,I283027);
DFFARX1 I_16480 (I78690,I2859,I282840,I283067,);
nor I_16481 (I283075,I283067,I282934);
not I_16482 (I283092,I283075);
not I_16483 (I283109,I283067);
nor I_16484 (I283126,I283109,I283010);
DFFARX1 I_16485 (I283126,I2859,I282840,I282826,);
nand I_16486 (I283157,I78675,I78678);
and I_16487 (I283174,I283157,I78687);
DFFARX1 I_16488 (I283174,I2859,I282840,I283200,);
nor I_16489 (I283208,I283200,I283067);
DFFARX1 I_16490 (I283208,I2859,I282840,I282808,);
nand I_16491 (I283239,I283200,I283109);
nand I_16492 (I282817,I283092,I283239);
not I_16493 (I283270,I283200);
nor I_16494 (I283287,I283270,I283010);
DFFARX1 I_16495 (I283287,I2859,I282840,I282829,);
nor I_16496 (I283318,I78693,I78678);
or I_16497 (I282820,I283067,I283318);
nor I_16498 (I282811,I283200,I283318);
or I_16499 (I282814,I282934,I283318);
DFFARX1 I_16500 (I283318,I2859,I282840,I282832,);
not I_16501 (I283418,I2866);
DFFARX1 I_16502 (I1684,I2859,I283418,I283444,);
not I_16503 (I283452,I283444);
nand I_16504 (I283469,I2052,I1548);
and I_16505 (I283486,I283469,I2476);
DFFARX1 I_16506 (I283486,I2859,I283418,I283512,);
not I_16507 (I283520,I2852);
DFFARX1 I_16508 (I1372,I2859,I283418,I283546,);
not I_16509 (I283554,I283546);
nor I_16510 (I283571,I283554,I283452);
and I_16511 (I283588,I283571,I2852);
nor I_16512 (I283605,I283554,I283520);
nor I_16513 (I283401,I283512,I283605);
DFFARX1 I_16514 (I1868,I2859,I283418,I283645,);
nor I_16515 (I283653,I283645,I283512);
not I_16516 (I283670,I283653);
not I_16517 (I283687,I283645);
nor I_16518 (I283704,I283687,I283588);
DFFARX1 I_16519 (I283704,I2859,I283418,I283404,);
nand I_16520 (I283735,I2100,I1652);
and I_16521 (I283752,I283735,I2676);
DFFARX1 I_16522 (I283752,I2859,I283418,I283778,);
nor I_16523 (I283786,I283778,I283645);
DFFARX1 I_16524 (I283786,I2859,I283418,I283386,);
nand I_16525 (I283817,I283778,I283687);
nand I_16526 (I283395,I283670,I283817);
not I_16527 (I283848,I283778);
nor I_16528 (I283865,I283848,I283588);
DFFARX1 I_16529 (I283865,I2859,I283418,I283407,);
nor I_16530 (I283896,I2388,I1652);
or I_16531 (I283398,I283645,I283896);
nor I_16532 (I283389,I283778,I283896);
or I_16533 (I283392,I283512,I283896);
DFFARX1 I_16534 (I283896,I2859,I283418,I283410,);
not I_16535 (I283996,I2866);
DFFARX1 I_16536 (I5255,I2859,I283996,I284022,);
not I_16537 (I284030,I284022);
nand I_16538 (I284047,I5258,I5270);
and I_16539 (I284064,I284047,I5249);
DFFARX1 I_16540 (I284064,I2859,I283996,I284090,);
not I_16541 (I284098,I5249);
DFFARX1 I_16542 (I5252,I2859,I283996,I284124,);
not I_16543 (I284132,I284124);
nor I_16544 (I284149,I284132,I284030);
and I_16545 (I284166,I284149,I5249);
nor I_16546 (I284183,I284132,I284098);
nor I_16547 (I283979,I284090,I284183);
DFFARX1 I_16548 (I5264,I2859,I283996,I284223,);
nor I_16549 (I284231,I284223,I284090);
not I_16550 (I284248,I284231);
not I_16551 (I284265,I284223);
nor I_16552 (I284282,I284265,I284166);
DFFARX1 I_16553 (I284282,I2859,I283996,I283982,);
nand I_16554 (I284313,I5267,I5252);
and I_16555 (I284330,I284313,I5261);
DFFARX1 I_16556 (I284330,I2859,I283996,I284356,);
nor I_16557 (I284364,I284356,I284223);
DFFARX1 I_16558 (I284364,I2859,I283996,I283964,);
nand I_16559 (I284395,I284356,I284265);
nand I_16560 (I283973,I284248,I284395);
not I_16561 (I284426,I284356);
nor I_16562 (I284443,I284426,I284166);
DFFARX1 I_16563 (I284443,I2859,I283996,I283985,);
nor I_16564 (I284474,I5255,I5252);
or I_16565 (I283976,I284223,I284474);
nor I_16566 (I283967,I284356,I284474);
or I_16567 (I283970,I284090,I284474);
DFFARX1 I_16568 (I284474,I2859,I283996,I283988,);
not I_16569 (I284574,I2866);
DFFARX1 I_16570 (I375397,I2859,I284574,I284600,);
not I_16571 (I284608,I284600);
nand I_16572 (I284625,I375373,I375388);
and I_16573 (I284642,I284625,I375400);
DFFARX1 I_16574 (I284642,I2859,I284574,I284668,);
not I_16575 (I284676,I375385);
DFFARX1 I_16576 (I375376,I2859,I284574,I284702,);
not I_16577 (I284710,I284702);
nor I_16578 (I284727,I284710,I284608);
and I_16579 (I284744,I284727,I375385);
nor I_16580 (I284761,I284710,I284676);
nor I_16581 (I284557,I284668,I284761);
DFFARX1 I_16582 (I375373,I2859,I284574,I284801,);
nor I_16583 (I284809,I284801,I284668);
not I_16584 (I284826,I284809);
not I_16585 (I284843,I284801);
nor I_16586 (I284860,I284843,I284744);
DFFARX1 I_16587 (I284860,I2859,I284574,I284560,);
nand I_16588 (I284891,I375391,I375382);
and I_16589 (I284908,I284891,I375394);
DFFARX1 I_16590 (I284908,I2859,I284574,I284934,);
nor I_16591 (I284942,I284934,I284801);
DFFARX1 I_16592 (I284942,I2859,I284574,I284542,);
nand I_16593 (I284973,I284934,I284843);
nand I_16594 (I284551,I284826,I284973);
not I_16595 (I285004,I284934);
nor I_16596 (I285021,I285004,I284744);
DFFARX1 I_16597 (I285021,I2859,I284574,I284563,);
nor I_16598 (I285052,I375379,I375382);
or I_16599 (I284554,I284801,I285052);
nor I_16600 (I284545,I284934,I285052);
or I_16601 (I284548,I284668,I285052);
DFFARX1 I_16602 (I285052,I2859,I284574,I284566,);
not I_16603 (I285152,I2866);
DFFARX1 I_16604 (I151473,I2859,I285152,I285178,);
not I_16605 (I285186,I285178);
nand I_16606 (I285203,I151476,I151452);
and I_16607 (I285220,I285203,I151449);
DFFARX1 I_16608 (I285220,I2859,I285152,I285246,);
not I_16609 (I285254,I151455);
DFFARX1 I_16610 (I151449,I2859,I285152,I285280,);
not I_16611 (I285288,I285280);
nor I_16612 (I285305,I285288,I285186);
and I_16613 (I285322,I285305,I151455);
nor I_16614 (I285339,I285288,I285254);
nor I_16615 (I285135,I285246,I285339);
DFFARX1 I_16616 (I151458,I2859,I285152,I285379,);
nor I_16617 (I285387,I285379,I285246);
not I_16618 (I285404,I285387);
not I_16619 (I285421,I285379);
nor I_16620 (I285438,I285421,I285322);
DFFARX1 I_16621 (I285438,I2859,I285152,I285138,);
nand I_16622 (I285469,I151461,I151470);
and I_16623 (I285486,I285469,I151467);
DFFARX1 I_16624 (I285486,I2859,I285152,I285512,);
nor I_16625 (I285520,I285512,I285379);
DFFARX1 I_16626 (I285520,I2859,I285152,I285120,);
nand I_16627 (I285551,I285512,I285421);
nand I_16628 (I285129,I285404,I285551);
not I_16629 (I285582,I285512);
nor I_16630 (I285599,I285582,I285322);
DFFARX1 I_16631 (I285599,I2859,I285152,I285141,);
nor I_16632 (I285630,I151464,I151470);
or I_16633 (I285132,I285379,I285630);
nor I_16634 (I285123,I285512,I285630);
or I_16635 (I285126,I285246,I285630);
DFFARX1 I_16636 (I285630,I2859,I285152,I285144,);
not I_16637 (I285730,I2866);
DFFARX1 I_16638 (I7964,I2859,I285730,I285756,);
not I_16639 (I285764,I285756);
nand I_16640 (I285781,I7961,I7952);
and I_16641 (I285798,I285781,I7952);
DFFARX1 I_16642 (I285798,I2859,I285730,I285824,);
not I_16643 (I285832,I7955);
DFFARX1 I_16644 (I7970,I2859,I285730,I285858,);
not I_16645 (I285866,I285858);
nor I_16646 (I285883,I285866,I285764);
and I_16647 (I285900,I285883,I7955);
nor I_16648 (I285917,I285866,I285832);
nor I_16649 (I285713,I285824,I285917);
DFFARX1 I_16650 (I7955,I2859,I285730,I285957,);
nor I_16651 (I285965,I285957,I285824);
not I_16652 (I285982,I285965);
not I_16653 (I285999,I285957);
nor I_16654 (I286016,I285999,I285900);
DFFARX1 I_16655 (I286016,I2859,I285730,I285716,);
nand I_16656 (I286047,I7973,I7958);
and I_16657 (I286064,I286047,I7976);
DFFARX1 I_16658 (I286064,I2859,I285730,I286090,);
nor I_16659 (I286098,I286090,I285957);
DFFARX1 I_16660 (I286098,I2859,I285730,I285698,);
nand I_16661 (I286129,I286090,I285999);
nand I_16662 (I285707,I285982,I286129);
not I_16663 (I286160,I286090);
nor I_16664 (I286177,I286160,I285900);
DFFARX1 I_16665 (I286177,I2859,I285730,I285719,);
nor I_16666 (I286208,I7967,I7958);
or I_16667 (I285710,I285957,I286208);
nor I_16668 (I285701,I286090,I286208);
or I_16669 (I285704,I285824,I286208);
DFFARX1 I_16670 (I286208,I2859,I285730,I285722,);
not I_16671 (I286308,I2866);
DFFARX1 I_16672 (I383795,I2859,I286308,I286334,);
not I_16673 (I286342,I286334);
nand I_16674 (I286359,I383771,I383786);
and I_16675 (I286376,I286359,I383798);
DFFARX1 I_16676 (I286376,I2859,I286308,I286402,);
not I_16677 (I286410,I383783);
DFFARX1 I_16678 (I383774,I2859,I286308,I286436,);
not I_16679 (I286444,I286436);
nor I_16680 (I286461,I286444,I286342);
and I_16681 (I286478,I286461,I383783);
nor I_16682 (I286495,I286444,I286410);
nor I_16683 (I286291,I286402,I286495);
DFFARX1 I_16684 (I383771,I2859,I286308,I286535,);
nor I_16685 (I286543,I286535,I286402);
not I_16686 (I286560,I286543);
not I_16687 (I286577,I286535);
nor I_16688 (I286594,I286577,I286478);
DFFARX1 I_16689 (I286594,I2859,I286308,I286294,);
nand I_16690 (I286625,I383789,I383780);
and I_16691 (I286642,I286625,I383792);
DFFARX1 I_16692 (I286642,I2859,I286308,I286668,);
nor I_16693 (I286676,I286668,I286535);
DFFARX1 I_16694 (I286676,I2859,I286308,I286276,);
nand I_16695 (I286707,I286668,I286577);
nand I_16696 (I286285,I286560,I286707);
not I_16697 (I286738,I286668);
nor I_16698 (I286755,I286738,I286478);
DFFARX1 I_16699 (I286755,I2859,I286308,I286297,);
nor I_16700 (I286786,I383777,I383780);
or I_16701 (I286288,I286535,I286786);
nor I_16702 (I286279,I286668,I286786);
or I_16703 (I286282,I286402,I286786);
DFFARX1 I_16704 (I286786,I2859,I286308,I286300,);
not I_16705 (I286886,I2866);
DFFARX1 I_16706 (I12180,I2859,I286886,I286912,);
not I_16707 (I286920,I286912);
nand I_16708 (I286937,I12177,I12168);
and I_16709 (I286954,I286937,I12168);
DFFARX1 I_16710 (I286954,I2859,I286886,I286980,);
not I_16711 (I286988,I12171);
DFFARX1 I_16712 (I12186,I2859,I286886,I287014,);
not I_16713 (I287022,I287014);
nor I_16714 (I287039,I287022,I286920);
and I_16715 (I287056,I287039,I12171);
nor I_16716 (I287073,I287022,I286988);
nor I_16717 (I286869,I286980,I287073);
DFFARX1 I_16718 (I12171,I2859,I286886,I287113,);
nor I_16719 (I287121,I287113,I286980);
not I_16720 (I287138,I287121);
not I_16721 (I287155,I287113);
nor I_16722 (I287172,I287155,I287056);
DFFARX1 I_16723 (I287172,I2859,I286886,I286872,);
nand I_16724 (I287203,I12189,I12174);
and I_16725 (I287220,I287203,I12192);
DFFARX1 I_16726 (I287220,I2859,I286886,I287246,);
nor I_16727 (I287254,I287246,I287113);
DFFARX1 I_16728 (I287254,I2859,I286886,I286854,);
nand I_16729 (I287285,I287246,I287155);
nand I_16730 (I286863,I287138,I287285);
not I_16731 (I287316,I287246);
nor I_16732 (I287333,I287316,I287056);
DFFARX1 I_16733 (I287333,I2859,I286886,I286875,);
nor I_16734 (I287364,I12183,I12174);
or I_16735 (I286866,I287113,I287364);
nor I_16736 (I286857,I287246,I287364);
or I_16737 (I286860,I286980,I287364);
DFFARX1 I_16738 (I287364,I2859,I286886,I286878,);
not I_16739 (I287464,I2866);
DFFARX1 I_16740 (I227320,I2859,I287464,I287490,);
not I_16741 (I287498,I287490);
nand I_16742 (I287515,I227329,I227338);
and I_16743 (I287532,I287515,I227344);
DFFARX1 I_16744 (I287532,I2859,I287464,I287558,);
not I_16745 (I287566,I227341);
DFFARX1 I_16746 (I227326,I2859,I287464,I287592,);
not I_16747 (I287600,I287592);
nor I_16748 (I287617,I287600,I287498);
and I_16749 (I287634,I287617,I227341);
nor I_16750 (I287651,I287600,I287566);
nor I_16751 (I287447,I287558,I287651);
DFFARX1 I_16752 (I227335,I2859,I287464,I287691,);
nor I_16753 (I287699,I287691,I287558);
not I_16754 (I287716,I287699);
not I_16755 (I287733,I287691);
nor I_16756 (I287750,I287733,I287634);
DFFARX1 I_16757 (I287750,I2859,I287464,I287450,);
nand I_16758 (I287781,I227332,I227323);
and I_16759 (I287798,I287781,I227320);
DFFARX1 I_16760 (I287798,I2859,I287464,I287824,);
nor I_16761 (I287832,I287824,I287691);
DFFARX1 I_16762 (I287832,I2859,I287464,I287432,);
nand I_16763 (I287863,I287824,I287733);
nand I_16764 (I287441,I287716,I287863);
not I_16765 (I287894,I287824);
nor I_16766 (I287911,I287894,I287634);
DFFARX1 I_16767 (I287911,I2859,I287464,I287453,);
nor I_16768 (I287942,I227323,I227323);
or I_16769 (I287444,I287691,I287942);
nor I_16770 (I287435,I287824,I287942);
or I_16771 (I287438,I287558,I287942);
DFFARX1 I_16772 (I287942,I2859,I287464,I287456,);
not I_16773 (I288042,I2866);
DFFARX1 I_16774 (I234834,I2859,I288042,I288068,);
not I_16775 (I288076,I288068);
nand I_16776 (I288093,I234843,I234852);
and I_16777 (I288110,I288093,I234858);
DFFARX1 I_16778 (I288110,I2859,I288042,I288136,);
not I_16779 (I288144,I234855);
DFFARX1 I_16780 (I234840,I2859,I288042,I288170,);
not I_16781 (I288178,I288170);
nor I_16782 (I288195,I288178,I288076);
and I_16783 (I288212,I288195,I234855);
nor I_16784 (I288229,I288178,I288144);
nor I_16785 (I288025,I288136,I288229);
DFFARX1 I_16786 (I234849,I2859,I288042,I288269,);
nor I_16787 (I288277,I288269,I288136);
not I_16788 (I288294,I288277);
not I_16789 (I288311,I288269);
nor I_16790 (I288328,I288311,I288212);
DFFARX1 I_16791 (I288328,I2859,I288042,I288028,);
nand I_16792 (I288359,I234846,I234837);
and I_16793 (I288376,I288359,I234834);
DFFARX1 I_16794 (I288376,I2859,I288042,I288402,);
nor I_16795 (I288410,I288402,I288269);
DFFARX1 I_16796 (I288410,I2859,I288042,I288010,);
nand I_16797 (I288441,I288402,I288311);
nand I_16798 (I288019,I288294,I288441);
not I_16799 (I288472,I288402);
nor I_16800 (I288489,I288472,I288212);
DFFARX1 I_16801 (I288489,I2859,I288042,I288031,);
nor I_16802 (I288520,I234837,I234837);
or I_16803 (I288022,I288269,I288520);
nor I_16804 (I288013,I288402,I288520);
or I_16805 (I288016,I288136,I288520);
DFFARX1 I_16806 (I288520,I2859,I288042,I288034,);
not I_16807 (I288620,I2866);
DFFARX1 I_16808 (I464352,I2859,I288620,I288646,);
not I_16809 (I288654,I288646);
nand I_16810 (I288671,I464334,I464346);
and I_16811 (I288688,I288671,I464349);
DFFARX1 I_16812 (I288688,I2859,I288620,I288714,);
not I_16813 (I288722,I464343);
DFFARX1 I_16814 (I464340,I2859,I288620,I288748,);
not I_16815 (I288756,I288748);
nor I_16816 (I288773,I288756,I288654);
and I_16817 (I288790,I288773,I464343);
nor I_16818 (I288807,I288756,I288722);
nor I_16819 (I288603,I288714,I288807);
DFFARX1 I_16820 (I464358,I2859,I288620,I288847,);
nor I_16821 (I288855,I288847,I288714);
not I_16822 (I288872,I288855);
not I_16823 (I288889,I288847);
nor I_16824 (I288906,I288889,I288790);
DFFARX1 I_16825 (I288906,I2859,I288620,I288606,);
nand I_16826 (I288937,I464337,I464337);
and I_16827 (I288954,I288937,I464334);
DFFARX1 I_16828 (I288954,I2859,I288620,I288980,);
nor I_16829 (I288988,I288980,I288847);
DFFARX1 I_16830 (I288988,I2859,I288620,I288588,);
nand I_16831 (I289019,I288980,I288889);
nand I_16832 (I288597,I288872,I289019);
not I_16833 (I289050,I288980);
nor I_16834 (I289067,I289050,I288790);
DFFARX1 I_16835 (I289067,I2859,I288620,I288609,);
nor I_16836 (I289098,I464355,I464337);
or I_16837 (I288600,I288847,I289098);
nor I_16838 (I288591,I288980,I289098);
or I_16839 (I288594,I288714,I289098);
DFFARX1 I_16840 (I289098,I2859,I288620,I288612,);
not I_16841 (I289198,I2866);
DFFARX1 I_16842 (I106637,I2859,I289198,I289224,);
not I_16843 (I289232,I289224);
nand I_16844 (I289249,I106640,I106661);
and I_16845 (I289266,I289249,I106649);
DFFARX1 I_16846 (I289266,I2859,I289198,I289292,);
not I_16847 (I289300,I106646);
DFFARX1 I_16848 (I106637,I2859,I289198,I289326,);
not I_16849 (I289334,I289326);
nor I_16850 (I289351,I289334,I289232);
and I_16851 (I289368,I289351,I106646);
nor I_16852 (I289385,I289334,I289300);
nor I_16853 (I289181,I289292,I289385);
DFFARX1 I_16854 (I106655,I2859,I289198,I289425,);
nor I_16855 (I289433,I289425,I289292);
not I_16856 (I289450,I289433);
not I_16857 (I289467,I289425);
nor I_16858 (I289484,I289467,I289368);
DFFARX1 I_16859 (I289484,I2859,I289198,I289184,);
nand I_16860 (I289515,I106640,I106643);
and I_16861 (I289532,I289515,I106652);
DFFARX1 I_16862 (I289532,I2859,I289198,I289558,);
nor I_16863 (I289566,I289558,I289425);
DFFARX1 I_16864 (I289566,I2859,I289198,I289166,);
nand I_16865 (I289597,I289558,I289467);
nand I_16866 (I289175,I289450,I289597);
not I_16867 (I289628,I289558);
nor I_16868 (I289645,I289628,I289368);
DFFARX1 I_16869 (I289645,I2859,I289198,I289187,);
nor I_16870 (I289676,I106658,I106643);
or I_16871 (I289178,I289425,I289676);
nor I_16872 (I289169,I289558,I289676);
or I_16873 (I289172,I289292,I289676);
DFFARX1 I_16874 (I289676,I2859,I289198,I289190,);
not I_16875 (I289776,I2866);
DFFARX1 I_16876 (I397361,I2859,I289776,I289802,);
not I_16877 (I289810,I289802);
nand I_16878 (I289827,I397337,I397352);
and I_16879 (I289844,I289827,I397364);
DFFARX1 I_16880 (I289844,I2859,I289776,I289870,);
not I_16881 (I289878,I397349);
DFFARX1 I_16882 (I397340,I2859,I289776,I289904,);
not I_16883 (I289912,I289904);
nor I_16884 (I289929,I289912,I289810);
and I_16885 (I289946,I289929,I397349);
nor I_16886 (I289963,I289912,I289878);
nor I_16887 (I289759,I289870,I289963);
DFFARX1 I_16888 (I397337,I2859,I289776,I290003,);
nor I_16889 (I290011,I290003,I289870);
not I_16890 (I290028,I290011);
not I_16891 (I290045,I290003);
nor I_16892 (I290062,I290045,I289946);
DFFARX1 I_16893 (I290062,I2859,I289776,I289762,);
nand I_16894 (I290093,I397355,I397346);
and I_16895 (I290110,I290093,I397358);
DFFARX1 I_16896 (I290110,I2859,I289776,I290136,);
nor I_16897 (I290144,I290136,I290003);
DFFARX1 I_16898 (I290144,I2859,I289776,I289744,);
nand I_16899 (I290175,I290136,I290045);
nand I_16900 (I289753,I290028,I290175);
not I_16901 (I290206,I290136);
nor I_16902 (I290223,I290206,I289946);
DFFARX1 I_16903 (I290223,I2859,I289776,I289765,);
nor I_16904 (I290254,I397343,I397346);
or I_16905 (I289756,I290003,I290254);
nor I_16906 (I289747,I290136,I290254);
or I_16907 (I289750,I289870,I290254);
DFFARX1 I_16908 (I290254,I2859,I289776,I289768,);
not I_16909 (I290354,I2866);
DFFARX1 I_16910 (I347066,I2859,I290354,I290380,);
not I_16911 (I290388,I290380);
nand I_16912 (I290405,I347054,I347072);
and I_16913 (I290422,I290405,I347069);
DFFARX1 I_16914 (I290422,I2859,I290354,I290448,);
not I_16915 (I290456,I347060);
DFFARX1 I_16916 (I347057,I2859,I290354,I290482,);
not I_16917 (I290490,I290482);
nor I_16918 (I290507,I290490,I290388);
and I_16919 (I290524,I290507,I347060);
nor I_16920 (I290541,I290490,I290456);
nor I_16921 (I290337,I290448,I290541);
DFFARX1 I_16922 (I347051,I2859,I290354,I290581,);
nor I_16923 (I290589,I290581,I290448);
not I_16924 (I290606,I290589);
not I_16925 (I290623,I290581);
nor I_16926 (I290640,I290623,I290524);
DFFARX1 I_16927 (I290640,I2859,I290354,I290340,);
nand I_16928 (I290671,I347051,I347054);
and I_16929 (I290688,I290671,I347057);
DFFARX1 I_16930 (I290688,I2859,I290354,I290714,);
nor I_16931 (I290722,I290714,I290581);
DFFARX1 I_16932 (I290722,I2859,I290354,I290322,);
nand I_16933 (I290753,I290714,I290623);
nand I_16934 (I290331,I290606,I290753);
not I_16935 (I290784,I290714);
nor I_16936 (I290801,I290784,I290524);
DFFARX1 I_16937 (I290801,I2859,I290354,I290343,);
nor I_16938 (I290832,I347063,I347054);
or I_16939 (I290334,I290581,I290832);
nor I_16940 (I290325,I290714,I290832);
or I_16941 (I290328,I290448,I290832);
DFFARX1 I_16942 (I290832,I2859,I290354,I290346,);
not I_16943 (I290932,I2866);
DFFARX1 I_16944 (I331256,I2859,I290932,I290958,);
not I_16945 (I290966,I290958);
nand I_16946 (I290983,I331244,I331262);
and I_16947 (I291000,I290983,I331259);
DFFARX1 I_16948 (I291000,I2859,I290932,I291026,);
not I_16949 (I291034,I331250);
DFFARX1 I_16950 (I331247,I2859,I290932,I291060,);
not I_16951 (I291068,I291060);
nor I_16952 (I291085,I291068,I290966);
and I_16953 (I291102,I291085,I331250);
nor I_16954 (I291119,I291068,I291034);
nor I_16955 (I290915,I291026,I291119);
DFFARX1 I_16956 (I331241,I2859,I290932,I291159,);
nor I_16957 (I291167,I291159,I291026);
not I_16958 (I291184,I291167);
not I_16959 (I291201,I291159);
nor I_16960 (I291218,I291201,I291102);
DFFARX1 I_16961 (I291218,I2859,I290932,I290918,);
nand I_16962 (I291249,I331241,I331244);
and I_16963 (I291266,I291249,I331247);
DFFARX1 I_16964 (I291266,I2859,I290932,I291292,);
nor I_16965 (I291300,I291292,I291159);
DFFARX1 I_16966 (I291300,I2859,I290932,I290900,);
nand I_16967 (I291331,I291292,I291201);
nand I_16968 (I290909,I291184,I291331);
not I_16969 (I291362,I291292);
nor I_16970 (I291379,I291362,I291102);
DFFARX1 I_16971 (I291379,I2859,I290932,I290921,);
nor I_16972 (I291410,I331253,I331244);
or I_16973 (I290912,I291159,I291410);
nor I_16974 (I290903,I291292,I291410);
or I_16975 (I290906,I291026,I291410);
DFFARX1 I_16976 (I291410,I2859,I290932,I290924,);
not I_16977 (I291510,I2866);
DFFARX1 I_16978 (I456260,I2859,I291510,I291536,);
not I_16979 (I291544,I291536);
nand I_16980 (I291561,I456242,I456254);
and I_16981 (I291578,I291561,I456257);
DFFARX1 I_16982 (I291578,I2859,I291510,I291604,);
not I_16983 (I291612,I456251);
DFFARX1 I_16984 (I456248,I2859,I291510,I291638,);
not I_16985 (I291646,I291638);
nor I_16986 (I291663,I291646,I291544);
and I_16987 (I291680,I291663,I456251);
nor I_16988 (I291697,I291646,I291612);
nor I_16989 (I291493,I291604,I291697);
DFFARX1 I_16990 (I456266,I2859,I291510,I291737,);
nor I_16991 (I291745,I291737,I291604);
not I_16992 (I291762,I291745);
not I_16993 (I291779,I291737);
nor I_16994 (I291796,I291779,I291680);
DFFARX1 I_16995 (I291796,I2859,I291510,I291496,);
nand I_16996 (I291827,I456245,I456245);
and I_16997 (I291844,I291827,I456242);
DFFARX1 I_16998 (I291844,I2859,I291510,I291870,);
nor I_16999 (I291878,I291870,I291737);
DFFARX1 I_17000 (I291878,I2859,I291510,I291478,);
nand I_17001 (I291909,I291870,I291779);
nand I_17002 (I291487,I291762,I291909);
not I_17003 (I291940,I291870);
nor I_17004 (I291957,I291940,I291680);
DFFARX1 I_17005 (I291957,I2859,I291510,I291499,);
nor I_17006 (I291988,I456263,I456245);
or I_17007 (I291490,I291737,I291988);
nor I_17008 (I291481,I291870,I291988);
or I_17009 (I291484,I291604,I291988);
DFFARX1 I_17010 (I291988,I2859,I291510,I291502,);
not I_17011 (I292088,I2866);
DFFARX1 I_17012 (I376043,I2859,I292088,I292114,);
not I_17013 (I292122,I292114);
nand I_17014 (I292139,I376019,I376034);
and I_17015 (I292156,I292139,I376046);
DFFARX1 I_17016 (I292156,I2859,I292088,I292182,);
not I_17017 (I292190,I376031);
DFFARX1 I_17018 (I376022,I2859,I292088,I292216,);
not I_17019 (I292224,I292216);
nor I_17020 (I292241,I292224,I292122);
and I_17021 (I292258,I292241,I376031);
nor I_17022 (I292275,I292224,I292190);
nor I_17023 (I292071,I292182,I292275);
DFFARX1 I_17024 (I376019,I2859,I292088,I292315,);
nor I_17025 (I292323,I292315,I292182);
not I_17026 (I292340,I292323);
not I_17027 (I292357,I292315);
nor I_17028 (I292374,I292357,I292258);
DFFARX1 I_17029 (I292374,I2859,I292088,I292074,);
nand I_17030 (I292405,I376037,I376028);
and I_17031 (I292422,I292405,I376040);
DFFARX1 I_17032 (I292422,I2859,I292088,I292448,);
nor I_17033 (I292456,I292448,I292315);
DFFARX1 I_17034 (I292456,I2859,I292088,I292056,);
nand I_17035 (I292487,I292448,I292357);
nand I_17036 (I292065,I292340,I292487);
not I_17037 (I292518,I292448);
nor I_17038 (I292535,I292518,I292258);
DFFARX1 I_17039 (I292535,I2859,I292088,I292077,);
nor I_17040 (I292566,I376025,I376028);
or I_17041 (I292068,I292315,I292566);
nor I_17042 (I292059,I292448,I292566);
or I_17043 (I292062,I292182,I292566);
DFFARX1 I_17044 (I292566,I2859,I292088,I292080,);
not I_17045 (I292666,I2866);
DFFARX1 I_17046 (I422078,I2859,I292666,I292692,);
not I_17047 (I292700,I292692);
nand I_17048 (I292717,I422075,I422093);
and I_17049 (I292734,I292717,I422090);
DFFARX1 I_17050 (I292734,I2859,I292666,I292760,);
not I_17051 (I292768,I422072);
DFFARX1 I_17052 (I422075,I2859,I292666,I292794,);
not I_17053 (I292802,I292794);
nor I_17054 (I292819,I292802,I292700);
and I_17055 (I292836,I292819,I422072);
nor I_17056 (I292853,I292802,I292768);
nor I_17057 (I292649,I292760,I292853);
DFFARX1 I_17058 (I422084,I2859,I292666,I292893,);
nor I_17059 (I292901,I292893,I292760);
not I_17060 (I292918,I292901);
not I_17061 (I292935,I292893);
nor I_17062 (I292952,I292935,I292836);
DFFARX1 I_17063 (I292952,I2859,I292666,I292652,);
nand I_17064 (I292983,I422087,I422072);
and I_17065 (I293000,I292983,I422078);
DFFARX1 I_17066 (I293000,I2859,I292666,I293026,);
nor I_17067 (I293034,I293026,I292893);
DFFARX1 I_17068 (I293034,I2859,I292666,I292634,);
nand I_17069 (I293065,I293026,I292935);
nand I_17070 (I292643,I292918,I293065);
not I_17071 (I293096,I293026);
nor I_17072 (I293113,I293096,I292836);
DFFARX1 I_17073 (I293113,I2859,I292666,I292655,);
nor I_17074 (I293144,I422081,I422072);
or I_17075 (I292646,I292893,I293144);
nor I_17076 (I292637,I293026,I293144);
or I_17077 (I292640,I292760,I293144);
DFFARX1 I_17078 (I293144,I2859,I292666,I292658,);
not I_17079 (I293244,I2866);
DFFARX1 I_17080 (I141987,I2859,I293244,I293270,);
not I_17081 (I293278,I293270);
nand I_17082 (I293295,I141990,I141966);
and I_17083 (I293312,I293295,I141963);
DFFARX1 I_17084 (I293312,I2859,I293244,I293338,);
not I_17085 (I293346,I141969);
DFFARX1 I_17086 (I141963,I2859,I293244,I293372,);
not I_17087 (I293380,I293372);
nor I_17088 (I293397,I293380,I293278);
and I_17089 (I293414,I293397,I141969);
nor I_17090 (I293431,I293380,I293346);
nor I_17091 (I293227,I293338,I293431);
DFFARX1 I_17092 (I141972,I2859,I293244,I293471,);
nor I_17093 (I293479,I293471,I293338);
not I_17094 (I293496,I293479);
not I_17095 (I293513,I293471);
nor I_17096 (I293530,I293513,I293414);
DFFARX1 I_17097 (I293530,I2859,I293244,I293230,);
nand I_17098 (I293561,I141975,I141984);
and I_17099 (I293578,I293561,I141981);
DFFARX1 I_17100 (I293578,I2859,I293244,I293604,);
nor I_17101 (I293612,I293604,I293471);
DFFARX1 I_17102 (I293612,I2859,I293244,I293212,);
nand I_17103 (I293643,I293604,I293513);
nand I_17104 (I293221,I293496,I293643);
not I_17105 (I293674,I293604);
nor I_17106 (I293691,I293674,I293414);
DFFARX1 I_17107 (I293691,I2859,I293244,I293233,);
nor I_17108 (I293722,I141978,I141984);
or I_17109 (I293224,I293471,I293722);
nor I_17110 (I293215,I293604,I293722);
or I_17111 (I293218,I293338,I293722);
DFFARX1 I_17112 (I293722,I2859,I293244,I293236,);
not I_17113 (I293822,I2866);
DFFARX1 I_17114 (I505746,I2859,I293822,I293848,);
not I_17115 (I293856,I293848);
nand I_17116 (I293873,I505749,I505758);
and I_17117 (I293890,I293873,I505761);
DFFARX1 I_17118 (I293890,I2859,I293822,I293916,);
not I_17119 (I293924,I505770);
DFFARX1 I_17120 (I505752,I2859,I293822,I293950,);
not I_17121 (I293958,I293950);
nor I_17122 (I293975,I293958,I293856);
and I_17123 (I293992,I293975,I505770);
nor I_17124 (I294009,I293958,I293924);
nor I_17125 (I293805,I293916,I294009);
DFFARX1 I_17126 (I505749,I2859,I293822,I294049,);
nor I_17127 (I294057,I294049,I293916);
not I_17128 (I294074,I294057);
not I_17129 (I294091,I294049);
nor I_17130 (I294108,I294091,I293992);
DFFARX1 I_17131 (I294108,I2859,I293822,I293808,);
nand I_17132 (I294139,I505767,I505746);
and I_17133 (I294156,I294139,I505764);
DFFARX1 I_17134 (I294156,I2859,I293822,I294182,);
nor I_17135 (I294190,I294182,I294049);
DFFARX1 I_17136 (I294190,I2859,I293822,I293790,);
nand I_17137 (I294221,I294182,I294091);
nand I_17138 (I293799,I294074,I294221);
not I_17139 (I294252,I294182);
nor I_17140 (I294269,I294252,I293992);
DFFARX1 I_17141 (I294269,I2859,I293822,I293811,);
nor I_17142 (I294300,I505755,I505746);
or I_17143 (I293802,I294049,I294300);
nor I_17144 (I293793,I294182,I294300);
or I_17145 (I293796,I293916,I294300);
DFFARX1 I_17146 (I294300,I2859,I293822,I293814,);
not I_17147 (I294400,I2866);
DFFARX1 I_17148 (I93547,I2859,I294400,I294426,);
not I_17149 (I294434,I294426);
nand I_17150 (I294451,I93550,I93571);
and I_17151 (I294468,I294451,I93559);
DFFARX1 I_17152 (I294468,I2859,I294400,I294494,);
not I_17153 (I294502,I93556);
DFFARX1 I_17154 (I93547,I2859,I294400,I294528,);
not I_17155 (I294536,I294528);
nor I_17156 (I294553,I294536,I294434);
and I_17157 (I294570,I294553,I93556);
nor I_17158 (I294587,I294536,I294502);
nor I_17159 (I294383,I294494,I294587);
DFFARX1 I_17160 (I93565,I2859,I294400,I294627,);
nor I_17161 (I294635,I294627,I294494);
not I_17162 (I294652,I294635);
not I_17163 (I294669,I294627);
nor I_17164 (I294686,I294669,I294570);
DFFARX1 I_17165 (I294686,I2859,I294400,I294386,);
nand I_17166 (I294717,I93550,I93553);
and I_17167 (I294734,I294717,I93562);
DFFARX1 I_17168 (I294734,I2859,I294400,I294760,);
nor I_17169 (I294768,I294760,I294627);
DFFARX1 I_17170 (I294768,I2859,I294400,I294368,);
nand I_17171 (I294799,I294760,I294669);
nand I_17172 (I294377,I294652,I294799);
not I_17173 (I294830,I294760);
nor I_17174 (I294847,I294830,I294570);
DFFARX1 I_17175 (I294847,I2859,I294400,I294389,);
nor I_17176 (I294878,I93568,I93553);
or I_17177 (I294380,I294627,I294878);
nor I_17178 (I294371,I294760,I294878);
or I_17179 (I294374,I294494,I294878);
DFFARX1 I_17180 (I294878,I2859,I294400,I294392,);
not I_17181 (I294978,I2866);
DFFARX1 I_17182 (I102472,I2859,I294978,I295004,);
not I_17183 (I295012,I295004);
nand I_17184 (I295029,I102475,I102496);
and I_17185 (I295046,I295029,I102484);
DFFARX1 I_17186 (I295046,I2859,I294978,I295072,);
not I_17187 (I295080,I102481);
DFFARX1 I_17188 (I102472,I2859,I294978,I295106,);
not I_17189 (I295114,I295106);
nor I_17190 (I295131,I295114,I295012);
and I_17191 (I295148,I295131,I102481);
nor I_17192 (I295165,I295114,I295080);
nor I_17193 (I294961,I295072,I295165);
DFFARX1 I_17194 (I102490,I2859,I294978,I295205,);
nor I_17195 (I295213,I295205,I295072);
not I_17196 (I295230,I295213);
not I_17197 (I295247,I295205);
nor I_17198 (I295264,I295247,I295148);
DFFARX1 I_17199 (I295264,I2859,I294978,I294964,);
nand I_17200 (I295295,I102475,I102478);
and I_17201 (I295312,I295295,I102487);
DFFARX1 I_17202 (I295312,I2859,I294978,I295338,);
nor I_17203 (I295346,I295338,I295205);
DFFARX1 I_17204 (I295346,I2859,I294978,I294946,);
nand I_17205 (I295377,I295338,I295247);
nand I_17206 (I294955,I295230,I295377);
not I_17207 (I295408,I295338);
nor I_17208 (I295425,I295408,I295148);
DFFARX1 I_17209 (I295425,I2859,I294978,I294967,);
nor I_17210 (I295456,I102493,I102478);
or I_17211 (I294958,I295205,I295456);
nor I_17212 (I294949,I295338,I295456);
or I_17213 (I294952,I295072,I295456);
DFFARX1 I_17214 (I295456,I2859,I294978,I294970,);
not I_17215 (I295556,I2866);
DFFARX1 I_17216 (I233678,I2859,I295556,I295582,);
not I_17217 (I295590,I295582);
nand I_17218 (I295607,I233687,I233696);
and I_17219 (I295624,I295607,I233702);
DFFARX1 I_17220 (I295624,I2859,I295556,I295650,);
not I_17221 (I295658,I233699);
DFFARX1 I_17222 (I233684,I2859,I295556,I295684,);
not I_17223 (I295692,I295684);
nor I_17224 (I295709,I295692,I295590);
and I_17225 (I295726,I295709,I233699);
nor I_17226 (I295743,I295692,I295658);
nor I_17227 (I295539,I295650,I295743);
DFFARX1 I_17228 (I233693,I2859,I295556,I295783,);
nor I_17229 (I295791,I295783,I295650);
not I_17230 (I295808,I295791);
not I_17231 (I295825,I295783);
nor I_17232 (I295842,I295825,I295726);
DFFARX1 I_17233 (I295842,I2859,I295556,I295542,);
nand I_17234 (I295873,I233690,I233681);
and I_17235 (I295890,I295873,I233678);
DFFARX1 I_17236 (I295890,I2859,I295556,I295916,);
nor I_17237 (I295924,I295916,I295783);
DFFARX1 I_17238 (I295924,I2859,I295556,I295524,);
nand I_17239 (I295955,I295916,I295825);
nand I_17240 (I295533,I295808,I295955);
not I_17241 (I295986,I295916);
nor I_17242 (I296003,I295986,I295726);
DFFARX1 I_17243 (I296003,I2859,I295556,I295545,);
nor I_17244 (I296034,I233681,I233681);
or I_17245 (I295536,I295783,I296034);
nor I_17246 (I295527,I295916,I296034);
or I_17247 (I295530,I295650,I296034);
DFFARX1 I_17248 (I296034,I2859,I295556,I295548,);
not I_17249 (I296134,I2866);
DFFARX1 I_17250 (I557062,I2859,I296134,I296160,);
not I_17251 (I296168,I296160);
nand I_17252 (I296185,I557047,I557035);
and I_17253 (I296202,I296185,I557050);
DFFARX1 I_17254 (I296202,I2859,I296134,I296228,);
not I_17255 (I296236,I557035);
DFFARX1 I_17256 (I557053,I2859,I296134,I296262,);
not I_17257 (I296270,I296262);
nor I_17258 (I296287,I296270,I296168);
and I_17259 (I296304,I296287,I557035);
nor I_17260 (I296321,I296270,I296236);
nor I_17261 (I296117,I296228,I296321);
DFFARX1 I_17262 (I557041,I2859,I296134,I296361,);
nor I_17263 (I296369,I296361,I296228);
not I_17264 (I296386,I296369);
not I_17265 (I296403,I296361);
nor I_17266 (I296420,I296403,I296304);
DFFARX1 I_17267 (I296420,I2859,I296134,I296120,);
nand I_17268 (I296451,I557038,I557044);
and I_17269 (I296468,I296451,I557059);
DFFARX1 I_17270 (I296468,I2859,I296134,I296494,);
nor I_17271 (I296502,I296494,I296361);
DFFARX1 I_17272 (I296502,I2859,I296134,I296102,);
nand I_17273 (I296533,I296494,I296403);
nand I_17274 (I296111,I296386,I296533);
not I_17275 (I296564,I296494);
nor I_17276 (I296581,I296564,I296304);
DFFARX1 I_17277 (I296581,I2859,I296134,I296123,);
nor I_17278 (I296612,I557056,I557044);
or I_17279 (I296114,I296361,I296612);
nor I_17280 (I296105,I296494,I296612);
or I_17281 (I296108,I296228,I296612);
DFFARX1 I_17282 (I296612,I2859,I296134,I296126,);
not I_17283 (I296712,I2866);
DFFARX1 I_17284 (I424322,I2859,I296712,I296738,);
not I_17285 (I296746,I296738);
nand I_17286 (I296763,I424319,I424337);
and I_17287 (I296780,I296763,I424334);
DFFARX1 I_17288 (I296780,I2859,I296712,I296806,);
not I_17289 (I296814,I424316);
DFFARX1 I_17290 (I424319,I2859,I296712,I296840,);
not I_17291 (I296848,I296840);
nor I_17292 (I296865,I296848,I296746);
and I_17293 (I296882,I296865,I424316);
nor I_17294 (I296899,I296848,I296814);
nor I_17295 (I296695,I296806,I296899);
DFFARX1 I_17296 (I424328,I2859,I296712,I296939,);
nor I_17297 (I296947,I296939,I296806);
not I_17298 (I296964,I296947);
not I_17299 (I296981,I296939);
nor I_17300 (I296998,I296981,I296882);
DFFARX1 I_17301 (I296998,I2859,I296712,I296698,);
nand I_17302 (I297029,I424331,I424316);
and I_17303 (I297046,I297029,I424322);
DFFARX1 I_17304 (I297046,I2859,I296712,I297072,);
nor I_17305 (I297080,I297072,I296939);
DFFARX1 I_17306 (I297080,I2859,I296712,I296680,);
nand I_17307 (I297111,I297072,I296981);
nand I_17308 (I296689,I296964,I297111);
not I_17309 (I297142,I297072);
nor I_17310 (I297159,I297142,I296882);
DFFARX1 I_17311 (I297159,I2859,I296712,I296701,);
nor I_17312 (I297190,I424325,I424316);
or I_17313 (I296692,I296939,I297190);
nor I_17314 (I296683,I297072,I297190);
or I_17315 (I296686,I296806,I297190);
DFFARX1 I_17316 (I297190,I2859,I296712,I296704,);
not I_17317 (I297290,I2866);
DFFARX1 I_17318 (I340215,I2859,I297290,I297316,);
not I_17319 (I297324,I297316);
nand I_17320 (I297341,I340203,I340221);
and I_17321 (I297358,I297341,I340218);
DFFARX1 I_17322 (I297358,I2859,I297290,I297384,);
not I_17323 (I297392,I340209);
DFFARX1 I_17324 (I340206,I2859,I297290,I297418,);
not I_17325 (I297426,I297418);
nor I_17326 (I297443,I297426,I297324);
and I_17327 (I297460,I297443,I340209);
nor I_17328 (I297477,I297426,I297392);
nor I_17329 (I297273,I297384,I297477);
DFFARX1 I_17330 (I340200,I2859,I297290,I297517,);
nor I_17331 (I297525,I297517,I297384);
not I_17332 (I297542,I297525);
not I_17333 (I297559,I297517);
nor I_17334 (I297576,I297559,I297460);
DFFARX1 I_17335 (I297576,I2859,I297290,I297276,);
nand I_17336 (I297607,I340200,I340203);
and I_17337 (I297624,I297607,I340206);
DFFARX1 I_17338 (I297624,I2859,I297290,I297650,);
nor I_17339 (I297658,I297650,I297517);
DFFARX1 I_17340 (I297658,I2859,I297290,I297258,);
nand I_17341 (I297689,I297650,I297559);
nand I_17342 (I297267,I297542,I297689);
not I_17343 (I297720,I297650);
nor I_17344 (I297737,I297720,I297460);
DFFARX1 I_17345 (I297737,I2859,I297290,I297279,);
nor I_17346 (I297768,I340212,I340203);
or I_17347 (I297270,I297517,I297768);
nor I_17348 (I297261,I297650,I297768);
or I_17349 (I297264,I297384,I297768);
DFFARX1 I_17350 (I297768,I2859,I297290,I297282,);
not I_17351 (I297868,I2866);
DFFARX1 I_17352 (I180001,I2859,I297868,I297894,);
not I_17353 (I297902,I297894);
nand I_17354 (I297919,I179992,I180010);
and I_17355 (I297936,I297919,I180013);
DFFARX1 I_17356 (I297936,I2859,I297868,I297962,);
not I_17357 (I297970,I180007);
DFFARX1 I_17358 (I179995,I2859,I297868,I297996,);
not I_17359 (I298004,I297996);
nor I_17360 (I298021,I298004,I297902);
and I_17361 (I298038,I298021,I180007);
nor I_17362 (I298055,I298004,I297970);
nor I_17363 (I297851,I297962,I298055);
DFFARX1 I_17364 (I180004,I2859,I297868,I298095,);
nor I_17365 (I298103,I298095,I297962);
not I_17366 (I298120,I298103);
not I_17367 (I298137,I298095);
nor I_17368 (I298154,I298137,I298038);
DFFARX1 I_17369 (I298154,I2859,I297868,I297854,);
nand I_17370 (I298185,I180019,I180016);
and I_17371 (I298202,I298185,I179998);
DFFARX1 I_17372 (I298202,I2859,I297868,I298228,);
nor I_17373 (I298236,I298228,I298095);
DFFARX1 I_17374 (I298236,I2859,I297868,I297836,);
nand I_17375 (I298267,I298228,I298137);
nand I_17376 (I297845,I298120,I298267);
not I_17377 (I298298,I298228);
nor I_17378 (I298315,I298298,I298038);
DFFARX1 I_17379 (I298315,I2859,I297868,I297857,);
nor I_17380 (I298346,I179992,I180016);
or I_17381 (I297848,I298095,I298346);
nor I_17382 (I297839,I298228,I298346);
or I_17383 (I297842,I297962,I298346);
DFFARX1 I_17384 (I298346,I2859,I297868,I297860,);
not I_17385 (I298446,I2866);
DFFARX1 I_17386 (I241770,I2859,I298446,I298472,);
not I_17387 (I298480,I298472);
nand I_17388 (I298497,I241779,I241788);
and I_17389 (I298514,I298497,I241794);
DFFARX1 I_17390 (I298514,I2859,I298446,I298540,);
not I_17391 (I298548,I241791);
DFFARX1 I_17392 (I241776,I2859,I298446,I298574,);
not I_17393 (I298582,I298574);
nor I_17394 (I298599,I298582,I298480);
and I_17395 (I298616,I298599,I241791);
nor I_17396 (I298633,I298582,I298548);
nor I_17397 (I298429,I298540,I298633);
DFFARX1 I_17398 (I241785,I2859,I298446,I298673,);
nor I_17399 (I298681,I298673,I298540);
not I_17400 (I298698,I298681);
not I_17401 (I298715,I298673);
nor I_17402 (I298732,I298715,I298616);
DFFARX1 I_17403 (I298732,I2859,I298446,I298432,);
nand I_17404 (I298763,I241782,I241773);
and I_17405 (I298780,I298763,I241770);
DFFARX1 I_17406 (I298780,I2859,I298446,I298806,);
nor I_17407 (I298814,I298806,I298673);
DFFARX1 I_17408 (I298814,I2859,I298446,I298414,);
nand I_17409 (I298845,I298806,I298715);
nand I_17410 (I298423,I298698,I298845);
not I_17411 (I298876,I298806);
nor I_17412 (I298893,I298876,I298616);
DFFARX1 I_17413 (I298893,I2859,I298446,I298435,);
nor I_17414 (I298924,I241773,I241773);
or I_17415 (I298426,I298673,I298924);
nor I_17416 (I298417,I298806,I298924);
or I_17417 (I298420,I298540,I298924);
DFFARX1 I_17418 (I298924,I2859,I298446,I298438,);
not I_17419 (I299024,I2866);
DFFARX1 I_17420 (I248706,I2859,I299024,I299050,);
not I_17421 (I299058,I299050);
nand I_17422 (I299075,I248715,I248724);
and I_17423 (I299092,I299075,I248730);
DFFARX1 I_17424 (I299092,I2859,I299024,I299118,);
not I_17425 (I299126,I248727);
DFFARX1 I_17426 (I248712,I2859,I299024,I299152,);
not I_17427 (I299160,I299152);
nor I_17428 (I299177,I299160,I299058);
and I_17429 (I299194,I299177,I248727);
nor I_17430 (I299211,I299160,I299126);
nor I_17431 (I299007,I299118,I299211);
DFFARX1 I_17432 (I248721,I2859,I299024,I299251,);
nor I_17433 (I299259,I299251,I299118);
not I_17434 (I299276,I299259);
not I_17435 (I299293,I299251);
nor I_17436 (I299310,I299293,I299194);
DFFARX1 I_17437 (I299310,I2859,I299024,I299010,);
nand I_17438 (I299341,I248718,I248709);
and I_17439 (I299358,I299341,I248706);
DFFARX1 I_17440 (I299358,I2859,I299024,I299384,);
nor I_17441 (I299392,I299384,I299251);
DFFARX1 I_17442 (I299392,I2859,I299024,I298992,);
nand I_17443 (I299423,I299384,I299293);
nand I_17444 (I299001,I299276,I299423);
not I_17445 (I299454,I299384);
nor I_17446 (I299471,I299454,I299194);
DFFARX1 I_17447 (I299471,I2859,I299024,I299013,);
nor I_17448 (I299502,I248709,I248709);
or I_17449 (I299004,I299251,I299502);
nor I_17450 (I298995,I299384,I299502);
or I_17451 (I298998,I299118,I299502);
DFFARX1 I_17452 (I299502,I2859,I299024,I299016,);
not I_17453 (I299602,I2866);
DFFARX1 I_17454 (I559442,I2859,I299602,I299628,);
not I_17455 (I299636,I299628);
nand I_17456 (I299653,I559427,I559415);
and I_17457 (I299670,I299653,I559430);
DFFARX1 I_17458 (I299670,I2859,I299602,I299696,);
not I_17459 (I299704,I559415);
DFFARX1 I_17460 (I559433,I2859,I299602,I299730,);
not I_17461 (I299738,I299730);
nor I_17462 (I299755,I299738,I299636);
and I_17463 (I299772,I299755,I559415);
nor I_17464 (I299789,I299738,I299704);
nor I_17465 (I299585,I299696,I299789);
DFFARX1 I_17466 (I559421,I2859,I299602,I299829,);
nor I_17467 (I299837,I299829,I299696);
not I_17468 (I299854,I299837);
not I_17469 (I299871,I299829);
nor I_17470 (I299888,I299871,I299772);
DFFARX1 I_17471 (I299888,I2859,I299602,I299588,);
nand I_17472 (I299919,I559418,I559424);
and I_17473 (I299936,I299919,I559439);
DFFARX1 I_17474 (I299936,I2859,I299602,I299962,);
nor I_17475 (I299970,I299962,I299829);
DFFARX1 I_17476 (I299970,I2859,I299602,I299570,);
nand I_17477 (I300001,I299962,I299871);
nand I_17478 (I299579,I299854,I300001);
not I_17479 (I300032,I299962);
nor I_17480 (I300049,I300032,I299772);
DFFARX1 I_17481 (I300049,I2859,I299602,I299591,);
nor I_17482 (I300080,I559436,I559424);
or I_17483 (I299582,I299829,I300080);
nor I_17484 (I299573,I299962,I300080);
or I_17485 (I299576,I299696,I300080);
DFFARX1 I_17486 (I300080,I2859,I299602,I299594,);
not I_17487 (I300180,I2866);
DFFARX1 I_17488 (I135663,I2859,I300180,I300206,);
not I_17489 (I300214,I300206);
nand I_17490 (I300231,I135666,I135642);
and I_17491 (I300248,I300231,I135639);
DFFARX1 I_17492 (I300248,I2859,I300180,I300274,);
not I_17493 (I300282,I135645);
DFFARX1 I_17494 (I135639,I2859,I300180,I300308,);
not I_17495 (I300316,I300308);
nor I_17496 (I300333,I300316,I300214);
and I_17497 (I300350,I300333,I135645);
nor I_17498 (I300367,I300316,I300282);
nor I_17499 (I300163,I300274,I300367);
DFFARX1 I_17500 (I135648,I2859,I300180,I300407,);
nor I_17501 (I300415,I300407,I300274);
not I_17502 (I300432,I300415);
not I_17503 (I300449,I300407);
nor I_17504 (I300466,I300449,I300350);
DFFARX1 I_17505 (I300466,I2859,I300180,I300166,);
nand I_17506 (I300497,I135651,I135660);
and I_17507 (I300514,I300497,I135657);
DFFARX1 I_17508 (I300514,I2859,I300180,I300540,);
nor I_17509 (I300548,I300540,I300407);
DFFARX1 I_17510 (I300548,I2859,I300180,I300148,);
nand I_17511 (I300579,I300540,I300449);
nand I_17512 (I300157,I300432,I300579);
not I_17513 (I300610,I300540);
nor I_17514 (I300627,I300610,I300350);
DFFARX1 I_17515 (I300627,I2859,I300180,I300169,);
nor I_17516 (I300658,I135654,I135660);
or I_17517 (I300160,I300407,I300658);
nor I_17518 (I300151,I300540,I300658);
or I_17519 (I300154,I300274,I300658);
DFFARX1 I_17520 (I300658,I2859,I300180,I300172,);
not I_17521 (I300758,I2866);
DFFARX1 I_17522 (I334945,I2859,I300758,I300784,);
not I_17523 (I300792,I300784);
nand I_17524 (I300809,I334933,I334951);
and I_17525 (I300826,I300809,I334948);
DFFARX1 I_17526 (I300826,I2859,I300758,I300852,);
not I_17527 (I300860,I334939);
DFFARX1 I_17528 (I334936,I2859,I300758,I300886,);
not I_17529 (I300894,I300886);
nor I_17530 (I300911,I300894,I300792);
and I_17531 (I300928,I300911,I334939);
nor I_17532 (I300945,I300894,I300860);
nor I_17533 (I300741,I300852,I300945);
DFFARX1 I_17534 (I334930,I2859,I300758,I300985,);
nor I_17535 (I300993,I300985,I300852);
not I_17536 (I301010,I300993);
not I_17537 (I301027,I300985);
nor I_17538 (I301044,I301027,I300928);
DFFARX1 I_17539 (I301044,I2859,I300758,I300744,);
nand I_17540 (I301075,I334930,I334933);
and I_17541 (I301092,I301075,I334936);
DFFARX1 I_17542 (I301092,I2859,I300758,I301118,);
nor I_17543 (I301126,I301118,I300985);
DFFARX1 I_17544 (I301126,I2859,I300758,I300726,);
nand I_17545 (I301157,I301118,I301027);
nand I_17546 (I300735,I301010,I301157);
not I_17547 (I301188,I301118);
nor I_17548 (I301205,I301188,I300928);
DFFARX1 I_17549 (I301205,I2859,I300758,I300747,);
nor I_17550 (I301236,I334942,I334933);
or I_17551 (I300738,I300985,I301236);
nor I_17552 (I300729,I301118,I301236);
or I_17553 (I300732,I300852,I301236);
DFFARX1 I_17554 (I301236,I2859,I300758,I300750,);
not I_17555 (I301336,I2866);
DFFARX1 I_17556 (I110207,I2859,I301336,I301362,);
not I_17557 (I301370,I301362);
nand I_17558 (I301387,I110210,I110231);
and I_17559 (I301404,I301387,I110219);
DFFARX1 I_17560 (I301404,I2859,I301336,I301430,);
not I_17561 (I301438,I110216);
DFFARX1 I_17562 (I110207,I2859,I301336,I301464,);
not I_17563 (I301472,I301464);
nor I_17564 (I301489,I301472,I301370);
and I_17565 (I301506,I301489,I110216);
nor I_17566 (I301523,I301472,I301438);
nor I_17567 (I301319,I301430,I301523);
DFFARX1 I_17568 (I110225,I2859,I301336,I301563,);
nor I_17569 (I301571,I301563,I301430);
not I_17570 (I301588,I301571);
not I_17571 (I301605,I301563);
nor I_17572 (I301622,I301605,I301506);
DFFARX1 I_17573 (I301622,I2859,I301336,I301322,);
nand I_17574 (I301653,I110210,I110213);
and I_17575 (I301670,I301653,I110222);
DFFARX1 I_17576 (I301670,I2859,I301336,I301696,);
nor I_17577 (I301704,I301696,I301563);
DFFARX1 I_17578 (I301704,I2859,I301336,I301304,);
nand I_17579 (I301735,I301696,I301605);
nand I_17580 (I301313,I301588,I301735);
not I_17581 (I301766,I301696);
nor I_17582 (I301783,I301766,I301506);
DFFARX1 I_17583 (I301783,I2859,I301336,I301325,);
nor I_17584 (I301814,I110228,I110213);
or I_17585 (I301316,I301563,I301814);
nor I_17586 (I301307,I301696,I301814);
or I_17587 (I301310,I301430,I301814);
DFFARX1 I_17588 (I301814,I2859,I301336,I301328,);
not I_17589 (I301914,I2866);
DFFARX1 I_17590 (I195233,I2859,I301914,I301940,);
not I_17591 (I301948,I301940);
nand I_17592 (I301965,I195224,I195242);
and I_17593 (I301982,I301965,I195245);
DFFARX1 I_17594 (I301982,I2859,I301914,I302008,);
not I_17595 (I302016,I195239);
DFFARX1 I_17596 (I195227,I2859,I301914,I302042,);
not I_17597 (I302050,I302042);
nor I_17598 (I302067,I302050,I301948);
and I_17599 (I302084,I302067,I195239);
nor I_17600 (I302101,I302050,I302016);
nor I_17601 (I301897,I302008,I302101);
DFFARX1 I_17602 (I195236,I2859,I301914,I302141,);
nor I_17603 (I302149,I302141,I302008);
not I_17604 (I302166,I302149);
not I_17605 (I302183,I302141);
nor I_17606 (I302200,I302183,I302084);
DFFARX1 I_17607 (I302200,I2859,I301914,I301900,);
nand I_17608 (I302231,I195251,I195248);
and I_17609 (I302248,I302231,I195230);
DFFARX1 I_17610 (I302248,I2859,I301914,I302274,);
nor I_17611 (I302282,I302274,I302141);
DFFARX1 I_17612 (I302282,I2859,I301914,I301882,);
nand I_17613 (I302313,I302274,I302183);
nand I_17614 (I301891,I302166,I302313);
not I_17615 (I302344,I302274);
nor I_17616 (I302361,I302344,I302084);
DFFARX1 I_17617 (I302361,I2859,I301914,I301903,);
nor I_17618 (I302392,I195224,I195248);
or I_17619 (I301894,I302141,I302392);
nor I_17620 (I301885,I302274,I302392);
or I_17621 (I301888,I302008,I302392);
DFFARX1 I_17622 (I302392,I2859,I301914,I301906,);
not I_17623 (I302492,I2866);
DFFARX1 I_17624 (I52504,I2859,I302492,I302518,);
not I_17625 (I302526,I302518);
nand I_17626 (I302543,I52519,I52492);
and I_17627 (I302560,I302543,I52507);
DFFARX1 I_17628 (I302560,I2859,I302492,I302586,);
not I_17629 (I302594,I52510);
DFFARX1 I_17630 (I52495,I2859,I302492,I302620,);
not I_17631 (I302628,I302620);
nor I_17632 (I302645,I302628,I302526);
and I_17633 (I302662,I302645,I52510);
nor I_17634 (I302679,I302628,I302594);
nor I_17635 (I302475,I302586,I302679);
DFFARX1 I_17636 (I52501,I2859,I302492,I302719,);
nor I_17637 (I302727,I302719,I302586);
not I_17638 (I302744,I302727);
not I_17639 (I302761,I302719);
nor I_17640 (I302778,I302761,I302662);
DFFARX1 I_17641 (I302778,I2859,I302492,I302478,);
nand I_17642 (I302809,I52516,I52498);
and I_17643 (I302826,I302809,I52513);
DFFARX1 I_17644 (I302826,I2859,I302492,I302852,);
nor I_17645 (I302860,I302852,I302719);
DFFARX1 I_17646 (I302860,I2859,I302492,I302460,);
nand I_17647 (I302891,I302852,I302761);
nand I_17648 (I302469,I302744,I302891);
not I_17649 (I302922,I302852);
nor I_17650 (I302939,I302922,I302662);
DFFARX1 I_17651 (I302939,I2859,I302492,I302481,);
nor I_17652 (I302970,I52492,I52498);
or I_17653 (I302472,I302719,I302970);
nor I_17654 (I302463,I302852,I302970);
or I_17655 (I302466,I302586,I302970);
DFFARX1 I_17656 (I302970,I2859,I302492,I302484,);
not I_17657 (I303070,I2866);
DFFARX1 I_17658 (I422639,I2859,I303070,I303096,);
not I_17659 (I303104,I303096);
nand I_17660 (I303121,I422636,I422654);
and I_17661 (I303138,I303121,I422651);
DFFARX1 I_17662 (I303138,I2859,I303070,I303164,);
not I_17663 (I303172,I422633);
DFFARX1 I_17664 (I422636,I2859,I303070,I303198,);
not I_17665 (I303206,I303198);
nor I_17666 (I303223,I303206,I303104);
and I_17667 (I303240,I303223,I422633);
nor I_17668 (I303257,I303206,I303172);
nor I_17669 (I303053,I303164,I303257);
DFFARX1 I_17670 (I422645,I2859,I303070,I303297,);
nor I_17671 (I303305,I303297,I303164);
not I_17672 (I303322,I303305);
not I_17673 (I303339,I303297);
nor I_17674 (I303356,I303339,I303240);
DFFARX1 I_17675 (I303356,I2859,I303070,I303056,);
nand I_17676 (I303387,I422648,I422633);
and I_17677 (I303404,I303387,I422639);
DFFARX1 I_17678 (I303404,I2859,I303070,I303430,);
nor I_17679 (I303438,I303430,I303297);
DFFARX1 I_17680 (I303438,I2859,I303070,I303038,);
nand I_17681 (I303469,I303430,I303339);
nand I_17682 (I303047,I303322,I303469);
not I_17683 (I303500,I303430);
nor I_17684 (I303517,I303500,I303240);
DFFARX1 I_17685 (I303517,I2859,I303070,I303059,);
nor I_17686 (I303548,I422642,I422633);
or I_17687 (I303050,I303297,I303548);
nor I_17688 (I303041,I303430,I303548);
or I_17689 (I303044,I303164,I303548);
DFFARX1 I_17690 (I303548,I2859,I303070,I303062,);
not I_17691 (I303648,I2866);
DFFARX1 I_17692 (I386379,I2859,I303648,I303674,);
not I_17693 (I303682,I303674);
nand I_17694 (I303699,I386355,I386370);
and I_17695 (I303716,I303699,I386382);
DFFARX1 I_17696 (I303716,I2859,I303648,I303742,);
not I_17697 (I303750,I386367);
DFFARX1 I_17698 (I386358,I2859,I303648,I303776,);
not I_17699 (I303784,I303776);
nor I_17700 (I303801,I303784,I303682);
and I_17701 (I303818,I303801,I386367);
nor I_17702 (I303835,I303784,I303750);
nor I_17703 (I303631,I303742,I303835);
DFFARX1 I_17704 (I386355,I2859,I303648,I303875,);
nor I_17705 (I303883,I303875,I303742);
not I_17706 (I303900,I303883);
not I_17707 (I303917,I303875);
nor I_17708 (I303934,I303917,I303818);
DFFARX1 I_17709 (I303934,I2859,I303648,I303634,);
nand I_17710 (I303965,I386373,I386364);
and I_17711 (I303982,I303965,I386376);
DFFARX1 I_17712 (I303982,I2859,I303648,I304008,);
nor I_17713 (I304016,I304008,I303875);
DFFARX1 I_17714 (I304016,I2859,I303648,I303616,);
nand I_17715 (I304047,I304008,I303917);
nand I_17716 (I303625,I303900,I304047);
not I_17717 (I304078,I304008);
nor I_17718 (I304095,I304078,I303818);
DFFARX1 I_17719 (I304095,I2859,I303648,I303637,);
nor I_17720 (I304126,I386361,I386364);
or I_17721 (I303628,I303875,I304126);
nor I_17722 (I303619,I304008,I304126);
or I_17723 (I303622,I303742,I304126);
DFFARX1 I_17724 (I304126,I2859,I303648,I303640,);
not I_17725 (I304226,I2866);
DFFARX1 I_17726 (I25346,I2859,I304226,I304252,);
not I_17727 (I304260,I304252);
nand I_17728 (I304277,I25355,I25364);
and I_17729 (I304294,I304277,I25343);
DFFARX1 I_17730 (I304294,I2859,I304226,I304320,);
not I_17731 (I304328,I25346);
DFFARX1 I_17732 (I25361,I2859,I304226,I304354,);
not I_17733 (I304362,I304354);
nor I_17734 (I304379,I304362,I304260);
and I_17735 (I304396,I304379,I25346);
nor I_17736 (I304413,I304362,I304328);
nor I_17737 (I304209,I304320,I304413);
DFFARX1 I_17738 (I25352,I2859,I304226,I304453,);
nor I_17739 (I304461,I304453,I304320);
not I_17740 (I304478,I304461);
not I_17741 (I304495,I304453);
nor I_17742 (I304512,I304495,I304396);
DFFARX1 I_17743 (I304512,I2859,I304226,I304212,);
nand I_17744 (I304543,I25367,I25343);
and I_17745 (I304560,I304543,I25349);
DFFARX1 I_17746 (I304560,I2859,I304226,I304586,);
nor I_17747 (I304594,I304586,I304453);
DFFARX1 I_17748 (I304594,I2859,I304226,I304194,);
nand I_17749 (I304625,I304586,I304495);
nand I_17750 (I304203,I304478,I304625);
not I_17751 (I304656,I304586);
nor I_17752 (I304673,I304656,I304396);
DFFARX1 I_17753 (I304673,I2859,I304226,I304215,);
nor I_17754 (I304704,I25358,I25343);
or I_17755 (I304206,I304453,I304704);
nor I_17756 (I304197,I304586,I304704);
or I_17757 (I304200,I304320,I304704);
DFFARX1 I_17758 (I304704,I2859,I304226,I304218,);
not I_17759 (I304804,I2866);
DFFARX1 I_17760 (I449902,I2859,I304804,I304830,);
not I_17761 (I304838,I304830);
nand I_17762 (I304855,I449884,I449896);
and I_17763 (I304872,I304855,I449899);
DFFARX1 I_17764 (I304872,I2859,I304804,I304898,);
not I_17765 (I304906,I449893);
DFFARX1 I_17766 (I449890,I2859,I304804,I304932,);
not I_17767 (I304940,I304932);
nor I_17768 (I304957,I304940,I304838);
and I_17769 (I304974,I304957,I449893);
nor I_17770 (I304991,I304940,I304906);
nor I_17771 (I304787,I304898,I304991);
DFFARX1 I_17772 (I449908,I2859,I304804,I305031,);
nor I_17773 (I305039,I305031,I304898);
not I_17774 (I305056,I305039);
not I_17775 (I305073,I305031);
nor I_17776 (I305090,I305073,I304974);
DFFARX1 I_17777 (I305090,I2859,I304804,I304790,);
nand I_17778 (I305121,I449887,I449887);
and I_17779 (I305138,I305121,I449884);
DFFARX1 I_17780 (I305138,I2859,I304804,I305164,);
nor I_17781 (I305172,I305164,I305031);
DFFARX1 I_17782 (I305172,I2859,I304804,I304772,);
nand I_17783 (I305203,I305164,I305073);
nand I_17784 (I304781,I305056,I305203);
not I_17785 (I305234,I305164);
nor I_17786 (I305251,I305234,I304974);
DFFARX1 I_17787 (I305251,I2859,I304804,I304793,);
nor I_17788 (I305282,I449905,I449887);
or I_17789 (I304784,I305031,I305282);
nor I_17790 (I304775,I305164,I305282);
or I_17791 (I304778,I304898,I305282);
DFFARX1 I_17792 (I305282,I2859,I304804,I304796,);
not I_17793 (I305382,I2866);
DFFARX1 I_17794 (I119853,I2859,I305382,I305408,);
not I_17795 (I305416,I305408);
nand I_17796 (I305433,I119856,I119832);
and I_17797 (I305450,I305433,I119829);
DFFARX1 I_17798 (I305450,I2859,I305382,I305476,);
not I_17799 (I305484,I119835);
DFFARX1 I_17800 (I119829,I2859,I305382,I305510,);
not I_17801 (I305518,I305510);
nor I_17802 (I305535,I305518,I305416);
and I_17803 (I305552,I305535,I119835);
nor I_17804 (I305569,I305518,I305484);
nor I_17805 (I305365,I305476,I305569);
DFFARX1 I_17806 (I119838,I2859,I305382,I305609,);
nor I_17807 (I305617,I305609,I305476);
not I_17808 (I305634,I305617);
not I_17809 (I305651,I305609);
nor I_17810 (I305668,I305651,I305552);
DFFARX1 I_17811 (I305668,I2859,I305382,I305368,);
nand I_17812 (I305699,I119841,I119850);
and I_17813 (I305716,I305699,I119847);
DFFARX1 I_17814 (I305716,I2859,I305382,I305742,);
nor I_17815 (I305750,I305742,I305609);
DFFARX1 I_17816 (I305750,I2859,I305382,I305350,);
nand I_17817 (I305781,I305742,I305651);
nand I_17818 (I305359,I305634,I305781);
not I_17819 (I305812,I305742);
nor I_17820 (I305829,I305812,I305552);
DFFARX1 I_17821 (I305829,I2859,I305382,I305371,);
nor I_17822 (I305860,I119844,I119850);
or I_17823 (I305362,I305609,I305860);
nor I_17824 (I305353,I305742,I305860);
or I_17825 (I305356,I305476,I305860);
DFFARX1 I_17826 (I305860,I2859,I305382,I305374,);
not I_17827 (I305960,I2866);
DFFARX1 I_17828 (I32197,I2859,I305960,I305986,);
not I_17829 (I305994,I305986);
nand I_17830 (I306011,I32206,I32215);
and I_17831 (I306028,I306011,I32194);
DFFARX1 I_17832 (I306028,I2859,I305960,I306054,);
not I_17833 (I306062,I32197);
DFFARX1 I_17834 (I32212,I2859,I305960,I306088,);
not I_17835 (I306096,I306088);
nor I_17836 (I306113,I306096,I305994);
and I_17837 (I306130,I306113,I32197);
nor I_17838 (I306147,I306096,I306062);
nor I_17839 (I305943,I306054,I306147);
DFFARX1 I_17840 (I32203,I2859,I305960,I306187,);
nor I_17841 (I306195,I306187,I306054);
not I_17842 (I306212,I306195);
not I_17843 (I306229,I306187);
nor I_17844 (I306246,I306229,I306130);
DFFARX1 I_17845 (I306246,I2859,I305960,I305946,);
nand I_17846 (I306277,I32218,I32194);
and I_17847 (I306294,I306277,I32200);
DFFARX1 I_17848 (I306294,I2859,I305960,I306320,);
nor I_17849 (I306328,I306320,I306187);
DFFARX1 I_17850 (I306328,I2859,I305960,I305928,);
nand I_17851 (I306359,I306320,I306229);
nand I_17852 (I305937,I306212,I306359);
not I_17853 (I306390,I306320);
nor I_17854 (I306407,I306390,I306130);
DFFARX1 I_17855 (I306407,I2859,I305960,I305949,);
nor I_17856 (I306438,I32209,I32194);
or I_17857 (I305940,I306187,I306438);
nor I_17858 (I305931,I306320,I306438);
or I_17859 (I305934,I306054,I306438);
DFFARX1 I_17860 (I306438,I2859,I305960,I305952,);
not I_17861 (I306538,I2866);
DFFARX1 I_17862 (I352336,I2859,I306538,I306564,);
not I_17863 (I306572,I306564);
nand I_17864 (I306589,I352324,I352342);
and I_17865 (I306606,I306589,I352339);
DFFARX1 I_17866 (I306606,I2859,I306538,I306632,);
not I_17867 (I306640,I352330);
DFFARX1 I_17868 (I352327,I2859,I306538,I306666,);
not I_17869 (I306674,I306666);
nor I_17870 (I306691,I306674,I306572);
and I_17871 (I306708,I306691,I352330);
nor I_17872 (I306725,I306674,I306640);
nor I_17873 (I306521,I306632,I306725);
DFFARX1 I_17874 (I352321,I2859,I306538,I306765,);
nor I_17875 (I306773,I306765,I306632);
not I_17876 (I306790,I306773);
not I_17877 (I306807,I306765);
nor I_17878 (I306824,I306807,I306708);
DFFARX1 I_17879 (I306824,I2859,I306538,I306524,);
nand I_17880 (I306855,I352321,I352324);
and I_17881 (I306872,I306855,I352327);
DFFARX1 I_17882 (I306872,I2859,I306538,I306898,);
nor I_17883 (I306906,I306898,I306765);
DFFARX1 I_17884 (I306906,I2859,I306538,I306506,);
nand I_17885 (I306937,I306898,I306807);
nand I_17886 (I306515,I306790,I306937);
not I_17887 (I306968,I306898);
nor I_17888 (I306985,I306968,I306708);
DFFARX1 I_17889 (I306985,I2859,I306538,I306527,);
nor I_17890 (I307016,I352333,I352324);
or I_17891 (I306518,I306765,I307016);
nor I_17892 (I306509,I306898,I307016);
or I_17893 (I306512,I306632,I307016);
DFFARX1 I_17894 (I307016,I2859,I306538,I306530,);
not I_17895 (I307116,I2866);
DFFARX1 I_17896 (I238302,I2859,I307116,I307142,);
not I_17897 (I307150,I307142);
nand I_17898 (I307167,I238311,I238320);
and I_17899 (I307184,I307167,I238326);
DFFARX1 I_17900 (I307184,I2859,I307116,I307210,);
not I_17901 (I307218,I238323);
DFFARX1 I_17902 (I238308,I2859,I307116,I307244,);
not I_17903 (I307252,I307244);
nor I_17904 (I307269,I307252,I307150);
and I_17905 (I307286,I307269,I238323);
nor I_17906 (I307303,I307252,I307218);
nor I_17907 (I307099,I307210,I307303);
DFFARX1 I_17908 (I238317,I2859,I307116,I307343,);
nor I_17909 (I307351,I307343,I307210);
not I_17910 (I307368,I307351);
not I_17911 (I307385,I307343);
nor I_17912 (I307402,I307385,I307286);
DFFARX1 I_17913 (I307402,I2859,I307116,I307102,);
nand I_17914 (I307433,I238314,I238305);
and I_17915 (I307450,I307433,I238302);
DFFARX1 I_17916 (I307450,I2859,I307116,I307476,);
nor I_17917 (I307484,I307476,I307343);
DFFARX1 I_17918 (I307484,I2859,I307116,I307084,);
nand I_17919 (I307515,I307476,I307385);
nand I_17920 (I307093,I307368,I307515);
not I_17921 (I307546,I307476);
nor I_17922 (I307563,I307546,I307286);
DFFARX1 I_17923 (I307563,I2859,I307116,I307105,);
nor I_17924 (I307594,I238305,I238305);
or I_17925 (I307096,I307343,I307594);
nor I_17926 (I307087,I307476,I307594);
or I_17927 (I307090,I307210,I307594);
DFFARX1 I_17928 (I307594,I2859,I307116,I307108,);
not I_17929 (I307694,I2866);
DFFARX1 I_17930 (I334418,I2859,I307694,I307720,);
not I_17931 (I307728,I307720);
nand I_17932 (I307745,I334406,I334424);
and I_17933 (I307762,I307745,I334421);
DFFARX1 I_17934 (I307762,I2859,I307694,I307788,);
not I_17935 (I307796,I334412);
DFFARX1 I_17936 (I334409,I2859,I307694,I307822,);
not I_17937 (I307830,I307822);
nor I_17938 (I307847,I307830,I307728);
and I_17939 (I307864,I307847,I334412);
nor I_17940 (I307881,I307830,I307796);
nor I_17941 (I307677,I307788,I307881);
DFFARX1 I_17942 (I334403,I2859,I307694,I307921,);
nor I_17943 (I307929,I307921,I307788);
not I_17944 (I307946,I307929);
not I_17945 (I307963,I307921);
nor I_17946 (I307980,I307963,I307864);
DFFARX1 I_17947 (I307980,I2859,I307694,I307680,);
nand I_17948 (I308011,I334403,I334406);
and I_17949 (I308028,I308011,I334409);
DFFARX1 I_17950 (I308028,I2859,I307694,I308054,);
nor I_17951 (I308062,I308054,I307921);
DFFARX1 I_17952 (I308062,I2859,I307694,I307662,);
nand I_17953 (I308093,I308054,I307963);
nand I_17954 (I307671,I307946,I308093);
not I_17955 (I308124,I308054);
nor I_17956 (I308141,I308124,I307864);
DFFARX1 I_17957 (I308141,I2859,I307694,I307683,);
nor I_17958 (I308172,I334415,I334406);
or I_17959 (I307674,I307921,I308172);
nor I_17960 (I307665,I308054,I308172);
or I_17961 (I307668,I307788,I308172);
DFFARX1 I_17962 (I308172,I2859,I307694,I307686,);
not I_17963 (I308272,I2866);
DFFARX1 I_17964 (I26927,I2859,I308272,I308298,);
not I_17965 (I308306,I308298);
nand I_17966 (I308323,I26936,I26945);
and I_17967 (I308340,I308323,I26924);
DFFARX1 I_17968 (I308340,I2859,I308272,I308366,);
not I_17969 (I308374,I26927);
DFFARX1 I_17970 (I26942,I2859,I308272,I308400,);
not I_17971 (I308408,I308400);
nor I_17972 (I308425,I308408,I308306);
and I_17973 (I308442,I308425,I26927);
nor I_17974 (I308459,I308408,I308374);
nor I_17975 (I308255,I308366,I308459);
DFFARX1 I_17976 (I26933,I2859,I308272,I308499,);
nor I_17977 (I308507,I308499,I308366);
not I_17978 (I308524,I308507);
not I_17979 (I308541,I308499);
nor I_17980 (I308558,I308541,I308442);
DFFARX1 I_17981 (I308558,I2859,I308272,I308258,);
nand I_17982 (I308589,I26948,I26924);
and I_17983 (I308606,I308589,I26930);
DFFARX1 I_17984 (I308606,I2859,I308272,I308632,);
nor I_17985 (I308640,I308632,I308499);
DFFARX1 I_17986 (I308640,I2859,I308272,I308240,);
nand I_17987 (I308671,I308632,I308541);
nand I_17988 (I308249,I308524,I308671);
not I_17989 (I308702,I308632);
nor I_17990 (I308719,I308702,I308442);
DFFARX1 I_17991 (I308719,I2859,I308272,I308261,);
nor I_17992 (I308750,I26939,I26924);
or I_17993 (I308252,I308499,I308750);
nor I_17994 (I308243,I308632,I308750);
or I_17995 (I308246,I308366,I308750);
DFFARX1 I_17996 (I308750,I2859,I308272,I308264,);
not I_17997 (I308850,I2866);
DFFARX1 I_17998 (I329675,I2859,I308850,I308876,);
not I_17999 (I308884,I308876);
nand I_18000 (I308901,I329663,I329681);
and I_18001 (I308918,I308901,I329678);
DFFARX1 I_18002 (I308918,I2859,I308850,I308944,);
not I_18003 (I308952,I329669);
DFFARX1 I_18004 (I329666,I2859,I308850,I308978,);
not I_18005 (I308986,I308978);
nor I_18006 (I309003,I308986,I308884);
and I_18007 (I309020,I309003,I329669);
nor I_18008 (I309037,I308986,I308952);
nor I_18009 (I308833,I308944,I309037);
DFFARX1 I_18010 (I329660,I2859,I308850,I309077,);
nor I_18011 (I309085,I309077,I308944);
not I_18012 (I309102,I309085);
not I_18013 (I309119,I309077);
nor I_18014 (I309136,I309119,I309020);
DFFARX1 I_18015 (I309136,I2859,I308850,I308836,);
nand I_18016 (I309167,I329660,I329663);
and I_18017 (I309184,I309167,I329666);
DFFARX1 I_18018 (I309184,I2859,I308850,I309210,);
nor I_18019 (I309218,I309210,I309077);
DFFARX1 I_18020 (I309218,I2859,I308850,I308818,);
nand I_18021 (I309249,I309210,I309119);
nand I_18022 (I308827,I309102,I309249);
not I_18023 (I309280,I309210);
nor I_18024 (I309297,I309280,I309020);
DFFARX1 I_18025 (I309297,I2859,I308850,I308839,);
nor I_18026 (I309328,I329672,I329663);
or I_18027 (I308830,I309077,I309328);
nor I_18028 (I308821,I309210,I309328);
or I_18029 (I308824,I308944,I309328);
DFFARX1 I_18030 (I309328,I2859,I308850,I308842,);
not I_18031 (I309428,I2866);
DFFARX1 I_18032 (I113529,I2859,I309428,I309454,);
not I_18033 (I309462,I309454);
nand I_18034 (I309479,I113532,I113508);
and I_18035 (I309496,I309479,I113505);
DFFARX1 I_18036 (I309496,I2859,I309428,I309522,);
not I_18037 (I309530,I113511);
DFFARX1 I_18038 (I113505,I2859,I309428,I309556,);
not I_18039 (I309564,I309556);
nor I_18040 (I309581,I309564,I309462);
and I_18041 (I309598,I309581,I113511);
nor I_18042 (I309615,I309564,I309530);
nor I_18043 (I309411,I309522,I309615);
DFFARX1 I_18044 (I113514,I2859,I309428,I309655,);
nor I_18045 (I309663,I309655,I309522);
not I_18046 (I309680,I309663);
not I_18047 (I309697,I309655);
nor I_18048 (I309714,I309697,I309598);
DFFARX1 I_18049 (I309714,I2859,I309428,I309414,);
nand I_18050 (I309745,I113517,I113526);
and I_18051 (I309762,I309745,I113523);
DFFARX1 I_18052 (I309762,I2859,I309428,I309788,);
nor I_18053 (I309796,I309788,I309655);
DFFARX1 I_18054 (I309796,I2859,I309428,I309396,);
nand I_18055 (I309827,I309788,I309697);
nand I_18056 (I309405,I309680,I309827);
not I_18057 (I309858,I309788);
nor I_18058 (I309875,I309858,I309598);
DFFARX1 I_18059 (I309875,I2859,I309428,I309417,);
nor I_18060 (I309906,I113520,I113526);
or I_18061 (I309408,I309655,I309906);
nor I_18062 (I309399,I309788,I309906);
or I_18063 (I309402,I309522,I309906);
DFFARX1 I_18064 (I309906,I2859,I309428,I309420,);
not I_18065 (I310006,I2866);
DFFARX1 I_18066 (I417590,I2859,I310006,I310032,);
not I_18067 (I310040,I310032);
nand I_18068 (I310057,I417587,I417605);
and I_18069 (I310074,I310057,I417602);
DFFARX1 I_18070 (I310074,I2859,I310006,I310100,);
not I_18071 (I310108,I417584);
DFFARX1 I_18072 (I417587,I2859,I310006,I310134,);
not I_18073 (I310142,I310134);
nor I_18074 (I310159,I310142,I310040);
and I_18075 (I310176,I310159,I417584);
nor I_18076 (I310193,I310142,I310108);
nor I_18077 (I309989,I310100,I310193);
DFFARX1 I_18078 (I417596,I2859,I310006,I310233,);
nor I_18079 (I310241,I310233,I310100);
not I_18080 (I310258,I310241);
not I_18081 (I310275,I310233);
nor I_18082 (I310292,I310275,I310176);
DFFARX1 I_18083 (I310292,I2859,I310006,I309992,);
nand I_18084 (I310323,I417599,I417584);
and I_18085 (I310340,I310323,I417590);
DFFARX1 I_18086 (I310340,I2859,I310006,I310366,);
nor I_18087 (I310374,I310366,I310233);
DFFARX1 I_18088 (I310374,I2859,I310006,I309974,);
nand I_18089 (I310405,I310366,I310275);
nand I_18090 (I309983,I310258,I310405);
not I_18091 (I310436,I310366);
nor I_18092 (I310453,I310436,I310176);
DFFARX1 I_18093 (I310453,I2859,I310006,I309995,);
nor I_18094 (I310484,I417593,I417584);
or I_18095 (I309986,I310233,I310484);
nor I_18096 (I309977,I310366,I310484);
or I_18097 (I309980,I310100,I310484);
DFFARX1 I_18098 (I310484,I2859,I310006,I309998,);
not I_18099 (I310584,I2866);
DFFARX1 I_18100 (I561227,I2859,I310584,I310610,);
not I_18101 (I310618,I310610);
nand I_18102 (I310635,I561212,I561200);
and I_18103 (I310652,I310635,I561215);
DFFARX1 I_18104 (I310652,I2859,I310584,I310678,);
not I_18105 (I310686,I561200);
DFFARX1 I_18106 (I561218,I2859,I310584,I310712,);
not I_18107 (I310720,I310712);
nor I_18108 (I310737,I310720,I310618);
and I_18109 (I310754,I310737,I561200);
nor I_18110 (I310771,I310720,I310686);
nor I_18111 (I310567,I310678,I310771);
DFFARX1 I_18112 (I561206,I2859,I310584,I310811,);
nor I_18113 (I310819,I310811,I310678);
not I_18114 (I310836,I310819);
not I_18115 (I310853,I310811);
nor I_18116 (I310870,I310853,I310754);
DFFARX1 I_18117 (I310870,I2859,I310584,I310570,);
nand I_18118 (I310901,I561203,I561209);
and I_18119 (I310918,I310901,I561224);
DFFARX1 I_18120 (I310918,I2859,I310584,I310944,);
nor I_18121 (I310952,I310944,I310811);
DFFARX1 I_18122 (I310952,I2859,I310584,I310552,);
nand I_18123 (I310983,I310944,I310853);
nand I_18124 (I310561,I310836,I310983);
not I_18125 (I311014,I310944);
nor I_18126 (I311031,I311014,I310754);
DFFARX1 I_18127 (I311031,I2859,I310584,I310573,);
nor I_18128 (I311062,I561221,I561209);
or I_18129 (I310564,I310811,I311062);
nor I_18130 (I310555,I310944,I311062);
or I_18131 (I310558,I310678,I311062);
DFFARX1 I_18132 (I311062,I2859,I310584,I310576,);
not I_18133 (I311162,I2866);
DFFARX1 I_18134 (I185441,I2859,I311162,I311188,);
not I_18135 (I311196,I311188);
nand I_18136 (I311213,I185432,I185450);
and I_18137 (I311230,I311213,I185453);
DFFARX1 I_18138 (I311230,I2859,I311162,I311256,);
not I_18139 (I311264,I185447);
DFFARX1 I_18140 (I185435,I2859,I311162,I311290,);
not I_18141 (I311298,I311290);
nor I_18142 (I311315,I311298,I311196);
and I_18143 (I311332,I311315,I185447);
nor I_18144 (I311349,I311298,I311264);
nor I_18145 (I311145,I311256,I311349);
DFFARX1 I_18146 (I185444,I2859,I311162,I311389,);
nor I_18147 (I311397,I311389,I311256);
not I_18148 (I311414,I311397);
not I_18149 (I311431,I311389);
nor I_18150 (I311448,I311431,I311332);
DFFARX1 I_18151 (I311448,I2859,I311162,I311148,);
nand I_18152 (I311479,I185459,I185456);
and I_18153 (I311496,I311479,I185438);
DFFARX1 I_18154 (I311496,I2859,I311162,I311522,);
nor I_18155 (I311530,I311522,I311389);
DFFARX1 I_18156 (I311530,I2859,I311162,I311130,);
nand I_18157 (I311561,I311522,I311431);
nand I_18158 (I311139,I311414,I311561);
not I_18159 (I311592,I311522);
nor I_18160 (I311609,I311592,I311332);
DFFARX1 I_18161 (I311609,I2859,I311162,I311151,);
nor I_18162 (I311640,I185432,I185456);
or I_18163 (I311142,I311389,I311640);
nor I_18164 (I311133,I311522,I311640);
or I_18165 (I311136,I311256,I311640);
DFFARX1 I_18166 (I311640,I2859,I311162,I311154,);
not I_18167 (I311740,I2866);
DFFARX1 I_18168 (I87002,I2859,I311740,I311766,);
not I_18169 (I311774,I311766);
nand I_18170 (I311791,I87005,I87026);
and I_18171 (I311808,I311791,I87014);
DFFARX1 I_18172 (I311808,I2859,I311740,I311834,);
not I_18173 (I311842,I87011);
DFFARX1 I_18174 (I87002,I2859,I311740,I311868,);
not I_18175 (I311876,I311868);
nor I_18176 (I311893,I311876,I311774);
and I_18177 (I311910,I311893,I87011);
nor I_18178 (I311927,I311876,I311842);
nor I_18179 (I311723,I311834,I311927);
DFFARX1 I_18180 (I87020,I2859,I311740,I311967,);
nor I_18181 (I311975,I311967,I311834);
not I_18182 (I311992,I311975);
not I_18183 (I312009,I311967);
nor I_18184 (I312026,I312009,I311910);
DFFARX1 I_18185 (I312026,I2859,I311740,I311726,);
nand I_18186 (I312057,I87005,I87008);
and I_18187 (I312074,I312057,I87017);
DFFARX1 I_18188 (I312074,I2859,I311740,I312100,);
nor I_18189 (I312108,I312100,I311967);
DFFARX1 I_18190 (I312108,I2859,I311740,I311708,);
nand I_18191 (I312139,I312100,I312009);
nand I_18192 (I311717,I311992,I312139);
not I_18193 (I312170,I312100);
nor I_18194 (I312187,I312170,I311910);
DFFARX1 I_18195 (I312187,I2859,I311740,I311729,);
nor I_18196 (I312218,I87023,I87008);
or I_18197 (I311720,I311967,I312218);
nor I_18198 (I311711,I312100,I312218);
or I_18199 (I311714,I311834,I312218);
DFFARX1 I_18200 (I312218,I2859,I311740,I311732,);
not I_18201 (I312318,I2866);
DFFARX1 I_18202 (I80457,I2859,I312318,I312344,);
not I_18203 (I312352,I312344);
nand I_18204 (I312369,I80460,I80481);
and I_18205 (I312386,I312369,I80469);
DFFARX1 I_18206 (I312386,I2859,I312318,I312412,);
not I_18207 (I312420,I80466);
DFFARX1 I_18208 (I80457,I2859,I312318,I312446,);
not I_18209 (I312454,I312446);
nor I_18210 (I312471,I312454,I312352);
and I_18211 (I312488,I312471,I80466);
nor I_18212 (I312505,I312454,I312420);
nor I_18213 (I312301,I312412,I312505);
DFFARX1 I_18214 (I80475,I2859,I312318,I312545,);
nor I_18215 (I312553,I312545,I312412);
not I_18216 (I312570,I312553);
not I_18217 (I312587,I312545);
nor I_18218 (I312604,I312587,I312488);
DFFARX1 I_18219 (I312604,I2859,I312318,I312304,);
nand I_18220 (I312635,I80460,I80463);
and I_18221 (I312652,I312635,I80472);
DFFARX1 I_18222 (I312652,I2859,I312318,I312678,);
nor I_18223 (I312686,I312678,I312545);
DFFARX1 I_18224 (I312686,I2859,I312318,I312286,);
nand I_18225 (I312717,I312678,I312587);
nand I_18226 (I312295,I312570,I312717);
not I_18227 (I312748,I312678);
nor I_18228 (I312765,I312748,I312488);
DFFARX1 I_18229 (I312765,I2859,I312318,I312307,);
nor I_18230 (I312796,I80478,I80463);
or I_18231 (I312298,I312545,I312796);
nor I_18232 (I312289,I312678,I312796);
or I_18233 (I312292,I312412,I312796);
DFFARX1 I_18234 (I312796,I2859,I312318,I312310,);
not I_18235 (I312896,I2866);
DFFARX1 I_18236 (I39048,I2859,I312896,I312922,);
not I_18237 (I312930,I312922);
nand I_18238 (I312947,I39057,I39066);
and I_18239 (I312964,I312947,I39045);
DFFARX1 I_18240 (I312964,I2859,I312896,I312990,);
not I_18241 (I312998,I39048);
DFFARX1 I_18242 (I39063,I2859,I312896,I313024,);
not I_18243 (I313032,I313024);
nor I_18244 (I313049,I313032,I312930);
and I_18245 (I313066,I313049,I39048);
nor I_18246 (I313083,I313032,I312998);
nor I_18247 (I312879,I312990,I313083);
DFFARX1 I_18248 (I39054,I2859,I312896,I313123,);
nor I_18249 (I313131,I313123,I312990);
not I_18250 (I313148,I313131);
not I_18251 (I313165,I313123);
nor I_18252 (I313182,I313165,I313066);
DFFARX1 I_18253 (I313182,I2859,I312896,I312882,);
nand I_18254 (I313213,I39069,I39045);
and I_18255 (I313230,I313213,I39051);
DFFARX1 I_18256 (I313230,I2859,I312896,I313256,);
nor I_18257 (I313264,I313256,I313123);
DFFARX1 I_18258 (I313264,I2859,I312896,I312864,);
nand I_18259 (I313295,I313256,I313165);
nand I_18260 (I312873,I313148,I313295);
not I_18261 (I313326,I313256);
nor I_18262 (I313343,I313326,I313066);
DFFARX1 I_18263 (I313343,I2859,I312896,I312885,);
nor I_18264 (I313374,I39060,I39045);
or I_18265 (I312876,I313123,I313374);
nor I_18266 (I312867,I313256,I313374);
or I_18267 (I312870,I312990,I313374);
DFFARX1 I_18268 (I313374,I2859,I312896,I312888,);
not I_18269 (I313474,I2866);
DFFARX1 I_18270 (I506834,I2859,I313474,I313500,);
not I_18271 (I313508,I313500);
nand I_18272 (I313525,I506837,I506846);
and I_18273 (I313542,I313525,I506849);
DFFARX1 I_18274 (I313542,I2859,I313474,I313568,);
not I_18275 (I313576,I506858);
DFFARX1 I_18276 (I506840,I2859,I313474,I313602,);
not I_18277 (I313610,I313602);
nor I_18278 (I313627,I313610,I313508);
and I_18279 (I313644,I313627,I506858);
nor I_18280 (I313661,I313610,I313576);
nor I_18281 (I313457,I313568,I313661);
DFFARX1 I_18282 (I506837,I2859,I313474,I313701,);
nor I_18283 (I313709,I313701,I313568);
not I_18284 (I313726,I313709);
not I_18285 (I313743,I313701);
nor I_18286 (I313760,I313743,I313644);
DFFARX1 I_18287 (I313760,I2859,I313474,I313460,);
nand I_18288 (I313791,I506855,I506834);
and I_18289 (I313808,I313791,I506852);
DFFARX1 I_18290 (I313808,I2859,I313474,I313834,);
nor I_18291 (I313842,I313834,I313701);
DFFARX1 I_18292 (I313842,I2859,I313474,I313442,);
nand I_18293 (I313873,I313834,I313743);
nand I_18294 (I313451,I313726,I313873);
not I_18295 (I313904,I313834);
nor I_18296 (I313921,I313904,I313644);
DFFARX1 I_18297 (I313921,I2859,I313474,I313463,);
nor I_18298 (I313952,I506843,I506834);
or I_18299 (I313454,I313701,I313952);
nor I_18300 (I313445,I313834,I313952);
or I_18301 (I313448,I313568,I313952);
DFFARX1 I_18302 (I313952,I2859,I313474,I313466,);
not I_18303 (I314052,I2866);
DFFARX1 I_18304 (I361831,I2859,I314052,I314078,);
not I_18305 (I314086,I314078);
nand I_18306 (I314103,I361807,I361822);
and I_18307 (I314120,I314103,I361834);
DFFARX1 I_18308 (I314120,I2859,I314052,I314146,);
not I_18309 (I314154,I361819);
DFFARX1 I_18310 (I361810,I2859,I314052,I314180,);
not I_18311 (I314188,I314180);
nor I_18312 (I314205,I314188,I314086);
and I_18313 (I314222,I314205,I361819);
nor I_18314 (I314239,I314188,I314154);
nor I_18315 (I314035,I314146,I314239);
DFFARX1 I_18316 (I361807,I2859,I314052,I314279,);
nor I_18317 (I314287,I314279,I314146);
not I_18318 (I314304,I314287);
not I_18319 (I314321,I314279);
nor I_18320 (I314338,I314321,I314222);
DFFARX1 I_18321 (I314338,I2859,I314052,I314038,);
nand I_18322 (I314369,I361825,I361816);
and I_18323 (I314386,I314369,I361828);
DFFARX1 I_18324 (I314386,I2859,I314052,I314412,);
nor I_18325 (I314420,I314412,I314279);
DFFARX1 I_18326 (I314420,I2859,I314052,I314020,);
nand I_18327 (I314451,I314412,I314321);
nand I_18328 (I314029,I314304,I314451);
not I_18329 (I314482,I314412);
nor I_18330 (I314499,I314482,I314222);
DFFARX1 I_18331 (I314499,I2859,I314052,I314041,);
nor I_18332 (I314530,I361813,I361816);
or I_18333 (I314032,I314279,I314530);
nor I_18334 (I314023,I314412,I314530);
or I_18335 (I314026,I314146,I314530);
DFFARX1 I_18336 (I314530,I2859,I314052,I314044,);
not I_18337 (I314630,I2866);
DFFARX1 I_18338 (I178369,I2859,I314630,I314656,);
not I_18339 (I314664,I314656);
nand I_18340 (I314681,I178360,I178378);
and I_18341 (I314698,I314681,I178381);
DFFARX1 I_18342 (I314698,I2859,I314630,I314724,);
not I_18343 (I314732,I178375);
DFFARX1 I_18344 (I178363,I2859,I314630,I314758,);
not I_18345 (I314766,I314758);
nor I_18346 (I314783,I314766,I314664);
and I_18347 (I314800,I314783,I178375);
nor I_18348 (I314817,I314766,I314732);
nor I_18349 (I314613,I314724,I314817);
DFFARX1 I_18350 (I178372,I2859,I314630,I314857,);
nor I_18351 (I314865,I314857,I314724);
not I_18352 (I314882,I314865);
not I_18353 (I314899,I314857);
nor I_18354 (I314916,I314899,I314800);
DFFARX1 I_18355 (I314916,I2859,I314630,I314616,);
nand I_18356 (I314947,I178387,I178384);
and I_18357 (I314964,I314947,I178366);
DFFARX1 I_18358 (I314964,I2859,I314630,I314990,);
nor I_18359 (I314998,I314990,I314857);
DFFARX1 I_18360 (I314998,I2859,I314630,I314598,);
nand I_18361 (I315029,I314990,I314899);
nand I_18362 (I314607,I314882,I315029);
not I_18363 (I315060,I314990);
nor I_18364 (I315077,I315060,I314800);
DFFARX1 I_18365 (I315077,I2859,I314630,I314619,);
nor I_18366 (I315108,I178360,I178384);
or I_18367 (I314610,I314857,I315108);
nor I_18368 (I314601,I314990,I315108);
or I_18369 (I314604,I314724,I315108);
DFFARX1 I_18370 (I315108,I2859,I314630,I314622,);
not I_18371 (I315208,I2866);
DFFARX1 I_18372 (I401883,I2859,I315208,I315234,);
not I_18373 (I315242,I315234);
nand I_18374 (I315259,I401859,I401874);
and I_18375 (I315276,I315259,I401886);
DFFARX1 I_18376 (I315276,I2859,I315208,I315302,);
not I_18377 (I315310,I401871);
DFFARX1 I_18378 (I401862,I2859,I315208,I315336,);
not I_18379 (I315344,I315336);
nor I_18380 (I315361,I315344,I315242);
and I_18381 (I315378,I315361,I401871);
nor I_18382 (I315395,I315344,I315310);
nor I_18383 (I315191,I315302,I315395);
DFFARX1 I_18384 (I401859,I2859,I315208,I315435,);
nor I_18385 (I315443,I315435,I315302);
not I_18386 (I315460,I315443);
not I_18387 (I315477,I315435);
nor I_18388 (I315494,I315477,I315378);
DFFARX1 I_18389 (I315494,I2859,I315208,I315194,);
nand I_18390 (I315525,I401877,I401868);
and I_18391 (I315542,I315525,I401880);
DFFARX1 I_18392 (I315542,I2859,I315208,I315568,);
nor I_18393 (I315576,I315568,I315435);
DFFARX1 I_18394 (I315576,I2859,I315208,I315176,);
nand I_18395 (I315607,I315568,I315477);
nand I_18396 (I315185,I315460,I315607);
not I_18397 (I315638,I315568);
nor I_18398 (I315655,I315638,I315378);
DFFARX1 I_18399 (I315655,I2859,I315208,I315197,);
nor I_18400 (I315686,I401865,I401868);
or I_18401 (I315188,I315435,I315686);
nor I_18402 (I315179,I315568,I315686);
or I_18403 (I315182,I315302,I315686);
DFFARX1 I_18404 (I315686,I2859,I315208,I315200,);
not I_18405 (I315786,I2866);
DFFARX1 I_18406 (I430493,I2859,I315786,I315812,);
not I_18407 (I315820,I315812);
nand I_18408 (I315837,I430490,I430508);
and I_18409 (I315854,I315837,I430505);
DFFARX1 I_18410 (I315854,I2859,I315786,I315880,);
not I_18411 (I315888,I430487);
DFFARX1 I_18412 (I430490,I2859,I315786,I315914,);
not I_18413 (I315922,I315914);
nor I_18414 (I315939,I315922,I315820);
and I_18415 (I315956,I315939,I430487);
nor I_18416 (I315973,I315922,I315888);
nor I_18417 (I315769,I315880,I315973);
DFFARX1 I_18418 (I430499,I2859,I315786,I316013,);
nor I_18419 (I316021,I316013,I315880);
not I_18420 (I316038,I316021);
not I_18421 (I316055,I316013);
nor I_18422 (I316072,I316055,I315956);
DFFARX1 I_18423 (I316072,I2859,I315786,I315772,);
nand I_18424 (I316103,I430502,I430487);
and I_18425 (I316120,I316103,I430493);
DFFARX1 I_18426 (I316120,I2859,I315786,I316146,);
nor I_18427 (I316154,I316146,I316013);
DFFARX1 I_18428 (I316154,I2859,I315786,I315754,);
nand I_18429 (I316185,I316146,I316055);
nand I_18430 (I315763,I316038,I316185);
not I_18431 (I316216,I316146);
nor I_18432 (I316233,I316216,I315956);
DFFARX1 I_18433 (I316233,I2859,I315786,I315775,);
nor I_18434 (I316264,I430496,I430487);
or I_18435 (I315766,I316013,I316264);
nor I_18436 (I315757,I316146,I316264);
or I_18437 (I315760,I315880,I316264);
DFFARX1 I_18438 (I316264,I2859,I315786,I315778,);
not I_18439 (I316364,I2866);
DFFARX1 I_18440 (I75102,I2859,I316364,I316390,);
not I_18441 (I316398,I316390);
nand I_18442 (I316415,I75105,I75126);
and I_18443 (I316432,I316415,I75114);
DFFARX1 I_18444 (I316432,I2859,I316364,I316458,);
not I_18445 (I316466,I75111);
DFFARX1 I_18446 (I75102,I2859,I316364,I316492,);
not I_18447 (I316500,I316492);
nor I_18448 (I316517,I316500,I316398);
and I_18449 (I316534,I316517,I75111);
nor I_18450 (I316551,I316500,I316466);
nor I_18451 (I316347,I316458,I316551);
DFFARX1 I_18452 (I75120,I2859,I316364,I316591,);
nor I_18453 (I316599,I316591,I316458);
not I_18454 (I316616,I316599);
not I_18455 (I316633,I316591);
nor I_18456 (I316650,I316633,I316534);
DFFARX1 I_18457 (I316650,I2859,I316364,I316350,);
nand I_18458 (I316681,I75105,I75108);
and I_18459 (I316698,I316681,I75117);
DFFARX1 I_18460 (I316698,I2859,I316364,I316724,);
nor I_18461 (I316732,I316724,I316591);
DFFARX1 I_18462 (I316732,I2859,I316364,I316332,);
nand I_18463 (I316763,I316724,I316633);
nand I_18464 (I316341,I316616,I316763);
not I_18465 (I316794,I316724);
nor I_18466 (I316811,I316794,I316534);
DFFARX1 I_18467 (I316811,I2859,I316364,I316353,);
nor I_18468 (I316842,I75123,I75108);
or I_18469 (I316344,I316591,I316842);
nor I_18470 (I316335,I316724,I316842);
or I_18471 (I316338,I316458,I316842);
DFFARX1 I_18472 (I316842,I2859,I316364,I316356,);
not I_18473 (I316942,I2866);
DFFARX1 I_18474 (I36413,I2859,I316942,I316968,);
not I_18475 (I316976,I316968);
nand I_18476 (I316993,I36422,I36431);
and I_18477 (I317010,I316993,I36410);
DFFARX1 I_18478 (I317010,I2859,I316942,I317036,);
not I_18479 (I317044,I36413);
DFFARX1 I_18480 (I36428,I2859,I316942,I317070,);
not I_18481 (I317078,I317070);
nor I_18482 (I317095,I317078,I316976);
and I_18483 (I317112,I317095,I36413);
nor I_18484 (I317129,I317078,I317044);
nor I_18485 (I316925,I317036,I317129);
DFFARX1 I_18486 (I36419,I2859,I316942,I317169,);
nor I_18487 (I317177,I317169,I317036);
not I_18488 (I317194,I317177);
not I_18489 (I317211,I317169);
nor I_18490 (I317228,I317211,I317112);
DFFARX1 I_18491 (I317228,I2859,I316942,I316928,);
nand I_18492 (I317259,I36434,I36410);
and I_18493 (I317276,I317259,I36416);
DFFARX1 I_18494 (I317276,I2859,I316942,I317302,);
nor I_18495 (I317310,I317302,I317169);
DFFARX1 I_18496 (I317310,I2859,I316942,I316910,);
nand I_18497 (I317341,I317302,I317211);
nand I_18498 (I316919,I317194,I317341);
not I_18499 (I317372,I317302);
nor I_18500 (I317389,I317372,I317112);
DFFARX1 I_18501 (I317389,I2859,I316942,I316931,);
nor I_18502 (I317420,I36425,I36410);
or I_18503 (I316922,I317169,I317420);
nor I_18504 (I316913,I317302,I317420);
or I_18505 (I316916,I317036,I317420);
DFFARX1 I_18506 (I317420,I2859,I316942,I316934,);
not I_18507 (I317520,I2866);
DFFARX1 I_18508 (I322297,I2859,I317520,I317546,);
not I_18509 (I317554,I317546);
nand I_18510 (I317571,I322285,I322303);
and I_18511 (I317588,I317571,I322300);
DFFARX1 I_18512 (I317588,I2859,I317520,I317614,);
not I_18513 (I317622,I322291);
DFFARX1 I_18514 (I322288,I2859,I317520,I317648,);
not I_18515 (I317656,I317648);
nor I_18516 (I317673,I317656,I317554);
and I_18517 (I317690,I317673,I322291);
nor I_18518 (I317707,I317656,I317622);
nor I_18519 (I317503,I317614,I317707);
DFFARX1 I_18520 (I322282,I2859,I317520,I317747,);
nor I_18521 (I317755,I317747,I317614);
not I_18522 (I317772,I317755);
not I_18523 (I317789,I317747);
nor I_18524 (I317806,I317789,I317690);
DFFARX1 I_18525 (I317806,I2859,I317520,I317506,);
nand I_18526 (I317837,I322282,I322285);
and I_18527 (I317854,I317837,I322288);
DFFARX1 I_18528 (I317854,I2859,I317520,I317880,);
nor I_18529 (I317888,I317880,I317747);
DFFARX1 I_18530 (I317888,I2859,I317520,I317488,);
nand I_18531 (I317919,I317880,I317789);
nand I_18532 (I317497,I317772,I317919);
not I_18533 (I317950,I317880);
nor I_18534 (I317967,I317950,I317690);
DFFARX1 I_18535 (I317967,I2859,I317520,I317509,);
nor I_18536 (I317998,I322294,I322285);
or I_18537 (I317500,I317747,I317998);
nor I_18538 (I317491,I317880,I317998);
or I_18539 (I317494,I317614,I317998);
DFFARX1 I_18540 (I317998,I2859,I317520,I317512,);
not I_18541 (I318095,I2866);
DFFARX1 I_18542 (I497298,I2859,I318095,I318121,);
not I_18543 (I318129,I318121);
nand I_18544 (I318146,I497280,I497280);
and I_18545 (I318163,I318146,I497286);
DFFARX1 I_18546 (I318163,I2859,I318095,I318189,);
DFFARX1 I_18547 (I318189,I2859,I318095,I318084,);
DFFARX1 I_18548 (I497283,I2859,I318095,I318220,);
nand I_18549 (I318228,I318220,I497292);
not I_18550 (I318245,I318228);
DFFARX1 I_18551 (I318245,I2859,I318095,I318271,);
not I_18552 (I318279,I318271);
nor I_18553 (I318087,I318129,I318279);
DFFARX1 I_18554 (I497304,I2859,I318095,I318319,);
nor I_18555 (I318078,I318319,I318189);
nor I_18556 (I318069,I318319,I318245);
nand I_18557 (I318355,I497295,I497289);
and I_18558 (I318372,I318355,I497283);
DFFARX1 I_18559 (I318372,I2859,I318095,I318398,);
not I_18560 (I318406,I318398);
nand I_18561 (I318423,I318406,I318319);
nand I_18562 (I318072,I318406,I318228);
nor I_18563 (I318454,I497301,I497289);
and I_18564 (I318471,I318319,I318454);
nor I_18565 (I318488,I318406,I318471);
DFFARX1 I_18566 (I318488,I2859,I318095,I318081,);
nor I_18567 (I318519,I318121,I318454);
DFFARX1 I_18568 (I318519,I2859,I318095,I318066,);
nor I_18569 (I318550,I318398,I318454);
not I_18570 (I318567,I318550);
nand I_18571 (I318075,I318567,I318423);
not I_18572 (I318622,I2866);
DFFARX1 I_18573 (I396048,I2859,I318622,I318648,);
not I_18574 (I318656,I318648);
nand I_18575 (I318673,I396063,I396045);
and I_18576 (I318690,I318673,I396045);
DFFARX1 I_18577 (I318690,I2859,I318622,I318716,);
DFFARX1 I_18578 (I318716,I2859,I318622,I318611,);
DFFARX1 I_18579 (I396054,I2859,I318622,I318747,);
nand I_18580 (I318755,I318747,I396072);
not I_18581 (I318772,I318755);
DFFARX1 I_18582 (I318772,I2859,I318622,I318798,);
not I_18583 (I318806,I318798);
nor I_18584 (I318614,I318656,I318806);
DFFARX1 I_18585 (I396069,I2859,I318622,I318846,);
nor I_18586 (I318605,I318846,I318716);
nor I_18587 (I318596,I318846,I318772);
nand I_18588 (I318882,I396066,I396057);
and I_18589 (I318899,I318882,I396051);
DFFARX1 I_18590 (I318899,I2859,I318622,I318925,);
not I_18591 (I318933,I318925);
nand I_18592 (I318950,I318933,I318846);
nand I_18593 (I318599,I318933,I318755);
nor I_18594 (I318981,I396060,I396057);
and I_18595 (I318998,I318846,I318981);
nor I_18596 (I319015,I318933,I318998);
DFFARX1 I_18597 (I319015,I2859,I318622,I318608,);
nor I_18598 (I319046,I318648,I318981);
DFFARX1 I_18599 (I319046,I2859,I318622,I318593,);
nor I_18600 (I319077,I318925,I318981);
not I_18601 (I319094,I319077);
nand I_18602 (I318602,I319094,I318950);
not I_18603 (I319149,I2866);
DFFARX1 I_18604 (I184350,I2859,I319149,I319175,);
not I_18605 (I319183,I319175);
nand I_18606 (I319200,I184347,I184356);
and I_18607 (I319217,I319200,I184365);
DFFARX1 I_18608 (I319217,I2859,I319149,I319243,);
DFFARX1 I_18609 (I319243,I2859,I319149,I319138,);
DFFARX1 I_18610 (I184368,I2859,I319149,I319274,);
nand I_18611 (I319282,I319274,I184371);
not I_18612 (I319299,I319282);
DFFARX1 I_18613 (I319299,I2859,I319149,I319325,);
not I_18614 (I319333,I319325);
nor I_18615 (I319141,I319183,I319333);
DFFARX1 I_18616 (I184344,I2859,I319149,I319373,);
nor I_18617 (I319132,I319373,I319243);
nor I_18618 (I319123,I319373,I319299);
nand I_18619 (I319409,I184359,I184362);
and I_18620 (I319426,I319409,I184353);
DFFARX1 I_18621 (I319426,I2859,I319149,I319452,);
not I_18622 (I319460,I319452);
nand I_18623 (I319477,I319460,I319373);
nand I_18624 (I319126,I319460,I319282);
nor I_18625 (I319508,I184344,I184362);
and I_18626 (I319525,I319373,I319508);
nor I_18627 (I319542,I319460,I319525);
DFFARX1 I_18628 (I319542,I2859,I319149,I319135,);
nor I_18629 (I319573,I319175,I319508);
DFFARX1 I_18630 (I319573,I2859,I319149,I319120,);
nor I_18631 (I319604,I319452,I319508);
not I_18632 (I319621,I319604);
nand I_18633 (I319129,I319621,I319477);
not I_18634 (I319676,I2866);
DFFARX1 I_18635 (I257954,I2859,I319676,I319702,);
not I_18636 (I319710,I319702);
nand I_18637 (I319727,I257957,I257954);
and I_18638 (I319744,I319727,I257966);
DFFARX1 I_18639 (I319744,I2859,I319676,I319770,);
DFFARX1 I_18640 (I319770,I2859,I319676,I319665,);
DFFARX1 I_18641 (I257963,I2859,I319676,I319801,);
nand I_18642 (I319809,I319801,I257969);
not I_18643 (I319826,I319809);
DFFARX1 I_18644 (I319826,I2859,I319676,I319852,);
not I_18645 (I319860,I319852);
nor I_18646 (I319668,I319710,I319860);
DFFARX1 I_18647 (I257978,I2859,I319676,I319900,);
nor I_18648 (I319659,I319900,I319770);
nor I_18649 (I319650,I319900,I319826);
nand I_18650 (I319936,I257972,I257960);
and I_18651 (I319953,I319936,I257957);
DFFARX1 I_18652 (I319953,I2859,I319676,I319979,);
not I_18653 (I319987,I319979);
nand I_18654 (I320004,I319987,I319900);
nand I_18655 (I319653,I319987,I319809);
nor I_18656 (I320035,I257975,I257960);
and I_18657 (I320052,I319900,I320035);
nor I_18658 (I320069,I319987,I320052);
DFFARX1 I_18659 (I320069,I2859,I319676,I319662,);
nor I_18660 (I320100,I319702,I320035);
DFFARX1 I_18661 (I320100,I2859,I319676,I319647,);
nor I_18662 (I320131,I319979,I320035);
not I_18663 (I320148,I320131);
nand I_18664 (I319656,I320148,I320004);
not I_18665 (I320203,I2866);
DFFARX1 I_18666 (I259110,I2859,I320203,I320229,);
not I_18667 (I320237,I320229);
nand I_18668 (I320254,I259113,I259110);
and I_18669 (I320271,I320254,I259122);
DFFARX1 I_18670 (I320271,I2859,I320203,I320297,);
DFFARX1 I_18671 (I320297,I2859,I320203,I320192,);
DFFARX1 I_18672 (I259119,I2859,I320203,I320328,);
nand I_18673 (I320336,I320328,I259125);
not I_18674 (I320353,I320336);
DFFARX1 I_18675 (I320353,I2859,I320203,I320379,);
not I_18676 (I320387,I320379);
nor I_18677 (I320195,I320237,I320387);
DFFARX1 I_18678 (I259134,I2859,I320203,I320427,);
nor I_18679 (I320186,I320427,I320297);
nor I_18680 (I320177,I320427,I320353);
nand I_18681 (I320463,I259128,I259116);
and I_18682 (I320480,I320463,I259113);
DFFARX1 I_18683 (I320480,I2859,I320203,I320506,);
not I_18684 (I320514,I320506);
nand I_18685 (I320531,I320514,I320427);
nand I_18686 (I320180,I320514,I320336);
nor I_18687 (I320562,I259131,I259116);
and I_18688 (I320579,I320427,I320562);
nor I_18689 (I320596,I320514,I320579);
DFFARX1 I_18690 (I320596,I2859,I320203,I320189,);
nor I_18691 (I320627,I320229,I320562);
DFFARX1 I_18692 (I320627,I2859,I320203,I320174,);
nor I_18693 (I320658,I320506,I320562);
not I_18694 (I320675,I320658);
nand I_18695 (I320183,I320675,I320531);
not I_18696 (I320730,I2866);
DFFARX1 I_18697 (I419837,I2859,I320730,I320756,);
not I_18698 (I320764,I320756);
nand I_18699 (I320781,I419846,I419834);
and I_18700 (I320798,I320781,I419831);
DFFARX1 I_18701 (I320798,I2859,I320730,I320824,);
DFFARX1 I_18702 (I320824,I2859,I320730,I320719,);
DFFARX1 I_18703 (I419831,I2859,I320730,I320855,);
nand I_18704 (I320863,I320855,I419828);
not I_18705 (I320880,I320863);
DFFARX1 I_18706 (I320880,I2859,I320730,I320906,);
not I_18707 (I320914,I320906);
nor I_18708 (I320722,I320764,I320914);
DFFARX1 I_18709 (I419834,I2859,I320730,I320954,);
nor I_18710 (I320713,I320954,I320824);
nor I_18711 (I320704,I320954,I320880);
nand I_18712 (I320990,I419849,I419840);
and I_18713 (I321007,I320990,I419843);
DFFARX1 I_18714 (I321007,I2859,I320730,I321033,);
not I_18715 (I321041,I321033);
nand I_18716 (I321058,I321041,I320954);
nand I_18717 (I320707,I321041,I320863);
nor I_18718 (I321089,I419828,I419840);
and I_18719 (I321106,I320954,I321089);
nor I_18720 (I321123,I321041,I321106);
DFFARX1 I_18721 (I321123,I2859,I320730,I320716,);
nor I_18722 (I321154,I320756,I321089);
DFFARX1 I_18723 (I321154,I2859,I320730,I320701,);
nor I_18724 (I321185,I321033,I321089);
not I_18725 (I321202,I321185);
nand I_18726 (I320710,I321202,I321058);
not I_18727 (I321257,I2866);
DFFARX1 I_18728 (I200721,I2859,I321257,I321283,);
not I_18729 (I321291,I321283);
nand I_18730 (I321308,I200739,I200730);
and I_18731 (I321325,I321308,I200733);
DFFARX1 I_18732 (I321325,I2859,I321257,I321351,);
DFFARX1 I_18733 (I321351,I2859,I321257,I321246,);
DFFARX1 I_18734 (I200727,I2859,I321257,I321382,);
nand I_18735 (I321390,I321382,I200718);
not I_18736 (I321407,I321390);
DFFARX1 I_18737 (I321407,I2859,I321257,I321433,);
not I_18738 (I321441,I321433);
nor I_18739 (I321249,I321291,I321441);
DFFARX1 I_18740 (I200724,I2859,I321257,I321481,);
nor I_18741 (I321240,I321481,I321351);
nor I_18742 (I321231,I321481,I321407);
nand I_18743 (I321517,I200718,I200715);
and I_18744 (I321534,I321517,I200736);
DFFARX1 I_18745 (I321534,I2859,I321257,I321560,);
not I_18746 (I321568,I321560);
nand I_18747 (I321585,I321568,I321481);
nand I_18748 (I321234,I321568,I321390);
nor I_18749 (I321616,I200715,I200715);
and I_18750 (I321633,I321481,I321616);
nor I_18751 (I321650,I321568,I321633);
DFFARX1 I_18752 (I321650,I2859,I321257,I321243,);
nor I_18753 (I321681,I321283,I321616);
DFFARX1 I_18754 (I321681,I2859,I321257,I321228,);
nor I_18755 (I321712,I321560,I321616);
not I_18756 (I321729,I321712);
nand I_18757 (I321237,I321729,I321585);
not I_18758 (I321784,I2866);
DFFARX1 I_18759 (I30637,I2859,I321784,I321810,);
not I_18760 (I321818,I321810);
nand I_18761 (I321835,I30613,I30622);
and I_18762 (I321852,I321835,I30616);
DFFARX1 I_18763 (I321852,I2859,I321784,I321878,);
DFFARX1 I_18764 (I321878,I2859,I321784,I321773,);
DFFARX1 I_18765 (I30634,I2859,I321784,I321909,);
nand I_18766 (I321917,I321909,I30625);
not I_18767 (I321934,I321917);
DFFARX1 I_18768 (I321934,I2859,I321784,I321960,);
not I_18769 (I321968,I321960);
nor I_18770 (I321776,I321818,I321968);
DFFARX1 I_18771 (I30619,I2859,I321784,I322008,);
nor I_18772 (I321767,I322008,I321878);
nor I_18773 (I321758,I322008,I321934);
nand I_18774 (I322044,I30631,I30628);
and I_18775 (I322061,I322044,I30616);
DFFARX1 I_18776 (I322061,I2859,I321784,I322087,);
not I_18777 (I322095,I322087);
nand I_18778 (I322112,I322095,I322008);
nand I_18779 (I321761,I322095,I321917);
nor I_18780 (I322143,I30613,I30628);
and I_18781 (I322160,I322008,I322143);
nor I_18782 (I322177,I322095,I322160);
DFFARX1 I_18783 (I322177,I2859,I321784,I321770,);
nor I_18784 (I322208,I321810,I322143);
DFFARX1 I_18785 (I322208,I2859,I321784,I321755,);
nor I_18786 (I322239,I322087,I322143);
not I_18787 (I322256,I322239);
nand I_18788 (I321764,I322256,I322112);
not I_18789 (I322311,I2866);
DFFARX1 I_18790 (I64993,I2859,I322311,I322337,);
not I_18791 (I322345,I322337);
nand I_18792 (I322362,I64990,I65008);
and I_18793 (I322379,I322362,I64999);
DFFARX1 I_18794 (I322379,I2859,I322311,I322405,);
DFFARX1 I_18795 (I322405,I2859,I322311,I322300,);
DFFARX1 I_18796 (I65005,I2859,I322311,I322436,);
nand I_18797 (I322444,I322436,I65002);
not I_18798 (I322461,I322444);
DFFARX1 I_18799 (I322461,I2859,I322311,I322487,);
not I_18800 (I322495,I322487);
nor I_18801 (I322303,I322345,I322495);
DFFARX1 I_18802 (I64996,I2859,I322311,I322535,);
nor I_18803 (I322294,I322535,I322405);
nor I_18804 (I322285,I322535,I322461);
nand I_18805 (I322571,I64987,I65011);
and I_18806 (I322588,I322571,I64990);
DFFARX1 I_18807 (I322588,I2859,I322311,I322614,);
not I_18808 (I322622,I322614);
nand I_18809 (I322639,I322622,I322535);
nand I_18810 (I322288,I322622,I322444);
nor I_18811 (I322670,I64987,I65011);
and I_18812 (I322687,I322535,I322670);
nor I_18813 (I322704,I322622,I322687);
DFFARX1 I_18814 (I322704,I2859,I322311,I322297,);
nor I_18815 (I322735,I322337,I322670);
DFFARX1 I_18816 (I322735,I2859,I322311,I322282,);
nor I_18817 (I322766,I322614,I322670);
not I_18818 (I322783,I322766);
nand I_18819 (I322291,I322783,I322639);
not I_18820 (I322838,I2866);
DFFARX1 I_18821 (I542175,I2859,I322838,I322864,);
not I_18822 (I322872,I322864);
nand I_18823 (I322889,I542172,I542181);
and I_18824 (I322906,I322889,I542160);
DFFARX1 I_18825 (I322906,I2859,I322838,I322932,);
DFFARX1 I_18826 (I322932,I2859,I322838,I322827,);
DFFARX1 I_18827 (I542163,I2859,I322838,I322963,);
nand I_18828 (I322971,I322963,I542178);
not I_18829 (I322988,I322971);
DFFARX1 I_18830 (I322988,I2859,I322838,I323014,);
not I_18831 (I323022,I323014);
nor I_18832 (I322830,I322872,I323022);
DFFARX1 I_18833 (I542184,I2859,I322838,I323062,);
nor I_18834 (I322821,I323062,I322932);
nor I_18835 (I322812,I323062,I322988);
nand I_18836 (I323098,I542166,I542187);
and I_18837 (I323115,I323098,I542169);
DFFARX1 I_18838 (I323115,I2859,I322838,I323141,);
not I_18839 (I323149,I323141);
nand I_18840 (I323166,I323149,I323062);
nand I_18841 (I322815,I323149,I322971);
nor I_18842 (I323197,I542160,I542187);
and I_18843 (I323214,I323062,I323197);
nor I_18844 (I323231,I323149,I323214);
DFFARX1 I_18845 (I323231,I2859,I322838,I322824,);
nor I_18846 (I323262,I322864,I323197);
DFFARX1 I_18847 (I323262,I2859,I322838,I322809,);
nor I_18848 (I323293,I323141,I323197);
not I_18849 (I323310,I323293);
nand I_18850 (I322818,I323310,I323166);
not I_18851 (I323365,I2866);
DFFARX1 I_18852 (I104263,I2859,I323365,I323391,);
not I_18853 (I323399,I323391);
nand I_18854 (I323416,I104260,I104278);
and I_18855 (I323433,I323416,I104269);
DFFARX1 I_18856 (I323433,I2859,I323365,I323459,);
DFFARX1 I_18857 (I323459,I2859,I323365,I323354,);
DFFARX1 I_18858 (I104275,I2859,I323365,I323490,);
nand I_18859 (I323498,I323490,I104272);
not I_18860 (I323515,I323498);
DFFARX1 I_18861 (I323515,I2859,I323365,I323541,);
not I_18862 (I323549,I323541);
nor I_18863 (I323357,I323399,I323549);
DFFARX1 I_18864 (I104266,I2859,I323365,I323589,);
nor I_18865 (I323348,I323589,I323459);
nor I_18866 (I323339,I323589,I323515);
nand I_18867 (I323625,I104257,I104281);
and I_18868 (I323642,I323625,I104260);
DFFARX1 I_18869 (I323642,I2859,I323365,I323668,);
not I_18870 (I323676,I323668);
nand I_18871 (I323693,I323676,I323589);
nand I_18872 (I323342,I323676,I323498);
nor I_18873 (I323724,I104257,I104281);
and I_18874 (I323741,I323589,I323724);
nor I_18875 (I323758,I323676,I323741);
DFFARX1 I_18876 (I323758,I2859,I323365,I323351,);
nor I_18877 (I323789,I323391,I323724);
DFFARX1 I_18878 (I323789,I2859,I323365,I323336,);
nor I_18879 (I323820,I323668,I323724);
not I_18880 (I323837,I323820);
nand I_18881 (I323345,I323837,I323693);
not I_18882 (I323892,I2866);
DFFARX1 I_18883 (I283386,I2859,I323892,I323918,);
not I_18884 (I323926,I323918);
nand I_18885 (I323943,I283389,I283386);
and I_18886 (I323960,I323943,I283398);
DFFARX1 I_18887 (I323960,I2859,I323892,I323986,);
DFFARX1 I_18888 (I323986,I2859,I323892,I323881,);
DFFARX1 I_18889 (I283395,I2859,I323892,I324017,);
nand I_18890 (I324025,I324017,I283401);
not I_18891 (I324042,I324025);
DFFARX1 I_18892 (I324042,I2859,I323892,I324068,);
not I_18893 (I324076,I324068);
nor I_18894 (I323884,I323926,I324076);
DFFARX1 I_18895 (I283410,I2859,I323892,I324116,);
nor I_18896 (I323875,I324116,I323986);
nor I_18897 (I323866,I324116,I324042);
nand I_18898 (I324152,I283404,I283392);
and I_18899 (I324169,I324152,I283389);
DFFARX1 I_18900 (I324169,I2859,I323892,I324195,);
not I_18901 (I324203,I324195);
nand I_18902 (I324220,I324203,I324116);
nand I_18903 (I323869,I324203,I324025);
nor I_18904 (I324251,I283407,I283392);
and I_18905 (I324268,I324116,I324251);
nor I_18906 (I324285,I324203,I324268);
DFFARX1 I_18907 (I324285,I2859,I323892,I323878,);
nor I_18908 (I324316,I323918,I324251);
DFFARX1 I_18909 (I324316,I2859,I323892,I323863,);
nor I_18910 (I324347,I324195,I324251);
not I_18911 (I324364,I324347);
nand I_18912 (I323872,I324364,I324220);
not I_18913 (I324419,I2866);
DFFARX1 I_18914 (I247565,I2859,I324419,I324445,);
not I_18915 (I324453,I324445);
nand I_18916 (I324470,I247550,I247571);
and I_18917 (I324487,I324470,I247559);
DFFARX1 I_18918 (I324487,I2859,I324419,I324513,);
DFFARX1 I_18919 (I324513,I2859,I324419,I324408,);
DFFARX1 I_18920 (I247553,I2859,I324419,I324544,);
nand I_18921 (I324552,I324544,I247562);
not I_18922 (I324569,I324552);
DFFARX1 I_18923 (I324569,I2859,I324419,I324595,);
not I_18924 (I324603,I324595);
nor I_18925 (I324411,I324453,I324603);
DFFARX1 I_18926 (I247568,I2859,I324419,I324643,);
nor I_18927 (I324402,I324643,I324513);
nor I_18928 (I324393,I324643,I324569);
nand I_18929 (I324679,I247550,I247553);
and I_18930 (I324696,I324679,I247574);
DFFARX1 I_18931 (I324696,I2859,I324419,I324722,);
not I_18932 (I324730,I324722);
nand I_18933 (I324747,I324730,I324643);
nand I_18934 (I324396,I324730,I324552);
nor I_18935 (I324778,I247556,I247553);
and I_18936 (I324795,I324643,I324778);
nor I_18937 (I324812,I324730,I324795);
DFFARX1 I_18938 (I324812,I2859,I324419,I324405,);
nor I_18939 (I324843,I324445,I324778);
DFFARX1 I_18940 (I324843,I2859,I324419,I324390,);
nor I_18941 (I324874,I324722,I324778);
not I_18942 (I324891,I324874);
nand I_18943 (I324399,I324891,I324747);
not I_18944 (I324946,I2866);
DFFARX1 I_18945 (I473600,I2859,I324946,I324972,);
not I_18946 (I324980,I324972);
nand I_18947 (I324997,I473582,I473582);
and I_18948 (I325014,I324997,I473588);
DFFARX1 I_18949 (I325014,I2859,I324946,I325040,);
DFFARX1 I_18950 (I325040,I2859,I324946,I324935,);
DFFARX1 I_18951 (I473585,I2859,I324946,I325071,);
nand I_18952 (I325079,I325071,I473594);
not I_18953 (I325096,I325079);
DFFARX1 I_18954 (I325096,I2859,I324946,I325122,);
not I_18955 (I325130,I325122);
nor I_18956 (I324938,I324980,I325130);
DFFARX1 I_18957 (I473606,I2859,I324946,I325170,);
nor I_18958 (I324929,I325170,I325040);
nor I_18959 (I324920,I325170,I325096);
nand I_18960 (I325206,I473597,I473591);
and I_18961 (I325223,I325206,I473585);
DFFARX1 I_18962 (I325223,I2859,I324946,I325249,);
not I_18963 (I325257,I325249);
nand I_18964 (I325274,I325257,I325170);
nand I_18965 (I324923,I325257,I325079);
nor I_18966 (I325305,I473603,I473591);
and I_18967 (I325322,I325170,I325305);
nor I_18968 (I325339,I325257,I325322);
DFFARX1 I_18969 (I325339,I2859,I324946,I324932,);
nor I_18970 (I325370,I324972,I325305);
DFFARX1 I_18971 (I325370,I2859,I324946,I324917,);
nor I_18972 (I325401,I325249,I325305);
not I_18973 (I325418,I325401);
nand I_18974 (I324926,I325418,I325274);
not I_18975 (I325473,I2866);
DFFARX1 I_18976 (I565380,I2859,I325473,I325499,);
not I_18977 (I325507,I325499);
nand I_18978 (I325524,I565377,I565386);
and I_18979 (I325541,I325524,I565365);
DFFARX1 I_18980 (I325541,I2859,I325473,I325567,);
DFFARX1 I_18981 (I325567,I2859,I325473,I325462,);
DFFARX1 I_18982 (I565368,I2859,I325473,I325598,);
nand I_18983 (I325606,I325598,I565383);
not I_18984 (I325623,I325606);
DFFARX1 I_18985 (I325623,I2859,I325473,I325649,);
not I_18986 (I325657,I325649);
nor I_18987 (I325465,I325507,I325657);
DFFARX1 I_18988 (I565389,I2859,I325473,I325697,);
nor I_18989 (I325456,I325697,I325567);
nor I_18990 (I325447,I325697,I325623);
nand I_18991 (I325733,I565371,I565392);
and I_18992 (I325750,I325733,I565374);
DFFARX1 I_18993 (I325750,I2859,I325473,I325776,);
not I_18994 (I325784,I325776);
nand I_18995 (I325801,I325784,I325697);
nand I_18996 (I325450,I325784,I325606);
nor I_18997 (I325832,I565365,I565392);
and I_18998 (I325849,I325697,I325832);
nor I_18999 (I325866,I325784,I325849);
DFFARX1 I_19000 (I325866,I2859,I325473,I325459,);
nor I_19001 (I325897,I325499,I325832);
DFFARX1 I_19002 (I325897,I2859,I325473,I325444,);
nor I_19003 (I325928,I325776,I325832);
not I_19004 (I325945,I325928);
nand I_19005 (I325453,I325945,I325801);
not I_19006 (I326000,I2866);
DFFARX1 I_19007 (I284542,I2859,I326000,I326026,);
not I_19008 (I326034,I326026);
nand I_19009 (I326051,I284545,I284542);
and I_19010 (I326068,I326051,I284554);
DFFARX1 I_19011 (I326068,I2859,I326000,I326094,);
DFFARX1 I_19012 (I326094,I2859,I326000,I325989,);
DFFARX1 I_19013 (I284551,I2859,I326000,I326125,);
nand I_19014 (I326133,I326125,I284557);
not I_19015 (I326150,I326133);
DFFARX1 I_19016 (I326150,I2859,I326000,I326176,);
not I_19017 (I326184,I326176);
nor I_19018 (I325992,I326034,I326184);
DFFARX1 I_19019 (I284566,I2859,I326000,I326224,);
nor I_19020 (I325983,I326224,I326094);
nor I_19021 (I325974,I326224,I326150);
nand I_19022 (I326260,I284560,I284548);
and I_19023 (I326277,I326260,I284545);
DFFARX1 I_19024 (I326277,I2859,I326000,I326303,);
not I_19025 (I326311,I326303);
nand I_19026 (I326328,I326311,I326224);
nand I_19027 (I325977,I326311,I326133);
nor I_19028 (I326359,I284563,I284548);
and I_19029 (I326376,I326224,I326359);
nor I_19030 (I326393,I326311,I326376);
DFFARX1 I_19031 (I326393,I2859,I326000,I325986,);
nor I_19032 (I326424,I326026,I326359);
DFFARX1 I_19033 (I326424,I2859,I326000,I325971,);
nor I_19034 (I326455,I326303,I326359);
not I_19035 (I326472,I326455);
nand I_19036 (I325980,I326472,I326328);
not I_19037 (I326527,I2866);
DFFARX1 I_19038 (I178910,I2859,I326527,I326553,);
not I_19039 (I326561,I326553);
nand I_19040 (I326578,I178907,I178916);
and I_19041 (I326595,I326578,I178925);
DFFARX1 I_19042 (I326595,I2859,I326527,I326621,);
DFFARX1 I_19043 (I326621,I2859,I326527,I326516,);
DFFARX1 I_19044 (I178928,I2859,I326527,I326652,);
nand I_19045 (I326660,I326652,I178931);
not I_19046 (I326677,I326660);
DFFARX1 I_19047 (I326677,I2859,I326527,I326703,);
not I_19048 (I326711,I326703);
nor I_19049 (I326519,I326561,I326711);
DFFARX1 I_19050 (I178904,I2859,I326527,I326751,);
nor I_19051 (I326510,I326751,I326621);
nor I_19052 (I326501,I326751,I326677);
nand I_19053 (I326787,I178919,I178922);
and I_19054 (I326804,I326787,I178913);
DFFARX1 I_19055 (I326804,I2859,I326527,I326830,);
not I_19056 (I326838,I326830);
nand I_19057 (I326855,I326838,I326751);
nand I_19058 (I326504,I326838,I326660);
nor I_19059 (I326886,I178904,I178922);
and I_19060 (I326903,I326751,I326886);
nor I_19061 (I326920,I326838,I326903);
DFFARX1 I_19062 (I326920,I2859,I326527,I326513,);
nor I_19063 (I326951,I326553,I326886);
DFFARX1 I_19064 (I326951,I2859,I326527,I326498,);
nor I_19065 (I326982,I326830,I326886);
not I_19066 (I326999,I326982);
nand I_19067 (I326507,I326999,I326855);
not I_19068 (I327054,I2866);
DFFARX1 I_19069 (I45393,I2859,I327054,I327080,);
not I_19070 (I327088,I327080);
nand I_19071 (I327105,I45369,I45378);
and I_19072 (I327122,I327105,I45372);
DFFARX1 I_19073 (I327122,I2859,I327054,I327148,);
DFFARX1 I_19074 (I327148,I2859,I327054,I327043,);
DFFARX1 I_19075 (I45390,I2859,I327054,I327179,);
nand I_19076 (I327187,I327179,I45381);
not I_19077 (I327204,I327187);
DFFARX1 I_19078 (I327204,I2859,I327054,I327230,);
not I_19079 (I327238,I327230);
nor I_19080 (I327046,I327088,I327238);
DFFARX1 I_19081 (I45375,I2859,I327054,I327278,);
nor I_19082 (I327037,I327278,I327148);
nor I_19083 (I327028,I327278,I327204);
nand I_19084 (I327314,I45387,I45384);
and I_19085 (I327331,I327314,I45372);
DFFARX1 I_19086 (I327331,I2859,I327054,I327357,);
not I_19087 (I327365,I327357);
nand I_19088 (I327382,I327365,I327278);
nand I_19089 (I327031,I327365,I327187);
nor I_19090 (I327413,I45369,I45384);
and I_19091 (I327430,I327278,I327413);
nor I_19092 (I327447,I327365,I327430);
DFFARX1 I_19093 (I327447,I2859,I327054,I327040,);
nor I_19094 (I327478,I327080,I327413);
DFFARX1 I_19095 (I327478,I2859,I327054,I327025,);
nor I_19096 (I327509,I327357,I327413);
not I_19097 (I327526,I327509);
nand I_19098 (I327034,I327526,I327382);
not I_19099 (I327581,I2866);
DFFARX1 I_19100 (I563000,I2859,I327581,I327607,);
not I_19101 (I327615,I327607);
nand I_19102 (I327632,I562997,I563006);
and I_19103 (I327649,I327632,I562985);
DFFARX1 I_19104 (I327649,I2859,I327581,I327675,);
DFFARX1 I_19105 (I327675,I2859,I327581,I327570,);
DFFARX1 I_19106 (I562988,I2859,I327581,I327706,);
nand I_19107 (I327714,I327706,I563003);
not I_19108 (I327731,I327714);
DFFARX1 I_19109 (I327731,I2859,I327581,I327757,);
not I_19110 (I327765,I327757);
nor I_19111 (I327573,I327615,I327765);
DFFARX1 I_19112 (I563009,I2859,I327581,I327805,);
nor I_19113 (I327564,I327805,I327675);
nor I_19114 (I327555,I327805,I327731);
nand I_19115 (I327841,I562991,I563012);
and I_19116 (I327858,I327841,I562994);
DFFARX1 I_19117 (I327858,I2859,I327581,I327884,);
not I_19118 (I327892,I327884);
nand I_19119 (I327909,I327892,I327805);
nand I_19120 (I327558,I327892,I327714);
nor I_19121 (I327940,I562985,I563012);
and I_19122 (I327957,I327805,I327940);
nor I_19123 (I327974,I327892,I327957);
DFFARX1 I_19124 (I327974,I2859,I327581,I327567,);
nor I_19125 (I328005,I327607,I327940);
DFFARX1 I_19126 (I328005,I2859,I327581,I327552,);
nor I_19127 (I328036,I327884,I327940);
not I_19128 (I328053,I328036);
nand I_19129 (I327561,I328053,I327909);
not I_19130 (I328108,I2866);
DFFARX1 I_19131 (I385712,I2859,I328108,I328134,);
not I_19132 (I328142,I328134);
nand I_19133 (I328159,I385727,I385709);
and I_19134 (I328176,I328159,I385709);
DFFARX1 I_19135 (I328176,I2859,I328108,I328202,);
DFFARX1 I_19136 (I328202,I2859,I328108,I328097,);
DFFARX1 I_19137 (I385718,I2859,I328108,I328233,);
nand I_19138 (I328241,I328233,I385736);
not I_19139 (I328258,I328241);
DFFARX1 I_19140 (I328258,I2859,I328108,I328284,);
not I_19141 (I328292,I328284);
nor I_19142 (I328100,I328142,I328292);
DFFARX1 I_19143 (I385733,I2859,I328108,I328332,);
nor I_19144 (I328091,I328332,I328202);
nor I_19145 (I328082,I328332,I328258);
nand I_19146 (I328368,I385730,I385721);
and I_19147 (I328385,I328368,I385715);
DFFARX1 I_19148 (I328385,I2859,I328108,I328411,);
not I_19149 (I328419,I328411);
nand I_19150 (I328436,I328419,I328332);
nand I_19151 (I328085,I328419,I328241);
nor I_19152 (I328467,I385724,I385721);
and I_19153 (I328484,I328332,I328467);
nor I_19154 (I328501,I328419,I328484);
DFFARX1 I_19155 (I328501,I2859,I328108,I328094,);
nor I_19156 (I328532,I328134,I328467);
DFFARX1 I_19157 (I328532,I2859,I328108,I328079,);
nor I_19158 (I328563,I328411,I328467);
not I_19159 (I328580,I328563);
nand I_19160 (I328088,I328580,I328436);
not I_19161 (I328635,I2866);
DFFARX1 I_19162 (I547530,I2859,I328635,I328661,);
not I_19163 (I328669,I328661);
nand I_19164 (I328686,I547527,I547536);
and I_19165 (I328703,I328686,I547515);
DFFARX1 I_19166 (I328703,I2859,I328635,I328729,);
DFFARX1 I_19167 (I328729,I2859,I328635,I328624,);
DFFARX1 I_19168 (I547518,I2859,I328635,I328760,);
nand I_19169 (I328768,I328760,I547533);
not I_19170 (I328785,I328768);
DFFARX1 I_19171 (I328785,I2859,I328635,I328811,);
not I_19172 (I328819,I328811);
nor I_19173 (I328627,I328669,I328819);
DFFARX1 I_19174 (I547539,I2859,I328635,I328859,);
nor I_19175 (I328618,I328859,I328729);
nor I_19176 (I328609,I328859,I328785);
nand I_19177 (I328895,I547521,I547542);
and I_19178 (I328912,I328895,I547524);
DFFARX1 I_19179 (I328912,I2859,I328635,I328938,);
not I_19180 (I328946,I328938);
nand I_19181 (I328963,I328946,I328859);
nand I_19182 (I328612,I328946,I328768);
nor I_19183 (I328994,I547515,I547542);
and I_19184 (I329011,I328859,I328994);
nor I_19185 (I329028,I328946,I329011);
DFFARX1 I_19186 (I329028,I2859,I328635,I328621,);
nor I_19187 (I329059,I328661,I328994);
DFFARX1 I_19188 (I329059,I2859,I328635,I328606,);
nor I_19189 (I329090,I328938,I328994);
not I_19190 (I329107,I329090);
nand I_19191 (I328615,I329107,I328963);
not I_19192 (I329162,I2866);
DFFARX1 I_19193 (I50136,I2859,I329162,I329188,);
not I_19194 (I329196,I329188);
nand I_19195 (I329213,I50112,I50130);
and I_19196 (I329230,I329213,I50118);
DFFARX1 I_19197 (I329230,I2859,I329162,I329256,);
DFFARX1 I_19198 (I329256,I2859,I329162,I329151,);
DFFARX1 I_19199 (I50127,I2859,I329162,I329287,);
nand I_19200 (I329295,I329287,I50133);
not I_19201 (I329312,I329295);
DFFARX1 I_19202 (I329312,I2859,I329162,I329338,);
not I_19203 (I329346,I329338);
nor I_19204 (I329154,I329196,I329346);
DFFARX1 I_19205 (I50112,I2859,I329162,I329386,);
nor I_19206 (I329145,I329386,I329256);
nor I_19207 (I329136,I329386,I329312);
nand I_19208 (I329422,I50124,I50115);
and I_19209 (I329439,I329422,I50139);
DFFARX1 I_19210 (I329439,I2859,I329162,I329465,);
not I_19211 (I329473,I329465);
nand I_19212 (I329490,I329473,I329386);
nand I_19213 (I329139,I329473,I329295);
nor I_19214 (I329521,I50121,I50115);
and I_19215 (I329538,I329386,I329521);
nor I_19216 (I329555,I329473,I329538);
DFFARX1 I_19217 (I329555,I2859,I329162,I329148,);
nor I_19218 (I329586,I329188,I329521);
DFFARX1 I_19219 (I329586,I2859,I329162,I329133,);
nor I_19220 (I329617,I329465,I329521);
not I_19221 (I329634,I329617);
nand I_19222 (I329142,I329634,I329490);
not I_19223 (I329689,I2866);
DFFARX1 I_19224 (I2492,I2859,I329689,I329715,);
not I_19225 (I329723,I329715);
nand I_19226 (I329740,I1908,I1676);
and I_19227 (I329757,I329740,I2564);
DFFARX1 I_19228 (I329757,I2859,I329689,I329783,);
DFFARX1 I_19229 (I329783,I2859,I329689,I329678,);
DFFARX1 I_19230 (I2844,I2859,I329689,I329814,);
nand I_19231 (I329822,I329814,I2220);
not I_19232 (I329839,I329822);
DFFARX1 I_19233 (I329839,I2859,I329689,I329865,);
not I_19234 (I329873,I329865);
nor I_19235 (I329681,I329723,I329873);
DFFARX1 I_19236 (I2580,I2859,I329689,I329913,);
nor I_19237 (I329672,I329913,I329783);
nor I_19238 (I329663,I329913,I329839);
nand I_19239 (I329949,I2028,I1900);
and I_19240 (I329966,I329949,I1452);
DFFARX1 I_19241 (I329966,I2859,I329689,I329992,);
not I_19242 (I330000,I329992);
nand I_19243 (I330017,I330000,I329913);
nand I_19244 (I329666,I330000,I329822);
nor I_19245 (I330048,I2228,I1900);
and I_19246 (I330065,I329913,I330048);
nor I_19247 (I330082,I330000,I330065);
DFFARX1 I_19248 (I330082,I2859,I329689,I329675,);
nor I_19249 (I330113,I329715,I330048);
DFFARX1 I_19250 (I330113,I2859,I329689,I329660,);
nor I_19251 (I330144,I329992,I330048);
not I_19252 (I330161,I330144);
nand I_19253 (I329669,I330161,I330017);
not I_19254 (I330216,I2866);
DFFARX1 I_19255 (I427691,I2859,I330216,I330242,);
not I_19256 (I330250,I330242);
nand I_19257 (I330267,I427700,I427688);
and I_19258 (I330284,I330267,I427685);
DFFARX1 I_19259 (I330284,I2859,I330216,I330310,);
DFFARX1 I_19260 (I330310,I2859,I330216,I330205,);
DFFARX1 I_19261 (I427685,I2859,I330216,I330341,);
nand I_19262 (I330349,I330341,I427682);
not I_19263 (I330366,I330349);
DFFARX1 I_19264 (I330366,I2859,I330216,I330392,);
not I_19265 (I330400,I330392);
nor I_19266 (I330208,I330250,I330400);
DFFARX1 I_19267 (I427688,I2859,I330216,I330440,);
nor I_19268 (I330199,I330440,I330310);
nor I_19269 (I330190,I330440,I330366);
nand I_19270 (I330476,I427703,I427694);
and I_19271 (I330493,I330476,I427697);
DFFARX1 I_19272 (I330493,I2859,I330216,I330519,);
not I_19273 (I330527,I330519);
nand I_19274 (I330544,I330527,I330440);
nand I_19275 (I330193,I330527,I330349);
nor I_19276 (I330575,I427682,I427694);
and I_19277 (I330592,I330440,I330575);
nor I_19278 (I330609,I330527,I330592);
DFFARX1 I_19279 (I330609,I2859,I330216,I330202,);
nor I_19280 (I330640,I330242,I330575);
DFFARX1 I_19281 (I330640,I2859,I330216,I330187,);
nor I_19282 (I330671,I330519,I330575);
not I_19283 (I330688,I330671);
nand I_19284 (I330196,I330688,I330544);
not I_19285 (I330743,I2866);
DFFARX1 I_19286 (I216786,I2859,I330743,I330769,);
not I_19287 (I330777,I330769);
nand I_19288 (I330794,I216804,I216795);
and I_19289 (I330811,I330794,I216798);
DFFARX1 I_19290 (I330811,I2859,I330743,I330837,);
DFFARX1 I_19291 (I330837,I2859,I330743,I330732,);
DFFARX1 I_19292 (I216792,I2859,I330743,I330868,);
nand I_19293 (I330876,I330868,I216783);
not I_19294 (I330893,I330876);
DFFARX1 I_19295 (I330893,I2859,I330743,I330919,);
not I_19296 (I330927,I330919);
nor I_19297 (I330735,I330777,I330927);
DFFARX1 I_19298 (I216789,I2859,I330743,I330967,);
nor I_19299 (I330726,I330967,I330837);
nor I_19300 (I330717,I330967,I330893);
nand I_19301 (I331003,I216783,I216780);
and I_19302 (I331020,I331003,I216801);
DFFARX1 I_19303 (I331020,I2859,I330743,I331046,);
not I_19304 (I331054,I331046);
nand I_19305 (I331071,I331054,I330967);
nand I_19306 (I330720,I331054,I330876);
nor I_19307 (I331102,I216780,I216780);
and I_19308 (I331119,I330967,I331102);
nor I_19309 (I331136,I331054,I331119);
DFFARX1 I_19310 (I331136,I2859,I330743,I330729,);
nor I_19311 (I331167,I330769,I331102);
DFFARX1 I_19312 (I331167,I2859,I330743,I330714,);
nor I_19313 (I331198,I331046,I331102);
not I_19314 (I331215,I331198);
nand I_19315 (I330723,I331215,I331071);
not I_19316 (I331270,I2866);
DFFARX1 I_19317 (I309974,I2859,I331270,I331296,);
not I_19318 (I331304,I331296);
nand I_19319 (I331321,I309977,I309974);
and I_19320 (I331338,I331321,I309986);
DFFARX1 I_19321 (I331338,I2859,I331270,I331364,);
DFFARX1 I_19322 (I331364,I2859,I331270,I331259,);
DFFARX1 I_19323 (I309983,I2859,I331270,I331395,);
nand I_19324 (I331403,I331395,I309989);
not I_19325 (I331420,I331403);
DFFARX1 I_19326 (I331420,I2859,I331270,I331446,);
not I_19327 (I331454,I331446);
nor I_19328 (I331262,I331304,I331454);
DFFARX1 I_19329 (I309998,I2859,I331270,I331494,);
nor I_19330 (I331253,I331494,I331364);
nor I_19331 (I331244,I331494,I331420);
nand I_19332 (I331530,I309992,I309980);
and I_19333 (I331547,I331530,I309977);
DFFARX1 I_19334 (I331547,I2859,I331270,I331573,);
not I_19335 (I331581,I331573);
nand I_19336 (I331598,I331581,I331494);
nand I_19337 (I331247,I331581,I331403);
nor I_19338 (I331629,I309995,I309980);
and I_19339 (I331646,I331494,I331629);
nor I_19340 (I331663,I331581,I331646);
DFFARX1 I_19341 (I331663,I2859,I331270,I331256,);
nor I_19342 (I331694,I331296,I331629);
DFFARX1 I_19343 (I331694,I2859,I331270,I331241,);
nor I_19344 (I331725,I331573,I331629);
not I_19345 (I331742,I331725);
nand I_19346 (I331250,I331742,I331598);
not I_19347 (I331797,I2866);
DFFARX1 I_19348 (I573115,I2859,I331797,I331823,);
not I_19349 (I331831,I331823);
nand I_19350 (I331848,I573112,I573121);
and I_19351 (I331865,I331848,I573100);
DFFARX1 I_19352 (I331865,I2859,I331797,I331891,);
DFFARX1 I_19353 (I331891,I2859,I331797,I331786,);
DFFARX1 I_19354 (I573103,I2859,I331797,I331922,);
nand I_19355 (I331930,I331922,I573118);
not I_19356 (I331947,I331930);
DFFARX1 I_19357 (I331947,I2859,I331797,I331973,);
not I_19358 (I331981,I331973);
nor I_19359 (I331789,I331831,I331981);
DFFARX1 I_19360 (I573124,I2859,I331797,I332021,);
nor I_19361 (I331780,I332021,I331891);
nor I_19362 (I331771,I332021,I331947);
nand I_19363 (I332057,I573106,I573127);
and I_19364 (I332074,I332057,I573109);
DFFARX1 I_19365 (I332074,I2859,I331797,I332100,);
not I_19366 (I332108,I332100);
nand I_19367 (I332125,I332108,I332021);
nand I_19368 (I331774,I332108,I331930);
nor I_19369 (I332156,I573100,I573127);
and I_19370 (I332173,I332021,I332156);
nor I_19371 (I332190,I332108,I332173);
DFFARX1 I_19372 (I332190,I2859,I331797,I331783,);
nor I_19373 (I332221,I331823,I332156);
DFFARX1 I_19374 (I332221,I2859,I331797,I331768,);
nor I_19375 (I332252,I332100,I332156);
not I_19376 (I332269,I332252);
nand I_19377 (I331777,I332269,I332125);
not I_19378 (I332324,I2866);
DFFARX1 I_19379 (I60828,I2859,I332324,I332350,);
not I_19380 (I332358,I332350);
nand I_19381 (I332375,I60825,I60843);
and I_19382 (I332392,I332375,I60834);
DFFARX1 I_19383 (I332392,I2859,I332324,I332418,);
DFFARX1 I_19384 (I332418,I2859,I332324,I332313,);
DFFARX1 I_19385 (I60840,I2859,I332324,I332449,);
nand I_19386 (I332457,I332449,I60837);
not I_19387 (I332474,I332457);
DFFARX1 I_19388 (I332474,I2859,I332324,I332500,);
not I_19389 (I332508,I332500);
nor I_19390 (I332316,I332358,I332508);
DFFARX1 I_19391 (I60831,I2859,I332324,I332548,);
nor I_19392 (I332307,I332548,I332418);
nor I_19393 (I332298,I332548,I332474);
nand I_19394 (I332584,I60822,I60846);
and I_19395 (I332601,I332584,I60825);
DFFARX1 I_19396 (I332601,I2859,I332324,I332627,);
not I_19397 (I332635,I332627);
nand I_19398 (I332652,I332635,I332548);
nand I_19399 (I332301,I332635,I332457);
nor I_19400 (I332683,I60822,I60846);
and I_19401 (I332700,I332548,I332683);
nor I_19402 (I332717,I332635,I332700);
DFFARX1 I_19403 (I332717,I2859,I332324,I332310,);
nor I_19404 (I332748,I332350,I332683);
DFFARX1 I_19405 (I332748,I2859,I332324,I332295,);
nor I_19406 (I332779,I332627,I332683);
not I_19407 (I332796,I332779);
nand I_19408 (I332304,I332796,I332652);
not I_19409 (I332851,I2866);
DFFARX1 I_19410 (I220356,I2859,I332851,I332877,);
not I_19411 (I332885,I332877);
nand I_19412 (I332902,I220374,I220365);
and I_19413 (I332919,I332902,I220368);
DFFARX1 I_19414 (I332919,I2859,I332851,I332945,);
DFFARX1 I_19415 (I332945,I2859,I332851,I332840,);
DFFARX1 I_19416 (I220362,I2859,I332851,I332976,);
nand I_19417 (I332984,I332976,I220353);
not I_19418 (I333001,I332984);
DFFARX1 I_19419 (I333001,I2859,I332851,I333027,);
not I_19420 (I333035,I333027);
nor I_19421 (I332843,I332885,I333035);
DFFARX1 I_19422 (I220359,I2859,I332851,I333075,);
nor I_19423 (I332834,I333075,I332945);
nor I_19424 (I332825,I333075,I333001);
nand I_19425 (I333111,I220353,I220350);
and I_19426 (I333128,I333111,I220371);
DFFARX1 I_19427 (I333128,I2859,I332851,I333154,);
not I_19428 (I333162,I333154);
nand I_19429 (I333179,I333162,I333075);
nand I_19430 (I332828,I333162,I332984);
nor I_19431 (I333210,I220350,I220350);
and I_19432 (I333227,I333075,I333210);
nor I_19433 (I333244,I333162,I333227);
DFFARX1 I_19434 (I333244,I2859,I332851,I332837,);
nor I_19435 (I333275,I332877,I333210);
DFFARX1 I_19436 (I333275,I2859,I332851,I332822,);
nor I_19437 (I333306,I333154,I333210);
not I_19438 (I333323,I333306);
nand I_19439 (I332831,I333323,I333179);
not I_19440 (I333378,I2866);
DFFARX1 I_19441 (I480536,I2859,I333378,I333404,);
not I_19442 (I333412,I333404);
nand I_19443 (I333429,I480518,I480518);
and I_19444 (I333446,I333429,I480524);
DFFARX1 I_19445 (I333446,I2859,I333378,I333472,);
DFFARX1 I_19446 (I333472,I2859,I333378,I333367,);
DFFARX1 I_19447 (I480521,I2859,I333378,I333503,);
nand I_19448 (I333511,I333503,I480530);
not I_19449 (I333528,I333511);
DFFARX1 I_19450 (I333528,I2859,I333378,I333554,);
not I_19451 (I333562,I333554);
nor I_19452 (I333370,I333412,I333562);
DFFARX1 I_19453 (I480542,I2859,I333378,I333602,);
nor I_19454 (I333361,I333602,I333472);
nor I_19455 (I333352,I333602,I333528);
nand I_19456 (I333638,I480533,I480527);
and I_19457 (I333655,I333638,I480521);
DFFARX1 I_19458 (I333655,I2859,I333378,I333681,);
not I_19459 (I333689,I333681);
nand I_19460 (I333706,I333689,I333602);
nand I_19461 (I333355,I333689,I333511);
nor I_19462 (I333737,I480539,I480527);
and I_19463 (I333754,I333602,I333737);
nor I_19464 (I333771,I333689,I333754);
DFFARX1 I_19465 (I333771,I2859,I333378,I333364,);
nor I_19466 (I333802,I333404,I333737);
DFFARX1 I_19467 (I333802,I2859,I333378,I333349,);
nor I_19468 (I333833,I333681,I333737);
not I_19469 (I333850,I333833);
nand I_19470 (I333358,I333850,I333706);
not I_19471 (I333905,I2866);
DFFARX1 I_19472 (I546340,I2859,I333905,I333931,);
not I_19473 (I333939,I333931);
nand I_19474 (I333956,I546337,I546346);
and I_19475 (I333973,I333956,I546325);
DFFARX1 I_19476 (I333973,I2859,I333905,I333999,);
DFFARX1 I_19477 (I333999,I2859,I333905,I333894,);
DFFARX1 I_19478 (I546328,I2859,I333905,I334030,);
nand I_19479 (I334038,I334030,I546343);
not I_19480 (I334055,I334038);
DFFARX1 I_19481 (I334055,I2859,I333905,I334081,);
not I_19482 (I334089,I334081);
nor I_19483 (I333897,I333939,I334089);
DFFARX1 I_19484 (I546349,I2859,I333905,I334129,);
nor I_19485 (I333888,I334129,I333999);
nor I_19486 (I333879,I334129,I334055);
nand I_19487 (I334165,I546331,I546352);
and I_19488 (I334182,I334165,I546334);
DFFARX1 I_19489 (I334182,I2859,I333905,I334208,);
not I_19490 (I334216,I334208);
nand I_19491 (I334233,I334216,I334129);
nand I_19492 (I333882,I334216,I334038);
nor I_19493 (I334264,I546325,I546352);
and I_19494 (I334281,I334129,I334264);
nor I_19495 (I334298,I334216,I334281);
DFFARX1 I_19496 (I334298,I2859,I333905,I333891,);
nor I_19497 (I334329,I333931,I334264);
DFFARX1 I_19498 (I334329,I2859,I333905,I333876,);
nor I_19499 (I334360,I334208,I334264);
not I_19500 (I334377,I334360);
nand I_19501 (I333885,I334377,I334233);
not I_19502 (I334432,I2866);
DFFARX1 I_19503 (I379898,I2859,I334432,I334458,);
not I_19504 (I334466,I334458);
nand I_19505 (I334483,I379913,I379895);
and I_19506 (I334500,I334483,I379895);
DFFARX1 I_19507 (I334500,I2859,I334432,I334526,);
DFFARX1 I_19508 (I334526,I2859,I334432,I334421,);
DFFARX1 I_19509 (I379904,I2859,I334432,I334557,);
nand I_19510 (I334565,I334557,I379922);
not I_19511 (I334582,I334565);
DFFARX1 I_19512 (I334582,I2859,I334432,I334608,);
not I_19513 (I334616,I334608);
nor I_19514 (I334424,I334466,I334616);
DFFARX1 I_19515 (I379919,I2859,I334432,I334656,);
nor I_19516 (I334415,I334656,I334526);
nor I_19517 (I334406,I334656,I334582);
nand I_19518 (I334692,I379916,I379907);
and I_19519 (I334709,I334692,I379901);
DFFARX1 I_19520 (I334709,I2859,I334432,I334735,);
not I_19521 (I334743,I334735);
nand I_19522 (I334760,I334743,I334656);
nand I_19523 (I334409,I334743,I334565);
nor I_19524 (I334791,I379910,I379907);
and I_19525 (I334808,I334656,I334791);
nor I_19526 (I334825,I334743,I334808);
DFFARX1 I_19527 (I334825,I2859,I334432,I334418,);
nor I_19528 (I334856,I334458,I334791);
DFFARX1 I_19529 (I334856,I2859,I334432,I334403,);
nor I_19530 (I334887,I334735,I334791);
not I_19531 (I334904,I334887);
nand I_19532 (I334412,I334904,I334760);
not I_19533 (I334959,I2866);
DFFARX1 I_19534 (I154093,I2859,I334959,I334985,);
not I_19535 (I334993,I334985);
nand I_19536 (I335010,I154084,I154084);
and I_19537 (I335027,I335010,I154102);
DFFARX1 I_19538 (I335027,I2859,I334959,I335053,);
DFFARX1 I_19539 (I335053,I2859,I334959,I334948,);
DFFARX1 I_19540 (I154105,I2859,I334959,I335084,);
nand I_19541 (I335092,I335084,I154087);
not I_19542 (I335109,I335092);
DFFARX1 I_19543 (I335109,I2859,I334959,I335135,);
not I_19544 (I335143,I335135);
nor I_19545 (I334951,I334993,I335143);
DFFARX1 I_19546 (I154099,I2859,I334959,I335183,);
nor I_19547 (I334942,I335183,I335053);
nor I_19548 (I334933,I335183,I335109);
nand I_19549 (I335219,I154111,I154090);
and I_19550 (I335236,I335219,I154096);
DFFARX1 I_19551 (I335236,I2859,I334959,I335262,);
not I_19552 (I335270,I335262);
nand I_19553 (I335287,I335270,I335183);
nand I_19554 (I334936,I335270,I335092);
nor I_19555 (I335318,I154108,I154090);
and I_19556 (I335335,I335183,I335318);
nor I_19557 (I335352,I335270,I335335);
DFFARX1 I_19558 (I335352,I2859,I334959,I334945,);
nor I_19559 (I335383,I334985,I335318);
DFFARX1 I_19560 (I335383,I2859,I334959,I334930,);
nor I_19561 (I335414,I335262,I335318);
not I_19562 (I335431,I335414);
nand I_19563 (I334939,I335431,I335287);
not I_19564 (I335486,I2866);
DFFARX1 I_19565 (I408968,I2859,I335486,I335512,);
not I_19566 (I335520,I335512);
nand I_19567 (I335537,I408983,I408965);
and I_19568 (I335554,I335537,I408965);
DFFARX1 I_19569 (I335554,I2859,I335486,I335580,);
DFFARX1 I_19570 (I335580,I2859,I335486,I335475,);
DFFARX1 I_19571 (I408974,I2859,I335486,I335611,);
nand I_19572 (I335619,I335611,I408992);
not I_19573 (I335636,I335619);
DFFARX1 I_19574 (I335636,I2859,I335486,I335662,);
not I_19575 (I335670,I335662);
nor I_19576 (I335478,I335520,I335670);
DFFARX1 I_19577 (I408989,I2859,I335486,I335710,);
nor I_19578 (I335469,I335710,I335580);
nor I_19579 (I335460,I335710,I335636);
nand I_19580 (I335746,I408986,I408977);
and I_19581 (I335763,I335746,I408971);
DFFARX1 I_19582 (I335763,I2859,I335486,I335789,);
not I_19583 (I335797,I335789);
nand I_19584 (I335814,I335797,I335710);
nand I_19585 (I335463,I335797,I335619);
nor I_19586 (I335845,I408980,I408977);
and I_19587 (I335862,I335710,I335845);
nor I_19588 (I335879,I335797,I335862);
DFFARX1 I_19589 (I335879,I2859,I335486,I335472,);
nor I_19590 (I335910,I335512,I335845);
DFFARX1 I_19591 (I335910,I2859,I335486,I335457,);
nor I_19592 (I335941,I335789,I335845);
not I_19593 (I335958,I335941);
nand I_19594 (I335466,I335958,I335814);
not I_19595 (I336013,I2866);
DFFARX1 I_19596 (I44339,I2859,I336013,I336039,);
not I_19597 (I336047,I336039);
nand I_19598 (I336064,I44315,I44324);
and I_19599 (I336081,I336064,I44318);
DFFARX1 I_19600 (I336081,I2859,I336013,I336107,);
DFFARX1 I_19601 (I336107,I2859,I336013,I336002,);
DFFARX1 I_19602 (I44336,I2859,I336013,I336138,);
nand I_19603 (I336146,I336138,I44327);
not I_19604 (I336163,I336146);
DFFARX1 I_19605 (I336163,I2859,I336013,I336189,);
not I_19606 (I336197,I336189);
nor I_19607 (I336005,I336047,I336197);
DFFARX1 I_19608 (I44321,I2859,I336013,I336237,);
nor I_19609 (I335996,I336237,I336107);
nor I_19610 (I335987,I336237,I336163);
nand I_19611 (I336273,I44333,I44330);
and I_19612 (I336290,I336273,I44318);
DFFARX1 I_19613 (I336290,I2859,I336013,I336316,);
not I_19614 (I336324,I336316);
nand I_19615 (I336341,I336324,I336237);
nand I_19616 (I335990,I336324,I336146);
nor I_19617 (I336372,I44315,I44330);
and I_19618 (I336389,I336237,I336372);
nor I_19619 (I336406,I336324,I336389);
DFFARX1 I_19620 (I336406,I2859,I336013,I335999,);
nor I_19621 (I336437,I336039,I336372);
DFFARX1 I_19622 (I336437,I2859,I336013,I335984,);
nor I_19623 (I336468,I336316,I336372);
not I_19624 (I336485,I336468);
nand I_19625 (I335993,I336485,I336341);
not I_19626 (I336540,I2866);
DFFARX1 I_19627 (I275294,I2859,I336540,I336566,);
not I_19628 (I336574,I336566);
nand I_19629 (I336591,I275297,I275294);
and I_19630 (I336608,I336591,I275306);
DFFARX1 I_19631 (I336608,I2859,I336540,I336634,);
DFFARX1 I_19632 (I336634,I2859,I336540,I336529,);
DFFARX1 I_19633 (I275303,I2859,I336540,I336665,);
nand I_19634 (I336673,I336665,I275309);
not I_19635 (I336690,I336673);
DFFARX1 I_19636 (I336690,I2859,I336540,I336716,);
not I_19637 (I336724,I336716);
nor I_19638 (I336532,I336574,I336724);
DFFARX1 I_19639 (I275318,I2859,I336540,I336764,);
nor I_19640 (I336523,I336764,I336634);
nor I_19641 (I336514,I336764,I336690);
nand I_19642 (I336800,I275312,I275300);
and I_19643 (I336817,I336800,I275297);
DFFARX1 I_19644 (I336817,I2859,I336540,I336843,);
not I_19645 (I336851,I336843);
nand I_19646 (I336868,I336851,I336764);
nand I_19647 (I336517,I336851,I336673);
nor I_19648 (I336899,I275315,I275300);
and I_19649 (I336916,I336764,I336899);
nor I_19650 (I336933,I336851,I336916);
DFFARX1 I_19651 (I336933,I2859,I336540,I336526,);
nor I_19652 (I336964,I336566,I336899);
DFFARX1 I_19653 (I336964,I2859,I336540,I336511,);
nor I_19654 (I336995,I336843,I336899);
not I_19655 (I337012,I336995);
nand I_19656 (I336520,I337012,I336868);
not I_19657 (I337067,I2866);
DFFARX1 I_19658 (I525858,I2859,I337067,I337093,);
not I_19659 (I337101,I337093);
nand I_19660 (I337118,I525840,I525843);
and I_19661 (I337135,I337118,I525855);
DFFARX1 I_19662 (I337135,I2859,I337067,I337161,);
DFFARX1 I_19663 (I337161,I2859,I337067,I337056,);
DFFARX1 I_19664 (I525864,I2859,I337067,I337192,);
nand I_19665 (I337200,I337192,I525849);
not I_19666 (I337217,I337200);
DFFARX1 I_19667 (I337217,I2859,I337067,I337243,);
not I_19668 (I337251,I337243);
nor I_19669 (I337059,I337101,I337251);
DFFARX1 I_19670 (I525861,I2859,I337067,I337291,);
nor I_19671 (I337050,I337291,I337161);
nor I_19672 (I337041,I337291,I337217);
nand I_19673 (I337327,I525852,I525846);
and I_19674 (I337344,I337327,I525840);
DFFARX1 I_19675 (I337344,I2859,I337067,I337370,);
not I_19676 (I337378,I337370);
nand I_19677 (I337395,I337378,I337291);
nand I_19678 (I337044,I337378,I337200);
nor I_19679 (I337426,I525843,I525846);
and I_19680 (I337443,I337291,I337426);
nor I_19681 (I337460,I337378,I337443);
DFFARX1 I_19682 (I337460,I2859,I337067,I337053,);
nor I_19683 (I337491,I337093,I337426);
DFFARX1 I_19684 (I337491,I2859,I337067,I337038,);
nor I_19685 (I337522,I337370,I337426);
not I_19686 (I337539,I337522);
nand I_19687 (I337047,I337539,I337395);
not I_19688 (I337594,I2866);
DFFARX1 I_19689 (I170750,I2859,I337594,I337620,);
not I_19690 (I337628,I337620);
nand I_19691 (I337645,I170747,I170756);
and I_19692 (I337662,I337645,I170765);
DFFARX1 I_19693 (I337662,I2859,I337594,I337688,);
DFFARX1 I_19694 (I337688,I2859,I337594,I337583,);
DFFARX1 I_19695 (I170768,I2859,I337594,I337719,);
nand I_19696 (I337727,I337719,I170771);
not I_19697 (I337744,I337727);
DFFARX1 I_19698 (I337744,I2859,I337594,I337770,);
not I_19699 (I337778,I337770);
nor I_19700 (I337586,I337628,I337778);
DFFARX1 I_19701 (I170744,I2859,I337594,I337818,);
nor I_19702 (I337577,I337818,I337688);
nor I_19703 (I337568,I337818,I337744);
nand I_19704 (I337854,I170759,I170762);
and I_19705 (I337871,I337854,I170753);
DFFARX1 I_19706 (I337871,I2859,I337594,I337897,);
not I_19707 (I337905,I337897);
nand I_19708 (I337922,I337905,I337818);
nand I_19709 (I337571,I337905,I337727);
nor I_19710 (I337953,I170744,I170762);
and I_19711 (I337970,I337818,I337953);
nor I_19712 (I337987,I337905,I337970);
DFFARX1 I_19713 (I337987,I2859,I337594,I337580,);
nor I_19714 (I338018,I337620,I337953);
DFFARX1 I_19715 (I338018,I2859,I337594,I337565,);
nor I_19716 (I338049,I337897,I337953);
not I_19717 (I338066,I338049);
nand I_19718 (I337574,I338066,I337922);
not I_19719 (I338121,I2866);
DFFARX1 I_19720 (I490362,I2859,I338121,I338147,);
not I_19721 (I338155,I338147);
nand I_19722 (I338172,I490344,I490344);
and I_19723 (I338189,I338172,I490350);
DFFARX1 I_19724 (I338189,I2859,I338121,I338215,);
DFFARX1 I_19725 (I338215,I2859,I338121,I338110,);
DFFARX1 I_19726 (I490347,I2859,I338121,I338246,);
nand I_19727 (I338254,I338246,I490356);
not I_19728 (I338271,I338254);
DFFARX1 I_19729 (I338271,I2859,I338121,I338297,);
not I_19730 (I338305,I338297);
nor I_19731 (I338113,I338155,I338305);
DFFARX1 I_19732 (I490368,I2859,I338121,I338345,);
nor I_19733 (I338104,I338345,I338215);
nor I_19734 (I338095,I338345,I338271);
nand I_19735 (I338381,I490359,I490353);
and I_19736 (I338398,I338381,I490347);
DFFARX1 I_19737 (I338398,I2859,I338121,I338424,);
not I_19738 (I338432,I338424);
nand I_19739 (I338449,I338432,I338345);
nand I_19740 (I338098,I338432,I338254);
nor I_19741 (I338480,I490365,I490353);
and I_19742 (I338497,I338345,I338480);
nor I_19743 (I338514,I338432,I338497);
DFFARX1 I_19744 (I338514,I2859,I338121,I338107,);
nor I_19745 (I338545,I338147,I338480);
DFFARX1 I_19746 (I338545,I2859,I338121,I338092,);
nor I_19747 (I338576,I338424,I338480);
not I_19748 (I338593,I338576);
nand I_19749 (I338101,I338593,I338449);
not I_19750 (I338648,I2866);
DFFARX1 I_19751 (I388296,I2859,I338648,I338674,);
not I_19752 (I338682,I338674);
nand I_19753 (I338699,I388311,I388293);
and I_19754 (I338716,I338699,I388293);
DFFARX1 I_19755 (I338716,I2859,I338648,I338742,);
DFFARX1 I_19756 (I338742,I2859,I338648,I338637,);
DFFARX1 I_19757 (I388302,I2859,I338648,I338773,);
nand I_19758 (I338781,I338773,I388320);
not I_19759 (I338798,I338781);
DFFARX1 I_19760 (I338798,I2859,I338648,I338824,);
not I_19761 (I338832,I338824);
nor I_19762 (I338640,I338682,I338832);
DFFARX1 I_19763 (I388317,I2859,I338648,I338872,);
nor I_19764 (I338631,I338872,I338742);
nor I_19765 (I338622,I338872,I338798);
nand I_19766 (I338908,I388314,I388305);
and I_19767 (I338925,I338908,I388299);
DFFARX1 I_19768 (I338925,I2859,I338648,I338951,);
not I_19769 (I338959,I338951);
nand I_19770 (I338976,I338959,I338872);
nand I_19771 (I338625,I338959,I338781);
nor I_19772 (I339007,I388308,I388305);
and I_19773 (I339024,I338872,I339007);
nor I_19774 (I339041,I338959,I339024);
DFFARX1 I_19775 (I339041,I2859,I338648,I338634,);
nor I_19776 (I339072,I338674,I339007);
DFFARX1 I_19777 (I339072,I2859,I338648,I338619,);
nor I_19778 (I339103,I338951,I339007);
not I_19779 (I339120,I339103);
nand I_19780 (I338628,I339120,I338976);
not I_19781 (I339175,I2866);
DFFARX1 I_19782 (I8488,I2859,I339175,I339201,);
not I_19783 (I339209,I339201);
nand I_19784 (I339226,I8500,I8503);
and I_19785 (I339243,I339226,I8479);
DFFARX1 I_19786 (I339243,I2859,I339175,I339269,);
DFFARX1 I_19787 (I339269,I2859,I339175,I339164,);
DFFARX1 I_19788 (I8497,I2859,I339175,I339300,);
nand I_19789 (I339308,I339300,I8485);
not I_19790 (I339325,I339308);
DFFARX1 I_19791 (I339325,I2859,I339175,I339351,);
not I_19792 (I339359,I339351);
nor I_19793 (I339167,I339209,I339359);
DFFARX1 I_19794 (I8482,I2859,I339175,I339399,);
nor I_19795 (I339158,I339399,I339269);
nor I_19796 (I339149,I339399,I339325);
nand I_19797 (I339435,I8491,I8482);
and I_19798 (I339452,I339435,I8479);
DFFARX1 I_19799 (I339452,I2859,I339175,I339478,);
not I_19800 (I339486,I339478);
nand I_19801 (I339503,I339486,I339399);
nand I_19802 (I339152,I339486,I339308);
nor I_19803 (I339534,I8494,I8482);
and I_19804 (I339551,I339399,I339534);
nor I_19805 (I339568,I339486,I339551);
DFFARX1 I_19806 (I339568,I2859,I339175,I339161,);
nor I_19807 (I339599,I339201,I339534);
DFFARX1 I_19808 (I339599,I2859,I339175,I339146,);
nor I_19809 (I339630,I339478,I339534);
not I_19810 (I339647,I339630);
nand I_19811 (I339155,I339647,I339503);
not I_19812 (I339702,I2866);
DFFARX1 I_19813 (I14285,I2859,I339702,I339728,);
not I_19814 (I339736,I339728);
nand I_19815 (I339753,I14297,I14300);
and I_19816 (I339770,I339753,I14276);
DFFARX1 I_19817 (I339770,I2859,I339702,I339796,);
DFFARX1 I_19818 (I339796,I2859,I339702,I339691,);
DFFARX1 I_19819 (I14294,I2859,I339702,I339827,);
nand I_19820 (I339835,I339827,I14282);
not I_19821 (I339852,I339835);
DFFARX1 I_19822 (I339852,I2859,I339702,I339878,);
not I_19823 (I339886,I339878);
nor I_19824 (I339694,I339736,I339886);
DFFARX1 I_19825 (I14279,I2859,I339702,I339926,);
nor I_19826 (I339685,I339926,I339796);
nor I_19827 (I339676,I339926,I339852);
nand I_19828 (I339962,I14288,I14279);
and I_19829 (I339979,I339962,I14276);
DFFARX1 I_19830 (I339979,I2859,I339702,I340005,);
not I_19831 (I340013,I340005);
nand I_19832 (I340030,I340013,I339926);
nand I_19833 (I339679,I340013,I339835);
nor I_19834 (I340061,I14291,I14279);
and I_19835 (I340078,I339926,I340061);
nor I_19836 (I340095,I340013,I340078);
DFFARX1 I_19837 (I340095,I2859,I339702,I339688,);
nor I_19838 (I340126,I339728,I340061);
DFFARX1 I_19839 (I340126,I2859,I339702,I339673,);
nor I_19840 (I340157,I340005,I340061);
not I_19841 (I340174,I340157);
nand I_19842 (I339682,I340174,I340030);
not I_19843 (I340229,I2866);
DFFARX1 I_19844 (I471288,I2859,I340229,I340255,);
not I_19845 (I340263,I340255);
nand I_19846 (I340280,I471270,I471270);
and I_19847 (I340297,I340280,I471276);
DFFARX1 I_19848 (I340297,I2859,I340229,I340323,);
DFFARX1 I_19849 (I340323,I2859,I340229,I340218,);
DFFARX1 I_19850 (I471273,I2859,I340229,I340354,);
nand I_19851 (I340362,I340354,I471282);
not I_19852 (I340379,I340362);
DFFARX1 I_19853 (I340379,I2859,I340229,I340405,);
not I_19854 (I340413,I340405);
nor I_19855 (I340221,I340263,I340413);
DFFARX1 I_19856 (I471294,I2859,I340229,I340453,);
nor I_19857 (I340212,I340453,I340323);
nor I_19858 (I340203,I340453,I340379);
nand I_19859 (I340489,I471285,I471279);
and I_19860 (I340506,I340489,I471273);
DFFARX1 I_19861 (I340506,I2859,I340229,I340532,);
not I_19862 (I340540,I340532);
nand I_19863 (I340557,I340540,I340453);
nand I_19864 (I340206,I340540,I340362);
nor I_19865 (I340588,I471291,I471279);
and I_19866 (I340605,I340453,I340588);
nor I_19867 (I340622,I340540,I340605);
DFFARX1 I_19868 (I340622,I2859,I340229,I340215,);
nor I_19869 (I340653,I340255,I340588);
DFFARX1 I_19870 (I340653,I2859,I340229,I340200,);
nor I_19871 (I340684,I340532,I340588);
not I_19872 (I340701,I340684);
nand I_19873 (I340209,I340701,I340557);
not I_19874 (I340756,I2866);
DFFARX1 I_19875 (I419276,I2859,I340756,I340782,);
not I_19876 (I340790,I340782);
nand I_19877 (I340807,I419285,I419273);
and I_19878 (I340824,I340807,I419270);
DFFARX1 I_19879 (I340824,I2859,I340756,I340850,);
DFFARX1 I_19880 (I340850,I2859,I340756,I340745,);
DFFARX1 I_19881 (I419270,I2859,I340756,I340881,);
nand I_19882 (I340889,I340881,I419267);
not I_19883 (I340906,I340889);
DFFARX1 I_19884 (I340906,I2859,I340756,I340932,);
not I_19885 (I340940,I340932);
nor I_19886 (I340748,I340790,I340940);
DFFARX1 I_19887 (I419273,I2859,I340756,I340980,);
nor I_19888 (I340739,I340980,I340850);
nor I_19889 (I340730,I340980,I340906);
nand I_19890 (I341016,I419288,I419279);
and I_19891 (I341033,I341016,I419282);
DFFARX1 I_19892 (I341033,I2859,I340756,I341059,);
not I_19893 (I341067,I341059);
nand I_19894 (I341084,I341067,I340980);
nand I_19895 (I340733,I341067,I340889);
nor I_19896 (I341115,I419267,I419279);
and I_19897 (I341132,I340980,I341115);
nor I_19898 (I341149,I341067,I341132);
DFFARX1 I_19899 (I341149,I2859,I340756,I340742,);
nor I_19900 (I341180,I340782,I341115);
DFFARX1 I_19901 (I341180,I2859,I340756,I340727,);
nor I_19902 (I341211,I341059,I341115);
not I_19903 (I341228,I341211);
nand I_19904 (I340736,I341228,I341084);
not I_19905 (I341283,I2866);
DFFARX1 I_19906 (I260266,I2859,I341283,I341309,);
not I_19907 (I341317,I341309);
nand I_19908 (I341334,I260269,I260266);
and I_19909 (I341351,I341334,I260278);
DFFARX1 I_19910 (I341351,I2859,I341283,I341377,);
DFFARX1 I_19911 (I341377,I2859,I341283,I341272,);
DFFARX1 I_19912 (I260275,I2859,I341283,I341408,);
nand I_19913 (I341416,I341408,I260281);
not I_19914 (I341433,I341416);
DFFARX1 I_19915 (I341433,I2859,I341283,I341459,);
not I_19916 (I341467,I341459);
nor I_19917 (I341275,I341317,I341467);
DFFARX1 I_19918 (I260290,I2859,I341283,I341507,);
nor I_19919 (I341266,I341507,I341377);
nor I_19920 (I341257,I341507,I341433);
nand I_19921 (I341543,I260284,I260272);
and I_19922 (I341560,I341543,I260269);
DFFARX1 I_19923 (I341560,I2859,I341283,I341586,);
not I_19924 (I341594,I341586);
nand I_19925 (I341611,I341594,I341507);
nand I_19926 (I341260,I341594,I341416);
nor I_19927 (I341642,I260287,I260272);
and I_19928 (I341659,I341507,I341642);
nor I_19929 (I341676,I341594,I341659);
DFFARX1 I_19930 (I341676,I2859,I341283,I341269,);
nor I_19931 (I341707,I341309,I341642);
DFFARX1 I_19932 (I341707,I2859,I341283,I341254,);
nor I_19933 (I341738,I341586,I341642);
not I_19934 (I341755,I341738);
nand I_19935 (I341263,I341755,I341611);
not I_19936 (I341810,I2866);
DFFARX1 I_19937 (I436667,I2859,I341810,I341836,);
not I_19938 (I341844,I341836);
nand I_19939 (I341861,I436676,I436664);
and I_19940 (I341878,I341861,I436661);
DFFARX1 I_19941 (I341878,I2859,I341810,I341904,);
DFFARX1 I_19942 (I341904,I2859,I341810,I341799,);
DFFARX1 I_19943 (I436661,I2859,I341810,I341935,);
nand I_19944 (I341943,I341935,I436658);
not I_19945 (I341960,I341943);
DFFARX1 I_19946 (I341960,I2859,I341810,I341986,);
not I_19947 (I341994,I341986);
nor I_19948 (I341802,I341844,I341994);
DFFARX1 I_19949 (I436664,I2859,I341810,I342034,);
nor I_19950 (I341793,I342034,I341904);
nor I_19951 (I341784,I342034,I341960);
nand I_19952 (I342070,I436679,I436670);
and I_19953 (I342087,I342070,I436673);
DFFARX1 I_19954 (I342087,I2859,I341810,I342113,);
not I_19955 (I342121,I342113);
nand I_19956 (I342138,I342121,I342034);
nand I_19957 (I341787,I342121,I341943);
nor I_19958 (I342169,I436658,I436670);
and I_19959 (I342186,I342034,I342169);
nor I_19960 (I342203,I342121,I342186);
DFFARX1 I_19961 (I342203,I2859,I341810,I341796,);
nor I_19962 (I342234,I341836,I342169);
DFFARX1 I_19963 (I342234,I2859,I341810,I341781,);
nor I_19964 (I342265,I342113,I342169);
not I_19965 (I342282,I342265);
nand I_19966 (I341790,I342282,I342138);
not I_19967 (I342337,I2866);
DFFARX1 I_19968 (I18516,I2859,I342337,I342363,);
not I_19969 (I342371,I342363);
nand I_19970 (I342388,I18492,I18501);
and I_19971 (I342405,I342388,I18495);
DFFARX1 I_19972 (I342405,I2859,I342337,I342431,);
DFFARX1 I_19973 (I342431,I2859,I342337,I342326,);
DFFARX1 I_19974 (I18513,I2859,I342337,I342462,);
nand I_19975 (I342470,I342462,I18504);
not I_19976 (I342487,I342470);
DFFARX1 I_19977 (I342487,I2859,I342337,I342513,);
not I_19978 (I342521,I342513);
nor I_19979 (I342329,I342371,I342521);
DFFARX1 I_19980 (I18498,I2859,I342337,I342561,);
nor I_19981 (I342320,I342561,I342431);
nor I_19982 (I342311,I342561,I342487);
nand I_19983 (I342597,I18510,I18507);
and I_19984 (I342614,I342597,I18495);
DFFARX1 I_19985 (I342614,I2859,I342337,I342640,);
not I_19986 (I342648,I342640);
nand I_19987 (I342665,I342648,I342561);
nand I_19988 (I342314,I342648,I342470);
nor I_19989 (I342696,I18492,I18507);
and I_19990 (I342713,I342561,I342696);
nor I_19991 (I342730,I342648,I342713);
DFFARX1 I_19992 (I342730,I2859,I342337,I342323,);
nor I_19993 (I342761,I342363,I342696);
DFFARX1 I_19994 (I342761,I2859,I342337,I342308,);
nor I_19995 (I342792,I342640,I342696);
not I_19996 (I342809,I342792);
nand I_19997 (I342317,I342809,I342665);
not I_19998 (I342864,I2866);
DFFARX1 I_19999 (I282808,I2859,I342864,I342890,);
not I_20000 (I342898,I342890);
nand I_20001 (I342915,I282811,I282808);
and I_20002 (I342932,I342915,I282820);
DFFARX1 I_20003 (I342932,I2859,I342864,I342958,);
DFFARX1 I_20004 (I342958,I2859,I342864,I342853,);
DFFARX1 I_20005 (I282817,I2859,I342864,I342989,);
nand I_20006 (I342997,I342989,I282823);
not I_20007 (I343014,I342997);
DFFARX1 I_20008 (I343014,I2859,I342864,I343040,);
not I_20009 (I343048,I343040);
nor I_20010 (I342856,I342898,I343048);
DFFARX1 I_20011 (I282832,I2859,I342864,I343088,);
nor I_20012 (I342847,I343088,I342958);
nor I_20013 (I342838,I343088,I343014);
nand I_20014 (I343124,I282826,I282814);
and I_20015 (I343141,I343124,I282811);
DFFARX1 I_20016 (I343141,I2859,I342864,I343167,);
not I_20017 (I343175,I343167);
nand I_20018 (I343192,I343175,I343088);
nand I_20019 (I342841,I343175,I342997);
nor I_20020 (I343223,I282829,I282814);
and I_20021 (I343240,I343088,I343223);
nor I_20022 (I343257,I343175,I343240);
DFFARX1 I_20023 (I343257,I2859,I342864,I342850,);
nor I_20024 (I343288,I342890,I343223);
DFFARX1 I_20025 (I343288,I2859,I342864,I342835,);
nor I_20026 (I343319,I343167,I343223);
not I_20027 (I343336,I343319);
nand I_20028 (I342844,I343336,I343192);
not I_20029 (I343391,I2866);
DFFARX1 I_20030 (I165310,I2859,I343391,I343417,);
not I_20031 (I343425,I343417);
nand I_20032 (I343442,I165307,I165316);
and I_20033 (I343459,I343442,I165325);
DFFARX1 I_20034 (I343459,I2859,I343391,I343485,);
DFFARX1 I_20035 (I343485,I2859,I343391,I343380,);
DFFARX1 I_20036 (I165328,I2859,I343391,I343516,);
nand I_20037 (I343524,I343516,I165331);
not I_20038 (I343541,I343524);
DFFARX1 I_20039 (I343541,I2859,I343391,I343567,);
not I_20040 (I343575,I343567);
nor I_20041 (I343383,I343425,I343575);
DFFARX1 I_20042 (I165304,I2859,I343391,I343615,);
nor I_20043 (I343374,I343615,I343485);
nor I_20044 (I343365,I343615,I343541);
nand I_20045 (I343651,I165319,I165322);
and I_20046 (I343668,I343651,I165313);
DFFARX1 I_20047 (I343668,I2859,I343391,I343694,);
not I_20048 (I343702,I343694);
nand I_20049 (I343719,I343702,I343615);
nand I_20050 (I343368,I343702,I343524);
nor I_20051 (I343750,I165304,I165322);
and I_20052 (I343767,I343615,I343750);
nor I_20053 (I343784,I343702,I343767);
DFFARX1 I_20054 (I343784,I2859,I343391,I343377,);
nor I_20055 (I343815,I343417,I343750);
DFFARX1 I_20056 (I343815,I2859,I343391,I343362,);
nor I_20057 (I343846,I343694,I343750);
not I_20058 (I343863,I343846);
nand I_20059 (I343371,I343863,I343719);
not I_20060 (I343918,I2866);
DFFARX1 I_20061 (I16920,I2859,I343918,I343944,);
not I_20062 (I343952,I343944);
nand I_20063 (I343969,I16932,I16935);
and I_20064 (I343986,I343969,I16911);
DFFARX1 I_20065 (I343986,I2859,I343918,I344012,);
DFFARX1 I_20066 (I344012,I2859,I343918,I343907,);
DFFARX1 I_20067 (I16929,I2859,I343918,I344043,);
nand I_20068 (I344051,I344043,I16917);
not I_20069 (I344068,I344051);
DFFARX1 I_20070 (I344068,I2859,I343918,I344094,);
not I_20071 (I344102,I344094);
nor I_20072 (I343910,I343952,I344102);
DFFARX1 I_20073 (I16914,I2859,I343918,I344142,);
nor I_20074 (I343901,I344142,I344012);
nor I_20075 (I343892,I344142,I344068);
nand I_20076 (I344178,I16923,I16914);
and I_20077 (I344195,I344178,I16911);
DFFARX1 I_20078 (I344195,I2859,I343918,I344221,);
not I_20079 (I344229,I344221);
nand I_20080 (I344246,I344229,I344142);
nand I_20081 (I343895,I344229,I344051);
nor I_20082 (I344277,I16926,I16914);
and I_20083 (I344294,I344142,I344277);
nor I_20084 (I344311,I344229,I344294);
DFFARX1 I_20085 (I344311,I2859,I343918,I343904,);
nor I_20086 (I344342,I343944,I344277);
DFFARX1 I_20087 (I344342,I2859,I343918,I343889,);
nor I_20088 (I344373,I344221,I344277);
not I_20089 (I344390,I344373);
nand I_20090 (I343898,I344390,I344246);
not I_20091 (I344445,I2866);
DFFARX1 I_20092 (I271248,I2859,I344445,I344471,);
not I_20093 (I344479,I344471);
nand I_20094 (I344496,I271251,I271248);
and I_20095 (I344513,I344496,I271260);
DFFARX1 I_20096 (I344513,I2859,I344445,I344539,);
DFFARX1 I_20097 (I344539,I2859,I344445,I344434,);
DFFARX1 I_20098 (I271257,I2859,I344445,I344570,);
nand I_20099 (I344578,I344570,I271263);
not I_20100 (I344595,I344578);
DFFARX1 I_20101 (I344595,I2859,I344445,I344621,);
not I_20102 (I344629,I344621);
nor I_20103 (I344437,I344479,I344629);
DFFARX1 I_20104 (I271272,I2859,I344445,I344669,);
nor I_20105 (I344428,I344669,I344539);
nor I_20106 (I344419,I344669,I344595);
nand I_20107 (I344705,I271266,I271254);
and I_20108 (I344722,I344705,I271251);
DFFARX1 I_20109 (I344722,I2859,I344445,I344748,);
not I_20110 (I344756,I344748);
nand I_20111 (I344773,I344756,I344669);
nand I_20112 (I344422,I344756,I344578);
nor I_20113 (I344804,I271269,I271254);
and I_20114 (I344821,I344669,I344804);
nor I_20115 (I344838,I344756,I344821);
DFFARX1 I_20116 (I344838,I2859,I344445,I344431,);
nor I_20117 (I344869,I344471,I344804);
DFFARX1 I_20118 (I344869,I2859,I344445,I344416,);
nor I_20119 (I344900,I344748,I344804);
not I_20120 (I344917,I344900);
nand I_20121 (I344425,I344917,I344773);
not I_20122 (I344972,I2866);
DFFARX1 I_20123 (I305928,I2859,I344972,I344998,);
not I_20124 (I345006,I344998);
nand I_20125 (I345023,I305931,I305928);
and I_20126 (I345040,I345023,I305940);
DFFARX1 I_20127 (I345040,I2859,I344972,I345066,);
DFFARX1 I_20128 (I345066,I2859,I344972,I344961,);
DFFARX1 I_20129 (I305937,I2859,I344972,I345097,);
nand I_20130 (I345105,I345097,I305943);
not I_20131 (I345122,I345105);
DFFARX1 I_20132 (I345122,I2859,I344972,I345148,);
not I_20133 (I345156,I345148);
nor I_20134 (I344964,I345006,I345156);
DFFARX1 I_20135 (I305952,I2859,I344972,I345196,);
nor I_20136 (I344955,I345196,I345066);
nor I_20137 (I344946,I345196,I345122);
nand I_20138 (I345232,I305946,I305934);
and I_20139 (I345249,I345232,I305931);
DFFARX1 I_20140 (I345249,I2859,I344972,I345275,);
not I_20141 (I345283,I345275);
nand I_20142 (I345300,I345283,I345196);
nand I_20143 (I344949,I345283,I345105);
nor I_20144 (I345331,I305949,I305934);
and I_20145 (I345348,I345196,I345331);
nor I_20146 (I345365,I345283,I345348);
DFFARX1 I_20147 (I345365,I2859,I344972,I344958,);
nor I_20148 (I345396,I344998,I345331);
DFFARX1 I_20149 (I345396,I2859,I344972,I344943,);
nor I_20150 (I345427,I345275,I345331);
not I_20151 (I345444,I345427);
nand I_20152 (I344952,I345444,I345300);
not I_20153 (I345499,I2866);
DFFARX1 I_20154 (I1820,I2859,I345499,I345525,);
not I_20155 (I345533,I345525);
nand I_20156 (I345550,I2436,I1388);
and I_20157 (I345567,I345550,I2796);
DFFARX1 I_20158 (I345567,I2859,I345499,I345593,);
DFFARX1 I_20159 (I345593,I2859,I345499,I345488,);
DFFARX1 I_20160 (I1516,I2859,I345499,I345624,);
nand I_20161 (I345632,I345624,I1596);
not I_20162 (I345649,I345632);
DFFARX1 I_20163 (I345649,I2859,I345499,I345675,);
not I_20164 (I345683,I345675);
nor I_20165 (I345491,I345533,I345683);
DFFARX1 I_20166 (I1948,I2859,I345499,I345723,);
nor I_20167 (I345482,I345723,I345593);
nor I_20168 (I345473,I345723,I345649);
nand I_20169 (I345759,I2116,I1956);
and I_20170 (I345776,I345759,I2548);
DFFARX1 I_20171 (I345776,I2859,I345499,I345802,);
not I_20172 (I345810,I345802);
nand I_20173 (I345827,I345810,I345723);
nand I_20174 (I345476,I345810,I345632);
nor I_20175 (I345858,I2260,I1956);
and I_20176 (I345875,I345723,I345858);
nor I_20177 (I345892,I345810,I345875);
DFFARX1 I_20178 (I345892,I2859,I345499,I345485,);
nor I_20179 (I345923,I345525,I345858);
DFFARX1 I_20180 (I345923,I2859,I345499,I345470,);
nor I_20181 (I345954,I345802,I345858);
not I_20182 (I345971,I345954);
nand I_20183 (I345479,I345971,I345827);
not I_20184 (I346026,I2866);
DFFARX1 I_20185 (I466086,I2859,I346026,I346052,);
not I_20186 (I346060,I346052);
nand I_20187 (I346077,I466068,I466068);
and I_20188 (I346094,I346077,I466074);
DFFARX1 I_20189 (I346094,I2859,I346026,I346120,);
DFFARX1 I_20190 (I346120,I2859,I346026,I346015,);
DFFARX1 I_20191 (I466071,I2859,I346026,I346151,);
nand I_20192 (I346159,I346151,I466080);
not I_20193 (I346176,I346159);
DFFARX1 I_20194 (I346176,I2859,I346026,I346202,);
not I_20195 (I346210,I346202);
nor I_20196 (I346018,I346060,I346210);
DFFARX1 I_20197 (I466092,I2859,I346026,I346250,);
nor I_20198 (I346009,I346250,I346120);
nor I_20199 (I346000,I346250,I346176);
nand I_20200 (I346286,I466083,I466077);
and I_20201 (I346303,I346286,I466071);
DFFARX1 I_20202 (I346303,I2859,I346026,I346329,);
not I_20203 (I346337,I346329);
nand I_20204 (I346354,I346337,I346250);
nand I_20205 (I346003,I346337,I346159);
nor I_20206 (I346385,I466089,I466077);
and I_20207 (I346402,I346250,I346385);
nor I_20208 (I346419,I346337,I346402);
DFFARX1 I_20209 (I346419,I2859,I346026,I346012,);
nor I_20210 (I346450,I346052,I346385);
DFFARX1 I_20211 (I346450,I2859,I346026,I345997,);
nor I_20212 (I346481,I346329,I346385);
not I_20213 (I346498,I346481);
nand I_20214 (I346006,I346498,I346354);
not I_20215 (I346553,I2866);
DFFARX1 I_20216 (I301304,I2859,I346553,I346579,);
not I_20217 (I346587,I346579);
nand I_20218 (I346604,I301307,I301304);
and I_20219 (I346621,I346604,I301316);
DFFARX1 I_20220 (I346621,I2859,I346553,I346647,);
DFFARX1 I_20221 (I346647,I2859,I346553,I346542,);
DFFARX1 I_20222 (I301313,I2859,I346553,I346678,);
nand I_20223 (I346686,I346678,I301319);
not I_20224 (I346703,I346686);
DFFARX1 I_20225 (I346703,I2859,I346553,I346729,);
not I_20226 (I346737,I346729);
nor I_20227 (I346545,I346587,I346737);
DFFARX1 I_20228 (I301328,I2859,I346553,I346777,);
nor I_20229 (I346536,I346777,I346647);
nor I_20230 (I346527,I346777,I346703);
nand I_20231 (I346813,I301322,I301310);
and I_20232 (I346830,I346813,I301307);
DFFARX1 I_20233 (I346830,I2859,I346553,I346856,);
not I_20234 (I346864,I346856);
nand I_20235 (I346881,I346864,I346777);
nand I_20236 (I346530,I346864,I346686);
nor I_20237 (I346912,I301325,I301310);
and I_20238 (I346929,I346777,I346912);
nor I_20239 (I346946,I346864,I346929);
DFFARX1 I_20240 (I346946,I2859,I346553,I346539,);
nor I_20241 (I346977,I346579,I346912);
DFFARX1 I_20242 (I346977,I2859,I346553,I346524,);
nor I_20243 (I347008,I346856,I346912);
not I_20244 (I347025,I347008);
nand I_20245 (I346533,I347025,I346881);
not I_20246 (I347080,I2866);
DFFARX1 I_20247 (I543365,I2859,I347080,I347106,);
not I_20248 (I347114,I347106);
nand I_20249 (I347131,I543362,I543371);
and I_20250 (I347148,I347131,I543350);
DFFARX1 I_20251 (I347148,I2859,I347080,I347174,);
DFFARX1 I_20252 (I347174,I2859,I347080,I347069,);
DFFARX1 I_20253 (I543353,I2859,I347080,I347205,);
nand I_20254 (I347213,I347205,I543368);
not I_20255 (I347230,I347213);
DFFARX1 I_20256 (I347230,I2859,I347080,I347256,);
not I_20257 (I347264,I347256);
nor I_20258 (I347072,I347114,I347264);
DFFARX1 I_20259 (I543374,I2859,I347080,I347304,);
nor I_20260 (I347063,I347304,I347174);
nor I_20261 (I347054,I347304,I347230);
nand I_20262 (I347340,I543356,I543377);
and I_20263 (I347357,I347340,I543359);
DFFARX1 I_20264 (I347357,I2859,I347080,I347383,);
not I_20265 (I347391,I347383);
nand I_20266 (I347408,I347391,I347304);
nand I_20267 (I347057,I347391,I347213);
nor I_20268 (I347439,I543350,I543377);
and I_20269 (I347456,I347304,I347439);
nor I_20270 (I347473,I347391,I347456);
DFFARX1 I_20271 (I347473,I2859,I347080,I347066,);
nor I_20272 (I347504,I347106,I347439);
DFFARX1 I_20273 (I347504,I2859,I347080,I347051,);
nor I_20274 (I347535,I347383,I347439);
not I_20275 (I347552,I347535);
nand I_20276 (I347060,I347552,I347408);
not I_20277 (I347607,I2866);
DFFARX1 I_20278 (I475912,I2859,I347607,I347633,);
not I_20279 (I347641,I347633);
nand I_20280 (I347658,I475894,I475894);
and I_20281 (I347675,I347658,I475900);
DFFARX1 I_20282 (I347675,I2859,I347607,I347701,);
DFFARX1 I_20283 (I347701,I2859,I347607,I347596,);
DFFARX1 I_20284 (I475897,I2859,I347607,I347732,);
nand I_20285 (I347740,I347732,I475906);
not I_20286 (I347757,I347740);
DFFARX1 I_20287 (I347757,I2859,I347607,I347783,);
not I_20288 (I347791,I347783);
nor I_20289 (I347599,I347641,I347791);
DFFARX1 I_20290 (I475918,I2859,I347607,I347831,);
nor I_20291 (I347590,I347831,I347701);
nor I_20292 (I347581,I347831,I347757);
nand I_20293 (I347867,I475909,I475903);
and I_20294 (I347884,I347867,I475897);
DFFARX1 I_20295 (I347884,I2859,I347607,I347910,);
not I_20296 (I347918,I347910);
nand I_20297 (I347935,I347918,I347831);
nand I_20298 (I347584,I347918,I347740);
nor I_20299 (I347966,I475915,I475903);
and I_20300 (I347983,I347831,I347966);
nor I_20301 (I348000,I347918,I347983);
DFFARX1 I_20302 (I348000,I2859,I347607,I347593,);
nor I_20303 (I348031,I347633,I347966);
DFFARX1 I_20304 (I348031,I2859,I347607,I347578,);
nor I_20305 (I348062,I347910,I347966);
not I_20306 (I348079,I348062);
nand I_20307 (I347587,I348079,I347935);
not I_20308 (I348134,I2866);
DFFARX1 I_20309 (I229647,I2859,I348134,I348160,);
not I_20310 (I348168,I348160);
nand I_20311 (I348185,I229632,I229653);
and I_20312 (I348202,I348185,I229641);
DFFARX1 I_20313 (I348202,I2859,I348134,I348228,);
DFFARX1 I_20314 (I348228,I2859,I348134,I348123,);
DFFARX1 I_20315 (I229635,I2859,I348134,I348259,);
nand I_20316 (I348267,I348259,I229644);
not I_20317 (I348284,I348267);
DFFARX1 I_20318 (I348284,I2859,I348134,I348310,);
not I_20319 (I348318,I348310);
nor I_20320 (I348126,I348168,I348318);
DFFARX1 I_20321 (I229650,I2859,I348134,I348358,);
nor I_20322 (I348117,I348358,I348228);
nor I_20323 (I348108,I348358,I348284);
nand I_20324 (I348394,I229632,I229635);
and I_20325 (I348411,I348394,I229656);
DFFARX1 I_20326 (I348411,I2859,I348134,I348437,);
not I_20327 (I348445,I348437);
nand I_20328 (I348462,I348445,I348358);
nand I_20329 (I348111,I348445,I348267);
nor I_20330 (I348493,I229638,I229635);
and I_20331 (I348510,I348358,I348493);
nor I_20332 (I348527,I348445,I348510);
DFFARX1 I_20333 (I348527,I2859,I348134,I348120,);
nor I_20334 (I348558,I348160,I348493);
DFFARX1 I_20335 (I348558,I2859,I348134,I348105,);
nor I_20336 (I348589,I348437,I348493);
not I_20337 (I348606,I348589);
nand I_20338 (I348114,I348606,I348462);
not I_20339 (I348661,I2866);
DFFARX1 I_20340 (I460884,I2859,I348661,I348687,);
not I_20341 (I348695,I348687);
nand I_20342 (I348712,I460866,I460866);
and I_20343 (I348729,I348712,I460872);
DFFARX1 I_20344 (I348729,I2859,I348661,I348755,);
DFFARX1 I_20345 (I348755,I2859,I348661,I348650,);
DFFARX1 I_20346 (I460869,I2859,I348661,I348786,);
nand I_20347 (I348794,I348786,I460878);
not I_20348 (I348811,I348794);
DFFARX1 I_20349 (I348811,I2859,I348661,I348837,);
not I_20350 (I348845,I348837);
nor I_20351 (I348653,I348695,I348845);
DFFARX1 I_20352 (I460890,I2859,I348661,I348885,);
nor I_20353 (I348644,I348885,I348755);
nor I_20354 (I348635,I348885,I348811);
nand I_20355 (I348921,I460881,I460875);
and I_20356 (I348938,I348921,I460869);
DFFARX1 I_20357 (I348938,I2859,I348661,I348964,);
not I_20358 (I348972,I348964);
nand I_20359 (I348989,I348972,I348885);
nand I_20360 (I348638,I348972,I348794);
nor I_20361 (I349020,I460887,I460875);
and I_20362 (I349037,I348885,I349020);
nor I_20363 (I349054,I348972,I349037);
DFFARX1 I_20364 (I349054,I2859,I348661,I348647,);
nor I_20365 (I349085,I348687,I349020);
DFFARX1 I_20366 (I349085,I2859,I348661,I348632,);
nor I_20367 (I349116,I348964,I349020);
not I_20368 (I349133,I349116);
nand I_20369 (I348641,I349133,I348989);
not I_20370 (I349188,I2866);
DFFARX1 I_20371 (I470132,I2859,I349188,I349214,);
not I_20372 (I349222,I349214);
nand I_20373 (I349239,I470114,I470114);
and I_20374 (I349256,I349239,I470120);
DFFARX1 I_20375 (I349256,I2859,I349188,I349282,);
DFFARX1 I_20376 (I349282,I2859,I349188,I349177,);
DFFARX1 I_20377 (I470117,I2859,I349188,I349313,);
nand I_20378 (I349321,I349313,I470126);
not I_20379 (I349338,I349321);
DFFARX1 I_20380 (I349338,I2859,I349188,I349364,);
not I_20381 (I349372,I349364);
nor I_20382 (I349180,I349222,I349372);
DFFARX1 I_20383 (I470138,I2859,I349188,I349412,);
nor I_20384 (I349171,I349412,I349282);
nor I_20385 (I349162,I349412,I349338);
nand I_20386 (I349448,I470129,I470123);
and I_20387 (I349465,I349448,I470117);
DFFARX1 I_20388 (I349465,I2859,I349188,I349491,);
not I_20389 (I349499,I349491);
nand I_20390 (I349516,I349499,I349412);
nand I_20391 (I349165,I349499,I349321);
nor I_20392 (I349547,I470135,I470123);
and I_20393 (I349564,I349412,I349547);
nor I_20394 (I349581,I349499,I349564);
DFFARX1 I_20395 (I349581,I2859,I349188,I349174,);
nor I_20396 (I349612,I349214,I349547);
DFFARX1 I_20397 (I349612,I2859,I349188,I349159,);
nor I_20398 (I349643,I349491,I349547);
not I_20399 (I349660,I349643);
nand I_20400 (I349168,I349660,I349516);
not I_20401 (I349715,I2866);
DFFARX1 I_20402 (I76893,I2859,I349715,I349741,);
not I_20403 (I349749,I349741);
nand I_20404 (I349766,I76890,I76908);
and I_20405 (I349783,I349766,I76899);
DFFARX1 I_20406 (I349783,I2859,I349715,I349809,);
DFFARX1 I_20407 (I349809,I2859,I349715,I349704,);
DFFARX1 I_20408 (I76905,I2859,I349715,I349840,);
nand I_20409 (I349848,I349840,I76902);
not I_20410 (I349865,I349848);
DFFARX1 I_20411 (I349865,I2859,I349715,I349891,);
not I_20412 (I349899,I349891);
nor I_20413 (I349707,I349749,I349899);
DFFARX1 I_20414 (I76896,I2859,I349715,I349939,);
nor I_20415 (I349698,I349939,I349809);
nor I_20416 (I349689,I349939,I349865);
nand I_20417 (I349975,I76887,I76911);
and I_20418 (I349992,I349975,I76890);
DFFARX1 I_20419 (I349992,I2859,I349715,I350018,);
not I_20420 (I350026,I350018);
nand I_20421 (I350043,I350026,I349939);
nand I_20422 (I349692,I350026,I349848);
nor I_20423 (I350074,I76887,I76911);
and I_20424 (I350091,I349939,I350074);
nor I_20425 (I350108,I350026,I350091);
DFFARX1 I_20426 (I350108,I2859,I349715,I349701,);
nor I_20427 (I350139,I349741,I350074);
DFFARX1 I_20428 (I350139,I2859,I349715,I349686,);
nor I_20429 (I350170,I350018,I350074);
not I_20430 (I350187,I350170);
nand I_20431 (I349695,I350187,I350043);
not I_20432 (I350242,I2866);
DFFARX1 I_20433 (I380544,I2859,I350242,I350268,);
not I_20434 (I350276,I350268);
nand I_20435 (I350293,I380559,I380541);
and I_20436 (I350310,I350293,I380541);
DFFARX1 I_20437 (I350310,I2859,I350242,I350336,);
DFFARX1 I_20438 (I350336,I2859,I350242,I350231,);
DFFARX1 I_20439 (I380550,I2859,I350242,I350367,);
nand I_20440 (I350375,I350367,I380568);
not I_20441 (I350392,I350375);
DFFARX1 I_20442 (I350392,I2859,I350242,I350418,);
not I_20443 (I350426,I350418);
nor I_20444 (I350234,I350276,I350426);
DFFARX1 I_20445 (I380565,I2859,I350242,I350466,);
nor I_20446 (I350225,I350466,I350336);
nor I_20447 (I350216,I350466,I350392);
nand I_20448 (I350502,I380562,I380553);
and I_20449 (I350519,I350502,I380547);
DFFARX1 I_20450 (I350519,I2859,I350242,I350545,);
not I_20451 (I350553,I350545);
nand I_20452 (I350570,I350553,I350466);
nand I_20453 (I350219,I350553,I350375);
nor I_20454 (I350601,I380556,I380553);
and I_20455 (I350618,I350466,I350601);
nor I_20456 (I350635,I350553,I350618);
DFFARX1 I_20457 (I350635,I2859,I350242,I350228,);
nor I_20458 (I350666,I350268,I350601);
DFFARX1 I_20459 (I350666,I2859,I350242,I350213,);
nor I_20460 (I350697,I350545,I350601);
not I_20461 (I350714,I350697);
nand I_20462 (I350222,I350714,I350570);
not I_20463 (I350769,I2866);
DFFARX1 I_20464 (I157255,I2859,I350769,I350795,);
not I_20465 (I350803,I350795);
nand I_20466 (I350820,I157246,I157246);
and I_20467 (I350837,I350820,I157264);
DFFARX1 I_20468 (I350837,I2859,I350769,I350863,);
DFFARX1 I_20469 (I350863,I2859,I350769,I350758,);
DFFARX1 I_20470 (I157267,I2859,I350769,I350894,);
nand I_20471 (I350902,I350894,I157249);
not I_20472 (I350919,I350902);
DFFARX1 I_20473 (I350919,I2859,I350769,I350945,);
not I_20474 (I350953,I350945);
nor I_20475 (I350761,I350803,I350953);
DFFARX1 I_20476 (I157261,I2859,I350769,I350993,);
nor I_20477 (I350752,I350993,I350863);
nor I_20478 (I350743,I350993,I350919);
nand I_20479 (I351029,I157273,I157252);
and I_20480 (I351046,I351029,I157258);
DFFARX1 I_20481 (I351046,I2859,I350769,I351072,);
not I_20482 (I351080,I351072);
nand I_20483 (I351097,I351080,I350993);
nand I_20484 (I350746,I351080,I350902);
nor I_20485 (I351128,I157270,I157252);
and I_20486 (I351145,I350993,I351128);
nor I_20487 (I351162,I351080,I351145);
DFFARX1 I_20488 (I351162,I2859,I350769,I350755,);
nor I_20489 (I351193,I350795,I351128);
DFFARX1 I_20490 (I351193,I2859,I350769,I350740,);
nor I_20491 (I351224,I351072,I351128);
not I_20492 (I351241,I351224);
nand I_20493 (I350749,I351241,I351097);
not I_20494 (I351296,I2866);
DFFARX1 I_20495 (I121946,I2859,I351296,I351322,);
not I_20496 (I351330,I351322);
nand I_20497 (I351347,I121937,I121937);
and I_20498 (I351364,I351347,I121955);
DFFARX1 I_20499 (I351364,I2859,I351296,I351390,);
DFFARX1 I_20500 (I351390,I2859,I351296,I351285,);
DFFARX1 I_20501 (I121958,I2859,I351296,I351421,);
nand I_20502 (I351429,I351421,I121940);
not I_20503 (I351446,I351429);
DFFARX1 I_20504 (I351446,I2859,I351296,I351472,);
not I_20505 (I351480,I351472);
nor I_20506 (I351288,I351330,I351480);
DFFARX1 I_20507 (I121952,I2859,I351296,I351520,);
nor I_20508 (I351279,I351520,I351390);
nor I_20509 (I351270,I351520,I351446);
nand I_20510 (I351556,I121964,I121943);
and I_20511 (I351573,I351556,I121949);
DFFARX1 I_20512 (I351573,I2859,I351296,I351599,);
not I_20513 (I351607,I351599);
nand I_20514 (I351624,I351607,I351520);
nand I_20515 (I351273,I351607,I351429);
nor I_20516 (I351655,I121961,I121943);
and I_20517 (I351672,I351520,I351655);
nor I_20518 (I351689,I351607,I351672);
DFFARX1 I_20519 (I351689,I2859,I351296,I351282,);
nor I_20520 (I351720,I351322,I351655);
DFFARX1 I_20521 (I351720,I2859,I351296,I351267,);
nor I_20522 (I351751,I351599,I351655);
not I_20523 (I351768,I351751);
nand I_20524 (I351276,I351768,I351624);
not I_20525 (I351823,I2866);
DFFARX1 I_20526 (I43812,I2859,I351823,I351849,);
not I_20527 (I351857,I351849);
nand I_20528 (I351874,I43788,I43797);
and I_20529 (I351891,I351874,I43791);
DFFARX1 I_20530 (I351891,I2859,I351823,I351917,);
DFFARX1 I_20531 (I351917,I2859,I351823,I351812,);
DFFARX1 I_20532 (I43809,I2859,I351823,I351948,);
nand I_20533 (I351956,I351948,I43800);
not I_20534 (I351973,I351956);
DFFARX1 I_20535 (I351973,I2859,I351823,I351999,);
not I_20536 (I352007,I351999);
nor I_20537 (I351815,I351857,I352007);
DFFARX1 I_20538 (I43794,I2859,I351823,I352047,);
nor I_20539 (I351806,I352047,I351917);
nor I_20540 (I351797,I352047,I351973);
nand I_20541 (I352083,I43806,I43803);
and I_20542 (I352100,I352083,I43791);
DFFARX1 I_20543 (I352100,I2859,I351823,I352126,);
not I_20544 (I352134,I352126);
nand I_20545 (I352151,I352134,I352047);
nand I_20546 (I351800,I352134,I351956);
nor I_20547 (I352182,I43788,I43803);
and I_20548 (I352199,I352047,I352182);
nor I_20549 (I352216,I352134,I352199);
DFFARX1 I_20550 (I352216,I2859,I351823,I351809,);
nor I_20551 (I352247,I351849,I352182);
DFFARX1 I_20552 (I352247,I2859,I351823,I351794,);
nor I_20553 (I352278,I352126,I352182);
not I_20554 (I352295,I352278);
nand I_20555 (I351803,I352295,I352151);
not I_20556 (I352350,I2866);
DFFARX1 I_20557 (I193054,I2859,I352350,I352376,);
not I_20558 (I352384,I352376);
nand I_20559 (I352401,I193051,I193060);
and I_20560 (I352418,I352401,I193069);
DFFARX1 I_20561 (I352418,I2859,I352350,I352444,);
DFFARX1 I_20562 (I352444,I2859,I352350,I352339,);
DFFARX1 I_20563 (I193072,I2859,I352350,I352475,);
nand I_20564 (I352483,I352475,I193075);
not I_20565 (I352500,I352483);
DFFARX1 I_20566 (I352500,I2859,I352350,I352526,);
not I_20567 (I352534,I352526);
nor I_20568 (I352342,I352384,I352534);
DFFARX1 I_20569 (I193048,I2859,I352350,I352574,);
nor I_20570 (I352333,I352574,I352444);
nor I_20571 (I352324,I352574,I352500);
nand I_20572 (I352610,I193063,I193066);
and I_20573 (I352627,I352610,I193057);
DFFARX1 I_20574 (I352627,I2859,I352350,I352653,);
not I_20575 (I352661,I352653);
nand I_20576 (I352678,I352661,I352574);
nand I_20577 (I352327,I352661,I352483);
nor I_20578 (I352709,I193048,I193066);
and I_20579 (I352726,I352574,I352709);
nor I_20580 (I352743,I352661,I352726);
DFFARX1 I_20581 (I352743,I2859,I352350,I352336,);
nor I_20582 (I352774,I352376,I352709);
DFFARX1 I_20583 (I352774,I2859,I352350,I352321,);
nor I_20584 (I352805,I352653,I352709);
not I_20585 (I352822,I352805);
nand I_20586 (I352330,I352822,I352678);
not I_20587 (I352877,I2866);
DFFARX1 I_20588 (I538010,I2859,I352877,I352903,);
not I_20589 (I352911,I352903);
nand I_20590 (I352928,I538007,I538016);
and I_20591 (I352945,I352928,I537995);
DFFARX1 I_20592 (I352945,I2859,I352877,I352971,);
DFFARX1 I_20593 (I352971,I2859,I352877,I352866,);
DFFARX1 I_20594 (I537998,I2859,I352877,I353002,);
nand I_20595 (I353010,I353002,I538013);
not I_20596 (I353027,I353010);
DFFARX1 I_20597 (I353027,I2859,I352877,I353053,);
not I_20598 (I353061,I353053);
nor I_20599 (I352869,I352911,I353061);
DFFARX1 I_20600 (I538019,I2859,I352877,I353101,);
nor I_20601 (I352860,I353101,I352971);
nor I_20602 (I352851,I353101,I353027);
nand I_20603 (I353137,I538001,I538022);
and I_20604 (I353154,I353137,I538004);
DFFARX1 I_20605 (I353154,I2859,I352877,I353180,);
not I_20606 (I353188,I353180);
nand I_20607 (I353205,I353188,I353101);
nand I_20608 (I352854,I353188,I353010);
nor I_20609 (I353236,I537995,I538022);
and I_20610 (I353253,I353101,I353236);
nor I_20611 (I353270,I353188,I353253);
DFFARX1 I_20612 (I353270,I2859,I352877,I352863,);
nor I_20613 (I353301,I352903,I353236);
DFFARX1 I_20614 (I353301,I2859,I352877,I352848,);
nor I_20615 (I353332,I353180,I353236);
not I_20616 (I353349,I353332);
nand I_20617 (I352857,I353349,I353205);
not I_20618 (I353404,I2866);
DFFARX1 I_20619 (I137756,I2859,I353404,I353430,);
not I_20620 (I353438,I353430);
nand I_20621 (I353455,I137747,I137747);
and I_20622 (I353472,I353455,I137765);
DFFARX1 I_20623 (I353472,I2859,I353404,I353498,);
DFFARX1 I_20624 (I353498,I2859,I353404,I353393,);
DFFARX1 I_20625 (I137768,I2859,I353404,I353529,);
nand I_20626 (I353537,I353529,I137750);
not I_20627 (I353554,I353537);
DFFARX1 I_20628 (I353554,I2859,I353404,I353580,);
not I_20629 (I353588,I353580);
nor I_20630 (I353396,I353438,I353588);
DFFARX1 I_20631 (I137762,I2859,I353404,I353628,);
nor I_20632 (I353387,I353628,I353498);
nor I_20633 (I353378,I353628,I353554);
nand I_20634 (I353664,I137774,I137753);
and I_20635 (I353681,I353664,I137759);
DFFARX1 I_20636 (I353681,I2859,I353404,I353707,);
not I_20637 (I353715,I353707);
nand I_20638 (I353732,I353715,I353628);
nand I_20639 (I353381,I353715,I353537);
nor I_20640 (I353763,I137771,I137753);
and I_20641 (I353780,I353628,I353763);
nor I_20642 (I353797,I353715,I353780);
DFFARX1 I_20643 (I353797,I2859,I353404,I353390,);
nor I_20644 (I353828,I353430,I353763);
DFFARX1 I_20645 (I353828,I2859,I353404,I353375,);
nor I_20646 (I353859,I353707,I353763);
not I_20647 (I353876,I353859);
nand I_20648 (I353384,I353876,I353732);
not I_20649 (I353931,I2866);
DFFARX1 I_20650 (I252189,I2859,I353931,I353957,);
not I_20651 (I353965,I353957);
nand I_20652 (I353982,I252174,I252195);
and I_20653 (I353999,I353982,I252183);
DFFARX1 I_20654 (I353999,I2859,I353931,I354025,);
DFFARX1 I_20655 (I354025,I2859,I353931,I353920,);
DFFARX1 I_20656 (I252177,I2859,I353931,I354056,);
nand I_20657 (I354064,I354056,I252186);
not I_20658 (I354081,I354064);
DFFARX1 I_20659 (I354081,I2859,I353931,I354107,);
not I_20660 (I354115,I354107);
nor I_20661 (I353923,I353965,I354115);
DFFARX1 I_20662 (I252192,I2859,I353931,I354155,);
nor I_20663 (I353914,I354155,I354025);
nor I_20664 (I353905,I354155,I354081);
nand I_20665 (I354191,I252174,I252177);
and I_20666 (I354208,I354191,I252198);
DFFARX1 I_20667 (I354208,I2859,I353931,I354234,);
not I_20668 (I354242,I354234);
nand I_20669 (I354259,I354242,I354155);
nand I_20670 (I353908,I354242,I354064);
nor I_20671 (I354290,I252180,I252177);
and I_20672 (I354307,I354155,I354290);
nor I_20673 (I354324,I354242,I354307);
DFFARX1 I_20674 (I354324,I2859,I353931,I353917,);
nor I_20675 (I354355,I353957,I354290);
DFFARX1 I_20676 (I354355,I2859,I353931,I353902,);
nor I_20677 (I354386,I354234,I354290);
not I_20678 (I354403,I354386);
nand I_20679 (I353911,I354403,I354259);
not I_20680 (I354458,I2866);
DFFARX1 I_20681 (I228491,I2859,I354458,I354484,);
not I_20682 (I354492,I354484);
nand I_20683 (I354509,I228476,I228497);
and I_20684 (I354526,I354509,I228485);
DFFARX1 I_20685 (I354526,I2859,I354458,I354552,);
DFFARX1 I_20686 (I354552,I2859,I354458,I354447,);
DFFARX1 I_20687 (I228479,I2859,I354458,I354583,);
nand I_20688 (I354591,I354583,I228488);
not I_20689 (I354608,I354591);
DFFARX1 I_20690 (I354608,I2859,I354458,I354634,);
not I_20691 (I354642,I354634);
nor I_20692 (I354450,I354492,I354642);
DFFARX1 I_20693 (I228494,I2859,I354458,I354682,);
nor I_20694 (I354441,I354682,I354552);
nor I_20695 (I354432,I354682,I354608);
nand I_20696 (I354718,I228476,I228479);
and I_20697 (I354735,I354718,I228500);
DFFARX1 I_20698 (I354735,I2859,I354458,I354761,);
not I_20699 (I354769,I354761);
nand I_20700 (I354786,I354769,I354682);
nand I_20701 (I354435,I354769,I354591);
nor I_20702 (I354817,I228482,I228479);
and I_20703 (I354834,I354682,I354817);
nor I_20704 (I354851,I354769,I354834);
DFFARX1 I_20705 (I354851,I2859,I354458,I354444,);
nor I_20706 (I354882,I354484,I354817);
DFFARX1 I_20707 (I354882,I2859,I354458,I354429,);
nor I_20708 (I354913,I354761,I354817);
not I_20709 (I354930,I354913);
nand I_20710 (I354438,I354930,I354786);
not I_20711 (I354985,I2866);
DFFARX1 I_20712 (I273560,I2859,I354985,I355011,);
not I_20713 (I355019,I355011);
nand I_20714 (I355036,I273563,I273560);
and I_20715 (I355053,I355036,I273572);
DFFARX1 I_20716 (I355053,I2859,I354985,I355079,);
DFFARX1 I_20717 (I355079,I2859,I354985,I354974,);
DFFARX1 I_20718 (I273569,I2859,I354985,I355110,);
nand I_20719 (I355118,I355110,I273575);
not I_20720 (I355135,I355118);
DFFARX1 I_20721 (I355135,I2859,I354985,I355161,);
not I_20722 (I355169,I355161);
nor I_20723 (I354977,I355019,I355169);
DFFARX1 I_20724 (I273584,I2859,I354985,I355209,);
nor I_20725 (I354968,I355209,I355079);
nor I_20726 (I354959,I355209,I355135);
nand I_20727 (I355245,I273578,I273566);
and I_20728 (I355262,I355245,I273563);
DFFARX1 I_20729 (I355262,I2859,I354985,I355288,);
not I_20730 (I355296,I355288);
nand I_20731 (I355313,I355296,I355209);
nand I_20732 (I354962,I355296,I355118);
nor I_20733 (I355344,I273581,I273566);
and I_20734 (I355361,I355209,I355344);
nor I_20735 (I355378,I355296,I355361);
DFFARX1 I_20736 (I355378,I2859,I354985,I354971,);
nor I_20737 (I355409,I355011,I355344);
DFFARX1 I_20738 (I355409,I2859,I354985,I354956,);
nor I_20739 (I355440,I355288,I355344);
not I_20740 (I355457,I355440);
nand I_20741 (I354965,I355457,I355313);
not I_20742 (I355512,I2866);
DFFARX1 I_20743 (I164766,I2859,I355512,I355538,);
not I_20744 (I355546,I355538);
nand I_20745 (I355563,I164763,I164772);
and I_20746 (I355580,I355563,I164781);
DFFARX1 I_20747 (I355580,I2859,I355512,I355606,);
DFFARX1 I_20748 (I355606,I2859,I355512,I355501,);
DFFARX1 I_20749 (I164784,I2859,I355512,I355637,);
nand I_20750 (I355645,I355637,I164787);
not I_20751 (I355662,I355645);
DFFARX1 I_20752 (I355662,I2859,I355512,I355688,);
not I_20753 (I355696,I355688);
nor I_20754 (I355504,I355546,I355696);
DFFARX1 I_20755 (I164760,I2859,I355512,I355736,);
nor I_20756 (I355495,I355736,I355606);
nor I_20757 (I355486,I355736,I355662);
nand I_20758 (I355772,I164775,I164778);
and I_20759 (I355789,I355772,I164769);
DFFARX1 I_20760 (I355789,I2859,I355512,I355815,);
not I_20761 (I355823,I355815);
nand I_20762 (I355840,I355823,I355736);
nand I_20763 (I355489,I355823,I355645);
nor I_20764 (I355871,I164760,I164778);
and I_20765 (I355888,I355736,I355871);
nor I_20766 (I355905,I355823,I355888);
DFFARX1 I_20767 (I355905,I2859,I355512,I355498,);
nor I_20768 (I355936,I355538,I355871);
DFFARX1 I_20769 (I355936,I2859,I355512,I355483,);
nor I_20770 (I355967,I355815,I355871);
not I_20771 (I355984,I355967);
nand I_20772 (I355492,I355984,I355840);
not I_20773 (I356039,I2866);
DFFARX1 I_20774 (I316332,I2859,I356039,I356065,);
not I_20775 (I356073,I356065);
nand I_20776 (I356090,I316335,I316332);
and I_20777 (I356107,I356090,I316344);
DFFARX1 I_20778 (I356107,I2859,I356039,I356133,);
DFFARX1 I_20779 (I356133,I2859,I356039,I356028,);
DFFARX1 I_20780 (I316341,I2859,I356039,I356164,);
nand I_20781 (I356172,I356164,I316347);
not I_20782 (I356189,I356172);
DFFARX1 I_20783 (I356189,I2859,I356039,I356215,);
not I_20784 (I356223,I356215);
nor I_20785 (I356031,I356073,I356223);
DFFARX1 I_20786 (I316356,I2859,I356039,I356263,);
nor I_20787 (I356022,I356263,I356133);
nor I_20788 (I356013,I356263,I356189);
nand I_20789 (I356299,I316350,I316338);
and I_20790 (I356316,I356299,I316335);
DFFARX1 I_20791 (I356316,I2859,I356039,I356342,);
not I_20792 (I356350,I356342);
nand I_20793 (I356367,I356350,I356263);
nand I_20794 (I356016,I356350,I356172);
nor I_20795 (I356398,I316353,I316338);
and I_20796 (I356415,I356263,I356398);
nor I_20797 (I356432,I356350,I356415);
DFFARX1 I_20798 (I356432,I2859,I356039,I356025,);
nor I_20799 (I356463,I356065,I356398);
DFFARX1 I_20800 (I356463,I2859,I356039,I356010,);
nor I_20801 (I356494,I356342,I356398);
not I_20802 (I356511,I356494);
nand I_20803 (I356019,I356511,I356367);
not I_20804 (I356566,I2866);
DFFARX1 I_20805 (I544555,I2859,I356566,I356592,);
not I_20806 (I356600,I356592);
nand I_20807 (I356617,I544552,I544561);
and I_20808 (I356634,I356617,I544540);
DFFARX1 I_20809 (I356634,I2859,I356566,I356660,);
DFFARX1 I_20810 (I356660,I2859,I356566,I356555,);
DFFARX1 I_20811 (I544543,I2859,I356566,I356691,);
nand I_20812 (I356699,I356691,I544558);
not I_20813 (I356716,I356699);
DFFARX1 I_20814 (I356716,I2859,I356566,I356742,);
not I_20815 (I356750,I356742);
nor I_20816 (I356558,I356600,I356750);
DFFARX1 I_20817 (I544564,I2859,I356566,I356790,);
nor I_20818 (I356549,I356790,I356660);
nor I_20819 (I356540,I356790,I356716);
nand I_20820 (I356826,I544546,I544567);
and I_20821 (I356843,I356826,I544549);
DFFARX1 I_20822 (I356843,I2859,I356566,I356869,);
not I_20823 (I356877,I356869);
nand I_20824 (I356894,I356877,I356790);
nand I_20825 (I356543,I356877,I356699);
nor I_20826 (I356925,I544540,I544567);
and I_20827 (I356942,I356790,I356925);
nor I_20828 (I356959,I356877,I356942);
DFFARX1 I_20829 (I356959,I2859,I356566,I356552,);
nor I_20830 (I356990,I356592,I356925);
DFFARX1 I_20831 (I356990,I2859,I356566,I356537,);
nor I_20832 (I357021,I356869,I356925);
not I_20833 (I357038,I357021);
nand I_20834 (I356546,I357038,I356894);
not I_20835 (I357093,I2866);
DFFARX1 I_20836 (I286854,I2859,I357093,I357119,);
not I_20837 (I357127,I357119);
nand I_20838 (I357144,I286857,I286854);
and I_20839 (I357161,I357144,I286866);
DFFARX1 I_20840 (I357161,I2859,I357093,I357187,);
DFFARX1 I_20841 (I357187,I2859,I357093,I357082,);
DFFARX1 I_20842 (I286863,I2859,I357093,I357218,);
nand I_20843 (I357226,I357218,I286869);
not I_20844 (I357243,I357226);
DFFARX1 I_20845 (I357243,I2859,I357093,I357269,);
not I_20846 (I357277,I357269);
nor I_20847 (I357085,I357127,I357277);
DFFARX1 I_20848 (I286878,I2859,I357093,I357317,);
nor I_20849 (I357076,I357317,I357187);
nor I_20850 (I357067,I357317,I357243);
nand I_20851 (I357353,I286872,I286860);
and I_20852 (I357370,I357353,I286857);
DFFARX1 I_20853 (I357370,I2859,I357093,I357396,);
not I_20854 (I357404,I357396);
nand I_20855 (I357421,I357404,I357317);
nand I_20856 (I357070,I357404,I357226);
nor I_20857 (I357452,I286875,I286860);
and I_20858 (I357469,I357317,I357452);
nor I_20859 (I357486,I357404,I357469);
DFFARX1 I_20860 (I357486,I2859,I357093,I357079,);
nor I_20861 (I357517,I357119,I357452);
DFFARX1 I_20862 (I357517,I2859,I357093,I357064,);
nor I_20863 (I357548,I357396,I357452);
not I_20864 (I357565,I357548);
nand I_20865 (I357073,I357565,I357421);
not I_20866 (I357620,I2866);
DFFARX1 I_20867 (I122473,I2859,I357620,I357646,);
not I_20868 (I357654,I357646);
nand I_20869 (I357671,I122464,I122464);
and I_20870 (I357688,I357671,I122482);
DFFARX1 I_20871 (I357688,I2859,I357620,I357714,);
DFFARX1 I_20872 (I357714,I2859,I357620,I357609,);
DFFARX1 I_20873 (I122485,I2859,I357620,I357745,);
nand I_20874 (I357753,I357745,I122467);
not I_20875 (I357770,I357753);
DFFARX1 I_20876 (I357770,I2859,I357620,I357796,);
not I_20877 (I357804,I357796);
nor I_20878 (I357612,I357654,I357804);
DFFARX1 I_20879 (I122479,I2859,I357620,I357844,);
nor I_20880 (I357603,I357844,I357714);
nor I_20881 (I357594,I357844,I357770);
nand I_20882 (I357880,I122491,I122470);
and I_20883 (I357897,I357880,I122476);
DFFARX1 I_20884 (I357897,I2859,I357620,I357923,);
not I_20885 (I357931,I357923);
nand I_20886 (I357948,I357931,I357844);
nand I_20887 (I357597,I357931,I357753);
nor I_20888 (I357979,I122488,I122470);
and I_20889 (I357996,I357844,I357979);
nor I_20890 (I358013,I357931,I357996);
DFFARX1 I_20891 (I358013,I2859,I357620,I357606,);
nor I_20892 (I358044,I357646,I357979);
DFFARX1 I_20893 (I358044,I2859,I357620,I357591,);
nor I_20894 (I358075,I357923,I357979);
not I_20895 (I358092,I358075);
nand I_20896 (I357600,I358092,I357948);
not I_20897 (I358147,I2866);
DFFARX1 I_20898 (I127216,I2859,I358147,I358173,);
not I_20899 (I358181,I358173);
nand I_20900 (I358198,I127207,I127207);
and I_20901 (I358215,I358198,I127225);
DFFARX1 I_20902 (I358215,I2859,I358147,I358241,);
DFFARX1 I_20903 (I358241,I2859,I358147,I358136,);
DFFARX1 I_20904 (I127228,I2859,I358147,I358272,);
nand I_20905 (I358280,I358272,I127210);
not I_20906 (I358297,I358280);
DFFARX1 I_20907 (I358297,I2859,I358147,I358323,);
not I_20908 (I358331,I358323);
nor I_20909 (I358139,I358181,I358331);
DFFARX1 I_20910 (I127222,I2859,I358147,I358371,);
nor I_20911 (I358130,I358371,I358241);
nor I_20912 (I358121,I358371,I358297);
nand I_20913 (I358407,I127234,I127213);
and I_20914 (I358424,I358407,I127219);
DFFARX1 I_20915 (I358424,I2859,I358147,I358450,);
not I_20916 (I358458,I358450);
nand I_20917 (I358475,I358458,I358371);
nand I_20918 (I358124,I358458,I358280);
nor I_20919 (I358506,I127231,I127213);
and I_20920 (I358523,I358371,I358506);
nor I_20921 (I358540,I358458,I358523);
DFFARX1 I_20922 (I358540,I2859,I358147,I358133,);
nor I_20923 (I358571,I358173,I358506);
DFFARX1 I_20924 (I358571,I2859,I358147,I358118,);
nor I_20925 (I358602,I358450,I358506);
not I_20926 (I358619,I358602);
nand I_20927 (I358127,I358619,I358475);
not I_20928 (I358674,I2866);
DFFARX1 I_20929 (I474178,I2859,I358674,I358700,);
not I_20930 (I358708,I358700);
nand I_20931 (I358725,I474160,I474160);
and I_20932 (I358742,I358725,I474166);
DFFARX1 I_20933 (I358742,I2859,I358674,I358768,);
DFFARX1 I_20934 (I358768,I2859,I358674,I358663,);
DFFARX1 I_20935 (I474163,I2859,I358674,I358799,);
nand I_20936 (I358807,I358799,I474172);
not I_20937 (I358824,I358807);
DFFARX1 I_20938 (I358824,I2859,I358674,I358850,);
not I_20939 (I358858,I358850);
nor I_20940 (I358666,I358708,I358858);
DFFARX1 I_20941 (I474184,I2859,I358674,I358898,);
nor I_20942 (I358657,I358898,I358768);
nor I_20943 (I358648,I358898,I358824);
nand I_20944 (I358934,I474175,I474169);
and I_20945 (I358951,I358934,I474163);
DFFARX1 I_20946 (I358951,I2859,I358674,I358977,);
not I_20947 (I358985,I358977);
nand I_20948 (I359002,I358985,I358898);
nand I_20949 (I358651,I358985,I358807);
nor I_20950 (I359033,I474181,I474169);
and I_20951 (I359050,I358898,I359033);
nor I_20952 (I359067,I358985,I359050);
DFFARX1 I_20953 (I359067,I2859,I358674,I358660,);
nor I_20954 (I359098,I358700,I359033);
DFFARX1 I_20955 (I359098,I2859,I358674,I358645,);
nor I_20956 (I359129,I358977,I359033);
not I_20957 (I359146,I359129);
nand I_20958 (I358654,I359146,I359002);
not I_20959 (I359201,I2866);
DFFARX1 I_20960 (I457416,I2859,I359201,I359227,);
not I_20961 (I359235,I359227);
nand I_20962 (I359252,I457398,I457398);
and I_20963 (I359269,I359252,I457404);
DFFARX1 I_20964 (I359269,I2859,I359201,I359295,);
DFFARX1 I_20965 (I359295,I2859,I359201,I359190,);
DFFARX1 I_20966 (I457401,I2859,I359201,I359326,);
nand I_20967 (I359334,I359326,I457410);
not I_20968 (I359351,I359334);
DFFARX1 I_20969 (I359351,I2859,I359201,I359377,);
not I_20970 (I359385,I359377);
nor I_20971 (I359193,I359235,I359385);
DFFARX1 I_20972 (I457422,I2859,I359201,I359425,);
nor I_20973 (I359184,I359425,I359295);
nor I_20974 (I359175,I359425,I359351);
nand I_20975 (I359461,I457413,I457407);
and I_20976 (I359478,I359461,I457401);
DFFARX1 I_20977 (I359478,I2859,I359201,I359504,);
not I_20978 (I359512,I359504);
nand I_20979 (I359529,I359512,I359425);
nand I_20980 (I359178,I359512,I359334);
nor I_20981 (I359560,I457419,I457407);
and I_20982 (I359577,I359425,I359560);
nor I_20983 (I359594,I359512,I359577);
DFFARX1 I_20984 (I359594,I2859,I359201,I359187,);
nor I_20985 (I359625,I359227,I359560);
DFFARX1 I_20986 (I359625,I2859,I359201,I359172,);
nor I_20987 (I359656,I359504,I359560);
not I_20988 (I359673,I359656);
nand I_20989 (I359181,I359673,I359529);
not I_20990 (I359728,I2866);
DFFARX1 I_20991 (I100098,I2859,I359728,I359754,);
not I_20992 (I359762,I359754);
nand I_20993 (I359779,I100095,I100113);
and I_20994 (I359796,I359779,I100104);
DFFARX1 I_20995 (I359796,I2859,I359728,I359822,);
DFFARX1 I_20996 (I359822,I2859,I359728,I359717,);
DFFARX1 I_20997 (I100110,I2859,I359728,I359853,);
nand I_20998 (I359861,I359853,I100107);
not I_20999 (I359878,I359861);
DFFARX1 I_21000 (I359878,I2859,I359728,I359904,);
not I_21001 (I359912,I359904);
nor I_21002 (I359720,I359762,I359912);
DFFARX1 I_21003 (I100101,I2859,I359728,I359952,);
nor I_21004 (I359711,I359952,I359822);
nor I_21005 (I359702,I359952,I359878);
nand I_21006 (I359988,I100092,I100116);
and I_21007 (I360005,I359988,I100095);
DFFARX1 I_21008 (I360005,I2859,I359728,I360031,);
not I_21009 (I360039,I360031);
nand I_21010 (I360056,I360039,I359952);
nand I_21011 (I359705,I360039,I359861);
nor I_21012 (I360087,I100092,I100116);
and I_21013 (I360104,I359952,I360087);
nor I_21014 (I360121,I360039,I360104);
DFFARX1 I_21015 (I360121,I2859,I359728,I359714,);
nor I_21016 (I360152,I359754,I360087);
DFFARX1 I_21017 (I360152,I2859,I359728,I359699,);
nor I_21018 (I360183,I360031,I360087);
not I_21019 (I360200,I360183);
nand I_21020 (I359708,I360200,I360056);
not I_21021 (I360255,I2866);
DFFARX1 I_21022 (I381190,I2859,I360255,I360281,);
not I_21023 (I360289,I360281);
nand I_21024 (I360306,I381205,I381187);
and I_21025 (I360323,I360306,I381187);
DFFARX1 I_21026 (I360323,I2859,I360255,I360349,);
DFFARX1 I_21027 (I360349,I2859,I360255,I360244,);
DFFARX1 I_21028 (I381196,I2859,I360255,I360380,);
nand I_21029 (I360388,I360380,I381214);
not I_21030 (I360405,I360388);
DFFARX1 I_21031 (I360405,I2859,I360255,I360431,);
not I_21032 (I360439,I360431);
nor I_21033 (I360247,I360289,I360439);
DFFARX1 I_21034 (I381211,I2859,I360255,I360479,);
nor I_21035 (I360238,I360479,I360349);
nor I_21036 (I360229,I360479,I360405);
nand I_21037 (I360515,I381208,I381199);
and I_21038 (I360532,I360515,I381193);
DFFARX1 I_21039 (I360532,I2859,I360255,I360558,);
not I_21040 (I360566,I360558);
nand I_21041 (I360583,I360566,I360479);
nand I_21042 (I360232,I360566,I360388);
nor I_21043 (I360614,I381202,I381199);
and I_21044 (I360631,I360479,I360614);
nor I_21045 (I360648,I360566,I360631);
DFFARX1 I_21046 (I360648,I2859,I360255,I360241,);
nor I_21047 (I360679,I360281,I360614);
DFFARX1 I_21048 (I360679,I2859,I360255,I360226,);
nor I_21049 (I360710,I360558,I360614);
not I_21050 (I360727,I360710);
nand I_21051 (I360235,I360727,I360583);
not I_21052 (I360782,I2866);
DFFARX1 I_21053 (I503582,I2859,I360782,I360808,);
not I_21054 (I360816,I360808);
nand I_21055 (I360833,I503588,I503570);
and I_21056 (I360850,I360833,I503579);
DFFARX1 I_21057 (I360850,I2859,I360782,I360876,);
DFFARX1 I_21058 (I360876,I2859,I360782,I360771,);
DFFARX1 I_21059 (I503585,I2859,I360782,I360907,);
nand I_21060 (I360915,I360907,I503573);
not I_21061 (I360932,I360915);
DFFARX1 I_21062 (I360932,I2859,I360782,I360958,);
not I_21063 (I360966,I360958);
nor I_21064 (I360774,I360816,I360966);
DFFARX1 I_21065 (I503591,I2859,I360782,I361006,);
nor I_21066 (I360765,I361006,I360876);
nor I_21067 (I360756,I361006,I360932);
nand I_21068 (I361042,I503570,I503576);
and I_21069 (I361059,I361042,I503594);
DFFARX1 I_21070 (I361059,I2859,I360782,I361085,);
not I_21071 (I361093,I361085);
nand I_21072 (I361110,I361093,I361006);
nand I_21073 (I360759,I361093,I360915);
nor I_21074 (I361141,I503573,I503576);
and I_21075 (I361158,I361006,I361141);
nor I_21076 (I361175,I361093,I361158);
DFFARX1 I_21077 (I361175,I2859,I360782,I360768,);
nor I_21078 (I361206,I360808,I361141);
DFFARX1 I_21079 (I361206,I2859,I360782,I360753,);
nor I_21080 (I361237,I361085,I361141);
not I_21081 (I361254,I361237);
nand I_21082 (I360762,I361254,I361110);
not I_21083 (I361309,I2866);
DFFARX1 I_21084 (I48028,I2859,I361309,I361335,);
not I_21085 (I361343,I361335);
nand I_21086 (I361360,I48004,I48013);
and I_21087 (I361377,I361360,I48007);
DFFARX1 I_21088 (I361377,I2859,I361309,I361403,);
DFFARX1 I_21089 (I361403,I2859,I361309,I361298,);
DFFARX1 I_21090 (I48025,I2859,I361309,I361434,);
nand I_21091 (I361442,I361434,I48016);
not I_21092 (I361459,I361442);
DFFARX1 I_21093 (I361459,I2859,I361309,I361485,);
not I_21094 (I361493,I361485);
nor I_21095 (I361301,I361343,I361493);
DFFARX1 I_21096 (I48010,I2859,I361309,I361533,);
nor I_21097 (I361292,I361533,I361403);
nor I_21098 (I361283,I361533,I361459);
nand I_21099 (I361569,I48022,I48019);
and I_21100 (I361586,I361569,I48007);
DFFARX1 I_21101 (I361586,I2859,I361309,I361612,);
not I_21102 (I361620,I361612);
nand I_21103 (I361637,I361620,I361533);
nand I_21104 (I361286,I361620,I361442);
nor I_21105 (I361668,I48004,I48019);
and I_21106 (I361685,I361533,I361668);
nor I_21107 (I361702,I361620,I361685);
DFFARX1 I_21108 (I361702,I2859,I361309,I361295,);
nor I_21109 (I361733,I361335,I361668);
DFFARX1 I_21110 (I361733,I2859,I361309,I361280,);
nor I_21111 (I361764,I361612,I361668);
not I_21112 (I361781,I361764);
nand I_21113 (I361289,I361781,I361637);
not I_21114 (I361842,I2866);
DFFARX1 I_21115 (I128788,I2859,I361842,I361868,);
DFFARX1 I_21116 (I128794,I2859,I361842,I361885,);
not I_21117 (I361893,I361885);
not I_21118 (I361910,I128815);
nor I_21119 (I361927,I361910,I128803);
not I_21120 (I361944,I128812);
nor I_21121 (I361961,I361927,I128797);
nor I_21122 (I361978,I361885,I361961);
DFFARX1 I_21123 (I361978,I2859,I361842,I361828,);
nor I_21124 (I362009,I128797,I128803);
nand I_21125 (I362026,I362009,I128815);
DFFARX1 I_21126 (I362026,I2859,I361842,I361831,);
nor I_21127 (I362057,I361944,I128797);
nand I_21128 (I362074,I362057,I128788);
nor I_21129 (I362091,I361868,I362074);
DFFARX1 I_21130 (I362091,I2859,I361842,I361807,);
not I_21131 (I362122,I362074);
nand I_21132 (I361819,I361885,I362122);
DFFARX1 I_21133 (I362074,I2859,I361842,I362162,);
not I_21134 (I362170,I362162);
not I_21135 (I362187,I128797);
not I_21136 (I362204,I128800);
nor I_21137 (I362221,I362204,I128812);
nor I_21138 (I361834,I362170,I362221);
nor I_21139 (I362252,I362204,I128809);
and I_21140 (I362269,I362252,I128791);
or I_21141 (I362286,I362269,I128806);
DFFARX1 I_21142 (I362286,I2859,I361842,I362312,);
nor I_21143 (I361822,I362312,I361868);
not I_21144 (I362334,I362312);
and I_21145 (I362351,I362334,I361868);
nor I_21146 (I361816,I361893,I362351);
nand I_21147 (I362382,I362334,I361944);
nor I_21148 (I361810,I362204,I362382);
nand I_21149 (I361813,I362334,I362122);
nand I_21150 (I362427,I361944,I128800);
nor I_21151 (I361825,I362187,I362427);
not I_21152 (I362488,I2866);
DFFARX1 I_21153 (I90578,I2859,I362488,I362514,);
DFFARX1 I_21154 (I90590,I2859,I362488,I362531,);
not I_21155 (I362539,I362531);
not I_21156 (I362556,I90596);
nor I_21157 (I362573,I362556,I90581);
not I_21158 (I362590,I90572);
nor I_21159 (I362607,I362573,I90593);
nor I_21160 (I362624,I362531,I362607);
DFFARX1 I_21161 (I362624,I2859,I362488,I362474,);
nor I_21162 (I362655,I90593,I90581);
nand I_21163 (I362672,I362655,I90596);
DFFARX1 I_21164 (I362672,I2859,I362488,I362477,);
nor I_21165 (I362703,I362590,I90593);
nand I_21166 (I362720,I362703,I90575);
nor I_21167 (I362737,I362514,I362720);
DFFARX1 I_21168 (I362737,I2859,I362488,I362453,);
not I_21169 (I362768,I362720);
nand I_21170 (I362465,I362531,I362768);
DFFARX1 I_21171 (I362720,I2859,I362488,I362808,);
not I_21172 (I362816,I362808);
not I_21173 (I362833,I90593);
not I_21174 (I362850,I90584);
nor I_21175 (I362867,I362850,I90572);
nor I_21176 (I362480,I362816,I362867);
nor I_21177 (I362898,I362850,I90587);
and I_21178 (I362915,I362898,I90575);
or I_21179 (I362932,I362915,I90572);
DFFARX1 I_21180 (I362932,I2859,I362488,I362958,);
nor I_21181 (I362468,I362958,I362514);
not I_21182 (I362980,I362958);
and I_21183 (I362997,I362980,I362514);
nor I_21184 (I362462,I362539,I362997);
nand I_21185 (I363028,I362980,I362590);
nor I_21186 (I362456,I362850,I363028);
nand I_21187 (I362459,I362980,I362768);
nand I_21188 (I363073,I362590,I90584);
nor I_21189 (I362471,I362833,I363073);
not I_21190 (I363134,I2866);
DFFARX1 I_21191 (I467820,I2859,I363134,I363160,);
DFFARX1 I_21192 (I467802,I2859,I363134,I363177,);
not I_21193 (I363185,I363177);
not I_21194 (I363202,I467811);
nor I_21195 (I363219,I363202,I467823);
not I_21196 (I363236,I467805);
nor I_21197 (I363253,I363219,I467814);
nor I_21198 (I363270,I363177,I363253);
DFFARX1 I_21199 (I363270,I2859,I363134,I363120,);
nor I_21200 (I363301,I467814,I467823);
nand I_21201 (I363318,I363301,I467811);
DFFARX1 I_21202 (I363318,I2859,I363134,I363123,);
nor I_21203 (I363349,I363236,I467814);
nand I_21204 (I363366,I363349,I467826);
nor I_21205 (I363383,I363160,I363366);
DFFARX1 I_21206 (I363383,I2859,I363134,I363099,);
not I_21207 (I363414,I363366);
nand I_21208 (I363111,I363177,I363414);
DFFARX1 I_21209 (I363366,I2859,I363134,I363454,);
not I_21210 (I363462,I363454);
not I_21211 (I363479,I467814);
not I_21212 (I363496,I467802);
nor I_21213 (I363513,I363496,I467805);
nor I_21214 (I363126,I363462,I363513);
nor I_21215 (I363544,I363496,I467808);
and I_21216 (I363561,I363544,I467817);
or I_21217 (I363578,I363561,I467805);
DFFARX1 I_21218 (I363578,I2859,I363134,I363604,);
nor I_21219 (I363114,I363604,I363160);
not I_21220 (I363626,I363604);
and I_21221 (I363643,I363626,I363160);
nor I_21222 (I363108,I363185,I363643);
nand I_21223 (I363674,I363626,I363236);
nor I_21224 (I363102,I363496,I363674);
nand I_21225 (I363105,I363626,I363414);
nand I_21226 (I363719,I363236,I467802);
nor I_21227 (I363117,I363479,I363719);
not I_21228 (I363780,I2866);
DFFARX1 I_21229 (I87603,I2859,I363780,I363806,);
DFFARX1 I_21230 (I87615,I2859,I363780,I363823,);
not I_21231 (I363831,I363823);
not I_21232 (I363848,I87621);
nor I_21233 (I363865,I363848,I87606);
not I_21234 (I363882,I87597);
nor I_21235 (I363899,I363865,I87618);
nor I_21236 (I363916,I363823,I363899);
DFFARX1 I_21237 (I363916,I2859,I363780,I363766,);
nor I_21238 (I363947,I87618,I87606);
nand I_21239 (I363964,I363947,I87621);
DFFARX1 I_21240 (I363964,I2859,I363780,I363769,);
nor I_21241 (I363995,I363882,I87618);
nand I_21242 (I364012,I363995,I87600);
nor I_21243 (I364029,I363806,I364012);
DFFARX1 I_21244 (I364029,I2859,I363780,I363745,);
not I_21245 (I364060,I364012);
nand I_21246 (I363757,I363823,I364060);
DFFARX1 I_21247 (I364012,I2859,I363780,I364100,);
not I_21248 (I364108,I364100);
not I_21249 (I364125,I87618);
not I_21250 (I364142,I87609);
nor I_21251 (I364159,I364142,I87597);
nor I_21252 (I363772,I364108,I364159);
nor I_21253 (I364190,I364142,I87612);
and I_21254 (I364207,I364190,I87600);
or I_21255 (I364224,I364207,I87597);
DFFARX1 I_21256 (I364224,I2859,I363780,I364250,);
nor I_21257 (I363760,I364250,I363806);
not I_21258 (I364272,I364250);
and I_21259 (I364289,I364272,I363806);
nor I_21260 (I363754,I363831,I364289);
nand I_21261 (I364320,I364272,I363882);
nor I_21262 (I363748,I364142,I364320);
nand I_21263 (I363751,I364272,I364060);
nand I_21264 (I364365,I363882,I87609);
nor I_21265 (I363763,I364125,I364365);
not I_21266 (I364426,I2866);
DFFARX1 I_21267 (I240617,I2859,I364426,I364452,);
DFFARX1 I_21268 (I240629,I2859,I364426,I364469,);
not I_21269 (I364477,I364469);
not I_21270 (I364494,I240638);
nor I_21271 (I364511,I364494,I240614);
not I_21272 (I364528,I240632);
nor I_21273 (I364545,I364511,I240626);
nor I_21274 (I364562,I364469,I364545);
DFFARX1 I_21275 (I364562,I2859,I364426,I364412,);
nor I_21276 (I364593,I240626,I240614);
nand I_21277 (I364610,I364593,I240638);
DFFARX1 I_21278 (I364610,I2859,I364426,I364415,);
nor I_21279 (I364641,I364528,I240626);
nand I_21280 (I364658,I364641,I240620);
nor I_21281 (I364675,I364452,I364658);
DFFARX1 I_21282 (I364675,I2859,I364426,I364391,);
not I_21283 (I364706,I364658);
nand I_21284 (I364403,I364469,I364706);
DFFARX1 I_21285 (I364658,I2859,I364426,I364746,);
not I_21286 (I364754,I364746);
not I_21287 (I364771,I240626);
not I_21288 (I364788,I240635);
nor I_21289 (I364805,I364788,I240632);
nor I_21290 (I364418,I364754,I364805);
nor I_21291 (I364836,I364788,I240617);
and I_21292 (I364853,I364836,I240614);
or I_21293 (I364870,I364853,I240623);
DFFARX1 I_21294 (I364870,I2859,I364426,I364896,);
nor I_21295 (I364406,I364896,I364452);
not I_21296 (I364918,I364896);
and I_21297 (I364935,I364918,I364452);
nor I_21298 (I364400,I364477,I364935);
nand I_21299 (I364966,I364918,I364528);
nor I_21300 (I364394,I364788,I364966);
nand I_21301 (I364397,I364918,I364706);
nand I_21302 (I365011,I364528,I240635);
nor I_21303 (I364409,I364771,I365011);
not I_21304 (I365072,I2866);
DFFARX1 I_21305 (I13749,I2859,I365072,I365098,);
DFFARX1 I_21306 (I13755,I2859,I365072,I365115,);
not I_21307 (I365123,I365115);
not I_21308 (I365140,I13749);
nor I_21309 (I365157,I365140,I13761);
not I_21310 (I365174,I13773);
nor I_21311 (I365191,I365157,I13767);
nor I_21312 (I365208,I365115,I365191);
DFFARX1 I_21313 (I365208,I2859,I365072,I365058,);
nor I_21314 (I365239,I13767,I13761);
nand I_21315 (I365256,I365239,I13749);
DFFARX1 I_21316 (I365256,I2859,I365072,I365061,);
nor I_21317 (I365287,I365174,I13767);
nand I_21318 (I365304,I365287,I13752);
nor I_21319 (I365321,I365098,I365304);
DFFARX1 I_21320 (I365321,I2859,I365072,I365037,);
not I_21321 (I365352,I365304);
nand I_21322 (I365049,I365115,I365352);
DFFARX1 I_21323 (I365304,I2859,I365072,I365392,);
not I_21324 (I365400,I365392);
not I_21325 (I365417,I13767);
not I_21326 (I365434,I13752);
nor I_21327 (I365451,I365434,I13773);
nor I_21328 (I365064,I365400,I365451);
nor I_21329 (I365482,I365434,I13770);
and I_21330 (I365499,I365482,I13764);
or I_21331 (I365516,I365499,I13758);
DFFARX1 I_21332 (I365516,I2859,I365072,I365542,);
nor I_21333 (I365052,I365542,I365098);
not I_21334 (I365564,I365542);
and I_21335 (I365581,I365564,I365098);
nor I_21336 (I365046,I365123,I365581);
nand I_21337 (I365612,I365564,I365174);
nor I_21338 (I365040,I365434,I365612);
nand I_21339 (I365043,I365564,I365352);
nand I_21340 (I365657,I365174,I13752);
nor I_21341 (I365055,I365417,I365657);
not I_21342 (I365718,I2866);
DFFARX1 I_21343 (I57853,I2859,I365718,I365744,);
DFFARX1 I_21344 (I57865,I2859,I365718,I365761,);
not I_21345 (I365769,I365761);
not I_21346 (I365786,I57871);
nor I_21347 (I365803,I365786,I57856);
not I_21348 (I365820,I57847);
nor I_21349 (I365837,I365803,I57868);
nor I_21350 (I365854,I365761,I365837);
DFFARX1 I_21351 (I365854,I2859,I365718,I365704,);
nor I_21352 (I365885,I57868,I57856);
nand I_21353 (I365902,I365885,I57871);
DFFARX1 I_21354 (I365902,I2859,I365718,I365707,);
nor I_21355 (I365933,I365820,I57868);
nand I_21356 (I365950,I365933,I57850);
nor I_21357 (I365967,I365744,I365950);
DFFARX1 I_21358 (I365967,I2859,I365718,I365683,);
not I_21359 (I365998,I365950);
nand I_21360 (I365695,I365761,I365998);
DFFARX1 I_21361 (I365950,I2859,I365718,I366038,);
not I_21362 (I366046,I366038);
not I_21363 (I366063,I57868);
not I_21364 (I366080,I57859);
nor I_21365 (I366097,I366080,I57847);
nor I_21366 (I365710,I366046,I366097);
nor I_21367 (I366128,I366080,I57862);
and I_21368 (I366145,I366128,I57850);
or I_21369 (I366162,I366145,I57847);
DFFARX1 I_21370 (I366162,I2859,I365718,I366188,);
nor I_21371 (I365698,I366188,I365744);
not I_21372 (I366210,I366188);
and I_21373 (I366227,I366210,I365744);
nor I_21374 (I365692,I365769,I366227);
nand I_21375 (I366258,I366210,I365820);
nor I_21376 (I365686,I366080,I366258);
nand I_21377 (I365689,I366210,I365998);
nand I_21378 (I366303,I365820,I57859);
nor I_21379 (I365701,I366063,I366303);
not I_21380 (I366364,I2866);
DFFARX1 I_21381 (I219163,I2859,I366364,I366390,);
DFFARX1 I_21382 (I219175,I2859,I366364,I366407,);
not I_21383 (I366415,I366407);
not I_21384 (I366432,I219160);
nor I_21385 (I366449,I366432,I219178);
not I_21386 (I366466,I219184);
nor I_21387 (I366483,I366449,I219166);
nor I_21388 (I366500,I366407,I366483);
DFFARX1 I_21389 (I366500,I2859,I366364,I366350,);
nor I_21390 (I366531,I219166,I219178);
nand I_21391 (I366548,I366531,I219160);
DFFARX1 I_21392 (I366548,I2859,I366364,I366353,);
nor I_21393 (I366579,I366466,I219166);
nand I_21394 (I366596,I366579,I219169);
nor I_21395 (I366613,I366390,I366596);
DFFARX1 I_21396 (I366613,I2859,I366364,I366329,);
not I_21397 (I366644,I366596);
nand I_21398 (I366341,I366407,I366644);
DFFARX1 I_21399 (I366596,I2859,I366364,I366684,);
not I_21400 (I366692,I366684);
not I_21401 (I366709,I219166);
not I_21402 (I366726,I219172);
nor I_21403 (I366743,I366726,I219184);
nor I_21404 (I366356,I366692,I366743);
nor I_21405 (I366774,I366726,I219181);
and I_21406 (I366791,I366774,I219160);
or I_21407 (I366808,I366791,I219163);
DFFARX1 I_21408 (I366808,I2859,I366364,I366834,);
nor I_21409 (I366344,I366834,I366390);
not I_21410 (I366856,I366834);
and I_21411 (I366873,I366856,I366390);
nor I_21412 (I366338,I366415,I366873);
nand I_21413 (I366904,I366856,I366466);
nor I_21414 (I366332,I366726,I366904);
nand I_21415 (I366335,I366856,I366644);
nand I_21416 (I366949,I366466,I219172);
nor I_21417 (I366347,I366709,I366949);
not I_21418 (I367010,I2866);
DFFARX1 I_21419 (I21654,I2859,I367010,I367036,);
DFFARX1 I_21420 (I21660,I2859,I367010,I367053,);
not I_21421 (I367061,I367053);
not I_21422 (I367078,I21678);
nor I_21423 (I367095,I367078,I21657);
not I_21424 (I367112,I21663);
nor I_21425 (I367129,I367095,I21669);
nor I_21426 (I367146,I367053,I367129);
DFFARX1 I_21427 (I367146,I2859,I367010,I366996,);
nor I_21428 (I367177,I21669,I21657);
nand I_21429 (I367194,I367177,I21678);
DFFARX1 I_21430 (I367194,I2859,I367010,I366999,);
nor I_21431 (I367225,I367112,I21669);
nand I_21432 (I367242,I367225,I21675);
nor I_21433 (I367259,I367036,I367242);
DFFARX1 I_21434 (I367259,I2859,I367010,I366975,);
not I_21435 (I367290,I367242);
nand I_21436 (I366987,I367053,I367290);
DFFARX1 I_21437 (I367242,I2859,I367010,I367330,);
not I_21438 (I367338,I367330);
not I_21439 (I367355,I21669);
not I_21440 (I367372,I21657);
nor I_21441 (I367389,I367372,I21663);
nor I_21442 (I367002,I367338,I367389);
nor I_21443 (I367420,I367372,I21666);
and I_21444 (I367437,I367420,I21654);
or I_21445 (I367454,I367437,I21672);
DFFARX1 I_21446 (I367454,I2859,I367010,I367480,);
nor I_21447 (I366990,I367480,I367036);
not I_21448 (I367502,I367480);
and I_21449 (I367519,I367502,I367036);
nor I_21450 (I366984,I367061,I367519);
nand I_21451 (I367550,I367502,I367112);
nor I_21452 (I366978,I367372,I367550);
nand I_21453 (I366981,I367502,I367290);
nand I_21454 (I367595,I367112,I21657);
nor I_21455 (I366993,I367355,I367595);
not I_21456 (I367656,I2866);
DFFARX1 I_21457 (I252755,I2859,I367656,I367682,);
DFFARX1 I_21458 (I252767,I2859,I367656,I367699,);
not I_21459 (I367707,I367699);
not I_21460 (I367724,I252776);
nor I_21461 (I367741,I367724,I252752);
not I_21462 (I367758,I252770);
nor I_21463 (I367775,I367741,I252764);
nor I_21464 (I367792,I367699,I367775);
DFFARX1 I_21465 (I367792,I2859,I367656,I367642,);
nor I_21466 (I367823,I252764,I252752);
nand I_21467 (I367840,I367823,I252776);
DFFARX1 I_21468 (I367840,I2859,I367656,I367645,);
nor I_21469 (I367871,I367758,I252764);
nand I_21470 (I367888,I367871,I252758);
nor I_21471 (I367905,I367682,I367888);
DFFARX1 I_21472 (I367905,I2859,I367656,I367621,);
not I_21473 (I367936,I367888);
nand I_21474 (I367633,I367699,I367936);
DFFARX1 I_21475 (I367888,I2859,I367656,I367976,);
not I_21476 (I367984,I367976);
not I_21477 (I368001,I252764);
not I_21478 (I368018,I252773);
nor I_21479 (I368035,I368018,I252770);
nor I_21480 (I367648,I367984,I368035);
nor I_21481 (I368066,I368018,I252755);
and I_21482 (I368083,I368066,I252752);
or I_21483 (I368100,I368083,I252761);
DFFARX1 I_21484 (I368100,I2859,I367656,I368126,);
nor I_21485 (I367636,I368126,I367682);
not I_21486 (I368148,I368126);
and I_21487 (I368165,I368148,I367682);
nor I_21488 (I367630,I367707,I368165);
nand I_21489 (I368196,I368148,I367758);
nor I_21490 (I367624,I368018,I368196);
nand I_21491 (I367627,I368148,I367936);
nand I_21492 (I368241,I367758,I252773);
nor I_21493 (I367639,I368001,I368241);
not I_21494 (I368302,I2866);
DFFARX1 I_21495 (I270098,I2859,I368302,I368328,);
DFFARX1 I_21496 (I270092,I2859,I368302,I368345,);
not I_21497 (I368353,I368345);
not I_21498 (I368370,I270107);
nor I_21499 (I368387,I368370,I270092);
not I_21500 (I368404,I270101);
nor I_21501 (I368421,I368387,I270110);
nor I_21502 (I368438,I368345,I368421);
DFFARX1 I_21503 (I368438,I2859,I368302,I368288,);
nor I_21504 (I368469,I270110,I270092);
nand I_21505 (I368486,I368469,I270107);
DFFARX1 I_21506 (I368486,I2859,I368302,I368291,);
nor I_21507 (I368517,I368404,I270110);
nand I_21508 (I368534,I368517,I270095);
nor I_21509 (I368551,I368328,I368534);
DFFARX1 I_21510 (I368551,I2859,I368302,I368267,);
not I_21511 (I368582,I368534);
nand I_21512 (I368279,I368345,I368582);
DFFARX1 I_21513 (I368534,I2859,I368302,I368622,);
not I_21514 (I368630,I368622);
not I_21515 (I368647,I270110);
not I_21516 (I368664,I270104);
nor I_21517 (I368681,I368664,I270101);
nor I_21518 (I368294,I368630,I368681);
nor I_21519 (I368712,I368664,I270113);
and I_21520 (I368729,I368712,I270116);
or I_21521 (I368746,I368729,I270095);
DFFARX1 I_21522 (I368746,I2859,I368302,I368772,);
nor I_21523 (I368282,I368772,I368328);
not I_21524 (I368794,I368772);
and I_21525 (I368811,I368794,I368328);
nor I_21526 (I368276,I368353,I368811);
nand I_21527 (I368842,I368794,I368404);
nor I_21528 (I368270,I368664,I368842);
nand I_21529 (I368273,I368794,I368582);
nand I_21530 (I368887,I368404,I270104);
nor I_21531 (I368285,I368647,I368887);
not I_21532 (I368948,I2866);
DFFARX1 I_21533 (I453948,I2859,I368948,I368974,);
DFFARX1 I_21534 (I453930,I2859,I368948,I368991,);
not I_21535 (I368999,I368991);
not I_21536 (I369016,I453939);
nor I_21537 (I369033,I369016,I453951);
not I_21538 (I369050,I453933);
nor I_21539 (I369067,I369033,I453942);
nor I_21540 (I369084,I368991,I369067);
DFFARX1 I_21541 (I369084,I2859,I368948,I368934,);
nor I_21542 (I369115,I453942,I453951);
nand I_21543 (I369132,I369115,I453939);
DFFARX1 I_21544 (I369132,I2859,I368948,I368937,);
nor I_21545 (I369163,I369050,I453942);
nand I_21546 (I369180,I369163,I453954);
nor I_21547 (I369197,I368974,I369180);
DFFARX1 I_21548 (I369197,I2859,I368948,I368913,);
not I_21549 (I369228,I369180);
nand I_21550 (I368925,I368991,I369228);
DFFARX1 I_21551 (I369180,I2859,I368948,I369268,);
not I_21552 (I369276,I369268);
not I_21553 (I369293,I453942);
not I_21554 (I369310,I453930);
nor I_21555 (I369327,I369310,I453933);
nor I_21556 (I368940,I369276,I369327);
nor I_21557 (I369358,I369310,I453936);
and I_21558 (I369375,I369358,I453945);
or I_21559 (I369392,I369375,I453933);
DFFARX1 I_21560 (I369392,I2859,I368948,I369418,);
nor I_21561 (I368928,I369418,I368974);
not I_21562 (I369440,I369418);
and I_21563 (I369457,I369440,I368974);
nor I_21564 (I368922,I368999,I369457);
nand I_21565 (I369488,I369440,I369050);
nor I_21566 (I368916,I369310,I369488);
nand I_21567 (I368919,I369440,I369228);
nand I_21568 (I369533,I369050,I453930);
nor I_21569 (I368931,I369293,I369533);
not I_21570 (I369594,I2866);
DFFARX1 I_21571 (I297842,I2859,I369594,I369620,);
DFFARX1 I_21572 (I297836,I2859,I369594,I369637,);
not I_21573 (I369645,I369637);
not I_21574 (I369662,I297851);
nor I_21575 (I369679,I369662,I297836);
not I_21576 (I369696,I297845);
nor I_21577 (I369713,I369679,I297854);
nor I_21578 (I369730,I369637,I369713);
DFFARX1 I_21579 (I369730,I2859,I369594,I369580,);
nor I_21580 (I369761,I297854,I297836);
nand I_21581 (I369778,I369761,I297851);
DFFARX1 I_21582 (I369778,I2859,I369594,I369583,);
nor I_21583 (I369809,I369696,I297854);
nand I_21584 (I369826,I369809,I297839);
nor I_21585 (I369843,I369620,I369826);
DFFARX1 I_21586 (I369843,I2859,I369594,I369559,);
not I_21587 (I369874,I369826);
nand I_21588 (I369571,I369637,I369874);
DFFARX1 I_21589 (I369826,I2859,I369594,I369914,);
not I_21590 (I369922,I369914);
not I_21591 (I369939,I297854);
not I_21592 (I369956,I297848);
nor I_21593 (I369973,I369956,I297845);
nor I_21594 (I369586,I369922,I369973);
nor I_21595 (I370004,I369956,I297857);
and I_21596 (I370021,I370004,I297860);
or I_21597 (I370038,I370021,I297839);
DFFARX1 I_21598 (I370038,I2859,I369594,I370064,);
nor I_21599 (I369574,I370064,I369620);
not I_21600 (I370086,I370064);
and I_21601 (I370103,I370086,I369620);
nor I_21602 (I369568,I369645,I370103);
nand I_21603 (I370134,I370086,I369696);
nor I_21604 (I369562,I369956,I370134);
nand I_21605 (I369565,I370086,I369874);
nand I_21606 (I370179,I369696,I297848);
nor I_21607 (I369577,I369939,I370179);
not I_21608 (I370240,I2866);
DFFARX1 I_21609 (I278190,I2859,I370240,I370266,);
DFFARX1 I_21610 (I278184,I2859,I370240,I370283,);
not I_21611 (I370291,I370283);
not I_21612 (I370308,I278199);
nor I_21613 (I370325,I370308,I278184);
not I_21614 (I370342,I278193);
nor I_21615 (I370359,I370325,I278202);
nor I_21616 (I370376,I370283,I370359);
DFFARX1 I_21617 (I370376,I2859,I370240,I370226,);
nor I_21618 (I370407,I278202,I278184);
nand I_21619 (I370424,I370407,I278199);
DFFARX1 I_21620 (I370424,I2859,I370240,I370229,);
nor I_21621 (I370455,I370342,I278202);
nand I_21622 (I370472,I370455,I278187);
nor I_21623 (I370489,I370266,I370472);
DFFARX1 I_21624 (I370489,I2859,I370240,I370205,);
not I_21625 (I370520,I370472);
nand I_21626 (I370217,I370283,I370520);
DFFARX1 I_21627 (I370472,I2859,I370240,I370560,);
not I_21628 (I370568,I370560);
not I_21629 (I370585,I278202);
not I_21630 (I370602,I278196);
nor I_21631 (I370619,I370602,I278193);
nor I_21632 (I370232,I370568,I370619);
nor I_21633 (I370650,I370602,I278205);
and I_21634 (I370667,I370650,I278208);
or I_21635 (I370684,I370667,I278187);
DFFARX1 I_21636 (I370684,I2859,I370240,I370710,);
nor I_21637 (I370220,I370710,I370266);
not I_21638 (I370732,I370710);
and I_21639 (I370749,I370732,I370266);
nor I_21640 (I370214,I370291,I370749);
nand I_21641 (I370780,I370732,I370342);
nor I_21642 (I370208,I370602,I370780);
nand I_21643 (I370211,I370732,I370520);
nand I_21644 (I370825,I370342,I278196);
nor I_21645 (I370223,I370585,I370825);
not I_21646 (I370886,I2866);
DFFARX1 I_21647 (I462618,I2859,I370886,I370912,);
DFFARX1 I_21648 (I462600,I2859,I370886,I370929,);
not I_21649 (I370937,I370929);
not I_21650 (I370954,I462609);
nor I_21651 (I370971,I370954,I462621);
not I_21652 (I370988,I462603);
nor I_21653 (I371005,I370971,I462612);
nor I_21654 (I371022,I370929,I371005);
DFFARX1 I_21655 (I371022,I2859,I370886,I370872,);
nor I_21656 (I371053,I462612,I462621);
nand I_21657 (I371070,I371053,I462609);
DFFARX1 I_21658 (I371070,I2859,I370886,I370875,);
nor I_21659 (I371101,I370988,I462612);
nand I_21660 (I371118,I371101,I462624);
nor I_21661 (I371135,I370912,I371118);
DFFARX1 I_21662 (I371135,I2859,I370886,I370851,);
not I_21663 (I371166,I371118);
nand I_21664 (I370863,I370929,I371166);
DFFARX1 I_21665 (I371118,I2859,I370886,I371206,);
not I_21666 (I371214,I371206);
not I_21667 (I371231,I462612);
not I_21668 (I371248,I462600);
nor I_21669 (I371265,I371248,I462603);
nor I_21670 (I370878,I371214,I371265);
nor I_21671 (I371296,I371248,I462606);
and I_21672 (I371313,I371296,I462615);
or I_21673 (I371330,I371313,I462603);
DFFARX1 I_21674 (I371330,I2859,I370886,I371356,);
nor I_21675 (I370866,I371356,I370912);
not I_21676 (I371378,I371356);
and I_21677 (I371395,I371378,I370912);
nor I_21678 (I370860,I370937,I371395);
nand I_21679 (I371426,I371378,I370988);
nor I_21680 (I370854,I371248,I371426);
nand I_21681 (I370857,I371378,I371166);
nand I_21682 (I371471,I370988,I462600);
nor I_21683 (I370869,I371231,I371471);
not I_21684 (I371532,I2866);
DFFARX1 I_21685 (I98908,I2859,I371532,I371558,);
DFFARX1 I_21686 (I98920,I2859,I371532,I371575,);
not I_21687 (I371583,I371575);
not I_21688 (I371600,I98926);
nor I_21689 (I371617,I371600,I98911);
not I_21690 (I371634,I98902);
nor I_21691 (I371651,I371617,I98923);
nor I_21692 (I371668,I371575,I371651);
DFFARX1 I_21693 (I371668,I2859,I371532,I371518,);
nor I_21694 (I371699,I98923,I98911);
nand I_21695 (I371716,I371699,I98926);
DFFARX1 I_21696 (I371716,I2859,I371532,I371521,);
nor I_21697 (I371747,I371634,I98923);
nand I_21698 (I371764,I371747,I98905);
nor I_21699 (I371781,I371558,I371764);
DFFARX1 I_21700 (I371781,I2859,I371532,I371497,);
not I_21701 (I371812,I371764);
nand I_21702 (I371509,I371575,I371812);
DFFARX1 I_21703 (I371764,I2859,I371532,I371852,);
not I_21704 (I371860,I371852);
not I_21705 (I371877,I98923);
not I_21706 (I371894,I98914);
nor I_21707 (I371911,I371894,I98902);
nor I_21708 (I371524,I371860,I371911);
nor I_21709 (I371942,I371894,I98917);
and I_21710 (I371959,I371942,I98905);
or I_21711 (I371976,I371959,I98902);
DFFARX1 I_21712 (I371976,I2859,I371532,I372002,);
nor I_21713 (I371512,I372002,I371558);
not I_21714 (I372024,I372002);
and I_21715 (I372041,I372024,I371558);
nor I_21716 (I371506,I371583,I372041);
nand I_21717 (I372072,I372024,I371634);
nor I_21718 (I371500,I371894,I372072);
nand I_21719 (I371503,I372024,I371812);
nand I_21720 (I372117,I371634,I98914);
nor I_21721 (I371515,I371877,I372117);
not I_21722 (I372178,I2866);
DFFARX1 I_21723 (I44842,I2859,I372178,I372204,);
DFFARX1 I_21724 (I44848,I2859,I372178,I372221,);
not I_21725 (I372229,I372221);
not I_21726 (I372246,I44866);
nor I_21727 (I372263,I372246,I44845);
not I_21728 (I372280,I44851);
nor I_21729 (I372297,I372263,I44857);
nor I_21730 (I372314,I372221,I372297);
DFFARX1 I_21731 (I372314,I2859,I372178,I372164,);
nor I_21732 (I372345,I44857,I44845);
nand I_21733 (I372362,I372345,I44866);
DFFARX1 I_21734 (I372362,I2859,I372178,I372167,);
nor I_21735 (I372393,I372280,I44857);
nand I_21736 (I372410,I372393,I44863);
nor I_21737 (I372427,I372204,I372410);
DFFARX1 I_21738 (I372427,I2859,I372178,I372143,);
not I_21739 (I372458,I372410);
nand I_21740 (I372155,I372221,I372458);
DFFARX1 I_21741 (I372410,I2859,I372178,I372498,);
not I_21742 (I372506,I372498);
not I_21743 (I372523,I44857);
not I_21744 (I372540,I44845);
nor I_21745 (I372557,I372540,I44851);
nor I_21746 (I372170,I372506,I372557);
nor I_21747 (I372588,I372540,I44854);
and I_21748 (I372605,I372588,I44842);
or I_21749 (I372622,I372605,I44860);
DFFARX1 I_21750 (I372622,I2859,I372178,I372648,);
nor I_21751 (I372158,I372648,I372204);
not I_21752 (I372670,I372648);
and I_21753 (I372687,I372670,I372204);
nor I_21754 (I372152,I372229,I372687);
nand I_21755 (I372718,I372670,I372280);
nor I_21756 (I372146,I372540,I372718);
nand I_21757 (I372149,I372670,I372458);
nand I_21758 (I372763,I372280,I44845);
nor I_21759 (I372161,I372523,I372763);
not I_21760 (I372824,I2866);
DFFARX1 I_21761 (I204288,I2859,I372824,I372850,);
DFFARX1 I_21762 (I204300,I2859,I372824,I372867,);
not I_21763 (I372875,I372867);
not I_21764 (I372892,I204285);
nor I_21765 (I372909,I372892,I204303);
not I_21766 (I372926,I204309);
nor I_21767 (I372943,I372909,I204291);
nor I_21768 (I372960,I372867,I372943);
DFFARX1 I_21769 (I372960,I2859,I372824,I372810,);
nor I_21770 (I372991,I204291,I204303);
nand I_21771 (I373008,I372991,I204285);
DFFARX1 I_21772 (I373008,I2859,I372824,I372813,);
nor I_21773 (I373039,I372926,I204291);
nand I_21774 (I373056,I373039,I204294);
nor I_21775 (I373073,I372850,I373056);
DFFARX1 I_21776 (I373073,I2859,I372824,I372789,);
not I_21777 (I373104,I373056);
nand I_21778 (I372801,I372867,I373104);
DFFARX1 I_21779 (I373056,I2859,I372824,I373144,);
not I_21780 (I373152,I373144);
not I_21781 (I373169,I204291);
not I_21782 (I373186,I204297);
nor I_21783 (I373203,I373186,I204309);
nor I_21784 (I372816,I373152,I373203);
nor I_21785 (I373234,I373186,I204306);
and I_21786 (I373251,I373234,I204285);
or I_21787 (I373268,I373251,I204288);
DFFARX1 I_21788 (I373268,I2859,I372824,I373294,);
nor I_21789 (I372804,I373294,I372850);
not I_21790 (I373316,I373294);
and I_21791 (I373333,I373316,I372850);
nor I_21792 (I372798,I372875,I373333);
nand I_21793 (I373364,I373316,I372926);
nor I_21794 (I372792,I373186,I373364);
nand I_21795 (I372795,I373316,I373104);
nand I_21796 (I373409,I372926,I204297);
nor I_21797 (I372807,I373169,I373409);
not I_21798 (I373470,I2866);
DFFARX1 I_21799 (I175102,I2859,I373470,I373496,);
DFFARX1 I_21800 (I175099,I2859,I373470,I373513,);
not I_21801 (I373521,I373513);
not I_21802 (I373538,I175114);
nor I_21803 (I373555,I373538,I175117);
not I_21804 (I373572,I175105);
nor I_21805 (I373589,I373555,I175111);
nor I_21806 (I373606,I373513,I373589);
DFFARX1 I_21807 (I373606,I2859,I373470,I373456,);
nor I_21808 (I373637,I175111,I175117);
nand I_21809 (I373654,I373637,I175114);
DFFARX1 I_21810 (I373654,I2859,I373470,I373459,);
nor I_21811 (I373685,I373572,I175111);
nand I_21812 (I373702,I373685,I175123);
nor I_21813 (I373719,I373496,I373702);
DFFARX1 I_21814 (I373719,I2859,I373470,I373435,);
not I_21815 (I373750,I373702);
nand I_21816 (I373447,I373513,I373750);
DFFARX1 I_21817 (I373702,I2859,I373470,I373790,);
not I_21818 (I373798,I373790);
not I_21819 (I373815,I175111);
not I_21820 (I373832,I175096);
nor I_21821 (I373849,I373832,I175105);
nor I_21822 (I373462,I373798,I373849);
nor I_21823 (I373880,I373832,I175108);
and I_21824 (I373897,I373880,I175096);
or I_21825 (I373914,I373897,I175120);
DFFARX1 I_21826 (I373914,I2859,I373470,I373940,);
nor I_21827 (I373450,I373940,I373496);
not I_21828 (I373962,I373940);
and I_21829 (I373979,I373962,I373496);
nor I_21830 (I373444,I373521,I373979);
nand I_21831 (I374010,I373962,I373572);
nor I_21832 (I373438,I373832,I374010);
nand I_21833 (I373441,I373962,I373750);
nand I_21834 (I374055,I373572,I175096);
nor I_21835 (I373453,I373815,I374055);
not I_21836 (I374116,I2866);
DFFARX1 I_21837 (I133004,I2859,I374116,I374142,);
DFFARX1 I_21838 (I133010,I2859,I374116,I374159,);
not I_21839 (I374167,I374159);
not I_21840 (I374184,I133031);
nor I_21841 (I374201,I374184,I133019);
not I_21842 (I374218,I133028);
nor I_21843 (I374235,I374201,I133013);
nor I_21844 (I374252,I374159,I374235);
DFFARX1 I_21845 (I374252,I2859,I374116,I374102,);
nor I_21846 (I374283,I133013,I133019);
nand I_21847 (I374300,I374283,I133031);
DFFARX1 I_21848 (I374300,I2859,I374116,I374105,);
nor I_21849 (I374331,I374218,I133013);
nand I_21850 (I374348,I374331,I133004);
nor I_21851 (I374365,I374142,I374348);
DFFARX1 I_21852 (I374365,I2859,I374116,I374081,);
not I_21853 (I374396,I374348);
nand I_21854 (I374093,I374159,I374396);
DFFARX1 I_21855 (I374348,I2859,I374116,I374436,);
not I_21856 (I374444,I374436);
not I_21857 (I374461,I133013);
not I_21858 (I374478,I133016);
nor I_21859 (I374495,I374478,I133028);
nor I_21860 (I374108,I374444,I374495);
nor I_21861 (I374526,I374478,I133025);
and I_21862 (I374543,I374526,I133007);
or I_21863 (I374560,I374543,I133022);
DFFARX1 I_21864 (I374560,I2859,I374116,I374586,);
nor I_21865 (I374096,I374586,I374142);
not I_21866 (I374608,I374586);
and I_21867 (I374625,I374608,I374142);
nor I_21868 (I374090,I374167,I374625);
nand I_21869 (I374656,I374608,I374218);
nor I_21870 (I374084,I374478,I374656);
nand I_21871 (I374087,I374608,I374396);
nand I_21872 (I374701,I374218,I133016);
nor I_21873 (I374099,I374461,I374701);
not I_21874 (I374762,I2866);
DFFARX1 I_21875 (I212023,I2859,I374762,I374788,);
DFFARX1 I_21876 (I212035,I2859,I374762,I374805,);
not I_21877 (I374813,I374805);
not I_21878 (I374830,I212020);
nor I_21879 (I374847,I374830,I212038);
not I_21880 (I374864,I212044);
nor I_21881 (I374881,I374847,I212026);
nor I_21882 (I374898,I374805,I374881);
DFFARX1 I_21883 (I374898,I2859,I374762,I374748,);
nor I_21884 (I374929,I212026,I212038);
nand I_21885 (I374946,I374929,I212020);
DFFARX1 I_21886 (I374946,I2859,I374762,I374751,);
nor I_21887 (I374977,I374864,I212026);
nand I_21888 (I374994,I374977,I212029);
nor I_21889 (I375011,I374788,I374994);
DFFARX1 I_21890 (I375011,I2859,I374762,I374727,);
not I_21891 (I375042,I374994);
nand I_21892 (I374739,I374805,I375042);
DFFARX1 I_21893 (I374994,I2859,I374762,I375082,);
not I_21894 (I375090,I375082);
not I_21895 (I375107,I212026);
not I_21896 (I375124,I212032);
nor I_21897 (I375141,I375124,I212044);
nor I_21898 (I374754,I375090,I375141);
nor I_21899 (I375172,I375124,I212041);
and I_21900 (I375189,I375172,I212020);
or I_21901 (I375206,I375189,I212023);
DFFARX1 I_21902 (I375206,I2859,I374762,I375232,);
nor I_21903 (I374742,I375232,I374788);
not I_21904 (I375254,I375232);
and I_21905 (I375271,I375254,I374788);
nor I_21906 (I374736,I374813,I375271);
nand I_21907 (I375302,I375254,I374864);
nor I_21908 (I374730,I375124,I375302);
nand I_21909 (I374733,I375254,I375042);
nand I_21910 (I375347,I374864,I212032);
nor I_21911 (I374745,I375107,I375347);
not I_21912 (I375408,I2866);
DFFARX1 I_21913 (I55473,I2859,I375408,I375434,);
DFFARX1 I_21914 (I55485,I2859,I375408,I375451,);
not I_21915 (I375459,I375451);
not I_21916 (I375476,I55491);
nor I_21917 (I375493,I375476,I55476);
not I_21918 (I375510,I55467);
nor I_21919 (I375527,I375493,I55488);
nor I_21920 (I375544,I375451,I375527);
DFFARX1 I_21921 (I375544,I2859,I375408,I375394,);
nor I_21922 (I375575,I55488,I55476);
nand I_21923 (I375592,I375575,I55491);
DFFARX1 I_21924 (I375592,I2859,I375408,I375397,);
nor I_21925 (I375623,I375510,I55488);
nand I_21926 (I375640,I375623,I55470);
nor I_21927 (I375657,I375434,I375640);
DFFARX1 I_21928 (I375657,I2859,I375408,I375373,);
not I_21929 (I375688,I375640);
nand I_21930 (I375385,I375451,I375688);
DFFARX1 I_21931 (I375640,I2859,I375408,I375728,);
not I_21932 (I375736,I375728);
not I_21933 (I375753,I55488);
not I_21934 (I375770,I55479);
nor I_21935 (I375787,I375770,I55467);
nor I_21936 (I375400,I375736,I375787);
nor I_21937 (I375818,I375770,I55482);
and I_21938 (I375835,I375818,I55470);
or I_21939 (I375852,I375835,I55467);
DFFARX1 I_21940 (I375852,I2859,I375408,I375878,);
nor I_21941 (I375388,I375878,I375434);
not I_21942 (I375900,I375878);
and I_21943 (I375917,I375900,I375434);
nor I_21944 (I375382,I375459,I375917);
nand I_21945 (I375948,I375900,I375510);
nor I_21946 (I375376,I375770,I375948);
nand I_21947 (I375379,I375900,I375688);
nand I_21948 (I375993,I375510,I55479);
nor I_21949 (I375391,I375753,I375993);
not I_21950 (I376054,I2866);
DFFARX1 I_21951 (I92363,I2859,I376054,I376080,);
DFFARX1 I_21952 (I92375,I2859,I376054,I376097,);
not I_21953 (I376105,I376097);
not I_21954 (I376122,I92381);
nor I_21955 (I376139,I376122,I92366);
not I_21956 (I376156,I92357);
nor I_21957 (I376173,I376139,I92378);
nor I_21958 (I376190,I376097,I376173);
DFFARX1 I_21959 (I376190,I2859,I376054,I376040,);
nor I_21960 (I376221,I92378,I92366);
nand I_21961 (I376238,I376221,I92381);
DFFARX1 I_21962 (I376238,I2859,I376054,I376043,);
nor I_21963 (I376269,I376156,I92378);
nand I_21964 (I376286,I376269,I92360);
nor I_21965 (I376303,I376080,I376286);
DFFARX1 I_21966 (I376303,I2859,I376054,I376019,);
not I_21967 (I376334,I376286);
nand I_21968 (I376031,I376097,I376334);
DFFARX1 I_21969 (I376286,I2859,I376054,I376374,);
not I_21970 (I376382,I376374);
not I_21971 (I376399,I92378);
not I_21972 (I376416,I92369);
nor I_21973 (I376433,I376416,I92357);
nor I_21974 (I376046,I376382,I376433);
nor I_21975 (I376464,I376416,I92372);
and I_21976 (I376481,I376464,I92360);
or I_21977 (I376498,I376481,I92357);
DFFARX1 I_21978 (I376498,I2859,I376054,I376524,);
nor I_21979 (I376034,I376524,I376080);
not I_21980 (I376546,I376524);
and I_21981 (I376563,I376546,I376080);
nor I_21982 (I376028,I376105,I376563);
nand I_21983 (I376594,I376546,I376156);
nor I_21984 (I376022,I376416,I376594);
nand I_21985 (I376025,I376546,I376334);
nand I_21986 (I376639,I376156,I92369);
nor I_21987 (I376037,I376399,I376639);
not I_21988 (I376700,I2866);
DFFARX1 I_21989 (I515556,I2859,I376700,I376726,);
DFFARX1 I_21990 (I515562,I2859,I376700,I376743,);
not I_21991 (I376751,I376743);
not I_21992 (I376768,I515559);
nor I_21993 (I376785,I376768,I515538);
not I_21994 (I376802,I515541);
nor I_21995 (I376819,I376785,I515547);
nor I_21996 (I376836,I376743,I376819);
DFFARX1 I_21997 (I376836,I2859,I376700,I376686,);
nor I_21998 (I376867,I515547,I515538);
nand I_21999 (I376884,I376867,I515559);
DFFARX1 I_22000 (I376884,I2859,I376700,I376689,);
nor I_22001 (I376915,I376802,I515547);
nand I_22002 (I376932,I376915,I515541);
nor I_22003 (I376949,I376726,I376932);
DFFARX1 I_22004 (I376949,I2859,I376700,I376665,);
not I_22005 (I376980,I376932);
nand I_22006 (I376677,I376743,I376980);
DFFARX1 I_22007 (I376932,I2859,I376700,I377020,);
not I_22008 (I377028,I377020);
not I_22009 (I377045,I515547);
not I_22010 (I377062,I515550);
nor I_22011 (I377079,I377062,I515541);
nor I_22012 (I376692,I377028,I377079);
nor I_22013 (I377110,I377062,I515538);
and I_22014 (I377127,I377110,I515544);
or I_22015 (I377144,I377127,I515553);
DFFARX1 I_22016 (I377144,I2859,I376700,I377170,);
nor I_22017 (I376680,I377170,I376726);
not I_22018 (I377192,I377170);
and I_22019 (I377209,I377192,I376726);
nor I_22020 (I376674,I376751,I377209);
nand I_22021 (I377240,I377192,I376802);
nor I_22022 (I376668,I377062,I377240);
nand I_22023 (I376671,I377192,I376980);
nand I_22024 (I377285,I376802,I515550);
nor I_22025 (I376683,I377045,I377285);
not I_22026 (I377346,I2866);
DFFARX1 I_22027 (I129315,I2859,I377346,I377372,);
DFFARX1 I_22028 (I129321,I2859,I377346,I377389,);
not I_22029 (I377397,I377389);
not I_22030 (I377414,I129342);
nor I_22031 (I377431,I377414,I129330);
not I_22032 (I377448,I129339);
nor I_22033 (I377465,I377431,I129324);
nor I_22034 (I377482,I377389,I377465);
DFFARX1 I_22035 (I377482,I2859,I377346,I377332,);
nor I_22036 (I377513,I129324,I129330);
nand I_22037 (I377530,I377513,I129342);
DFFARX1 I_22038 (I377530,I2859,I377346,I377335,);
nor I_22039 (I377561,I377448,I129324);
nand I_22040 (I377578,I377561,I129315);
nor I_22041 (I377595,I377372,I377578);
DFFARX1 I_22042 (I377595,I2859,I377346,I377311,);
not I_22043 (I377626,I377578);
nand I_22044 (I377323,I377389,I377626);
DFFARX1 I_22045 (I377578,I2859,I377346,I377666,);
not I_22046 (I377674,I377666);
not I_22047 (I377691,I129324);
not I_22048 (I377708,I129327);
nor I_22049 (I377725,I377708,I129339);
nor I_22050 (I377338,I377674,I377725);
nor I_22051 (I377756,I377708,I129336);
and I_22052 (I377773,I377756,I129318);
or I_22053 (I377790,I377773,I129333);
DFFARX1 I_22054 (I377790,I2859,I377346,I377816,);
nor I_22055 (I377326,I377816,I377372);
not I_22056 (I377838,I377816);
and I_22057 (I377855,I377838,I377372);
nor I_22058 (I377320,I377397,I377855);
nand I_22059 (I377886,I377838,I377448);
nor I_22060 (I377314,I377708,I377886);
nand I_22061 (I377317,I377838,I377626);
nand I_22062 (I377931,I377448,I129327);
nor I_22063 (I377329,I377691,I377931);
not I_22064 (I377992,I2866);
DFFARX1 I_22065 (I35883,I2859,I377992,I378018,);
DFFARX1 I_22066 (I35889,I2859,I377992,I378035,);
not I_22067 (I378043,I378035);
not I_22068 (I378060,I35907);
nor I_22069 (I378077,I378060,I35886);
not I_22070 (I378094,I35892);
nor I_22071 (I378111,I378077,I35898);
nor I_22072 (I378128,I378035,I378111);
DFFARX1 I_22073 (I378128,I2859,I377992,I377978,);
nor I_22074 (I378159,I35898,I35886);
nand I_22075 (I378176,I378159,I35907);
DFFARX1 I_22076 (I378176,I2859,I377992,I377981,);
nor I_22077 (I378207,I378094,I35898);
nand I_22078 (I378224,I378207,I35904);
nor I_22079 (I378241,I378018,I378224);
DFFARX1 I_22080 (I378241,I2859,I377992,I377957,);
not I_22081 (I378272,I378224);
nand I_22082 (I377969,I378035,I378272);
DFFARX1 I_22083 (I378224,I2859,I377992,I378312,);
not I_22084 (I378320,I378312);
not I_22085 (I378337,I35898);
not I_22086 (I378354,I35886);
nor I_22087 (I378371,I378354,I35892);
nor I_22088 (I377984,I378320,I378371);
nor I_22089 (I378402,I378354,I35895);
and I_22090 (I378419,I378402,I35883);
or I_22091 (I378436,I378419,I35901);
DFFARX1 I_22092 (I378436,I2859,I377992,I378462,);
nor I_22093 (I377972,I378462,I378018);
not I_22094 (I378484,I378462);
and I_22095 (I378501,I378484,I378018);
nor I_22096 (I377966,I378043,I378501);
nand I_22097 (I378532,I378484,I378094);
nor I_22098 (I377960,I378354,I378532);
nand I_22099 (I377963,I378484,I378272);
nand I_22100 (I378577,I378094,I35886);
nor I_22101 (I377975,I378337,I378577);
not I_22102 (I378638,I2866);
DFFARX1 I_22103 (I11641,I2859,I378638,I378664,);
DFFARX1 I_22104 (I11647,I2859,I378638,I378681,);
not I_22105 (I378689,I378681);
not I_22106 (I378706,I11641);
nor I_22107 (I378723,I378706,I11653);
not I_22108 (I378740,I11665);
nor I_22109 (I378757,I378723,I11659);
nor I_22110 (I378774,I378681,I378757);
DFFARX1 I_22111 (I378774,I2859,I378638,I378624,);
nor I_22112 (I378805,I11659,I11653);
nand I_22113 (I378822,I378805,I11641);
DFFARX1 I_22114 (I378822,I2859,I378638,I378627,);
nor I_22115 (I378853,I378740,I11659);
nand I_22116 (I378870,I378853,I11644);
nor I_22117 (I378887,I378664,I378870);
DFFARX1 I_22118 (I378887,I2859,I378638,I378603,);
not I_22119 (I378918,I378870);
nand I_22120 (I378615,I378681,I378918);
DFFARX1 I_22121 (I378870,I2859,I378638,I378958,);
not I_22122 (I378966,I378958);
not I_22123 (I378983,I11659);
not I_22124 (I379000,I11644);
nor I_22125 (I379017,I379000,I11665);
nor I_22126 (I378630,I378966,I379017);
nor I_22127 (I379048,I379000,I11662);
and I_22128 (I379065,I379048,I11656);
or I_22129 (I379082,I379065,I11650);
DFFARX1 I_22130 (I379082,I2859,I378638,I379108,);
nor I_22131 (I378618,I379108,I378664);
not I_22132 (I379130,I379108);
and I_22133 (I379147,I379130,I378664);
nor I_22134 (I378612,I378689,I379147);
nand I_22135 (I379178,I379130,I378740);
nor I_22136 (I378606,I379000,I379178);
nand I_22137 (I378609,I379130,I378918);
nand I_22138 (I379223,I378740,I11644);
nor I_22139 (I378621,I378983,I379223);
not I_22140 (I379284,I2866);
DFFARX1 I_22141 (I48531,I2859,I379284,I379310,);
DFFARX1 I_22142 (I48537,I2859,I379284,I379327,);
not I_22143 (I379335,I379327);
not I_22144 (I379352,I48555);
nor I_22145 (I379369,I379352,I48534);
not I_22146 (I379386,I48540);
nor I_22147 (I379403,I379369,I48546);
nor I_22148 (I379420,I379327,I379403);
DFFARX1 I_22149 (I379420,I2859,I379284,I379270,);
nor I_22150 (I379451,I48546,I48534);
nand I_22151 (I379468,I379451,I48555);
DFFARX1 I_22152 (I379468,I2859,I379284,I379273,);
nor I_22153 (I379499,I379386,I48546);
nand I_22154 (I379516,I379499,I48552);
nor I_22155 (I379533,I379310,I379516);
DFFARX1 I_22156 (I379533,I2859,I379284,I379249,);
not I_22157 (I379564,I379516);
nand I_22158 (I379261,I379327,I379564);
DFFARX1 I_22159 (I379516,I2859,I379284,I379604,);
not I_22160 (I379612,I379604);
not I_22161 (I379629,I48546);
not I_22162 (I379646,I48534);
nor I_22163 (I379663,I379646,I48540);
nor I_22164 (I379276,I379612,I379663);
nor I_22165 (I379694,I379646,I48543);
and I_22166 (I379711,I379694,I48531);
or I_22167 (I379728,I379711,I48549);
DFFARX1 I_22168 (I379728,I2859,I379284,I379754,);
nor I_22169 (I379264,I379754,I379310);
not I_22170 (I379776,I379754);
and I_22171 (I379793,I379776,I379310);
nor I_22172 (I379258,I379335,I379793);
nand I_22173 (I379824,I379776,I379386);
nor I_22174 (I379252,I379646,I379824);
nand I_22175 (I379255,I379776,I379564);
nand I_22176 (I379869,I379386,I48534);
nor I_22177 (I379267,I379629,I379869);
not I_22178 (I379930,I2866);
DFFARX1 I_22179 (I285126,I2859,I379930,I379956,);
DFFARX1 I_22180 (I285120,I2859,I379930,I379973,);
not I_22181 (I379981,I379973);
not I_22182 (I379998,I285135);
nor I_22183 (I380015,I379998,I285120);
not I_22184 (I380032,I285129);
nor I_22185 (I380049,I380015,I285138);
nor I_22186 (I380066,I379973,I380049);
DFFARX1 I_22187 (I380066,I2859,I379930,I379916,);
nor I_22188 (I380097,I285138,I285120);
nand I_22189 (I380114,I380097,I285135);
DFFARX1 I_22190 (I380114,I2859,I379930,I379919,);
nor I_22191 (I380145,I380032,I285138);
nand I_22192 (I380162,I380145,I285123);
nor I_22193 (I380179,I379956,I380162);
DFFARX1 I_22194 (I380179,I2859,I379930,I379895,);
not I_22195 (I380210,I380162);
nand I_22196 (I379907,I379973,I380210);
DFFARX1 I_22197 (I380162,I2859,I379930,I380250,);
not I_22198 (I380258,I380250);
not I_22199 (I380275,I285138);
not I_22200 (I380292,I285132);
nor I_22201 (I380309,I380292,I285129);
nor I_22202 (I379922,I380258,I380309);
nor I_22203 (I380340,I380292,I285141);
and I_22204 (I380357,I380340,I285144);
or I_22205 (I380374,I380357,I285123);
DFFARX1 I_22206 (I380374,I2859,I379930,I380400,);
nor I_22207 (I379910,I380400,I379956);
not I_22208 (I380422,I380400);
and I_22209 (I380439,I380422,I379956);
nor I_22210 (I379904,I379981,I380439);
nand I_22211 (I380470,I380422,I380032);
nor I_22212 (I379898,I380292,I380470);
nand I_22213 (I379901,I380422,I380210);
nand I_22214 (I380515,I380032,I285132);
nor I_22215 (I379913,I380275,I380515);
not I_22216 (I380576,I2866);
DFFARX1 I_22217 (I303044,I2859,I380576,I380602,);
DFFARX1 I_22218 (I303038,I2859,I380576,I380619,);
not I_22219 (I380627,I380619);
not I_22220 (I380644,I303053);
nor I_22221 (I380661,I380644,I303038);
not I_22222 (I380678,I303047);
nor I_22223 (I380695,I380661,I303056);
nor I_22224 (I380712,I380619,I380695);
DFFARX1 I_22225 (I380712,I2859,I380576,I380562,);
nor I_22226 (I380743,I303056,I303038);
nand I_22227 (I380760,I380743,I303053);
DFFARX1 I_22228 (I380760,I2859,I380576,I380565,);
nor I_22229 (I380791,I380678,I303056);
nand I_22230 (I380808,I380791,I303041);
nor I_22231 (I380825,I380602,I380808);
DFFARX1 I_22232 (I380825,I2859,I380576,I380541,);
not I_22233 (I380856,I380808);
nand I_22234 (I380553,I380619,I380856);
DFFARX1 I_22235 (I380808,I2859,I380576,I380896,);
not I_22236 (I380904,I380896);
not I_22237 (I380921,I303056);
not I_22238 (I380938,I303050);
nor I_22239 (I380955,I380938,I303047);
nor I_22240 (I380568,I380904,I380955);
nor I_22241 (I380986,I380938,I303059);
and I_22242 (I381003,I380986,I303062);
or I_22243 (I381020,I381003,I303041);
DFFARX1 I_22244 (I381020,I2859,I380576,I381046,);
nor I_22245 (I380556,I381046,I380602);
not I_22246 (I381068,I381046);
and I_22247 (I381085,I381068,I380602);
nor I_22248 (I380550,I380627,I381085);
nand I_22249 (I381116,I381068,I380678);
nor I_22250 (I380544,I380938,I381116);
nand I_22251 (I380547,I381068,I380856);
nand I_22252 (I381161,I380678,I303050);
nor I_22253 (I380559,I380921,I381161);
not I_22254 (I381222,I2866);
DFFARX1 I_22255 (I266630,I2859,I381222,I381248,);
DFFARX1 I_22256 (I266624,I2859,I381222,I381265,);
not I_22257 (I381273,I381265);
not I_22258 (I381290,I266639);
nor I_22259 (I381307,I381290,I266624);
not I_22260 (I381324,I266633);
nor I_22261 (I381341,I381307,I266642);
nor I_22262 (I381358,I381265,I381341);
DFFARX1 I_22263 (I381358,I2859,I381222,I381208,);
nor I_22264 (I381389,I266642,I266624);
nand I_22265 (I381406,I381389,I266639);
DFFARX1 I_22266 (I381406,I2859,I381222,I381211,);
nor I_22267 (I381437,I381324,I266642);
nand I_22268 (I381454,I381437,I266627);
nor I_22269 (I381471,I381248,I381454);
DFFARX1 I_22270 (I381471,I2859,I381222,I381187,);
not I_22271 (I381502,I381454);
nand I_22272 (I381199,I381265,I381502);
DFFARX1 I_22273 (I381454,I2859,I381222,I381542,);
not I_22274 (I381550,I381542);
not I_22275 (I381567,I266642);
not I_22276 (I381584,I266636);
nor I_22277 (I381601,I381584,I266633);
nor I_22278 (I381214,I381550,I381601);
nor I_22279 (I381632,I381584,I266645);
and I_22280 (I381649,I381632,I266648);
or I_22281 (I381666,I381649,I266627);
DFFARX1 I_22282 (I381666,I2859,I381222,I381692,);
nor I_22283 (I381202,I381692,I381248);
not I_22284 (I381714,I381692);
and I_22285 (I381731,I381714,I381248);
nor I_22286 (I381196,I381273,I381731);
nand I_22287 (I381762,I381714,I381324);
nor I_22288 (I381190,I381584,I381762);
nand I_22289 (I381193,I381714,I381502);
nand I_22290 (I381807,I381324,I266636);
nor I_22291 (I381205,I381567,I381807);
not I_22292 (I381868,I2866);
DFFARX1 I_22293 (I114559,I2859,I381868,I381894,);
DFFARX1 I_22294 (I114565,I2859,I381868,I381911,);
not I_22295 (I381919,I381911);
not I_22296 (I381936,I114586);
nor I_22297 (I381953,I381936,I114574);
not I_22298 (I381970,I114583);
nor I_22299 (I381987,I381953,I114568);
nor I_22300 (I382004,I381911,I381987);
DFFARX1 I_22301 (I382004,I2859,I381868,I381854,);
nor I_22302 (I382035,I114568,I114574);
nand I_22303 (I382052,I382035,I114586);
DFFARX1 I_22304 (I382052,I2859,I381868,I381857,);
nor I_22305 (I382083,I381970,I114568);
nand I_22306 (I382100,I382083,I114559);
nor I_22307 (I382117,I381894,I382100);
DFFARX1 I_22308 (I382117,I2859,I381868,I381833,);
not I_22309 (I382148,I382100);
nand I_22310 (I381845,I381911,I382148);
DFFARX1 I_22311 (I382100,I2859,I381868,I382188,);
not I_22312 (I382196,I382188);
not I_22313 (I382213,I114568);
not I_22314 (I382230,I114571);
nor I_22315 (I382247,I382230,I114583);
nor I_22316 (I381860,I382196,I382247);
nor I_22317 (I382278,I382230,I114580);
and I_22318 (I382295,I382278,I114562);
or I_22319 (I382312,I382295,I114577);
DFFARX1 I_22320 (I382312,I2859,I381868,I382338,);
nor I_22321 (I381848,I382338,I381894);
not I_22322 (I382360,I382338);
and I_22323 (I382377,I382360,I381894);
nor I_22324 (I381842,I381919,I382377);
nand I_22325 (I382408,I382360,I381970);
nor I_22326 (I381836,I382230,I382408);
nand I_22327 (I381839,I382360,I382148);
nand I_22328 (I382453,I381970,I114571);
nor I_22329 (I381851,I382213,I382453);
not I_22330 (I382514,I2866);
DFFARX1 I_22331 (I153557,I2859,I382514,I382540,);
DFFARX1 I_22332 (I153563,I2859,I382514,I382557,);
not I_22333 (I382565,I382557);
not I_22334 (I382582,I153584);
nor I_22335 (I382599,I382582,I153572);
not I_22336 (I382616,I153581);
nor I_22337 (I382633,I382599,I153566);
nor I_22338 (I382650,I382557,I382633);
DFFARX1 I_22339 (I382650,I2859,I382514,I382500,);
nor I_22340 (I382681,I153566,I153572);
nand I_22341 (I382698,I382681,I153584);
DFFARX1 I_22342 (I382698,I2859,I382514,I382503,);
nor I_22343 (I382729,I382616,I153566);
nand I_22344 (I382746,I382729,I153557);
nor I_22345 (I382763,I382540,I382746);
DFFARX1 I_22346 (I382763,I2859,I382514,I382479,);
not I_22347 (I382794,I382746);
nand I_22348 (I382491,I382557,I382794);
DFFARX1 I_22349 (I382746,I2859,I382514,I382834,);
not I_22350 (I382842,I382834);
not I_22351 (I382859,I153566);
not I_22352 (I382876,I153569);
nor I_22353 (I382893,I382876,I153581);
nor I_22354 (I382506,I382842,I382893);
nor I_22355 (I382924,I382876,I153578);
and I_22356 (I382941,I382924,I153560);
or I_22357 (I382958,I382941,I153575);
DFFARX1 I_22358 (I382958,I2859,I382514,I382984,);
nor I_22359 (I382494,I382984,I382540);
not I_22360 (I383006,I382984);
and I_22361 (I383023,I383006,I382540);
nor I_22362 (I382488,I382565,I383023);
nand I_22363 (I383054,I383006,I382616);
nor I_22364 (I382482,I382876,I383054);
nand I_22365 (I382485,I383006,I382794);
nand I_22366 (I383099,I382616,I153569);
nor I_22367 (I382497,I382859,I383099);
not I_22368 (I383160,I2866);
DFFARX1 I_22369 (I300154,I2859,I383160,I383186,);
DFFARX1 I_22370 (I300148,I2859,I383160,I383203,);
not I_22371 (I383211,I383203);
not I_22372 (I383228,I300163);
nor I_22373 (I383245,I383228,I300148);
not I_22374 (I383262,I300157);
nor I_22375 (I383279,I383245,I300166);
nor I_22376 (I383296,I383203,I383279);
DFFARX1 I_22377 (I383296,I2859,I383160,I383146,);
nor I_22378 (I383327,I300166,I300148);
nand I_22379 (I383344,I383327,I300163);
DFFARX1 I_22380 (I383344,I2859,I383160,I383149,);
nor I_22381 (I383375,I383262,I300166);
nand I_22382 (I383392,I383375,I300151);
nor I_22383 (I383409,I383186,I383392);
DFFARX1 I_22384 (I383409,I2859,I383160,I383125,);
not I_22385 (I383440,I383392);
nand I_22386 (I383137,I383203,I383440);
DFFARX1 I_22387 (I383392,I2859,I383160,I383480,);
not I_22388 (I383488,I383480);
not I_22389 (I383505,I300166);
not I_22390 (I383522,I300160);
nor I_22391 (I383539,I383522,I300157);
nor I_22392 (I383152,I383488,I383539);
nor I_22393 (I383570,I383522,I300169);
and I_22394 (I383587,I383570,I300172);
or I_22395 (I383604,I383587,I300151);
DFFARX1 I_22396 (I383604,I2859,I383160,I383630,);
nor I_22397 (I383140,I383630,I383186);
not I_22398 (I383652,I383630);
and I_22399 (I383669,I383652,I383186);
nor I_22400 (I383134,I383211,I383669);
nand I_22401 (I383700,I383652,I383262);
nor I_22402 (I383128,I383522,I383700);
nand I_22403 (I383131,I383652,I383440);
nand I_22404 (I383745,I383262,I300160);
nor I_22405 (I383143,I383505,I383745);
not I_22406 (I383806,I2866);
DFFARX1 I_22407 (I2132,I2859,I383806,I383832,);
DFFARX1 I_22408 (I1988,I2859,I383806,I383849,);
not I_22409 (I383857,I383849);
not I_22410 (I383874,I2180);
nor I_22411 (I383891,I383874,I2172);
not I_22412 (I383908,I2508);
nor I_22413 (I383925,I383891,I2484);
nor I_22414 (I383942,I383849,I383925);
DFFARX1 I_22415 (I383942,I2859,I383806,I383792,);
nor I_22416 (I383973,I2484,I2172);
nand I_22417 (I383990,I383973,I2180);
DFFARX1 I_22418 (I383990,I2859,I383806,I383795,);
nor I_22419 (I384021,I383908,I2484);
nand I_22420 (I384038,I384021,I2692);
nor I_22421 (I384055,I383832,I384038);
DFFARX1 I_22422 (I384055,I2859,I383806,I383771,);
not I_22423 (I384086,I384038);
nand I_22424 (I383783,I383849,I384086);
DFFARX1 I_22425 (I384038,I2859,I383806,I384126,);
not I_22426 (I384134,I384126);
not I_22427 (I384151,I2484);
not I_22428 (I384168,I2644);
nor I_22429 (I384185,I384168,I2508);
nor I_22430 (I383798,I384134,I384185);
nor I_22431 (I384216,I384168,I2068);
and I_22432 (I384233,I384216,I2276);
or I_22433 (I384250,I384233,I1740);
DFFARX1 I_22434 (I384250,I2859,I383806,I384276,);
nor I_22435 (I383786,I384276,I383832);
not I_22436 (I384298,I384276);
and I_22437 (I384315,I384298,I383832);
nor I_22438 (I383780,I383857,I384315);
nand I_22439 (I384346,I384298,I383908);
nor I_22440 (I383774,I384168,I384346);
nand I_22441 (I383777,I384298,I384086);
nand I_22442 (I384391,I383908,I2644);
nor I_22443 (I383789,I384151,I384391);
not I_22444 (I384452,I2866);
DFFARX1 I_22445 (I440654,I2859,I384452,I384478,);
DFFARX1 I_22446 (I440636,I2859,I384452,I384495,);
not I_22447 (I384503,I384495);
not I_22448 (I384520,I440645);
nor I_22449 (I384537,I384520,I440657);
not I_22450 (I384554,I440639);
nor I_22451 (I384571,I384537,I440648);
nor I_22452 (I384588,I384495,I384571);
DFFARX1 I_22453 (I384588,I2859,I384452,I384438,);
nor I_22454 (I384619,I440648,I440657);
nand I_22455 (I384636,I384619,I440645);
DFFARX1 I_22456 (I384636,I2859,I384452,I384441,);
nor I_22457 (I384667,I384554,I440648);
nand I_22458 (I384684,I384667,I440660);
nor I_22459 (I384701,I384478,I384684);
DFFARX1 I_22460 (I384701,I2859,I384452,I384417,);
not I_22461 (I384732,I384684);
nand I_22462 (I384429,I384495,I384732);
DFFARX1 I_22463 (I384684,I2859,I384452,I384772,);
not I_22464 (I384780,I384772);
not I_22465 (I384797,I440648);
not I_22466 (I384814,I440636);
nor I_22467 (I384831,I384814,I440639);
nor I_22468 (I384444,I384780,I384831);
nor I_22469 (I384862,I384814,I440642);
and I_22470 (I384879,I384862,I440651);
or I_22471 (I384896,I384879,I440639);
DFFARX1 I_22472 (I384896,I2859,I384452,I384922,);
nor I_22473 (I384432,I384922,I384478);
not I_22474 (I384944,I384922);
and I_22475 (I384961,I384944,I384478);
nor I_22476 (I384426,I384503,I384961);
nand I_22477 (I384992,I384944,I384554);
nor I_22478 (I384420,I384814,I384992);
nand I_22479 (I384423,I384944,I384732);
nand I_22480 (I385037,I384554,I440636);
nor I_22481 (I384435,I384797,I385037);
not I_22482 (I385098,I2866);
DFFARX1 I_22483 (I463774,I2859,I385098,I385124,);
DFFARX1 I_22484 (I463756,I2859,I385098,I385141,);
not I_22485 (I385149,I385141);
not I_22486 (I385166,I463765);
nor I_22487 (I385183,I385166,I463777);
not I_22488 (I385200,I463759);
nor I_22489 (I385217,I385183,I463768);
nor I_22490 (I385234,I385141,I385217);
DFFARX1 I_22491 (I385234,I2859,I385098,I385084,);
nor I_22492 (I385265,I463768,I463777);
nand I_22493 (I385282,I385265,I463765);
DFFARX1 I_22494 (I385282,I2859,I385098,I385087,);
nor I_22495 (I385313,I385200,I463768);
nand I_22496 (I385330,I385313,I463780);
nor I_22497 (I385347,I385124,I385330);
DFFARX1 I_22498 (I385347,I2859,I385098,I385063,);
not I_22499 (I385378,I385330);
nand I_22500 (I385075,I385141,I385378);
DFFARX1 I_22501 (I385330,I2859,I385098,I385418,);
not I_22502 (I385426,I385418);
not I_22503 (I385443,I463768);
not I_22504 (I385460,I463756);
nor I_22505 (I385477,I385460,I463759);
nor I_22506 (I385090,I385426,I385477);
nor I_22507 (I385508,I385460,I463762);
and I_22508 (I385525,I385508,I463771);
or I_22509 (I385542,I385525,I463759);
DFFARX1 I_22510 (I385542,I2859,I385098,I385568,);
nor I_22511 (I385078,I385568,I385124);
not I_22512 (I385590,I385568);
and I_22513 (I385607,I385590,I385124);
nor I_22514 (I385072,I385149,I385607);
nand I_22515 (I385638,I385590,I385200);
nor I_22516 (I385066,I385460,I385638);
nand I_22517 (I385069,I385590,I385378);
nand I_22518 (I385683,I385200,I463756);
nor I_22519 (I385081,I385443,I385683);
not I_22520 (I385744,I2866);
DFFARX1 I_22521 (I138274,I2859,I385744,I385770,);
DFFARX1 I_22522 (I138280,I2859,I385744,I385787,);
not I_22523 (I385795,I385787);
not I_22524 (I385812,I138301);
nor I_22525 (I385829,I385812,I138289);
not I_22526 (I385846,I138298);
nor I_22527 (I385863,I385829,I138283);
nor I_22528 (I385880,I385787,I385863);
DFFARX1 I_22529 (I385880,I2859,I385744,I385730,);
nor I_22530 (I385911,I138283,I138289);
nand I_22531 (I385928,I385911,I138301);
DFFARX1 I_22532 (I385928,I2859,I385744,I385733,);
nor I_22533 (I385959,I385846,I138283);
nand I_22534 (I385976,I385959,I138274);
nor I_22535 (I385993,I385770,I385976);
DFFARX1 I_22536 (I385993,I2859,I385744,I385709,);
not I_22537 (I386024,I385976);
nand I_22538 (I385721,I385787,I386024);
DFFARX1 I_22539 (I385976,I2859,I385744,I386064,);
not I_22540 (I386072,I386064);
not I_22541 (I386089,I138283);
not I_22542 (I386106,I138286);
nor I_22543 (I386123,I386106,I138298);
nor I_22544 (I385736,I386072,I386123);
nor I_22545 (I386154,I386106,I138295);
and I_22546 (I386171,I386154,I138277);
or I_22547 (I386188,I386171,I138292);
DFFARX1 I_22548 (I386188,I2859,I385744,I386214,);
nor I_22549 (I385724,I386214,I385770);
not I_22550 (I386236,I386214);
and I_22551 (I386253,I386236,I385770);
nor I_22552 (I385718,I385795,I386253);
nand I_22553 (I386284,I386236,I385846);
nor I_22554 (I385712,I386106,I386284);
nand I_22555 (I385715,I386236,I386024);
nand I_22556 (I386329,I385846,I138286);
nor I_22557 (I385727,I386089,I386329);
not I_22558 (I386390,I2866);
DFFARX1 I_22559 (I484582,I2859,I386390,I386416,);
DFFARX1 I_22560 (I484564,I2859,I386390,I386433,);
not I_22561 (I386441,I386433);
not I_22562 (I386458,I484573);
nor I_22563 (I386475,I386458,I484585);
not I_22564 (I386492,I484567);
nor I_22565 (I386509,I386475,I484576);
nor I_22566 (I386526,I386433,I386509);
DFFARX1 I_22567 (I386526,I2859,I386390,I386376,);
nor I_22568 (I386557,I484576,I484585);
nand I_22569 (I386574,I386557,I484573);
DFFARX1 I_22570 (I386574,I2859,I386390,I386379,);
nor I_22571 (I386605,I386492,I484576);
nand I_22572 (I386622,I386605,I484588);
nor I_22573 (I386639,I386416,I386622);
DFFARX1 I_22574 (I386639,I2859,I386390,I386355,);
not I_22575 (I386670,I386622);
nand I_22576 (I386367,I386433,I386670);
DFFARX1 I_22577 (I386622,I2859,I386390,I386710,);
not I_22578 (I386718,I386710);
not I_22579 (I386735,I484576);
not I_22580 (I386752,I484564);
nor I_22581 (I386769,I386752,I484567);
nor I_22582 (I386382,I386718,I386769);
nor I_22583 (I386800,I386752,I484570);
and I_22584 (I386817,I386800,I484579);
or I_22585 (I386834,I386817,I484567);
DFFARX1 I_22586 (I386834,I2859,I386390,I386860,);
nor I_22587 (I386370,I386860,I386416);
not I_22588 (I386882,I386860);
and I_22589 (I386899,I386882,I386416);
nor I_22590 (I386364,I386441,I386899);
nand I_22591 (I386930,I386882,I386492);
nor I_22592 (I386358,I386752,I386930);
nand I_22593 (I386361,I386882,I386670);
nand I_22594 (I386975,I386492,I484564);
nor I_22595 (I386373,I386735,I386975);
not I_22596 (I387036,I2866);
DFFARX1 I_22597 (I1412,I2859,I387036,I387062,);
DFFARX1 I_22598 (I2788,I2859,I387036,I387079,);
not I_22599 (I387087,I387079);
not I_22600 (I387104,I1524);
nor I_22601 (I387121,I387104,I2092);
not I_22602 (I387138,I1764);
nor I_22603 (I387155,I387121,I1812);
nor I_22604 (I387172,I387079,I387155);
DFFARX1 I_22605 (I387172,I2859,I387036,I387022,);
nor I_22606 (I387203,I1812,I2092);
nand I_22607 (I387220,I387203,I1524);
DFFARX1 I_22608 (I387220,I2859,I387036,I387025,);
nor I_22609 (I387251,I387138,I1812);
nand I_22610 (I387268,I387251,I2332);
nor I_22611 (I387285,I387062,I387268);
DFFARX1 I_22612 (I387285,I2859,I387036,I387001,);
not I_22613 (I387316,I387268);
nand I_22614 (I387013,I387079,I387316);
DFFARX1 I_22615 (I387268,I2859,I387036,I387356,);
not I_22616 (I387364,I387356);
not I_22617 (I387381,I1812);
not I_22618 (I387398,I1732);
nor I_22619 (I387415,I387398,I1764);
nor I_22620 (I387028,I387364,I387415);
nor I_22621 (I387446,I387398,I2556);
and I_22622 (I387463,I387446,I2188);
or I_22623 (I387480,I387463,I1588);
DFFARX1 I_22624 (I387480,I2859,I387036,I387506,);
nor I_22625 (I387016,I387506,I387062);
not I_22626 (I387528,I387506);
and I_22627 (I387545,I387528,I387062);
nor I_22628 (I387010,I387087,I387545);
nand I_22629 (I387576,I387528,I387138);
nor I_22630 (I387004,I387398,I387576);
nand I_22631 (I387007,I387528,I387316);
nand I_22632 (I387621,I387138,I1732);
nor I_22633 (I387019,I387381,I387621);
not I_22634 (I387682,I2866);
DFFARX1 I_22635 (I68563,I2859,I387682,I387708,);
DFFARX1 I_22636 (I68575,I2859,I387682,I387725,);
not I_22637 (I387733,I387725);
not I_22638 (I387750,I68581);
nor I_22639 (I387767,I387750,I68566);
not I_22640 (I387784,I68557);
nor I_22641 (I387801,I387767,I68578);
nor I_22642 (I387818,I387725,I387801);
DFFARX1 I_22643 (I387818,I2859,I387682,I387668,);
nor I_22644 (I387849,I68578,I68566);
nand I_22645 (I387866,I387849,I68581);
DFFARX1 I_22646 (I387866,I2859,I387682,I387671,);
nor I_22647 (I387897,I387784,I68578);
nand I_22648 (I387914,I387897,I68560);
nor I_22649 (I387931,I387708,I387914);
DFFARX1 I_22650 (I387931,I2859,I387682,I387647,);
not I_22651 (I387962,I387914);
nand I_22652 (I387659,I387725,I387962);
DFFARX1 I_22653 (I387914,I2859,I387682,I388002,);
not I_22654 (I388010,I388002);
not I_22655 (I388027,I68578);
not I_22656 (I388044,I68569);
nor I_22657 (I388061,I388044,I68557);
nor I_22658 (I387674,I388010,I388061);
nor I_22659 (I388092,I388044,I68572);
and I_22660 (I388109,I388092,I68560);
or I_22661 (I388126,I388109,I68557);
DFFARX1 I_22662 (I388126,I2859,I387682,I388152,);
nor I_22663 (I387662,I388152,I387708);
not I_22664 (I388174,I388152);
and I_22665 (I388191,I388174,I387708);
nor I_22666 (I387656,I387733,I388191);
nand I_22667 (I388222,I388174,I387784);
nor I_22668 (I387650,I388044,I388222);
nand I_22669 (I387653,I388174,I387962);
nand I_22670 (I388267,I387784,I68569);
nor I_22671 (I387665,I388027,I388267);
not I_22672 (I388328,I2866);
DFFARX1 I_22673 (I489206,I2859,I388328,I388354,);
DFFARX1 I_22674 (I489188,I2859,I388328,I388371,);
not I_22675 (I388379,I388371);
not I_22676 (I388396,I489197);
nor I_22677 (I388413,I388396,I489209);
not I_22678 (I388430,I489191);
nor I_22679 (I388447,I388413,I489200);
nor I_22680 (I388464,I388371,I388447);
DFFARX1 I_22681 (I388464,I2859,I388328,I388314,);
nor I_22682 (I388495,I489200,I489209);
nand I_22683 (I388512,I388495,I489197);
DFFARX1 I_22684 (I388512,I2859,I388328,I388317,);
nor I_22685 (I388543,I388430,I489200);
nand I_22686 (I388560,I388543,I489212);
nor I_22687 (I388577,I388354,I388560);
DFFARX1 I_22688 (I388577,I2859,I388328,I388293,);
not I_22689 (I388608,I388560);
nand I_22690 (I388305,I388371,I388608);
DFFARX1 I_22691 (I388560,I2859,I388328,I388648,);
not I_22692 (I388656,I388648);
not I_22693 (I388673,I489200);
not I_22694 (I388690,I489188);
nor I_22695 (I388707,I388690,I489191);
nor I_22696 (I388320,I388656,I388707);
nor I_22697 (I388738,I388690,I489194);
and I_22698 (I388755,I388738,I489203);
or I_22699 (I388772,I388755,I489191);
DFFARX1 I_22700 (I388772,I2859,I388328,I388798,);
nor I_22701 (I388308,I388798,I388354);
not I_22702 (I388820,I388798);
and I_22703 (I388837,I388820,I388354);
nor I_22704 (I388302,I388379,I388837);
nand I_22705 (I388868,I388820,I388430);
nor I_22706 (I388296,I388690,I388868);
nand I_22707 (I388299,I388820,I388608);
nand I_22708 (I388913,I388430,I489188);
nor I_22709 (I388311,I388673,I388913);
not I_22710 (I388974,I2866);
DFFARX1 I_22711 (I42207,I2859,I388974,I389000,);
DFFARX1 I_22712 (I42213,I2859,I388974,I389017,);
not I_22713 (I389025,I389017);
not I_22714 (I389042,I42231);
nor I_22715 (I389059,I389042,I42210);
not I_22716 (I389076,I42216);
nor I_22717 (I389093,I389059,I42222);
nor I_22718 (I389110,I389017,I389093);
DFFARX1 I_22719 (I389110,I2859,I388974,I388960,);
nor I_22720 (I389141,I42222,I42210);
nand I_22721 (I389158,I389141,I42231);
DFFARX1 I_22722 (I389158,I2859,I388974,I388963,);
nor I_22723 (I389189,I389076,I42222);
nand I_22724 (I389206,I389189,I42228);
nor I_22725 (I389223,I389000,I389206);
DFFARX1 I_22726 (I389223,I2859,I388974,I388939,);
not I_22727 (I389254,I389206);
nand I_22728 (I388951,I389017,I389254);
DFFARX1 I_22729 (I389206,I2859,I388974,I389294,);
not I_22730 (I389302,I389294);
not I_22731 (I389319,I42222);
not I_22732 (I389336,I42210);
nor I_22733 (I389353,I389336,I42216);
nor I_22734 (I388966,I389302,I389353);
nor I_22735 (I389384,I389336,I42219);
and I_22736 (I389401,I389384,I42207);
or I_22737 (I389418,I389401,I42225);
DFFARX1 I_22738 (I389418,I2859,I388974,I389444,);
nor I_22739 (I388954,I389444,I389000);
not I_22740 (I389466,I389444);
and I_22741 (I389483,I389466,I389000);
nor I_22742 (I388948,I389025,I389483);
nand I_22743 (I389514,I389466,I389076);
nor I_22744 (I388942,I389336,I389514);
nand I_22745 (I388945,I389466,I389254);
nand I_22746 (I389559,I389076,I42210);
nor I_22747 (I388957,I389319,I389559);
not I_22748 (I389620,I2866);
DFFARX1 I_22749 (I554060,I2859,I389620,I389646,);
DFFARX1 I_22750 (I554084,I2859,I389620,I389663,);
not I_22751 (I389671,I389663);
not I_22752 (I389688,I554066);
nor I_22753 (I389705,I389688,I554075);
not I_22754 (I389722,I554060);
nor I_22755 (I389739,I389705,I554081);
nor I_22756 (I389756,I389663,I389739);
DFFARX1 I_22757 (I389756,I2859,I389620,I389606,);
nor I_22758 (I389787,I554081,I554075);
nand I_22759 (I389804,I389787,I554066);
DFFARX1 I_22760 (I389804,I2859,I389620,I389609,);
nor I_22761 (I389835,I389722,I554081);
nand I_22762 (I389852,I389835,I554078);
nor I_22763 (I389869,I389646,I389852);
DFFARX1 I_22764 (I389869,I2859,I389620,I389585,);
not I_22765 (I389900,I389852);
nand I_22766 (I389597,I389663,I389900);
DFFARX1 I_22767 (I389852,I2859,I389620,I389940,);
not I_22768 (I389948,I389940);
not I_22769 (I389965,I554081);
not I_22770 (I389982,I554072);
nor I_22771 (I389999,I389982,I554060);
nor I_22772 (I389612,I389948,I389999);
nor I_22773 (I390030,I389982,I554063);
and I_22774 (I390047,I390030,I554087);
or I_22775 (I390064,I390047,I554069);
DFFARX1 I_22776 (I390064,I2859,I389620,I390090,);
nor I_22777 (I389600,I390090,I389646);
not I_22778 (I390112,I390090);
and I_22779 (I390129,I390112,I389646);
nor I_22780 (I389594,I389671,I390129);
nand I_22781 (I390160,I390112,I389722);
nor I_22782 (I389588,I389982,I390160);
nand I_22783 (I389591,I390112,I389900);
nand I_22784 (I390205,I389722,I554072);
nor I_22785 (I389603,I389965,I390205);
not I_22786 (I390266,I2866);
DFFARX1 I_22787 (I230213,I2859,I390266,I390292,);
DFFARX1 I_22788 (I230225,I2859,I390266,I390309,);
not I_22789 (I390317,I390309);
not I_22790 (I390334,I230234);
nor I_22791 (I390351,I390334,I230210);
not I_22792 (I390368,I230228);
nor I_22793 (I390385,I390351,I230222);
nor I_22794 (I390402,I390309,I390385);
DFFARX1 I_22795 (I390402,I2859,I390266,I390252,);
nor I_22796 (I390433,I230222,I230210);
nand I_22797 (I390450,I390433,I230234);
DFFARX1 I_22798 (I390450,I2859,I390266,I390255,);
nor I_22799 (I390481,I390368,I230222);
nand I_22800 (I390498,I390481,I230216);
nor I_22801 (I390515,I390292,I390498);
DFFARX1 I_22802 (I390515,I2859,I390266,I390231,);
not I_22803 (I390546,I390498);
nand I_22804 (I390243,I390309,I390546);
DFFARX1 I_22805 (I390498,I2859,I390266,I390586,);
not I_22806 (I390594,I390586);
not I_22807 (I390611,I230222);
not I_22808 (I390628,I230231);
nor I_22809 (I390645,I390628,I230228);
nor I_22810 (I390258,I390594,I390645);
nor I_22811 (I390676,I390628,I230213);
and I_22812 (I390693,I390676,I230210);
or I_22813 (I390710,I390693,I230219);
DFFARX1 I_22814 (I390710,I2859,I390266,I390736,);
nor I_22815 (I390246,I390736,I390292);
not I_22816 (I390758,I390736);
and I_22817 (I390775,I390758,I390292);
nor I_22818 (I390240,I390317,I390775);
nand I_22819 (I390806,I390758,I390368);
nor I_22820 (I390234,I390628,I390806);
nand I_22821 (I390237,I390758,I390546);
nand I_22822 (I390851,I390368,I230231);
nor I_22823 (I390249,I390611,I390851);
not I_22824 (I390912,I2866);
DFFARX1 I_22825 (I504676,I2859,I390912,I390938,);
DFFARX1 I_22826 (I504682,I2859,I390912,I390955,);
not I_22827 (I390963,I390955);
not I_22828 (I390980,I504679);
nor I_22829 (I390997,I390980,I504658);
not I_22830 (I391014,I504661);
nor I_22831 (I391031,I390997,I504667);
nor I_22832 (I391048,I390955,I391031);
DFFARX1 I_22833 (I391048,I2859,I390912,I390898,);
nor I_22834 (I391079,I504667,I504658);
nand I_22835 (I391096,I391079,I504679);
DFFARX1 I_22836 (I391096,I2859,I390912,I390901,);
nor I_22837 (I391127,I391014,I504667);
nand I_22838 (I391144,I391127,I504661);
nor I_22839 (I391161,I390938,I391144);
DFFARX1 I_22840 (I391161,I2859,I390912,I390877,);
not I_22841 (I391192,I391144);
nand I_22842 (I390889,I390955,I391192);
DFFARX1 I_22843 (I391144,I2859,I390912,I391232,);
not I_22844 (I391240,I391232);
not I_22845 (I391257,I504667);
not I_22846 (I391274,I504670);
nor I_22847 (I391291,I391274,I504661);
nor I_22848 (I390904,I391240,I391291);
nor I_22849 (I391322,I391274,I504658);
and I_22850 (I391339,I391322,I504664);
or I_22851 (I391356,I391339,I504673);
DFFARX1 I_22852 (I391356,I2859,I390912,I391382,);
nor I_22853 (I390892,I391382,I390938);
not I_22854 (I391404,I391382);
and I_22855 (I391421,I391404,I390938);
nor I_22856 (I390886,I390963,I391421);
nand I_22857 (I391452,I391404,I391014);
nor I_22858 (I390880,I391274,I391452);
nand I_22859 (I390883,I391404,I391192);
nand I_22860 (I391497,I391014,I504670);
nor I_22861 (I390895,I391257,I391497);
not I_22862 (I391558,I2866);
DFFARX1 I_22863 (I143544,I2859,I391558,I391584,);
DFFARX1 I_22864 (I143550,I2859,I391558,I391601,);
not I_22865 (I391609,I391601);
not I_22866 (I391626,I143571);
nor I_22867 (I391643,I391626,I143559);
not I_22868 (I391660,I143568);
nor I_22869 (I391677,I391643,I143553);
nor I_22870 (I391694,I391601,I391677);
DFFARX1 I_22871 (I391694,I2859,I391558,I391544,);
nor I_22872 (I391725,I143553,I143559);
nand I_22873 (I391742,I391725,I143571);
DFFARX1 I_22874 (I391742,I2859,I391558,I391547,);
nor I_22875 (I391773,I391660,I143553);
nand I_22876 (I391790,I391773,I143544);
nor I_22877 (I391807,I391584,I391790);
DFFARX1 I_22878 (I391807,I2859,I391558,I391523,);
not I_22879 (I391838,I391790);
nand I_22880 (I391535,I391601,I391838);
DFFARX1 I_22881 (I391790,I2859,I391558,I391878,);
not I_22882 (I391886,I391878);
not I_22883 (I391903,I143553);
not I_22884 (I391920,I143556);
nor I_22885 (I391937,I391920,I143568);
nor I_22886 (I391550,I391886,I391937);
nor I_22887 (I391968,I391920,I143565);
and I_22888 (I391985,I391968,I143547);
or I_22889 (I392002,I391985,I143562);
DFFARX1 I_22890 (I392002,I2859,I391558,I392028,);
nor I_22891 (I391538,I392028,I391584);
not I_22892 (I392050,I392028);
and I_22893 (I392067,I392050,I391584);
nor I_22894 (I391532,I391609,I392067);
nand I_22895 (I392098,I392050,I391660);
nor I_22896 (I391526,I391920,I392098);
nand I_22897 (I391529,I392050,I391838);
nand I_22898 (I392143,I391660,I143556);
nor I_22899 (I391541,I391903,I392143);
not I_22900 (I392204,I2866);
DFFARX1 I_22901 (I17965,I2859,I392204,I392230,);
DFFARX1 I_22902 (I17971,I2859,I392204,I392247,);
not I_22903 (I392255,I392247);
not I_22904 (I392272,I17965);
nor I_22905 (I392289,I392272,I17977);
not I_22906 (I392306,I17989);
nor I_22907 (I392323,I392289,I17983);
nor I_22908 (I392340,I392247,I392323);
DFFARX1 I_22909 (I392340,I2859,I392204,I392190,);
nor I_22910 (I392371,I17983,I17977);
nand I_22911 (I392388,I392371,I17965);
DFFARX1 I_22912 (I392388,I2859,I392204,I392193,);
nor I_22913 (I392419,I392306,I17983);
nand I_22914 (I392436,I392419,I17968);
nor I_22915 (I392453,I392230,I392436);
DFFARX1 I_22916 (I392453,I2859,I392204,I392169,);
not I_22917 (I392484,I392436);
nand I_22918 (I392181,I392247,I392484);
DFFARX1 I_22919 (I392436,I2859,I392204,I392524,);
not I_22920 (I392532,I392524);
not I_22921 (I392549,I17983);
not I_22922 (I392566,I17968);
nor I_22923 (I392583,I392566,I17989);
nor I_22924 (I392196,I392532,I392583);
nor I_22925 (I392614,I392566,I17986);
and I_22926 (I392631,I392614,I17980);
or I_22927 (I392648,I392631,I17974);
DFFARX1 I_22928 (I392648,I2859,I392204,I392674,);
nor I_22929 (I392184,I392674,I392230);
not I_22930 (I392696,I392674);
and I_22931 (I392713,I392696,I392230);
nor I_22932 (I392178,I392255,I392713);
nand I_22933 (I392744,I392696,I392306);
nor I_22934 (I392172,I392566,I392744);
nand I_22935 (I392175,I392696,I392484);
nand I_22936 (I392789,I392306,I17968);
nor I_22937 (I392187,I392549,I392789);
not I_22938 (I392850,I2866);
DFFARX1 I_22939 (I346003,I2859,I392850,I392876,);
DFFARX1 I_22940 (I346000,I2859,I392850,I392893,);
not I_22941 (I392901,I392893);
not I_22942 (I392918,I346000);
nor I_22943 (I392935,I392918,I346003);
not I_22944 (I392952,I346015);
nor I_22945 (I392969,I392935,I346009);
nor I_22946 (I392986,I392893,I392969);
DFFARX1 I_22947 (I392986,I2859,I392850,I392836,);
nor I_22948 (I393017,I346009,I346003);
nand I_22949 (I393034,I393017,I346000);
DFFARX1 I_22950 (I393034,I2859,I392850,I392839,);
nor I_22951 (I393065,I392952,I346009);
nand I_22952 (I393082,I393065,I345997);
nor I_22953 (I393099,I392876,I393082);
DFFARX1 I_22954 (I393099,I2859,I392850,I392815,);
not I_22955 (I393130,I393082);
nand I_22956 (I392827,I392893,I393130);
DFFARX1 I_22957 (I393082,I2859,I392850,I393170,);
not I_22958 (I393178,I393170);
not I_22959 (I393195,I346009);
not I_22960 (I393212,I346006);
nor I_22961 (I393229,I393212,I346015);
nor I_22962 (I392842,I393178,I393229);
nor I_22963 (I393260,I393212,I346012);
and I_22964 (I393277,I393260,I346018);
or I_22965 (I393294,I393277,I345997);
DFFARX1 I_22966 (I393294,I2859,I392850,I393320,);
nor I_22967 (I392830,I393320,I392876);
not I_22968 (I393342,I393320);
and I_22969 (I393359,I393342,I392876);
nor I_22970 (I392824,I392901,I393359);
nand I_22971 (I393390,I393342,I392952);
nor I_22972 (I392818,I393212,I393390);
nand I_22973 (I392821,I393342,I393130);
nand I_22974 (I393435,I392952,I346006);
nor I_22975 (I392833,I393195,I393435);
not I_22976 (I393496,I2866);
DFFARX1 I_22977 (I301888,I2859,I393496,I393522,);
DFFARX1 I_22978 (I301882,I2859,I393496,I393539,);
not I_22979 (I393547,I393539);
not I_22980 (I393564,I301897);
nor I_22981 (I393581,I393564,I301882);
not I_22982 (I393598,I301891);
nor I_22983 (I393615,I393581,I301900);
nor I_22984 (I393632,I393539,I393615);
DFFARX1 I_22985 (I393632,I2859,I393496,I393482,);
nor I_22986 (I393663,I301900,I301882);
nand I_22987 (I393680,I393663,I301897);
DFFARX1 I_22988 (I393680,I2859,I393496,I393485,);
nor I_22989 (I393711,I393598,I301900);
nand I_22990 (I393728,I393711,I301885);
nor I_22991 (I393745,I393522,I393728);
DFFARX1 I_22992 (I393745,I2859,I393496,I393461,);
not I_22993 (I393776,I393728);
nand I_22994 (I393473,I393539,I393776);
DFFARX1 I_22995 (I393728,I2859,I393496,I393816,);
not I_22996 (I393824,I393816);
not I_22997 (I393841,I301900);
not I_22998 (I393858,I301894);
nor I_22999 (I393875,I393858,I301891);
nor I_23000 (I393488,I393824,I393875);
nor I_23001 (I393906,I393858,I301903);
and I_23002 (I393923,I393906,I301906);
or I_23003 (I393940,I393923,I301885);
DFFARX1 I_23004 (I393940,I2859,I393496,I393966,);
nor I_23005 (I393476,I393966,I393522);
not I_23006 (I393988,I393966);
and I_23007 (I394005,I393988,I393522);
nor I_23008 (I393470,I393547,I394005);
nand I_23009 (I394036,I393988,I393598);
nor I_23010 (I393464,I393858,I394036);
nand I_23011 (I393467,I393988,I393776);
nand I_23012 (I394081,I393598,I301894);
nor I_23013 (I393479,I393841,I394081);
not I_23014 (I394142,I2866);
DFFARX1 I_23015 (I258538,I2859,I394142,I394168,);
DFFARX1 I_23016 (I258532,I2859,I394142,I394185,);
not I_23017 (I394193,I394185);
not I_23018 (I394210,I258547);
nor I_23019 (I394227,I394210,I258532);
not I_23020 (I394244,I258541);
nor I_23021 (I394261,I394227,I258550);
nor I_23022 (I394278,I394185,I394261);
DFFARX1 I_23023 (I394278,I2859,I394142,I394128,);
nor I_23024 (I394309,I258550,I258532);
nand I_23025 (I394326,I394309,I258547);
DFFARX1 I_23026 (I394326,I2859,I394142,I394131,);
nor I_23027 (I394357,I394244,I258550);
nand I_23028 (I394374,I394357,I258535);
nor I_23029 (I394391,I394168,I394374);
DFFARX1 I_23030 (I394391,I2859,I394142,I394107,);
not I_23031 (I394422,I394374);
nand I_23032 (I394119,I394185,I394422);
DFFARX1 I_23033 (I394374,I2859,I394142,I394462,);
not I_23034 (I394470,I394462);
not I_23035 (I394487,I258550);
not I_23036 (I394504,I258544);
nor I_23037 (I394521,I394504,I258541);
nor I_23038 (I394134,I394470,I394521);
nor I_23039 (I394552,I394504,I258553);
and I_23040 (I394569,I394552,I258556);
or I_23041 (I394586,I394569,I258535);
DFFARX1 I_23042 (I394586,I2859,I394142,I394612,);
nor I_23043 (I394122,I394612,I394168);
not I_23044 (I394634,I394612);
and I_23045 (I394651,I394634,I394168);
nor I_23046 (I394116,I394193,I394651);
nand I_23047 (I394682,I394634,I394244);
nor I_23048 (I394110,I394504,I394682);
nand I_23049 (I394113,I394634,I394422);
nand I_23050 (I394727,I394244,I258544);
nor I_23051 (I394125,I394487,I394727);
not I_23052 (I394788,I2866);
DFFARX1 I_23053 (I182718,I2859,I394788,I394814,);
DFFARX1 I_23054 (I182715,I2859,I394788,I394831,);
not I_23055 (I394839,I394831);
not I_23056 (I394856,I182730);
nor I_23057 (I394873,I394856,I182733);
not I_23058 (I394890,I182721);
nor I_23059 (I394907,I394873,I182727);
nor I_23060 (I394924,I394831,I394907);
DFFARX1 I_23061 (I394924,I2859,I394788,I394774,);
nor I_23062 (I394955,I182727,I182733);
nand I_23063 (I394972,I394955,I182730);
DFFARX1 I_23064 (I394972,I2859,I394788,I394777,);
nor I_23065 (I395003,I394890,I182727);
nand I_23066 (I395020,I395003,I182739);
nor I_23067 (I395037,I394814,I395020);
DFFARX1 I_23068 (I395037,I2859,I394788,I394753,);
not I_23069 (I395068,I395020);
nand I_23070 (I394765,I394831,I395068);
DFFARX1 I_23071 (I395020,I2859,I394788,I395108,);
not I_23072 (I395116,I395108);
not I_23073 (I395133,I182727);
not I_23074 (I395150,I182712);
nor I_23075 (I395167,I395150,I182721);
nor I_23076 (I394780,I395116,I395167);
nor I_23077 (I395198,I395150,I182724);
and I_23078 (I395215,I395198,I182712);
or I_23079 (I395232,I395215,I182736);
DFFARX1 I_23080 (I395232,I2859,I394788,I395258,);
nor I_23081 (I394768,I395258,I394814);
not I_23082 (I395280,I395258);
and I_23083 (I395297,I395280,I394814);
nor I_23084 (I394762,I394839,I395297);
nand I_23085 (I395328,I395280,I394890);
nor I_23086 (I394756,I395150,I395328);
nand I_23087 (I394759,I395280,I395068);
nand I_23088 (I395373,I394890,I182712);
nor I_23089 (I394771,I395133,I395373);
not I_23090 (I395434,I2866);
DFFARX1 I_23091 (I329139,I2859,I395434,I395460,);
DFFARX1 I_23092 (I329136,I2859,I395434,I395477,);
not I_23093 (I395485,I395477);
not I_23094 (I395502,I329136);
nor I_23095 (I395519,I395502,I329139);
not I_23096 (I395536,I329151);
nor I_23097 (I395553,I395519,I329145);
nor I_23098 (I395570,I395477,I395553);
DFFARX1 I_23099 (I395570,I2859,I395434,I395420,);
nor I_23100 (I395601,I329145,I329139);
nand I_23101 (I395618,I395601,I329136);
DFFARX1 I_23102 (I395618,I2859,I395434,I395423,);
nor I_23103 (I395649,I395536,I329145);
nand I_23104 (I395666,I395649,I329133);
nor I_23105 (I395683,I395460,I395666);
DFFARX1 I_23106 (I395683,I2859,I395434,I395399,);
not I_23107 (I395714,I395666);
nand I_23108 (I395411,I395477,I395714);
DFFARX1 I_23109 (I395666,I2859,I395434,I395754,);
not I_23110 (I395762,I395754);
not I_23111 (I395779,I329145);
not I_23112 (I395796,I329142);
nor I_23113 (I395813,I395796,I329151);
nor I_23114 (I395426,I395762,I395813);
nor I_23115 (I395844,I395796,I329148);
and I_23116 (I395861,I395844,I329154);
or I_23117 (I395878,I395861,I329133);
DFFARX1 I_23118 (I395878,I2859,I395434,I395904,);
nor I_23119 (I395414,I395904,I395460);
not I_23120 (I395926,I395904);
and I_23121 (I395943,I395926,I395460);
nor I_23122 (I395408,I395485,I395943);
nand I_23123 (I395974,I395926,I395536);
nor I_23124 (I395402,I395796,I395974);
nand I_23125 (I395405,I395926,I395714);
nand I_23126 (I396019,I395536,I329142);
nor I_23127 (I395417,I395779,I396019);
not I_23128 (I396080,I2866);
DFFARX1 I_23129 (I2268,I2859,I396080,I396106,);
DFFARX1 I_23130 (I1468,I2859,I396080,I396123,);
not I_23131 (I396131,I396123);
not I_23132 (I396148,I1788);
nor I_23133 (I396165,I396148,I1700);
not I_23134 (I396182,I1756);
nor I_23135 (I396199,I396165,I1708);
nor I_23136 (I396216,I396123,I396199);
DFFARX1 I_23137 (I396216,I2859,I396080,I396066,);
nor I_23138 (I396247,I1708,I1700);
nand I_23139 (I396264,I396247,I1788);
DFFARX1 I_23140 (I396264,I2859,I396080,I396069,);
nor I_23141 (I396295,I396182,I1708);
nand I_23142 (I396312,I396295,I2364);
nor I_23143 (I396329,I396106,I396312);
DFFARX1 I_23144 (I396329,I2859,I396080,I396045,);
not I_23145 (I396360,I396312);
nand I_23146 (I396057,I396123,I396360);
DFFARX1 I_23147 (I396312,I2859,I396080,I396400,);
not I_23148 (I396408,I396400);
not I_23149 (I396425,I1708);
not I_23150 (I396442,I1484);
nor I_23151 (I396459,I396442,I1756);
nor I_23152 (I396072,I396408,I396459);
nor I_23153 (I396490,I396442,I2716);
and I_23154 (I396507,I396490,I2292);
or I_23155 (I396524,I396507,I2604);
DFFARX1 I_23156 (I396524,I2859,I396080,I396550,);
nor I_23157 (I396060,I396550,I396106);
not I_23158 (I396572,I396550);
and I_23159 (I396589,I396572,I396106);
nor I_23160 (I396054,I396131,I396589);
nand I_23161 (I396620,I396572,I396182);
nor I_23162 (I396048,I396442,I396620);
nand I_23163 (I396051,I396572,I396360);
nand I_23164 (I396665,I396182,I1484);
nor I_23165 (I396063,I396425,I396665);
not I_23166 (I396726,I2866);
DFFARX1 I_23167 (I183262,I2859,I396726,I396752,);
DFFARX1 I_23168 (I183259,I2859,I396726,I396769,);
not I_23169 (I396777,I396769);
not I_23170 (I396794,I183274);
nor I_23171 (I396811,I396794,I183277);
not I_23172 (I396828,I183265);
nor I_23173 (I396845,I396811,I183271);
nor I_23174 (I396862,I396769,I396845);
DFFARX1 I_23175 (I396862,I2859,I396726,I396712,);
nor I_23176 (I396893,I183271,I183277);
nand I_23177 (I396910,I396893,I183274);
DFFARX1 I_23178 (I396910,I2859,I396726,I396715,);
nor I_23179 (I396941,I396828,I183271);
nand I_23180 (I396958,I396941,I183283);
nor I_23181 (I396975,I396752,I396958);
DFFARX1 I_23182 (I396975,I2859,I396726,I396691,);
not I_23183 (I397006,I396958);
nand I_23184 (I396703,I396769,I397006);
DFFARX1 I_23185 (I396958,I2859,I396726,I397046,);
not I_23186 (I397054,I397046);
not I_23187 (I397071,I183271);
not I_23188 (I397088,I183256);
nor I_23189 (I397105,I397088,I183265);
nor I_23190 (I396718,I397054,I397105);
nor I_23191 (I397136,I397088,I183268);
and I_23192 (I397153,I397136,I183256);
or I_23193 (I397170,I397153,I183280);
DFFARX1 I_23194 (I397170,I2859,I396726,I397196,);
nor I_23195 (I396706,I397196,I396752);
not I_23196 (I397218,I397196);
and I_23197 (I397235,I397218,I396752);
nor I_23198 (I396700,I396777,I397235);
nand I_23199 (I397266,I397218,I396828);
nor I_23200 (I396694,I397088,I397266);
nand I_23201 (I396697,I397218,I397006);
nand I_23202 (I397311,I396828,I183256);
nor I_23203 (I396709,I397071,I397311);
not I_23204 (I397372,I2866);
DFFARX1 I_23205 (I246975,I2859,I397372,I397398,);
DFFARX1 I_23206 (I246987,I2859,I397372,I397415,);
not I_23207 (I397423,I397415);
not I_23208 (I397440,I246996);
nor I_23209 (I397457,I397440,I246972);
not I_23210 (I397474,I246990);
nor I_23211 (I397491,I397457,I246984);
nor I_23212 (I397508,I397415,I397491);
DFFARX1 I_23213 (I397508,I2859,I397372,I397358,);
nor I_23214 (I397539,I246984,I246972);
nand I_23215 (I397556,I397539,I246996);
DFFARX1 I_23216 (I397556,I2859,I397372,I397361,);
nor I_23217 (I397587,I397474,I246984);
nand I_23218 (I397604,I397587,I246978);
nor I_23219 (I397621,I397398,I397604);
DFFARX1 I_23220 (I397621,I2859,I397372,I397337,);
not I_23221 (I397652,I397604);
nand I_23222 (I397349,I397415,I397652);
DFFARX1 I_23223 (I397604,I2859,I397372,I397692,);
not I_23224 (I397700,I397692);
not I_23225 (I397717,I246984);
not I_23226 (I397734,I246993);
nor I_23227 (I397751,I397734,I246990);
nor I_23228 (I397364,I397700,I397751);
nor I_23229 (I397782,I397734,I246975);
and I_23230 (I397799,I397782,I246972);
or I_23231 (I397816,I397799,I246981);
DFFARX1 I_23232 (I397816,I2859,I397372,I397842,);
nor I_23233 (I397352,I397842,I397398);
not I_23234 (I397864,I397842);
and I_23235 (I397881,I397864,I397398);
nor I_23236 (I397346,I397423,I397881);
nand I_23237 (I397912,I397864,I397474);
nor I_23238 (I397340,I397734,I397912);
nand I_23239 (I397343,I397864,I397652);
nand I_23240 (I397957,I397474,I246993);
nor I_23241 (I397355,I397717,I397957);
not I_23242 (I398018,I2866);
DFFARX1 I_23243 (I23235,I2859,I398018,I398044,);
DFFARX1 I_23244 (I23241,I2859,I398018,I398061,);
not I_23245 (I398069,I398061);
not I_23246 (I398086,I23259);
nor I_23247 (I398103,I398086,I23238);
not I_23248 (I398120,I23244);
nor I_23249 (I398137,I398103,I23250);
nor I_23250 (I398154,I398061,I398137);
DFFARX1 I_23251 (I398154,I2859,I398018,I398004,);
nor I_23252 (I398185,I23250,I23238);
nand I_23253 (I398202,I398185,I23259);
DFFARX1 I_23254 (I398202,I2859,I398018,I398007,);
nor I_23255 (I398233,I398120,I23250);
nand I_23256 (I398250,I398233,I23256);
nor I_23257 (I398267,I398044,I398250);
DFFARX1 I_23258 (I398267,I2859,I398018,I397983,);
not I_23259 (I398298,I398250);
nand I_23260 (I397995,I398061,I398298);
DFFARX1 I_23261 (I398250,I2859,I398018,I398338,);
not I_23262 (I398346,I398338);
not I_23263 (I398363,I23250);
not I_23264 (I398380,I23238);
nor I_23265 (I398397,I398380,I23244);
nor I_23266 (I398010,I398346,I398397);
nor I_23267 (I398428,I398380,I23247);
and I_23268 (I398445,I398428,I23235);
or I_23269 (I398462,I398445,I23253);
DFFARX1 I_23270 (I398462,I2859,I398018,I398488,);
nor I_23271 (I397998,I398488,I398044);
not I_23272 (I398510,I398488);
and I_23273 (I398527,I398510,I398044);
nor I_23274 (I397992,I398069,I398527);
nand I_23275 (I398558,I398510,I398120);
nor I_23276 (I397986,I398380,I398558);
nand I_23277 (I397989,I398510,I398298);
nand I_23278 (I398603,I398120,I23238);
nor I_23279 (I398001,I398363,I398603);
not I_23280 (I398664,I2866);
DFFARX1 I_23281 (I278768,I2859,I398664,I398690,);
DFFARX1 I_23282 (I278762,I2859,I398664,I398707,);
not I_23283 (I398715,I398707);
not I_23284 (I398732,I278777);
nor I_23285 (I398749,I398732,I278762);
not I_23286 (I398766,I278771);
nor I_23287 (I398783,I398749,I278780);
nor I_23288 (I398800,I398707,I398783);
DFFARX1 I_23289 (I398800,I2859,I398664,I398650,);
nor I_23290 (I398831,I278780,I278762);
nand I_23291 (I398848,I398831,I278777);
DFFARX1 I_23292 (I398848,I2859,I398664,I398653,);
nor I_23293 (I398879,I398766,I278780);
nand I_23294 (I398896,I398879,I278765);
nor I_23295 (I398913,I398690,I398896);
DFFARX1 I_23296 (I398913,I2859,I398664,I398629,);
not I_23297 (I398944,I398896);
nand I_23298 (I398641,I398707,I398944);
DFFARX1 I_23299 (I398896,I2859,I398664,I398984,);
not I_23300 (I398992,I398984);
not I_23301 (I399009,I278780);
not I_23302 (I399026,I278774);
nor I_23303 (I399043,I399026,I278771);
nor I_23304 (I398656,I398992,I399043);
nor I_23305 (I399074,I399026,I278783);
and I_23306 (I399091,I399074,I278786);
or I_23307 (I399108,I399091,I278765);
DFFARX1 I_23308 (I399108,I2859,I398664,I399134,);
nor I_23309 (I398644,I399134,I398690);
not I_23310 (I399156,I399134);
and I_23311 (I399173,I399156,I398690);
nor I_23312 (I398638,I398715,I399173);
nand I_23313 (I399204,I399156,I398766);
nor I_23314 (I398632,I399026,I399204);
nand I_23315 (I398635,I399156,I398944);
nand I_23316 (I399249,I398766,I278774);
nor I_23317 (I398647,I399009,I399249);
not I_23318 (I399310,I2866);
DFFARX1 I_23319 (I213808,I2859,I399310,I399336,);
DFFARX1 I_23320 (I213820,I2859,I399310,I399353,);
not I_23321 (I399361,I399353);
not I_23322 (I399378,I213805);
nor I_23323 (I399395,I399378,I213823);
not I_23324 (I399412,I213829);
nor I_23325 (I399429,I399395,I213811);
nor I_23326 (I399446,I399353,I399429);
DFFARX1 I_23327 (I399446,I2859,I399310,I399296,);
nor I_23328 (I399477,I213811,I213823);
nand I_23329 (I399494,I399477,I213805);
DFFARX1 I_23330 (I399494,I2859,I399310,I399299,);
nor I_23331 (I399525,I399412,I213811);
nand I_23332 (I399542,I399525,I213814);
nor I_23333 (I399559,I399336,I399542);
DFFARX1 I_23334 (I399559,I2859,I399310,I399275,);
not I_23335 (I399590,I399542);
nand I_23336 (I399287,I399353,I399590);
DFFARX1 I_23337 (I399542,I2859,I399310,I399630,);
not I_23338 (I399638,I399630);
not I_23339 (I399655,I213811);
not I_23340 (I399672,I213817);
nor I_23341 (I399689,I399672,I213829);
nor I_23342 (I399302,I399638,I399689);
nor I_23343 (I399720,I399672,I213826);
and I_23344 (I399737,I399720,I213805);
or I_23345 (I399754,I399737,I213808);
DFFARX1 I_23346 (I399754,I2859,I399310,I399780,);
nor I_23347 (I399290,I399780,I399336);
not I_23348 (I399802,I399780);
and I_23349 (I399819,I399802,I399336);
nor I_23350 (I399284,I399361,I399819);
nand I_23351 (I399850,I399802,I399412);
nor I_23352 (I399278,I399672,I399850);
nand I_23353 (I399281,I399802,I399590);
nand I_23354 (I399895,I399412,I213817);
nor I_23355 (I399293,I399655,I399895);
not I_23356 (I399956,I2866);
DFFARX1 I_23357 (I349165,I2859,I399956,I399982,);
DFFARX1 I_23358 (I349162,I2859,I399956,I399999,);
not I_23359 (I400007,I399999);
not I_23360 (I400024,I349162);
nor I_23361 (I400041,I400024,I349165);
not I_23362 (I400058,I349177);
nor I_23363 (I400075,I400041,I349171);
nor I_23364 (I400092,I399999,I400075);
DFFARX1 I_23365 (I400092,I2859,I399956,I399942,);
nor I_23366 (I400123,I349171,I349165);
nand I_23367 (I400140,I400123,I349162);
DFFARX1 I_23368 (I400140,I2859,I399956,I399945,);
nor I_23369 (I400171,I400058,I349171);
nand I_23370 (I400188,I400171,I349159);
nor I_23371 (I400205,I399982,I400188);
DFFARX1 I_23372 (I400205,I2859,I399956,I399921,);
not I_23373 (I400236,I400188);
nand I_23374 (I399933,I399999,I400236);
DFFARX1 I_23375 (I400188,I2859,I399956,I400276,);
not I_23376 (I400284,I400276);
not I_23377 (I400301,I349171);
not I_23378 (I400318,I349168);
nor I_23379 (I400335,I400318,I349177);
nor I_23380 (I399948,I400284,I400335);
nor I_23381 (I400366,I400318,I349174);
and I_23382 (I400383,I400366,I349180);
or I_23383 (I400400,I400383,I349159);
DFFARX1 I_23384 (I400400,I2859,I399956,I400426,);
nor I_23385 (I399936,I400426,I399982);
not I_23386 (I400448,I400426);
and I_23387 (I400465,I400448,I399982);
nor I_23388 (I399930,I400007,I400465);
nand I_23389 (I400496,I400448,I400058);
nor I_23390 (I399924,I400318,I400496);
nand I_23391 (I399927,I400448,I400236);
nand I_23392 (I400541,I400058,I349168);
nor I_23393 (I399939,I400301,I400541);
not I_23394 (I400602,I2866);
DFFARX1 I_23395 (I97123,I2859,I400602,I400628,);
DFFARX1 I_23396 (I97135,I2859,I400602,I400645,);
not I_23397 (I400653,I400645);
not I_23398 (I400670,I97141);
nor I_23399 (I400687,I400670,I97126);
not I_23400 (I400704,I97117);
nor I_23401 (I400721,I400687,I97138);
nor I_23402 (I400738,I400645,I400721);
DFFARX1 I_23403 (I400738,I2859,I400602,I400588,);
nor I_23404 (I400769,I97138,I97126);
nand I_23405 (I400786,I400769,I97141);
DFFARX1 I_23406 (I400786,I2859,I400602,I400591,);
nor I_23407 (I400817,I400704,I97138);
nand I_23408 (I400834,I400817,I97120);
nor I_23409 (I400851,I400628,I400834);
DFFARX1 I_23410 (I400851,I2859,I400602,I400567,);
not I_23411 (I400882,I400834);
nand I_23412 (I400579,I400645,I400882);
DFFARX1 I_23413 (I400834,I2859,I400602,I400922,);
not I_23414 (I400930,I400922);
not I_23415 (I400947,I97138);
not I_23416 (I400964,I97129);
nor I_23417 (I400981,I400964,I97117);
nor I_23418 (I400594,I400930,I400981);
nor I_23419 (I401012,I400964,I97132);
and I_23420 (I401029,I401012,I97120);
or I_23421 (I401046,I401029,I97117);
DFFARX1 I_23422 (I401046,I2859,I400602,I401072,);
nor I_23423 (I400582,I401072,I400628);
not I_23424 (I401094,I401072);
and I_23425 (I401111,I401094,I400628);
nor I_23426 (I400576,I400653,I401111);
nand I_23427 (I401142,I401094,I400704);
nor I_23428 (I400570,I400964,I401142);
nand I_23429 (I400573,I401094,I400882);
nand I_23430 (I401187,I400704,I97129);
nor I_23431 (I400585,I400947,I401187);
not I_23432 (I401248,I2866);
DFFARX1 I_23433 (I138801,I2859,I401248,I401274,);
DFFARX1 I_23434 (I138807,I2859,I401248,I401291,);
not I_23435 (I401299,I401291);
not I_23436 (I401316,I138828);
nor I_23437 (I401333,I401316,I138816);
not I_23438 (I401350,I138825);
nor I_23439 (I401367,I401333,I138810);
nor I_23440 (I401384,I401291,I401367);
DFFARX1 I_23441 (I401384,I2859,I401248,I401234,);
nor I_23442 (I401415,I138810,I138816);
nand I_23443 (I401432,I401415,I138828);
DFFARX1 I_23444 (I401432,I2859,I401248,I401237,);
nor I_23445 (I401463,I401350,I138810);
nand I_23446 (I401480,I401463,I138801);
nor I_23447 (I401497,I401274,I401480);
DFFARX1 I_23448 (I401497,I2859,I401248,I401213,);
not I_23449 (I401528,I401480);
nand I_23450 (I401225,I401291,I401528);
DFFARX1 I_23451 (I401480,I2859,I401248,I401568,);
not I_23452 (I401576,I401568);
not I_23453 (I401593,I138810);
not I_23454 (I401610,I138813);
nor I_23455 (I401627,I401610,I138825);
nor I_23456 (I401240,I401576,I401627);
nor I_23457 (I401658,I401610,I138822);
and I_23458 (I401675,I401658,I138804);
or I_23459 (I401692,I401675,I138819);
DFFARX1 I_23460 (I401692,I2859,I401248,I401718,);
nor I_23461 (I401228,I401718,I401274);
not I_23462 (I401740,I401718);
and I_23463 (I401757,I401740,I401274);
nor I_23464 (I401222,I401299,I401757);
nand I_23465 (I401788,I401740,I401350);
nor I_23466 (I401216,I401610,I401788);
nand I_23467 (I401219,I401740,I401528);
nand I_23468 (I401833,I401350,I138813);
nor I_23469 (I401231,I401593,I401833);
not I_23470 (I401894,I2866);
DFFARX1 I_23471 (I455682,I2859,I401894,I401920,);
DFFARX1 I_23472 (I455664,I2859,I401894,I401937,);
not I_23473 (I401945,I401937);
not I_23474 (I401962,I455673);
nor I_23475 (I401979,I401962,I455685);
not I_23476 (I401996,I455667);
nor I_23477 (I402013,I401979,I455676);
nor I_23478 (I402030,I401937,I402013);
DFFARX1 I_23479 (I402030,I2859,I401894,I401880,);
nor I_23480 (I402061,I455676,I455685);
nand I_23481 (I402078,I402061,I455673);
DFFARX1 I_23482 (I402078,I2859,I401894,I401883,);
nor I_23483 (I402109,I401996,I455676);
nand I_23484 (I402126,I402109,I455688);
nor I_23485 (I402143,I401920,I402126);
DFFARX1 I_23486 (I402143,I2859,I401894,I401859,);
not I_23487 (I402174,I402126);
nand I_23488 (I401871,I401937,I402174);
DFFARX1 I_23489 (I402126,I2859,I401894,I402214,);
not I_23490 (I402222,I402214);
not I_23491 (I402239,I455676);
not I_23492 (I402256,I455664);
nor I_23493 (I402273,I402256,I455667);
nor I_23494 (I401886,I402222,I402273);
nor I_23495 (I402304,I402256,I455670);
and I_23496 (I402321,I402304,I455679);
or I_23497 (I402338,I402321,I455667);
DFFARX1 I_23498 (I402338,I2859,I401894,I402364,);
nor I_23499 (I401874,I402364,I401920);
not I_23500 (I402386,I402364);
and I_23501 (I402403,I402386,I401920);
nor I_23502 (I401868,I401945,I402403);
nand I_23503 (I402434,I402386,I401996);
nor I_23504 (I401862,I402256,I402434);
nand I_23505 (I401865,I402386,I402174);
nand I_23506 (I402479,I401996,I455664);
nor I_23507 (I401877,I402239,I402479);
not I_23508 (I402540,I2866);
DFFARX1 I_23509 (I242929,I2859,I402540,I402566,);
DFFARX1 I_23510 (I242941,I2859,I402540,I402583,);
not I_23511 (I402591,I402583);
not I_23512 (I402608,I242950);
nor I_23513 (I402625,I402608,I242926);
not I_23514 (I402642,I242944);
nor I_23515 (I402659,I402625,I242938);
nor I_23516 (I402676,I402583,I402659);
DFFARX1 I_23517 (I402676,I2859,I402540,I402526,);
nor I_23518 (I402707,I242938,I242926);
nand I_23519 (I402724,I402707,I242950);
DFFARX1 I_23520 (I402724,I2859,I402540,I402529,);
nor I_23521 (I402755,I402642,I242938);
nand I_23522 (I402772,I402755,I242932);
nor I_23523 (I402789,I402566,I402772);
DFFARX1 I_23524 (I402789,I2859,I402540,I402505,);
not I_23525 (I402820,I402772);
nand I_23526 (I402517,I402583,I402820);
DFFARX1 I_23527 (I402772,I2859,I402540,I402860,);
not I_23528 (I402868,I402860);
not I_23529 (I402885,I242938);
not I_23530 (I402902,I242947);
nor I_23531 (I402919,I402902,I242944);
nor I_23532 (I402532,I402868,I402919);
nor I_23533 (I402950,I402902,I242929);
and I_23534 (I402967,I402950,I242926);
or I_23535 (I402984,I402967,I242935);
DFFARX1 I_23536 (I402984,I2859,I402540,I403010,);
nor I_23537 (I402520,I403010,I402566);
not I_23538 (I403032,I403010);
and I_23539 (I403049,I403032,I402566);
nor I_23540 (I402514,I402591,I403049);
nand I_23541 (I403080,I403032,I402642);
nor I_23542 (I402508,I402902,I403080);
nand I_23543 (I402511,I403032,I402820);
nand I_23544 (I403125,I402642,I242947);
nor I_23545 (I402523,I402885,I403125);
not I_23546 (I403186,I2866);
DFFARX1 I_23547 (I70943,I2859,I403186,I403212,);
DFFARX1 I_23548 (I70955,I2859,I403186,I403229,);
not I_23549 (I403237,I403229);
not I_23550 (I403254,I70961);
nor I_23551 (I403271,I403254,I70946);
not I_23552 (I403288,I70937);
nor I_23553 (I403305,I403271,I70958);
nor I_23554 (I403322,I403229,I403305);
DFFARX1 I_23555 (I403322,I2859,I403186,I403172,);
nor I_23556 (I403353,I70958,I70946);
nand I_23557 (I403370,I403353,I70961);
DFFARX1 I_23558 (I403370,I2859,I403186,I403175,);
nor I_23559 (I403401,I403288,I70958);
nand I_23560 (I403418,I403401,I70940);
nor I_23561 (I403435,I403212,I403418);
DFFARX1 I_23562 (I403435,I2859,I403186,I403151,);
not I_23563 (I403466,I403418);
nand I_23564 (I403163,I403229,I403466);
DFFARX1 I_23565 (I403418,I2859,I403186,I403506,);
not I_23566 (I403514,I403506);
not I_23567 (I403531,I70958);
not I_23568 (I403548,I70949);
nor I_23569 (I403565,I403548,I70937);
nor I_23570 (I403178,I403514,I403565);
nor I_23571 (I403596,I403548,I70952);
and I_23572 (I403613,I403596,I70940);
or I_23573 (I403630,I403613,I70937);
DFFARX1 I_23574 (I403630,I2859,I403186,I403656,);
nor I_23575 (I403166,I403656,I403212);
not I_23576 (I403678,I403656);
and I_23577 (I403695,I403678,I403212);
nor I_23578 (I403160,I403237,I403695);
nand I_23579 (I403726,I403678,I403288);
nor I_23580 (I403154,I403548,I403726);
nand I_23581 (I403157,I403678,I403466);
nand I_23582 (I403771,I403288,I70949);
nor I_23583 (I403169,I403531,I403771);
not I_23584 (I403832,I2866);
DFFARX1 I_23585 (I285704,I2859,I403832,I403858,);
DFFARX1 I_23586 (I285698,I2859,I403832,I403875,);
not I_23587 (I403883,I403875);
not I_23588 (I403900,I285713);
nor I_23589 (I403917,I403900,I285698);
not I_23590 (I403934,I285707);
nor I_23591 (I403951,I403917,I285716);
nor I_23592 (I403968,I403875,I403951);
DFFARX1 I_23593 (I403968,I2859,I403832,I403818,);
nor I_23594 (I403999,I285716,I285698);
nand I_23595 (I404016,I403999,I285713);
DFFARX1 I_23596 (I404016,I2859,I403832,I403821,);
nor I_23597 (I404047,I403934,I285716);
nand I_23598 (I404064,I404047,I285701);
nor I_23599 (I404081,I403858,I404064);
DFFARX1 I_23600 (I404081,I2859,I403832,I403797,);
not I_23601 (I404112,I404064);
nand I_23602 (I403809,I403875,I404112);
DFFARX1 I_23603 (I404064,I2859,I403832,I404152,);
not I_23604 (I404160,I404152);
not I_23605 (I404177,I285716);
not I_23606 (I404194,I285710);
nor I_23607 (I404211,I404194,I285707);
nor I_23608 (I403824,I404160,I404211);
nor I_23609 (I404242,I404194,I285719);
and I_23610 (I404259,I404242,I285722);
or I_23611 (I404276,I404259,I285701);
DFFARX1 I_23612 (I404276,I2859,I403832,I404302,);
nor I_23613 (I403812,I404302,I403858);
not I_23614 (I404324,I404302);
and I_23615 (I404341,I404324,I403858);
nor I_23616 (I403806,I403883,I404341);
nand I_23617 (I404372,I404324,I403934);
nor I_23618 (I403800,I404194,I404372);
nand I_23619 (I403803,I404324,I404112);
nand I_23620 (I404417,I403934,I285710);
nor I_23621 (I403815,I404177,I404417);
not I_23622 (I404478,I2866);
DFFARX1 I_23623 (I488628,I2859,I404478,I404504,);
DFFARX1 I_23624 (I488610,I2859,I404478,I404521,);
not I_23625 (I404529,I404521);
not I_23626 (I404546,I488619);
nor I_23627 (I404563,I404546,I488631);
not I_23628 (I404580,I488613);
nor I_23629 (I404597,I404563,I488622);
nor I_23630 (I404614,I404521,I404597);
DFFARX1 I_23631 (I404614,I2859,I404478,I404464,);
nor I_23632 (I404645,I488622,I488631);
nand I_23633 (I404662,I404645,I488619);
DFFARX1 I_23634 (I404662,I2859,I404478,I404467,);
nor I_23635 (I404693,I404580,I488622);
nand I_23636 (I404710,I404693,I488634);
nor I_23637 (I404727,I404504,I404710);
DFFARX1 I_23638 (I404727,I2859,I404478,I404443,);
not I_23639 (I404758,I404710);
nand I_23640 (I404455,I404521,I404758);
DFFARX1 I_23641 (I404710,I2859,I404478,I404798,);
not I_23642 (I404806,I404798);
not I_23643 (I404823,I488622);
not I_23644 (I404840,I488610);
nor I_23645 (I404857,I404840,I488613);
nor I_23646 (I404470,I404806,I404857);
nor I_23647 (I404888,I404840,I488616);
and I_23648 (I404905,I404888,I488625);
or I_23649 (I404922,I404905,I488613);
DFFARX1 I_23650 (I404922,I2859,I404478,I404948,);
nor I_23651 (I404458,I404948,I404504);
not I_23652 (I404970,I404948);
and I_23653 (I404987,I404970,I404504);
nor I_23654 (I404452,I404529,I404987);
nand I_23655 (I405018,I404970,I404580);
nor I_23656 (I404446,I404840,I405018);
nand I_23657 (I404449,I404970,I404758);
nand I_23658 (I405063,I404580,I488610);
nor I_23659 (I404461,I404823,I405063);
not I_23660 (I405124,I2866);
DFFARX1 I_23661 (I356543,I2859,I405124,I405150,);
DFFARX1 I_23662 (I356540,I2859,I405124,I405167,);
not I_23663 (I405175,I405167);
not I_23664 (I405192,I356540);
nor I_23665 (I405209,I405192,I356543);
not I_23666 (I405226,I356555);
nor I_23667 (I405243,I405209,I356549);
nor I_23668 (I405260,I405167,I405243);
DFFARX1 I_23669 (I405260,I2859,I405124,I405110,);
nor I_23670 (I405291,I356549,I356543);
nand I_23671 (I405308,I405291,I356540);
DFFARX1 I_23672 (I405308,I2859,I405124,I405113,);
nor I_23673 (I405339,I405226,I356549);
nand I_23674 (I405356,I405339,I356537);
nor I_23675 (I405373,I405150,I405356);
DFFARX1 I_23676 (I405373,I2859,I405124,I405089,);
not I_23677 (I405404,I405356);
nand I_23678 (I405101,I405167,I405404);
DFFARX1 I_23679 (I405356,I2859,I405124,I405444,);
not I_23680 (I405452,I405444);
not I_23681 (I405469,I356549);
not I_23682 (I405486,I356546);
nor I_23683 (I405503,I405486,I356555);
nor I_23684 (I405116,I405452,I405503);
nor I_23685 (I405534,I405486,I356552);
and I_23686 (I405551,I405534,I356558);
or I_23687 (I405568,I405551,I356537);
DFFARX1 I_23688 (I405568,I2859,I405124,I405594,);
nor I_23689 (I405104,I405594,I405150);
not I_23690 (I405616,I405594);
and I_23691 (I405633,I405616,I405150);
nor I_23692 (I405098,I405175,I405633);
nand I_23693 (I405664,I405616,I405226);
nor I_23694 (I405092,I405486,I405664);
nand I_23695 (I405095,I405616,I405404);
nand I_23696 (I405709,I405226,I356546);
nor I_23697 (I405107,I405469,I405709);
not I_23698 (I405770,I2866);
DFFARX1 I_23699 (I136166,I2859,I405770,I405796,);
DFFARX1 I_23700 (I136172,I2859,I405770,I405813,);
not I_23701 (I405821,I405813);
not I_23702 (I405838,I136193);
nor I_23703 (I405855,I405838,I136181);
not I_23704 (I405872,I136190);
nor I_23705 (I405889,I405855,I136175);
nor I_23706 (I405906,I405813,I405889);
DFFARX1 I_23707 (I405906,I2859,I405770,I405756,);
nor I_23708 (I405937,I136175,I136181);
nand I_23709 (I405954,I405937,I136193);
DFFARX1 I_23710 (I405954,I2859,I405770,I405759,);
nor I_23711 (I405985,I405872,I136175);
nand I_23712 (I406002,I405985,I136166);
nor I_23713 (I406019,I405796,I406002);
DFFARX1 I_23714 (I406019,I2859,I405770,I405735,);
not I_23715 (I406050,I406002);
nand I_23716 (I405747,I405813,I406050);
DFFARX1 I_23717 (I406002,I2859,I405770,I406090,);
not I_23718 (I406098,I406090);
not I_23719 (I406115,I136175);
not I_23720 (I406132,I136178);
nor I_23721 (I406149,I406132,I136190);
nor I_23722 (I405762,I406098,I406149);
nor I_23723 (I406180,I406132,I136187);
and I_23724 (I406197,I406180,I136169);
or I_23725 (I406214,I406197,I136184);
DFFARX1 I_23726 (I406214,I2859,I405770,I406240,);
nor I_23727 (I405750,I406240,I405796);
not I_23728 (I406262,I406240);
and I_23729 (I406279,I406262,I405796);
nor I_23730 (I405744,I405821,I406279);
nand I_23731 (I406310,I406262,I405872);
nor I_23732 (I405738,I406132,I406310);
nand I_23733 (I405741,I406262,I406050);
nand I_23734 (I406355,I405872,I136178);
nor I_23735 (I405753,I406115,I406355);
not I_23736 (I406416,I2866);
DFFARX1 I_23737 (I88198,I2859,I406416,I406442,);
DFFARX1 I_23738 (I88210,I2859,I406416,I406459,);
not I_23739 (I406467,I406459);
not I_23740 (I406484,I88216);
nor I_23741 (I406501,I406484,I88201);
not I_23742 (I406518,I88192);
nor I_23743 (I406535,I406501,I88213);
nor I_23744 (I406552,I406459,I406535);
DFFARX1 I_23745 (I406552,I2859,I406416,I406402,);
nor I_23746 (I406583,I88213,I88201);
nand I_23747 (I406600,I406583,I88216);
DFFARX1 I_23748 (I406600,I2859,I406416,I406405,);
nor I_23749 (I406631,I406518,I88213);
nand I_23750 (I406648,I406631,I88195);
nor I_23751 (I406665,I406442,I406648);
DFFARX1 I_23752 (I406665,I2859,I406416,I406381,);
not I_23753 (I406696,I406648);
nand I_23754 (I406393,I406459,I406696);
DFFARX1 I_23755 (I406648,I2859,I406416,I406736,);
not I_23756 (I406744,I406736);
not I_23757 (I406761,I88213);
not I_23758 (I406778,I88204);
nor I_23759 (I406795,I406778,I88192);
nor I_23760 (I406408,I406744,I406795);
nor I_23761 (I406826,I406778,I88207);
and I_23762 (I406843,I406826,I88195);
or I_23763 (I406860,I406843,I88192);
DFFARX1 I_23764 (I406860,I2859,I406416,I406886,);
nor I_23765 (I406396,I406886,I406442);
not I_23766 (I406908,I406886);
and I_23767 (I406925,I406908,I406442);
nor I_23768 (I406390,I406467,I406925);
nand I_23769 (I406956,I406908,I406518);
nor I_23770 (I406384,I406778,I406956);
nand I_23771 (I406387,I406908,I406696);
nand I_23772 (I407001,I406518,I88204);
nor I_23773 (I406399,I406761,I407001);
not I_23774 (I407062,I2866);
DFFARX1 I_23775 (I347584,I2859,I407062,I407088,);
DFFARX1 I_23776 (I347581,I2859,I407062,I407105,);
not I_23777 (I407113,I407105);
not I_23778 (I407130,I347581);
nor I_23779 (I407147,I407130,I347584);
not I_23780 (I407164,I347596);
nor I_23781 (I407181,I407147,I347590);
nor I_23782 (I407198,I407105,I407181);
DFFARX1 I_23783 (I407198,I2859,I407062,I407048,);
nor I_23784 (I407229,I347590,I347584);
nand I_23785 (I407246,I407229,I347581);
DFFARX1 I_23786 (I407246,I2859,I407062,I407051,);
nor I_23787 (I407277,I407164,I347590);
nand I_23788 (I407294,I407277,I347578);
nor I_23789 (I407311,I407088,I407294);
DFFARX1 I_23790 (I407311,I2859,I407062,I407027,);
not I_23791 (I407342,I407294);
nand I_23792 (I407039,I407105,I407342);
DFFARX1 I_23793 (I407294,I2859,I407062,I407382,);
not I_23794 (I407390,I407382);
not I_23795 (I407407,I347590);
not I_23796 (I407424,I347587);
nor I_23797 (I407441,I407424,I347596);
nor I_23798 (I407054,I407390,I407441);
nor I_23799 (I407472,I407424,I347593);
and I_23800 (I407489,I407472,I347599);
or I_23801 (I407506,I407489,I347578);
DFFARX1 I_23802 (I407506,I2859,I407062,I407532,);
nor I_23803 (I407042,I407532,I407088);
not I_23804 (I407554,I407532);
and I_23805 (I407571,I407554,I407088);
nor I_23806 (I407036,I407113,I407571);
nand I_23807 (I407602,I407554,I407164);
nor I_23808 (I407030,I407424,I407602);
nand I_23809 (I407033,I407554,I407342);
nand I_23810 (I407647,I407164,I347587);
nor I_23811 (I407045,I407407,I407647);
not I_23812 (I407708,I2866);
DFFARX1 I_23813 (I217973,I2859,I407708,I407734,);
DFFARX1 I_23814 (I217985,I2859,I407708,I407751,);
not I_23815 (I407759,I407751);
not I_23816 (I407776,I217970);
nor I_23817 (I407793,I407776,I217988);
not I_23818 (I407810,I217994);
nor I_23819 (I407827,I407793,I217976);
nor I_23820 (I407844,I407751,I407827);
DFFARX1 I_23821 (I407844,I2859,I407708,I407694,);
nor I_23822 (I407875,I217976,I217988);
nand I_23823 (I407892,I407875,I217970);
DFFARX1 I_23824 (I407892,I2859,I407708,I407697,);
nor I_23825 (I407923,I407810,I217976);
nand I_23826 (I407940,I407923,I217979);
nor I_23827 (I407957,I407734,I407940);
DFFARX1 I_23828 (I407957,I2859,I407708,I407673,);
not I_23829 (I407988,I407940);
nand I_23830 (I407685,I407751,I407988);
DFFARX1 I_23831 (I407940,I2859,I407708,I408028,);
not I_23832 (I408036,I408028);
not I_23833 (I408053,I217976);
not I_23834 (I408070,I217982);
nor I_23835 (I408087,I408070,I217994);
nor I_23836 (I407700,I408036,I408087);
nor I_23837 (I408118,I408070,I217991);
and I_23838 (I408135,I408118,I217970);
or I_23839 (I408152,I408135,I217973);
DFFARX1 I_23840 (I408152,I2859,I407708,I408178,);
nor I_23841 (I407688,I408178,I407734);
not I_23842 (I408200,I408178);
and I_23843 (I408217,I408200,I407734);
nor I_23844 (I407682,I407759,I408217);
nand I_23845 (I408248,I408200,I407810);
nor I_23846 (I407676,I408070,I408248);
nand I_23847 (I407679,I408200,I407988);
nand I_23848 (I408293,I407810,I217982);
nor I_23849 (I407691,I408053,I408293);
not I_23850 (I408354,I2866);
DFFARX1 I_23851 (I208453,I2859,I408354,I408380,);
DFFARX1 I_23852 (I208465,I2859,I408354,I408397,);
not I_23853 (I408405,I408397);
not I_23854 (I408422,I208450);
nor I_23855 (I408439,I408422,I208468);
not I_23856 (I408456,I208474);
nor I_23857 (I408473,I408439,I208456);
nor I_23858 (I408490,I408397,I408473);
DFFARX1 I_23859 (I408490,I2859,I408354,I408340,);
nor I_23860 (I408521,I208456,I208468);
nand I_23861 (I408538,I408521,I208450);
DFFARX1 I_23862 (I408538,I2859,I408354,I408343,);
nor I_23863 (I408569,I408456,I208456);
nand I_23864 (I408586,I408569,I208459);
nor I_23865 (I408603,I408380,I408586);
DFFARX1 I_23866 (I408603,I2859,I408354,I408319,);
not I_23867 (I408634,I408586);
nand I_23868 (I408331,I408397,I408634);
DFFARX1 I_23869 (I408586,I2859,I408354,I408674,);
not I_23870 (I408682,I408674);
not I_23871 (I408699,I208456);
not I_23872 (I408716,I208462);
nor I_23873 (I408733,I408716,I208474);
nor I_23874 (I408346,I408682,I408733);
nor I_23875 (I408764,I408716,I208471);
and I_23876 (I408781,I408764,I208450);
or I_23877 (I408798,I408781,I208453);
DFFARX1 I_23878 (I408798,I2859,I408354,I408824,);
nor I_23879 (I408334,I408824,I408380);
not I_23880 (I408846,I408824);
and I_23881 (I408863,I408846,I408380);
nor I_23882 (I408328,I408405,I408863);
nand I_23883 (I408894,I408846,I408456);
nor I_23884 (I408322,I408716,I408894);
nand I_23885 (I408325,I408846,I408634);
nand I_23886 (I408939,I408456,I208462);
nor I_23887 (I408337,I408699,I408939);
not I_23888 (I409000,I2866);
DFFARX1 I_23889 (I438920,I2859,I409000,I409026,);
DFFARX1 I_23890 (I438902,I2859,I409000,I409043,);
not I_23891 (I409051,I409043);
not I_23892 (I409068,I438911);
nor I_23893 (I409085,I409068,I438923);
not I_23894 (I409102,I438905);
nor I_23895 (I409119,I409085,I438914);
nor I_23896 (I409136,I409043,I409119);
DFFARX1 I_23897 (I409136,I2859,I409000,I408986,);
nor I_23898 (I409167,I438914,I438923);
nand I_23899 (I409184,I409167,I438911);
DFFARX1 I_23900 (I409184,I2859,I409000,I408989,);
nor I_23901 (I409215,I409102,I438914);
nand I_23902 (I409232,I409215,I438926);
nor I_23903 (I409249,I409026,I409232);
DFFARX1 I_23904 (I409249,I2859,I409000,I408965,);
not I_23905 (I409280,I409232);
nand I_23906 (I408977,I409043,I409280);
DFFARX1 I_23907 (I409232,I2859,I409000,I409320,);
not I_23908 (I409328,I409320);
not I_23909 (I409345,I438914);
not I_23910 (I409362,I438902);
nor I_23911 (I409379,I409362,I438905);
nor I_23912 (I408992,I409328,I409379);
nor I_23913 (I409410,I409362,I438908);
and I_23914 (I409427,I409410,I438917);
or I_23915 (I409444,I409427,I438905);
DFFARX1 I_23916 (I409444,I2859,I409000,I409470,);
nor I_23917 (I408980,I409470,I409026);
not I_23918 (I409492,I409470);
and I_23919 (I409509,I409492,I409026);
nor I_23920 (I408974,I409051,I409509);
nand I_23921 (I409540,I409492,I409102);
nor I_23922 (I408968,I409362,I409540);
nand I_23923 (I408971,I409492,I409280);
nand I_23924 (I409585,I409102,I438902);
nor I_23925 (I408983,I409345,I409585);
not I_23926 (I409646,I2866);
DFFARX1 I_23927 (I106048,I2859,I409646,I409672,);
DFFARX1 I_23928 (I106060,I2859,I409646,I409689,);
not I_23929 (I409697,I409689);
not I_23930 (I409714,I106066);
nor I_23931 (I409731,I409714,I106051);
not I_23932 (I409748,I106042);
nor I_23933 (I409765,I409731,I106063);
nor I_23934 (I409782,I409689,I409765);
DFFARX1 I_23935 (I409782,I2859,I409646,I409632,);
nor I_23936 (I409813,I106063,I106051);
nand I_23937 (I409830,I409813,I106066);
DFFARX1 I_23938 (I409830,I2859,I409646,I409635,);
nor I_23939 (I409861,I409748,I106063);
nand I_23940 (I409878,I409861,I106045);
nor I_23941 (I409895,I409672,I409878);
DFFARX1 I_23942 (I409895,I2859,I409646,I409611,);
not I_23943 (I409926,I409878);
nand I_23944 (I409623,I409689,I409926);
DFFARX1 I_23945 (I409878,I2859,I409646,I409966,);
not I_23946 (I409974,I409966);
not I_23947 (I409991,I106063);
not I_23948 (I410008,I106054);
nor I_23949 (I410025,I410008,I106042);
nor I_23950 (I409638,I409974,I410025);
nor I_23951 (I410056,I410008,I106057);
and I_23952 (I410073,I410056,I106045);
or I_23953 (I410090,I410073,I106042);
DFFARX1 I_23954 (I410090,I2859,I409646,I410116,);
nor I_23955 (I409626,I410116,I409672);
not I_23956 (I410138,I410116);
and I_23957 (I410155,I410138,I409672);
nor I_23958 (I409620,I409697,I410155);
nand I_23959 (I410186,I410138,I409748);
nor I_23960 (I409614,I410008,I410186);
nand I_23961 (I409617,I410138,I409926);
nand I_23962 (I410231,I409748,I106054);
nor I_23963 (I409629,I409991,I410231);
not I_23964 (I410292,I2866);
DFFARX1 I_23965 (I418145,I2859,I410292,I410318,);
DFFARX1 I_23966 (I418148,I2859,I410292,I410335,);
not I_23967 (I410343,I410335);
not I_23968 (I410360,I418145);
nor I_23969 (I410377,I410360,I418157);
not I_23970 (I410394,I418166);
nor I_23971 (I410411,I410377,I418154);
nor I_23972 (I410428,I410335,I410411);
DFFARX1 I_23973 (I410428,I2859,I410292,I410278,);
nor I_23974 (I410459,I418154,I418157);
nand I_23975 (I410476,I410459,I418145);
DFFARX1 I_23976 (I410476,I2859,I410292,I410281,);
nor I_23977 (I410507,I410394,I418154);
nand I_23978 (I410524,I410507,I418160);
nor I_23979 (I410541,I410318,I410524);
DFFARX1 I_23980 (I410541,I2859,I410292,I410257,);
not I_23981 (I410572,I410524);
nand I_23982 (I410269,I410335,I410572);
DFFARX1 I_23983 (I410524,I2859,I410292,I410612,);
not I_23984 (I410620,I410612);
not I_23985 (I410637,I418154);
not I_23986 (I410654,I418151);
nor I_23987 (I410671,I410654,I418166);
nor I_23988 (I410284,I410620,I410671);
nor I_23989 (I410702,I410654,I418163);
and I_23990 (I410719,I410702,I418151);
or I_23991 (I410736,I410719,I418148);
DFFARX1 I_23992 (I410736,I2859,I410292,I410762,);
nor I_23993 (I410272,I410762,I410318);
not I_23994 (I410784,I410762);
and I_23995 (I410801,I410784,I410318);
nor I_23996 (I410266,I410343,I410801);
nand I_23997 (I410832,I410784,I410394);
nor I_23998 (I410260,I410654,I410832);
nand I_23999 (I410263,I410784,I410572);
nand I_24000 (I410877,I410394,I418151);
nor I_24001 (I410275,I410637,I410877);
not I_24002 (I410938,I2866);
DFFARX1 I_24003 (I32721,I2859,I410938,I410964,);
DFFARX1 I_24004 (I32727,I2859,I410938,I410981,);
not I_24005 (I410989,I410981);
not I_24006 (I411006,I32745);
nor I_24007 (I411023,I411006,I32724);
not I_24008 (I411040,I32730);
nor I_24009 (I411057,I411023,I32736);
nor I_24010 (I411074,I410981,I411057);
DFFARX1 I_24011 (I411074,I2859,I410938,I410924,);
nor I_24012 (I411105,I32736,I32724);
nand I_24013 (I411122,I411105,I32745);
DFFARX1 I_24014 (I411122,I2859,I410938,I410927,);
nor I_24015 (I411153,I411040,I32736);
nand I_24016 (I411170,I411153,I32742);
nor I_24017 (I411187,I410964,I411170);
DFFARX1 I_24018 (I411187,I2859,I410938,I410903,);
not I_24019 (I411218,I411170);
nand I_24020 (I410915,I410981,I411218);
DFFARX1 I_24021 (I411170,I2859,I410938,I411258,);
not I_24022 (I411266,I411258);
not I_24023 (I411283,I32736);
not I_24024 (I411300,I32724);
nor I_24025 (I411317,I411300,I32730);
nor I_24026 (I410930,I411266,I411317);
nor I_24027 (I411348,I411300,I32733);
and I_24028 (I411365,I411348,I32721);
or I_24029 (I411382,I411365,I32739);
DFFARX1 I_24030 (I411382,I2859,I410938,I411408,);
nor I_24031 (I410918,I411408,I410964);
not I_24032 (I411430,I411408);
and I_24033 (I411447,I411430,I410964);
nor I_24034 (I410912,I410989,I411447);
nand I_24035 (I411478,I411430,I411040);
nor I_24036 (I410906,I411300,I411478);
nand I_24037 (I410909,I411430,I411218);
nand I_24038 (I411523,I411040,I32724);
nor I_24039 (I410921,I411283,I411523);
not I_24040 (I411584,I2866);
DFFARX1 I_24041 (I518335,I2859,I411584,I411610,);
DFFARX1 I_24042 (I518329,I2859,I411584,I411627,);
not I_24043 (I411635,I411627);
not I_24044 (I411652,I518338);
nor I_24045 (I411669,I411652,I518350);
not I_24046 (I411686,I518332);
nor I_24047 (I411703,I411669,I518329);
nor I_24048 (I411720,I411627,I411703);
DFFARX1 I_24049 (I411720,I2859,I411584,I411570,);
nor I_24050 (I411751,I518329,I518350);
nand I_24051 (I411768,I411751,I518338);
DFFARX1 I_24052 (I411768,I2859,I411584,I411573,);
nor I_24053 (I411799,I411686,I518329);
nand I_24054 (I411816,I411799,I518326);
nor I_24055 (I411833,I411610,I411816);
DFFARX1 I_24056 (I411833,I2859,I411584,I411549,);
not I_24057 (I411864,I411816);
nand I_24058 (I411561,I411627,I411864);
DFFARX1 I_24059 (I411816,I2859,I411584,I411904,);
not I_24060 (I411912,I411904);
not I_24061 (I411929,I518329);
not I_24062 (I411946,I518347);
nor I_24063 (I411963,I411946,I518332);
nor I_24064 (I411576,I411912,I411963);
nor I_24065 (I411994,I411946,I518341);
and I_24066 (I412011,I411994,I518326);
or I_24067 (I412028,I412011,I518344);
DFFARX1 I_24068 (I412028,I2859,I411584,I412054,);
nor I_24069 (I411564,I412054,I411610);
not I_24070 (I412076,I412054);
and I_24071 (I412093,I412076,I411610);
nor I_24072 (I411558,I411635,I412093);
nand I_24073 (I412124,I412076,I411686);
nor I_24074 (I411552,I411946,I412124);
nand I_24075 (I411555,I412076,I411864);
nand I_24076 (I412169,I411686,I518347);
nor I_24077 (I411567,I411929,I412169);
not I_24078 (I412230,I2866);
DFFARX1 I_24079 (I49585,I2859,I412230,I412256,);
DFFARX1 I_24080 (I49591,I2859,I412230,I412273,);
not I_24081 (I412281,I412273);
not I_24082 (I412298,I49609);
nor I_24083 (I412315,I412298,I49588);
not I_24084 (I412332,I49594);
nor I_24085 (I412349,I412315,I49600);
nor I_24086 (I412366,I412273,I412349);
DFFARX1 I_24087 (I412366,I2859,I412230,I412216,);
nor I_24088 (I412397,I49600,I49588);
nand I_24089 (I412414,I412397,I49609);
DFFARX1 I_24090 (I412414,I2859,I412230,I412219,);
nor I_24091 (I412445,I412332,I49600);
nand I_24092 (I412462,I412445,I49606);
nor I_24093 (I412479,I412256,I412462);
DFFARX1 I_24094 (I412479,I2859,I412230,I412195,);
not I_24095 (I412510,I412462);
nand I_24096 (I412207,I412273,I412510);
DFFARX1 I_24097 (I412462,I2859,I412230,I412550,);
not I_24098 (I412558,I412550);
not I_24099 (I412575,I49600);
not I_24100 (I412592,I49588);
nor I_24101 (I412609,I412592,I49594);
nor I_24102 (I412222,I412558,I412609);
nor I_24103 (I412640,I412592,I49597);
and I_24104 (I412657,I412640,I49585);
or I_24105 (I412674,I412657,I49603);
DFFARX1 I_24106 (I412674,I2859,I412230,I412700,);
nor I_24107 (I412210,I412700,I412256);
not I_24108 (I412722,I412700);
and I_24109 (I412739,I412722,I412256);
nor I_24110 (I412204,I412281,I412739);
nand I_24111 (I412770,I412722,I412332);
nor I_24112 (I412198,I412592,I412770);
nand I_24113 (I412201,I412722,I412510);
nand I_24114 (I412815,I412332,I49588);
nor I_24115 (I412213,I412575,I412815);
not I_24116 (I412876,I2866);
DFFARX1 I_24117 (I224433,I2859,I412876,I412902,);
DFFARX1 I_24118 (I224445,I2859,I412876,I412919,);
not I_24119 (I412927,I412919);
not I_24120 (I412944,I224454);
nor I_24121 (I412961,I412944,I224430);
not I_24122 (I412978,I224448);
nor I_24123 (I412995,I412961,I224442);
nor I_24124 (I413012,I412919,I412995);
DFFARX1 I_24125 (I413012,I2859,I412876,I412862,);
nor I_24126 (I413043,I224442,I224430);
nand I_24127 (I413060,I413043,I224454);
DFFARX1 I_24128 (I413060,I2859,I412876,I412865,);
nor I_24129 (I413091,I412978,I224442);
nand I_24130 (I413108,I413091,I224436);
nor I_24131 (I413125,I412902,I413108);
DFFARX1 I_24132 (I413125,I2859,I412876,I412841,);
not I_24133 (I413156,I413108);
nand I_24134 (I412853,I412919,I413156);
DFFARX1 I_24135 (I413108,I2859,I412876,I413196,);
not I_24136 (I413204,I413196);
not I_24137 (I413221,I224442);
not I_24138 (I413238,I224451);
nor I_24139 (I413255,I413238,I224448);
nor I_24140 (I412868,I413204,I413255);
nor I_24141 (I413286,I413238,I224433);
and I_24142 (I413303,I413286,I224430);
or I_24143 (I413320,I413303,I224439);
DFFARX1 I_24144 (I413320,I2859,I412876,I413346,);
nor I_24145 (I412856,I413346,I412902);
not I_24146 (I413368,I413346);
and I_24147 (I413385,I413368,I412902);
nor I_24148 (I412850,I412927,I413385);
nand I_24149 (I413416,I413368,I412978);
nor I_24150 (I412844,I413238,I413416);
nand I_24151 (I412847,I413368,I413156);
nand I_24152 (I413461,I412978,I224451);
nor I_24153 (I412859,I413221,I413461);
not I_24154 (I413522,I2866);
DFFARX1 I_24155 (I339152,I2859,I413522,I413548,);
DFFARX1 I_24156 (I339149,I2859,I413522,I413565,);
not I_24157 (I413573,I413565);
not I_24158 (I413590,I339149);
nor I_24159 (I413607,I413590,I339152);
not I_24160 (I413624,I339164);
nor I_24161 (I413641,I413607,I339158);
nor I_24162 (I413658,I413565,I413641);
DFFARX1 I_24163 (I413658,I2859,I413522,I413508,);
nor I_24164 (I413689,I339158,I339152);
nand I_24165 (I413706,I413689,I339149);
DFFARX1 I_24166 (I413706,I2859,I413522,I413511,);
nor I_24167 (I413737,I413624,I339158);
nand I_24168 (I413754,I413737,I339146);
nor I_24169 (I413771,I413548,I413754);
DFFARX1 I_24170 (I413771,I2859,I413522,I413487,);
not I_24171 (I413802,I413754);
nand I_24172 (I413499,I413565,I413802);
DFFARX1 I_24173 (I413754,I2859,I413522,I413842,);
not I_24174 (I413850,I413842);
not I_24175 (I413867,I339158);
not I_24176 (I413884,I339155);
nor I_24177 (I413901,I413884,I339164);
nor I_24178 (I413514,I413850,I413901);
nor I_24179 (I413932,I413884,I339161);
and I_24180 (I413949,I413932,I339167);
or I_24181 (I413966,I413949,I339146);
DFFARX1 I_24182 (I413966,I2859,I413522,I413992,);
nor I_24183 (I413502,I413992,I413548);
not I_24184 (I414014,I413992);
and I_24185 (I414031,I414014,I413548);
nor I_24186 (I413496,I413573,I414031);
nand I_24187 (I414062,I414014,I413624);
nor I_24188 (I413490,I413884,I414062);
nand I_24189 (I413493,I414014,I413802);
nand I_24190 (I414107,I413624,I339155);
nor I_24191 (I413505,I413867,I414107);
not I_24192 (I414168,I2866);
DFFARX1 I_24193 (I41153,I2859,I414168,I414194,);
DFFARX1 I_24194 (I41159,I2859,I414168,I414211,);
not I_24195 (I414219,I414211);
not I_24196 (I414236,I41177);
nor I_24197 (I414253,I414236,I41156);
not I_24198 (I414270,I41162);
nor I_24199 (I414287,I414253,I41168);
nor I_24200 (I414304,I414211,I414287);
DFFARX1 I_24201 (I414304,I2859,I414168,I414154,);
nor I_24202 (I414335,I41168,I41156);
nand I_24203 (I414352,I414335,I41177);
DFFARX1 I_24204 (I414352,I2859,I414168,I414157,);
nor I_24205 (I414383,I414270,I41168);
nand I_24206 (I414400,I414383,I41174);
nor I_24207 (I414417,I414194,I414400);
DFFARX1 I_24208 (I414417,I2859,I414168,I414133,);
not I_24209 (I414448,I414400);
nand I_24210 (I414145,I414211,I414448);
DFFARX1 I_24211 (I414400,I2859,I414168,I414488,);
not I_24212 (I414496,I414488);
not I_24213 (I414513,I41168);
not I_24214 (I414530,I41156);
nor I_24215 (I414547,I414530,I41162);
nor I_24216 (I414160,I414496,I414547);
nor I_24217 (I414578,I414530,I41165);
and I_24218 (I414595,I414578,I41153);
or I_24219 (I414612,I414595,I41171);
DFFARX1 I_24220 (I414612,I2859,I414168,I414638,);
nor I_24221 (I414148,I414638,I414194);
not I_24222 (I414660,I414638);
and I_24223 (I414677,I414660,I414194);
nor I_24224 (I414142,I414219,I414677);
nand I_24225 (I414708,I414660,I414270);
nor I_24226 (I414136,I414530,I414708);
nand I_24227 (I414139,I414660,I414448);
nand I_24228 (I414753,I414270,I41156);
nor I_24229 (I414151,I414513,I414753);
not I_24230 (I414808,I2866);
DFFARX1 I_24231 (I314023,I2859,I414808,I414834,);
DFFARX1 I_24232 (I414834,I2859,I414808,I414851,);
not I_24233 (I414800,I414851);
not I_24234 (I414873,I414834);
DFFARX1 I_24235 (I314035,I2859,I414808,I414899,);
nand I_24236 (I414907,I414899,I314044);
not I_24237 (I414924,I314044);
not I_24238 (I414941,I314026);
nand I_24239 (I414958,I314029,I314020);
and I_24240 (I414975,I314029,I314020);
not I_24241 (I414992,I314038);
nand I_24242 (I415009,I414992,I414941);
nor I_24243 (I414782,I415009,I414907);
nor I_24244 (I415040,I414924,I415009);
nand I_24245 (I414785,I414975,I415040);
not I_24246 (I415071,I314041);
nor I_24247 (I415088,I415071,I314029);
nor I_24248 (I415105,I415088,I314038);
nor I_24249 (I415122,I414873,I415105);
DFFARX1 I_24250 (I415122,I2859,I414808,I414794,);
not I_24251 (I415153,I415088);
DFFARX1 I_24252 (I415153,I2859,I414808,I414797,);
and I_24253 (I414791,I414899,I415088);
nor I_24254 (I415198,I415071,I314020);
and I_24255 (I415215,I415198,I314032);
or I_24256 (I415232,I415215,I314023);
DFFARX1 I_24257 (I415232,I2859,I414808,I415258,);
nor I_24258 (I415266,I415258,I414992);
DFFARX1 I_24259 (I415266,I2859,I414808,I414779,);
nand I_24260 (I415297,I415258,I414899);
nand I_24261 (I415314,I414992,I415297);
nor I_24262 (I414788,I415314,I414958);
not I_24263 (I415369,I2866);
DFFARX1 I_24264 (I358127,I2859,I415369,I415395,);
DFFARX1 I_24265 (I415395,I2859,I415369,I415412,);
not I_24266 (I415361,I415412);
not I_24267 (I415434,I415395);
DFFARX1 I_24268 (I358124,I2859,I415369,I415460,);
nand I_24269 (I415468,I415460,I358139);
not I_24270 (I415485,I358139);
not I_24271 (I415502,I358136);
nand I_24272 (I415519,I358133,I358121);
and I_24273 (I415536,I358133,I358121);
not I_24274 (I415553,I358118);
nand I_24275 (I415570,I415553,I415502);
nor I_24276 (I415343,I415570,I415468);
nor I_24277 (I415601,I415485,I415570);
nand I_24278 (I415346,I415536,I415601);
not I_24279 (I415632,I358124);
nor I_24280 (I415649,I415632,I358133);
nor I_24281 (I415666,I415649,I358118);
nor I_24282 (I415683,I415434,I415666);
DFFARX1 I_24283 (I415683,I2859,I415369,I415355,);
not I_24284 (I415714,I415649);
DFFARX1 I_24285 (I415714,I2859,I415369,I415358,);
and I_24286 (I415352,I415460,I415649);
nor I_24287 (I415759,I415632,I358130);
and I_24288 (I415776,I415759,I358118);
or I_24289 (I415793,I415776,I358121);
DFFARX1 I_24290 (I415793,I2859,I415369,I415819,);
nor I_24291 (I415827,I415819,I415553);
DFFARX1 I_24292 (I415827,I2859,I415369,I415340,);
nand I_24293 (I415858,I415819,I415460);
nand I_24294 (I415875,I415553,I415858);
nor I_24295 (I415349,I415875,I415519);
not I_24296 (I415930,I2866);
DFFARX1 I_24297 (I194704,I2859,I415930,I415956,);
DFFARX1 I_24298 (I415956,I2859,I415930,I415973,);
not I_24299 (I415922,I415973);
not I_24300 (I415995,I415956);
DFFARX1 I_24301 (I194692,I2859,I415930,I416021,);
nand I_24302 (I416029,I416021,I194698);
not I_24303 (I416046,I194698);
not I_24304 (I416063,I194695);
nand I_24305 (I416080,I194683,I194680);
and I_24306 (I416097,I194683,I194680);
not I_24307 (I416114,I194707);
nand I_24308 (I416131,I416114,I416063);
nor I_24309 (I415904,I416131,I416029);
nor I_24310 (I416162,I416046,I416131);
nand I_24311 (I415907,I416097,I416162);
not I_24312 (I416193,I194680);
nor I_24313 (I416210,I416193,I194683);
nor I_24314 (I416227,I416210,I194707);
nor I_24315 (I416244,I415995,I416227);
DFFARX1 I_24316 (I416244,I2859,I415930,I415916,);
not I_24317 (I416275,I416210);
DFFARX1 I_24318 (I416275,I2859,I415930,I415919,);
and I_24319 (I415913,I416021,I416210);
nor I_24320 (I416320,I416193,I194689);
and I_24321 (I416337,I416320,I194686);
or I_24322 (I416354,I416337,I194701);
DFFARX1 I_24323 (I416354,I2859,I415930,I416380,);
nor I_24324 (I416388,I416380,I416114);
DFFARX1 I_24325 (I416388,I2859,I415930,I415901,);
nand I_24326 (I416419,I416380,I416021);
nand I_24327 (I416436,I416114,I416419);
nor I_24328 (I415910,I416436,I416080);
not I_24329 (I416491,I2866);
DFFARX1 I_24330 (I293793,I2859,I416491,I416517,);
DFFARX1 I_24331 (I416517,I2859,I416491,I416534,);
not I_24332 (I416483,I416534);
not I_24333 (I416556,I416517);
DFFARX1 I_24334 (I293805,I2859,I416491,I416582,);
nand I_24335 (I416590,I416582,I293814);
not I_24336 (I416607,I293814);
not I_24337 (I416624,I293796);
nand I_24338 (I416641,I293799,I293790);
and I_24339 (I416658,I293799,I293790);
not I_24340 (I416675,I293808);
nand I_24341 (I416692,I416675,I416624);
nor I_24342 (I416465,I416692,I416590);
nor I_24343 (I416723,I416607,I416692);
nand I_24344 (I416468,I416658,I416723);
not I_24345 (I416754,I293811);
nor I_24346 (I416771,I416754,I293799);
nor I_24347 (I416788,I416771,I293808);
nor I_24348 (I416805,I416556,I416788);
DFFARX1 I_24349 (I416805,I2859,I416491,I416477,);
not I_24350 (I416836,I416771);
DFFARX1 I_24351 (I416836,I2859,I416491,I416480,);
and I_24352 (I416474,I416582,I416771);
nor I_24353 (I416881,I416754,I293790);
and I_24354 (I416898,I416881,I293802);
or I_24355 (I416915,I416898,I293793);
DFFARX1 I_24356 (I416915,I2859,I416491,I416941,);
nor I_24357 (I416949,I416941,I416675);
DFFARX1 I_24358 (I416949,I2859,I416491,I416462,);
nand I_24359 (I416980,I416941,I416582);
nand I_24360 (I416997,I416675,I416980);
nor I_24361 (I416471,I416997,I416641);
not I_24362 (I417052,I2866);
DFFARX1 I_24363 (I342317,I2859,I417052,I417078,);
DFFARX1 I_24364 (I417078,I2859,I417052,I417095,);
not I_24365 (I417044,I417095);
not I_24366 (I417117,I417078);
DFFARX1 I_24367 (I342314,I2859,I417052,I417143,);
nand I_24368 (I417151,I417143,I342329);
not I_24369 (I417168,I342329);
not I_24370 (I417185,I342326);
nand I_24371 (I417202,I342323,I342311);
and I_24372 (I417219,I342323,I342311);
not I_24373 (I417236,I342308);
nand I_24374 (I417253,I417236,I417185);
nor I_24375 (I417026,I417253,I417151);
nor I_24376 (I417284,I417168,I417253);
nand I_24377 (I417029,I417219,I417284);
not I_24378 (I417315,I342314);
nor I_24379 (I417332,I417315,I342323);
nor I_24380 (I417349,I417332,I342308);
nor I_24381 (I417366,I417117,I417349);
DFFARX1 I_24382 (I417366,I2859,I417052,I417038,);
not I_24383 (I417397,I417332);
DFFARX1 I_24384 (I417397,I2859,I417052,I417041,);
and I_24385 (I417035,I417143,I417332);
nor I_24386 (I417442,I417315,I342320);
and I_24387 (I417459,I417442,I342308);
or I_24388 (I417476,I417459,I342311);
DFFARX1 I_24389 (I417476,I2859,I417052,I417502,);
nor I_24390 (I417510,I417502,I417236);
DFFARX1 I_24391 (I417510,I2859,I417052,I417023,);
nand I_24392 (I417541,I417502,I417143);
nand I_24393 (I417558,I417236,I417541);
nor I_24394 (I417032,I417558,I417202);
not I_24395 (I417613,I2866);
DFFARX1 I_24396 (I560620,I2859,I417613,I417639,);
DFFARX1 I_24397 (I417639,I2859,I417613,I417656,);
not I_24398 (I417605,I417656);
not I_24399 (I417678,I417639);
DFFARX1 I_24400 (I560614,I2859,I417613,I417704,);
nand I_24401 (I417712,I417704,I560605);
not I_24402 (I417729,I560605);
not I_24403 (I417746,I560632);
nand I_24404 (I417763,I560617,I560626);
and I_24405 (I417780,I560617,I560626);
not I_24406 (I417797,I560611);
nand I_24407 (I417814,I417797,I417746);
nor I_24408 (I417587,I417814,I417712);
nor I_24409 (I417845,I417729,I417814);
nand I_24410 (I417590,I417780,I417845);
not I_24411 (I417876,I560629);
nor I_24412 (I417893,I417876,I560617);
nor I_24413 (I417910,I417893,I560611);
nor I_24414 (I417927,I417678,I417910);
DFFARX1 I_24415 (I417927,I2859,I417613,I417599,);
not I_24416 (I417958,I417893);
DFFARX1 I_24417 (I417958,I2859,I417613,I417602,);
and I_24418 (I417596,I417704,I417893);
nor I_24419 (I418003,I417876,I560623);
and I_24420 (I418020,I418003,I560605);
or I_24421 (I418037,I418020,I560608);
DFFARX1 I_24422 (I418037,I2859,I417613,I418063,);
nor I_24423 (I418071,I418063,I417797);
DFFARX1 I_24424 (I418071,I2859,I417613,I417584,);
nand I_24425 (I418102,I418063,I417704);
nand I_24426 (I418119,I417797,I418102);
nor I_24427 (I417593,I418119,I417763);
not I_24428 (I418174,I2866);
DFFARX1 I_24429 (I124066,I2859,I418174,I418200,);
DFFARX1 I_24430 (I418200,I2859,I418174,I418217,);
not I_24431 (I418166,I418217);
not I_24432 (I418239,I418200);
DFFARX1 I_24433 (I124063,I2859,I418174,I418265,);
nand I_24434 (I418273,I418265,I124057);
not I_24435 (I418290,I124057);
not I_24436 (I418307,I124054);
nand I_24437 (I418324,I124048,I124045);
and I_24438 (I418341,I124048,I124045);
not I_24439 (I418358,I124060);
nand I_24440 (I418375,I418358,I418307);
nor I_24441 (I418148,I418375,I418273);
nor I_24442 (I418406,I418290,I418375);
nand I_24443 (I418151,I418341,I418406);
not I_24444 (I418437,I124072);
nor I_24445 (I418454,I418437,I124048);
nor I_24446 (I418471,I418454,I124060);
nor I_24447 (I418488,I418239,I418471);
DFFARX1 I_24448 (I418488,I2859,I418174,I418160,);
not I_24449 (I418519,I418454);
DFFARX1 I_24450 (I418519,I2859,I418174,I418163,);
and I_24451 (I418157,I418265,I418454);
nor I_24452 (I418564,I418437,I124069);
and I_24453 (I418581,I418564,I124045);
or I_24454 (I418598,I418581,I124051);
DFFARX1 I_24455 (I418598,I2859,I418174,I418624,);
nor I_24456 (I418632,I418624,I418358);
DFFARX1 I_24457 (I418632,I2859,I418174,I418145,);
nand I_24458 (I418663,I418624,I418265);
nand I_24459 (I418680,I418358,I418663);
nor I_24460 (I418154,I418680,I418324);
not I_24461 (I418735,I2866);
DFFARX1 I_24462 (I156213,I2859,I418735,I418761,);
DFFARX1 I_24463 (I418761,I2859,I418735,I418778,);
not I_24464 (I418727,I418778);
not I_24465 (I418800,I418761);
DFFARX1 I_24466 (I156210,I2859,I418735,I418826,);
nand I_24467 (I418834,I418826,I156204);
not I_24468 (I418851,I156204);
not I_24469 (I418868,I156201);
nand I_24470 (I418885,I156195,I156192);
and I_24471 (I418902,I156195,I156192);
not I_24472 (I418919,I156207);
nand I_24473 (I418936,I418919,I418868);
nor I_24474 (I418709,I418936,I418834);
nor I_24475 (I418967,I418851,I418936);
nand I_24476 (I418712,I418902,I418967);
not I_24477 (I418998,I156219);
nor I_24478 (I419015,I418998,I156195);
nor I_24479 (I419032,I419015,I156207);
nor I_24480 (I419049,I418800,I419032);
DFFARX1 I_24481 (I419049,I2859,I418735,I418721,);
not I_24482 (I419080,I419015);
DFFARX1 I_24483 (I419080,I2859,I418735,I418724,);
and I_24484 (I418718,I418826,I419015);
nor I_24485 (I419125,I418998,I156216);
and I_24486 (I419142,I419125,I156192);
or I_24487 (I419159,I419142,I156198);
DFFARX1 I_24488 (I419159,I2859,I418735,I419185,);
nor I_24489 (I419193,I419185,I418919);
DFFARX1 I_24490 (I419193,I2859,I418735,I418706,);
nand I_24491 (I419224,I419185,I418826);
nand I_24492 (I419241,I418919,I419224);
nor I_24493 (I418715,I419241,I418885);
not I_24494 (I419296,I2866);
DFFARX1 I_24495 (I186544,I2859,I419296,I419322,);
DFFARX1 I_24496 (I419322,I2859,I419296,I419339,);
not I_24497 (I419288,I419339);
not I_24498 (I419361,I419322);
DFFARX1 I_24499 (I186532,I2859,I419296,I419387,);
nand I_24500 (I419395,I419387,I186538);
not I_24501 (I419412,I186538);
not I_24502 (I419429,I186535);
nand I_24503 (I419446,I186523,I186520);
and I_24504 (I419463,I186523,I186520);
not I_24505 (I419480,I186547);
nand I_24506 (I419497,I419480,I419429);
nor I_24507 (I419270,I419497,I419395);
nor I_24508 (I419528,I419412,I419497);
nand I_24509 (I419273,I419463,I419528);
not I_24510 (I419559,I186520);
nor I_24511 (I419576,I419559,I186523);
nor I_24512 (I419593,I419576,I186547);
nor I_24513 (I419610,I419361,I419593);
DFFARX1 I_24514 (I419610,I2859,I419296,I419282,);
not I_24515 (I419641,I419576);
DFFARX1 I_24516 (I419641,I2859,I419296,I419285,);
and I_24517 (I419279,I419387,I419576);
nor I_24518 (I419686,I419559,I186529);
and I_24519 (I419703,I419686,I186526);
or I_24520 (I419720,I419703,I186541);
DFFARX1 I_24521 (I419720,I2859,I419296,I419746,);
nor I_24522 (I419754,I419746,I419480);
DFFARX1 I_24523 (I419754,I2859,I419296,I419267,);
nand I_24524 (I419785,I419746,I419387);
nand I_24525 (I419802,I419480,I419785);
nor I_24526 (I419276,I419802,I419446);
not I_24527 (I419857,I2866);
DFFARX1 I_24528 (I459147,I2859,I419857,I419883,);
DFFARX1 I_24529 (I419883,I2859,I419857,I419900,);
not I_24530 (I419849,I419900);
not I_24531 (I419922,I419883);
DFFARX1 I_24532 (I459138,I2859,I419857,I419948,);
nand I_24533 (I419956,I419948,I459135);
not I_24534 (I419973,I459135);
not I_24535 (I419990,I459144);
nand I_24536 (I420007,I459153,I459135);
and I_24537 (I420024,I459153,I459135);
not I_24538 (I420041,I459132);
nand I_24539 (I420058,I420041,I419990);
nor I_24540 (I419831,I420058,I419956);
nor I_24541 (I420089,I419973,I420058);
nand I_24542 (I419834,I420024,I420089);
not I_24543 (I420120,I459141);
nor I_24544 (I420137,I420120,I459153);
nor I_24545 (I420154,I420137,I459132);
nor I_24546 (I420171,I419922,I420154);
DFFARX1 I_24547 (I420171,I2859,I419857,I419843,);
not I_24548 (I420202,I420137);
DFFARX1 I_24549 (I420202,I2859,I419857,I419846,);
and I_24550 (I419840,I419948,I420137);
nor I_24551 (I420247,I420120,I459156);
and I_24552 (I420264,I420247,I459132);
or I_24553 (I420281,I420264,I459150);
DFFARX1 I_24554 (I420281,I2859,I419857,I420307,);
nor I_24555 (I420315,I420307,I420041);
DFFARX1 I_24556 (I420315,I2859,I419857,I419828,);
nand I_24557 (I420346,I420307,I419948);
nand I_24558 (I420363,I420041,I420346);
nor I_24559 (I419837,I420363,I420007);
not I_24560 (I420418,I2866);
DFFARX1 I_24561 (I151997,I2859,I420418,I420444,);
DFFARX1 I_24562 (I420444,I2859,I420418,I420461,);
not I_24563 (I420410,I420461);
not I_24564 (I420483,I420444);
DFFARX1 I_24565 (I151994,I2859,I420418,I420509,);
nand I_24566 (I420517,I420509,I151988);
not I_24567 (I420534,I151988);
not I_24568 (I420551,I151985);
nand I_24569 (I420568,I151979,I151976);
and I_24570 (I420585,I151979,I151976);
not I_24571 (I420602,I151991);
nand I_24572 (I420619,I420602,I420551);
nor I_24573 (I420392,I420619,I420517);
nor I_24574 (I420650,I420534,I420619);
nand I_24575 (I420395,I420585,I420650);
not I_24576 (I420681,I152003);
nor I_24577 (I420698,I420681,I151979);
nor I_24578 (I420715,I420698,I151991);
nor I_24579 (I420732,I420483,I420715);
DFFARX1 I_24580 (I420732,I2859,I420418,I420404,);
not I_24581 (I420763,I420698);
DFFARX1 I_24582 (I420763,I2859,I420418,I420407,);
and I_24583 (I420401,I420509,I420698);
nor I_24584 (I420808,I420681,I152000);
and I_24585 (I420825,I420808,I151976);
or I_24586 (I420842,I420825,I151982);
DFFARX1 I_24587 (I420842,I2859,I420418,I420868,);
nor I_24588 (I420876,I420868,I420602);
DFFARX1 I_24589 (I420876,I2859,I420418,I420389,);
nand I_24590 (I420907,I420868,I420509);
nand I_24591 (I420924,I420602,I420907);
nor I_24592 (I420398,I420924,I420568);
not I_24593 (I420979,I2866);
DFFARX1 I_24594 (I464927,I2859,I420979,I421005,);
DFFARX1 I_24595 (I421005,I2859,I420979,I421022,);
not I_24596 (I420971,I421022);
not I_24597 (I421044,I421005);
DFFARX1 I_24598 (I464918,I2859,I420979,I421070,);
nand I_24599 (I421078,I421070,I464915);
not I_24600 (I421095,I464915);
not I_24601 (I421112,I464924);
nand I_24602 (I421129,I464933,I464915);
and I_24603 (I421146,I464933,I464915);
not I_24604 (I421163,I464912);
nand I_24605 (I421180,I421163,I421112);
nor I_24606 (I420953,I421180,I421078);
nor I_24607 (I421211,I421095,I421180);
nand I_24608 (I420956,I421146,I421211);
not I_24609 (I421242,I464921);
nor I_24610 (I421259,I421242,I464933);
nor I_24611 (I421276,I421259,I464912);
nor I_24612 (I421293,I421044,I421276);
DFFARX1 I_24613 (I421293,I2859,I420979,I420965,);
not I_24614 (I421324,I421259);
DFFARX1 I_24615 (I421324,I2859,I420979,I420968,);
and I_24616 (I420962,I421070,I421259);
nor I_24617 (I421369,I421242,I464936);
and I_24618 (I421386,I421369,I464912);
or I_24619 (I421403,I421386,I464930);
DFFARX1 I_24620 (I421403,I2859,I420979,I421429,);
nor I_24621 (I421437,I421429,I421163);
DFFARX1 I_24622 (I421437,I2859,I420979,I420950,);
nand I_24623 (I421468,I421429,I421070);
nand I_24624 (I421485,I421163,I421468);
nor I_24625 (I420959,I421485,I421129);
not I_24626 (I421540,I2866);
DFFARX1 I_24627 (I215013,I2859,I421540,I421566,);
DFFARX1 I_24628 (I421566,I2859,I421540,I421583,);
not I_24629 (I421532,I421583);
not I_24630 (I421605,I421566);
DFFARX1 I_24631 (I215010,I2859,I421540,I421631,);
nand I_24632 (I421639,I421631,I215004);
not I_24633 (I421656,I215004);
not I_24634 (I421673,I215016);
nand I_24635 (I421690,I215019,I214998);
and I_24636 (I421707,I215019,I214998);
not I_24637 (I421724,I214995);
nand I_24638 (I421741,I421724,I421673);
nor I_24639 (I421514,I421741,I421639);
nor I_24640 (I421772,I421656,I421741);
nand I_24641 (I421517,I421707,I421772);
not I_24642 (I421803,I215001);
nor I_24643 (I421820,I421803,I215019);
nor I_24644 (I421837,I421820,I214995);
nor I_24645 (I421854,I421605,I421837);
DFFARX1 I_24646 (I421854,I2859,I421540,I421526,);
not I_24647 (I421885,I421820);
DFFARX1 I_24648 (I421885,I2859,I421540,I421529,);
and I_24649 (I421523,I421631,I421820);
nor I_24650 (I421930,I421803,I214995);
and I_24651 (I421947,I421930,I215007);
or I_24652 (I421964,I421947,I214998);
DFFARX1 I_24653 (I421964,I2859,I421540,I421990,);
nor I_24654 (I421998,I421990,I421724);
DFFARX1 I_24655 (I421998,I2859,I421540,I421511,);
nand I_24656 (I422029,I421990,I421631);
nand I_24657 (I422046,I421724,I422029);
nor I_24658 (I421520,I422046,I421690);
not I_24659 (I422101,I2866);
DFFARX1 I_24660 (I149362,I2859,I422101,I422127,);
DFFARX1 I_24661 (I422127,I2859,I422101,I422144,);
not I_24662 (I422093,I422144);
not I_24663 (I422166,I422127);
DFFARX1 I_24664 (I149359,I2859,I422101,I422192,);
nand I_24665 (I422200,I422192,I149353);
not I_24666 (I422217,I149353);
not I_24667 (I422234,I149350);
nand I_24668 (I422251,I149344,I149341);
and I_24669 (I422268,I149344,I149341);
not I_24670 (I422285,I149356);
nand I_24671 (I422302,I422285,I422234);
nor I_24672 (I422075,I422302,I422200);
nor I_24673 (I422333,I422217,I422302);
nand I_24674 (I422078,I422268,I422333);
not I_24675 (I422364,I149368);
nor I_24676 (I422381,I422364,I149344);
nor I_24677 (I422398,I422381,I149356);
nor I_24678 (I422415,I422166,I422398);
DFFARX1 I_24679 (I422415,I2859,I422101,I422087,);
not I_24680 (I422446,I422381);
DFFARX1 I_24681 (I422446,I2859,I422101,I422090,);
and I_24682 (I422084,I422192,I422381);
nor I_24683 (I422491,I422364,I149365);
and I_24684 (I422508,I422491,I149341);
or I_24685 (I422525,I422508,I149347);
DFFARX1 I_24686 (I422525,I2859,I422101,I422551,);
nor I_24687 (I422559,I422551,I422285);
DFFARX1 I_24688 (I422559,I2859,I422101,I422072,);
nand I_24689 (I422590,I422551,I422192);
nand I_24690 (I422607,I422285,I422590);
nor I_24691 (I422081,I422607,I422251);
not I_24692 (I422662,I2866);
DFFARX1 I_24693 (I401213,I2859,I422662,I422688,);
DFFARX1 I_24694 (I422688,I2859,I422662,I422705,);
not I_24695 (I422654,I422705);
not I_24696 (I422727,I422688);
DFFARX1 I_24697 (I401240,I2859,I422662,I422753,);
nand I_24698 (I422761,I422753,I401231);
not I_24699 (I422778,I401231);
not I_24700 (I422795,I401213);
nand I_24701 (I422812,I401225,I401228);
and I_24702 (I422829,I401225,I401228);
not I_24703 (I422846,I401237);
nand I_24704 (I422863,I422846,I422795);
nor I_24705 (I422636,I422863,I422761);
nor I_24706 (I422894,I422778,I422863);
nand I_24707 (I422639,I422829,I422894);
not I_24708 (I422925,I401222);
nor I_24709 (I422942,I422925,I401225);
nor I_24710 (I422959,I422942,I401237);
nor I_24711 (I422976,I422727,I422959);
DFFARX1 I_24712 (I422976,I2859,I422662,I422648,);
not I_24713 (I423007,I422942);
DFFARX1 I_24714 (I423007,I2859,I422662,I422651,);
and I_24715 (I422645,I422753,I422942);
nor I_24716 (I423052,I422925,I401216);
and I_24717 (I423069,I423052,I401219);
or I_24718 (I423086,I423069,I401234);
DFFARX1 I_24719 (I423086,I2859,I422662,I423112,);
nor I_24720 (I423120,I423112,I422846);
DFFARX1 I_24721 (I423120,I2859,I422662,I422633,);
nand I_24722 (I423151,I423112,I422753);
nand I_24723 (I423168,I422846,I423151);
nor I_24724 (I422642,I423168,I422812);
not I_24725 (I423223,I2866);
DFFARX1 I_24726 (I482845,I2859,I423223,I423249,);
DFFARX1 I_24727 (I423249,I2859,I423223,I423266,);
not I_24728 (I423215,I423266);
not I_24729 (I423288,I423249);
DFFARX1 I_24730 (I482836,I2859,I423223,I423314,);
nand I_24731 (I423322,I423314,I482833);
not I_24732 (I423339,I482833);
not I_24733 (I423356,I482842);
nand I_24734 (I423373,I482851,I482833);
and I_24735 (I423390,I482851,I482833);
not I_24736 (I423407,I482830);
nand I_24737 (I423424,I423407,I423356);
nor I_24738 (I423197,I423424,I423322);
nor I_24739 (I423455,I423339,I423424);
nand I_24740 (I423200,I423390,I423455);
not I_24741 (I423486,I482839);
nor I_24742 (I423503,I423486,I482851);
nor I_24743 (I423520,I423503,I482830);
nor I_24744 (I423537,I423288,I423520);
DFFARX1 I_24745 (I423537,I2859,I423223,I423209,);
not I_24746 (I423568,I423503);
DFFARX1 I_24747 (I423568,I2859,I423223,I423212,);
and I_24748 (I423206,I423314,I423503);
nor I_24749 (I423613,I423486,I482854);
and I_24750 (I423630,I423613,I482830);
or I_24751 (I423647,I423630,I482848);
DFFARX1 I_24752 (I423647,I2859,I423223,I423673,);
nor I_24753 (I423681,I423673,I423407);
DFFARX1 I_24754 (I423681,I2859,I423223,I423194,);
nand I_24755 (I423712,I423673,I423314);
nand I_24756 (I423729,I423407,I423712);
nor I_24757 (I423203,I423729,I423373);
not I_24758 (I423784,I2866);
DFFARX1 I_24759 (I190352,I2859,I423784,I423810,);
DFFARX1 I_24760 (I423810,I2859,I423784,I423827,);
not I_24761 (I423776,I423827);
not I_24762 (I423849,I423810);
DFFARX1 I_24763 (I190340,I2859,I423784,I423875,);
nand I_24764 (I423883,I423875,I190346);
not I_24765 (I423900,I190346);
not I_24766 (I423917,I190343);
nand I_24767 (I423934,I190331,I190328);
and I_24768 (I423951,I190331,I190328);
not I_24769 (I423968,I190355);
nand I_24770 (I423985,I423968,I423917);
nor I_24771 (I423758,I423985,I423883);
nor I_24772 (I424016,I423900,I423985);
nand I_24773 (I423761,I423951,I424016);
not I_24774 (I424047,I190328);
nor I_24775 (I424064,I424047,I190331);
nor I_24776 (I424081,I424064,I190355);
nor I_24777 (I424098,I423849,I424081);
DFFARX1 I_24778 (I424098,I2859,I423784,I423770,);
not I_24779 (I424129,I424064);
DFFARX1 I_24780 (I424129,I2859,I423784,I423773,);
and I_24781 (I423767,I423875,I424064);
nor I_24782 (I424174,I424047,I190337);
and I_24783 (I424191,I424174,I190334);
or I_24784 (I424208,I424191,I190349);
DFFARX1 I_24785 (I424208,I2859,I423784,I424234,);
nor I_24786 (I424242,I424234,I423968);
DFFARX1 I_24787 (I424242,I2859,I423784,I423755,);
nand I_24788 (I424273,I424234,I423875);
nand I_24789 (I424290,I423968,I424273);
nor I_24790 (I423764,I424290,I423934);
not I_24791 (I424345,I2866);
DFFARX1 I_24792 (I491515,I2859,I424345,I424371,);
DFFARX1 I_24793 (I424371,I2859,I424345,I424388,);
not I_24794 (I424337,I424388);
not I_24795 (I424410,I424371);
DFFARX1 I_24796 (I491506,I2859,I424345,I424436,);
nand I_24797 (I424444,I424436,I491503);
not I_24798 (I424461,I491503);
not I_24799 (I424478,I491512);
nand I_24800 (I424495,I491521,I491503);
and I_24801 (I424512,I491521,I491503);
not I_24802 (I424529,I491500);
nand I_24803 (I424546,I424529,I424478);
nor I_24804 (I424319,I424546,I424444);
nor I_24805 (I424577,I424461,I424546);
nand I_24806 (I424322,I424512,I424577);
not I_24807 (I424608,I491509);
nor I_24808 (I424625,I424608,I491521);
nor I_24809 (I424642,I424625,I491500);
nor I_24810 (I424659,I424410,I424642);
DFFARX1 I_24811 (I424659,I2859,I424345,I424331,);
not I_24812 (I424690,I424625);
DFFARX1 I_24813 (I424690,I2859,I424345,I424334,);
and I_24814 (I424328,I424436,I424625);
nor I_24815 (I424735,I424608,I491524);
and I_24816 (I424752,I424735,I491500);
or I_24817 (I424769,I424752,I491518);
DFFARX1 I_24818 (I424769,I2859,I424345,I424795,);
nor I_24819 (I424803,I424795,I424529);
DFFARX1 I_24820 (I424803,I2859,I424345,I424316,);
nand I_24821 (I424834,I424795,I424436);
nand I_24822 (I424851,I424529,I424834);
nor I_24823 (I424325,I424851,I424495);
not I_24824 (I424906,I2866);
DFFARX1 I_24825 (I130917,I2859,I424906,I424932,);
DFFARX1 I_24826 (I424932,I2859,I424906,I424949,);
not I_24827 (I424898,I424949);
not I_24828 (I424971,I424932);
DFFARX1 I_24829 (I130914,I2859,I424906,I424997,);
nand I_24830 (I425005,I424997,I130908);
not I_24831 (I425022,I130908);
not I_24832 (I425039,I130905);
nand I_24833 (I425056,I130899,I130896);
and I_24834 (I425073,I130899,I130896);
not I_24835 (I425090,I130911);
nand I_24836 (I425107,I425090,I425039);
nor I_24837 (I424880,I425107,I425005);
nor I_24838 (I425138,I425022,I425107);
nand I_24839 (I424883,I425073,I425138);
not I_24840 (I425169,I130923);
nor I_24841 (I425186,I425169,I130899);
nor I_24842 (I425203,I425186,I130911);
nor I_24843 (I425220,I424971,I425203);
DFFARX1 I_24844 (I425220,I2859,I424906,I424892,);
not I_24845 (I425251,I425186);
DFFARX1 I_24846 (I425251,I2859,I424906,I424895,);
and I_24847 (I424889,I424997,I425186);
nor I_24848 (I425296,I425169,I130920);
and I_24849 (I425313,I425296,I130896);
or I_24850 (I425330,I425313,I130902);
DFFARX1 I_24851 (I425330,I2859,I424906,I425356,);
nor I_24852 (I425364,I425356,I425090);
DFFARX1 I_24853 (I425364,I2859,I424906,I424877,);
nand I_24854 (I425395,I425356,I424997);
nand I_24855 (I425412,I425090,I425395);
nor I_24856 (I424886,I425412,I425056);
not I_24857 (I425467,I2866);
DFFARX1 I_24858 (I354965,I2859,I425467,I425493,);
DFFARX1 I_24859 (I425493,I2859,I425467,I425510,);
not I_24860 (I425459,I425510);
not I_24861 (I425532,I425493);
DFFARX1 I_24862 (I354962,I2859,I425467,I425558,);
nand I_24863 (I425566,I425558,I354977);
not I_24864 (I425583,I354977);
not I_24865 (I425600,I354974);
nand I_24866 (I425617,I354971,I354959);
and I_24867 (I425634,I354971,I354959);
not I_24868 (I425651,I354956);
nand I_24869 (I425668,I425651,I425600);
nor I_24870 (I425441,I425668,I425566);
nor I_24871 (I425699,I425583,I425668);
nand I_24872 (I425444,I425634,I425699);
not I_24873 (I425730,I354962);
nor I_24874 (I425747,I425730,I354971);
nor I_24875 (I425764,I425747,I354956);
nor I_24876 (I425781,I425532,I425764);
DFFARX1 I_24877 (I425781,I2859,I425467,I425453,);
not I_24878 (I425812,I425747);
DFFARX1 I_24879 (I425812,I2859,I425467,I425456,);
and I_24880 (I425450,I425558,I425747);
nor I_24881 (I425857,I425730,I354968);
and I_24882 (I425874,I425857,I354956);
or I_24883 (I425891,I425874,I354959);
DFFARX1 I_24884 (I425891,I2859,I425467,I425917,);
nor I_24885 (I425925,I425917,I425651);
DFFARX1 I_24886 (I425925,I2859,I425467,I425438,);
nand I_24887 (I425956,I425917,I425558);
nand I_24888 (I425973,I425651,I425956);
nor I_24889 (I425447,I425973,I425617);
not I_24890 (I426028,I2866);
DFFARX1 I_24891 (I344425,I2859,I426028,I426054,);
DFFARX1 I_24892 (I426054,I2859,I426028,I426071,);
not I_24893 (I426020,I426071);
not I_24894 (I426093,I426054);
DFFARX1 I_24895 (I344422,I2859,I426028,I426119,);
nand I_24896 (I426127,I426119,I344437);
not I_24897 (I426144,I344437);
not I_24898 (I426161,I344434);
nand I_24899 (I426178,I344431,I344419);
and I_24900 (I426195,I344431,I344419);
not I_24901 (I426212,I344416);
nand I_24902 (I426229,I426212,I426161);
nor I_24903 (I426002,I426229,I426127);
nor I_24904 (I426260,I426144,I426229);
nand I_24905 (I426005,I426195,I426260);
not I_24906 (I426291,I344422);
nor I_24907 (I426308,I426291,I344431);
nor I_24908 (I426325,I426308,I344416);
nor I_24909 (I426342,I426093,I426325);
DFFARX1 I_24910 (I426342,I2859,I426028,I426014,);
not I_24911 (I426373,I426308);
DFFARX1 I_24912 (I426373,I2859,I426028,I426017,);
and I_24913 (I426011,I426119,I426308);
nor I_24914 (I426418,I426291,I344428);
and I_24915 (I426435,I426418,I344416);
or I_24916 (I426452,I426435,I344419);
DFFARX1 I_24917 (I426452,I2859,I426028,I426478,);
nor I_24918 (I426486,I426478,I426212);
DFFARX1 I_24919 (I426486,I2859,I426028,I425999,);
nand I_24920 (I426517,I426478,I426119);
nand I_24921 (I426534,I426212,I426517);
nor I_24922 (I426008,I426534,I426178);
not I_24923 (I426589,I2866);
DFFARX1 I_24924 (I304197,I2859,I426589,I426615,);
DFFARX1 I_24925 (I426615,I2859,I426589,I426632,);
not I_24926 (I426581,I426632);
not I_24927 (I426654,I426615);
DFFARX1 I_24928 (I304209,I2859,I426589,I426680,);
nand I_24929 (I426688,I426680,I304218);
not I_24930 (I426705,I304218);
not I_24931 (I426722,I304200);
nand I_24932 (I426739,I304203,I304194);
and I_24933 (I426756,I304203,I304194);
not I_24934 (I426773,I304212);
nand I_24935 (I426790,I426773,I426722);
nor I_24936 (I426563,I426790,I426688);
nor I_24937 (I426821,I426705,I426790);
nand I_24938 (I426566,I426756,I426821);
not I_24939 (I426852,I304215);
nor I_24940 (I426869,I426852,I304203);
nor I_24941 (I426886,I426869,I304212);
nor I_24942 (I426903,I426654,I426886);
DFFARX1 I_24943 (I426903,I2859,I426589,I426575,);
not I_24944 (I426934,I426869);
DFFARX1 I_24945 (I426934,I2859,I426589,I426578,);
and I_24946 (I426572,I426680,I426869);
nor I_24947 (I426979,I426852,I304194);
and I_24948 (I426996,I426979,I304206);
or I_24949 (I427013,I426996,I304197);
DFFARX1 I_24950 (I427013,I2859,I426589,I427039,);
nor I_24951 (I427047,I427039,I426773);
DFFARX1 I_24952 (I427047,I2859,I426589,I426560,);
nand I_24953 (I427078,I427039,I426680);
nand I_24954 (I427095,I426773,I427078);
nor I_24955 (I426569,I427095,I426739);
not I_24956 (I427150,I2866);
DFFARX1 I_24957 (I452789,I2859,I427150,I427176,);
DFFARX1 I_24958 (I427176,I2859,I427150,I427193,);
not I_24959 (I427142,I427193);
not I_24960 (I427215,I427176);
DFFARX1 I_24961 (I452780,I2859,I427150,I427241,);
nand I_24962 (I427249,I427241,I452777);
not I_24963 (I427266,I452777);
not I_24964 (I427283,I452786);
nand I_24965 (I427300,I452795,I452777);
and I_24966 (I427317,I452795,I452777);
not I_24967 (I427334,I452774);
nand I_24968 (I427351,I427334,I427283);
nor I_24969 (I427124,I427351,I427249);
nor I_24970 (I427382,I427266,I427351);
nand I_24971 (I427127,I427317,I427382);
not I_24972 (I427413,I452783);
nor I_24973 (I427430,I427413,I452795);
nor I_24974 (I427447,I427430,I452774);
nor I_24975 (I427464,I427215,I427447);
DFFARX1 I_24976 (I427464,I2859,I427150,I427136,);
not I_24977 (I427495,I427430);
DFFARX1 I_24978 (I427495,I2859,I427150,I427139,);
and I_24979 (I427133,I427241,I427430);
nor I_24980 (I427540,I427413,I452798);
and I_24981 (I427557,I427540,I452774);
or I_24982 (I427574,I427557,I452792);
DFFARX1 I_24983 (I427574,I2859,I427150,I427600,);
nor I_24984 (I427608,I427600,I427334);
DFFARX1 I_24985 (I427608,I2859,I427150,I427121,);
nand I_24986 (I427639,I427600,I427241);
nand I_24987 (I427656,I427334,I427639);
nor I_24988 (I427130,I427656,I427300);
not I_24989 (I427711,I2866);
DFFARX1 I_24990 (I485157,I2859,I427711,I427737,);
DFFARX1 I_24991 (I427737,I2859,I427711,I427754,);
not I_24992 (I427703,I427754);
not I_24993 (I427776,I427737);
DFFARX1 I_24994 (I485148,I2859,I427711,I427802,);
nand I_24995 (I427810,I427802,I485145);
not I_24996 (I427827,I485145);
not I_24997 (I427844,I485154);
nand I_24998 (I427861,I485163,I485145);
and I_24999 (I427878,I485163,I485145);
not I_25000 (I427895,I485142);
nand I_25001 (I427912,I427895,I427844);
nor I_25002 (I427685,I427912,I427810);
nor I_25003 (I427943,I427827,I427912);
nand I_25004 (I427688,I427878,I427943);
not I_25005 (I427974,I485151);
nor I_25006 (I427991,I427974,I485163);
nor I_25007 (I428008,I427991,I485142);
nor I_25008 (I428025,I427776,I428008);
DFFARX1 I_25009 (I428025,I2859,I427711,I427697,);
not I_25010 (I428056,I427991);
DFFARX1 I_25011 (I428056,I2859,I427711,I427700,);
and I_25012 (I427694,I427802,I427991);
nor I_25013 (I428101,I427974,I485166);
and I_25014 (I428118,I428101,I485142);
or I_25015 (I428135,I428118,I485160);
DFFARX1 I_25016 (I428135,I2859,I427711,I428161,);
nor I_25017 (I428169,I428161,I427895);
DFFARX1 I_25018 (I428169,I2859,I427711,I427682,);
nand I_25019 (I428200,I428161,I427802);
nand I_25020 (I428217,I427895,I428200);
nor I_25021 (I427691,I428217,I427861);
not I_25022 (I428272,I2866);
DFFARX1 I_25023 (I355492,I2859,I428272,I428298,);
DFFARX1 I_25024 (I428298,I2859,I428272,I428315,);
not I_25025 (I428264,I428315);
not I_25026 (I428337,I428298);
DFFARX1 I_25027 (I355489,I2859,I428272,I428363,);
nand I_25028 (I428371,I428363,I355504);
not I_25029 (I428388,I355504);
not I_25030 (I428405,I355501);
nand I_25031 (I428422,I355498,I355486);
and I_25032 (I428439,I355498,I355486);
not I_25033 (I428456,I355483);
nand I_25034 (I428473,I428456,I428405);
nor I_25035 (I428246,I428473,I428371);
nor I_25036 (I428504,I428388,I428473);
nand I_25037 (I428249,I428439,I428504);
not I_25038 (I428535,I355489);
nor I_25039 (I428552,I428535,I355498);
nor I_25040 (I428569,I428552,I355483);
nor I_25041 (I428586,I428337,I428569);
DFFARX1 I_25042 (I428586,I2859,I428272,I428258,);
not I_25043 (I428617,I428552);
DFFARX1 I_25044 (I428617,I2859,I428272,I428261,);
and I_25045 (I428255,I428363,I428552);
nor I_25046 (I428662,I428535,I355495);
and I_25047 (I428679,I428662,I355483);
or I_25048 (I428696,I428679,I355486);
DFFARX1 I_25049 (I428696,I2859,I428272,I428722,);
nor I_25050 (I428730,I428722,I428456);
DFFARX1 I_25051 (I428730,I2859,I428272,I428243,);
nand I_25052 (I428761,I428722,I428363);
nand I_25053 (I428778,I428456,I428761);
nor I_25054 (I428252,I428778,I428422);
not I_25055 (I428833,I2866);
DFFARX1 I_25056 (I144619,I2859,I428833,I428859,);
DFFARX1 I_25057 (I428859,I2859,I428833,I428876,);
not I_25058 (I428825,I428876);
not I_25059 (I428898,I428859);
DFFARX1 I_25060 (I144616,I2859,I428833,I428924,);
nand I_25061 (I428932,I428924,I144610);
not I_25062 (I428949,I144610);
not I_25063 (I428966,I144607);
nand I_25064 (I428983,I144601,I144598);
and I_25065 (I429000,I144601,I144598);
not I_25066 (I429017,I144613);
nand I_25067 (I429034,I429017,I428966);
nor I_25068 (I428807,I429034,I428932);
nor I_25069 (I429065,I428949,I429034);
nand I_25070 (I428810,I429000,I429065);
not I_25071 (I429096,I144625);
nor I_25072 (I429113,I429096,I144601);
nor I_25073 (I429130,I429113,I144613);
nor I_25074 (I429147,I428898,I429130);
DFFARX1 I_25075 (I429147,I2859,I428833,I428819,);
not I_25076 (I429178,I429113);
DFFARX1 I_25077 (I429178,I2859,I428833,I428822,);
and I_25078 (I428816,I428924,I429113);
nor I_25079 (I429223,I429096,I144622);
and I_25080 (I429240,I429223,I144598);
or I_25081 (I429257,I429240,I144604);
DFFARX1 I_25082 (I429257,I2859,I428833,I429283,);
nor I_25083 (I429291,I429283,I429017);
DFFARX1 I_25084 (I429291,I2859,I428833,I428804,);
nand I_25085 (I429322,I429283,I428924);
nand I_25086 (I429339,I429017,I429322);
nor I_25087 (I428813,I429339,I428983);
not I_25088 (I429394,I2866);
DFFARX1 I_25089 (I58445,I2859,I429394,I429420,);
DFFARX1 I_25090 (I429420,I2859,I429394,I429437,);
not I_25091 (I429386,I429437);
not I_25092 (I429459,I429420);
DFFARX1 I_25093 (I58460,I2859,I429394,I429485,);
nand I_25094 (I429493,I429485,I58442);
not I_25095 (I429510,I58442);
not I_25096 (I429527,I58451);
nand I_25097 (I429544,I58457,I58448);
and I_25098 (I429561,I58457,I58448);
not I_25099 (I429578,I58445);
nand I_25100 (I429595,I429578,I429527);
nor I_25101 (I429368,I429595,I429493);
nor I_25102 (I429626,I429510,I429595);
nand I_25103 (I429371,I429561,I429626);
not I_25104 (I429657,I58442);
nor I_25105 (I429674,I429657,I58457);
nor I_25106 (I429691,I429674,I58445);
nor I_25107 (I429708,I429459,I429691);
DFFARX1 I_25108 (I429708,I2859,I429394,I429380,);
not I_25109 (I429739,I429674);
DFFARX1 I_25110 (I429739,I2859,I429394,I429383,);
and I_25111 (I429377,I429485,I429674);
nor I_25112 (I429784,I429657,I58466);
and I_25113 (I429801,I429784,I58463);
or I_25114 (I429818,I429801,I58454);
DFFARX1 I_25115 (I429818,I2859,I429394,I429844,);
nor I_25116 (I429852,I429844,I429578);
DFFARX1 I_25117 (I429852,I2859,I429394,I429365,);
nand I_25118 (I429883,I429844,I429485);
nand I_25119 (I429900,I429578,I429883);
nor I_25120 (I429374,I429900,I429544);
not I_25121 (I429955,I2866);
DFFARX1 I_25122 (I489781,I2859,I429955,I429981,);
DFFARX1 I_25123 (I429981,I2859,I429955,I429998,);
not I_25124 (I429947,I429998);
not I_25125 (I430020,I429981);
DFFARX1 I_25126 (I489772,I2859,I429955,I430046,);
nand I_25127 (I430054,I430046,I489769);
not I_25128 (I430071,I489769);
not I_25129 (I430088,I489778);
nand I_25130 (I430105,I489787,I489769);
and I_25131 (I430122,I489787,I489769);
not I_25132 (I430139,I489766);
nand I_25133 (I430156,I430139,I430088);
nor I_25134 (I429929,I430156,I430054);
nor I_25135 (I430187,I430071,I430156);
nand I_25136 (I429932,I430122,I430187);
not I_25137 (I430218,I489775);
nor I_25138 (I430235,I430218,I489787);
nor I_25139 (I430252,I430235,I489766);
nor I_25140 (I430269,I430020,I430252);
DFFARX1 I_25141 (I430269,I2859,I429955,I429941,);
not I_25142 (I430300,I430235);
DFFARX1 I_25143 (I430300,I2859,I429955,I429944,);
and I_25144 (I429938,I430046,I430235);
nor I_25145 (I430345,I430218,I489790);
and I_25146 (I430362,I430345,I489766);
or I_25147 (I430379,I430362,I489784);
DFFARX1 I_25148 (I430379,I2859,I429955,I430405,);
nor I_25149 (I430413,I430405,I430139);
DFFARX1 I_25150 (I430413,I2859,I429955,I429926,);
nand I_25151 (I430444,I430405,I430046);
nand I_25152 (I430461,I430139,I430444);
nor I_25153 (I429935,I430461,I430105);
not I_25154 (I430516,I2866);
DFFARX1 I_25155 (I520063,I2859,I430516,I430542,);
DFFARX1 I_25156 (I430542,I2859,I430516,I430559,);
not I_25157 (I430508,I430559);
not I_25158 (I430581,I430542);
DFFARX1 I_25159 (I520060,I2859,I430516,I430607,);
nand I_25160 (I430615,I430607,I520066);
not I_25161 (I430632,I520066);
not I_25162 (I430649,I520075);
nand I_25163 (I430666,I520069,I520063);
and I_25164 (I430683,I520069,I520063);
not I_25165 (I430700,I520081);
nand I_25166 (I430717,I430700,I430649);
nor I_25167 (I430490,I430717,I430615);
nor I_25168 (I430748,I430632,I430717);
nand I_25169 (I430493,I430683,I430748);
not I_25170 (I430779,I520078);
nor I_25171 (I430796,I430779,I520069);
nor I_25172 (I430813,I430796,I520081);
nor I_25173 (I430830,I430581,I430813);
DFFARX1 I_25174 (I430830,I2859,I430516,I430502,);
not I_25175 (I430861,I430796);
DFFARX1 I_25176 (I430861,I2859,I430516,I430505,);
and I_25177 (I430499,I430607,I430796);
nor I_25178 (I430906,I430779,I520072);
and I_25179 (I430923,I430906,I520084);
or I_25180 (I430940,I430923,I520060);
DFFARX1 I_25181 (I430940,I2859,I430516,I430966,);
nor I_25182 (I430974,I430966,I430700);
DFFARX1 I_25183 (I430974,I2859,I430516,I430487,);
nand I_25184 (I431005,I430966,I430607);
nand I_25185 (I431022,I430700,I431005);
nor I_25186 (I430496,I431022,I430666);
not I_25187 (I431077,I2866);
DFFARX1 I_25188 (I372143,I2859,I431077,I431103,);
DFFARX1 I_25189 (I431103,I2859,I431077,I431120,);
not I_25190 (I431069,I431120);
not I_25191 (I431142,I431103);
DFFARX1 I_25192 (I372170,I2859,I431077,I431168,);
nand I_25193 (I431176,I431168,I372161);
not I_25194 (I431193,I372161);
not I_25195 (I431210,I372143);
nand I_25196 (I431227,I372155,I372158);
and I_25197 (I431244,I372155,I372158);
not I_25198 (I431261,I372167);
nand I_25199 (I431278,I431261,I431210);
nor I_25200 (I431051,I431278,I431176);
nor I_25201 (I431309,I431193,I431278);
nand I_25202 (I431054,I431244,I431309);
not I_25203 (I431340,I372152);
nor I_25204 (I431357,I431340,I372155);
nor I_25205 (I431374,I431357,I372167);
nor I_25206 (I431391,I431142,I431374);
DFFARX1 I_25207 (I431391,I2859,I431077,I431063,);
not I_25208 (I431422,I431357);
DFFARX1 I_25209 (I431422,I2859,I431077,I431066,);
and I_25210 (I431060,I431168,I431357);
nor I_25211 (I431467,I431340,I372146);
and I_25212 (I431484,I431467,I372149);
or I_25213 (I431501,I431484,I372164);
DFFARX1 I_25214 (I431501,I2859,I431077,I431527,);
nor I_25215 (I431535,I431527,I431261);
DFFARX1 I_25216 (I431535,I2859,I431077,I431048,);
nand I_25217 (I431566,I431527,I431168);
nand I_25218 (I431583,I431261,I431566);
nor I_25219 (I431057,I431583,I431227);
not I_25220 (I431638,I2866);
DFFARX1 I_25221 (I526421,I2859,I431638,I431664,);
DFFARX1 I_25222 (I431664,I2859,I431638,I431681,);
not I_25223 (I431630,I431681);
not I_25224 (I431703,I431664);
DFFARX1 I_25225 (I526418,I2859,I431638,I431729,);
nand I_25226 (I431737,I431729,I526424);
not I_25227 (I431754,I526424);
not I_25228 (I431771,I526433);
nand I_25229 (I431788,I526427,I526421);
and I_25230 (I431805,I526427,I526421);
not I_25231 (I431822,I526439);
nand I_25232 (I431839,I431822,I431771);
nor I_25233 (I431612,I431839,I431737);
nor I_25234 (I431870,I431754,I431839);
nand I_25235 (I431615,I431805,I431870);
not I_25236 (I431901,I526436);
nor I_25237 (I431918,I431901,I526427);
nor I_25238 (I431935,I431918,I526439);
nor I_25239 (I431952,I431703,I431935);
DFFARX1 I_25240 (I431952,I2859,I431638,I431624,);
not I_25241 (I431983,I431918);
DFFARX1 I_25242 (I431983,I2859,I431638,I431627,);
and I_25243 (I431621,I431729,I431918);
nor I_25244 (I432028,I431901,I526430);
and I_25245 (I432045,I432028,I526442);
or I_25246 (I432062,I432045,I526418);
DFFARX1 I_25247 (I432062,I2859,I431638,I432088,);
nor I_25248 (I432096,I432088,I431822);
DFFARX1 I_25249 (I432096,I2859,I431638,I431609,);
nand I_25250 (I432127,I432088,I431729);
nand I_25251 (I432144,I431822,I432127);
nor I_25252 (I431618,I432144,I431788);
not I_25253 (I432199,I2866);
DFFARX1 I_25254 (I163152,I2859,I432199,I432225,);
DFFARX1 I_25255 (I432225,I2859,I432199,I432242,);
not I_25256 (I432191,I432242);
not I_25257 (I432264,I432225);
DFFARX1 I_25258 (I163140,I2859,I432199,I432290,);
nand I_25259 (I432298,I432290,I163146);
not I_25260 (I432315,I163146);
not I_25261 (I432332,I163143);
nand I_25262 (I432349,I163131,I163128);
and I_25263 (I432366,I163131,I163128);
not I_25264 (I432383,I163155);
nand I_25265 (I432400,I432383,I432332);
nor I_25266 (I432173,I432400,I432298);
nor I_25267 (I432431,I432315,I432400);
nand I_25268 (I432176,I432366,I432431);
not I_25269 (I432462,I163128);
nor I_25270 (I432479,I432462,I163131);
nor I_25271 (I432496,I432479,I163155);
nor I_25272 (I432513,I432264,I432496);
DFFARX1 I_25273 (I432513,I2859,I432199,I432185,);
not I_25274 (I432544,I432479);
DFFARX1 I_25275 (I432544,I2859,I432199,I432188,);
and I_25276 (I432182,I432290,I432479);
nor I_25277 (I432589,I432462,I163137);
and I_25278 (I432606,I432589,I163134);
or I_25279 (I432623,I432606,I163149);
DFFARX1 I_25280 (I432623,I2859,I432199,I432649,);
nor I_25281 (I432657,I432649,I432383);
DFFARX1 I_25282 (I432657,I2859,I432199,I432170,);
nand I_25283 (I432688,I432649,I432290);
nand I_25284 (I432705,I432383,I432688);
nor I_25285 (I432179,I432705,I432349);
not I_25286 (I432760,I2866);
DFFARX1 I_25287 (I83435,I2859,I432760,I432786,);
DFFARX1 I_25288 (I432786,I2859,I432760,I432803,);
not I_25289 (I432752,I432803);
not I_25290 (I432825,I432786);
DFFARX1 I_25291 (I83450,I2859,I432760,I432851,);
nand I_25292 (I432859,I432851,I83432);
not I_25293 (I432876,I83432);
not I_25294 (I432893,I83441);
nand I_25295 (I432910,I83447,I83438);
and I_25296 (I432927,I83447,I83438);
not I_25297 (I432944,I83435);
nand I_25298 (I432961,I432944,I432893);
nor I_25299 (I432734,I432961,I432859);
nor I_25300 (I432992,I432876,I432961);
nand I_25301 (I432737,I432927,I432992);
not I_25302 (I433023,I83432);
nor I_25303 (I433040,I433023,I83447);
nor I_25304 (I433057,I433040,I83435);
nor I_25305 (I433074,I432825,I433057);
DFFARX1 I_25306 (I433074,I2859,I432760,I432746,);
not I_25307 (I433105,I433040);
DFFARX1 I_25308 (I433105,I2859,I432760,I432749,);
and I_25309 (I432743,I432851,I433040);
nor I_25310 (I433150,I433023,I83456);
and I_25311 (I433167,I433150,I83453);
or I_25312 (I433184,I433167,I83444);
DFFARX1 I_25313 (I433184,I2859,I432760,I433210,);
nor I_25314 (I433218,I433210,I432944);
DFFARX1 I_25315 (I433218,I2859,I432760,I432731,);
nand I_25316 (I433249,I433210,I432851);
nand I_25317 (I433266,I432944,I433249);
nor I_25318 (I432740,I433266,I432910);
not I_25319 (I433321,I2866);
DFFARX1 I_25320 (I359708,I2859,I433321,I433347,);
DFFARX1 I_25321 (I433347,I2859,I433321,I433364,);
not I_25322 (I433313,I433364);
not I_25323 (I433386,I433347);
DFFARX1 I_25324 (I359705,I2859,I433321,I433412,);
nand I_25325 (I433420,I433412,I359720);
not I_25326 (I433437,I359720);
not I_25327 (I433454,I359717);
nand I_25328 (I433471,I359714,I359702);
and I_25329 (I433488,I359714,I359702);
not I_25330 (I433505,I359699);
nand I_25331 (I433522,I433505,I433454);
nor I_25332 (I433295,I433522,I433420);
nor I_25333 (I433553,I433437,I433522);
nand I_25334 (I433298,I433488,I433553);
not I_25335 (I433584,I359705);
nor I_25336 (I433601,I433584,I359714);
nor I_25337 (I433618,I433601,I359699);
nor I_25338 (I433635,I433386,I433618);
DFFARX1 I_25339 (I433635,I2859,I433321,I433307,);
not I_25340 (I433666,I433601);
DFFARX1 I_25341 (I433666,I2859,I433321,I433310,);
and I_25342 (I433304,I433412,I433601);
nor I_25343 (I433711,I433584,I359711);
and I_25344 (I433728,I433711,I359699);
or I_25345 (I433745,I433728,I359702);
DFFARX1 I_25346 (I433745,I2859,I433321,I433771,);
nor I_25347 (I433779,I433771,I433505);
DFFARX1 I_25348 (I433779,I2859,I433321,I433292,);
nand I_25349 (I433810,I433771,I433412);
nand I_25350 (I433827,I433505,I433810);
nor I_25351 (I433301,I433827,I433471);
not I_25352 (I433882,I2866);
DFFARX1 I_25353 (I286279,I2859,I433882,I433908,);
DFFARX1 I_25354 (I433908,I2859,I433882,I433925,);
not I_25355 (I433874,I433925);
not I_25356 (I433947,I433908);
DFFARX1 I_25357 (I286291,I2859,I433882,I433973,);
nand I_25358 (I433981,I433973,I286300);
not I_25359 (I433998,I286300);
not I_25360 (I434015,I286282);
nand I_25361 (I434032,I286285,I286276);
and I_25362 (I434049,I286285,I286276);
not I_25363 (I434066,I286294);
nand I_25364 (I434083,I434066,I434015);
nor I_25365 (I433856,I434083,I433981);
nor I_25366 (I434114,I433998,I434083);
nand I_25367 (I433859,I434049,I434114);
not I_25368 (I434145,I286297);
nor I_25369 (I434162,I434145,I286285);
nor I_25370 (I434179,I434162,I286294);
nor I_25371 (I434196,I433947,I434179);
DFFARX1 I_25372 (I434196,I2859,I433882,I433868,);
not I_25373 (I434227,I434162);
DFFARX1 I_25374 (I434227,I2859,I433882,I433871,);
and I_25375 (I433865,I433973,I434162);
nor I_25376 (I434272,I434145,I286276);
and I_25377 (I434289,I434272,I286288);
or I_25378 (I434306,I434289,I286279);
DFFARX1 I_25379 (I434306,I2859,I433882,I434332,);
nor I_25380 (I434340,I434332,I434066);
DFFARX1 I_25381 (I434340,I2859,I433882,I433853,);
nand I_25382 (I434371,I434332,I433973);
nand I_25383 (I434388,I434066,I434371);
nor I_25384 (I433862,I434388,I434032);
not I_25385 (I434443,I2866);
DFFARX1 I_25386 (I150943,I2859,I434443,I434469,);
DFFARX1 I_25387 (I434469,I2859,I434443,I434486,);
not I_25388 (I434435,I434486);
not I_25389 (I434508,I434469);
DFFARX1 I_25390 (I150940,I2859,I434443,I434534,);
nand I_25391 (I434542,I434534,I150934);
not I_25392 (I434559,I150934);
not I_25393 (I434576,I150931);
nand I_25394 (I434593,I150925,I150922);
and I_25395 (I434610,I150925,I150922);
not I_25396 (I434627,I150937);
nand I_25397 (I434644,I434627,I434576);
nor I_25398 (I434417,I434644,I434542);
nor I_25399 (I434675,I434559,I434644);
nand I_25400 (I434420,I434610,I434675);
not I_25401 (I434706,I150949);
nor I_25402 (I434723,I434706,I150925);
nor I_25403 (I434740,I434723,I150937);
nor I_25404 (I434757,I434508,I434740);
DFFARX1 I_25405 (I434757,I2859,I434443,I434429,);
not I_25406 (I434788,I434723);
DFFARX1 I_25407 (I434788,I2859,I434443,I434432,);
and I_25408 (I434426,I434534,I434723);
nor I_25409 (I434833,I434706,I150946);
and I_25410 (I434850,I434833,I150922);
or I_25411 (I434867,I434850,I150928);
DFFARX1 I_25412 (I434867,I2859,I434443,I434893,);
nor I_25413 (I434901,I434893,I434627);
DFFARX1 I_25414 (I434901,I2859,I434443,I434414,);
nand I_25415 (I434932,I434893,I434534);
nand I_25416 (I434949,I434627,I434932);
nor I_25417 (I434423,I434949,I434593);
not I_25418 (I435004,I2866);
DFFARX1 I_25419 (I250440,I2859,I435004,I435030,);
DFFARX1 I_25420 (I435030,I2859,I435004,I435047,);
not I_25421 (I434996,I435047);
not I_25422 (I435069,I435030);
DFFARX1 I_25423 (I250455,I2859,I435004,I435095,);
nand I_25424 (I435103,I435095,I250446);
not I_25425 (I435120,I250446);
not I_25426 (I435137,I250452);
nand I_25427 (I435154,I250449,I250458);
and I_25428 (I435171,I250449,I250458);
not I_25429 (I435188,I250443);
nand I_25430 (I435205,I435188,I435137);
nor I_25431 (I434978,I435205,I435103);
nor I_25432 (I435236,I435120,I435205);
nand I_25433 (I434981,I435171,I435236);
not I_25434 (I435267,I250440);
nor I_25435 (I435284,I435267,I250449);
nor I_25436 (I435301,I435284,I250443);
nor I_25437 (I435318,I435069,I435301);
DFFARX1 I_25438 (I435318,I2859,I435004,I434990,);
not I_25439 (I435349,I435284);
DFFARX1 I_25440 (I435349,I2859,I435004,I434993,);
and I_25441 (I434987,I435095,I435284);
nor I_25442 (I435394,I435267,I250464);
and I_25443 (I435411,I435394,I250443);
or I_25444 (I435428,I435411,I250461);
DFFARX1 I_25445 (I435428,I2859,I435004,I435454,);
nor I_25446 (I435462,I435454,I435188);
DFFARX1 I_25447 (I435462,I2859,I435004,I434975,);
nand I_25448 (I435493,I435454,I435095);
nand I_25449 (I435510,I435188,I435493);
nor I_25450 (I434984,I435510,I435154);
not I_25451 (I435565,I2866);
DFFARX1 I_25452 (I370205,I2859,I435565,I435591,);
DFFARX1 I_25453 (I435591,I2859,I435565,I435608,);
not I_25454 (I435557,I435608);
not I_25455 (I435630,I435591);
DFFARX1 I_25456 (I370232,I2859,I435565,I435656,);
nand I_25457 (I435664,I435656,I370223);
not I_25458 (I435681,I370223);
not I_25459 (I435698,I370205);
nand I_25460 (I435715,I370217,I370220);
and I_25461 (I435732,I370217,I370220);
not I_25462 (I435749,I370229);
nand I_25463 (I435766,I435749,I435698);
nor I_25464 (I435539,I435766,I435664);
nor I_25465 (I435797,I435681,I435766);
nand I_25466 (I435542,I435732,I435797);
not I_25467 (I435828,I370214);
nor I_25468 (I435845,I435828,I370217);
nor I_25469 (I435862,I435845,I370229);
nor I_25470 (I435879,I435630,I435862);
DFFARX1 I_25471 (I435879,I2859,I435565,I435551,);
not I_25472 (I435910,I435845);
DFFARX1 I_25473 (I435910,I2859,I435565,I435554,);
and I_25474 (I435548,I435656,I435845);
nor I_25475 (I435955,I435828,I370208);
and I_25476 (I435972,I435955,I370211);
or I_25477 (I435989,I435972,I370226);
DFFARX1 I_25478 (I435989,I2859,I435565,I436015,);
nor I_25479 (I436023,I436015,I435749);
DFFARX1 I_25480 (I436023,I2859,I435565,I435536,);
nand I_25481 (I436054,I436015,I435656);
nand I_25482 (I436071,I435749,I436054);
nor I_25483 (I435545,I436071,I435715);
not I_25484 (I436126,I2866);
DFFARX1 I_25485 (I451633,I2859,I436126,I436152,);
DFFARX1 I_25486 (I436152,I2859,I436126,I436169,);
not I_25487 (I436118,I436169);
not I_25488 (I436191,I436152);
DFFARX1 I_25489 (I451624,I2859,I436126,I436217,);
nand I_25490 (I436225,I436217,I451621);
not I_25491 (I436242,I451621);
not I_25492 (I436259,I451630);
nand I_25493 (I436276,I451639,I451621);
and I_25494 (I436293,I451639,I451621);
not I_25495 (I436310,I451618);
nand I_25496 (I436327,I436310,I436259);
nor I_25497 (I436100,I436327,I436225);
nor I_25498 (I436358,I436242,I436327);
nand I_25499 (I436103,I436293,I436358);
not I_25500 (I436389,I451627);
nor I_25501 (I436406,I436389,I451639);
nor I_25502 (I436423,I436406,I451618);
nor I_25503 (I436440,I436191,I436423);
DFFARX1 I_25504 (I436440,I2859,I436126,I436112,);
not I_25505 (I436471,I436406);
DFFARX1 I_25506 (I436471,I2859,I436126,I436115,);
and I_25507 (I436109,I436217,I436406);
nor I_25508 (I436516,I436389,I451642);
and I_25509 (I436533,I436516,I451618);
or I_25510 (I436550,I436533,I451636);
DFFARX1 I_25511 (I436550,I2859,I436126,I436576,);
nor I_25512 (I436584,I436576,I436310);
DFFARX1 I_25513 (I436584,I2859,I436126,I436097,);
nand I_25514 (I436615,I436576,I436217);
nand I_25515 (I436632,I436310,I436615);
nor I_25516 (I436106,I436632,I436276);
not I_25517 (I436687,I2866);
DFFARX1 I_25518 (I570140,I2859,I436687,I436713,);
DFFARX1 I_25519 (I436713,I2859,I436687,I436730,);
not I_25520 (I436679,I436730);
not I_25521 (I436752,I436713);
DFFARX1 I_25522 (I570134,I2859,I436687,I436778,);
nand I_25523 (I436786,I436778,I570125);
not I_25524 (I436803,I570125);
not I_25525 (I436820,I570152);
nand I_25526 (I436837,I570137,I570146);
and I_25527 (I436854,I570137,I570146);
not I_25528 (I436871,I570131);
nand I_25529 (I436888,I436871,I436820);
nor I_25530 (I436661,I436888,I436786);
nor I_25531 (I436919,I436803,I436888);
nand I_25532 (I436664,I436854,I436919);
not I_25533 (I436950,I570149);
nor I_25534 (I436967,I436950,I570137);
nor I_25535 (I436984,I436967,I570131);
nor I_25536 (I437001,I436752,I436984);
DFFARX1 I_25537 (I437001,I2859,I436687,I436673,);
not I_25538 (I437032,I436967);
DFFARX1 I_25539 (I437032,I2859,I436687,I436676,);
and I_25540 (I436670,I436778,I436967);
nor I_25541 (I437077,I436950,I570143);
and I_25542 (I437094,I437077,I570125);
or I_25543 (I437111,I437094,I570128);
DFFARX1 I_25544 (I437111,I2859,I436687,I437137,);
nor I_25545 (I437145,I437137,I436871);
DFFARX1 I_25546 (I437145,I2859,I436687,I436658,);
nand I_25547 (I437176,I437137,I436778);
nand I_25548 (I437193,I436871,I437176);
nor I_25549 (I436667,I437193,I436837);
not I_25550 (I437248,I2866);
DFFARX1 I_25551 (I193616,I2859,I437248,I437274,);
DFFARX1 I_25552 (I437274,I2859,I437248,I437291,);
not I_25553 (I437240,I437291);
not I_25554 (I437313,I437274);
DFFARX1 I_25555 (I193604,I2859,I437248,I437339,);
nand I_25556 (I437347,I437339,I193610);
not I_25557 (I437364,I193610);
not I_25558 (I437381,I193607);
nand I_25559 (I437398,I193595,I193592);
and I_25560 (I437415,I193595,I193592);
not I_25561 (I437432,I193619);
nand I_25562 (I437449,I437432,I437381);
nor I_25563 (I437222,I437449,I437347);
nor I_25564 (I437480,I437364,I437449);
nand I_25565 (I437225,I437415,I437480);
not I_25566 (I437511,I193592);
nor I_25567 (I437528,I437511,I193595);
nor I_25568 (I437545,I437528,I193619);
nor I_25569 (I437562,I437313,I437545);
DFFARX1 I_25570 (I437562,I2859,I437248,I437234,);
not I_25571 (I437593,I437528);
DFFARX1 I_25572 (I437593,I2859,I437248,I437237,);
and I_25573 (I437231,I437339,I437528);
nor I_25574 (I437638,I437511,I193601);
and I_25575 (I437655,I437638,I193598);
or I_25576 (I437672,I437655,I193613);
DFFARX1 I_25577 (I437672,I2859,I437248,I437698,);
nor I_25578 (I437706,I437698,I437432);
DFFARX1 I_25579 (I437706,I2859,I437248,I437219,);
nand I_25580 (I437737,I437698,I437339);
nand I_25581 (I437754,I437432,I437737);
nor I_25582 (I437228,I437754,I437398);
not I_25583 (I437809,I2866);
DFFARX1 I_25584 (I149889,I2859,I437809,I437835,);
DFFARX1 I_25585 (I437835,I2859,I437809,I437852,);
not I_25586 (I437801,I437852);
not I_25587 (I437874,I437835);
DFFARX1 I_25588 (I149886,I2859,I437809,I437900,);
nand I_25589 (I437908,I437900,I149880);
not I_25590 (I437925,I149880);
not I_25591 (I437942,I149877);
nand I_25592 (I437959,I149871,I149868);
and I_25593 (I437976,I149871,I149868);
not I_25594 (I437993,I149883);
nand I_25595 (I438010,I437993,I437942);
nor I_25596 (I437783,I438010,I437908);
nor I_25597 (I438041,I437925,I438010);
nand I_25598 (I437786,I437976,I438041);
not I_25599 (I438072,I149895);
nor I_25600 (I438089,I438072,I149871);
nor I_25601 (I438106,I438089,I149883);
nor I_25602 (I438123,I437874,I438106);
DFFARX1 I_25603 (I438123,I2859,I437809,I437795,);
not I_25604 (I438154,I438089);
DFFARX1 I_25605 (I438154,I2859,I437809,I437798,);
and I_25606 (I437792,I437900,I438089);
nor I_25607 (I438199,I438072,I149892);
and I_25608 (I438216,I438199,I149868);
or I_25609 (I438233,I438216,I149874);
DFFARX1 I_25610 (I438233,I2859,I437809,I438259,);
nor I_25611 (I438267,I438259,I437993);
DFFARX1 I_25612 (I438267,I2859,I437809,I437780,);
nand I_25613 (I438298,I438259,I437900);
nand I_25614 (I438315,I437993,I438298);
nor I_25615 (I437789,I438315,I437959);
not I_25616 (I438370,I2866);
DFFARX1 I_25617 (I201328,I2859,I438370,I438396,);
DFFARX1 I_25618 (I438396,I2859,I438370,I438413,);
not I_25619 (I438362,I438413);
not I_25620 (I438435,I438396);
DFFARX1 I_25621 (I201325,I2859,I438370,I438461,);
nand I_25622 (I438469,I438461,I201319);
not I_25623 (I438486,I201319);
not I_25624 (I438503,I201331);
nand I_25625 (I438520,I201334,I201313);
and I_25626 (I438537,I201334,I201313);
not I_25627 (I438554,I201310);
nand I_25628 (I438571,I438554,I438503);
nor I_25629 (I438344,I438571,I438469);
nor I_25630 (I438602,I438486,I438571);
nand I_25631 (I438347,I438537,I438602);
not I_25632 (I438633,I201316);
nor I_25633 (I438650,I438633,I201334);
nor I_25634 (I438667,I438650,I201310);
nor I_25635 (I438684,I438435,I438667);
DFFARX1 I_25636 (I438684,I2859,I438370,I438356,);
not I_25637 (I438715,I438650);
DFFARX1 I_25638 (I438715,I2859,I438370,I438359,);
and I_25639 (I438353,I438461,I438650);
nor I_25640 (I438760,I438633,I201310);
and I_25641 (I438777,I438760,I201322);
or I_25642 (I438794,I438777,I201313);
DFFARX1 I_25643 (I438794,I2859,I438370,I438820,);
nor I_25644 (I438828,I438820,I438554);
DFFARX1 I_25645 (I438828,I2859,I438370,I438341,);
nand I_25646 (I438859,I438820,I438461);
nand I_25647 (I438876,I438554,I438859);
nor I_25648 (I438350,I438876,I438520);
not I_25649 (I438934,I2866);
DFFARX1 I_25650 (I370857,I2859,I438934,I438960,);
and I_25651 (I438968,I438960,I370851);
DFFARX1 I_25652 (I438968,I2859,I438934,I438917,);
DFFARX1 I_25653 (I370869,I2859,I438934,I439008,);
not I_25654 (I439016,I370860);
not I_25655 (I439033,I370872);
nand I_25656 (I439050,I439033,I439016);
nor I_25657 (I438905,I439008,I439050);
DFFARX1 I_25658 (I439050,I2859,I438934,I439090,);
not I_25659 (I438926,I439090);
not I_25660 (I439112,I370878);
nand I_25661 (I439129,I439033,I439112);
DFFARX1 I_25662 (I439129,I2859,I438934,I439155,);
not I_25663 (I439163,I439155);
not I_25664 (I439180,I370854);
nand I_25665 (I439197,I439180,I370875);
and I_25666 (I439214,I439016,I439197);
nor I_25667 (I439231,I439129,I439214);
DFFARX1 I_25668 (I439231,I2859,I438934,I438902,);
DFFARX1 I_25669 (I439214,I2859,I438934,I438923,);
nor I_25670 (I439276,I370854,I370866);
nor I_25671 (I438914,I439129,I439276);
or I_25672 (I439307,I370854,I370866);
nor I_25673 (I439324,I370851,I370863);
DFFARX1 I_25674 (I439324,I2859,I438934,I439350,);
not I_25675 (I439358,I439350);
nor I_25676 (I438920,I439358,I439163);
nand I_25677 (I439389,I439358,I439008);
not I_25678 (I439406,I370851);
nand I_25679 (I439423,I439406,I439112);
nand I_25680 (I439440,I439358,I439423);
nand I_25681 (I438911,I439440,I439389);
nand I_25682 (I438908,I439423,I439307);
not I_25683 (I439512,I2866);
DFFARX1 I_25684 (I23786,I2859,I439512,I439538,);
and I_25685 (I439546,I439538,I23762);
DFFARX1 I_25686 (I439546,I2859,I439512,I439495,);
DFFARX1 I_25687 (I23780,I2859,I439512,I439586,);
not I_25688 (I439594,I23768);
not I_25689 (I439611,I23765);
nand I_25690 (I439628,I439611,I439594);
nor I_25691 (I439483,I439586,I439628);
DFFARX1 I_25692 (I439628,I2859,I439512,I439668,);
not I_25693 (I439504,I439668);
not I_25694 (I439690,I23774);
nand I_25695 (I439707,I439611,I439690);
DFFARX1 I_25696 (I439707,I2859,I439512,I439733,);
not I_25697 (I439741,I439733);
not I_25698 (I439758,I23765);
nand I_25699 (I439775,I439758,I23783);
and I_25700 (I439792,I439594,I439775);
nor I_25701 (I439809,I439707,I439792);
DFFARX1 I_25702 (I439809,I2859,I439512,I439480,);
DFFARX1 I_25703 (I439792,I2859,I439512,I439501,);
nor I_25704 (I439854,I23765,I23777);
nor I_25705 (I439492,I439707,I439854);
or I_25706 (I439885,I23765,I23777);
nor I_25707 (I439902,I23771,I23762);
DFFARX1 I_25708 (I439902,I2859,I439512,I439928,);
not I_25709 (I439936,I439928);
nor I_25710 (I439498,I439936,I439741);
nand I_25711 (I439967,I439936,I439586);
not I_25712 (I439984,I23771);
nand I_25713 (I440001,I439984,I439690);
nand I_25714 (I440018,I439936,I440001);
nand I_25715 (I439489,I440018,I439967);
nand I_25716 (I439486,I440001,I439885);
not I_25717 (I440090,I2866);
DFFARX1 I_25718 (I246409,I2859,I440090,I440116,);
and I_25719 (I440124,I440116,I246397);
DFFARX1 I_25720 (I440124,I2859,I440090,I440073,);
DFFARX1 I_25721 (I246412,I2859,I440090,I440164,);
not I_25722 (I440172,I246403);
not I_25723 (I440189,I246394);
nand I_25724 (I440206,I440189,I440172);
nor I_25725 (I440061,I440164,I440206);
DFFARX1 I_25726 (I440206,I2859,I440090,I440246,);
not I_25727 (I440082,I440246);
not I_25728 (I440268,I246400);
nand I_25729 (I440285,I440189,I440268);
DFFARX1 I_25730 (I440285,I2859,I440090,I440311,);
not I_25731 (I440319,I440311);
not I_25732 (I440336,I246415);
nand I_25733 (I440353,I440336,I246418);
and I_25734 (I440370,I440172,I440353);
nor I_25735 (I440387,I440285,I440370);
DFFARX1 I_25736 (I440387,I2859,I440090,I440058,);
DFFARX1 I_25737 (I440370,I2859,I440090,I440079,);
nor I_25738 (I440432,I246415,I246394);
nor I_25739 (I440070,I440285,I440432);
or I_25740 (I440463,I246415,I246394);
nor I_25741 (I440480,I246406,I246397);
DFFARX1 I_25742 (I440480,I2859,I440090,I440506,);
not I_25743 (I440514,I440506);
nor I_25744 (I440076,I440514,I440319);
nand I_25745 (I440545,I440514,I440164);
not I_25746 (I440562,I246406);
nand I_25747 (I440579,I440562,I440268);
nand I_25748 (I440596,I440514,I440579);
nand I_25749 (I440067,I440596,I440545);
nand I_25750 (I440064,I440579,I440463);
not I_25751 (I440668,I2866);
DFFARX1 I_25752 (I209643,I2859,I440668,I440694,);
and I_25753 (I440702,I440694,I209658);
DFFARX1 I_25754 (I440702,I2859,I440668,I440651,);
DFFARX1 I_25755 (I209649,I2859,I440668,I440742,);
not I_25756 (I440750,I209643);
not I_25757 (I440767,I209661);
nand I_25758 (I440784,I440767,I440750);
nor I_25759 (I440639,I440742,I440784);
DFFARX1 I_25760 (I440784,I2859,I440668,I440824,);
not I_25761 (I440660,I440824);
not I_25762 (I440846,I209652);
nand I_25763 (I440863,I440767,I440846);
DFFARX1 I_25764 (I440863,I2859,I440668,I440889,);
not I_25765 (I440897,I440889);
not I_25766 (I440914,I209664);
nand I_25767 (I440931,I440914,I209640);
and I_25768 (I440948,I440750,I440931);
nor I_25769 (I440965,I440863,I440948);
DFFARX1 I_25770 (I440965,I2859,I440668,I440636,);
DFFARX1 I_25771 (I440948,I2859,I440668,I440657,);
nor I_25772 (I441010,I209664,I209640);
nor I_25773 (I440648,I440863,I441010);
or I_25774 (I441041,I209664,I209640);
nor I_25775 (I441058,I209646,I209655);
DFFARX1 I_25776 (I441058,I2859,I440668,I441084,);
not I_25777 (I441092,I441084);
nor I_25778 (I440654,I441092,I440897);
nand I_25779 (I441123,I441092,I440742);
not I_25780 (I441140,I209646);
nand I_25781 (I441157,I441140,I440846);
nand I_25782 (I441174,I441092,I441157);
nand I_25783 (I440645,I441174,I441123);
nand I_25784 (I440642,I441157,I441041);
not I_25785 (I441246,I2866);
DFFARX1 I_25786 (I318596,I2859,I441246,I441272,);
and I_25787 (I441280,I441272,I318602);
DFFARX1 I_25788 (I441280,I2859,I441246,I441229,);
DFFARX1 I_25789 (I318608,I2859,I441246,I441320,);
not I_25790 (I441328,I318593);
not I_25791 (I441345,I318593);
nand I_25792 (I441362,I441345,I441328);
nor I_25793 (I441217,I441320,I441362);
DFFARX1 I_25794 (I441362,I2859,I441246,I441402,);
not I_25795 (I441238,I441402);
not I_25796 (I441424,I318611);
nand I_25797 (I441441,I441345,I441424);
DFFARX1 I_25798 (I441441,I2859,I441246,I441467,);
not I_25799 (I441475,I441467);
not I_25800 (I441492,I318605);
nand I_25801 (I441509,I441492,I318596);
and I_25802 (I441526,I441328,I441509);
nor I_25803 (I441543,I441441,I441526);
DFFARX1 I_25804 (I441543,I2859,I441246,I441214,);
DFFARX1 I_25805 (I441526,I2859,I441246,I441235,);
nor I_25806 (I441588,I318605,I318614);
nor I_25807 (I441226,I441441,I441588);
or I_25808 (I441619,I318605,I318614);
nor I_25809 (I441636,I318599,I318599);
DFFARX1 I_25810 (I441636,I2859,I441246,I441662,);
not I_25811 (I441670,I441662);
nor I_25812 (I441232,I441670,I441475);
nand I_25813 (I441701,I441670,I441320);
not I_25814 (I441718,I318599);
nand I_25815 (I441735,I441718,I441424);
nand I_25816 (I441752,I441670,I441735);
nand I_25817 (I441223,I441752,I441701);
nand I_25818 (I441220,I441735,I441619);
not I_25819 (I441824,I2866);
DFFARX1 I_25820 (I141463,I2859,I441824,I441850,);
and I_25821 (I441858,I441850,I141448);
DFFARX1 I_25822 (I441858,I2859,I441824,I441807,);
DFFARX1 I_25823 (I141454,I2859,I441824,I441898,);
not I_25824 (I441906,I141436);
not I_25825 (I441923,I141457);
nand I_25826 (I441940,I441923,I441906);
nor I_25827 (I441795,I441898,I441940);
DFFARX1 I_25828 (I441940,I2859,I441824,I441980,);
not I_25829 (I441816,I441980);
not I_25830 (I442002,I141460);
nand I_25831 (I442019,I441923,I442002);
DFFARX1 I_25832 (I442019,I2859,I441824,I442045,);
not I_25833 (I442053,I442045);
not I_25834 (I442070,I141451);
nand I_25835 (I442087,I442070,I141439);
and I_25836 (I442104,I441906,I442087);
nor I_25837 (I442121,I442019,I442104);
DFFARX1 I_25838 (I442121,I2859,I441824,I441792,);
DFFARX1 I_25839 (I442104,I2859,I441824,I441813,);
nor I_25840 (I442166,I141451,I141445);
nor I_25841 (I441804,I442019,I442166);
or I_25842 (I442197,I141451,I141445);
nor I_25843 (I442214,I141442,I141436);
DFFARX1 I_25844 (I442214,I2859,I441824,I442240,);
not I_25845 (I442248,I442240);
nor I_25846 (I441810,I442248,I442053);
nand I_25847 (I442279,I442248,I441898);
not I_25848 (I442296,I141442);
nand I_25849 (I442313,I442296,I442002);
nand I_25850 (I442330,I442248,I442313);
nand I_25851 (I441801,I442330,I442279);
nand I_25852 (I441798,I442313,I442197);
not I_25853 (I442402,I2866);
DFFARX1 I_25854 (I552302,I2859,I442402,I442428,);
and I_25855 (I442436,I442428,I552284);
DFFARX1 I_25856 (I442436,I2859,I442402,I442385,);
DFFARX1 I_25857 (I552275,I2859,I442402,I442476,);
not I_25858 (I442484,I552290);
not I_25859 (I442501,I552278);
nand I_25860 (I442518,I442501,I442484);
nor I_25861 (I442373,I442476,I442518);
DFFARX1 I_25862 (I442518,I2859,I442402,I442558,);
not I_25863 (I442394,I442558);
not I_25864 (I442580,I552287);
nand I_25865 (I442597,I442501,I442580);
DFFARX1 I_25866 (I442597,I2859,I442402,I442623,);
not I_25867 (I442631,I442623);
not I_25868 (I442648,I552296);
nand I_25869 (I442665,I442648,I552275);
and I_25870 (I442682,I442484,I442665);
nor I_25871 (I442699,I442597,I442682);
DFFARX1 I_25872 (I442699,I2859,I442402,I442370,);
DFFARX1 I_25873 (I442682,I2859,I442402,I442391,);
nor I_25874 (I442744,I552296,I552299);
nor I_25875 (I442382,I442597,I442744);
or I_25876 (I442775,I552296,I552299);
nor I_25877 (I442792,I552293,I552281);
DFFARX1 I_25878 (I442792,I2859,I442402,I442818,);
not I_25879 (I442826,I442818);
nor I_25880 (I442388,I442826,I442631);
nand I_25881 (I442857,I442826,I442476);
not I_25882 (I442874,I552293);
nand I_25883 (I442891,I442874,I442580);
nand I_25884 (I442908,I442826,I442891);
nand I_25885 (I442379,I442908,I442857);
nand I_25886 (I442376,I442891,I442775);
not I_25887 (I442980,I2866);
DFFARX1 I_25888 (I345473,I2859,I442980,I443006,);
and I_25889 (I443014,I443006,I345479);
DFFARX1 I_25890 (I443014,I2859,I442980,I442963,);
DFFARX1 I_25891 (I345485,I2859,I442980,I443054,);
not I_25892 (I443062,I345470);
not I_25893 (I443079,I345470);
nand I_25894 (I443096,I443079,I443062);
nor I_25895 (I442951,I443054,I443096);
DFFARX1 I_25896 (I443096,I2859,I442980,I443136,);
not I_25897 (I442972,I443136);
not I_25898 (I443158,I345488);
nand I_25899 (I443175,I443079,I443158);
DFFARX1 I_25900 (I443175,I2859,I442980,I443201,);
not I_25901 (I443209,I443201);
not I_25902 (I443226,I345482);
nand I_25903 (I443243,I443226,I345473);
and I_25904 (I443260,I443062,I443243);
nor I_25905 (I443277,I443175,I443260);
DFFARX1 I_25906 (I443277,I2859,I442980,I442948,);
DFFARX1 I_25907 (I443260,I2859,I442980,I442969,);
nor I_25908 (I443322,I345482,I345491);
nor I_25909 (I442960,I443175,I443322);
or I_25910 (I443353,I345482,I345491);
nor I_25911 (I443370,I345476,I345476);
DFFARX1 I_25912 (I443370,I2859,I442980,I443396,);
not I_25913 (I443404,I443396);
nor I_25914 (I442966,I443404,I443209);
nand I_25915 (I443435,I443404,I443054);
not I_25916 (I443452,I345476);
nand I_25917 (I443469,I443452,I443158);
nand I_25918 (I443486,I443404,I443469);
nand I_25919 (I442957,I443486,I443435);
nand I_25920 (I442954,I443469,I443353);
not I_25921 (I443558,I2866);
DFFARX1 I_25922 (I181624,I2859,I443558,I443584,);
and I_25923 (I443592,I443584,I181639);
DFFARX1 I_25924 (I443592,I2859,I443558,I443541,);
DFFARX1 I_25925 (I181642,I2859,I443558,I443632,);
not I_25926 (I443640,I181636);
not I_25927 (I443657,I181651);
nand I_25928 (I443674,I443657,I443640);
nor I_25929 (I443529,I443632,I443674);
DFFARX1 I_25930 (I443674,I2859,I443558,I443714,);
not I_25931 (I443550,I443714);
not I_25932 (I443736,I181627);
nand I_25933 (I443753,I443657,I443736);
DFFARX1 I_25934 (I443753,I2859,I443558,I443779,);
not I_25935 (I443787,I443779);
not I_25936 (I443804,I181630);
nand I_25937 (I443821,I443804,I181624);
and I_25938 (I443838,I443640,I443821);
nor I_25939 (I443855,I443753,I443838);
DFFARX1 I_25940 (I443855,I2859,I443558,I443526,);
DFFARX1 I_25941 (I443838,I2859,I443558,I443547,);
nor I_25942 (I443900,I181630,I181633);
nor I_25943 (I443538,I443753,I443900);
or I_25944 (I443931,I181630,I181633);
nor I_25945 (I443948,I181648,I181645);
DFFARX1 I_25946 (I443948,I2859,I443558,I443974,);
not I_25947 (I443982,I443974);
nor I_25948 (I443544,I443982,I443787);
nand I_25949 (I444013,I443982,I443632);
not I_25950 (I444030,I181648);
nand I_25951 (I444047,I444030,I443736);
nand I_25952 (I444064,I443982,I444047);
nand I_25953 (I443535,I444064,I444013);
nand I_25954 (I443532,I444047,I443931);
not I_25955 (I444136,I2866);
DFFARX1 I_25956 (I327028,I2859,I444136,I444162,);
and I_25957 (I444170,I444162,I327034);
DFFARX1 I_25958 (I444170,I2859,I444136,I444119,);
DFFARX1 I_25959 (I327040,I2859,I444136,I444210,);
not I_25960 (I444218,I327025);
not I_25961 (I444235,I327025);
nand I_25962 (I444252,I444235,I444218);
nor I_25963 (I444107,I444210,I444252);
DFFARX1 I_25964 (I444252,I2859,I444136,I444292,);
not I_25965 (I444128,I444292);
not I_25966 (I444314,I327043);
nand I_25967 (I444331,I444235,I444314);
DFFARX1 I_25968 (I444331,I2859,I444136,I444357,);
not I_25969 (I444365,I444357);
not I_25970 (I444382,I327037);
nand I_25971 (I444399,I444382,I327028);
and I_25972 (I444416,I444218,I444399);
nor I_25973 (I444433,I444331,I444416);
DFFARX1 I_25974 (I444433,I2859,I444136,I444104,);
DFFARX1 I_25975 (I444416,I2859,I444136,I444125,);
nor I_25976 (I444478,I327037,I327046);
nor I_25977 (I444116,I444331,I444478);
or I_25978 (I444509,I327037,I327046);
nor I_25979 (I444526,I327031,I327031);
DFFARX1 I_25980 (I444526,I2859,I444136,I444552,);
not I_25981 (I444560,I444552);
nor I_25982 (I444122,I444560,I444365);
nand I_25983 (I444591,I444560,I444210);
not I_25984 (I444608,I327031);
nand I_25985 (I444625,I444608,I444314);
nand I_25986 (I444642,I444560,I444625);
nand I_25987 (I444113,I444642,I444591);
nand I_25988 (I444110,I444625,I444509);
not I_25989 (I444714,I2866);
DFFARX1 I_25990 (I561822,I2859,I444714,I444740,);
and I_25991 (I444748,I444740,I561804);
DFFARX1 I_25992 (I444748,I2859,I444714,I444697,);
DFFARX1 I_25993 (I561795,I2859,I444714,I444788,);
not I_25994 (I444796,I561810);
not I_25995 (I444813,I561798);
nand I_25996 (I444830,I444813,I444796);
nor I_25997 (I444685,I444788,I444830);
DFFARX1 I_25998 (I444830,I2859,I444714,I444870,);
not I_25999 (I444706,I444870);
not I_26000 (I444892,I561807);
nand I_26001 (I444909,I444813,I444892);
DFFARX1 I_26002 (I444909,I2859,I444714,I444935,);
not I_26003 (I444943,I444935);
not I_26004 (I444960,I561816);
nand I_26005 (I444977,I444960,I561795);
and I_26006 (I444994,I444796,I444977);
nor I_26007 (I445011,I444909,I444994);
DFFARX1 I_26008 (I445011,I2859,I444714,I444682,);
DFFARX1 I_26009 (I444994,I2859,I444714,I444703,);
nor I_26010 (I445056,I561816,I561819);
nor I_26011 (I444694,I444909,I445056);
or I_26012 (I445087,I561816,I561819);
nor I_26013 (I445104,I561813,I561801);
DFFARX1 I_26014 (I445104,I2859,I444714,I445130,);
not I_26015 (I445138,I445130);
nor I_26016 (I444700,I445138,I444943);
nand I_26017 (I445169,I445138,I444788);
not I_26018 (I445186,I561813);
nand I_26019 (I445203,I445186,I444892);
nand I_26020 (I445220,I445138,I445203);
nand I_26021 (I444691,I445220,I445169);
nand I_26022 (I444688,I445203,I445087);
not I_26023 (I445292,I2866);
DFFARX1 I_26024 (I1444,I2859,I445292,I445318,);
and I_26025 (I445326,I445318,I1796);
DFFARX1 I_26026 (I445326,I2859,I445292,I445275,);
DFFARX1 I_26027 (I1836,I2859,I445292,I445366,);
not I_26028 (I445374,I1612);
not I_26029 (I445391,I2684);
nand I_26030 (I445408,I445391,I445374);
nor I_26031 (I445263,I445366,I445408);
DFFARX1 I_26032 (I445408,I2859,I445292,I445448,);
not I_26033 (I445284,I445448);
not I_26034 (I445470,I2596);
nand I_26035 (I445487,I445391,I445470);
DFFARX1 I_26036 (I445487,I2859,I445292,I445513,);
not I_26037 (I445521,I445513);
not I_26038 (I445538,I2012);
nand I_26039 (I445555,I445538,I2316);
and I_26040 (I445572,I445374,I445555);
nor I_26041 (I445589,I445487,I445572);
DFFARX1 I_26042 (I445589,I2859,I445292,I445260,);
DFFARX1 I_26043 (I445572,I2859,I445292,I445281,);
nor I_26044 (I445634,I2012,I2308);
nor I_26045 (I445272,I445487,I445634);
or I_26046 (I445665,I2012,I2308);
nor I_26047 (I445682,I2204,I2396);
DFFARX1 I_26048 (I445682,I2859,I445292,I445708,);
not I_26049 (I445716,I445708);
nor I_26050 (I445278,I445716,I445521);
nand I_26051 (I445747,I445716,I445366);
not I_26052 (I445764,I2204);
nand I_26053 (I445781,I445764,I445470);
nand I_26054 (I445798,I445716,I445781);
nand I_26055 (I445269,I445798,I445747);
nand I_26056 (I445266,I445781,I445665);
not I_26057 (I445870,I2866);
DFFARX1 I_26058 (I82242,I2859,I445870,I445896,);
and I_26059 (I445904,I445896,I82245);
DFFARX1 I_26060 (I445904,I2859,I445870,I445853,);
DFFARX1 I_26061 (I82245,I2859,I445870,I445944,);
not I_26062 (I445952,I82260);
not I_26063 (I445969,I82266);
nand I_26064 (I445986,I445969,I445952);
nor I_26065 (I445841,I445944,I445986);
DFFARX1 I_26066 (I445986,I2859,I445870,I446026,);
not I_26067 (I445862,I446026);
not I_26068 (I446048,I82254);
nand I_26069 (I446065,I445969,I446048);
DFFARX1 I_26070 (I446065,I2859,I445870,I446091,);
not I_26071 (I446099,I446091);
not I_26072 (I446116,I82251);
nand I_26073 (I446133,I446116,I82248);
and I_26074 (I446150,I445952,I446133);
nor I_26075 (I446167,I446065,I446150);
DFFARX1 I_26076 (I446167,I2859,I445870,I445838,);
DFFARX1 I_26077 (I446150,I2859,I445870,I445859,);
nor I_26078 (I446212,I82251,I82242);
nor I_26079 (I445850,I446065,I446212);
or I_26080 (I446243,I82251,I82242);
nor I_26081 (I446260,I82257,I82263);
DFFARX1 I_26082 (I446260,I2859,I445870,I446286,);
not I_26083 (I446294,I446286);
nor I_26084 (I445856,I446294,I446099);
nand I_26085 (I446325,I446294,I445944);
not I_26086 (I446342,I82257);
nand I_26087 (I446359,I446342,I446048);
nand I_26088 (I446376,I446294,I446359);
nand I_26089 (I445847,I446376,I446325);
nand I_26090 (I445844,I446359,I446243);
not I_26091 (I446448,I2866);
DFFARX1 I_26092 (I269529,I2859,I446448,I446474,);
and I_26093 (I446482,I446474,I269517);
DFFARX1 I_26094 (I446482,I2859,I446448,I446431,);
DFFARX1 I_26095 (I269520,I2859,I446448,I446522,);
not I_26096 (I446530,I269514);
not I_26097 (I446547,I269538);
nand I_26098 (I446564,I446547,I446530);
nor I_26099 (I446419,I446522,I446564);
DFFARX1 I_26100 (I446564,I2859,I446448,I446604,);
not I_26101 (I446440,I446604);
not I_26102 (I446626,I269526);
nand I_26103 (I446643,I446547,I446626);
DFFARX1 I_26104 (I446643,I2859,I446448,I446669,);
not I_26105 (I446677,I446669);
not I_26106 (I446694,I269535);
nand I_26107 (I446711,I446694,I269532);
and I_26108 (I446728,I446530,I446711);
nor I_26109 (I446745,I446643,I446728);
DFFARX1 I_26110 (I446745,I2859,I446448,I446416,);
DFFARX1 I_26111 (I446728,I2859,I446448,I446437,);
nor I_26112 (I446790,I269535,I269523);
nor I_26113 (I446428,I446643,I446790);
or I_26114 (I446821,I269535,I269523);
nor I_26115 (I446838,I269514,I269517);
DFFARX1 I_26116 (I446838,I2859,I446448,I446864,);
not I_26117 (I446872,I446864);
nor I_26118 (I446434,I446872,I446677);
nand I_26119 (I446903,I446872,I446522);
not I_26120 (I446920,I269514);
nand I_26121 (I446937,I446920,I446626);
nand I_26122 (I446954,I446872,I446937);
nand I_26123 (I446425,I446954,I446903);
nand I_26124 (I446422,I446937,I446821);
not I_26125 (I447026,I2866);
DFFARX1 I_26126 (I192504,I2859,I447026,I447052,);
and I_26127 (I447060,I447052,I192519);
DFFARX1 I_26128 (I447060,I2859,I447026,I447009,);
DFFARX1 I_26129 (I192522,I2859,I447026,I447100,);
not I_26130 (I447108,I192516);
not I_26131 (I447125,I192531);
nand I_26132 (I447142,I447125,I447108);
nor I_26133 (I446997,I447100,I447142);
DFFARX1 I_26134 (I447142,I2859,I447026,I447182,);
not I_26135 (I447018,I447182);
not I_26136 (I447204,I192507);
nand I_26137 (I447221,I447125,I447204);
DFFARX1 I_26138 (I447221,I2859,I447026,I447247,);
not I_26139 (I447255,I447247);
not I_26140 (I447272,I192510);
nand I_26141 (I447289,I447272,I192504);
and I_26142 (I447306,I447108,I447289);
nor I_26143 (I447323,I447221,I447306);
DFFARX1 I_26144 (I447323,I2859,I447026,I446994,);
DFFARX1 I_26145 (I447306,I2859,I447026,I447015,);
nor I_26146 (I447368,I192510,I192513);
nor I_26147 (I447006,I447221,I447368);
or I_26148 (I447399,I192510,I192513);
nor I_26149 (I447416,I192528,I192525);
DFFARX1 I_26150 (I447416,I2859,I447026,I447442,);
not I_26151 (I447450,I447442);
nor I_26152 (I447012,I447450,I447255);
nand I_26153 (I447481,I447450,I447100);
not I_26154 (I447498,I192528);
nand I_26155 (I447515,I447498,I447204);
nand I_26156 (I447532,I447450,I447515);
nand I_26157 (I447003,I447532,I447481);
nand I_26158 (I447000,I447515,I447399);
not I_26159 (I447604,I2866);
DFFARX1 I_26160 (I3479,I2859,I447604,I447630,);
and I_26161 (I447638,I447630,I3485);
DFFARX1 I_26162 (I447638,I2859,I447604,I447587,);
DFFARX1 I_26163 (I3464,I2859,I447604,I447678,);
not I_26164 (I447686,I3470);
not I_26165 (I447703,I3476);
nand I_26166 (I447720,I447703,I447686);
nor I_26167 (I447575,I447678,I447720);
DFFARX1 I_26168 (I447720,I2859,I447604,I447760,);
not I_26169 (I447596,I447760);
not I_26170 (I447782,I3467);
nand I_26171 (I447799,I447703,I447782);
DFFARX1 I_26172 (I447799,I2859,I447604,I447825,);
not I_26173 (I447833,I447825);
not I_26174 (I447850,I3482);
nand I_26175 (I447867,I447850,I3467);
and I_26176 (I447884,I447686,I447867);
nor I_26177 (I447901,I447799,I447884);
DFFARX1 I_26178 (I447901,I2859,I447604,I447572,);
DFFARX1 I_26179 (I447884,I2859,I447604,I447593,);
nor I_26180 (I447946,I3482,I3470);
nor I_26181 (I447584,I447799,I447946);
or I_26182 (I447977,I3482,I3470);
nor I_26183 (I447994,I3473,I3464);
DFFARX1 I_26184 (I447994,I2859,I447604,I448020,);
not I_26185 (I448028,I448020);
nor I_26186 (I447590,I448028,I447833);
nand I_26187 (I448059,I448028,I447678);
not I_26188 (I448076,I3473);
nand I_26189 (I448093,I448076,I447782);
nand I_26190 (I448110,I448028,I448093);
nand I_26191 (I447581,I448110,I448059);
nand I_26192 (I447578,I448093,I447977);
not I_26193 (I448182,I2866);
DFFARX1 I_26194 (I378609,I2859,I448182,I448208,);
and I_26195 (I448216,I448208,I378603);
DFFARX1 I_26196 (I448216,I2859,I448182,I448165,);
DFFARX1 I_26197 (I378621,I2859,I448182,I448256,);
not I_26198 (I448264,I378612);
not I_26199 (I448281,I378624);
nand I_26200 (I448298,I448281,I448264);
nor I_26201 (I448153,I448256,I448298);
DFFARX1 I_26202 (I448298,I2859,I448182,I448338,);
not I_26203 (I448174,I448338);
not I_26204 (I448360,I378630);
nand I_26205 (I448377,I448281,I448360);
DFFARX1 I_26206 (I448377,I2859,I448182,I448403,);
not I_26207 (I448411,I448403);
not I_26208 (I448428,I378606);
nand I_26209 (I448445,I448428,I378627);
and I_26210 (I448462,I448264,I448445);
nor I_26211 (I448479,I448377,I448462);
DFFARX1 I_26212 (I448479,I2859,I448182,I448150,);
DFFARX1 I_26213 (I448462,I2859,I448182,I448171,);
nor I_26214 (I448524,I378606,I378618);
nor I_26215 (I448162,I448377,I448524);
or I_26216 (I448555,I378606,I378618);
nor I_26217 (I448572,I378603,I378615);
DFFARX1 I_26218 (I448572,I2859,I448182,I448598,);
not I_26219 (I448606,I448598);
nor I_26220 (I448168,I448606,I448411);
nand I_26221 (I448637,I448606,I448256);
not I_26222 (I448654,I378603);
nand I_26223 (I448671,I448654,I448360);
nand I_26224 (I448688,I448606,I448671);
nand I_26225 (I448159,I448688,I448637);
nand I_26226 (I448156,I448671,I448555);
not I_26227 (I448760,I2866);
DFFARX1 I_26228 (I118802,I2859,I448760,I448786,);
and I_26229 (I448794,I448786,I118787);
DFFARX1 I_26230 (I448794,I2859,I448760,I448743,);
DFFARX1 I_26231 (I118793,I2859,I448760,I448834,);
not I_26232 (I448842,I118775);
not I_26233 (I448859,I118796);
nand I_26234 (I448876,I448859,I448842);
nor I_26235 (I448731,I448834,I448876);
DFFARX1 I_26236 (I448876,I2859,I448760,I448916,);
not I_26237 (I448752,I448916);
not I_26238 (I448938,I118799);
nand I_26239 (I448955,I448859,I448938);
DFFARX1 I_26240 (I448955,I2859,I448760,I448981,);
not I_26241 (I448989,I448981);
not I_26242 (I449006,I118790);
nand I_26243 (I449023,I449006,I118778);
and I_26244 (I449040,I448842,I449023);
nor I_26245 (I449057,I448955,I449040);
DFFARX1 I_26246 (I449057,I2859,I448760,I448728,);
DFFARX1 I_26247 (I449040,I2859,I448760,I448749,);
nor I_26248 (I449102,I118790,I118784);
nor I_26249 (I448740,I448955,I449102);
or I_26250 (I449133,I118790,I118784);
nor I_26251 (I449150,I118781,I118775);
DFFARX1 I_26252 (I449150,I2859,I448760,I449176,);
not I_26253 (I449184,I449176);
nor I_26254 (I448746,I449184,I448989);
nand I_26255 (I449215,I449184,I448834);
not I_26256 (I449232,I118781);
nand I_26257 (I449249,I449232,I448938);
nand I_26258 (I449266,I449184,I449249);
nand I_26259 (I448737,I449266,I449215);
nand I_26260 (I448734,I449249,I449133);
not I_26261 (I449338,I2866);
DFFARX1 I_26262 (I166936,I2859,I449338,I449364,);
and I_26263 (I449372,I449364,I166951);
DFFARX1 I_26264 (I449372,I2859,I449338,I449321,);
DFFARX1 I_26265 (I166954,I2859,I449338,I449412,);
not I_26266 (I449420,I166948);
not I_26267 (I449437,I166963);
nand I_26268 (I449454,I449437,I449420);
nor I_26269 (I449309,I449412,I449454);
DFFARX1 I_26270 (I449454,I2859,I449338,I449494,);
not I_26271 (I449330,I449494);
not I_26272 (I449516,I166939);
nand I_26273 (I449533,I449437,I449516);
DFFARX1 I_26274 (I449533,I2859,I449338,I449559,);
not I_26275 (I449567,I449559);
not I_26276 (I449584,I166942);
nand I_26277 (I449601,I449584,I166936);
and I_26278 (I449618,I449420,I449601);
nor I_26279 (I449635,I449533,I449618);
DFFARX1 I_26280 (I449635,I2859,I449338,I449306,);
DFFARX1 I_26281 (I449618,I2859,I449338,I449327,);
nor I_26282 (I449680,I166942,I166945);
nor I_26283 (I449318,I449533,I449680);
or I_26284 (I449711,I166942,I166945);
nor I_26285 (I449728,I166960,I166957);
DFFARX1 I_26286 (I449728,I2859,I449338,I449754,);
not I_26287 (I449762,I449754);
nor I_26288 (I449324,I449762,I449567);
nand I_26289 (I449793,I449762,I449412);
not I_26290 (I449810,I166960);
nand I_26291 (I449827,I449810,I449516);
nand I_26292 (I449844,I449762,I449827);
nand I_26293 (I449315,I449844,I449793);
nand I_26294 (I449312,I449827,I449711);
not I_26295 (I449916,I2866);
DFFARX1 I_26296 (I156746,I2859,I449916,I449942,);
and I_26297 (I449950,I449942,I156731);
DFFARX1 I_26298 (I449950,I2859,I449916,I449899,);
DFFARX1 I_26299 (I156737,I2859,I449916,I449990,);
not I_26300 (I449998,I156719);
not I_26301 (I450015,I156740);
nand I_26302 (I450032,I450015,I449998);
nor I_26303 (I449887,I449990,I450032);
DFFARX1 I_26304 (I450032,I2859,I449916,I450072,);
not I_26305 (I449908,I450072);
not I_26306 (I450094,I156743);
nand I_26307 (I450111,I450015,I450094);
DFFARX1 I_26308 (I450111,I2859,I449916,I450137,);
not I_26309 (I450145,I450137);
not I_26310 (I450162,I156734);
nand I_26311 (I450179,I450162,I156722);
and I_26312 (I450196,I449998,I450179);
nor I_26313 (I450213,I450111,I450196);
DFFARX1 I_26314 (I450213,I2859,I449916,I449884,);
DFFARX1 I_26315 (I450196,I2859,I449916,I449905,);
nor I_26316 (I450258,I156734,I156728);
nor I_26317 (I449896,I450111,I450258);
or I_26318 (I450289,I156734,I156728);
nor I_26319 (I450306,I156725,I156719);
DFFARX1 I_26320 (I450306,I2859,I449916,I450332,);
not I_26321 (I450340,I450332);
nor I_26322 (I449902,I450340,I450145);
nand I_26323 (I450371,I450340,I449990);
not I_26324 (I450388,I156725);
nand I_26325 (I450405,I450388,I450094);
nand I_26326 (I450422,I450340,I450405);
nand I_26327 (I449893,I450422,I450371);
nand I_26328 (I449890,I450405,I450289);
not I_26329 (I450494,I2866);
DFFARX1 I_26330 (I318069,I2859,I450494,I450520,);
and I_26331 (I450528,I450520,I318075);
DFFARX1 I_26332 (I450528,I2859,I450494,I450477,);
DFFARX1 I_26333 (I318081,I2859,I450494,I450568,);
not I_26334 (I450576,I318066);
not I_26335 (I450593,I318066);
nand I_26336 (I450610,I450593,I450576);
nor I_26337 (I450465,I450568,I450610);
DFFARX1 I_26338 (I450610,I2859,I450494,I450650,);
not I_26339 (I450486,I450650);
not I_26340 (I450672,I318084);
nand I_26341 (I450689,I450593,I450672);
DFFARX1 I_26342 (I450689,I2859,I450494,I450715,);
not I_26343 (I450723,I450715);
not I_26344 (I450740,I318078);
nand I_26345 (I450757,I450740,I318069);
and I_26346 (I450774,I450576,I450757);
nor I_26347 (I450791,I450689,I450774);
DFFARX1 I_26348 (I450791,I2859,I450494,I450462,);
DFFARX1 I_26349 (I450774,I2859,I450494,I450483,);
nor I_26350 (I450836,I318078,I318087);
nor I_26351 (I450474,I450689,I450836);
or I_26352 (I450867,I318078,I318087);
nor I_26353 (I450884,I318072,I318072);
DFFARX1 I_26354 (I450884,I2859,I450494,I450910,);
not I_26355 (I450918,I450910);
nor I_26356 (I450480,I450918,I450723);
nand I_26357 (I450949,I450918,I450568);
not I_26358 (I450966,I318072);
nand I_26359 (I450983,I450966,I450672);
nand I_26360 (I451000,I450918,I450983);
nand I_26361 (I450471,I451000,I450949);
nand I_26362 (I450468,I450983,I450867);
not I_26363 (I451072,I2866);
DFFARX1 I_26364 (I230803,I2859,I451072,I451098,);
and I_26365 (I451106,I451098,I230791);
DFFARX1 I_26366 (I451106,I2859,I451072,I451055,);
DFFARX1 I_26367 (I230806,I2859,I451072,I451146,);
not I_26368 (I451154,I230797);
not I_26369 (I451171,I230788);
nand I_26370 (I451188,I451171,I451154);
nor I_26371 (I451043,I451146,I451188);
DFFARX1 I_26372 (I451188,I2859,I451072,I451228,);
not I_26373 (I451064,I451228);
not I_26374 (I451250,I230794);
nand I_26375 (I451267,I451171,I451250);
DFFARX1 I_26376 (I451267,I2859,I451072,I451293,);
not I_26377 (I451301,I451293);
not I_26378 (I451318,I230809);
nand I_26379 (I451335,I451318,I230812);
and I_26380 (I451352,I451154,I451335);
nor I_26381 (I451369,I451267,I451352);
DFFARX1 I_26382 (I451369,I2859,I451072,I451040,);
DFFARX1 I_26383 (I451352,I2859,I451072,I451061,);
nor I_26384 (I451414,I230809,I230788);
nor I_26385 (I451052,I451267,I451414);
or I_26386 (I451445,I230809,I230788);
nor I_26387 (I451462,I230800,I230791);
DFFARX1 I_26388 (I451462,I2859,I451072,I451488,);
not I_26389 (I451496,I451488);
nor I_26390 (I451058,I451496,I451301);
nand I_26391 (I451527,I451496,I451146);
not I_26392 (I451544,I230800);
nand I_26393 (I451561,I451544,I451250);
nand I_26394 (I451578,I451496,I451561);
nand I_26395 (I451049,I451578,I451527);
nand I_26396 (I451046,I451561,I451445);
not I_26397 (I451650,I2866);
DFFARX1 I_26398 (I555872,I2859,I451650,I451676,);
and I_26399 (I451684,I451676,I555854);
DFFARX1 I_26400 (I451684,I2859,I451650,I451633,);
DFFARX1 I_26401 (I555845,I2859,I451650,I451724,);
not I_26402 (I451732,I555860);
not I_26403 (I451749,I555848);
nand I_26404 (I451766,I451749,I451732);
nor I_26405 (I451621,I451724,I451766);
DFFARX1 I_26406 (I451766,I2859,I451650,I451806,);
not I_26407 (I451642,I451806);
not I_26408 (I451828,I555857);
nand I_26409 (I451845,I451749,I451828);
DFFARX1 I_26410 (I451845,I2859,I451650,I451871,);
not I_26411 (I451879,I451871);
not I_26412 (I451896,I555866);
nand I_26413 (I451913,I451896,I555845);
and I_26414 (I451930,I451732,I451913);
nor I_26415 (I451947,I451845,I451930);
DFFARX1 I_26416 (I451947,I2859,I451650,I451618,);
DFFARX1 I_26417 (I451930,I2859,I451650,I451639,);
nor I_26418 (I451992,I555866,I555869);
nor I_26419 (I451630,I451845,I451992);
or I_26420 (I452023,I555866,I555869);
nor I_26421 (I452040,I555863,I555851);
DFFARX1 I_26422 (I452040,I2859,I451650,I452066,);
not I_26423 (I452074,I452066);
nor I_26424 (I451636,I452074,I451879);
nand I_26425 (I452105,I452074,I451724);
not I_26426 (I452122,I555863);
nand I_26427 (I452139,I452122,I451828);
nand I_26428 (I452156,I452074,I452139);
nand I_26429 (I451627,I452156,I452105);
nand I_26430 (I451624,I452139,I452023);
not I_26431 (I452228,I2866);
DFFARX1 I_26432 (I212618,I2859,I452228,I452254,);
and I_26433 (I452262,I452254,I212633);
DFFARX1 I_26434 (I452262,I2859,I452228,I452211,);
DFFARX1 I_26435 (I212624,I2859,I452228,I452302,);
not I_26436 (I452310,I212618);
not I_26437 (I452327,I212636);
nand I_26438 (I452344,I452327,I452310);
nor I_26439 (I452199,I452302,I452344);
DFFARX1 I_26440 (I452344,I2859,I452228,I452384,);
not I_26441 (I452220,I452384);
not I_26442 (I452406,I212627);
nand I_26443 (I452423,I452327,I452406);
DFFARX1 I_26444 (I452423,I2859,I452228,I452449,);
not I_26445 (I452457,I452449);
not I_26446 (I452474,I212639);
nand I_26447 (I452491,I452474,I212615);
and I_26448 (I452508,I452310,I452491);
nor I_26449 (I452525,I452423,I452508);
DFFARX1 I_26450 (I452525,I2859,I452228,I452196,);
DFFARX1 I_26451 (I452508,I2859,I452228,I452217,);
nor I_26452 (I452570,I212639,I212615);
nor I_26453 (I452208,I452423,I452570);
or I_26454 (I452601,I212639,I212615);
nor I_26455 (I452618,I212621,I212630);
DFFARX1 I_26456 (I452618,I2859,I452228,I452644,);
not I_26457 (I452652,I452644);
nor I_26458 (I452214,I452652,I452457);
nand I_26459 (I452683,I452652,I452302);
not I_26460 (I452700,I212621);
nand I_26461 (I452717,I452700,I452406);
nand I_26462 (I452734,I452652,I452717);
nand I_26463 (I452205,I452734,I452683);
nand I_26464 (I452202,I452717,I452601);
not I_26465 (I452806,I2866);
DFFARX1 I_26466 (I222711,I2859,I452806,I452832,);
and I_26467 (I452840,I452832,I222699);
DFFARX1 I_26468 (I452840,I2859,I452806,I452789,);
DFFARX1 I_26469 (I222714,I2859,I452806,I452880,);
not I_26470 (I452888,I222705);
not I_26471 (I452905,I222696);
nand I_26472 (I452922,I452905,I452888);
nor I_26473 (I452777,I452880,I452922);
DFFARX1 I_26474 (I452922,I2859,I452806,I452962,);
not I_26475 (I452798,I452962);
not I_26476 (I452984,I222702);
nand I_26477 (I453001,I452905,I452984);
DFFARX1 I_26478 (I453001,I2859,I452806,I453027,);
not I_26479 (I453035,I453027);
not I_26480 (I453052,I222717);
nand I_26481 (I453069,I453052,I222720);
and I_26482 (I453086,I452888,I453069);
nor I_26483 (I453103,I453001,I453086);
DFFARX1 I_26484 (I453103,I2859,I452806,I452774,);
DFFARX1 I_26485 (I453086,I2859,I452806,I452795,);
nor I_26486 (I453148,I222717,I222696);
nor I_26487 (I452786,I453001,I453148);
or I_26488 (I453179,I222717,I222696);
nor I_26489 (I453196,I222708,I222699);
DFFARX1 I_26490 (I453196,I2859,I452806,I453222,);
not I_26491 (I453230,I453222);
nor I_26492 (I452792,I453230,I453035);
nand I_26493 (I453261,I453230,I452880);
not I_26494 (I453278,I222708);
nand I_26495 (I453295,I453278,I452984);
nand I_26496 (I453312,I453230,I453295);
nand I_26497 (I452783,I453312,I453261);
nand I_26498 (I452780,I453295,I453179);
not I_26499 (I453384,I2866);
DFFARX1 I_26500 (I272419,I2859,I453384,I453410,);
and I_26501 (I453418,I453410,I272407);
DFFARX1 I_26502 (I453418,I2859,I453384,I453367,);
DFFARX1 I_26503 (I272410,I2859,I453384,I453458,);
not I_26504 (I453466,I272404);
not I_26505 (I453483,I272428);
nand I_26506 (I453500,I453483,I453466);
nor I_26507 (I453355,I453458,I453500);
DFFARX1 I_26508 (I453500,I2859,I453384,I453540,);
not I_26509 (I453376,I453540);
not I_26510 (I453562,I272416);
nand I_26511 (I453579,I453483,I453562);
DFFARX1 I_26512 (I453579,I2859,I453384,I453605,);
not I_26513 (I453613,I453605);
not I_26514 (I453630,I272425);
nand I_26515 (I453647,I453630,I272422);
and I_26516 (I453664,I453466,I453647);
nor I_26517 (I453681,I453579,I453664);
DFFARX1 I_26518 (I453681,I2859,I453384,I453352,);
DFFARX1 I_26519 (I453664,I2859,I453384,I453373,);
nor I_26520 (I453726,I272425,I272413);
nor I_26521 (I453364,I453579,I453726);
or I_26522 (I453757,I272425,I272413);
nor I_26523 (I453774,I272404,I272407);
DFFARX1 I_26524 (I453774,I2859,I453384,I453800,);
not I_26525 (I453808,I453800);
nor I_26526 (I453370,I453808,I453613);
nand I_26527 (I453839,I453808,I453458);
not I_26528 (I453856,I272404);
nand I_26529 (I453873,I453856,I453562);
nand I_26530 (I453890,I453808,I453873);
nand I_26531 (I453361,I453890,I453839);
nand I_26532 (I453358,I453873,I453757);
not I_26533 (I453962,I2866);
DFFARX1 I_26534 (I251033,I2859,I453962,I453988,);
and I_26535 (I453996,I453988,I251021);
DFFARX1 I_26536 (I453996,I2859,I453962,I453945,);
DFFARX1 I_26537 (I251036,I2859,I453962,I454036,);
not I_26538 (I454044,I251027);
not I_26539 (I454061,I251018);
nand I_26540 (I454078,I454061,I454044);
nor I_26541 (I453933,I454036,I454078);
DFFARX1 I_26542 (I454078,I2859,I453962,I454118,);
not I_26543 (I453954,I454118);
not I_26544 (I454140,I251024);
nand I_26545 (I454157,I454061,I454140);
DFFARX1 I_26546 (I454157,I2859,I453962,I454183,);
not I_26547 (I454191,I454183);
not I_26548 (I454208,I251039);
nand I_26549 (I454225,I454208,I251042);
and I_26550 (I454242,I454044,I454225);
nor I_26551 (I454259,I454157,I454242);
DFFARX1 I_26552 (I454259,I2859,I453962,I453930,);
DFFARX1 I_26553 (I454242,I2859,I453962,I453951,);
nor I_26554 (I454304,I251039,I251018);
nor I_26555 (I453942,I454157,I454304);
or I_26556 (I454335,I251039,I251018);
nor I_26557 (I454352,I251030,I251021);
DFFARX1 I_26558 (I454352,I2859,I453962,I454378,);
not I_26559 (I454386,I454378);
nor I_26560 (I453948,I454386,I454191);
nand I_26561 (I454417,I454386,I454036);
not I_26562 (I454434,I251030);
nand I_26563 (I454451,I454434,I454140);
nand I_26564 (I454468,I454386,I454451);
nand I_26565 (I453939,I454468,I454417);
nand I_26566 (I453936,I454451,I454335);
not I_26567 (I454540,I2866);
DFFARX1 I_26568 (I95332,I2859,I454540,I454566,);
and I_26569 (I454574,I454566,I95335);
DFFARX1 I_26570 (I454574,I2859,I454540,I454523,);
DFFARX1 I_26571 (I95335,I2859,I454540,I454614,);
not I_26572 (I454622,I95350);
not I_26573 (I454639,I95356);
nand I_26574 (I454656,I454639,I454622);
nor I_26575 (I454511,I454614,I454656);
DFFARX1 I_26576 (I454656,I2859,I454540,I454696,);
not I_26577 (I454532,I454696);
not I_26578 (I454718,I95344);
nand I_26579 (I454735,I454639,I454718);
DFFARX1 I_26580 (I454735,I2859,I454540,I454761,);
not I_26581 (I454769,I454761);
not I_26582 (I454786,I95341);
nand I_26583 (I454803,I454786,I95338);
and I_26584 (I454820,I454622,I454803);
nor I_26585 (I454837,I454735,I454820);
DFFARX1 I_26586 (I454837,I2859,I454540,I454508,);
DFFARX1 I_26587 (I454820,I2859,I454540,I454529,);
nor I_26588 (I454882,I95341,I95332);
nor I_26589 (I454520,I454735,I454882);
or I_26590 (I454913,I95341,I95332);
nor I_26591 (I454930,I95347,I95353);
DFFARX1 I_26592 (I454930,I2859,I454540,I454956,);
not I_26593 (I454964,I454956);
nor I_26594 (I454526,I454964,I454769);
nand I_26595 (I454995,I454964,I454614);
not I_26596 (I455012,I95347);
nand I_26597 (I455029,I455012,I454718);
nand I_26598 (I455046,I454964,I455029);
nand I_26599 (I454517,I455046,I454995);
nand I_26600 (I454514,I455029,I454913);
not I_26601 (I455118,I2866);
DFFARX1 I_26602 (I131977,I2859,I455118,I455144,);
and I_26603 (I455152,I455144,I131962);
DFFARX1 I_26604 (I455152,I2859,I455118,I455101,);
DFFARX1 I_26605 (I131968,I2859,I455118,I455192,);
not I_26606 (I455200,I131950);
not I_26607 (I455217,I131971);
nand I_26608 (I455234,I455217,I455200);
nor I_26609 (I455089,I455192,I455234);
DFFARX1 I_26610 (I455234,I2859,I455118,I455274,);
not I_26611 (I455110,I455274);
not I_26612 (I455296,I131974);
nand I_26613 (I455313,I455217,I455296);
DFFARX1 I_26614 (I455313,I2859,I455118,I455339,);
not I_26615 (I455347,I455339);
not I_26616 (I455364,I131965);
nand I_26617 (I455381,I455364,I131953);
and I_26618 (I455398,I455200,I455381);
nor I_26619 (I455415,I455313,I455398);
DFFARX1 I_26620 (I455415,I2859,I455118,I455086,);
DFFARX1 I_26621 (I455398,I2859,I455118,I455107,);
nor I_26622 (I455460,I131965,I131959);
nor I_26623 (I455098,I455313,I455460);
or I_26624 (I455491,I131965,I131959);
nor I_26625 (I455508,I131956,I131950);
DFFARX1 I_26626 (I455508,I2859,I455118,I455534,);
not I_26627 (I455542,I455534);
nor I_26628 (I455104,I455542,I455347);
nand I_26629 (I455573,I455542,I455192);
not I_26630 (I455590,I131956);
nand I_26631 (I455607,I455590,I455296);
nand I_26632 (I455624,I455542,I455607);
nand I_26633 (I455095,I455624,I455573);
nand I_26634 (I455092,I455607,I455491);
not I_26635 (I455696,I2866);
DFFARX1 I_26636 (I226757,I2859,I455696,I455722,);
and I_26637 (I455730,I455722,I226745);
DFFARX1 I_26638 (I455730,I2859,I455696,I455679,);
DFFARX1 I_26639 (I226760,I2859,I455696,I455770,);
not I_26640 (I455778,I226751);
not I_26641 (I455795,I226742);
nand I_26642 (I455812,I455795,I455778);
nor I_26643 (I455667,I455770,I455812);
DFFARX1 I_26644 (I455812,I2859,I455696,I455852,);
not I_26645 (I455688,I455852);
not I_26646 (I455874,I226748);
nand I_26647 (I455891,I455795,I455874);
DFFARX1 I_26648 (I455891,I2859,I455696,I455917,);
not I_26649 (I455925,I455917);
not I_26650 (I455942,I226763);
nand I_26651 (I455959,I455942,I226766);
and I_26652 (I455976,I455778,I455959);
nor I_26653 (I455993,I455891,I455976);
DFFARX1 I_26654 (I455993,I2859,I455696,I455664,);
DFFARX1 I_26655 (I455976,I2859,I455696,I455685,);
nor I_26656 (I456038,I226763,I226742);
nor I_26657 (I455676,I455891,I456038);
or I_26658 (I456069,I226763,I226742);
nor I_26659 (I456086,I226754,I226745);
DFFARX1 I_26660 (I456086,I2859,I455696,I456112,);
not I_26661 (I456120,I456112);
nor I_26662 (I455682,I456120,I455925);
nand I_26663 (I456151,I456120,I455770);
not I_26664 (I456168,I226754);
nand I_26665 (I456185,I456168,I455874);
nand I_26666 (I456202,I456120,I456185);
nand I_26667 (I455673,I456202,I456151);
nand I_26668 (I455670,I456185,I456069);
not I_26669 (I456274,I2866);
DFFARX1 I_26670 (I226179,I2859,I456274,I456300,);
and I_26671 (I456308,I456300,I226167);
DFFARX1 I_26672 (I456308,I2859,I456274,I456257,);
DFFARX1 I_26673 (I226182,I2859,I456274,I456348,);
not I_26674 (I456356,I226173);
not I_26675 (I456373,I226164);
nand I_26676 (I456390,I456373,I456356);
nor I_26677 (I456245,I456348,I456390);
DFFARX1 I_26678 (I456390,I2859,I456274,I456430,);
not I_26679 (I456266,I456430);
not I_26680 (I456452,I226170);
nand I_26681 (I456469,I456373,I456452);
DFFARX1 I_26682 (I456469,I2859,I456274,I456495,);
not I_26683 (I456503,I456495);
not I_26684 (I456520,I226185);
nand I_26685 (I456537,I456520,I226188);
and I_26686 (I456554,I456356,I456537);
nor I_26687 (I456571,I456469,I456554);
DFFARX1 I_26688 (I456571,I2859,I456274,I456242,);
DFFARX1 I_26689 (I456554,I2859,I456274,I456263,);
nor I_26690 (I456616,I226185,I226164);
nor I_26691 (I456254,I456469,I456616);
or I_26692 (I456647,I226185,I226164);
nor I_26693 (I456664,I226176,I226167);
DFFARX1 I_26694 (I456664,I2859,I456274,I456690,);
not I_26695 (I456698,I456690);
nor I_26696 (I456260,I456698,I456503);
nand I_26697 (I456729,I456698,I456348);
not I_26698 (I456746,I226176);
nand I_26699 (I456763,I456746,I456452);
nand I_26700 (I456780,I456698,I456763);
nand I_26701 (I456251,I456780,I456729);
nand I_26702 (I456248,I456763,I456647);
not I_26703 (I456852,I2866);
DFFARX1 I_26704 (I337568,I2859,I456852,I456878,);
and I_26705 (I456886,I456878,I337574);
DFFARX1 I_26706 (I456886,I2859,I456852,I456835,);
DFFARX1 I_26707 (I337580,I2859,I456852,I456926,);
not I_26708 (I456934,I337565);
not I_26709 (I456951,I337565);
nand I_26710 (I456968,I456951,I456934);
nor I_26711 (I456823,I456926,I456968);
DFFARX1 I_26712 (I456968,I2859,I456852,I457008,);
not I_26713 (I456844,I457008);
not I_26714 (I457030,I337583);
nand I_26715 (I457047,I456951,I457030);
DFFARX1 I_26716 (I457047,I2859,I456852,I457073,);
not I_26717 (I457081,I457073);
not I_26718 (I457098,I337577);
nand I_26719 (I457115,I457098,I337568);
and I_26720 (I457132,I456934,I457115);
nor I_26721 (I457149,I457047,I457132);
DFFARX1 I_26722 (I457149,I2859,I456852,I456820,);
DFFARX1 I_26723 (I457132,I2859,I456852,I456841,);
nor I_26724 (I457194,I337577,I337586);
nor I_26725 (I456832,I457047,I457194);
or I_26726 (I457225,I337577,I337586);
nor I_26727 (I457242,I337571,I337571);
DFFARX1 I_26728 (I457242,I2859,I456852,I457268,);
not I_26729 (I457276,I457268);
nor I_26730 (I456838,I457276,I457081);
nand I_26731 (I457307,I457276,I456926);
not I_26732 (I457324,I337571);
nand I_26733 (I457341,I457324,I457030);
nand I_26734 (I457358,I457276,I457341);
nand I_26735 (I456829,I457358,I457307);
nand I_26736 (I456826,I457341,I457225);
not I_26737 (I457430,I2866);
DFFARX1 I_26738 (I154638,I2859,I457430,I457456,);
and I_26739 (I457464,I457456,I154623);
DFFARX1 I_26740 (I457464,I2859,I457430,I457413,);
DFFARX1 I_26741 (I154629,I2859,I457430,I457504,);
not I_26742 (I457512,I154611);
not I_26743 (I457529,I154632);
nand I_26744 (I457546,I457529,I457512);
nor I_26745 (I457401,I457504,I457546);
DFFARX1 I_26746 (I457546,I2859,I457430,I457586,);
not I_26747 (I457422,I457586);
not I_26748 (I457608,I154635);
nand I_26749 (I457625,I457529,I457608);
DFFARX1 I_26750 (I457625,I2859,I457430,I457651,);
not I_26751 (I457659,I457651);
not I_26752 (I457676,I154626);
nand I_26753 (I457693,I457676,I154614);
and I_26754 (I457710,I457512,I457693);
nor I_26755 (I457727,I457625,I457710);
DFFARX1 I_26756 (I457727,I2859,I457430,I457398,);
DFFARX1 I_26757 (I457710,I2859,I457430,I457419,);
nor I_26758 (I457772,I154626,I154620);
nor I_26759 (I457410,I457625,I457772);
or I_26760 (I457803,I154626,I154620);
nor I_26761 (I457820,I154617,I154611);
DFFARX1 I_26762 (I457820,I2859,I457430,I457846,);
not I_26763 (I457854,I457846);
nor I_26764 (I457416,I457854,I457659);
nand I_26765 (I457885,I457854,I457504);
not I_26766 (I457902,I154617);
nand I_26767 (I457919,I457902,I457608);
nand I_26768 (I457936,I457854,I457919);
nand I_26769 (I457407,I457936,I457885);
nand I_26770 (I457404,I457919,I457803);
not I_26771 (I458008,I2866);
DFFARX1 I_26772 (I20624,I2859,I458008,I458034,);
and I_26773 (I458042,I458034,I20600);
DFFARX1 I_26774 (I458042,I2859,I458008,I457991,);
DFFARX1 I_26775 (I20618,I2859,I458008,I458082,);
not I_26776 (I458090,I20606);
not I_26777 (I458107,I20603);
nand I_26778 (I458124,I458107,I458090);
nor I_26779 (I457979,I458082,I458124);
DFFARX1 I_26780 (I458124,I2859,I458008,I458164,);
not I_26781 (I458000,I458164);
not I_26782 (I458186,I20612);
nand I_26783 (I458203,I458107,I458186);
DFFARX1 I_26784 (I458203,I2859,I458008,I458229,);
not I_26785 (I458237,I458229);
not I_26786 (I458254,I20603);
nand I_26787 (I458271,I458254,I20621);
and I_26788 (I458288,I458090,I458271);
nor I_26789 (I458305,I458203,I458288);
DFFARX1 I_26790 (I458305,I2859,I458008,I457976,);
DFFARX1 I_26791 (I458288,I2859,I458008,I457997,);
nor I_26792 (I458350,I20603,I20615);
nor I_26793 (I457988,I458203,I458350);
or I_26794 (I458381,I20603,I20615);
nor I_26795 (I458398,I20609,I20600);
DFFARX1 I_26796 (I458398,I2859,I458008,I458424,);
not I_26797 (I458432,I458424);
nor I_26798 (I457994,I458432,I458237);
nand I_26799 (I458463,I458432,I458082);
not I_26800 (I458480,I20609);
nand I_26801 (I458497,I458480,I458186);
nand I_26802 (I458514,I458432,I458497);
nand I_26803 (I457985,I458514,I458463);
nand I_26804 (I457982,I458497,I458381);
not I_26805 (I458586,I2866);
DFFARX1 I_26806 (I516647,I2859,I458586,I458612,);
and I_26807 (I458620,I458612,I516641);
DFFARX1 I_26808 (I458620,I2859,I458586,I458569,);
DFFARX1 I_26809 (I516626,I2859,I458586,I458660,);
not I_26810 (I458668,I516632);
not I_26811 (I458685,I516644);
nand I_26812 (I458702,I458685,I458668);
nor I_26813 (I458557,I458660,I458702);
DFFARX1 I_26814 (I458702,I2859,I458586,I458742,);
not I_26815 (I458578,I458742);
not I_26816 (I458764,I516626);
nand I_26817 (I458781,I458685,I458764);
DFFARX1 I_26818 (I458781,I2859,I458586,I458807,);
not I_26819 (I458815,I458807);
not I_26820 (I458832,I516650);
nand I_26821 (I458849,I458832,I516638);
and I_26822 (I458866,I458668,I458849);
nor I_26823 (I458883,I458781,I458866);
DFFARX1 I_26824 (I458883,I2859,I458586,I458554,);
DFFARX1 I_26825 (I458866,I2859,I458586,I458575,);
nor I_26826 (I458928,I516650,I516629);
nor I_26827 (I458566,I458781,I458928);
or I_26828 (I458959,I516650,I516629);
nor I_26829 (I458976,I516635,I516629);
DFFARX1 I_26830 (I458976,I2859,I458586,I459002,);
not I_26831 (I459010,I459002);
nor I_26832 (I458572,I459010,I458815);
nand I_26833 (I459041,I459010,I458660);
not I_26834 (I459058,I516635);
nand I_26835 (I459075,I459058,I458764);
nand I_26836 (I459092,I459010,I459075);
nand I_26837 (I458563,I459092,I459041);
nand I_26838 (I458560,I459075,I458959);
not I_26839 (I459164,I2866);
DFFARX1 I_26840 (I118275,I2859,I459164,I459190,);
and I_26841 (I459198,I459190,I118260);
DFFARX1 I_26842 (I459198,I2859,I459164,I459147,);
DFFARX1 I_26843 (I118266,I2859,I459164,I459238,);
not I_26844 (I459246,I118248);
not I_26845 (I459263,I118269);
nand I_26846 (I459280,I459263,I459246);
nor I_26847 (I459135,I459238,I459280);
DFFARX1 I_26848 (I459280,I2859,I459164,I459320,);
not I_26849 (I459156,I459320);
not I_26850 (I459342,I118272);
nand I_26851 (I459359,I459263,I459342);
DFFARX1 I_26852 (I459359,I2859,I459164,I459385,);
not I_26853 (I459393,I459385);
not I_26854 (I459410,I118263);
nand I_26855 (I459427,I459410,I118251);
and I_26856 (I459444,I459246,I459427);
nor I_26857 (I459461,I459359,I459444);
DFFARX1 I_26858 (I459461,I2859,I459164,I459132,);
DFFARX1 I_26859 (I459444,I2859,I459164,I459153,);
nor I_26860 (I459506,I118263,I118257);
nor I_26861 (I459144,I459359,I459506);
or I_26862 (I459537,I118263,I118257);
nor I_26863 (I459554,I118254,I118248);
DFFARX1 I_26864 (I459554,I2859,I459164,I459580,);
not I_26865 (I459588,I459580);
nor I_26866 (I459150,I459588,I459393);
nand I_26867 (I459619,I459588,I459238);
not I_26868 (I459636,I118254);
nand I_26869 (I459653,I459636,I459342);
nand I_26870 (I459670,I459588,I459653);
nand I_26871 (I459141,I459670,I459619);
nand I_26872 (I459138,I459653,I459537);
not I_26873 (I459742,I2866);
DFFARX1 I_26874 (I244097,I2859,I459742,I459768,);
and I_26875 (I459776,I459768,I244085);
DFFARX1 I_26876 (I459776,I2859,I459742,I459725,);
DFFARX1 I_26877 (I244100,I2859,I459742,I459816,);
not I_26878 (I459824,I244091);
not I_26879 (I459841,I244082);
nand I_26880 (I459858,I459841,I459824);
nor I_26881 (I459713,I459816,I459858);
DFFARX1 I_26882 (I459858,I2859,I459742,I459898,);
not I_26883 (I459734,I459898);
not I_26884 (I459920,I244088);
nand I_26885 (I459937,I459841,I459920);
DFFARX1 I_26886 (I459937,I2859,I459742,I459963,);
not I_26887 (I459971,I459963);
not I_26888 (I459988,I244103);
nand I_26889 (I460005,I459988,I244106);
and I_26890 (I460022,I459824,I460005);
nor I_26891 (I460039,I459937,I460022);
DFFARX1 I_26892 (I460039,I2859,I459742,I459710,);
DFFARX1 I_26893 (I460022,I2859,I459742,I459731,);
nor I_26894 (I460084,I244103,I244082);
nor I_26895 (I459722,I459937,I460084);
or I_26896 (I460115,I244103,I244082);
nor I_26897 (I460132,I244094,I244085);
DFFARX1 I_26898 (I460132,I2859,I459742,I460158,);
not I_26899 (I460166,I460158);
nor I_26900 (I459728,I460166,I459971);
nand I_26901 (I460197,I460166,I459816);
not I_26902 (I460214,I244094);
nand I_26903 (I460231,I460214,I459920);
nand I_26904 (I460248,I460166,I460231);
nand I_26905 (I459719,I460248,I460197);
nand I_26906 (I459716,I460231,I460115);
not I_26907 (I460320,I2866);
DFFARX1 I_26908 (I436100,I2859,I460320,I460346,);
and I_26909 (I460354,I460346,I436097);
DFFARX1 I_26910 (I460354,I2859,I460320,I460303,);
DFFARX1 I_26911 (I436103,I2859,I460320,I460394,);
not I_26912 (I460402,I436106);
not I_26913 (I460419,I436100);
nand I_26914 (I460436,I460419,I460402);
nor I_26915 (I460291,I460394,I460436);
DFFARX1 I_26916 (I460436,I2859,I460320,I460476,);
not I_26917 (I460312,I460476);
not I_26918 (I460498,I436115);
nand I_26919 (I460515,I460419,I460498);
DFFARX1 I_26920 (I460515,I2859,I460320,I460541,);
not I_26921 (I460549,I460541);
not I_26922 (I460566,I436112);
nand I_26923 (I460583,I460566,I436118);
and I_26924 (I460600,I460402,I460583);
nor I_26925 (I460617,I460515,I460600);
DFFARX1 I_26926 (I460617,I2859,I460320,I460288,);
DFFARX1 I_26927 (I460600,I2859,I460320,I460309,);
nor I_26928 (I460662,I436112,I436097);
nor I_26929 (I460300,I460515,I460662);
or I_26930 (I460693,I436112,I436097);
nor I_26931 (I460710,I436109,I436103);
DFFARX1 I_26932 (I460710,I2859,I460320,I460736,);
not I_26933 (I460744,I460736);
nor I_26934 (I460306,I460744,I460549);
nand I_26935 (I460775,I460744,I460394);
not I_26936 (I460792,I436109);
nand I_26937 (I460809,I460792,I460498);
nand I_26938 (I460826,I460744,I460809);
nand I_26939 (I460297,I460826,I460775);
nand I_26940 (I460294,I460809,I460693);
not I_26941 (I460898,I2866);
DFFARX1 I_26942 (I162040,I2859,I460898,I460924,);
and I_26943 (I460932,I460924,I162055);
DFFARX1 I_26944 (I460932,I2859,I460898,I460881,);
DFFARX1 I_26945 (I162058,I2859,I460898,I460972,);
not I_26946 (I460980,I162052);
not I_26947 (I460997,I162067);
nand I_26948 (I461014,I460997,I460980);
nor I_26949 (I460869,I460972,I461014);
DFFARX1 I_26950 (I461014,I2859,I460898,I461054,);
not I_26951 (I460890,I461054);
not I_26952 (I461076,I162043);
nand I_26953 (I461093,I460997,I461076);
DFFARX1 I_26954 (I461093,I2859,I460898,I461119,);
not I_26955 (I461127,I461119);
not I_26956 (I461144,I162046);
nand I_26957 (I461161,I461144,I162040);
and I_26958 (I461178,I460980,I461161);
nor I_26959 (I461195,I461093,I461178);
DFFARX1 I_26960 (I461195,I2859,I460898,I460866,);
DFFARX1 I_26961 (I461178,I2859,I460898,I460887,);
nor I_26962 (I461240,I162046,I162049);
nor I_26963 (I460878,I461093,I461240);
or I_26964 (I461271,I162046,I162049);
nor I_26965 (I461288,I162064,I162061);
DFFARX1 I_26966 (I461288,I2859,I460898,I461314,);
not I_26967 (I461322,I461314);
nor I_26968 (I460884,I461322,I461127);
nand I_26969 (I461353,I461322,I460972);
not I_26970 (I461370,I162064);
nand I_26971 (I461387,I461370,I461076);
nand I_26972 (I461404,I461322,I461387);
nand I_26973 (I460875,I461404,I461353);
nand I_26974 (I460872,I461387,I461271);
not I_26975 (I461476,I2866);
DFFARX1 I_26976 (I314613,I2859,I461476,I461502,);
and I_26977 (I461510,I461502,I314601);
DFFARX1 I_26978 (I461510,I2859,I461476,I461459,);
DFFARX1 I_26979 (I314604,I2859,I461476,I461550,);
not I_26980 (I461558,I314598);
not I_26981 (I461575,I314622);
nand I_26982 (I461592,I461575,I461558);
nor I_26983 (I461447,I461550,I461592);
DFFARX1 I_26984 (I461592,I2859,I461476,I461632,);
not I_26985 (I461468,I461632);
not I_26986 (I461654,I314610);
nand I_26987 (I461671,I461575,I461654);
DFFARX1 I_26988 (I461671,I2859,I461476,I461697,);
not I_26989 (I461705,I461697);
not I_26990 (I461722,I314619);
nand I_26991 (I461739,I461722,I314616);
and I_26992 (I461756,I461558,I461739);
nor I_26993 (I461773,I461671,I461756);
DFFARX1 I_26994 (I461773,I2859,I461476,I461444,);
DFFARX1 I_26995 (I461756,I2859,I461476,I461465,);
nor I_26996 (I461818,I314619,I314607);
nor I_26997 (I461456,I461671,I461818);
or I_26998 (I461849,I314619,I314607);
nor I_26999 (I461866,I314598,I314601);
DFFARX1 I_27000 (I461866,I2859,I461476,I461892,);
not I_27001 (I461900,I461892);
nor I_27002 (I461462,I461900,I461705);
nand I_27003 (I461931,I461900,I461550);
not I_27004 (I461948,I314598);
nand I_27005 (I461965,I461948,I461654);
nand I_27006 (I461982,I461900,I461965);
nand I_27007 (I461453,I461982,I461931);
nand I_27008 (I461450,I461965,I461849);
not I_27009 (I462054,I2866);
DFFARX1 I_27010 (I196856,I2859,I462054,I462080,);
and I_27011 (I462088,I462080,I196871);
DFFARX1 I_27012 (I462088,I2859,I462054,I462037,);
DFFARX1 I_27013 (I196874,I2859,I462054,I462128,);
not I_27014 (I462136,I196868);
not I_27015 (I462153,I196883);
nand I_27016 (I462170,I462153,I462136);
nor I_27017 (I462025,I462128,I462170);
DFFARX1 I_27018 (I462170,I2859,I462054,I462210,);
not I_27019 (I462046,I462210);
not I_27020 (I462232,I196859);
nand I_27021 (I462249,I462153,I462232);
DFFARX1 I_27022 (I462249,I2859,I462054,I462275,);
not I_27023 (I462283,I462275);
not I_27024 (I462300,I196862);
nand I_27025 (I462317,I462300,I196856);
and I_27026 (I462334,I462136,I462317);
nor I_27027 (I462351,I462249,I462334);
DFFARX1 I_27028 (I462351,I2859,I462054,I462022,);
DFFARX1 I_27029 (I462334,I2859,I462054,I462043,);
nor I_27030 (I462396,I196862,I196865);
nor I_27031 (I462034,I462249,I462396);
or I_27032 (I462427,I196862,I196865);
nor I_27033 (I462444,I196880,I196877);
DFFARX1 I_27034 (I462444,I2859,I462054,I462470,);
not I_27035 (I462478,I462470);
nor I_27036 (I462040,I462478,I462283);
nand I_27037 (I462509,I462478,I462128);
not I_27038 (I462526,I196880);
nand I_27039 (I462543,I462526,I462232);
nand I_27040 (I462560,I462478,I462543);
nand I_27041 (I462031,I462560,I462509);
nand I_27042 (I462028,I462543,I462427);
not I_27043 (I462632,I2866);
DFFARX1 I_27044 (I271841,I2859,I462632,I462658,);
and I_27045 (I462666,I462658,I271829);
DFFARX1 I_27046 (I462666,I2859,I462632,I462615,);
DFFARX1 I_27047 (I271832,I2859,I462632,I462706,);
not I_27048 (I462714,I271826);
not I_27049 (I462731,I271850);
nand I_27050 (I462748,I462731,I462714);
nor I_27051 (I462603,I462706,I462748);
DFFARX1 I_27052 (I462748,I2859,I462632,I462788,);
not I_27053 (I462624,I462788);
not I_27054 (I462810,I271838);
nand I_27055 (I462827,I462731,I462810);
DFFARX1 I_27056 (I462827,I2859,I462632,I462853,);
not I_27057 (I462861,I462853);
not I_27058 (I462878,I271847);
nand I_27059 (I462895,I462878,I271844);
and I_27060 (I462912,I462714,I462895);
nor I_27061 (I462929,I462827,I462912);
DFFARX1 I_27062 (I462929,I2859,I462632,I462600,);
DFFARX1 I_27063 (I462912,I2859,I462632,I462621,);
nor I_27064 (I462974,I271847,I271835);
nor I_27065 (I462612,I462827,I462974);
or I_27066 (I463005,I271847,I271835);
nor I_27067 (I463022,I271826,I271829);
DFFARX1 I_27068 (I463022,I2859,I462632,I463048,);
not I_27069 (I463056,I463048);
nor I_27070 (I462618,I463056,I462861);
nand I_27071 (I463087,I463056,I462706);
not I_27072 (I463104,I271826);
nand I_27073 (I463121,I463104,I462810);
nand I_27074 (I463138,I463056,I463121);
nand I_27075 (I462609,I463138,I463087);
nand I_27076 (I462606,I463121,I463005);
not I_27077 (I463210,I2866);
DFFARX1 I_27078 (I340730,I2859,I463210,I463236,);
and I_27079 (I463244,I463236,I340736);
DFFARX1 I_27080 (I463244,I2859,I463210,I463193,);
DFFARX1 I_27081 (I340742,I2859,I463210,I463284,);
not I_27082 (I463292,I340727);
not I_27083 (I463309,I340727);
nand I_27084 (I463326,I463309,I463292);
nor I_27085 (I463181,I463284,I463326);
DFFARX1 I_27086 (I463326,I2859,I463210,I463366,);
not I_27087 (I463202,I463366);
not I_27088 (I463388,I340745);
nand I_27089 (I463405,I463309,I463388);
DFFARX1 I_27090 (I463405,I2859,I463210,I463431,);
not I_27091 (I463439,I463431);
not I_27092 (I463456,I340739);
nand I_27093 (I463473,I463456,I340730);
and I_27094 (I463490,I463292,I463473);
nor I_27095 (I463507,I463405,I463490);
DFFARX1 I_27096 (I463507,I2859,I463210,I463178,);
DFFARX1 I_27097 (I463490,I2859,I463210,I463199,);
nor I_27098 (I463552,I340739,I340748);
nor I_27099 (I463190,I463405,I463552);
or I_27100 (I463583,I340739,I340748);
nor I_27101 (I463600,I340733,I340733);
DFFARX1 I_27102 (I463600,I2859,I463210,I463626,);
not I_27103 (I463634,I463626);
nor I_27104 (I463196,I463634,I463439);
nand I_27105 (I463665,I463634,I463284);
not I_27106 (I463682,I340733);
nand I_27107 (I463699,I463682,I463388);
nand I_27108 (I463716,I463634,I463699);
nand I_27109 (I463187,I463716,I463665);
nand I_27110 (I463184,I463699,I463583);
not I_27111 (I463788,I2866);
DFFARX1 I_27112 (I572532,I2859,I463788,I463814,);
and I_27113 (I463822,I463814,I572514);
DFFARX1 I_27114 (I463822,I2859,I463788,I463771,);
DFFARX1 I_27115 (I572505,I2859,I463788,I463862,);
not I_27116 (I463870,I572520);
not I_27117 (I463887,I572508);
nand I_27118 (I463904,I463887,I463870);
nor I_27119 (I463759,I463862,I463904);
DFFARX1 I_27120 (I463904,I2859,I463788,I463944,);
not I_27121 (I463780,I463944);
not I_27122 (I463966,I572517);
nand I_27123 (I463983,I463887,I463966);
DFFARX1 I_27124 (I463983,I2859,I463788,I464009,);
not I_27125 (I464017,I464009);
not I_27126 (I464034,I572526);
nand I_27127 (I464051,I464034,I572505);
and I_27128 (I464068,I463870,I464051);
nor I_27129 (I464085,I463983,I464068);
DFFARX1 I_27130 (I464085,I2859,I463788,I463756,);
DFFARX1 I_27131 (I464068,I2859,I463788,I463777,);
nor I_27132 (I464130,I572526,I572529);
nor I_27133 (I463768,I463983,I464130);
or I_27134 (I464161,I572526,I572529);
nor I_27135 (I464178,I572523,I572511);
DFFARX1 I_27136 (I464178,I2859,I463788,I464204,);
not I_27137 (I464212,I464204);
nor I_27138 (I463774,I464212,I464017);
nand I_27139 (I464243,I464212,I463862);
not I_27140 (I464260,I572523);
nand I_27141 (I464277,I464260,I463966);
nand I_27142 (I464294,I464212,I464277);
nand I_27143 (I463765,I464294,I464243);
nand I_27144 (I463762,I464277,I464161);
not I_27145 (I464366,I2866);
DFFARX1 I_27146 (I280511,I2859,I464366,I464392,);
and I_27147 (I464400,I464392,I280499);
DFFARX1 I_27148 (I464400,I2859,I464366,I464349,);
DFFARX1 I_27149 (I280502,I2859,I464366,I464440,);
not I_27150 (I464448,I280496);
not I_27151 (I464465,I280520);
nand I_27152 (I464482,I464465,I464448);
nor I_27153 (I464337,I464440,I464482);
DFFARX1 I_27154 (I464482,I2859,I464366,I464522,);
not I_27155 (I464358,I464522);
not I_27156 (I464544,I280508);
nand I_27157 (I464561,I464465,I464544);
DFFARX1 I_27158 (I464561,I2859,I464366,I464587,);
not I_27159 (I464595,I464587);
not I_27160 (I464612,I280517);
nand I_27161 (I464629,I464612,I280514);
and I_27162 (I464646,I464448,I464629);
nor I_27163 (I464663,I464561,I464646);
DFFARX1 I_27164 (I464663,I2859,I464366,I464334,);
DFFARX1 I_27165 (I464646,I2859,I464366,I464355,);
nor I_27166 (I464708,I280517,I280505);
nor I_27167 (I464346,I464561,I464708);
or I_27168 (I464739,I280517,I280505);
nor I_27169 (I464756,I280496,I280499);
DFFARX1 I_27170 (I464756,I2859,I464366,I464782,);
not I_27171 (I464790,I464782);
nor I_27172 (I464352,I464790,I464595);
nand I_27173 (I464821,I464790,I464440);
not I_27174 (I464838,I280496);
nand I_27175 (I464855,I464838,I464544);
nand I_27176 (I464872,I464790,I464855);
nand I_27177 (I464343,I464872,I464821);
nand I_27178 (I464340,I464855,I464739);
not I_27179 (I464944,I2866);
DFFARX1 I_27180 (I117748,I2859,I464944,I464970,);
and I_27181 (I464978,I464970,I117733);
DFFARX1 I_27182 (I464978,I2859,I464944,I464927,);
DFFARX1 I_27183 (I117739,I2859,I464944,I465018,);
not I_27184 (I465026,I117721);
not I_27185 (I465043,I117742);
nand I_27186 (I465060,I465043,I465026);
nor I_27187 (I464915,I465018,I465060);
DFFARX1 I_27188 (I465060,I2859,I464944,I465100,);
not I_27189 (I464936,I465100);
not I_27190 (I465122,I117745);
nand I_27191 (I465139,I465043,I465122);
DFFARX1 I_27192 (I465139,I2859,I464944,I465165,);
not I_27193 (I465173,I465165);
not I_27194 (I465190,I117736);
nand I_27195 (I465207,I465190,I117724);
and I_27196 (I465224,I465026,I465207);
nor I_27197 (I465241,I465139,I465224);
DFFARX1 I_27198 (I465241,I2859,I464944,I464912,);
DFFARX1 I_27199 (I465224,I2859,I464944,I464933,);
nor I_27200 (I465286,I117736,I117730);
nor I_27201 (I464924,I465139,I465286);
or I_27202 (I465317,I117736,I117730);
nor I_27203 (I465334,I117727,I117721);
DFFARX1 I_27204 (I465334,I2859,I464944,I465360,);
not I_27205 (I465368,I465360);
nor I_27206 (I464930,I465368,I465173);
nand I_27207 (I465399,I465368,I465018);
not I_27208 (I465416,I117727);
nand I_27209 (I465433,I465416,I465122);
nand I_27210 (I465450,I465368,I465433);
nand I_27211 (I464921,I465450,I465399);
nand I_27212 (I464918,I465433,I465317);
not I_27213 (I465522,I2866);
DFFARX1 I_27214 (I201908,I2859,I465522,I465548,);
and I_27215 (I465556,I465548,I201923);
DFFARX1 I_27216 (I465556,I2859,I465522,I465505,);
DFFARX1 I_27217 (I201914,I2859,I465522,I465596,);
not I_27218 (I465604,I201908);
not I_27219 (I465621,I201926);
nand I_27220 (I465638,I465621,I465604);
nor I_27221 (I465493,I465596,I465638);
DFFARX1 I_27222 (I465638,I2859,I465522,I465678,);
not I_27223 (I465514,I465678);
not I_27224 (I465700,I201917);
nand I_27225 (I465717,I465621,I465700);
DFFARX1 I_27226 (I465717,I2859,I465522,I465743,);
not I_27227 (I465751,I465743);
not I_27228 (I465768,I201929);
nand I_27229 (I465785,I465768,I201905);
and I_27230 (I465802,I465604,I465785);
nor I_27231 (I465819,I465717,I465802);
DFFARX1 I_27232 (I465819,I2859,I465522,I465490,);
DFFARX1 I_27233 (I465802,I2859,I465522,I465511,);
nor I_27234 (I465864,I201929,I201905);
nor I_27235 (I465502,I465717,I465864);
or I_27236 (I465895,I201929,I201905);
nor I_27237 (I465912,I201911,I201920);
DFFARX1 I_27238 (I465912,I2859,I465522,I465938,);
not I_27239 (I465946,I465938);
nor I_27240 (I465508,I465946,I465751);
nand I_27241 (I465977,I465946,I465596);
not I_27242 (I465994,I201911);
nand I_27243 (I466011,I465994,I465700);
nand I_27244 (I466028,I465946,I466011);
nand I_27245 (I465499,I466028,I465977);
nand I_27246 (I465496,I466011,I465895);
not I_27247 (I466100,I2866);
DFFARX1 I_27248 (I299585,I2859,I466100,I466126,);
and I_27249 (I466134,I466126,I299573);
DFFARX1 I_27250 (I466134,I2859,I466100,I466083,);
DFFARX1 I_27251 (I299576,I2859,I466100,I466174,);
not I_27252 (I466182,I299570);
not I_27253 (I466199,I299594);
nand I_27254 (I466216,I466199,I466182);
nor I_27255 (I466071,I466174,I466216);
DFFARX1 I_27256 (I466216,I2859,I466100,I466256,);
not I_27257 (I466092,I466256);
not I_27258 (I466278,I299582);
nand I_27259 (I466295,I466199,I466278);
DFFARX1 I_27260 (I466295,I2859,I466100,I466321,);
not I_27261 (I466329,I466321);
not I_27262 (I466346,I299591);
nand I_27263 (I466363,I466346,I299588);
and I_27264 (I466380,I466182,I466363);
nor I_27265 (I466397,I466295,I466380);
DFFARX1 I_27266 (I466397,I2859,I466100,I466068,);
DFFARX1 I_27267 (I466380,I2859,I466100,I466089,);
nor I_27268 (I466442,I299591,I299579);
nor I_27269 (I466080,I466295,I466442);
or I_27270 (I466473,I299591,I299579);
nor I_27271 (I466490,I299570,I299573);
DFFARX1 I_27272 (I466490,I2859,I466100,I466516,);
not I_27273 (I466524,I466516);
nor I_27274 (I466086,I466524,I466329);
nand I_27275 (I466555,I466524,I466174);
not I_27276 (I466572,I299570);
nand I_27277 (I466589,I466572,I466278);
nand I_27278 (I466606,I466524,I466589);
nand I_27279 (I466077,I466606,I466555);
nand I_27280 (I466074,I466589,I466473);
not I_27281 (I466678,I2866);
DFFARX1 I_27282 (I189240,I2859,I466678,I466704,);
and I_27283 (I466712,I466704,I189255);
DFFARX1 I_27284 (I466712,I2859,I466678,I466661,);
DFFARX1 I_27285 (I189258,I2859,I466678,I466752,);
not I_27286 (I466760,I189252);
not I_27287 (I466777,I189267);
nand I_27288 (I466794,I466777,I466760);
nor I_27289 (I466649,I466752,I466794);
DFFARX1 I_27290 (I466794,I2859,I466678,I466834,);
not I_27291 (I466670,I466834);
not I_27292 (I466856,I189243);
nand I_27293 (I466873,I466777,I466856);
DFFARX1 I_27294 (I466873,I2859,I466678,I466899,);
not I_27295 (I466907,I466899);
not I_27296 (I466924,I189246);
nand I_27297 (I466941,I466924,I189240);
and I_27298 (I466958,I466760,I466941);
nor I_27299 (I466975,I466873,I466958);
DFFARX1 I_27300 (I466975,I2859,I466678,I466646,);
DFFARX1 I_27301 (I466958,I2859,I466678,I466667,);
nor I_27302 (I467020,I189246,I189249);
nor I_27303 (I466658,I466873,I467020);
or I_27304 (I467051,I189246,I189249);
nor I_27305 (I467068,I189264,I189261);
DFFARX1 I_27306 (I467068,I2859,I466678,I467094,);
not I_27307 (I467102,I467094);
nor I_27308 (I466664,I467102,I466907);
nand I_27309 (I467133,I467102,I466752);
not I_27310 (I467150,I189264);
nand I_27311 (I467167,I467150,I466856);
nand I_27312 (I467184,I467102,I467167);
nand I_27313 (I466655,I467184,I467133);
nand I_27314 (I466652,I467167,I467051);
not I_27315 (I467256,I2866);
DFFARX1 I_27316 (I394759,I2859,I467256,I467282,);
and I_27317 (I467290,I467282,I394753);
DFFARX1 I_27318 (I467290,I2859,I467256,I467239,);
DFFARX1 I_27319 (I394771,I2859,I467256,I467330,);
not I_27320 (I467338,I394762);
not I_27321 (I467355,I394774);
nand I_27322 (I467372,I467355,I467338);
nor I_27323 (I467227,I467330,I467372);
DFFARX1 I_27324 (I467372,I2859,I467256,I467412,);
not I_27325 (I467248,I467412);
not I_27326 (I467434,I394780);
nand I_27327 (I467451,I467355,I467434);
DFFARX1 I_27328 (I467451,I2859,I467256,I467477,);
not I_27329 (I467485,I467477);
not I_27330 (I467502,I394756);
nand I_27331 (I467519,I467502,I394777);
and I_27332 (I467536,I467338,I467519);
nor I_27333 (I467553,I467451,I467536);
DFFARX1 I_27334 (I467553,I2859,I467256,I467224,);
DFFARX1 I_27335 (I467536,I2859,I467256,I467245,);
nor I_27336 (I467598,I394756,I394768);
nor I_27337 (I467236,I467451,I467598);
or I_27338 (I467629,I394756,I394768);
nor I_27339 (I467646,I394753,I394765);
DFFARX1 I_27340 (I467646,I2859,I467256,I467672,);
not I_27341 (I467680,I467672);
nor I_27342 (I467242,I467680,I467485);
nand I_27343 (I467711,I467680,I467330);
not I_27344 (I467728,I394753);
nand I_27345 (I467745,I467728,I467434);
nand I_27346 (I467762,I467680,I467745);
nand I_27347 (I467233,I467762,I467711);
nand I_27348 (I467230,I467745,I467629);
not I_27349 (I467834,I2866);
DFFARX1 I_27350 (I275887,I2859,I467834,I467860,);
and I_27351 (I467868,I467860,I275875);
DFFARX1 I_27352 (I467868,I2859,I467834,I467817,);
DFFARX1 I_27353 (I275878,I2859,I467834,I467908,);
not I_27354 (I467916,I275872);
not I_27355 (I467933,I275896);
nand I_27356 (I467950,I467933,I467916);
nor I_27357 (I467805,I467908,I467950);
DFFARX1 I_27358 (I467950,I2859,I467834,I467990,);
not I_27359 (I467826,I467990);
not I_27360 (I468012,I275884);
nand I_27361 (I468029,I467933,I468012);
DFFARX1 I_27362 (I468029,I2859,I467834,I468055,);
not I_27363 (I468063,I468055);
not I_27364 (I468080,I275893);
nand I_27365 (I468097,I468080,I275890);
and I_27366 (I468114,I467916,I468097);
nor I_27367 (I468131,I468029,I468114);
DFFARX1 I_27368 (I468131,I2859,I467834,I467802,);
DFFARX1 I_27369 (I468114,I2859,I467834,I467823,);
nor I_27370 (I468176,I275893,I275881);
nor I_27371 (I467814,I468029,I468176);
or I_27372 (I468207,I275893,I275881);
nor I_27373 (I468224,I275872,I275875);
DFFARX1 I_27374 (I468224,I2859,I467834,I468250,);
not I_27375 (I468258,I468250);
nor I_27376 (I467820,I468258,I468063);
nand I_27377 (I468289,I468258,I467908);
not I_27378 (I468306,I275872);
nand I_27379 (I468323,I468306,I468012);
nand I_27380 (I468340,I468258,I468323);
nand I_27381 (I467811,I468340,I468289);
nand I_27382 (I467808,I468323,I468207);
not I_27383 (I468412,I2866);
DFFARX1 I_27384 (I94737,I2859,I468412,I468438,);
and I_27385 (I468446,I468438,I94740);
DFFARX1 I_27386 (I468446,I2859,I468412,I468395,);
DFFARX1 I_27387 (I94740,I2859,I468412,I468486,);
not I_27388 (I468494,I94755);
not I_27389 (I468511,I94761);
nand I_27390 (I468528,I468511,I468494);
nor I_27391 (I468383,I468486,I468528);
DFFARX1 I_27392 (I468528,I2859,I468412,I468568,);
not I_27393 (I468404,I468568);
not I_27394 (I468590,I94749);
nand I_27395 (I468607,I468511,I468590);
DFFARX1 I_27396 (I468607,I2859,I468412,I468633,);
not I_27397 (I468641,I468633);
not I_27398 (I468658,I94746);
nand I_27399 (I468675,I468658,I94743);
and I_27400 (I468692,I468494,I468675);
nor I_27401 (I468709,I468607,I468692);
DFFARX1 I_27402 (I468709,I2859,I468412,I468380,);
DFFARX1 I_27403 (I468692,I2859,I468412,I468401,);
nor I_27404 (I468754,I94746,I94737);
nor I_27405 (I468392,I468607,I468754);
or I_27406 (I468785,I94746,I94737);
nor I_27407 (I468802,I94752,I94758);
DFFARX1 I_27408 (I468802,I2859,I468412,I468828,);
not I_27409 (I468836,I468828);
nor I_27410 (I468398,I468836,I468641);
nand I_27411 (I468867,I468836,I468486);
not I_27412 (I468884,I94752);
nand I_27413 (I468901,I468884,I468590);
nand I_27414 (I468918,I468836,I468901);
nand I_27415 (I468389,I468918,I468867);
nand I_27416 (I468386,I468901,I468785);
not I_27417 (I468990,I2866);
DFFARX1 I_27418 (I54277,I2859,I468990,I469016,);
and I_27419 (I469024,I469016,I54280);
DFFARX1 I_27420 (I469024,I2859,I468990,I468973,);
DFFARX1 I_27421 (I54280,I2859,I468990,I469064,);
not I_27422 (I469072,I54295);
not I_27423 (I469089,I54301);
nand I_27424 (I469106,I469089,I469072);
nor I_27425 (I468961,I469064,I469106);
DFFARX1 I_27426 (I469106,I2859,I468990,I469146,);
not I_27427 (I468982,I469146);
not I_27428 (I469168,I54289);
nand I_27429 (I469185,I469089,I469168);
DFFARX1 I_27430 (I469185,I2859,I468990,I469211,);
not I_27431 (I469219,I469211);
not I_27432 (I469236,I54286);
nand I_27433 (I469253,I469236,I54283);
and I_27434 (I469270,I469072,I469253);
nor I_27435 (I469287,I469185,I469270);
DFFARX1 I_27436 (I469287,I2859,I468990,I468958,);
DFFARX1 I_27437 (I469270,I2859,I468990,I468979,);
nor I_27438 (I469332,I54286,I54277);
nor I_27439 (I468970,I469185,I469332);
or I_27440 (I469363,I54286,I54277);
nor I_27441 (I469380,I54292,I54298);
DFFARX1 I_27442 (I469380,I2859,I468990,I469406,);
not I_27443 (I469414,I469406);
nor I_27444 (I468976,I469414,I469219);
nand I_27445 (I469445,I469414,I469064);
not I_27446 (I469462,I54292);
nand I_27447 (I469479,I469462,I469168);
nand I_27448 (I469496,I469414,I469479);
nand I_27449 (I468967,I469496,I469445);
nand I_27450 (I468964,I469479,I469363);
not I_27451 (I469568,I2866);
DFFARX1 I_27452 (I125653,I2859,I469568,I469594,);
and I_27453 (I469602,I469594,I125638);
DFFARX1 I_27454 (I469602,I2859,I469568,I469551,);
DFFARX1 I_27455 (I125644,I2859,I469568,I469642,);
not I_27456 (I469650,I125626);
not I_27457 (I469667,I125647);
nand I_27458 (I469684,I469667,I469650);
nor I_27459 (I469539,I469642,I469684);
DFFARX1 I_27460 (I469684,I2859,I469568,I469724,);
not I_27461 (I469560,I469724);
not I_27462 (I469746,I125650);
nand I_27463 (I469763,I469667,I469746);
DFFARX1 I_27464 (I469763,I2859,I469568,I469789,);
not I_27465 (I469797,I469789);
not I_27466 (I469814,I125641);
nand I_27467 (I469831,I469814,I125629);
and I_27468 (I469848,I469650,I469831);
nor I_27469 (I469865,I469763,I469848);
DFFARX1 I_27470 (I469865,I2859,I469568,I469536,);
DFFARX1 I_27471 (I469848,I2859,I469568,I469557,);
nor I_27472 (I469910,I125641,I125635);
nor I_27473 (I469548,I469763,I469910);
or I_27474 (I469941,I125641,I125635);
nor I_27475 (I469958,I125632,I125626);
DFFARX1 I_27476 (I469958,I2859,I469568,I469984,);
not I_27477 (I469992,I469984);
nor I_27478 (I469554,I469992,I469797);
nand I_27479 (I470023,I469992,I469642);
not I_27480 (I470040,I125632);
nand I_27481 (I470057,I470040,I469746);
nand I_27482 (I470074,I469992,I470057);
nand I_27483 (I469545,I470074,I470023);
nand I_27484 (I469542,I470057,I469941);
not I_27485 (I470146,I2866);
DFFARX1 I_27486 (I26421,I2859,I470146,I470172,);
and I_27487 (I470180,I470172,I26397);
DFFARX1 I_27488 (I470180,I2859,I470146,I470129,);
DFFARX1 I_27489 (I26415,I2859,I470146,I470220,);
not I_27490 (I470228,I26403);
not I_27491 (I470245,I26400);
nand I_27492 (I470262,I470245,I470228);
nor I_27493 (I470117,I470220,I470262);
DFFARX1 I_27494 (I470262,I2859,I470146,I470302,);
not I_27495 (I470138,I470302);
not I_27496 (I470324,I26409);
nand I_27497 (I470341,I470245,I470324);
DFFARX1 I_27498 (I470341,I2859,I470146,I470367,);
not I_27499 (I470375,I470367);
not I_27500 (I470392,I26400);
nand I_27501 (I470409,I470392,I26418);
and I_27502 (I470426,I470228,I470409);
nor I_27503 (I470443,I470341,I470426);
DFFARX1 I_27504 (I470443,I2859,I470146,I470114,);
DFFARX1 I_27505 (I470426,I2859,I470146,I470135,);
nor I_27506 (I470488,I26400,I26412);
nor I_27507 (I470126,I470341,I470488);
or I_27508 (I470519,I26400,I26412);
nor I_27509 (I470536,I26406,I26397);
DFFARX1 I_27510 (I470536,I2859,I470146,I470562,);
not I_27511 (I470570,I470562);
nor I_27512 (I470132,I470570,I470375);
nand I_27513 (I470601,I470570,I470220);
not I_27514 (I470618,I26406);
nand I_27515 (I470635,I470618,I470324);
nand I_27516 (I470652,I470570,I470635);
nand I_27517 (I470123,I470652,I470601);
nand I_27518 (I470120,I470635,I470519);
not I_27519 (I470724,I2866);
DFFARX1 I_27520 (I534452,I2859,I470724,I470750,);
and I_27521 (I470758,I470750,I534434);
DFFARX1 I_27522 (I470758,I2859,I470724,I470707,);
DFFARX1 I_27523 (I534425,I2859,I470724,I470798,);
not I_27524 (I470806,I534440);
not I_27525 (I470823,I534428);
nand I_27526 (I470840,I470823,I470806);
nor I_27527 (I470695,I470798,I470840);
DFFARX1 I_27528 (I470840,I2859,I470724,I470880,);
not I_27529 (I470716,I470880);
not I_27530 (I470902,I534437);
nand I_27531 (I470919,I470823,I470902);
DFFARX1 I_27532 (I470919,I2859,I470724,I470945,);
not I_27533 (I470953,I470945);
not I_27534 (I470970,I534446);
nand I_27535 (I470987,I470970,I534425);
and I_27536 (I471004,I470806,I470987);
nor I_27537 (I471021,I470919,I471004);
DFFARX1 I_27538 (I471021,I2859,I470724,I470692,);
DFFARX1 I_27539 (I471004,I2859,I470724,I470713,);
nor I_27540 (I471066,I534446,I534449);
nor I_27541 (I470704,I470919,I471066);
or I_27542 (I471097,I534446,I534449);
nor I_27543 (I471114,I534443,I534431);
DFFARX1 I_27544 (I471114,I2859,I470724,I471140,);
not I_27545 (I471148,I471140);
nor I_27546 (I470710,I471148,I470953);
nand I_27547 (I471179,I471148,I470798);
not I_27548 (I471196,I534443);
nand I_27549 (I471213,I471196,I470902);
nand I_27550 (I471230,I471148,I471213);
nand I_27551 (I470701,I471230,I471179);
nand I_27552 (I470698,I471213,I471097);
not I_27553 (I471302,I2866);
DFFARX1 I_27554 (I538617,I2859,I471302,I471328,);
and I_27555 (I471336,I471328,I538599);
DFFARX1 I_27556 (I471336,I2859,I471302,I471285,);
DFFARX1 I_27557 (I538590,I2859,I471302,I471376,);
not I_27558 (I471384,I538605);
not I_27559 (I471401,I538593);
nand I_27560 (I471418,I471401,I471384);
nor I_27561 (I471273,I471376,I471418);
DFFARX1 I_27562 (I471418,I2859,I471302,I471458,);
not I_27563 (I471294,I471458);
not I_27564 (I471480,I538602);
nand I_27565 (I471497,I471401,I471480);
DFFARX1 I_27566 (I471497,I2859,I471302,I471523,);
not I_27567 (I471531,I471523);
not I_27568 (I471548,I538611);
nand I_27569 (I471565,I471548,I538590);
and I_27570 (I471582,I471384,I471565);
nor I_27571 (I471599,I471497,I471582);
DFFARX1 I_27572 (I471599,I2859,I471302,I471270,);
DFFARX1 I_27573 (I471582,I2859,I471302,I471291,);
nor I_27574 (I471644,I538611,I538614);
nor I_27575 (I471282,I471497,I471644);
or I_27576 (I471675,I538611,I538614);
nor I_27577 (I471692,I538608,I538596);
DFFARX1 I_27578 (I471692,I2859,I471302,I471718,);
not I_27579 (I471726,I471718);
nor I_27580 (I471288,I471726,I471531);
nand I_27581 (I471757,I471726,I471376);
not I_27582 (I471774,I538608);
nand I_27583 (I471791,I471774,I471480);
nand I_27584 (I471808,I471726,I471791);
nand I_27585 (I471279,I471808,I471757);
nand I_27586 (I471276,I471791,I471675);
not I_27587 (I471880,I2866);
DFFARX1 I_27588 (I81052,I2859,I471880,I471906,);
and I_27589 (I471914,I471906,I81055);
DFFARX1 I_27590 (I471914,I2859,I471880,I471863,);
DFFARX1 I_27591 (I81055,I2859,I471880,I471954,);
not I_27592 (I471962,I81070);
not I_27593 (I471979,I81076);
nand I_27594 (I471996,I471979,I471962);
nor I_27595 (I471851,I471954,I471996);
DFFARX1 I_27596 (I471996,I2859,I471880,I472036,);
not I_27597 (I471872,I472036);
not I_27598 (I472058,I81064);
nand I_27599 (I472075,I471979,I472058);
DFFARX1 I_27600 (I472075,I2859,I471880,I472101,);
not I_27601 (I472109,I472101);
not I_27602 (I472126,I81061);
nand I_27603 (I472143,I472126,I81058);
and I_27604 (I472160,I471962,I472143);
nor I_27605 (I472177,I472075,I472160);
DFFARX1 I_27606 (I472177,I2859,I471880,I471848,);
DFFARX1 I_27607 (I472160,I2859,I471880,I471869,);
nor I_27608 (I472222,I81061,I81052);
nor I_27609 (I471860,I472075,I472222);
or I_27610 (I472253,I81061,I81052);
nor I_27611 (I472270,I81067,I81073);
DFFARX1 I_27612 (I472270,I2859,I471880,I472296,);
not I_27613 (I472304,I472296);
nor I_27614 (I471866,I472304,I472109);
nand I_27615 (I472335,I472304,I471954);
not I_27616 (I472352,I81067);
nand I_27617 (I472369,I472352,I472058);
nand I_27618 (I472386,I472304,I472369);
nand I_27619 (I471857,I472386,I472335);
nand I_27620 (I471854,I472369,I472253);
not I_27621 (I472458,I2866);
DFFARX1 I_27622 (I414139,I2859,I472458,I472484,);
and I_27623 (I472492,I472484,I414133);
DFFARX1 I_27624 (I472492,I2859,I472458,I472441,);
DFFARX1 I_27625 (I414151,I2859,I472458,I472532,);
not I_27626 (I472540,I414142);
not I_27627 (I472557,I414154);
nand I_27628 (I472574,I472557,I472540);
nor I_27629 (I472429,I472532,I472574);
DFFARX1 I_27630 (I472574,I2859,I472458,I472614,);
not I_27631 (I472450,I472614);
not I_27632 (I472636,I414160);
nand I_27633 (I472653,I472557,I472636);
DFFARX1 I_27634 (I472653,I2859,I472458,I472679,);
not I_27635 (I472687,I472679);
not I_27636 (I472704,I414136);
nand I_27637 (I472721,I472704,I414157);
and I_27638 (I472738,I472540,I472721);
nor I_27639 (I472755,I472653,I472738);
DFFARX1 I_27640 (I472755,I2859,I472458,I472426,);
DFFARX1 I_27641 (I472738,I2859,I472458,I472447,);
nor I_27642 (I472800,I414136,I414148);
nor I_27643 (I472438,I472653,I472800);
or I_27644 (I472831,I414136,I414148);
nor I_27645 (I472848,I414133,I414145);
DFFARX1 I_27646 (I472848,I2859,I472458,I472874,);
not I_27647 (I472882,I472874);
nor I_27648 (I472444,I472882,I472687);
nand I_27649 (I472913,I472882,I472532);
not I_27650 (I472930,I414133);
nand I_27651 (I472947,I472930,I472636);
nand I_27652 (I472964,I472882,I472947);
nand I_27653 (I472435,I472964,I472913);
nand I_27654 (I472432,I472947,I472831);
not I_27655 (I473036,I2866);
DFFARX1 I_27656 (I225023,I2859,I473036,I473062,);
and I_27657 (I473070,I473062,I225011);
DFFARX1 I_27658 (I473070,I2859,I473036,I473019,);
DFFARX1 I_27659 (I225026,I2859,I473036,I473110,);
not I_27660 (I473118,I225017);
not I_27661 (I473135,I225008);
nand I_27662 (I473152,I473135,I473118);
nor I_27663 (I473007,I473110,I473152);
DFFARX1 I_27664 (I473152,I2859,I473036,I473192,);
not I_27665 (I473028,I473192);
not I_27666 (I473214,I225014);
nand I_27667 (I473231,I473135,I473214);
DFFARX1 I_27668 (I473231,I2859,I473036,I473257,);
not I_27669 (I473265,I473257);
not I_27670 (I473282,I225029);
nand I_27671 (I473299,I473282,I225032);
and I_27672 (I473316,I473118,I473299);
nor I_27673 (I473333,I473231,I473316);
DFFARX1 I_27674 (I473333,I2859,I473036,I473004,);
DFFARX1 I_27675 (I473316,I2859,I473036,I473025,);
nor I_27676 (I473378,I225029,I225008);
nor I_27677 (I473016,I473231,I473378);
or I_27678 (I473409,I225029,I225008);
nor I_27679 (I473426,I225020,I225011);
DFFARX1 I_27680 (I473426,I2859,I473036,I473452,);
not I_27681 (I473460,I473452);
nor I_27682 (I473022,I473460,I473265);
nand I_27683 (I473491,I473460,I473110);
not I_27684 (I473508,I225020);
nand I_27685 (I473525,I473508,I473214);
nand I_27686 (I473542,I473460,I473525);
nand I_27687 (I473013,I473542,I473491);
nand I_27688 (I473010,I473525,I473409);
not I_27689 (I473614,I2866);
DFFARX1 I_27690 (I207263,I2859,I473614,I473640,);
and I_27691 (I473648,I473640,I207278);
DFFARX1 I_27692 (I473648,I2859,I473614,I473597,);
DFFARX1 I_27693 (I207269,I2859,I473614,I473688,);
not I_27694 (I473696,I207263);
not I_27695 (I473713,I207281);
nand I_27696 (I473730,I473713,I473696);
nor I_27697 (I473585,I473688,I473730);
DFFARX1 I_27698 (I473730,I2859,I473614,I473770,);
not I_27699 (I473606,I473770);
not I_27700 (I473792,I207272);
nand I_27701 (I473809,I473713,I473792);
DFFARX1 I_27702 (I473809,I2859,I473614,I473835,);
not I_27703 (I473843,I473835);
not I_27704 (I473860,I207284);
nand I_27705 (I473877,I473860,I207260);
and I_27706 (I473894,I473696,I473877);
nor I_27707 (I473911,I473809,I473894);
DFFARX1 I_27708 (I473911,I2859,I473614,I473582,);
DFFARX1 I_27709 (I473894,I2859,I473614,I473603,);
nor I_27710 (I473956,I207284,I207260);
nor I_27711 (I473594,I473809,I473956);
or I_27712 (I473987,I207284,I207260);
nor I_27713 (I474004,I207266,I207275);
DFFARX1 I_27714 (I474004,I2859,I473614,I474030,);
not I_27715 (I474038,I474030);
nor I_27716 (I473600,I474038,I473843);
nand I_27717 (I474069,I474038,I473688);
not I_27718 (I474086,I207266);
nand I_27719 (I474103,I474086,I473792);
nand I_27720 (I474120,I474038,I474103);
nand I_27721 (I473591,I474120,I474069);
nand I_27722 (I473588,I474103,I473987);
not I_27723 (I474192,I2866);
DFFARX1 I_27724 (I400573,I2859,I474192,I474218,);
and I_27725 (I474226,I474218,I400567);
DFFARX1 I_27726 (I474226,I2859,I474192,I474175,);
DFFARX1 I_27727 (I400585,I2859,I474192,I474266,);
not I_27728 (I474274,I400576);
not I_27729 (I474291,I400588);
nand I_27730 (I474308,I474291,I474274);
nor I_27731 (I474163,I474266,I474308);
DFFARX1 I_27732 (I474308,I2859,I474192,I474348,);
not I_27733 (I474184,I474348);
not I_27734 (I474370,I400594);
nand I_27735 (I474387,I474291,I474370);
DFFARX1 I_27736 (I474387,I2859,I474192,I474413,);
not I_27737 (I474421,I474413);
not I_27738 (I474438,I400570);
nand I_27739 (I474455,I474438,I400591);
and I_27740 (I474472,I474274,I474455);
nor I_27741 (I474489,I474387,I474472);
DFFARX1 I_27742 (I474489,I2859,I474192,I474160,);
DFFARX1 I_27743 (I474472,I2859,I474192,I474181,);
nor I_27744 (I474534,I400570,I400582);
nor I_27745 (I474172,I474387,I474534);
or I_27746 (I474565,I400570,I400582);
nor I_27747 (I474582,I400567,I400579);
DFFARX1 I_27748 (I474582,I2859,I474192,I474608,);
not I_27749 (I474616,I474608);
nor I_27750 (I474178,I474616,I474421);
nand I_27751 (I474647,I474616,I474266);
not I_27752 (I474664,I400567);
nand I_27753 (I474681,I474664,I474370);
nand I_27754 (I474698,I474616,I474681);
nand I_27755 (I474169,I474698,I474647);
nand I_27756 (I474166,I474681,I474565);
not I_27757 (I474770,I2866);
DFFARX1 I_27758 (I262015,I2859,I474770,I474796,);
and I_27759 (I474804,I474796,I262003);
DFFARX1 I_27760 (I474804,I2859,I474770,I474753,);
DFFARX1 I_27761 (I262006,I2859,I474770,I474844,);
not I_27762 (I474852,I262000);
not I_27763 (I474869,I262024);
nand I_27764 (I474886,I474869,I474852);
nor I_27765 (I474741,I474844,I474886);
DFFARX1 I_27766 (I474886,I2859,I474770,I474926,);
not I_27767 (I474762,I474926);
not I_27768 (I474948,I262012);
nand I_27769 (I474965,I474869,I474948);
DFFARX1 I_27770 (I474965,I2859,I474770,I474991,);
not I_27771 (I474999,I474991);
not I_27772 (I475016,I262021);
nand I_27773 (I475033,I475016,I262018);
and I_27774 (I475050,I474852,I475033);
nor I_27775 (I475067,I474965,I475050);
DFFARX1 I_27776 (I475067,I2859,I474770,I474738,);
DFFARX1 I_27777 (I475050,I2859,I474770,I474759,);
nor I_27778 (I475112,I262021,I262009);
nor I_27779 (I474750,I474965,I475112);
or I_27780 (I475143,I262021,I262009);
nor I_27781 (I475160,I262000,I262003);
DFFARX1 I_27782 (I475160,I2859,I474770,I475186,);
not I_27783 (I475194,I475186);
nor I_27784 (I474756,I475194,I474999);
nand I_27785 (I475225,I475194,I474844);
not I_27786 (I475242,I262000);
nand I_27787 (I475259,I475242,I474948);
nand I_27788 (I475276,I475194,I475259);
nand I_27789 (I474747,I475276,I475225);
nand I_27790 (I474744,I475259,I475143);
not I_27791 (I475348,I2866);
DFFARX1 I_27792 (I298429,I2859,I475348,I475374,);
and I_27793 (I475382,I475374,I298417);
DFFARX1 I_27794 (I475382,I2859,I475348,I475331,);
DFFARX1 I_27795 (I298420,I2859,I475348,I475422,);
not I_27796 (I475430,I298414);
not I_27797 (I475447,I298438);
nand I_27798 (I475464,I475447,I475430);
nor I_27799 (I475319,I475422,I475464);
DFFARX1 I_27800 (I475464,I2859,I475348,I475504,);
not I_27801 (I475340,I475504);
not I_27802 (I475526,I298426);
nand I_27803 (I475543,I475447,I475526);
DFFARX1 I_27804 (I475543,I2859,I475348,I475569,);
not I_27805 (I475577,I475569);
not I_27806 (I475594,I298435);
nand I_27807 (I475611,I475594,I298432);
and I_27808 (I475628,I475430,I475611);
nor I_27809 (I475645,I475543,I475628);
DFFARX1 I_27810 (I475645,I2859,I475348,I475316,);
DFFARX1 I_27811 (I475628,I2859,I475348,I475337,);
nor I_27812 (I475690,I298435,I298423);
nor I_27813 (I475328,I475543,I475690);
or I_27814 (I475721,I298435,I298423);
nor I_27815 (I475738,I298414,I298417);
DFFARX1 I_27816 (I475738,I2859,I475348,I475764,);
not I_27817 (I475772,I475764);
nor I_27818 (I475334,I475772,I475577);
nand I_27819 (I475803,I475772,I475422);
not I_27820 (I475820,I298414);
nand I_27821 (I475837,I475820,I475526);
nand I_27822 (I475854,I475772,I475837);
nand I_27823 (I475325,I475854,I475803);
nand I_27824 (I475322,I475837,I475721);
not I_27825 (I475926,I2866);
DFFARX1 I_27826 (I553492,I2859,I475926,I475952,);
and I_27827 (I475960,I475952,I553474);
DFFARX1 I_27828 (I475960,I2859,I475926,I475909,);
DFFARX1 I_27829 (I553465,I2859,I475926,I476000,);
not I_27830 (I476008,I553480);
not I_27831 (I476025,I553468);
nand I_27832 (I476042,I476025,I476008);
nor I_27833 (I475897,I476000,I476042);
DFFARX1 I_27834 (I476042,I2859,I475926,I476082,);
not I_27835 (I475918,I476082);
not I_27836 (I476104,I553477);
nand I_27837 (I476121,I476025,I476104);
DFFARX1 I_27838 (I476121,I2859,I475926,I476147,);
not I_27839 (I476155,I476147);
not I_27840 (I476172,I553486);
nand I_27841 (I476189,I476172,I553465);
and I_27842 (I476206,I476008,I476189);
nor I_27843 (I476223,I476121,I476206);
DFFARX1 I_27844 (I476223,I2859,I475926,I475894,);
DFFARX1 I_27845 (I476206,I2859,I475926,I475915,);
nor I_27846 (I476268,I553486,I553489);
nor I_27847 (I475906,I476121,I476268);
or I_27848 (I476299,I553486,I553489);
nor I_27849 (I476316,I553483,I553471);
DFFARX1 I_27850 (I476316,I2859,I475926,I476342,);
not I_27851 (I476350,I476342);
nor I_27852 (I475912,I476350,I476155);
nand I_27853 (I476381,I476350,I476000);
not I_27854 (I476398,I553483);
nand I_27855 (I476415,I476398,I476104);
nand I_27856 (I476432,I476350,I476415);
nand I_27857 (I475903,I476432,I476381);
nand I_27858 (I475900,I476415,I476299);
not I_27859 (I476504,I2866);
DFFARX1 I_27860 (I503047,I2859,I476504,I476530,);
and I_27861 (I476538,I476530,I503041);
DFFARX1 I_27862 (I476538,I2859,I476504,I476487,);
DFFARX1 I_27863 (I503026,I2859,I476504,I476578,);
not I_27864 (I476586,I503032);
not I_27865 (I476603,I503044);
nand I_27866 (I476620,I476603,I476586);
nor I_27867 (I476475,I476578,I476620);
DFFARX1 I_27868 (I476620,I2859,I476504,I476660,);
not I_27869 (I476496,I476660);
not I_27870 (I476682,I503026);
nand I_27871 (I476699,I476603,I476682);
DFFARX1 I_27872 (I476699,I2859,I476504,I476725,);
not I_27873 (I476733,I476725);
not I_27874 (I476750,I503050);
nand I_27875 (I476767,I476750,I503038);
and I_27876 (I476784,I476586,I476767);
nor I_27877 (I476801,I476699,I476784);
DFFARX1 I_27878 (I476801,I2859,I476504,I476472,);
DFFARX1 I_27879 (I476784,I2859,I476504,I476493,);
nor I_27880 (I476846,I503050,I503029);
nor I_27881 (I476484,I476699,I476846);
or I_27882 (I476877,I503050,I503029);
nor I_27883 (I476894,I503035,I503029);
DFFARX1 I_27884 (I476894,I2859,I476504,I476920,);
not I_27885 (I476928,I476920);
nor I_27886 (I476490,I476928,I476733);
nand I_27887 (I476959,I476928,I476578);
not I_27888 (I476976,I503035);
nand I_27889 (I476993,I476976,I476682);
nand I_27890 (I477010,I476928,I476993);
nand I_27891 (I476481,I477010,I476959);
nand I_27892 (I476478,I476993,I476877);
not I_27893 (I477082,I2866);
DFFARX1 I_27894 (I27475,I2859,I477082,I477108,);
and I_27895 (I477116,I477108,I27451);
DFFARX1 I_27896 (I477116,I2859,I477082,I477065,);
DFFARX1 I_27897 (I27469,I2859,I477082,I477156,);
not I_27898 (I477164,I27457);
not I_27899 (I477181,I27454);
nand I_27900 (I477198,I477181,I477164);
nor I_27901 (I477053,I477156,I477198);
DFFARX1 I_27902 (I477198,I2859,I477082,I477238,);
not I_27903 (I477074,I477238);
not I_27904 (I477260,I27463);
nand I_27905 (I477277,I477181,I477260);
DFFARX1 I_27906 (I477277,I2859,I477082,I477303,);
not I_27907 (I477311,I477303);
not I_27908 (I477328,I27454);
nand I_27909 (I477345,I477328,I27472);
and I_27910 (I477362,I477164,I477345);
nor I_27911 (I477379,I477277,I477362);
DFFARX1 I_27912 (I477379,I2859,I477082,I477050,);
DFFARX1 I_27913 (I477362,I2859,I477082,I477071,);
nor I_27914 (I477424,I27454,I27466);
nor I_27915 (I477062,I477277,I477424);
or I_27916 (I477455,I27454,I27466);
nor I_27917 (I477472,I27460,I27451);
DFFARX1 I_27918 (I477472,I2859,I477082,I477498,);
not I_27919 (I477506,I477498);
nor I_27920 (I477068,I477506,I477311);
nand I_27921 (I477537,I477506,I477156);
not I_27922 (I477554,I27460);
nand I_27923 (I477571,I477554,I477260);
nand I_27924 (I477588,I477506,I477571);
nand I_27925 (I477059,I477588,I477537);
nand I_27926 (I477056,I477571,I477455);
not I_27927 (I477660,I2866);
DFFARX1 I_27928 (I152530,I2859,I477660,I477686,);
and I_27929 (I477694,I477686,I152515);
DFFARX1 I_27930 (I477694,I2859,I477660,I477643,);
DFFARX1 I_27931 (I152521,I2859,I477660,I477734,);
not I_27932 (I477742,I152503);
not I_27933 (I477759,I152524);
nand I_27934 (I477776,I477759,I477742);
nor I_27935 (I477631,I477734,I477776);
DFFARX1 I_27936 (I477776,I2859,I477660,I477816,);
not I_27937 (I477652,I477816);
not I_27938 (I477838,I152527);
nand I_27939 (I477855,I477759,I477838);
DFFARX1 I_27940 (I477855,I2859,I477660,I477881,);
not I_27941 (I477889,I477881);
not I_27942 (I477906,I152518);
nand I_27943 (I477923,I477906,I152506);
and I_27944 (I477940,I477742,I477923);
nor I_27945 (I477957,I477855,I477940);
DFFARX1 I_27946 (I477957,I2859,I477660,I477628,);
DFFARX1 I_27947 (I477940,I2859,I477660,I477649,);
nor I_27948 (I478002,I152518,I152512);
nor I_27949 (I477640,I477855,I478002);
or I_27950 (I478033,I152518,I152512);
nor I_27951 (I478050,I152509,I152503);
DFFARX1 I_27952 (I478050,I2859,I477660,I478076,);
not I_27953 (I478084,I478076);
nor I_27954 (I477646,I478084,I477889);
nand I_27955 (I478115,I478084,I477734);
not I_27956 (I478132,I152509);
nand I_27957 (I478149,I478132,I477838);
nand I_27958 (I478166,I478084,I478149);
nand I_27959 (I477637,I478166,I478115);
nand I_27960 (I477634,I478149,I478033);
not I_27961 (I478238,I2866);
DFFARX1 I_27962 (I121437,I2859,I478238,I478264,);
and I_27963 (I478272,I478264,I121422);
DFFARX1 I_27964 (I478272,I2859,I478238,I478221,);
DFFARX1 I_27965 (I121428,I2859,I478238,I478312,);
not I_27966 (I478320,I121410);
not I_27967 (I478337,I121431);
nand I_27968 (I478354,I478337,I478320);
nor I_27969 (I478209,I478312,I478354);
DFFARX1 I_27970 (I478354,I2859,I478238,I478394,);
not I_27971 (I478230,I478394);
not I_27972 (I478416,I121434);
nand I_27973 (I478433,I478337,I478416);
DFFARX1 I_27974 (I478433,I2859,I478238,I478459,);
not I_27975 (I478467,I478459);
not I_27976 (I478484,I121425);
nand I_27977 (I478501,I478484,I121413);
and I_27978 (I478518,I478320,I478501);
nor I_27979 (I478535,I478433,I478518);
DFFARX1 I_27980 (I478535,I2859,I478238,I478206,);
DFFARX1 I_27981 (I478518,I2859,I478238,I478227,);
nor I_27982 (I478580,I121425,I121419);
nor I_27983 (I478218,I478433,I478580);
or I_27984 (I478611,I121425,I121419);
nor I_27985 (I478628,I121416,I121410);
DFFARX1 I_27986 (I478628,I2859,I478238,I478654,);
not I_27987 (I478662,I478654);
nor I_27988 (I478224,I478662,I478467);
nand I_27989 (I478693,I478662,I478312);
not I_27990 (I478710,I121416);
nand I_27991 (I478727,I478710,I478416);
nand I_27992 (I478744,I478662,I478727);
nand I_27993 (I478215,I478744,I478693);
nand I_27994 (I478212,I478727,I478611);
not I_27995 (I478816,I2866);
DFFARX1 I_27996 (I223867,I2859,I478816,I478842,);
and I_27997 (I478850,I478842,I223855);
DFFARX1 I_27998 (I478850,I2859,I478816,I478799,);
DFFARX1 I_27999 (I223870,I2859,I478816,I478890,);
not I_28000 (I478898,I223861);
not I_28001 (I478915,I223852);
nand I_28002 (I478932,I478915,I478898);
nor I_28003 (I478787,I478890,I478932);
DFFARX1 I_28004 (I478932,I2859,I478816,I478972,);
not I_28005 (I478808,I478972);
not I_28006 (I478994,I223858);
nand I_28007 (I479011,I478915,I478994);
DFFARX1 I_28008 (I479011,I2859,I478816,I479037,);
not I_28009 (I479045,I479037);
not I_28010 (I479062,I223873);
nand I_28011 (I479079,I479062,I223876);
and I_28012 (I479096,I478898,I479079);
nor I_28013 (I479113,I479011,I479096);
DFFARX1 I_28014 (I479113,I2859,I478816,I478784,);
DFFARX1 I_28015 (I479096,I2859,I478816,I478805,);
nor I_28016 (I479158,I223873,I223852);
nor I_28017 (I478796,I479011,I479158);
or I_28018 (I479189,I223873,I223852);
nor I_28019 (I479206,I223864,I223855);
DFFARX1 I_28020 (I479206,I2859,I478816,I479232,);
not I_28021 (I479240,I479232);
nor I_28022 (I478802,I479240,I479045);
nand I_28023 (I479271,I479240,I478890);
not I_28024 (I479288,I223864);
nand I_28025 (I479305,I479288,I478994);
nand I_28026 (I479322,I479240,I479305);
nand I_28027 (I478793,I479322,I479271);
nand I_28028 (I478790,I479305,I479189);
not I_28029 (I479394,I2866);
DFFARX1 I_28030 (I307677,I2859,I479394,I479420,);
and I_28031 (I479428,I479420,I307665);
DFFARX1 I_28032 (I479428,I2859,I479394,I479377,);
DFFARX1 I_28033 (I307668,I2859,I479394,I479468,);
not I_28034 (I479476,I307662);
not I_28035 (I479493,I307686);
nand I_28036 (I479510,I479493,I479476);
nor I_28037 (I479365,I479468,I479510);
DFFARX1 I_28038 (I479510,I2859,I479394,I479550,);
not I_28039 (I479386,I479550);
not I_28040 (I479572,I307674);
nand I_28041 (I479589,I479493,I479572);
DFFARX1 I_28042 (I479589,I2859,I479394,I479615,);
not I_28043 (I479623,I479615);
not I_28044 (I479640,I307683);
nand I_28045 (I479657,I479640,I307680);
and I_28046 (I479674,I479476,I479657);
nor I_28047 (I479691,I479589,I479674);
DFFARX1 I_28048 (I479691,I2859,I479394,I479362,);
DFFARX1 I_28049 (I479674,I2859,I479394,I479383,);
nor I_28050 (I479736,I307683,I307671);
nor I_28051 (I479374,I479589,I479736);
or I_28052 (I479767,I307683,I307671);
nor I_28053 (I479784,I307662,I307665);
DFFARX1 I_28054 (I479784,I2859,I479394,I479810,);
not I_28055 (I479818,I479810);
nor I_28056 (I479380,I479818,I479623);
nand I_28057 (I479849,I479818,I479468);
not I_28058 (I479866,I307662);
nand I_28059 (I479883,I479866,I479572);
nand I_28060 (I479900,I479818,I479883);
nand I_28061 (I479371,I479900,I479849);
nand I_28062 (I479368,I479883,I479767);
not I_28063 (I479972,I2866);
DFFARX1 I_28064 (I123018,I2859,I479972,I479998,);
and I_28065 (I480006,I479998,I123003);
DFFARX1 I_28066 (I480006,I2859,I479972,I479955,);
DFFARX1 I_28067 (I123009,I2859,I479972,I480046,);
not I_28068 (I480054,I122991);
not I_28069 (I480071,I123012);
nand I_28070 (I480088,I480071,I480054);
nor I_28071 (I479943,I480046,I480088);
DFFARX1 I_28072 (I480088,I2859,I479972,I480128,);
not I_28073 (I479964,I480128);
not I_28074 (I480150,I123015);
nand I_28075 (I480167,I480071,I480150);
DFFARX1 I_28076 (I480167,I2859,I479972,I480193,);
not I_28077 (I480201,I480193);
not I_28078 (I480218,I123006);
nand I_28079 (I480235,I480218,I122994);
and I_28080 (I480252,I480054,I480235);
nor I_28081 (I480269,I480167,I480252);
DFFARX1 I_28082 (I480269,I2859,I479972,I479940,);
DFFARX1 I_28083 (I480252,I2859,I479972,I479961,);
nor I_28084 (I480314,I123006,I123000);
nor I_28085 (I479952,I480167,I480314);
or I_28086 (I480345,I123006,I123000);
nor I_28087 (I480362,I122997,I122991);
DFFARX1 I_28088 (I480362,I2859,I479972,I480388,);
not I_28089 (I480396,I480388);
nor I_28090 (I479958,I480396,I480201);
nand I_28091 (I480427,I480396,I480046);
not I_28092 (I480444,I122997);
nand I_28093 (I480461,I480444,I480150);
nand I_28094 (I480478,I480396,I480461);
nand I_28095 (I479949,I480478,I480427);
nand I_28096 (I479946,I480461,I480345);
not I_28097 (I480550,I2866);
DFFARX1 I_28098 (I433856,I2859,I480550,I480576,);
and I_28099 (I480584,I480576,I433853);
DFFARX1 I_28100 (I480584,I2859,I480550,I480533,);
DFFARX1 I_28101 (I433859,I2859,I480550,I480624,);
not I_28102 (I480632,I433862);
not I_28103 (I480649,I433856);
nand I_28104 (I480666,I480649,I480632);
nor I_28105 (I480521,I480624,I480666);
DFFARX1 I_28106 (I480666,I2859,I480550,I480706,);
not I_28107 (I480542,I480706);
not I_28108 (I480728,I433871);
nand I_28109 (I480745,I480649,I480728);
DFFARX1 I_28110 (I480745,I2859,I480550,I480771,);
not I_28111 (I480779,I480771);
not I_28112 (I480796,I433868);
nand I_28113 (I480813,I480796,I433874);
and I_28114 (I480830,I480632,I480813);
nor I_28115 (I480847,I480745,I480830);
DFFARX1 I_28116 (I480847,I2859,I480550,I480518,);
DFFARX1 I_28117 (I480830,I2859,I480550,I480539,);
nor I_28118 (I480892,I433868,I433853);
nor I_28119 (I480530,I480745,I480892);
or I_28120 (I480923,I433868,I433853);
nor I_28121 (I480940,I433865,I433859);
DFFARX1 I_28122 (I480940,I2859,I480550,I480966,);
not I_28123 (I480974,I480966);
nor I_28124 (I480536,I480974,I480779);
nand I_28125 (I481005,I480974,I480624);
not I_28126 (I481022,I433865);
nand I_28127 (I481039,I481022,I480728);
nand I_28128 (I481056,I480974,I481039);
nand I_28129 (I480527,I481056,I481005);
nand I_28130 (I480524,I481039,I480923);
not I_28131 (I481128,I2866);
DFFARX1 I_28132 (I549922,I2859,I481128,I481154,);
and I_28133 (I481162,I481154,I549904);
DFFARX1 I_28134 (I481162,I2859,I481128,I481111,);
DFFARX1 I_28135 (I549895,I2859,I481128,I481202,);
not I_28136 (I481210,I549910);
not I_28137 (I481227,I549898);
nand I_28138 (I481244,I481227,I481210);
nor I_28139 (I481099,I481202,I481244);
DFFARX1 I_28140 (I481244,I2859,I481128,I481284,);
not I_28141 (I481120,I481284);
not I_28142 (I481306,I549907);
nand I_28143 (I481323,I481227,I481306);
DFFARX1 I_28144 (I481323,I2859,I481128,I481349,);
not I_28145 (I481357,I481349);
not I_28146 (I481374,I549916);
nand I_28147 (I481391,I481374,I549895);
and I_28148 (I481408,I481210,I481391);
nor I_28149 (I481425,I481323,I481408);
DFFARX1 I_28150 (I481425,I2859,I481128,I481096,);
DFFARX1 I_28151 (I481408,I2859,I481128,I481117,);
nor I_28152 (I481470,I549916,I549919);
nor I_28153 (I481108,I481323,I481470);
or I_28154 (I481501,I549916,I549919);
nor I_28155 (I481518,I549913,I549901);
DFFARX1 I_28156 (I481518,I2859,I481128,I481544,);
not I_28157 (I481552,I481544);
nor I_28158 (I481114,I481552,I481357);
nand I_28159 (I481583,I481552,I481202);
not I_28160 (I481600,I549913);
nand I_28161 (I481617,I481600,I481306);
nand I_28162 (I481634,I481552,I481617);
nand I_28163 (I481105,I481634,I481583);
nand I_28164 (I481102,I481617,I481501);
not I_28165 (I481706,I2866);
DFFARX1 I_28166 (I326501,I2859,I481706,I481732,);
and I_28167 (I481740,I481732,I326507);
DFFARX1 I_28168 (I481740,I2859,I481706,I481689,);
DFFARX1 I_28169 (I326513,I2859,I481706,I481780,);
not I_28170 (I481788,I326498);
not I_28171 (I481805,I326498);
nand I_28172 (I481822,I481805,I481788);
nor I_28173 (I481677,I481780,I481822);
DFFARX1 I_28174 (I481822,I2859,I481706,I481862,);
not I_28175 (I481698,I481862);
not I_28176 (I481884,I326516);
nand I_28177 (I481901,I481805,I481884);
DFFARX1 I_28178 (I481901,I2859,I481706,I481927,);
not I_28179 (I481935,I481927);
not I_28180 (I481952,I326510);
nand I_28181 (I481969,I481952,I326501);
and I_28182 (I481986,I481788,I481969);
nor I_28183 (I482003,I481901,I481986);
DFFARX1 I_28184 (I482003,I2859,I481706,I481674,);
DFFARX1 I_28185 (I481986,I2859,I481706,I481695,);
nor I_28186 (I482048,I326510,I326519);
nor I_28187 (I481686,I481901,I482048);
or I_28188 (I482079,I326510,I326519);
nor I_28189 (I482096,I326504,I326504);
DFFARX1 I_28190 (I482096,I2859,I481706,I482122,);
not I_28191 (I482130,I482122);
nor I_28192 (I481692,I482130,I481935);
nand I_28193 (I482161,I482130,I481780);
not I_28194 (I482178,I326504);
nand I_28195 (I482195,I482178,I481884);
nand I_28196 (I482212,I482130,I482195);
nand I_28197 (I481683,I482212,I482161);
nand I_28198 (I481680,I482195,I482079);
not I_28199 (I482284,I2866);
DFFARX1 I_28200 (I545757,I2859,I482284,I482310,);
and I_28201 (I482318,I482310,I545739);
DFFARX1 I_28202 (I482318,I2859,I482284,I482267,);
DFFARX1 I_28203 (I545730,I2859,I482284,I482358,);
not I_28204 (I482366,I545745);
not I_28205 (I482383,I545733);
nand I_28206 (I482400,I482383,I482366);
nor I_28207 (I482255,I482358,I482400);
DFFARX1 I_28208 (I482400,I2859,I482284,I482440,);
not I_28209 (I482276,I482440);
not I_28210 (I482462,I545742);
nand I_28211 (I482479,I482383,I482462);
DFFARX1 I_28212 (I482479,I2859,I482284,I482505,);
not I_28213 (I482513,I482505);
not I_28214 (I482530,I545751);
nand I_28215 (I482547,I482530,I545730);
and I_28216 (I482564,I482366,I482547);
nor I_28217 (I482581,I482479,I482564);
DFFARX1 I_28218 (I482581,I2859,I482284,I482252,);
DFFARX1 I_28219 (I482564,I2859,I482284,I482273,);
nor I_28220 (I482626,I545751,I545754);
nor I_28221 (I482264,I482479,I482626);
or I_28222 (I482657,I545751,I545754);
nor I_28223 (I482674,I545748,I545736);
DFFARX1 I_28224 (I482674,I2859,I482284,I482700,);
not I_28225 (I482708,I482700);
nor I_28226 (I482270,I482708,I482513);
nand I_28227 (I482739,I482708,I482358);
not I_28228 (I482756,I545748);
nand I_28229 (I482773,I482756,I482462);
nand I_28230 (I482790,I482708,I482773);
nand I_28231 (I482261,I482790,I482739);
nand I_28232 (I482258,I482773,I482657);
not I_28233 (I482862,I2866);
DFFARX1 I_28234 (I289181,I2859,I482862,I482888,);
and I_28235 (I482896,I482888,I289169);
DFFARX1 I_28236 (I482896,I2859,I482862,I482845,);
DFFARX1 I_28237 (I289172,I2859,I482862,I482936,);
not I_28238 (I482944,I289166);
not I_28239 (I482961,I289190);
nand I_28240 (I482978,I482961,I482944);
nor I_28241 (I482833,I482936,I482978);
DFFARX1 I_28242 (I482978,I2859,I482862,I483018,);
not I_28243 (I482854,I483018);
not I_28244 (I483040,I289178);
nand I_28245 (I483057,I482961,I483040);
DFFARX1 I_28246 (I483057,I2859,I482862,I483083,);
not I_28247 (I483091,I483083);
not I_28248 (I483108,I289187);
nand I_28249 (I483125,I483108,I289184);
and I_28250 (I483142,I482944,I483125);
nor I_28251 (I483159,I483057,I483142);
DFFARX1 I_28252 (I483159,I2859,I482862,I482830,);
DFFARX1 I_28253 (I483142,I2859,I482862,I482851,);
nor I_28254 (I483204,I289187,I289175);
nor I_28255 (I482842,I483057,I483204);
or I_28256 (I483235,I289187,I289175);
nor I_28257 (I483252,I289166,I289169);
DFFARX1 I_28258 (I483252,I2859,I482862,I483278,);
not I_28259 (I483286,I483278);
nor I_28260 (I482848,I483286,I483091);
nand I_28261 (I483317,I483286,I482936);
not I_28262 (I483334,I289166);
nand I_28263 (I483351,I483334,I483040);
nand I_28264 (I483368,I483286,I483351);
nand I_28265 (I482839,I483368,I483317);
nand I_28266 (I482836,I483351,I483235);
not I_28267 (I483440,I2866);
DFFARX1 I_28268 (I416465,I2859,I483440,I483466,);
and I_28269 (I483474,I483466,I416462);
DFFARX1 I_28270 (I483474,I2859,I483440,I483423,);
DFFARX1 I_28271 (I416468,I2859,I483440,I483514,);
not I_28272 (I483522,I416471);
not I_28273 (I483539,I416465);
nand I_28274 (I483556,I483539,I483522);
nor I_28275 (I483411,I483514,I483556);
DFFARX1 I_28276 (I483556,I2859,I483440,I483596,);
not I_28277 (I483432,I483596);
not I_28278 (I483618,I416480);
nand I_28279 (I483635,I483539,I483618);
DFFARX1 I_28280 (I483635,I2859,I483440,I483661,);
not I_28281 (I483669,I483661);
not I_28282 (I483686,I416477);
nand I_28283 (I483703,I483686,I416483);
and I_28284 (I483720,I483522,I483703);
nor I_28285 (I483737,I483635,I483720);
DFFARX1 I_28286 (I483737,I2859,I483440,I483408,);
DFFARX1 I_28287 (I483720,I2859,I483440,I483429,);
nor I_28288 (I483782,I416477,I416462);
nor I_28289 (I483420,I483635,I483782);
or I_28290 (I483813,I416477,I416462);
nor I_28291 (I483830,I416474,I416468);
DFFARX1 I_28292 (I483830,I2859,I483440,I483856,);
not I_28293 (I483864,I483856);
nor I_28294 (I483426,I483864,I483669);
nand I_28295 (I483895,I483864,I483514);
not I_28296 (I483912,I416474);
nand I_28297 (I483929,I483912,I483618);
nand I_28298 (I483946,I483864,I483929);
nand I_28299 (I483417,I483946,I483895);
nand I_28300 (I483414,I483929,I483813);
not I_28301 (I484018,I2866);
DFFARX1 I_28302 (I158327,I2859,I484018,I484044,);
and I_28303 (I484052,I484044,I158312);
DFFARX1 I_28304 (I484052,I2859,I484018,I484001,);
DFFARX1 I_28305 (I158318,I2859,I484018,I484092,);
not I_28306 (I484100,I158300);
not I_28307 (I484117,I158321);
nand I_28308 (I484134,I484117,I484100);
nor I_28309 (I483989,I484092,I484134);
DFFARX1 I_28310 (I484134,I2859,I484018,I484174,);
not I_28311 (I484010,I484174);
not I_28312 (I484196,I158324);
nand I_28313 (I484213,I484117,I484196);
DFFARX1 I_28314 (I484213,I2859,I484018,I484239,);
not I_28315 (I484247,I484239);
not I_28316 (I484264,I158315);
nand I_28317 (I484281,I484264,I158303);
and I_28318 (I484298,I484100,I484281);
nor I_28319 (I484315,I484213,I484298);
DFFARX1 I_28320 (I484315,I2859,I484018,I483986,);
DFFARX1 I_28321 (I484298,I2859,I484018,I484007,);
nor I_28322 (I484360,I158315,I158309);
nor I_28323 (I483998,I484213,I484360);
or I_28324 (I484391,I158315,I158309);
nor I_28325 (I484408,I158306,I158300);
DFFARX1 I_28326 (I484408,I2859,I484018,I484434,);
not I_28327 (I484442,I484434);
nor I_28328 (I484004,I484442,I484247);
nand I_28329 (I484473,I484442,I484092);
not I_28330 (I484490,I158306);
nand I_28331 (I484507,I484490,I484196);
nand I_28332 (I484524,I484442,I484507);
nand I_28333 (I483995,I484524,I484473);
nand I_28334 (I483992,I484507,I484391);
not I_28335 (I484596,I2866);
DFFARX1 I_28336 (I555277,I2859,I484596,I484622,);
and I_28337 (I484630,I484622,I555259);
DFFARX1 I_28338 (I484630,I2859,I484596,I484579,);
DFFARX1 I_28339 (I555250,I2859,I484596,I484670,);
not I_28340 (I484678,I555265);
not I_28341 (I484695,I555253);
nand I_28342 (I484712,I484695,I484678);
nor I_28343 (I484567,I484670,I484712);
DFFARX1 I_28344 (I484712,I2859,I484596,I484752,);
not I_28345 (I484588,I484752);
not I_28346 (I484774,I555262);
nand I_28347 (I484791,I484695,I484774);
DFFARX1 I_28348 (I484791,I2859,I484596,I484817,);
not I_28349 (I484825,I484817);
not I_28350 (I484842,I555271);
nand I_28351 (I484859,I484842,I555250);
and I_28352 (I484876,I484678,I484859);
nor I_28353 (I484893,I484791,I484876);
DFFARX1 I_28354 (I484893,I2859,I484596,I484564,);
DFFARX1 I_28355 (I484876,I2859,I484596,I484585,);
nor I_28356 (I484938,I555271,I555274);
nor I_28357 (I484576,I484791,I484938);
or I_28358 (I484969,I555271,I555274);
nor I_28359 (I484986,I555268,I555256);
DFFARX1 I_28360 (I484986,I2859,I484596,I485012,);
not I_28361 (I485020,I485012);
nor I_28362 (I484582,I485020,I484825);
nand I_28363 (I485051,I485020,I484670);
not I_28364 (I485068,I555268);
nand I_28365 (I485085,I485068,I484774);
nand I_28366 (I485102,I485020,I485085);
nand I_28367 (I484573,I485102,I485051);
nand I_28368 (I484570,I485085,I484969);
not I_28369 (I485174,I2866);
DFFARX1 I_28370 (I429368,I2859,I485174,I485200,);
and I_28371 (I485208,I485200,I429365);
DFFARX1 I_28372 (I485208,I2859,I485174,I485157,);
DFFARX1 I_28373 (I429371,I2859,I485174,I485248,);
not I_28374 (I485256,I429374);
not I_28375 (I485273,I429368);
nand I_28376 (I485290,I485273,I485256);
nor I_28377 (I485145,I485248,I485290);
DFFARX1 I_28378 (I485290,I2859,I485174,I485330,);
not I_28379 (I485166,I485330);
not I_28380 (I485352,I429383);
nand I_28381 (I485369,I485273,I485352);
DFFARX1 I_28382 (I485369,I2859,I485174,I485395,);
not I_28383 (I485403,I485395);
not I_28384 (I485420,I429380);
nand I_28385 (I485437,I485420,I429386);
and I_28386 (I485454,I485256,I485437);
nor I_28387 (I485471,I485369,I485454);
DFFARX1 I_28388 (I485471,I2859,I485174,I485142,);
DFFARX1 I_28389 (I485454,I2859,I485174,I485163,);
nor I_28390 (I485516,I429380,I429365);
nor I_28391 (I485154,I485369,I485516);
or I_28392 (I485547,I429380,I429365);
nor I_28393 (I485564,I429377,I429371);
DFFARX1 I_28394 (I485564,I2859,I485174,I485590,);
not I_28395 (I485598,I485590);
nor I_28396 (I485160,I485598,I485403);
nand I_28397 (I485629,I485598,I485248);
not I_28398 (I485646,I429377);
nand I_28399 (I485663,I485646,I485352);
nand I_28400 (I485680,I485598,I485663);
nand I_28401 (I485151,I485680,I485629);
nand I_28402 (I485148,I485663,I485547);
not I_28403 (I485752,I2866);
DFFARX1 I_28404 (I35380,I2859,I485752,I485778,);
and I_28405 (I485786,I485778,I35356);
DFFARX1 I_28406 (I485786,I2859,I485752,I485735,);
DFFARX1 I_28407 (I35374,I2859,I485752,I485826,);
not I_28408 (I485834,I35362);
not I_28409 (I485851,I35359);
nand I_28410 (I485868,I485851,I485834);
nor I_28411 (I485723,I485826,I485868);
DFFARX1 I_28412 (I485868,I2859,I485752,I485908,);
not I_28413 (I485744,I485908);
not I_28414 (I485930,I35368);
nand I_28415 (I485947,I485851,I485930);
DFFARX1 I_28416 (I485947,I2859,I485752,I485973,);
not I_28417 (I485981,I485973);
not I_28418 (I485998,I35359);
nand I_28419 (I486015,I485998,I35377);
and I_28420 (I486032,I485834,I486015);
nor I_28421 (I486049,I485947,I486032);
DFFARX1 I_28422 (I486049,I2859,I485752,I485720,);
DFFARX1 I_28423 (I486032,I2859,I485752,I485741,);
nor I_28424 (I486094,I35359,I35371);
nor I_28425 (I485732,I485947,I486094);
or I_28426 (I486125,I35359,I35371);
nor I_28427 (I486142,I35365,I35356);
DFFARX1 I_28428 (I486142,I2859,I485752,I486168,);
not I_28429 (I486176,I486168);
nor I_28430 (I485738,I486176,I485981);
nand I_28431 (I486207,I486176,I485826);
not I_28432 (I486224,I35365);
nand I_28433 (I486241,I486224,I485930);
nand I_28434 (I486258,I486176,I486241);
nand I_28435 (I485729,I486258,I486207);
nand I_28436 (I485726,I486241,I486125);
not I_28437 (I486330,I2866);
DFFARX1 I_28438 (I297273,I2859,I486330,I486356,);
and I_28439 (I486364,I486356,I297261);
DFFARX1 I_28440 (I486364,I2859,I486330,I486313,);
DFFARX1 I_28441 (I297264,I2859,I486330,I486404,);
not I_28442 (I486412,I297258);
not I_28443 (I486429,I297282);
nand I_28444 (I486446,I486429,I486412);
nor I_28445 (I486301,I486404,I486446);
DFFARX1 I_28446 (I486446,I2859,I486330,I486486,);
not I_28447 (I486322,I486486);
not I_28448 (I486508,I297270);
nand I_28449 (I486525,I486429,I486508);
DFFARX1 I_28450 (I486525,I2859,I486330,I486551,);
not I_28451 (I486559,I486551);
not I_28452 (I486576,I297279);
nand I_28453 (I486593,I486576,I297276);
and I_28454 (I486610,I486412,I486593);
nor I_28455 (I486627,I486525,I486610);
DFFARX1 I_28456 (I486627,I2859,I486330,I486298,);
DFFARX1 I_28457 (I486610,I2859,I486330,I486319,);
nor I_28458 (I486672,I297279,I297267);
nor I_28459 (I486310,I486525,I486672);
or I_28460 (I486703,I297279,I297267);
nor I_28461 (I486720,I297258,I297261);
DFFARX1 I_28462 (I486720,I2859,I486330,I486746,);
not I_28463 (I486754,I486746);
nor I_28464 (I486316,I486754,I486559);
nand I_28465 (I486785,I486754,I486404);
not I_28466 (I486802,I297258);
nand I_28467 (I486819,I486802,I486508);
nand I_28468 (I486836,I486754,I486819);
nand I_28469 (I486307,I486836,I486785);
nand I_28470 (I486304,I486819,I486703);
not I_28471 (I486908,I2866);
DFFARX1 I_28472 (I365689,I2859,I486908,I486934,);
and I_28473 (I486942,I486934,I365683);
DFFARX1 I_28474 (I486942,I2859,I486908,I486891,);
DFFARX1 I_28475 (I365701,I2859,I486908,I486982,);
not I_28476 (I486990,I365692);
not I_28477 (I487007,I365704);
nand I_28478 (I487024,I487007,I486990);
nor I_28479 (I486879,I486982,I487024);
DFFARX1 I_28480 (I487024,I2859,I486908,I487064,);
not I_28481 (I486900,I487064);
not I_28482 (I487086,I365710);
nand I_28483 (I487103,I487007,I487086);
DFFARX1 I_28484 (I487103,I2859,I486908,I487129,);
not I_28485 (I487137,I487129);
not I_28486 (I487154,I365686);
nand I_28487 (I487171,I487154,I365707);
and I_28488 (I487188,I486990,I487171);
nor I_28489 (I487205,I487103,I487188);
DFFARX1 I_28490 (I487205,I2859,I486908,I486876,);
DFFARX1 I_28491 (I487188,I2859,I486908,I486897,);
nor I_28492 (I487250,I365686,I365698);
nor I_28493 (I486888,I487103,I487250);
or I_28494 (I487281,I365686,I365698);
nor I_28495 (I487298,I365683,I365695);
DFFARX1 I_28496 (I487298,I2859,I486908,I487324,);
not I_28497 (I487332,I487324);
nor I_28498 (I486894,I487332,I487137);
nand I_28499 (I487363,I487332,I486982);
not I_28500 (I487380,I365683);
nand I_28501 (I487397,I487380,I487086);
nand I_28502 (I487414,I487332,I487397);
nand I_28503 (I486885,I487414,I487363);
nand I_28504 (I486882,I487397,I487281);
not I_28505 (I487486,I2866);
DFFARX1 I_28506 (I172376,I2859,I487486,I487512,);
and I_28507 (I487520,I487512,I172391);
DFFARX1 I_28508 (I487520,I2859,I487486,I487469,);
DFFARX1 I_28509 (I172394,I2859,I487486,I487560,);
not I_28510 (I487568,I172388);
not I_28511 (I487585,I172403);
nand I_28512 (I487602,I487585,I487568);
nor I_28513 (I487457,I487560,I487602);
DFFARX1 I_28514 (I487602,I2859,I487486,I487642,);
not I_28515 (I487478,I487642);
not I_28516 (I487664,I172379);
nand I_28517 (I487681,I487585,I487664);
DFFARX1 I_28518 (I487681,I2859,I487486,I487707,);
not I_28519 (I487715,I487707);
not I_28520 (I487732,I172382);
nand I_28521 (I487749,I487732,I172376);
and I_28522 (I487766,I487568,I487749);
nor I_28523 (I487783,I487681,I487766);
DFFARX1 I_28524 (I487783,I2859,I487486,I487454,);
DFFARX1 I_28525 (I487766,I2859,I487486,I487475,);
nor I_28526 (I487828,I172382,I172385);
nor I_28527 (I487466,I487681,I487828);
or I_28528 (I487859,I172382,I172385);
nor I_28529 (I487876,I172400,I172397);
DFFARX1 I_28530 (I487876,I2859,I487486,I487902,);
not I_28531 (I487910,I487902);
nor I_28532 (I487472,I487910,I487715);
nand I_28533 (I487941,I487910,I487560);
not I_28534 (I487958,I172400);
nand I_28535 (I487975,I487958,I487664);
nand I_28536 (I487992,I487910,I487975);
nand I_28537 (I487463,I487992,I487941);
nand I_28538 (I487460,I487975,I487859);
not I_28539 (I488064,I2866);
DFFARX1 I_28540 (I507943,I2859,I488064,I488090,);
and I_28541 (I488098,I488090,I507937);
DFFARX1 I_28542 (I488098,I2859,I488064,I488047,);
DFFARX1 I_28543 (I507922,I2859,I488064,I488138,);
not I_28544 (I488146,I507928);
not I_28545 (I488163,I507940);
nand I_28546 (I488180,I488163,I488146);
nor I_28547 (I488035,I488138,I488180);
DFFARX1 I_28548 (I488180,I2859,I488064,I488220,);
not I_28549 (I488056,I488220);
not I_28550 (I488242,I507922);
nand I_28551 (I488259,I488163,I488242);
DFFARX1 I_28552 (I488259,I2859,I488064,I488285,);
not I_28553 (I488293,I488285);
not I_28554 (I488310,I507946);
nand I_28555 (I488327,I488310,I507934);
and I_28556 (I488344,I488146,I488327);
nor I_28557 (I488361,I488259,I488344);
DFFARX1 I_28558 (I488361,I2859,I488064,I488032,);
DFFARX1 I_28559 (I488344,I2859,I488064,I488053,);
nor I_28560 (I488406,I507946,I507925);
nor I_28561 (I488044,I488259,I488406);
or I_28562 (I488437,I507946,I507925);
nor I_28563 (I488454,I507931,I507925);
DFFARX1 I_28564 (I488454,I2859,I488064,I488480,);
not I_28565 (I488488,I488480);
nor I_28566 (I488050,I488488,I488293);
nand I_28567 (I488519,I488488,I488138);
not I_28568 (I488536,I507931);
nand I_28569 (I488553,I488536,I488242);
nand I_28570 (I488570,I488488,I488553);
nand I_28571 (I488041,I488570,I488519);
nand I_28572 (I488038,I488553,I488437);
not I_28573 (I488642,I2866);
DFFARX1 I_28574 (I147787,I2859,I488642,I488668,);
and I_28575 (I488676,I488668,I147772);
DFFARX1 I_28576 (I488676,I2859,I488642,I488625,);
DFFARX1 I_28577 (I147778,I2859,I488642,I488716,);
not I_28578 (I488724,I147760);
not I_28579 (I488741,I147781);
nand I_28580 (I488758,I488741,I488724);
nor I_28581 (I488613,I488716,I488758);
DFFARX1 I_28582 (I488758,I2859,I488642,I488798,);
not I_28583 (I488634,I488798);
not I_28584 (I488820,I147784);
nand I_28585 (I488837,I488741,I488820);
DFFARX1 I_28586 (I488837,I2859,I488642,I488863,);
not I_28587 (I488871,I488863);
not I_28588 (I488888,I147775);
nand I_28589 (I488905,I488888,I147763);
and I_28590 (I488922,I488724,I488905);
nor I_28591 (I488939,I488837,I488922);
DFFARX1 I_28592 (I488939,I2859,I488642,I488610,);
DFFARX1 I_28593 (I488922,I2859,I488642,I488631,);
nor I_28594 (I488984,I147775,I147769);
nor I_28595 (I488622,I488837,I488984);
or I_28596 (I489015,I147775,I147769);
nor I_28597 (I489032,I147766,I147760);
DFFARX1 I_28598 (I489032,I2859,I488642,I489058,);
not I_28599 (I489066,I489058);
nor I_28600 (I488628,I489066,I488871);
nand I_28601 (I489097,I489066,I488716);
not I_28602 (I489114,I147766);
nand I_28603 (I489131,I489114,I488820);
nand I_28604 (I489148,I489066,I489131);
nand I_28605 (I488619,I489148,I489097);
nand I_28606 (I488616,I489131,I489015);
not I_28607 (I489220,I2866);
DFFARX1 I_28608 (I399281,I2859,I489220,I489246,);
and I_28609 (I489254,I489246,I399275);
DFFARX1 I_28610 (I489254,I2859,I489220,I489203,);
DFFARX1 I_28611 (I399293,I2859,I489220,I489294,);
not I_28612 (I489302,I399284);
not I_28613 (I489319,I399296);
nand I_28614 (I489336,I489319,I489302);
nor I_28615 (I489191,I489294,I489336);
DFFARX1 I_28616 (I489336,I2859,I489220,I489376,);
not I_28617 (I489212,I489376);
not I_28618 (I489398,I399302);
nand I_28619 (I489415,I489319,I489398);
DFFARX1 I_28620 (I489415,I2859,I489220,I489441,);
not I_28621 (I489449,I489441);
not I_28622 (I489466,I399278);
nand I_28623 (I489483,I489466,I399299);
and I_28624 (I489500,I489302,I489483);
nor I_28625 (I489517,I489415,I489500);
DFFARX1 I_28626 (I489517,I2859,I489220,I489188,);
DFFARX1 I_28627 (I489500,I2859,I489220,I489209,);
nor I_28628 (I489562,I399278,I399290);
nor I_28629 (I489200,I489415,I489562);
or I_28630 (I489593,I399278,I399290);
nor I_28631 (I489610,I399275,I399287);
DFFARX1 I_28632 (I489610,I2859,I489220,I489636,);
not I_28633 (I489644,I489636);
nor I_28634 (I489206,I489644,I489449);
nand I_28635 (I489675,I489644,I489294);
not I_28636 (I489692,I399275);
nand I_28637 (I489709,I489692,I489398);
nand I_28638 (I489726,I489644,I489709);
nand I_28639 (I489197,I489726,I489675);
nand I_28640 (I489194,I489709,I489593);
not I_28641 (I489798,I2866);
DFFARX1 I_28642 (I403803,I2859,I489798,I489824,);
and I_28643 (I489832,I489824,I403797);
DFFARX1 I_28644 (I489832,I2859,I489798,I489781,);
DFFARX1 I_28645 (I403815,I2859,I489798,I489872,);
not I_28646 (I489880,I403806);
not I_28647 (I489897,I403818);
nand I_28648 (I489914,I489897,I489880);
nor I_28649 (I489769,I489872,I489914);
DFFARX1 I_28650 (I489914,I2859,I489798,I489954,);
not I_28651 (I489790,I489954);
not I_28652 (I489976,I403824);
nand I_28653 (I489993,I489897,I489976);
DFFARX1 I_28654 (I489993,I2859,I489798,I490019,);
not I_28655 (I490027,I490019);
not I_28656 (I490044,I403800);
nand I_28657 (I490061,I490044,I403821);
and I_28658 (I490078,I489880,I490061);
nor I_28659 (I490095,I489993,I490078);
DFFARX1 I_28660 (I490095,I2859,I489798,I489766,);
DFFARX1 I_28661 (I490078,I2859,I489798,I489787,);
nor I_28662 (I490140,I403800,I403812);
nor I_28663 (I489778,I489993,I490140);
or I_28664 (I490171,I403800,I403812);
nor I_28665 (I490188,I403797,I403809);
DFFARX1 I_28666 (I490188,I2859,I489798,I490214,);
not I_28667 (I490222,I490214);
nor I_28668 (I489784,I490222,I490027);
nand I_28669 (I490253,I490222,I489872);
not I_28670 (I490270,I403797);
nand I_28671 (I490287,I490270,I489976);
nand I_28672 (I490304,I490222,I490287);
nand I_28673 (I489775,I490304,I490253);
nand I_28674 (I489772,I490287,I490171);
not I_28675 (I490376,I2866);
DFFARX1 I_28676 (I13222,I2859,I490376,I490402,);
and I_28677 (I490410,I490402,I13225);
DFFARX1 I_28678 (I490410,I2859,I490376,I490359,);
DFFARX1 I_28679 (I13225,I2859,I490376,I490450,);
not I_28680 (I490458,I13228);
not I_28681 (I490475,I13243);
nand I_28682 (I490492,I490475,I490458);
nor I_28683 (I490347,I490450,I490492);
DFFARX1 I_28684 (I490492,I2859,I490376,I490532,);
not I_28685 (I490368,I490532);
not I_28686 (I490554,I13237);
nand I_28687 (I490571,I490475,I490554);
DFFARX1 I_28688 (I490571,I2859,I490376,I490597,);
not I_28689 (I490605,I490597);
not I_28690 (I490622,I13240);
nand I_28691 (I490639,I490622,I13222);
and I_28692 (I490656,I490458,I490639);
nor I_28693 (I490673,I490571,I490656);
DFFARX1 I_28694 (I490673,I2859,I490376,I490344,);
DFFARX1 I_28695 (I490656,I2859,I490376,I490365,);
nor I_28696 (I490718,I13240,I13234);
nor I_28697 (I490356,I490571,I490718);
or I_28698 (I490749,I13240,I13234);
nor I_28699 (I490766,I13231,I13246);
DFFARX1 I_28700 (I490766,I2859,I490376,I490792,);
not I_28701 (I490800,I490792);
nor I_28702 (I490362,I490800,I490605);
nand I_28703 (I490831,I490800,I490450);
not I_28704 (I490848,I13231);
nand I_28705 (I490865,I490848,I490554);
nand I_28706 (I490882,I490800,I490865);
nand I_28707 (I490353,I490882,I490831);
nand I_28708 (I490350,I490865,I490749);
not I_28709 (I490954,I2866);
DFFARX1 I_28710 (I189784,I2859,I490954,I490980,);
and I_28711 (I490988,I490980,I189799);
DFFARX1 I_28712 (I490988,I2859,I490954,I490937,);
DFFARX1 I_28713 (I189802,I2859,I490954,I491028,);
not I_28714 (I491036,I189796);
not I_28715 (I491053,I189811);
nand I_28716 (I491070,I491053,I491036);
nor I_28717 (I490925,I491028,I491070);
DFFARX1 I_28718 (I491070,I2859,I490954,I491110,);
not I_28719 (I490946,I491110);
not I_28720 (I491132,I189787);
nand I_28721 (I491149,I491053,I491132);
DFFARX1 I_28722 (I491149,I2859,I490954,I491175,);
not I_28723 (I491183,I491175);
not I_28724 (I491200,I189790);
nand I_28725 (I491217,I491200,I189784);
and I_28726 (I491234,I491036,I491217);
nor I_28727 (I491251,I491149,I491234);
DFFARX1 I_28728 (I491251,I2859,I490954,I490922,);
DFFARX1 I_28729 (I491234,I2859,I490954,I490943,);
nor I_28730 (I491296,I189790,I189793);
nor I_28731 (I490934,I491149,I491296);
or I_28732 (I491327,I189790,I189793);
nor I_28733 (I491344,I189808,I189805);
DFFARX1 I_28734 (I491344,I2859,I490954,I491370,);
not I_28735 (I491378,I491370);
nor I_28736 (I490940,I491378,I491183);
nand I_28737 (I491409,I491378,I491028);
not I_28738 (I491426,I189808);
nand I_28739 (I491443,I491426,I491132);
nand I_28740 (I491460,I491378,I491443);
nand I_28741 (I490931,I491460,I491409);
nand I_28742 (I490928,I491443,I491327);
not I_28743 (I491532,I2866);
DFFARX1 I_28744 (I85217,I2859,I491532,I491558,);
and I_28745 (I491566,I491558,I85220);
DFFARX1 I_28746 (I491566,I2859,I491532,I491515,);
DFFARX1 I_28747 (I85220,I2859,I491532,I491606,);
not I_28748 (I491614,I85235);
not I_28749 (I491631,I85241);
nand I_28750 (I491648,I491631,I491614);
nor I_28751 (I491503,I491606,I491648);
DFFARX1 I_28752 (I491648,I2859,I491532,I491688,);
not I_28753 (I491524,I491688);
not I_28754 (I491710,I85229);
nand I_28755 (I491727,I491631,I491710);
DFFARX1 I_28756 (I491727,I2859,I491532,I491753,);
not I_28757 (I491761,I491753);
not I_28758 (I491778,I85226);
nand I_28759 (I491795,I491778,I85223);
and I_28760 (I491812,I491614,I491795);
nor I_28761 (I491829,I491727,I491812);
DFFARX1 I_28762 (I491829,I2859,I491532,I491500,);
DFFARX1 I_28763 (I491812,I2859,I491532,I491521,);
nor I_28764 (I491874,I85226,I85217);
nor I_28765 (I491512,I491727,I491874);
or I_28766 (I491905,I85226,I85217);
nor I_28767 (I491922,I85232,I85238);
DFFARX1 I_28768 (I491922,I2859,I491532,I491948,);
not I_28769 (I491956,I491948);
nor I_28770 (I491518,I491956,I491761);
nand I_28771 (I491987,I491956,I491606);
not I_28772 (I492004,I85232);
nand I_28773 (I492021,I492004,I491710);
nand I_28774 (I492038,I491956,I492021);
nand I_28775 (I491509,I492038,I491987);
nand I_28776 (I491506,I492021,I491905);
not I_28777 (I492110,I2866);
DFFARX1 I_28778 (I29056,I2859,I492110,I492136,);
and I_28779 (I492144,I492136,I29032);
DFFARX1 I_28780 (I492144,I2859,I492110,I492093,);
DFFARX1 I_28781 (I29050,I2859,I492110,I492184,);
not I_28782 (I492192,I29038);
not I_28783 (I492209,I29035);
nand I_28784 (I492226,I492209,I492192);
nor I_28785 (I492081,I492184,I492226);
DFFARX1 I_28786 (I492226,I2859,I492110,I492266,);
not I_28787 (I492102,I492266);
not I_28788 (I492288,I29044);
nand I_28789 (I492305,I492209,I492288);
DFFARX1 I_28790 (I492305,I2859,I492110,I492331,);
not I_28791 (I492339,I492331);
not I_28792 (I492356,I29035);
nand I_28793 (I492373,I492356,I29053);
and I_28794 (I492390,I492192,I492373);
nor I_28795 (I492407,I492305,I492390);
DFFARX1 I_28796 (I492407,I2859,I492110,I492078,);
DFFARX1 I_28797 (I492390,I2859,I492110,I492099,);
nor I_28798 (I492452,I29035,I29047);
nor I_28799 (I492090,I492305,I492452);
or I_28800 (I492483,I29035,I29047);
nor I_28801 (I492500,I29041,I29032);
DFFARX1 I_28802 (I492500,I2859,I492110,I492526,);
not I_28803 (I492534,I492526);
nor I_28804 (I492096,I492534,I492339);
nand I_28805 (I492565,I492534,I492184);
not I_28806 (I492582,I29041);
nand I_28807 (I492599,I492582,I492288);
nand I_28808 (I492616,I492534,I492599);
nand I_28809 (I492087,I492616,I492565);
nand I_28810 (I492084,I492599,I492483);
not I_28811 (I492688,I2866);
DFFARX1 I_28812 (I509031,I2859,I492688,I492714,);
and I_28813 (I492722,I492714,I509025);
DFFARX1 I_28814 (I492722,I2859,I492688,I492671,);
DFFARX1 I_28815 (I509010,I2859,I492688,I492762,);
not I_28816 (I492770,I509016);
not I_28817 (I492787,I509028);
nand I_28818 (I492804,I492787,I492770);
nor I_28819 (I492659,I492762,I492804);
DFFARX1 I_28820 (I492804,I2859,I492688,I492844,);
not I_28821 (I492680,I492844);
not I_28822 (I492866,I509010);
nand I_28823 (I492883,I492787,I492866);
DFFARX1 I_28824 (I492883,I2859,I492688,I492909,);
not I_28825 (I492917,I492909);
not I_28826 (I492934,I509034);
nand I_28827 (I492951,I492934,I509022);
and I_28828 (I492968,I492770,I492951);
nor I_28829 (I492985,I492883,I492968);
DFFARX1 I_28830 (I492985,I2859,I492688,I492656,);
DFFARX1 I_28831 (I492968,I2859,I492688,I492677,);
nor I_28832 (I493030,I509034,I509013);
nor I_28833 (I492668,I492883,I493030);
or I_28834 (I493061,I509034,I509013);
nor I_28835 (I493078,I509019,I509013);
DFFARX1 I_28836 (I493078,I2859,I492688,I493104,);
not I_28837 (I493112,I493104);
nor I_28838 (I492674,I493112,I492917);
nand I_28839 (I493143,I493112,I492762);
not I_28840 (I493160,I509019);
nand I_28841 (I493177,I493160,I492866);
nand I_28842 (I493194,I493112,I493177);
nand I_28843 (I492665,I493194,I493143);
nand I_28844 (I492662,I493177,I493061);
not I_28845 (I493266,I2866);
DFFARX1 I_28846 (I313457,I2859,I493266,I493292,);
and I_28847 (I493300,I493292,I313445);
DFFARX1 I_28848 (I493300,I2859,I493266,I493249,);
DFFARX1 I_28849 (I313448,I2859,I493266,I493340,);
not I_28850 (I493348,I313442);
not I_28851 (I493365,I313466);
nand I_28852 (I493382,I493365,I493348);
nor I_28853 (I493237,I493340,I493382);
DFFARX1 I_28854 (I493382,I2859,I493266,I493422,);
not I_28855 (I493258,I493422);
not I_28856 (I493444,I313454);
nand I_28857 (I493461,I493365,I493444);
DFFARX1 I_28858 (I493461,I2859,I493266,I493487,);
not I_28859 (I493495,I493487);
not I_28860 (I493512,I313463);
nand I_28861 (I493529,I493512,I313460);
and I_28862 (I493546,I493348,I493529);
nor I_28863 (I493563,I493461,I493546);
DFFARX1 I_28864 (I493563,I2859,I493266,I493234,);
DFFARX1 I_28865 (I493546,I2859,I493266,I493255,);
nor I_28866 (I493608,I313463,I313451);
nor I_28867 (I493246,I493461,I493608);
or I_28868 (I493639,I313463,I313451);
nor I_28869 (I493656,I313442,I313445);
DFFARX1 I_28870 (I493656,I2859,I493266,I493682,);
not I_28871 (I493690,I493682);
nor I_28872 (I493252,I493690,I493495);
nand I_28873 (I493721,I493690,I493340);
not I_28874 (I493738,I313442);
nand I_28875 (I493755,I493738,I493444);
nand I_28876 (I493772,I493690,I493755);
nand I_28877 (I493243,I493772,I493721);
nand I_28878 (I493240,I493755,I493639);
not I_28879 (I493844,I2866);
DFFARX1 I_28880 (I521818,I2859,I493844,I493870,);
and I_28881 (I493878,I493870,I521800);
DFFARX1 I_28882 (I493878,I2859,I493844,I493827,);
DFFARX1 I_28883 (I521809,I2859,I493844,I493918,);
not I_28884 (I493926,I521794);
not I_28885 (I493943,I521806);
nand I_28886 (I493960,I493943,I493926);
nor I_28887 (I493815,I493918,I493960);
DFFARX1 I_28888 (I493960,I2859,I493844,I494000,);
not I_28889 (I493836,I494000);
not I_28890 (I494022,I521797);
nand I_28891 (I494039,I493943,I494022);
DFFARX1 I_28892 (I494039,I2859,I493844,I494065,);
not I_28893 (I494073,I494065);
not I_28894 (I494090,I521794);
nand I_28895 (I494107,I494090,I521797);
and I_28896 (I494124,I493926,I494107);
nor I_28897 (I494141,I494039,I494124);
DFFARX1 I_28898 (I494141,I2859,I493844,I493812,);
DFFARX1 I_28899 (I494124,I2859,I493844,I493833,);
nor I_28900 (I494186,I521794,I521815);
nor I_28901 (I493824,I494039,I494186);
or I_28902 (I494217,I521794,I521815);
nor I_28903 (I494234,I521803,I521812);
DFFARX1 I_28904 (I494234,I2859,I493844,I494260,);
not I_28905 (I494268,I494260);
nor I_28906 (I493830,I494268,I494073);
nand I_28907 (I494299,I494268,I493918);
not I_28908 (I494316,I521803);
nand I_28909 (I494333,I494316,I494022);
nand I_28910 (I494350,I494268,I494333);
nand I_28911 (I493821,I494350,I494299);
nand I_28912 (I493818,I494333,I494217);
not I_28913 (I494422,I2866);
DFFARX1 I_28914 (I562417,I2859,I494422,I494448,);
and I_28915 (I494456,I494448,I562399);
DFFARX1 I_28916 (I494456,I2859,I494422,I494405,);
DFFARX1 I_28917 (I562390,I2859,I494422,I494496,);
not I_28918 (I494504,I562405);
not I_28919 (I494521,I562393);
nand I_28920 (I494538,I494521,I494504);
nor I_28921 (I494393,I494496,I494538);
DFFARX1 I_28922 (I494538,I2859,I494422,I494578,);
not I_28923 (I494414,I494578);
not I_28924 (I494600,I562402);
nand I_28925 (I494617,I494521,I494600);
DFFARX1 I_28926 (I494617,I2859,I494422,I494643,);
not I_28927 (I494651,I494643);
not I_28928 (I494668,I562411);
nand I_28929 (I494685,I494668,I562390);
and I_28930 (I494702,I494504,I494685);
nor I_28931 (I494719,I494617,I494702);
DFFARX1 I_28932 (I494719,I2859,I494422,I494390,);
DFFARX1 I_28933 (I494702,I2859,I494422,I494411,);
nor I_28934 (I494764,I562411,I562414);
nor I_28935 (I494402,I494617,I494764);
or I_28936 (I494795,I562411,I562414);
nor I_28937 (I494812,I562408,I562396);
DFFARX1 I_28938 (I494812,I2859,I494422,I494838,);
not I_28939 (I494846,I494838);
nor I_28940 (I494408,I494846,I494651);
nand I_28941 (I494877,I494846,I494496);
not I_28942 (I494894,I562408);
nand I_28943 (I494911,I494894,I494600);
nand I_28944 (I494928,I494846,I494911);
nand I_28945 (I494399,I494928,I494877);
nand I_28946 (I494396,I494911,I494795);
not I_28947 (I495000,I2866);
DFFARX1 I_28948 (I319650,I2859,I495000,I495026,);
and I_28949 (I495034,I495026,I319656);
DFFARX1 I_28950 (I495034,I2859,I495000,I494983,);
DFFARX1 I_28951 (I319662,I2859,I495000,I495074,);
not I_28952 (I495082,I319647);
not I_28953 (I495099,I319647);
nand I_28954 (I495116,I495099,I495082);
nor I_28955 (I494971,I495074,I495116);
DFFARX1 I_28956 (I495116,I2859,I495000,I495156,);
not I_28957 (I494992,I495156);
not I_28958 (I495178,I319665);
nand I_28959 (I495195,I495099,I495178);
DFFARX1 I_28960 (I495195,I2859,I495000,I495221,);
not I_28961 (I495229,I495221);
not I_28962 (I495246,I319659);
nand I_28963 (I495263,I495246,I319650);
and I_28964 (I495280,I495082,I495263);
nor I_28965 (I495297,I495195,I495280);
DFFARX1 I_28966 (I495297,I2859,I495000,I494968,);
DFFARX1 I_28967 (I495280,I2859,I495000,I494989,);
nor I_28968 (I495342,I319659,I319668);
nor I_28969 (I494980,I495195,I495342);
or I_28970 (I495373,I319659,I319668);
nor I_28971 (I495390,I319653,I319653);
DFFARX1 I_28972 (I495390,I2859,I495000,I495416,);
not I_28973 (I495424,I495416);
nor I_28974 (I494986,I495424,I495229);
nand I_28975 (I495455,I495424,I495074);
not I_28976 (I495472,I319653);
nand I_28977 (I495489,I495472,I495178);
nand I_28978 (I495506,I495424,I495489);
nand I_28979 (I494977,I495506,I495455);
nand I_28980 (I494974,I495489,I495373);
not I_28981 (I495578,I2866);
DFFARX1 I_28982 (I84622,I2859,I495578,I495604,);
and I_28983 (I495612,I495604,I84625);
DFFARX1 I_28984 (I495612,I2859,I495578,I495561,);
DFFARX1 I_28985 (I84625,I2859,I495578,I495652,);
not I_28986 (I495660,I84640);
not I_28987 (I495677,I84646);
nand I_28988 (I495694,I495677,I495660);
nor I_28989 (I495549,I495652,I495694);
DFFARX1 I_28990 (I495694,I2859,I495578,I495734,);
not I_28991 (I495570,I495734);
not I_28992 (I495756,I84634);
nand I_28993 (I495773,I495677,I495756);
DFFARX1 I_28994 (I495773,I2859,I495578,I495799,);
not I_28995 (I495807,I495799);
not I_28996 (I495824,I84631);
nand I_28997 (I495841,I495824,I84628);
and I_28998 (I495858,I495660,I495841);
nor I_28999 (I495875,I495773,I495858);
DFFARX1 I_29000 (I495875,I2859,I495578,I495546,);
DFFARX1 I_29001 (I495858,I2859,I495578,I495567,);
nor I_29002 (I495920,I84631,I84622);
nor I_29003 (I495558,I495773,I495920);
or I_29004 (I495951,I84631,I84622);
nor I_29005 (I495968,I84637,I84643);
DFFARX1 I_29006 (I495968,I2859,I495578,I495994,);
not I_29007 (I496002,I495994);
nor I_29008 (I495564,I496002,I495807);
nand I_29009 (I496033,I496002,I495652);
not I_29010 (I496050,I84637);
nand I_29011 (I496067,I496050,I495756);
nand I_29012 (I496084,I496002,I496067);
nand I_29013 (I495555,I496084,I496033);
nand I_29014 (I495552,I496067,I495951);
not I_29015 (I496156,I2866);
DFFARX1 I_29016 (I144098,I2859,I496156,I496182,);
and I_29017 (I496190,I496182,I144083);
DFFARX1 I_29018 (I496190,I2859,I496156,I496139,);
DFFARX1 I_29019 (I144089,I2859,I496156,I496230,);
not I_29020 (I496238,I144071);
not I_29021 (I496255,I144092);
nand I_29022 (I496272,I496255,I496238);
nor I_29023 (I496127,I496230,I496272);
DFFARX1 I_29024 (I496272,I2859,I496156,I496312,);
not I_29025 (I496148,I496312);
not I_29026 (I496334,I144095);
nand I_29027 (I496351,I496255,I496334);
DFFARX1 I_29028 (I496351,I2859,I496156,I496377,);
not I_29029 (I496385,I496377);
not I_29030 (I496402,I144086);
nand I_29031 (I496419,I496402,I144074);
and I_29032 (I496436,I496238,I496419);
nor I_29033 (I496453,I496351,I496436);
DFFARX1 I_29034 (I496453,I2859,I496156,I496124,);
DFFARX1 I_29035 (I496436,I2859,I496156,I496145,);
nor I_29036 (I496498,I144086,I144080);
nor I_29037 (I496136,I496351,I496498);
or I_29038 (I496529,I144086,I144080);
nor I_29039 (I496546,I144077,I144071);
DFFARX1 I_29040 (I496546,I2859,I496156,I496572,);
not I_29041 (I496580,I496572);
nor I_29042 (I496142,I496580,I496385);
nand I_29043 (I496611,I496580,I496230);
not I_29044 (I496628,I144077);
nand I_29045 (I496645,I496628,I496334);
nand I_29046 (I496662,I496580,I496645);
nand I_29047 (I496133,I496662,I496611);
nand I_29048 (I496130,I496645,I496529);
not I_29049 (I496734,I2866);
DFFARX1 I_29050 (I263749,I2859,I496734,I496760,);
and I_29051 (I496768,I496760,I263737);
DFFARX1 I_29052 (I496768,I2859,I496734,I496717,);
DFFARX1 I_29053 (I263740,I2859,I496734,I496808,);
not I_29054 (I496816,I263734);
not I_29055 (I496833,I263758);
nand I_29056 (I496850,I496833,I496816);
nor I_29057 (I496705,I496808,I496850);
DFFARX1 I_29058 (I496850,I2859,I496734,I496890,);
not I_29059 (I496726,I496890);
not I_29060 (I496912,I263746);
nand I_29061 (I496929,I496833,I496912);
DFFARX1 I_29062 (I496929,I2859,I496734,I496955,);
not I_29063 (I496963,I496955);
not I_29064 (I496980,I263755);
nand I_29065 (I496997,I496980,I263752);
and I_29066 (I497014,I496816,I496997);
nor I_29067 (I497031,I496929,I497014);
DFFARX1 I_29068 (I497031,I2859,I496734,I496702,);
DFFARX1 I_29069 (I497014,I2859,I496734,I496723,);
nor I_29070 (I497076,I263755,I263743);
nor I_29071 (I496714,I496929,I497076);
or I_29072 (I497107,I263755,I263743);
nor I_29073 (I497124,I263734,I263737);
DFFARX1 I_29074 (I497124,I2859,I496734,I497150,);
not I_29075 (I497158,I497150);
nor I_29076 (I496720,I497158,I496963);
nand I_29077 (I497189,I497158,I496808);
not I_29078 (I497206,I263734);
nand I_29079 (I497223,I497206,I496912);
nand I_29080 (I497240,I497158,I497223);
nand I_29081 (I496711,I497240,I497189);
nand I_29082 (I496708,I497223,I497107);
not I_29083 (I497312,I2866);
DFFARX1 I_29084 (I147260,I2859,I497312,I497338,);
and I_29085 (I497346,I497338,I147245);
DFFARX1 I_29086 (I497346,I2859,I497312,I497295,);
DFFARX1 I_29087 (I147251,I2859,I497312,I497386,);
not I_29088 (I497394,I147233);
not I_29089 (I497411,I147254);
nand I_29090 (I497428,I497411,I497394);
nor I_29091 (I497283,I497386,I497428);
DFFARX1 I_29092 (I497428,I2859,I497312,I497468,);
not I_29093 (I497304,I497468);
not I_29094 (I497490,I147257);
nand I_29095 (I497507,I497411,I497490);
DFFARX1 I_29096 (I497507,I2859,I497312,I497533,);
not I_29097 (I497541,I497533);
not I_29098 (I497558,I147248);
nand I_29099 (I497575,I497558,I147236);
and I_29100 (I497592,I497394,I497575);
nor I_29101 (I497609,I497507,I497592);
DFFARX1 I_29102 (I497609,I2859,I497312,I497280,);
DFFARX1 I_29103 (I497592,I2859,I497312,I497301,);
nor I_29104 (I497654,I147248,I147242);
nor I_29105 (I497292,I497507,I497654);
or I_29106 (I497685,I147248,I147242);
nor I_29107 (I497702,I147239,I147233);
DFFARX1 I_29108 (I497702,I2859,I497312,I497728,);
not I_29109 (I497736,I497728);
nor I_29110 (I497298,I497736,I497541);
nand I_29111 (I497767,I497736,I497386);
not I_29112 (I497784,I147239);
nand I_29113 (I497801,I497784,I497490);
nand I_29114 (I497818,I497736,I497801);
nand I_29115 (I497289,I497818,I497767);
nand I_29116 (I497286,I497801,I497685);
not I_29117 (I497890,I2866);
DFFARX1 I_29118 (I140409,I2859,I497890,I497916,);
and I_29119 (I497924,I497916,I140394);
DFFARX1 I_29120 (I497924,I2859,I497890,I497873,);
DFFARX1 I_29121 (I140400,I2859,I497890,I497964,);
not I_29122 (I497972,I140382);
not I_29123 (I497989,I140403);
nand I_29124 (I498006,I497989,I497972);
nor I_29125 (I497861,I497964,I498006);
DFFARX1 I_29126 (I498006,I2859,I497890,I498046,);
not I_29127 (I497882,I498046);
not I_29128 (I498068,I140406);
nand I_29129 (I498085,I497989,I498068);
DFFARX1 I_29130 (I498085,I2859,I497890,I498111,);
not I_29131 (I498119,I498111);
not I_29132 (I498136,I140397);
nand I_29133 (I498153,I498136,I140385);
and I_29134 (I498170,I497972,I498153);
nor I_29135 (I498187,I498085,I498170);
DFFARX1 I_29136 (I498187,I2859,I497890,I497858,);
DFFARX1 I_29137 (I498170,I2859,I497890,I497879,);
nor I_29138 (I498232,I140397,I140391);
nor I_29139 (I497870,I498085,I498232);
or I_29140 (I498263,I140397,I140391);
nor I_29141 (I498280,I140388,I140382);
DFFARX1 I_29142 (I498280,I2859,I497890,I498306,);
not I_29143 (I498314,I498306);
nor I_29144 (I497876,I498314,I498119);
nand I_29145 (I498345,I498314,I497964);
not I_29146 (I498362,I140388);
nand I_29147 (I498379,I498362,I498068);
nand I_29148 (I498396,I498314,I498379);
nand I_29149 (I497867,I498396,I498345);
nand I_29150 (I497864,I498379,I498263);
not I_29151 (I498468,I2866);
DFFARX1 I_29152 (I510663,I2859,I498468,I498494,);
and I_29153 (I498502,I498494,I510657);
DFFARX1 I_29154 (I498502,I2859,I498468,I498451,);
DFFARX1 I_29155 (I510642,I2859,I498468,I498542,);
not I_29156 (I498550,I510648);
not I_29157 (I498567,I510660);
nand I_29158 (I498584,I498567,I498550);
nor I_29159 (I498439,I498542,I498584);
DFFARX1 I_29160 (I498584,I2859,I498468,I498624,);
not I_29161 (I498460,I498624);
not I_29162 (I498646,I510642);
nand I_29163 (I498663,I498567,I498646);
DFFARX1 I_29164 (I498663,I2859,I498468,I498689,);
not I_29165 (I498697,I498689);
not I_29166 (I498714,I510666);
nand I_29167 (I498731,I498714,I510654);
and I_29168 (I498748,I498550,I498731);
nor I_29169 (I498765,I498663,I498748);
DFFARX1 I_29170 (I498765,I2859,I498468,I498436,);
DFFARX1 I_29171 (I498748,I2859,I498468,I498457,);
nor I_29172 (I498810,I510666,I510645);
nor I_29173 (I498448,I498663,I498810);
or I_29174 (I498841,I510666,I510645);
nor I_29175 (I498858,I510651,I510645);
DFFARX1 I_29176 (I498858,I2859,I498468,I498884,);
not I_29177 (I498892,I498884);
nor I_29178 (I498454,I498892,I498697);
nand I_29179 (I498923,I498892,I498542);
not I_29180 (I498940,I510651);
nand I_29181 (I498957,I498940,I498646);
nand I_29182 (I498974,I498892,I498957);
nand I_29183 (I498445,I498974,I498923);
nand I_29184 (I498442,I498957,I498841);
not I_29185 (I499046,I2866);
DFFARX1 I_29186 (I281089,I2859,I499046,I499072,);
and I_29187 (I499080,I499072,I281077);
DFFARX1 I_29188 (I499080,I2859,I499046,I499029,);
DFFARX1 I_29189 (I281080,I2859,I499046,I499120,);
not I_29190 (I499128,I281074);
not I_29191 (I499145,I281098);
nand I_29192 (I499162,I499145,I499128);
nor I_29193 (I499017,I499120,I499162);
DFFARX1 I_29194 (I499162,I2859,I499046,I499202,);
not I_29195 (I499038,I499202);
not I_29196 (I499224,I281086);
nand I_29197 (I499241,I499145,I499224);
DFFARX1 I_29198 (I499241,I2859,I499046,I499267,);
not I_29199 (I499275,I499267);
not I_29200 (I499292,I281095);
nand I_29201 (I499309,I499292,I281092);
and I_29202 (I499326,I499128,I499309);
nor I_29203 (I499343,I499241,I499326);
DFFARX1 I_29204 (I499343,I2859,I499046,I499014,);
DFFARX1 I_29205 (I499326,I2859,I499046,I499035,);
nor I_29206 (I499388,I281095,I281083);
nor I_29207 (I499026,I499241,I499388);
or I_29208 (I499419,I281095,I281083);
nor I_29209 (I499436,I281074,I281077);
DFFARX1 I_29210 (I499436,I2859,I499046,I499462,);
not I_29211 (I499470,I499462);
nor I_29212 (I499032,I499470,I499275);
nand I_29213 (I499501,I499470,I499120);
not I_29214 (I499518,I281074);
nand I_29215 (I499535,I499518,I499224);
nand I_29216 (I499552,I499470,I499535);
nand I_29217 (I499023,I499552,I499501);
nand I_29218 (I499020,I499535,I499419);
not I_29219 (I499624,I2866);
DFFARX1 I_29220 (I50707,I2859,I499624,I499650,);
and I_29221 (I499658,I499650,I50731);
DFFARX1 I_29222 (I499658,I2859,I499624,I499607,);
DFFARX1 I_29223 (I50707,I2859,I499624,I499698,);
not I_29224 (I499706,I50725);
not I_29225 (I499723,I50710);
nand I_29226 (I499740,I499723,I499706);
nor I_29227 (I499595,I499698,I499740);
DFFARX1 I_29228 (I499740,I2859,I499624,I499780,);
not I_29229 (I499616,I499780);
not I_29230 (I499802,I50719);
nand I_29231 (I499819,I499723,I499802);
DFFARX1 I_29232 (I499819,I2859,I499624,I499845,);
not I_29233 (I499853,I499845);
not I_29234 (I499870,I50716);
nand I_29235 (I499887,I499870,I50713);
and I_29236 (I499904,I499706,I499887);
nor I_29237 (I499921,I499819,I499904);
DFFARX1 I_29238 (I499921,I2859,I499624,I499592,);
DFFARX1 I_29239 (I499904,I2859,I499624,I499613,);
nor I_29240 (I499966,I50716,I50722);
nor I_29241 (I499604,I499819,I499966);
or I_29242 (I499997,I50716,I50722);
nor I_29243 (I500014,I50728,I50734);
DFFARX1 I_29244 (I500014,I2859,I499624,I500040,);
not I_29245 (I500048,I500040);
nor I_29246 (I499610,I500048,I499853);
nand I_29247 (I500079,I500048,I499698);
not I_29248 (I500096,I50728);
nand I_29249 (I500113,I500096,I499802);
nand I_29250 (I500130,I500048,I500113);
nand I_29251 (I499601,I500130,I500079);
nand I_29252 (I499598,I500113,I499997);
not I_29253 (I500202,I2866);
DFFARX1 I_29254 (I2356,I2859,I500202,I500228,);
and I_29255 (I500236,I500228,I1604);
DFFARX1 I_29256 (I500236,I2859,I500202,I500185,);
DFFARX1 I_29257 (I2516,I2859,I500202,I500276,);
not I_29258 (I500284,I2124);
not I_29259 (I500301,I1436);
nand I_29260 (I500318,I500301,I500284);
nor I_29261 (I500173,I500276,I500318);
DFFARX1 I_29262 (I500318,I2859,I500202,I500358,);
not I_29263 (I500194,I500358);
not I_29264 (I500380,I2444);
nand I_29265 (I500397,I500301,I500380);
DFFARX1 I_29266 (I500397,I2859,I500202,I500423,);
not I_29267 (I500431,I500423);
not I_29268 (I500448,I2420);
nand I_29269 (I500465,I500448,I1780);
and I_29270 (I500482,I500284,I500465);
nor I_29271 (I500499,I500397,I500482);
DFFARX1 I_29272 (I500499,I2859,I500202,I500170,);
DFFARX1 I_29273 (I500482,I2859,I500202,I500191,);
nor I_29274 (I500544,I2420,I1572);
nor I_29275 (I500182,I500397,I500544);
or I_29276 (I500575,I2420,I1572);
nor I_29277 (I500592,I2732,I1532);
DFFARX1 I_29278 (I500592,I2859,I500202,I500618,);
not I_29279 (I500626,I500618);
nor I_29280 (I500188,I500626,I500431);
nand I_29281 (I500657,I500626,I500276);
not I_29282 (I500674,I2732);
nand I_29283 (I500691,I500674,I500380);
nand I_29284 (I500708,I500626,I500691);
nand I_29285 (I500179,I500708,I500657);
nand I_29286 (I500176,I500691,I500575);
not I_29287 (I500780,I2866);
DFFARX1 I_29288 (I399927,I2859,I500780,I500806,);
and I_29289 (I500814,I500806,I399921);
DFFARX1 I_29290 (I500814,I2859,I500780,I500763,);
DFFARX1 I_29291 (I399939,I2859,I500780,I500854,);
not I_29292 (I500862,I399930);
not I_29293 (I500879,I399942);
nand I_29294 (I500896,I500879,I500862);
nor I_29295 (I500751,I500854,I500896);
DFFARX1 I_29296 (I500896,I2859,I500780,I500936,);
not I_29297 (I500772,I500936);
not I_29298 (I500958,I399948);
nand I_29299 (I500975,I500879,I500958);
DFFARX1 I_29300 (I500975,I2859,I500780,I501001,);
not I_29301 (I501009,I501001);
not I_29302 (I501026,I399924);
nand I_29303 (I501043,I501026,I399945);
and I_29304 (I501060,I500862,I501043);
nor I_29305 (I501077,I500975,I501060);
DFFARX1 I_29306 (I501077,I2859,I500780,I500748,);
DFFARX1 I_29307 (I501060,I2859,I500780,I500769,);
nor I_29308 (I501122,I399924,I399936);
nor I_29309 (I500760,I500975,I501122);
or I_29310 (I501153,I399924,I399936);
nor I_29311 (I501170,I399921,I399933);
DFFARX1 I_29312 (I501170,I2859,I500780,I501196,);
not I_29313 (I501204,I501196);
nor I_29314 (I500766,I501204,I501009);
nand I_29315 (I501235,I501204,I500854);
not I_29316 (I501252,I399921);
nand I_29317 (I501269,I501252,I500958);
nand I_29318 (I501286,I501204,I501269);
nand I_29319 (I500757,I501286,I501235);
nand I_29320 (I500754,I501269,I501153);
not I_29321 (I501358,I2866);
DFFARX1 I_29322 (I133558,I2859,I501358,I501384,);
and I_29323 (I501392,I501384,I133543);
DFFARX1 I_29324 (I501392,I2859,I501358,I501341,);
DFFARX1 I_29325 (I133549,I2859,I501358,I501432,);
not I_29326 (I501440,I133531);
not I_29327 (I501457,I133552);
nand I_29328 (I501474,I501457,I501440);
nor I_29329 (I501329,I501432,I501474);
DFFARX1 I_29330 (I501474,I2859,I501358,I501514,);
not I_29331 (I501350,I501514);
not I_29332 (I501536,I133555);
nand I_29333 (I501553,I501457,I501536);
DFFARX1 I_29334 (I501553,I2859,I501358,I501579,);
not I_29335 (I501587,I501579);
not I_29336 (I501604,I133546);
nand I_29337 (I501621,I501604,I133534);
and I_29338 (I501638,I501440,I501621);
nor I_29339 (I501655,I501553,I501638);
DFFARX1 I_29340 (I501655,I2859,I501358,I501326,);
DFFARX1 I_29341 (I501638,I2859,I501358,I501347,);
nor I_29342 (I501700,I133546,I133540);
nor I_29343 (I501338,I501553,I501700);
or I_29344 (I501731,I133546,I133540);
nor I_29345 (I501748,I133537,I133531);
DFFARX1 I_29346 (I501748,I2859,I501358,I501774,);
not I_29347 (I501782,I501774);
nor I_29348 (I501344,I501782,I501587);
nand I_29349 (I501813,I501782,I501432);
not I_29350 (I501830,I133537);
nand I_29351 (I501847,I501830,I501536);
nand I_29352 (I501864,I501782,I501847);
nand I_29353 (I501335,I501864,I501813);
nand I_29354 (I501332,I501847,I501731);
not I_29355 (I501936,I2866);
DFFARX1 I_29356 (I70342,I2859,I501936,I501962,);
and I_29357 (I501970,I501962,I70345);
DFFARX1 I_29358 (I501970,I2859,I501936,I501919,);
DFFARX1 I_29359 (I70345,I2859,I501936,I502010,);
not I_29360 (I502018,I70360);
not I_29361 (I502035,I70366);
nand I_29362 (I502052,I502035,I502018);
nor I_29363 (I501907,I502010,I502052);
DFFARX1 I_29364 (I502052,I2859,I501936,I502092,);
not I_29365 (I501928,I502092);
not I_29366 (I502114,I70354);
nand I_29367 (I502131,I502035,I502114);
DFFARX1 I_29368 (I502131,I2859,I501936,I502157,);
not I_29369 (I502165,I502157);
not I_29370 (I502182,I70351);
nand I_29371 (I502199,I502182,I70348);
and I_29372 (I502216,I502018,I502199);
nor I_29373 (I502233,I502131,I502216);
DFFARX1 I_29374 (I502233,I2859,I501936,I501904,);
DFFARX1 I_29375 (I502216,I2859,I501936,I501925,);
nor I_29376 (I502278,I70351,I70342);
nor I_29377 (I501916,I502131,I502278);
or I_29378 (I502309,I70351,I70342);
nor I_29379 (I502326,I70357,I70363);
DFFARX1 I_29380 (I502326,I2859,I501936,I502352,);
not I_29381 (I502360,I502352);
nor I_29382 (I501922,I502360,I502165);
nand I_29383 (I502391,I502360,I502010);
not I_29384 (I502408,I70357);
nand I_29385 (I502425,I502408,I502114);
nand I_29386 (I502442,I502360,I502425);
nand I_29387 (I501913,I502442,I502391);
nand I_29388 (I501910,I502425,I502309);
not I_29389 (I502514,I2866);
DFFARX1 I_29390 (I120368,I2859,I502514,I502540,);
nand I_29391 (I502548,I502540,I120371);
DFFARX1 I_29392 (I120365,I2859,I502514,I502574,);
DFFARX1 I_29393 (I502574,I2859,I502514,I502591,);
not I_29394 (I502506,I502591);
not I_29395 (I502613,I120374);
nor I_29396 (I502630,I120374,I120359);
not I_29397 (I502647,I120383);
nand I_29398 (I502664,I502613,I502647);
nor I_29399 (I502681,I120383,I120374);
and I_29400 (I502485,I502681,I502548);
not I_29401 (I502712,I120362);
nand I_29402 (I502729,I502712,I120380);
nor I_29403 (I502746,I120362,I120356);
not I_29404 (I502763,I502746);
nand I_29405 (I502488,I502630,I502763);
DFFARX1 I_29406 (I502746,I2859,I502514,I502503,);
nor I_29407 (I502808,I120377,I120383);
nor I_29408 (I502825,I502808,I120359);
and I_29409 (I502842,I502825,I502729);
DFFARX1 I_29410 (I502842,I2859,I502514,I502500,);
nor I_29411 (I502497,I502808,I502664);
or I_29412 (I502494,I502746,I502808);
nor I_29413 (I502901,I120377,I120356);
DFFARX1 I_29414 (I502901,I2859,I502514,I502927,);
not I_29415 (I502935,I502927);
nand I_29416 (I502952,I502935,I502613);
nor I_29417 (I502969,I502952,I120359);
DFFARX1 I_29418 (I502969,I2859,I502514,I502482,);
nor I_29419 (I503000,I502935,I502664);
nor I_29420 (I502491,I502808,I503000);
not I_29421 (I503058,I2866);
DFFARX1 I_29422 (I531051,I2859,I503058,I503084,);
nand I_29423 (I503092,I503084,I531060);
DFFARX1 I_29424 (I531063,I2859,I503058,I503118,);
DFFARX1 I_29425 (I503118,I2859,I503058,I503135,);
not I_29426 (I503050,I503135);
not I_29427 (I503157,I531057);
nor I_29428 (I503174,I531057,I531054);
not I_29429 (I503191,I531048);
nand I_29430 (I503208,I503157,I503191);
nor I_29431 (I503225,I531048,I531057);
and I_29432 (I503029,I503225,I503092);
not I_29433 (I503256,I531045);
nand I_29434 (I503273,I503256,I531042);
nor I_29435 (I503290,I531045,I531042);
not I_29436 (I503307,I503290);
nand I_29437 (I503032,I503174,I503307);
DFFARX1 I_29438 (I503290,I2859,I503058,I503047,);
nor I_29439 (I503352,I531045,I531048);
nor I_29440 (I503369,I503352,I531054);
and I_29441 (I503386,I503369,I503273);
DFFARX1 I_29442 (I503386,I2859,I503058,I503044,);
nor I_29443 (I503041,I503352,I503208);
or I_29444 (I503038,I503290,I503352);
nor I_29445 (I503445,I531045,I531066);
DFFARX1 I_29446 (I503445,I2859,I503058,I503471,);
not I_29447 (I503479,I503471);
nand I_29448 (I503496,I503479,I503157);
nor I_29449 (I503513,I503496,I531054);
DFFARX1 I_29450 (I503513,I2859,I503058,I503026,);
nor I_29451 (I503544,I503479,I503208);
nor I_29452 (I503035,I503352,I503544);
not I_29453 (I503602,I2866);
DFFARX1 I_29454 (I477074,I2859,I503602,I503628,);
nand I_29455 (I503636,I503628,I477053);
DFFARX1 I_29456 (I477050,I2859,I503602,I503662,);
DFFARX1 I_29457 (I503662,I2859,I503602,I503679,);
not I_29458 (I503594,I503679);
not I_29459 (I503701,I477062);
nor I_29460 (I503718,I477062,I477071);
not I_29461 (I503735,I477059);
nand I_29462 (I503752,I503701,I503735);
nor I_29463 (I503769,I477059,I477062);
and I_29464 (I503573,I503769,I503636);
not I_29465 (I503800,I477068);
nand I_29466 (I503817,I503800,I477065);
nor I_29467 (I503834,I477068,I477050);
not I_29468 (I503851,I503834);
nand I_29469 (I503576,I503718,I503851);
DFFARX1 I_29470 (I503834,I2859,I503602,I503591,);
nor I_29471 (I503896,I477053,I477059);
nor I_29472 (I503913,I503896,I477071);
and I_29473 (I503930,I503913,I503817);
DFFARX1 I_29474 (I503930,I2859,I503602,I503588,);
nor I_29475 (I503585,I503896,I503752);
or I_29476 (I503582,I503834,I503896);
nor I_29477 (I503989,I477053,I477056);
DFFARX1 I_29478 (I503989,I2859,I503602,I504015,);
not I_29479 (I504023,I504015);
nand I_29480 (I504040,I504023,I503701);
nor I_29481 (I504057,I504040,I477071);
DFFARX1 I_29482 (I504057,I2859,I503602,I503570,);
nor I_29483 (I504088,I504023,I503752);
nor I_29484 (I503579,I503896,I504088);
not I_29485 (I504146,I2866);
DFFARX1 I_29486 (I557657,I2859,I504146,I504172,);
nand I_29487 (I504180,I504172,I557642);
DFFARX1 I_29488 (I557636,I2859,I504146,I504206,);
DFFARX1 I_29489 (I504206,I2859,I504146,I504223,);
not I_29490 (I504138,I504223);
not I_29491 (I504245,I557630);
nor I_29492 (I504262,I557630,I557651);
not I_29493 (I504279,I557639);
nand I_29494 (I504296,I504245,I504279);
nor I_29495 (I504313,I557639,I557630);
and I_29496 (I504117,I504313,I504180);
not I_29497 (I504344,I557648);
nand I_29498 (I504361,I504344,I557654);
nor I_29499 (I504378,I557648,I557645);
not I_29500 (I504395,I504378);
nand I_29501 (I504120,I504262,I504395);
DFFARX1 I_29502 (I504378,I2859,I504146,I504135,);
nor I_29503 (I504440,I557633,I557639);
nor I_29504 (I504457,I504440,I557651);
and I_29505 (I504474,I504457,I504361);
DFFARX1 I_29506 (I504474,I2859,I504146,I504132,);
nor I_29507 (I504129,I504440,I504296);
or I_29508 (I504126,I504378,I504440);
nor I_29509 (I504533,I557633,I557630);
DFFARX1 I_29510 (I504533,I2859,I504146,I504559,);
not I_29511 (I504567,I504559);
nand I_29512 (I504584,I504567,I504245);
nor I_29513 (I504601,I504584,I557651);
DFFARX1 I_29514 (I504601,I2859,I504146,I504114,);
nor I_29515 (I504632,I504567,I504296);
nor I_29516 (I504123,I504440,I504632);
not I_29517 (I504690,I2866);
DFFARX1 I_29518 (I259691,I2859,I504690,I504716,);
nand I_29519 (I504724,I504716,I259706);
DFFARX1 I_29520 (I259700,I2859,I504690,I504750,);
DFFARX1 I_29521 (I504750,I2859,I504690,I504767,);
not I_29522 (I504682,I504767);
not I_29523 (I504789,I259703);
nor I_29524 (I504806,I259703,I259709);
not I_29525 (I504823,I259691);
nand I_29526 (I504840,I504789,I504823);
nor I_29527 (I504857,I259691,I259703);
and I_29528 (I504661,I504857,I504724);
not I_29529 (I504888,I259688);
nand I_29530 (I504905,I504888,I259694);
nor I_29531 (I504922,I259688,I259688);
not I_29532 (I504939,I504922);
nand I_29533 (I504664,I504806,I504939);
DFFARX1 I_29534 (I504922,I2859,I504690,I504679,);
nor I_29535 (I504984,I259697,I259691);
nor I_29536 (I505001,I504984,I259709);
and I_29537 (I505018,I505001,I504905);
DFFARX1 I_29538 (I505018,I2859,I504690,I504676,);
nor I_29539 (I504673,I504984,I504840);
or I_29540 (I504670,I504922,I504984);
nor I_29541 (I505077,I259697,I259712);
DFFARX1 I_29542 (I505077,I2859,I504690,I505103,);
not I_29543 (I505111,I505103);
nand I_29544 (I505128,I505111,I504789);
nor I_29545 (I505145,I505128,I259709);
DFFARX1 I_29546 (I505145,I2859,I504690,I504658,);
nor I_29547 (I505176,I505111,I504840);
nor I_29548 (I504667,I504984,I505176);
not I_29549 (I505234,I2866);
DFFARX1 I_29550 (I67376,I2859,I505234,I505260,);
nand I_29551 (I505268,I505260,I67391);
DFFARX1 I_29552 (I67388,I2859,I505234,I505294,);
DFFARX1 I_29553 (I505294,I2859,I505234,I505311,);
not I_29554 (I505226,I505311);
not I_29555 (I505333,I67367);
nor I_29556 (I505350,I67367,I67373);
not I_29557 (I505367,I67379);
nand I_29558 (I505384,I505333,I505367);
nor I_29559 (I505401,I67379,I67367);
and I_29560 (I505205,I505401,I505268);
not I_29561 (I505432,I67385);
nand I_29562 (I505449,I505432,I67367);
nor I_29563 (I505466,I67385,I67370);
not I_29564 (I505483,I505466);
nand I_29565 (I505208,I505350,I505483);
DFFARX1 I_29566 (I505466,I2859,I505234,I505223,);
nor I_29567 (I505528,I67370,I67379);
nor I_29568 (I505545,I505528,I67373);
and I_29569 (I505562,I505545,I505449);
DFFARX1 I_29570 (I505562,I2859,I505234,I505220,);
nor I_29571 (I505217,I505528,I505384);
or I_29572 (I505214,I505466,I505528);
nor I_29573 (I505621,I67370,I67382);
DFFARX1 I_29574 (I505621,I2859,I505234,I505647,);
not I_29575 (I505655,I505647);
nand I_29576 (I505672,I505655,I505333);
nor I_29577 (I505689,I505672,I67373);
DFFARX1 I_29578 (I505689,I2859,I505234,I505202,);
nor I_29579 (I505720,I505655,I505384);
nor I_29580 (I505211,I505528,I505720);
not I_29581 (I505778,I2866);
DFFARX1 I_29582 (I540997,I2859,I505778,I505804,);
nand I_29583 (I505812,I505804,I540982);
DFFARX1 I_29584 (I540976,I2859,I505778,I505838,);
DFFARX1 I_29585 (I505838,I2859,I505778,I505855,);
not I_29586 (I505770,I505855);
not I_29587 (I505877,I540970);
nor I_29588 (I505894,I540970,I540991);
not I_29589 (I505911,I540979);
nand I_29590 (I505928,I505877,I505911);
nor I_29591 (I505945,I540979,I540970);
and I_29592 (I505749,I505945,I505812);
not I_29593 (I505976,I540988);
nand I_29594 (I505993,I505976,I540994);
nor I_29595 (I506010,I540988,I540985);
not I_29596 (I506027,I506010);
nand I_29597 (I505752,I505894,I506027);
DFFARX1 I_29598 (I506010,I2859,I505778,I505767,);
nor I_29599 (I506072,I540973,I540979);
nor I_29600 (I506089,I506072,I540991);
and I_29601 (I506106,I506089,I505993);
DFFARX1 I_29602 (I506106,I2859,I505778,I505764,);
nor I_29603 (I505761,I506072,I505928);
or I_29604 (I505758,I506010,I506072);
nor I_29605 (I506165,I540973,I540970);
DFFARX1 I_29606 (I506165,I2859,I505778,I506191,);
not I_29607 (I506199,I506191);
nand I_29608 (I506216,I506199,I505877);
nor I_29609 (I506233,I506216,I540991);
DFFARX1 I_29610 (I506233,I2859,I505778,I505746,);
nor I_29611 (I506264,I506199,I505928);
nor I_29612 (I505755,I506072,I506264);
not I_29613 (I506322,I2866);
DFFARX1 I_29614 (I573722,I2859,I506322,I506348,);
nand I_29615 (I506356,I506348,I573707);
DFFARX1 I_29616 (I573701,I2859,I506322,I506382,);
DFFARX1 I_29617 (I506382,I2859,I506322,I506399,);
not I_29618 (I506314,I506399);
not I_29619 (I506421,I573695);
nor I_29620 (I506438,I573695,I573716);
not I_29621 (I506455,I573704);
nand I_29622 (I506472,I506421,I506455);
nor I_29623 (I506489,I573704,I573695);
and I_29624 (I506293,I506489,I506356);
not I_29625 (I506520,I573713);
nand I_29626 (I506537,I506520,I573719);
nor I_29627 (I506554,I573713,I573710);
not I_29628 (I506571,I506554);
nand I_29629 (I506296,I506438,I506571);
DFFARX1 I_29630 (I506554,I2859,I506322,I506311,);
nor I_29631 (I506616,I573698,I573704);
nor I_29632 (I506633,I506616,I573716);
and I_29633 (I506650,I506633,I506537);
DFFARX1 I_29634 (I506650,I2859,I506322,I506308,);
nor I_29635 (I506305,I506616,I506472);
or I_29636 (I506302,I506554,I506616);
nor I_29637 (I506709,I573698,I573695);
DFFARX1 I_29638 (I506709,I2859,I506322,I506735,);
not I_29639 (I506743,I506735);
nand I_29640 (I506760,I506743,I506421);
nor I_29641 (I506777,I506760,I573716);
DFFARX1 I_29642 (I506777,I2859,I506322,I506290,);
nor I_29643 (I506808,I506743,I506472);
nor I_29644 (I506299,I506616,I506808);
not I_29645 (I506866,I2866);
DFFARX1 I_29646 (I539212,I2859,I506866,I506892,);
nand I_29647 (I506900,I506892,I539197);
DFFARX1 I_29648 (I539191,I2859,I506866,I506926,);
DFFARX1 I_29649 (I506926,I2859,I506866,I506943,);
not I_29650 (I506858,I506943);
not I_29651 (I506965,I539185);
nor I_29652 (I506982,I539185,I539206);
not I_29653 (I506999,I539194);
nand I_29654 (I507016,I506965,I506999);
nor I_29655 (I507033,I539194,I539185);
and I_29656 (I506837,I507033,I506900);
not I_29657 (I507064,I539203);
nand I_29658 (I507081,I507064,I539209);
nor I_29659 (I507098,I539203,I539200);
not I_29660 (I507115,I507098);
nand I_29661 (I506840,I506982,I507115);
DFFARX1 I_29662 (I507098,I2859,I506866,I506855,);
nor I_29663 (I507160,I539188,I539194);
nor I_29664 (I507177,I507160,I539206);
and I_29665 (I507194,I507177,I507081);
DFFARX1 I_29666 (I507194,I2859,I506866,I506852,);
nor I_29667 (I506849,I507160,I507016);
or I_29668 (I506846,I507098,I507160);
nor I_29669 (I507253,I539188,I539185);
DFFARX1 I_29670 (I507253,I2859,I506866,I507279,);
not I_29671 (I507287,I507279);
nand I_29672 (I507304,I507287,I506965);
nor I_29673 (I507321,I507304,I539206);
DFFARX1 I_29674 (I507321,I2859,I506866,I506834,);
nor I_29675 (I507352,I507287,I507016);
nor I_29676 (I506843,I507160,I507352);
not I_29677 (I507410,I2866);
DFFARX1 I_29678 (I343368,I2859,I507410,I507436,);
nand I_29679 (I507444,I507436,I343362);
DFFARX1 I_29680 (I343365,I2859,I507410,I507470,);
DFFARX1 I_29681 (I507470,I2859,I507410,I507487,);
not I_29682 (I507402,I507487);
not I_29683 (I507509,I343371);
nor I_29684 (I507526,I343371,I343365);
not I_29685 (I507543,I343374);
nand I_29686 (I507560,I507509,I507543);
nor I_29687 (I507577,I343374,I343371);
and I_29688 (I507381,I507577,I507444);
not I_29689 (I507608,I343383);
nand I_29690 (I507625,I507608,I343377);
nor I_29691 (I507642,I343383,I343380);
not I_29692 (I507659,I507642);
nand I_29693 (I507384,I507526,I507659);
DFFARX1 I_29694 (I507642,I2859,I507410,I507399,);
nor I_29695 (I507704,I343362,I343374);
nor I_29696 (I507721,I507704,I343365);
and I_29697 (I507738,I507721,I507625);
DFFARX1 I_29698 (I507738,I2859,I507410,I507396,);
nor I_29699 (I507393,I507704,I507560);
or I_29700 (I507390,I507642,I507704);
nor I_29701 (I507797,I343362,I343368);
DFFARX1 I_29702 (I507797,I2859,I507410,I507823,);
not I_29703 (I507831,I507823);
nand I_29704 (I507848,I507831,I507509);
nor I_29705 (I507865,I507848,I343365);
DFFARX1 I_29706 (I507865,I2859,I507410,I507378,);
nor I_29707 (I507896,I507831,I507560);
nor I_29708 (I507387,I507704,I507896);
not I_29709 (I507954,I2866);
DFFARX1 I_29710 (I169136,I2859,I507954,I507980,);
nand I_29711 (I507988,I507980,I169133);
DFFARX1 I_29712 (I169112,I2859,I507954,I508014,);
DFFARX1 I_29713 (I508014,I2859,I507954,I508031,);
not I_29714 (I507946,I508031);
not I_29715 (I508053,I169127);
nor I_29716 (I508070,I169127,I169130);
not I_29717 (I508087,I169121);
nand I_29718 (I508104,I508053,I508087);
nor I_29719 (I508121,I169121,I169127);
and I_29720 (I507925,I508121,I507988);
not I_29721 (I508152,I169118);
nand I_29722 (I508169,I508152,I169139);
nor I_29723 (I508186,I169118,I169115);
not I_29724 (I508203,I508186);
nand I_29725 (I507928,I508070,I508203);
DFFARX1 I_29726 (I508186,I2859,I507954,I507943,);
nor I_29727 (I508248,I169124,I169121);
nor I_29728 (I508265,I508248,I169130);
and I_29729 (I508282,I508265,I508169);
DFFARX1 I_29730 (I508282,I2859,I507954,I507940,);
nor I_29731 (I507937,I508248,I508104);
or I_29732 (I507934,I508186,I508248);
nor I_29733 (I508341,I169124,I169112);
DFFARX1 I_29734 (I508341,I2859,I507954,I508367,);
not I_29735 (I508375,I508367);
nand I_29736 (I508392,I508375,I508053);
nor I_29737 (I508409,I508392,I169130);
DFFARX1 I_29738 (I508409,I2859,I507954,I507922,);
nor I_29739 (I508440,I508375,I508104);
nor I_29740 (I507931,I508248,I508440);
not I_29741 (I508498,I2866);
DFFARX1 I_29742 (I295527,I2859,I508498,I508524,);
nand I_29743 (I508532,I508524,I295542);
DFFARX1 I_29744 (I295536,I2859,I508498,I508558,);
DFFARX1 I_29745 (I508558,I2859,I508498,I508575,);
not I_29746 (I508490,I508575);
not I_29747 (I508597,I295539);
nor I_29748 (I508614,I295539,I295545);
not I_29749 (I508631,I295527);
nand I_29750 (I508648,I508597,I508631);
nor I_29751 (I508665,I295527,I295539);
and I_29752 (I508469,I508665,I508532);
not I_29753 (I508696,I295524);
nand I_29754 (I508713,I508696,I295530);
nor I_29755 (I508730,I295524,I295524);
not I_29756 (I508747,I508730);
nand I_29757 (I508472,I508614,I508747);
DFFARX1 I_29758 (I508730,I2859,I508498,I508487,);
nor I_29759 (I508792,I295533,I295527);
nor I_29760 (I508809,I508792,I295545);
and I_29761 (I508826,I508809,I508713);
DFFARX1 I_29762 (I508826,I2859,I508498,I508484,);
nor I_29763 (I508481,I508792,I508648);
or I_29764 (I508478,I508730,I508792);
nor I_29765 (I508885,I295533,I295548);
DFFARX1 I_29766 (I508885,I2859,I508498,I508911,);
not I_29767 (I508919,I508911);
nand I_29768 (I508936,I508919,I508597);
nor I_29769 (I508953,I508936,I295545);
DFFARX1 I_29770 (I508953,I2859,I508498,I508466,);
nor I_29771 (I508984,I508919,I508648);
nor I_29772 (I508475,I508792,I508984);
not I_29773 (I509042,I2866);
DFFARX1 I_29774 (I268939,I2859,I509042,I509068,);
nand I_29775 (I509076,I509068,I268954);
DFFARX1 I_29776 (I268948,I2859,I509042,I509102,);
DFFARX1 I_29777 (I509102,I2859,I509042,I509119,);
not I_29778 (I509034,I509119);
not I_29779 (I509141,I268951);
nor I_29780 (I509158,I268951,I268957);
not I_29781 (I509175,I268939);
nand I_29782 (I509192,I509141,I509175);
nor I_29783 (I509209,I268939,I268951);
and I_29784 (I509013,I509209,I509076);
not I_29785 (I509240,I268936);
nand I_29786 (I509257,I509240,I268942);
nor I_29787 (I509274,I268936,I268936);
not I_29788 (I509291,I509274);
nand I_29789 (I509016,I509158,I509291);
DFFARX1 I_29790 (I509274,I2859,I509042,I509031,);
nor I_29791 (I509336,I268945,I268939);
nor I_29792 (I509353,I509336,I268957);
and I_29793 (I509370,I509353,I509257);
DFFARX1 I_29794 (I509370,I2859,I509042,I509028,);
nor I_29795 (I509025,I509336,I509192);
or I_29796 (I509022,I509274,I509336);
nor I_29797 (I509429,I268945,I268960);
DFFARX1 I_29798 (I509429,I2859,I509042,I509455,);
not I_29799 (I509463,I509455);
nand I_29800 (I509480,I509463,I509141);
nor I_29801 (I509497,I509480,I268957);
DFFARX1 I_29802 (I509497,I2859,I509042,I509010,);
nor I_29803 (I509528,I509463,I509192);
nor I_29804 (I509019,I509336,I509528);
not I_29805 (I509586,I2866);
DFFARX1 I_29806 (I65591,I2859,I509586,I509612,);
nand I_29807 (I509620,I509612,I65606);
DFFARX1 I_29808 (I65603,I2859,I509586,I509646,);
DFFARX1 I_29809 (I509646,I2859,I509586,I509663,);
not I_29810 (I509578,I509663);
not I_29811 (I509685,I65582);
nor I_29812 (I509702,I65582,I65588);
not I_29813 (I509719,I65594);
nand I_29814 (I509736,I509685,I509719);
nor I_29815 (I509753,I65594,I65582);
and I_29816 (I509557,I509753,I509620);
not I_29817 (I509784,I65600);
nand I_29818 (I509801,I509784,I65582);
nor I_29819 (I509818,I65600,I65585);
not I_29820 (I509835,I509818);
nand I_29821 (I509560,I509702,I509835);
DFFARX1 I_29822 (I509818,I2859,I509586,I509575,);
nor I_29823 (I509880,I65585,I65594);
nor I_29824 (I509897,I509880,I65588);
and I_29825 (I509914,I509897,I509801);
DFFARX1 I_29826 (I509914,I2859,I509586,I509572,);
nor I_29827 (I509569,I509880,I509736);
or I_29828 (I509566,I509818,I509880);
nor I_29829 (I509973,I65585,I65597);
DFFARX1 I_29830 (I509973,I2859,I509586,I509999,);
not I_29831 (I510007,I509999);
nand I_29832 (I510024,I510007,I509685);
nor I_29833 (I510041,I510024,I65588);
DFFARX1 I_29834 (I510041,I2859,I509586,I509554,);
nor I_29835 (I510072,I510007,I509736);
nor I_29836 (I509563,I509880,I510072);
not I_29837 (I510130,I2866);
DFFARX1 I_29838 (I344949,I2859,I510130,I510156,);
nand I_29839 (I510164,I510156,I344943);
DFFARX1 I_29840 (I344946,I2859,I510130,I510190,);
DFFARX1 I_29841 (I510190,I2859,I510130,I510207,);
not I_29842 (I510122,I510207);
not I_29843 (I510229,I344952);
nor I_29844 (I510246,I344952,I344946);
not I_29845 (I510263,I344955);
nand I_29846 (I510280,I510229,I510263);
nor I_29847 (I510297,I344955,I344952);
and I_29848 (I510101,I510297,I510164);
not I_29849 (I510328,I344964);
nand I_29850 (I510345,I510328,I344958);
nor I_29851 (I510362,I344964,I344961);
not I_29852 (I510379,I510362);
nand I_29853 (I510104,I510246,I510379);
DFFARX1 I_29854 (I510362,I2859,I510130,I510119,);
nor I_29855 (I510424,I344943,I344955);
nor I_29856 (I510441,I510424,I344946);
and I_29857 (I510458,I510441,I510345);
DFFARX1 I_29858 (I510458,I2859,I510130,I510116,);
nor I_29859 (I510113,I510424,I510280);
or I_29860 (I510110,I510362,I510424);
nor I_29861 (I510517,I344943,I344949);
DFFARX1 I_29862 (I510517,I2859,I510130,I510543,);
not I_29863 (I510551,I510543);
nand I_29864 (I510568,I510551,I510229);
nor I_29865 (I510585,I510568,I344946);
DFFARX1 I_29866 (I510585,I2859,I510130,I510098,);
nor I_29867 (I510616,I510551,I510280);
nor I_29868 (I510107,I510424,I510616);
not I_29869 (I510674,I2866);
DFFARX1 I_29870 (I225607,I2859,I510674,I510700,);
nand I_29871 (I510708,I510700,I225595);
DFFARX1 I_29872 (I225601,I2859,I510674,I510734,);
DFFARX1 I_29873 (I510734,I2859,I510674,I510751,);
not I_29874 (I510666,I510751);
not I_29875 (I510773,I225586);
nor I_29876 (I510790,I225586,I225598);
not I_29877 (I510807,I225589);
nand I_29878 (I510824,I510773,I510807);
nor I_29879 (I510841,I225589,I225586);
and I_29880 (I510645,I510841,I510708);
not I_29881 (I510872,I225604);
nand I_29882 (I510889,I510872,I225586);
nor I_29883 (I510906,I225604,I225610);
not I_29884 (I510923,I510906);
nand I_29885 (I510648,I510790,I510923);
DFFARX1 I_29886 (I510906,I2859,I510674,I510663,);
nor I_29887 (I510968,I225592,I225589);
nor I_29888 (I510985,I510968,I225598);
and I_29889 (I511002,I510985,I510889);
DFFARX1 I_29890 (I511002,I2859,I510674,I510660,);
nor I_29891 (I510657,I510968,I510824);
or I_29892 (I510654,I510906,I510968);
nor I_29893 (I511061,I225592,I225589);
DFFARX1 I_29894 (I511061,I2859,I510674,I511087,);
not I_29895 (I511095,I511087);
nand I_29896 (I511112,I511095,I510773);
nor I_29897 (I511129,I511112,I225598);
DFFARX1 I_29898 (I511129,I2859,I510674,I510642,);
nor I_29899 (I511160,I511095,I510824);
nor I_29900 (I510651,I510968,I511160);
not I_29901 (I511218,I2866);
DFFARX1 I_29902 (I2764,I2859,I511218,I511244,);
nand I_29903 (I511252,I511244,I1620);
DFFARX1 I_29904 (I2156,I2859,I511218,I511278,);
DFFARX1 I_29905 (I511278,I2859,I511218,I511295,);
not I_29906 (I511210,I511295);
not I_29907 (I511317,I2500);
nor I_29908 (I511334,I2500,I1428);
not I_29909 (I511351,I2452);
nand I_29910 (I511368,I511317,I511351);
nor I_29911 (I511385,I2452,I2500);
and I_29912 (I511189,I511385,I511252);
not I_29913 (I511416,I1932);
nand I_29914 (I511433,I511416,I1828);
nor I_29915 (I511450,I1932,I1636);
not I_29916 (I511467,I511450);
nand I_29917 (I511192,I511334,I511467);
DFFARX1 I_29918 (I511450,I2859,I511218,I511207,);
nor I_29919 (I511512,I2076,I2452);
nor I_29920 (I511529,I511512,I1428);
and I_29921 (I511546,I511529,I511433);
DFFARX1 I_29922 (I511546,I2859,I511218,I511204,);
nor I_29923 (I511201,I511512,I511368);
or I_29924 (I511198,I511450,I511512);
nor I_29925 (I511605,I2076,I1884);
DFFARX1 I_29926 (I511605,I2859,I511218,I511631,);
not I_29927 (I511639,I511631);
nand I_29928 (I511656,I511639,I511317);
nor I_29929 (I511673,I511656,I1428);
DFFARX1 I_29930 (I511673,I2859,I511218,I511186,);
nor I_29931 (I511704,I511639,I511368);
nor I_29932 (I511195,I511512,I511704);
not I_29933 (I511762,I2866);
DFFARX1 I_29934 (I558252,I2859,I511762,I511788,);
nand I_29935 (I511796,I511788,I558237);
DFFARX1 I_29936 (I558231,I2859,I511762,I511822,);
DFFARX1 I_29937 (I511822,I2859,I511762,I511839,);
not I_29938 (I511754,I511839);
not I_29939 (I511861,I558225);
nor I_29940 (I511878,I558225,I558246);
not I_29941 (I511895,I558234);
nand I_29942 (I511912,I511861,I511895);
nor I_29943 (I511929,I558234,I558225);
and I_29944 (I511733,I511929,I511796);
not I_29945 (I511960,I558243);
nand I_29946 (I511977,I511960,I558249);
nor I_29947 (I511994,I558243,I558240);
not I_29948 (I512011,I511994);
nand I_29949 (I511736,I511878,I512011);
DFFARX1 I_29950 (I511994,I2859,I511762,I511751,);
nor I_29951 (I512056,I558228,I558234);
nor I_29952 (I512073,I512056,I558246);
and I_29953 (I512090,I512073,I511977);
DFFARX1 I_29954 (I512090,I2859,I511762,I511748,);
nor I_29955 (I511745,I512056,I511912);
or I_29956 (I511742,I511994,I512056);
nor I_29957 (I512149,I558228,I558225);
DFFARX1 I_29958 (I512149,I2859,I511762,I512175,);
not I_29959 (I512183,I512175);
nand I_29960 (I512200,I512183,I511861);
nor I_29961 (I512217,I512200,I558246);
DFFARX1 I_29962 (I512217,I2859,I511762,I511730,);
nor I_29963 (I512248,I512183,I511912);
nor I_29964 (I511739,I512056,I512248);
not I_29965 (I512306,I2866);
DFFARX1 I_29966 (I393461,I2859,I512306,I512332,);
nand I_29967 (I512340,I512332,I393461);
DFFARX1 I_29968 (I393473,I2859,I512306,I512366,);
DFFARX1 I_29969 (I512366,I2859,I512306,I512383,);
not I_29970 (I512298,I512383);
not I_29971 (I512405,I393467);
nor I_29972 (I512422,I393467,I393488);
not I_29973 (I512439,I393476);
nand I_29974 (I512456,I512405,I512439);
nor I_29975 (I512473,I393476,I393467);
and I_29976 (I512277,I512473,I512340);
not I_29977 (I512504,I393470);
nand I_29978 (I512521,I512504,I393485);
nor I_29979 (I512538,I393470,I393479);
not I_29980 (I512555,I512538);
nand I_29981 (I512280,I512422,I512555);
DFFARX1 I_29982 (I512538,I2859,I512306,I512295,);
nor I_29983 (I512600,I393482,I393476);
nor I_29984 (I512617,I512600,I393488);
and I_29985 (I512634,I512617,I512521);
DFFARX1 I_29986 (I512634,I2859,I512306,I512292,);
nor I_29987 (I512289,I512600,I512456);
or I_29988 (I512286,I512538,I512600);
nor I_29989 (I512693,I393482,I393464);
DFFARX1 I_29990 (I512693,I2859,I512306,I512719,);
not I_29991 (I512727,I512719);
nand I_29992 (I512744,I512727,I512405);
nor I_29993 (I512761,I512744,I393488);
DFFARX1 I_29994 (I512761,I2859,I512306,I512274,);
nor I_29995 (I512792,I512727,I512456);
nor I_29996 (I512283,I512600,I512792);
not I_29997 (I512850,I2866);
DFFARX1 I_29998 (I300729,I2859,I512850,I512876,);
nand I_29999 (I512884,I512876,I300744);
DFFARX1 I_30000 (I300738,I2859,I512850,I512910,);
DFFARX1 I_30001 (I512910,I2859,I512850,I512927,);
not I_30002 (I512842,I512927);
not I_30003 (I512949,I300741);
nor I_30004 (I512966,I300741,I300747);
not I_30005 (I512983,I300729);
nand I_30006 (I513000,I512949,I512983);
nor I_30007 (I513017,I300729,I300741);
and I_30008 (I512821,I513017,I512884);
not I_30009 (I513048,I300726);
nand I_30010 (I513065,I513048,I300732);
nor I_30011 (I513082,I300726,I300726);
not I_30012 (I513099,I513082);
nand I_30013 (I512824,I512966,I513099);
DFFARX1 I_30014 (I513082,I2859,I512850,I512839,);
nor I_30015 (I513144,I300735,I300729);
nor I_30016 (I513161,I513144,I300747);
and I_30017 (I513178,I513161,I513065);
DFFARX1 I_30018 (I513178,I2859,I512850,I512836,);
nor I_30019 (I512833,I513144,I513000);
or I_30020 (I512830,I513082,I513144);
nor I_30021 (I513237,I300735,I300750);
DFFARX1 I_30022 (I513237,I2859,I512850,I513263,);
not I_30023 (I513271,I513263);
nand I_30024 (I513288,I513271,I512949);
nor I_30025 (I513305,I513288,I300747);
DFFARX1 I_30026 (I513305,I2859,I512850,I512818,);
nor I_30027 (I513336,I513271,I513000);
nor I_30028 (I512827,I513144,I513336);
not I_30029 (I513394,I2866);
DFFARX1 I_30030 (I187632,I2859,I513394,I513420,);
nand I_30031 (I513428,I513420,I187629);
DFFARX1 I_30032 (I187608,I2859,I513394,I513454,);
DFFARX1 I_30033 (I513454,I2859,I513394,I513471,);
not I_30034 (I513386,I513471);
not I_30035 (I513493,I187623);
nor I_30036 (I513510,I187623,I187626);
not I_30037 (I513527,I187617);
nand I_30038 (I513544,I513493,I513527);
nor I_30039 (I513561,I187617,I187623);
and I_30040 (I513365,I513561,I513428);
not I_30041 (I513592,I187614);
nand I_30042 (I513609,I513592,I187635);
nor I_30043 (I513626,I187614,I187611);
not I_30044 (I513643,I513626);
nand I_30045 (I513368,I513510,I513643);
DFFARX1 I_30046 (I513626,I2859,I513394,I513383,);
nor I_30047 (I513688,I187620,I187617);
nor I_30048 (I513705,I513688,I187626);
and I_30049 (I513722,I513705,I513609);
DFFARX1 I_30050 (I513722,I2859,I513394,I513380,);
nor I_30051 (I513377,I513688,I513544);
or I_30052 (I513374,I513626,I513688);
nor I_30053 (I513781,I187620,I187608);
DFFARX1 I_30054 (I513781,I2859,I513394,I513807,);
not I_30055 (I513815,I513807);
nand I_30056 (I513832,I513815,I513493);
nor I_30057 (I513849,I513832,I187626);
DFFARX1 I_30058 (I513849,I2859,I513394,I513362,);
nor I_30059 (I513880,I513815,I513544);
nor I_30060 (I513371,I513688,I513880);
not I_30061 (I513938,I2866);
DFFARX1 I_30062 (I88796,I2859,I513938,I513964,);
nand I_30063 (I513972,I513964,I88811);
DFFARX1 I_30064 (I88808,I2859,I513938,I513998,);
DFFARX1 I_30065 (I513998,I2859,I513938,I514015,);
not I_30066 (I513930,I514015);
not I_30067 (I514037,I88787);
nor I_30068 (I514054,I88787,I88793);
not I_30069 (I514071,I88799);
nand I_30070 (I514088,I514037,I514071);
nor I_30071 (I514105,I88799,I88787);
and I_30072 (I513909,I514105,I513972);
not I_30073 (I514136,I88805);
nand I_30074 (I514153,I514136,I88787);
nor I_30075 (I514170,I88805,I88790);
not I_30076 (I514187,I514170);
nand I_30077 (I513912,I514054,I514187);
DFFARX1 I_30078 (I514170,I2859,I513938,I513927,);
nor I_30079 (I514232,I88790,I88799);
nor I_30080 (I514249,I514232,I88793);
and I_30081 (I514266,I514249,I514153);
DFFARX1 I_30082 (I514266,I2859,I513938,I513924,);
nor I_30083 (I513921,I514232,I514088);
or I_30084 (I513918,I514170,I514232);
nor I_30085 (I514325,I88790,I88802);
DFFARX1 I_30086 (I514325,I2859,I513938,I514351,);
not I_30087 (I514359,I514351);
nand I_30088 (I514376,I514359,I514037);
nor I_30089 (I514393,I514376,I88793);
DFFARX1 I_30090 (I514393,I2859,I513938,I513906,);
nor I_30091 (I514424,I514359,I514088);
nor I_30092 (I513915,I514232,I514424);
not I_30093 (I514482,I2866);
DFFARX1 I_30094 (I498460,I2859,I514482,I514508,);
nand I_30095 (I514516,I514508,I498439);
DFFARX1 I_30096 (I498436,I2859,I514482,I514542,);
DFFARX1 I_30097 (I514542,I2859,I514482,I514559,);
not I_30098 (I514474,I514559);
not I_30099 (I514581,I498448);
nor I_30100 (I514598,I498448,I498457);
not I_30101 (I514615,I498445);
nand I_30102 (I514632,I514581,I514615);
nor I_30103 (I514649,I498445,I498448);
and I_30104 (I514453,I514649,I514516);
not I_30105 (I514680,I498454);
nand I_30106 (I514697,I514680,I498451);
nor I_30107 (I514714,I498454,I498436);
not I_30108 (I514731,I514714);
nand I_30109 (I514456,I514598,I514731);
DFFARX1 I_30110 (I514714,I2859,I514482,I514471,);
nor I_30111 (I514776,I498439,I498445);
nor I_30112 (I514793,I514776,I498457);
and I_30113 (I514810,I514793,I514697);
DFFARX1 I_30114 (I514810,I2859,I514482,I514468,);
nor I_30115 (I514465,I514776,I514632);
or I_30116 (I514462,I514714,I514776);
nor I_30117 (I514869,I498439,I498442);
DFFARX1 I_30118 (I514869,I2859,I514482,I514895,);
not I_30119 (I514903,I514895);
nand I_30120 (I514920,I514903,I514581);
nor I_30121 (I514937,I514920,I498457);
DFFARX1 I_30122 (I514937,I2859,I514482,I514450,);
nor I_30123 (I514968,I514903,I514632);
nor I_30124 (I514459,I514776,I514968);
not I_30125 (I515026,I2866);
DFFARX1 I_30126 (I159366,I2859,I515026,I515052,);
nand I_30127 (I515060,I515052,I159369);
DFFARX1 I_30128 (I159363,I2859,I515026,I515086,);
DFFARX1 I_30129 (I515086,I2859,I515026,I515103,);
not I_30130 (I515018,I515103);
not I_30131 (I515125,I159372);
nor I_30132 (I515142,I159372,I159357);
not I_30133 (I515159,I159381);
nand I_30134 (I515176,I515125,I515159);
nor I_30135 (I515193,I159381,I159372);
and I_30136 (I514997,I515193,I515060);
not I_30137 (I515224,I159360);
nand I_30138 (I515241,I515224,I159378);
nor I_30139 (I515258,I159360,I159354);
not I_30140 (I515275,I515258);
nand I_30141 (I515000,I515142,I515275);
DFFARX1 I_30142 (I515258,I2859,I515026,I515015,);
nor I_30143 (I515320,I159375,I159381);
nor I_30144 (I515337,I515320,I159357);
and I_30145 (I515354,I515337,I515241);
DFFARX1 I_30146 (I515354,I2859,I515026,I515012,);
nor I_30147 (I515009,I515320,I515176);
or I_30148 (I515006,I515258,I515320);
nor I_30149 (I515413,I159375,I159354);
DFFARX1 I_30150 (I515413,I2859,I515026,I515439,);
not I_30151 (I515447,I515439);
nand I_30152 (I515464,I515447,I515125);
nor I_30153 (I515481,I515464,I159357);
DFFARX1 I_30154 (I515481,I2859,I515026,I514994,);
nor I_30155 (I515512,I515447,I515176);
nor I_30156 (I515003,I515320,I515512);
not I_30157 (I515570,I2866);
DFFARX1 I_30158 (I221561,I2859,I515570,I515596,);
nand I_30159 (I515604,I515596,I221549);
DFFARX1 I_30160 (I221555,I2859,I515570,I515630,);
DFFARX1 I_30161 (I515630,I2859,I515570,I515647,);
not I_30162 (I515562,I515647);
not I_30163 (I515669,I221540);
nor I_30164 (I515686,I221540,I221552);
not I_30165 (I515703,I221543);
nand I_30166 (I515720,I515669,I515703);
nor I_30167 (I515737,I221543,I221540);
and I_30168 (I515541,I515737,I515604);
not I_30169 (I515768,I221558);
nand I_30170 (I515785,I515768,I221540);
nor I_30171 (I515802,I221558,I221564);
not I_30172 (I515819,I515802);
nand I_30173 (I515544,I515686,I515819);
DFFARX1 I_30174 (I515802,I2859,I515570,I515559,);
nor I_30175 (I515864,I221546,I221543);
nor I_30176 (I515881,I515864,I221552);
and I_30177 (I515898,I515881,I515785);
DFFARX1 I_30178 (I515898,I2859,I515570,I515556,);
nor I_30179 (I515553,I515864,I515720);
or I_30180 (I515550,I515802,I515864);
nor I_30181 (I515957,I221546,I221543);
DFFARX1 I_30182 (I515957,I2859,I515570,I515983,);
not I_30183 (I515991,I515983);
nand I_30184 (I516008,I515991,I515669);
nor I_30185 (I516025,I516008,I221552);
DFFARX1 I_30186 (I516025,I2859,I515570,I515538,);
nor I_30187 (I516056,I515991,I515720);
nor I_30188 (I515547,I515864,I516056);
not I_30189 (I516114,I2866);
DFFARX1 I_30190 (I472450,I2859,I516114,I516140,);
nand I_30191 (I516148,I516140,I472429);
DFFARX1 I_30192 (I472426,I2859,I516114,I516174,);
DFFARX1 I_30193 (I516174,I2859,I516114,I516191,);
not I_30194 (I516106,I516191);
not I_30195 (I516213,I472438);
nor I_30196 (I516230,I472438,I472447);
not I_30197 (I516247,I472435);
nand I_30198 (I516264,I516213,I516247);
nor I_30199 (I516281,I472435,I472438);
and I_30200 (I516085,I516281,I516148);
not I_30201 (I516312,I472444);
nand I_30202 (I516329,I516312,I472441);
nor I_30203 (I516346,I472444,I472426);
not I_30204 (I516363,I516346);
nand I_30205 (I516088,I516230,I516363);
DFFARX1 I_30206 (I516346,I2859,I516114,I516103,);
nor I_30207 (I516408,I472429,I472435);
nor I_30208 (I516425,I516408,I472447);
and I_30209 (I516442,I516425,I516329);
DFFARX1 I_30210 (I516442,I2859,I516114,I516100,);
nor I_30211 (I516097,I516408,I516264);
or I_30212 (I516094,I516346,I516408);
nor I_30213 (I516501,I472429,I472432);
DFFARX1 I_30214 (I516501,I2859,I516114,I516527,);
not I_30215 (I516535,I516527);
nand I_30216 (I516552,I516535,I516213);
nor I_30217 (I516569,I516552,I472447);
DFFARX1 I_30218 (I516569,I2859,I516114,I516082,);
nor I_30219 (I516600,I516535,I516264);
nor I_30220 (I516091,I516408,I516600);
not I_30221 (I516658,I2866);
DFFARX1 I_30222 (I145137,I2859,I516658,I516684,);
nand I_30223 (I516692,I516684,I145140);
DFFARX1 I_30224 (I145134,I2859,I516658,I516718,);
DFFARX1 I_30225 (I516718,I2859,I516658,I516735,);
not I_30226 (I516650,I516735);
not I_30227 (I516757,I145143);
nor I_30228 (I516774,I145143,I145128);
not I_30229 (I516791,I145152);
nand I_30230 (I516808,I516757,I516791);
nor I_30231 (I516825,I145152,I145143);
and I_30232 (I516629,I516825,I516692);
not I_30233 (I516856,I145131);
nand I_30234 (I516873,I516856,I145149);
nor I_30235 (I516890,I145131,I145125);
not I_30236 (I516907,I516890);
nand I_30237 (I516632,I516774,I516907);
DFFARX1 I_30238 (I516890,I2859,I516658,I516647,);
nor I_30239 (I516952,I145146,I145152);
nor I_30240 (I516969,I516952,I145128);
and I_30241 (I516986,I516969,I516873);
DFFARX1 I_30242 (I516986,I2859,I516658,I516644,);
nor I_30243 (I516641,I516952,I516808);
or I_30244 (I516638,I516890,I516952);
nor I_30245 (I517045,I145146,I145125);
DFFARX1 I_30246 (I517045,I2859,I516658,I517071,);
not I_30247 (I517079,I517071);
nand I_30248 (I517096,I517079,I516757);
nor I_30249 (I517113,I517096,I145128);
DFFARX1 I_30250 (I517113,I2859,I516658,I516626,);
nor I_30251 (I517144,I517079,I516808);
nor I_30252 (I516635,I516952,I517144);
not I_30253 (I517202,I2866);
DFFARX1 I_30254 (I512833,I2859,I517202,I517228,);
nand I_30255 (I517236,I517228,I512842);
not I_30256 (I517253,I517236);
DFFARX1 I_30257 (I512818,I2859,I517202,I517279,);
not I_30258 (I517287,I517279);
not I_30259 (I517304,I512821);
or I_30260 (I517321,I512818,I512821);
nor I_30261 (I517338,I512818,I512821);
or I_30262 (I517355,I512836,I512818);
DFFARX1 I_30263 (I517355,I2859,I517202,I517194,);
not I_30264 (I517386,I512824);
nand I_30265 (I517403,I517386,I512839);
nand I_30266 (I517420,I517304,I517403);
and I_30267 (I517173,I517287,I517420);
nor I_30268 (I517451,I512824,I512827);
and I_30269 (I517468,I517287,I517451);
nor I_30270 (I517179,I517253,I517468);
DFFARX1 I_30271 (I517451,I2859,I517202,I517508,);
not I_30272 (I517516,I517508);
nor I_30273 (I517188,I517287,I517516);
or I_30274 (I517547,I517355,I512830);
nor I_30275 (I517564,I512830,I512836);
nand I_30276 (I517581,I517420,I517564);
nand I_30277 (I517598,I517547,I517581);
DFFARX1 I_30278 (I517598,I2859,I517202,I517191,);
nor I_30279 (I517629,I517564,I517321);
DFFARX1 I_30280 (I517629,I2859,I517202,I517170,);
nor I_30281 (I517660,I512830,I512821);
DFFARX1 I_30282 (I517660,I2859,I517202,I517686,);
DFFARX1 I_30283 (I517686,I2859,I517202,I517185,);
not I_30284 (I517708,I517686);
nand I_30285 (I517182,I517708,I517236);
nand I_30286 (I517176,I517708,I517338);
not I_30287 (I517780,I2866);
DFFARX1 I_30288 (I235415,I2859,I517780,I517806,);
nand I_30289 (I517814,I517806,I235430);
not I_30290 (I517831,I517814);
DFFARX1 I_30291 (I235412,I2859,I517780,I517857,);
not I_30292 (I517865,I517857);
not I_30293 (I517882,I235421);
or I_30294 (I517899,I235415,I235421);
nor I_30295 (I517916,I235415,I235421);
or I_30296 (I517933,I235412,I235415);
DFFARX1 I_30297 (I517933,I2859,I517780,I517772,);
not I_30298 (I517964,I235433);
nand I_30299 (I517981,I517964,I235436);
nand I_30300 (I517998,I517882,I517981);
and I_30301 (I517751,I517865,I517998);
nor I_30302 (I518029,I235433,I235418);
and I_30303 (I518046,I517865,I518029);
nor I_30304 (I517757,I517831,I518046);
DFFARX1 I_30305 (I518029,I2859,I517780,I518086,);
not I_30306 (I518094,I518086);
nor I_30307 (I517766,I517865,I518094);
or I_30308 (I518125,I517933,I235424);
nor I_30309 (I518142,I235424,I235412);
nand I_30310 (I518159,I517998,I518142);
nand I_30311 (I518176,I518125,I518159);
DFFARX1 I_30312 (I518176,I2859,I517780,I517769,);
nor I_30313 (I518207,I518142,I517899);
DFFARX1 I_30314 (I518207,I2859,I517780,I517748,);
nor I_30315 (I518238,I235424,I235427);
DFFARX1 I_30316 (I518238,I2859,I517780,I518264,);
DFFARX1 I_30317 (I518264,I2859,I517780,I517763,);
not I_30318 (I518286,I518264);
nand I_30319 (I517760,I518286,I517814);
nand I_30320 (I517754,I518286,I517916);
not I_30321 (I518358,I2866);
DFFARX1 I_30322 (I428252,I2859,I518358,I518384,);
nand I_30323 (I518392,I518384,I428249);
not I_30324 (I518409,I518392);
DFFARX1 I_30325 (I428249,I2859,I518358,I518435,);
not I_30326 (I518443,I518435);
not I_30327 (I518460,I428246);
or I_30328 (I518477,I428255,I428246);
nor I_30329 (I518494,I428255,I428246);
or I_30330 (I518511,I428258,I428255);
DFFARX1 I_30331 (I518511,I2859,I518358,I518350,);
not I_30332 (I518542,I428246);
nand I_30333 (I518559,I518542,I428243);
nand I_30334 (I518576,I518460,I518559);
and I_30335 (I518329,I518443,I518576);
nor I_30336 (I518607,I428246,I428261);
and I_30337 (I518624,I518443,I518607);
nor I_30338 (I518335,I518409,I518624);
DFFARX1 I_30339 (I518607,I2859,I518358,I518664,);
not I_30340 (I518672,I518664);
nor I_30341 (I518344,I518443,I518672);
or I_30342 (I518703,I518511,I428264);
nor I_30343 (I518720,I428264,I428258);
nand I_30344 (I518737,I518576,I518720);
nand I_30345 (I518754,I518703,I518737);
DFFARX1 I_30346 (I518754,I2859,I518358,I518347,);
nor I_30347 (I518785,I518720,I518477);
DFFARX1 I_30348 (I518785,I2859,I518358,I518326,);
nor I_30349 (I518816,I428264,I428243);
DFFARX1 I_30350 (I518816,I2859,I518358,I518842,);
DFFARX1 I_30351 (I518842,I2859,I518358,I518341,);
not I_30352 (I518864,I518842);
nand I_30353 (I518338,I518864,I518392);
nand I_30354 (I518332,I518864,I518494);
not I_30355 (I518936,I2866);
DFFARX1 I_30356 (I263156,I2859,I518936,I518962,);
nand I_30357 (I518970,I518962,I263159);
not I_30358 (I518987,I518970);
DFFARX1 I_30359 (I263171,I2859,I518936,I519013,);
not I_30360 (I519021,I519013);
not I_30361 (I519038,I263156);
or I_30362 (I519055,I263165,I263156);
nor I_30363 (I519072,I263165,I263156);
or I_30364 (I519089,I263174,I263165);
DFFARX1 I_30365 (I519089,I2859,I518936,I518928,);
not I_30366 (I519120,I263177);
nand I_30367 (I519137,I519120,I263159);
nand I_30368 (I519154,I519038,I519137);
and I_30369 (I518907,I519021,I519154);
nor I_30370 (I519185,I263177,I263162);
and I_30371 (I519202,I519021,I519185);
nor I_30372 (I518913,I518987,I519202);
DFFARX1 I_30373 (I519185,I2859,I518936,I519242,);
not I_30374 (I519250,I519242);
nor I_30375 (I518922,I519021,I519250);
or I_30376 (I519281,I519089,I263168);
nor I_30377 (I519298,I263168,I263174);
nand I_30378 (I519315,I519154,I519298);
nand I_30379 (I519332,I519281,I519315);
DFFARX1 I_30380 (I519332,I2859,I518936,I518925,);
nor I_30381 (I519363,I519298,I519055);
DFFARX1 I_30382 (I519363,I2859,I518936,I518904,);
nor I_30383 (I519394,I263168,I263180);
DFFARX1 I_30384 (I519394,I2859,I518936,I519420,);
DFFARX1 I_30385 (I519420,I2859,I518936,I518919,);
not I_30386 (I519442,I519420);
nand I_30387 (I518916,I519442,I518970);
nand I_30388 (I518910,I519442,I519072);
not I_30389 (I519514,I2866);
DFFARX1 I_30390 (I4657,I2859,I519514,I519540,);
nand I_30391 (I519548,I519540,I4654);
not I_30392 (I519565,I519548);
DFFARX1 I_30393 (I4675,I2859,I519514,I519591,);
not I_30394 (I519599,I519591);
not I_30395 (I519616,I4660);
or I_30396 (I519633,I4669,I4660);
nor I_30397 (I519650,I4669,I4660);
or I_30398 (I519667,I4654,I4669);
DFFARX1 I_30399 (I519667,I2859,I519514,I519506,);
not I_30400 (I519698,I4666);
nand I_30401 (I519715,I519698,I4672);
nand I_30402 (I519732,I519616,I519715);
and I_30403 (I519485,I519599,I519732);
nor I_30404 (I519763,I4666,I4660);
and I_30405 (I519780,I519599,I519763);
nor I_30406 (I519491,I519565,I519780);
DFFARX1 I_30407 (I519763,I2859,I519514,I519820,);
not I_30408 (I519828,I519820);
nor I_30409 (I519500,I519599,I519828);
or I_30410 (I519859,I519667,I4657);
nor I_30411 (I519876,I4657,I4654);
nand I_30412 (I519893,I519732,I519876);
nand I_30413 (I519910,I519859,I519893);
DFFARX1 I_30414 (I519910,I2859,I519514,I519503,);
nor I_30415 (I519941,I519876,I519633);
DFFARX1 I_30416 (I519941,I2859,I519514,I519482,);
nor I_30417 (I519972,I4657,I4663);
DFFARX1 I_30418 (I519972,I2859,I519514,I519998,);
DFFARX1 I_30419 (I519998,I2859,I519514,I519497,);
not I_30420 (I520020,I519998);
nand I_30421 (I519494,I520020,I519548);
nand I_30422 (I519488,I520020,I519650);
not I_30423 (I520092,I2866);
DFFARX1 I_30424 (I292056,I2859,I520092,I520118,);
nand I_30425 (I520126,I520118,I292059);
not I_30426 (I520143,I520126);
DFFARX1 I_30427 (I292071,I2859,I520092,I520169,);
not I_30428 (I520177,I520169);
not I_30429 (I520194,I292056);
or I_30430 (I520211,I292065,I292056);
nor I_30431 (I520228,I292065,I292056);
or I_30432 (I520245,I292074,I292065);
DFFARX1 I_30433 (I520245,I2859,I520092,I520084,);
not I_30434 (I520276,I292077);
nand I_30435 (I520293,I520276,I292059);
nand I_30436 (I520310,I520194,I520293);
and I_30437 (I520063,I520177,I520310);
nor I_30438 (I520341,I292077,I292062);
and I_30439 (I520358,I520177,I520341);
nor I_30440 (I520069,I520143,I520358);
DFFARX1 I_30441 (I520341,I2859,I520092,I520398,);
not I_30442 (I520406,I520398);
nor I_30443 (I520078,I520177,I520406);
or I_30444 (I520437,I520245,I292068);
nor I_30445 (I520454,I292068,I292074);
nand I_30446 (I520471,I520310,I520454);
nand I_30447 (I520488,I520437,I520471);
DFFARX1 I_30448 (I520488,I2859,I520092,I520081,);
nor I_30449 (I520519,I520454,I520211);
DFFARX1 I_30450 (I520519,I2859,I520092,I520060,);
nor I_30451 (I520550,I292068,I292080);
DFFARX1 I_30452 (I520550,I2859,I520092,I520576,);
DFFARX1 I_30453 (I520576,I2859,I520092,I520075,);
not I_30454 (I520598,I520576);
nand I_30455 (I520072,I520598,I520126);
nand I_30456 (I520066,I520598,I520228);
not I_30457 (I520670,I2866);
DFFARX1 I_30458 (I73912,I2859,I520670,I520696,);
nand I_30459 (I520704,I520696,I73915);
not I_30460 (I520721,I520704);
DFFARX1 I_30461 (I73924,I2859,I520670,I520747,);
not I_30462 (I520755,I520747);
not I_30463 (I520772,I73927);
or I_30464 (I520789,I73918,I73927);
nor I_30465 (I520806,I73918,I73927);
or I_30466 (I520823,I73930,I73918);
DFFARX1 I_30467 (I520823,I2859,I520670,I520662,);
not I_30468 (I520854,I73915);
nand I_30469 (I520871,I520854,I73921);
nand I_30470 (I520888,I520772,I520871);
and I_30471 (I520641,I520755,I520888);
nor I_30472 (I520919,I73915,I73933);
and I_30473 (I520936,I520755,I520919);
nor I_30474 (I520647,I520721,I520936);
DFFARX1 I_30475 (I520919,I2859,I520670,I520976,);
not I_30476 (I520984,I520976);
nor I_30477 (I520656,I520755,I520984);
or I_30478 (I521015,I520823,I73912);
nor I_30479 (I521032,I73912,I73930);
nand I_30480 (I521049,I520888,I521032);
nand I_30481 (I521066,I521015,I521049);
DFFARX1 I_30482 (I521066,I2859,I520670,I520659,);
nor I_30483 (I521097,I521032,I520789);
DFFARX1 I_30484 (I521097,I2859,I520670,I520638,);
nor I_30485 (I521128,I73912,I73936);
DFFARX1 I_30486 (I521128,I2859,I520670,I521154,);
DFFARX1 I_30487 (I521154,I2859,I520670,I520653,);
not I_30488 (I521176,I521154);
nand I_30489 (I520650,I521176,I520704);
nand I_30490 (I520644,I521176,I520806);
not I_30491 (I521248,I2866);
DFFARX1 I_30492 (I435545,I2859,I521248,I521274,);
nand I_30493 (I521282,I521274,I435542);
not I_30494 (I521299,I521282);
DFFARX1 I_30495 (I435542,I2859,I521248,I521325,);
not I_30496 (I521333,I521325);
not I_30497 (I521350,I435539);
or I_30498 (I521367,I435548,I435539);
nor I_30499 (I521384,I435548,I435539);
or I_30500 (I521401,I435551,I435548);
DFFARX1 I_30501 (I521401,I2859,I521248,I521240,);
not I_30502 (I521432,I435539);
nand I_30503 (I521449,I521432,I435536);
nand I_30504 (I521466,I521350,I521449);
and I_30505 (I521219,I521333,I521466);
nor I_30506 (I521497,I435539,I435554);
and I_30507 (I521514,I521333,I521497);
nor I_30508 (I521225,I521299,I521514);
DFFARX1 I_30509 (I521497,I2859,I521248,I521554,);
not I_30510 (I521562,I521554);
nor I_30511 (I521234,I521333,I521562);
or I_30512 (I521593,I521401,I435557);
nor I_30513 (I521610,I435557,I435551);
nand I_30514 (I521627,I521466,I521610);
nand I_30515 (I521644,I521593,I521627);
DFFARX1 I_30516 (I521644,I2859,I521248,I521237,);
nor I_30517 (I521675,I521610,I521367);
DFFARX1 I_30518 (I521675,I2859,I521248,I521216,);
nor I_30519 (I521706,I435557,I435536);
DFFARX1 I_30520 (I521706,I2859,I521248,I521732,);
DFFARX1 I_30521 (I521732,I2859,I521248,I521231,);
not I_30522 (I521754,I521732);
nand I_30523 (I521228,I521754,I521282);
nand I_30524 (I521222,I521754,I521384);
not I_30525 (I521826,I2866);
DFFARX1 I_30526 (I445856,I2859,I521826,I521852,);
nand I_30527 (I521860,I521852,I445841);
not I_30528 (I521877,I521860);
DFFARX1 I_30529 (I445844,I2859,I521826,I521903,);
not I_30530 (I521911,I521903);
not I_30531 (I521928,I445859);
or I_30532 (I521945,I445862,I445859);
nor I_30533 (I521962,I445862,I445859);
or I_30534 (I521979,I445838,I445862);
DFFARX1 I_30535 (I521979,I2859,I521826,I521818,);
not I_30536 (I522010,I445850);
nand I_30537 (I522027,I522010,I445853);
nand I_30538 (I522044,I521928,I522027);
and I_30539 (I521797,I521911,I522044);
nor I_30540 (I522075,I445850,I445847);
and I_30541 (I522092,I521911,I522075);
nor I_30542 (I521803,I521877,I522092);
DFFARX1 I_30543 (I522075,I2859,I521826,I522132,);
not I_30544 (I522140,I522132);
nor I_30545 (I521812,I521911,I522140);
or I_30546 (I522171,I521979,I445838);
nor I_30547 (I522188,I445838,I445838);
nand I_30548 (I522205,I522044,I522188);
nand I_30549 (I522222,I522171,I522205);
DFFARX1 I_30550 (I522222,I2859,I521826,I521815,);
nor I_30551 (I522253,I522188,I521945);
DFFARX1 I_30552 (I522253,I2859,I521826,I521794,);
nor I_30553 (I522284,I445838,I445841);
DFFARX1 I_30554 (I522284,I2859,I521826,I522310,);
DFFARX1 I_30555 (I522310,I2859,I521826,I521809,);
not I_30556 (I522332,I522310);
nand I_30557 (I521806,I522332,I521860);
nand I_30558 (I521800,I522332,I521962);
not I_30559 (I522404,I2866);
DFFARX1 I_30560 (I457994,I2859,I522404,I522430,);
nand I_30561 (I522438,I522430,I457979);
not I_30562 (I522455,I522438);
DFFARX1 I_30563 (I457982,I2859,I522404,I522481,);
not I_30564 (I522489,I522481);
not I_30565 (I522506,I457997);
or I_30566 (I522523,I458000,I457997);
nor I_30567 (I522540,I458000,I457997);
or I_30568 (I522557,I457976,I458000);
DFFARX1 I_30569 (I522557,I2859,I522404,I522396,);
not I_30570 (I522588,I457988);
nand I_30571 (I522605,I522588,I457991);
nand I_30572 (I522622,I522506,I522605);
and I_30573 (I522375,I522489,I522622);
nor I_30574 (I522653,I457988,I457985);
and I_30575 (I522670,I522489,I522653);
nor I_30576 (I522381,I522455,I522670);
DFFARX1 I_30577 (I522653,I2859,I522404,I522710,);
not I_30578 (I522718,I522710);
nor I_30579 (I522390,I522489,I522718);
or I_30580 (I522749,I522557,I457976);
nor I_30581 (I522766,I457976,I457976);
nand I_30582 (I522783,I522622,I522766);
nand I_30583 (I522800,I522749,I522783);
DFFARX1 I_30584 (I522800,I2859,I522404,I522393,);
nor I_30585 (I522831,I522766,I522523);
DFFARX1 I_30586 (I522831,I2859,I522404,I522372,);
nor I_30587 (I522862,I457976,I457979);
DFFARX1 I_30588 (I522862,I2859,I522404,I522888,);
DFFARX1 I_30589 (I522888,I2859,I522404,I522387,);
not I_30590 (I522910,I522888);
nand I_30591 (I522384,I522910,I522438);
nand I_30592 (I522378,I522910,I522540);
not I_30593 (I522982,I2866);
DFFARX1 I_30594 (I179451,I2859,I522982,I523008,);
nand I_30595 (I523016,I523008,I179460);
not I_30596 (I523033,I523016);
DFFARX1 I_30597 (I179448,I2859,I522982,I523059,);
not I_30598 (I523067,I523059);
not I_30599 (I523084,I179454);
or I_30600 (I523101,I179448,I179454);
nor I_30601 (I523118,I179448,I179454);
or I_30602 (I523135,I179463,I179448);
DFFARX1 I_30603 (I523135,I2859,I522982,I522974,);
not I_30604 (I523166,I179457);
nand I_30605 (I523183,I523166,I179472);
nand I_30606 (I523200,I523084,I523183);
and I_30607 (I522953,I523067,I523200);
nor I_30608 (I523231,I179457,I179475);
and I_30609 (I523248,I523067,I523231);
nor I_30610 (I522959,I523033,I523248);
DFFARX1 I_30611 (I523231,I2859,I522982,I523288,);
not I_30612 (I523296,I523288);
nor I_30613 (I522968,I523067,I523296);
or I_30614 (I523327,I523135,I179466);
nor I_30615 (I523344,I179466,I179463);
nand I_30616 (I523361,I523200,I523344);
nand I_30617 (I523378,I523327,I523361);
DFFARX1 I_30618 (I523378,I2859,I522982,I522971,);
nor I_30619 (I523409,I523344,I523101);
DFFARX1 I_30620 (I523409,I2859,I522982,I522950,);
nor I_30621 (I523440,I179466,I179469);
DFFARX1 I_30622 (I523440,I2859,I522982,I523466,);
DFFARX1 I_30623 (I523466,I2859,I522982,I522965,);
not I_30624 (I523488,I523466);
nand I_30625 (I522962,I523488,I523016);
nand I_30626 (I522956,I523488,I523118);
not I_30627 (I523560,I2866);
DFFARX1 I_30628 (I407679,I2859,I523560,I523586,);
nand I_30629 (I523594,I523586,I407700);
not I_30630 (I523611,I523594);
DFFARX1 I_30631 (I407673,I2859,I523560,I523637,);
not I_30632 (I523645,I523637);
not I_30633 (I523662,I407694);
or I_30634 (I523679,I407685,I407694);
nor I_30635 (I523696,I407685,I407694);
or I_30636 (I523713,I407688,I407685);
DFFARX1 I_30637 (I523713,I2859,I523560,I523552,);
not I_30638 (I523744,I407676);
nand I_30639 (I523761,I523744,I407691);
nand I_30640 (I523778,I523662,I523761);
and I_30641 (I523531,I523645,I523778);
nor I_30642 (I523809,I407676,I407673);
and I_30643 (I523826,I523645,I523809);
nor I_30644 (I523537,I523611,I523826);
DFFARX1 I_30645 (I523809,I2859,I523560,I523866,);
not I_30646 (I523874,I523866);
nor I_30647 (I523546,I523645,I523874);
or I_30648 (I523905,I523713,I407697);
nor I_30649 (I523922,I407697,I407688);
nand I_30650 (I523939,I523778,I523922);
nand I_30651 (I523956,I523905,I523939);
DFFARX1 I_30652 (I523956,I2859,I523560,I523549,);
nor I_30653 (I523987,I523922,I523679);
DFFARX1 I_30654 (I523987,I2859,I523560,I523528,);
nor I_30655 (I524018,I407697,I407682);
DFFARX1 I_30656 (I524018,I2859,I523560,I524044,);
DFFARX1 I_30657 (I524044,I2859,I523560,I523543,);
not I_30658 (I524066,I524044);
nand I_30659 (I523540,I524066,I523594);
nand I_30660 (I523534,I524066,I523696);
not I_30661 (I524138,I2866);
DFFARX1 I_30662 (I53697,I2859,I524138,I524164,);
nand I_30663 (I524172,I524164,I53706);
not I_30664 (I524189,I524172);
DFFARX1 I_30665 (I53688,I2859,I524138,I524215,);
not I_30666 (I524223,I524215);
not I_30667 (I524240,I53694);
or I_30668 (I524257,I53703,I53694);
nor I_30669 (I524274,I53703,I53694);
or I_30670 (I524291,I53691,I53703);
DFFARX1 I_30671 (I524291,I2859,I524138,I524130,);
not I_30672 (I524322,I53709);
nand I_30673 (I524339,I524322,I53682);
nand I_30674 (I524356,I524240,I524339);
and I_30675 (I524109,I524223,I524356);
nor I_30676 (I524387,I53709,I53685);
and I_30677 (I524404,I524223,I524387);
nor I_30678 (I524115,I524189,I524404);
DFFARX1 I_30679 (I524387,I2859,I524138,I524444,);
not I_30680 (I524452,I524444);
nor I_30681 (I524124,I524223,I524452);
or I_30682 (I524483,I524291,I53700);
nor I_30683 (I524500,I53700,I53691);
nand I_30684 (I524517,I524356,I524500);
nand I_30685 (I524534,I524483,I524517);
DFFARX1 I_30686 (I524534,I2859,I524138,I524127,);
nor I_30687 (I524565,I524500,I524257);
DFFARX1 I_30688 (I524565,I2859,I524138,I524106,);
nor I_30689 (I524596,I53700,I53682);
DFFARX1 I_30690 (I524596,I2859,I524138,I524622,);
DFFARX1 I_30691 (I524622,I2859,I524138,I524121,);
not I_30692 (I524644,I524622);
nand I_30693 (I524118,I524644,I524172);
nand I_30694 (I524112,I524644,I524274);
not I_30695 (I524716,I2866);
DFFARX1 I_30696 (I405741,I2859,I524716,I524742,);
nand I_30697 (I524750,I524742,I405762);
not I_30698 (I524767,I524750);
DFFARX1 I_30699 (I405735,I2859,I524716,I524793,);
not I_30700 (I524801,I524793);
not I_30701 (I524818,I405756);
or I_30702 (I524835,I405747,I405756);
nor I_30703 (I524852,I405747,I405756);
or I_30704 (I524869,I405750,I405747);
DFFARX1 I_30705 (I524869,I2859,I524716,I524708,);
not I_30706 (I524900,I405738);
nand I_30707 (I524917,I524900,I405753);
nand I_30708 (I524934,I524818,I524917);
and I_30709 (I524687,I524801,I524934);
nor I_30710 (I524965,I405738,I405735);
and I_30711 (I524982,I524801,I524965);
nor I_30712 (I524693,I524767,I524982);
DFFARX1 I_30713 (I524965,I2859,I524716,I525022,);
not I_30714 (I525030,I525022);
nor I_30715 (I524702,I524801,I525030);
or I_30716 (I525061,I524869,I405759);
nor I_30717 (I525078,I405759,I405750);
nand I_30718 (I525095,I524934,I525078);
nand I_30719 (I525112,I525061,I525095);
DFFARX1 I_30720 (I525112,I2859,I524716,I524705,);
nor I_30721 (I525143,I525078,I524835);
DFFARX1 I_30722 (I525143,I2859,I524716,I524684,);
nor I_30723 (I525174,I405759,I405744);
DFFARX1 I_30724 (I525174,I2859,I524716,I525200,);
DFFARX1 I_30725 (I525200,I2859,I524716,I524699,);
not I_30726 (I525222,I525200);
nand I_30727 (I524696,I525222,I524750);
nand I_30728 (I524690,I525222,I524852);
not I_30729 (I525294,I2866);
DFFARX1 I_30730 (I231947,I2859,I525294,I525320,);
nand I_30731 (I525328,I525320,I231962);
not I_30732 (I525345,I525328);
DFFARX1 I_30733 (I231944,I2859,I525294,I525371,);
not I_30734 (I525379,I525371);
not I_30735 (I525396,I231953);
or I_30736 (I525413,I231947,I231953);
nor I_30737 (I525430,I231947,I231953);
or I_30738 (I525447,I231944,I231947);
DFFARX1 I_30739 (I525447,I2859,I525294,I525286,);
not I_30740 (I525478,I231965);
nand I_30741 (I525495,I525478,I231968);
nand I_30742 (I525512,I525396,I525495);
and I_30743 (I525265,I525379,I525512);
nor I_30744 (I525543,I231965,I231950);
and I_30745 (I525560,I525379,I525543);
nor I_30746 (I525271,I525345,I525560);
DFFARX1 I_30747 (I525543,I2859,I525294,I525600,);
not I_30748 (I525608,I525600);
nor I_30749 (I525280,I525379,I525608);
or I_30750 (I525639,I525447,I231956);
nor I_30751 (I525656,I231956,I231944);
nand I_30752 (I525673,I525512,I525656);
nand I_30753 (I525690,I525639,I525673);
DFFARX1 I_30754 (I525690,I2859,I525294,I525283,);
nor I_30755 (I525721,I525656,I525413);
DFFARX1 I_30756 (I525721,I2859,I525294,I525262,);
nor I_30757 (I525752,I231956,I231959);
DFFARX1 I_30758 (I525752,I2859,I525294,I525778,);
DFFARX1 I_30759 (I525778,I2859,I525294,I525277,);
not I_30760 (I525800,I525778);
nand I_30761 (I525274,I525800,I525328);
nand I_30762 (I525268,I525800,I525430);
not I_30763 (I525872,I2866);
DFFARX1 I_30764 (I560034,I2859,I525872,I525898,);
nand I_30765 (I525906,I525898,I560025);
not I_30766 (I525923,I525906);
DFFARX1 I_30767 (I560010,I2859,I525872,I525949,);
not I_30768 (I525957,I525949);
not I_30769 (I525974,I560013);
or I_30770 (I525991,I560022,I560013);
nor I_30771 (I526008,I560022,I560013);
or I_30772 (I526025,I560019,I560022);
DFFARX1 I_30773 (I526025,I2859,I525872,I525864,);
not I_30774 (I526056,I560031);
nand I_30775 (I526073,I526056,I560010);
nand I_30776 (I526090,I525974,I526073);
and I_30777 (I525843,I525957,I526090);
nor I_30778 (I526121,I560031,I560016);
and I_30779 (I526138,I525957,I526121);
nor I_30780 (I525849,I525923,I526138);
DFFARX1 I_30781 (I526121,I2859,I525872,I526178,);
not I_30782 (I526186,I526178);
nor I_30783 (I525858,I525957,I526186);
or I_30784 (I526217,I526025,I560037);
nor I_30785 (I526234,I560037,I560019);
nand I_30786 (I526251,I526090,I526234);
nand I_30787 (I526268,I526217,I526251);
DFFARX1 I_30788 (I526268,I2859,I525872,I525861,);
nor I_30789 (I526299,I526234,I525991);
DFFARX1 I_30790 (I526299,I2859,I525872,I525840,);
nor I_30791 (I526330,I560037,I560028);
DFFARX1 I_30792 (I526330,I2859,I525872,I526356,);
DFFARX1 I_30793 (I526356,I2859,I525872,I525855,);
not I_30794 (I526378,I526356);
nand I_30795 (I525852,I526378,I525906);
nand I_30796 (I525846,I526378,I526008);
not I_30797 (I526450,I2866);
DFFARX1 I_30798 (I409617,I2859,I526450,I526476,);
nand I_30799 (I526484,I526476,I409638);
not I_30800 (I526501,I526484);
DFFARX1 I_30801 (I409611,I2859,I526450,I526527,);
not I_30802 (I526535,I526527);
not I_30803 (I526552,I409632);
or I_30804 (I526569,I409623,I409632);
nor I_30805 (I526586,I409623,I409632);
or I_30806 (I526603,I409626,I409623);
DFFARX1 I_30807 (I526603,I2859,I526450,I526442,);
not I_30808 (I526634,I409614);
nand I_30809 (I526651,I526634,I409629);
nand I_30810 (I526668,I526552,I526651);
and I_30811 (I526421,I526535,I526668);
nor I_30812 (I526699,I409614,I409611);
and I_30813 (I526716,I526535,I526699);
nor I_30814 (I526427,I526501,I526716);
DFFARX1 I_30815 (I526699,I2859,I526450,I526756,);
not I_30816 (I526764,I526756);
nor I_30817 (I526436,I526535,I526764);
or I_30818 (I526795,I526603,I409635);
nor I_30819 (I526812,I409635,I409626);
nand I_30820 (I526829,I526668,I526812);
nand I_30821 (I526846,I526795,I526829);
DFFARX1 I_30822 (I526846,I2859,I526450,I526439,);
nor I_30823 (I526877,I526812,I526569);
DFFARX1 I_30824 (I526877,I2859,I526450,I526418,);
nor I_30825 (I526908,I409635,I409620);
DFFARX1 I_30826 (I526908,I2859,I526450,I526934,);
DFFARX1 I_30827 (I526934,I2859,I526450,I526433,);
not I_30828 (I526956,I526934);
nand I_30829 (I526430,I526956,I526484);
nand I_30830 (I526424,I526956,I526586);
not I_30831 (I527028,I2866);
DFFARX1 I_30832 (I2612,I2859,I527028,I527054,);
nand I_30833 (I527062,I527054,I2236);
not I_30834 (I527079,I527062);
DFFARX1 I_30835 (I2060,I2859,I527028,I527105,);
not I_30836 (I527113,I527105);
not I_30837 (I527130,I1996);
or I_30838 (I527147,I2524,I1996);
nor I_30839 (I527164,I2524,I1996);
or I_30840 (I527181,I1644,I2524);
DFFARX1 I_30841 (I527181,I2859,I527028,I527020,);
not I_30842 (I527212,I1924);
nand I_30843 (I527229,I527212,I2756);
nand I_30844 (I527246,I527130,I527229);
and I_30845 (I526999,I527113,I527246);
nor I_30846 (I527277,I1924,I2084);
and I_30847 (I527294,I527113,I527277);
nor I_30848 (I527005,I527079,I527294);
DFFARX1 I_30849 (I527277,I2859,I527028,I527334,);
not I_30850 (I527342,I527334);
nor I_30851 (I527014,I527113,I527342);
or I_30852 (I527373,I527181,I2300);
nor I_30853 (I527390,I2300,I1644);
nand I_30854 (I527407,I527246,I527390);
nand I_30855 (I527424,I527373,I527407);
DFFARX1 I_30856 (I527424,I2859,I527028,I527017,);
nor I_30857 (I527455,I527390,I527147);
DFFARX1 I_30858 (I527455,I2859,I527028,I526996,);
nor I_30859 (I527486,I2300,I2660);
DFFARX1 I_30860 (I527486,I2859,I527028,I527512,);
DFFARX1 I_30861 (I527512,I2859,I527028,I527011,);
not I_30862 (I527534,I527512);
nand I_30863 (I527008,I527534,I527062);
nand I_30864 (I527002,I527534,I527164);
not I_30865 (I527606,I2866);
DFFARX1 I_30866 (I261422,I2859,I527606,I527632,);
nand I_30867 (I527640,I527632,I261425);
not I_30868 (I527657,I527640);
DFFARX1 I_30869 (I261437,I2859,I527606,I527683,);
not I_30870 (I527691,I527683);
not I_30871 (I527708,I261422);
or I_30872 (I527725,I261431,I261422);
nor I_30873 (I527742,I261431,I261422);
or I_30874 (I527759,I261440,I261431);
DFFARX1 I_30875 (I527759,I2859,I527606,I527598,);
not I_30876 (I527790,I261443);
nand I_30877 (I527807,I527790,I261425);
nand I_30878 (I527824,I527708,I527807);
and I_30879 (I527577,I527691,I527824);
nor I_30880 (I527855,I261443,I261428);
and I_30881 (I527872,I527691,I527855);
nor I_30882 (I527583,I527657,I527872);
DFFARX1 I_30883 (I527855,I2859,I527606,I527912,);
not I_30884 (I527920,I527912);
nor I_30885 (I527592,I527691,I527920);
or I_30886 (I527951,I527759,I261434);
nor I_30887 (I527968,I261434,I261440);
nand I_30888 (I527985,I527824,I527968);
nand I_30889 (I528002,I527951,I527985);
DFFARX1 I_30890 (I528002,I2859,I527606,I527595,);
nor I_30891 (I528033,I527968,I527725);
DFFARX1 I_30892 (I528033,I2859,I527606,I527574,);
nor I_30893 (I528064,I261434,I261446);
DFFARX1 I_30894 (I528064,I2859,I527606,I528090,);
DFFARX1 I_30895 (I528090,I2859,I527606,I527589,);
not I_30896 (I528112,I528090);
nand I_30897 (I527586,I528112,I527640);
nand I_30898 (I527580,I528112,I527742);
not I_30899 (I528184,I2866);
DFFARX1 I_30900 (I303616,I2859,I528184,I528210,);
nand I_30901 (I528218,I528210,I303619);
not I_30902 (I528235,I528218);
DFFARX1 I_30903 (I303631,I2859,I528184,I528261,);
not I_30904 (I528269,I528261);
not I_30905 (I528286,I303616);
or I_30906 (I528303,I303625,I303616);
nor I_30907 (I528320,I303625,I303616);
or I_30908 (I528337,I303634,I303625);
DFFARX1 I_30909 (I528337,I2859,I528184,I528176,);
not I_30910 (I528368,I303637);
nand I_30911 (I528385,I528368,I303619);
nand I_30912 (I528402,I528286,I528385);
and I_30913 (I528155,I528269,I528402);
nor I_30914 (I528433,I303637,I303622);
and I_30915 (I528450,I528269,I528433);
nor I_30916 (I528161,I528235,I528450);
DFFARX1 I_30917 (I528433,I2859,I528184,I528490,);
not I_30918 (I528498,I528490);
nor I_30919 (I528170,I528269,I528498);
or I_30920 (I528529,I528337,I303628);
nor I_30921 (I528546,I303628,I303634);
nand I_30922 (I528563,I528402,I528546);
nand I_30923 (I528580,I528529,I528563);
DFFARX1 I_30924 (I528580,I2859,I528184,I528173,);
nor I_30925 (I528611,I528546,I528303);
DFFARX1 I_30926 (I528611,I2859,I528184,I528152,);
nor I_30927 (I528642,I303628,I303640);
DFFARX1 I_30928 (I528642,I2859,I528184,I528668,);
DFFARX1 I_30929 (I528668,I2859,I528184,I528167,);
not I_30930 (I528690,I528668);
nand I_30931 (I528164,I528690,I528218);
nand I_30932 (I528158,I528690,I528320);
not I_30933 (I528762,I2866);
DFFARX1 I_30934 (I86407,I2859,I528762,I528788,);
nand I_30935 (I528796,I528788,I86410);
not I_30936 (I528813,I528796);
DFFARX1 I_30937 (I86419,I2859,I528762,I528839,);
not I_30938 (I528847,I528839);
not I_30939 (I528864,I86422);
or I_30940 (I528881,I86413,I86422);
nor I_30941 (I528898,I86413,I86422);
or I_30942 (I528915,I86425,I86413);
DFFARX1 I_30943 (I528915,I2859,I528762,I528754,);
not I_30944 (I528946,I86410);
nand I_30945 (I528963,I528946,I86416);
nand I_30946 (I528980,I528864,I528963);
and I_30947 (I528733,I528847,I528980);
nor I_30948 (I529011,I86410,I86428);
and I_30949 (I529028,I528847,I529011);
nor I_30950 (I528739,I528813,I529028);
DFFARX1 I_30951 (I529011,I2859,I528762,I529068,);
not I_30952 (I529076,I529068);
nor I_30953 (I528748,I528847,I529076);
or I_30954 (I529107,I528915,I86407);
nor I_30955 (I529124,I86407,I86425);
nand I_30956 (I529141,I528980,I529124);
nand I_30957 (I529158,I529107,I529141);
DFFARX1 I_30958 (I529158,I2859,I528762,I528751,);
nor I_30959 (I529189,I529124,I528881);
DFFARX1 I_30960 (I529189,I2859,I528762,I528730,);
nor I_30961 (I529220,I86407,I86431);
DFFARX1 I_30962 (I529220,I2859,I528762,I529246,);
DFFARX1 I_30963 (I529246,I2859,I528762,I528745,);
not I_30964 (I529268,I529246);
nand I_30965 (I528742,I529268,I528796);
nand I_30966 (I528736,I529268,I528898);
not I_30967 (I529340,I2866);
DFFARX1 I_30968 (I28517,I2859,I529340,I529366,);
nand I_30969 (I529374,I529366,I28508);
not I_30970 (I529391,I529374);
DFFARX1 I_30971 (I28505,I2859,I529340,I529417,);
not I_30972 (I529425,I529417);
not I_30973 (I529442,I28514);
or I_30974 (I529459,I28505,I28514);
nor I_30975 (I529476,I28505,I28514);
or I_30976 (I529493,I28511,I28505);
DFFARX1 I_30977 (I529493,I2859,I529340,I529332,);
not I_30978 (I529524,I28520);
nand I_30979 (I529541,I529524,I28529);
nand I_30980 (I529558,I529442,I529541);
and I_30981 (I529311,I529425,I529558);
nor I_30982 (I529589,I28520,I28523);
and I_30983 (I529606,I529425,I529589);
nor I_30984 (I529317,I529391,I529606);
DFFARX1 I_30985 (I529589,I2859,I529340,I529646,);
not I_30986 (I529654,I529646);
nor I_30987 (I529326,I529425,I529654);
or I_30988 (I529685,I529493,I28508);
nor I_30989 (I529702,I28508,I28511);
nand I_30990 (I529719,I529558,I529702);
nand I_30991 (I529736,I529685,I529719);
DFFARX1 I_30992 (I529736,I2859,I529340,I529329,);
nor I_30993 (I529767,I529702,I529459);
DFFARX1 I_30994 (I529767,I2859,I529340,I529308,);
nor I_30995 (I529798,I28508,I28526);
DFFARX1 I_30996 (I529798,I2859,I529340,I529824,);
DFFARX1 I_30997 (I529824,I2859,I529340,I529323,);
not I_30998 (I529846,I529824);
nand I_30999 (I529320,I529846,I529374);
nand I_31000 (I529314,I529846,I529476);
not I_31001 (I529918,I2866);
DFFARX1 I_31002 (I6904,I2859,I529918,I529944,);
nand I_31003 (I529952,I529944,I6898);
not I_31004 (I529969,I529952);
DFFARX1 I_31005 (I6916,I2859,I529918,I529995,);
not I_31006 (I530003,I529995);
not I_31007 (I530020,I6919);
or I_31008 (I530037,I6922,I6919);
nor I_31009 (I530054,I6922,I6919);
or I_31010 (I530071,I6907,I6922);
DFFARX1 I_31011 (I530071,I2859,I529918,I529910,);
not I_31012 (I530102,I6910);
nand I_31013 (I530119,I530102,I6913);
nand I_31014 (I530136,I530020,I530119);
and I_31015 (I529889,I530003,I530136);
nor I_31016 (I530167,I6910,I6901);
and I_31017 (I530184,I530003,I530167);
nor I_31018 (I529895,I529969,I530184);
DFFARX1 I_31019 (I530167,I2859,I529918,I530224,);
not I_31020 (I530232,I530224);
nor I_31021 (I529904,I530003,I530232);
or I_31022 (I530263,I530071,I6901);
nor I_31023 (I530280,I6901,I6907);
nand I_31024 (I530297,I530136,I530280);
nand I_31025 (I530314,I530263,I530297);
DFFARX1 I_31026 (I530314,I2859,I529918,I529907,);
nor I_31027 (I530345,I530280,I530037);
DFFARX1 I_31028 (I530345,I2859,I529918,I529886,);
nor I_31029 (I530376,I6901,I6898);
DFFARX1 I_31030 (I530376,I2859,I529918,I530402,);
DFFARX1 I_31031 (I530402,I2859,I529918,I529901,);
not I_31032 (I530424,I530402);
nand I_31033 (I529898,I530424,I529952);
nand I_31034 (I529892,I530424,I530054);
not I_31035 (I530496,I2866);
DFFARX1 I_31036 (I177819,I2859,I530496,I530522,);
nand I_31037 (I530530,I530522,I177828);
not I_31038 (I530547,I530530);
DFFARX1 I_31039 (I177816,I2859,I530496,I530573,);
not I_31040 (I530581,I530573);
not I_31041 (I530598,I177822);
or I_31042 (I530615,I177816,I177822);
nor I_31043 (I530632,I177816,I177822);
or I_31044 (I530649,I177831,I177816);
DFFARX1 I_31045 (I530649,I2859,I530496,I530488,);
not I_31046 (I530680,I177825);
nand I_31047 (I530697,I530680,I177840);
nand I_31048 (I530714,I530598,I530697);
and I_31049 (I530467,I530581,I530714);
nor I_31050 (I530745,I177825,I177843);
and I_31051 (I530762,I530581,I530745);
nor I_31052 (I530473,I530547,I530762);
DFFARX1 I_31053 (I530745,I2859,I530496,I530802,);
not I_31054 (I530810,I530802);
nor I_31055 (I530482,I530581,I530810);
or I_31056 (I530841,I530649,I177834);
nor I_31057 (I530858,I177834,I177831);
nand I_31058 (I530875,I530714,I530858);
nand I_31059 (I530892,I530841,I530875);
DFFARX1 I_31060 (I530892,I2859,I530496,I530485,);
nor I_31061 (I530923,I530858,I530615);
DFFARX1 I_31062 (I530923,I2859,I530496,I530464,);
nor I_31063 (I530954,I177834,I177837);
DFFARX1 I_31064 (I530954,I2859,I530496,I530980,);
DFFARX1 I_31065 (I530980,I2859,I530496,I530479,);
not I_31066 (I531002,I530980);
nand I_31067 (I530476,I531002,I530530);
nand I_31068 (I530470,I531002,I530632);
not I_31069 (I531074,I2866);
DFFARX1 I_31070 (I570744,I2859,I531074,I531100,);
nand I_31071 (I531108,I531100,I570735);
not I_31072 (I531125,I531108);
DFFARX1 I_31073 (I570720,I2859,I531074,I531151,);
not I_31074 (I531159,I531151);
not I_31075 (I531176,I570723);
or I_31076 (I531193,I570732,I570723);
nor I_31077 (I531210,I570732,I570723);
or I_31078 (I531227,I570729,I570732);
DFFARX1 I_31079 (I531227,I2859,I531074,I531066,);
not I_31080 (I531258,I570741);
nand I_31081 (I531275,I531258,I570720);
nand I_31082 (I531292,I531176,I531275);
and I_31083 (I531045,I531159,I531292);
nor I_31084 (I531323,I570741,I570726);
and I_31085 (I531340,I531159,I531323);
nor I_31086 (I531051,I531125,I531340);
DFFARX1 I_31087 (I531323,I2859,I531074,I531380,);
not I_31088 (I531388,I531380);
nor I_31089 (I531060,I531159,I531388);
or I_31090 (I531419,I531227,I570747);
nor I_31091 (I531436,I570747,I570729);
nand I_31092 (I531453,I531292,I531436);
nand I_31093 (I531470,I531419,I531453);
DFFARX1 I_31094 (I531470,I2859,I531074,I531063,);
nor I_31095 (I531501,I531436,I531193);
DFFARX1 I_31096 (I531501,I2859,I531074,I531042,);
nor I_31097 (I531532,I570747,I570738);
DFFARX1 I_31098 (I531532,I2859,I531074,I531558,);
DFFARX1 I_31099 (I531558,I2859,I531074,I531057,);
not I_31100 (I531580,I531558);
nand I_31101 (I531054,I531580,I531108);
nand I_31102 (I531048,I531580,I531210);
not I_31103 (I531655,I2866);
DFFARX1 I_31104 (I236014,I2859,I531655,I531681,);
nand I_31105 (I531689,I531681,I235993);
not I_31106 (I531706,I531689);
DFFARX1 I_31107 (I236005,I2859,I531655,I531732,);
not I_31108 (I531740,I531732);
nor I_31109 (I531757,I235993,I236002);
not I_31110 (I531774,I531757);
DFFARX1 I_31111 (I531774,I2859,I531655,I531641,);
or I_31112 (I531805,I235996,I235993);
DFFARX1 I_31113 (I531805,I2859,I531655,I531644,);
not I_31114 (I531836,I235999);
nor I_31115 (I531853,I531836,I235990);
nor I_31116 (I531870,I531853,I236002);
nor I_31117 (I531887,I235990,I236008);
nor I_31118 (I531904,I531740,I531887);
nor I_31119 (I531629,I531706,I531904);
not I_31120 (I531935,I531887);
nand I_31121 (I531632,I531935,I531689);
nand I_31122 (I531626,I531935,I531757);
nor I_31123 (I531623,I531887,I531870);
nor I_31124 (I531994,I236011,I235996);
not I_31125 (I532011,I531994);
DFFARX1 I_31126 (I531994,I2859,I531655,I532037,);
not I_31127 (I531647,I532037);
nor I_31128 (I532059,I236011,I235990);
DFFARX1 I_31129 (I532059,I2859,I531655,I532085,);
and I_31130 (I532093,I532085,I235993);
nor I_31131 (I532110,I532093,I532011);
DFFARX1 I_31132 (I532110,I2859,I531655,I531638,);
nor I_31133 (I532141,I532085,I531870);
DFFARX1 I_31134 (I532141,I2859,I531655,I531620,);
nor I_31135 (I531635,I532085,I531774);
not I_31136 (I532216,I2866);
DFFARX1 I_31137 (I571925,I2859,I532216,I532242,);
nand I_31138 (I532250,I532242,I571919);
not I_31139 (I532267,I532250);
DFFARX1 I_31140 (I571937,I2859,I532216,I532293,);
not I_31141 (I532301,I532293);
nor I_31142 (I532318,I571922,I571913);
not I_31143 (I532335,I532318);
DFFARX1 I_31144 (I532335,I2859,I532216,I532202,);
or I_31145 (I532366,I571928,I571922);
DFFARX1 I_31146 (I532366,I2859,I532216,I532205,);
not I_31147 (I532397,I571931);
nor I_31148 (I532414,I532397,I571934);
nor I_31149 (I532431,I532414,I571913);
nor I_31150 (I532448,I571934,I571916);
nor I_31151 (I532465,I532301,I532448);
nor I_31152 (I532190,I532267,I532465);
not I_31153 (I532496,I532448);
nand I_31154 (I532193,I532496,I532250);
nand I_31155 (I532187,I532496,I532318);
nor I_31156 (I532184,I532448,I532431);
nor I_31157 (I532555,I571910,I571928);
not I_31158 (I532572,I532555);
DFFARX1 I_31159 (I532555,I2859,I532216,I532598,);
not I_31160 (I532208,I532598);
nor I_31161 (I532620,I571910,I571910);
DFFARX1 I_31162 (I532620,I2859,I532216,I532646,);
and I_31163 (I532654,I532646,I571922);
nor I_31164 (I532671,I532654,I532572);
DFFARX1 I_31165 (I532671,I2859,I532216,I532199,);
nor I_31166 (I532702,I532646,I532431);
DFFARX1 I_31167 (I532702,I2859,I532216,I532181,);
nor I_31168 (I532196,I532646,I532335);
not I_31169 (I532777,I2866);
DFFARX1 I_31170 (I197421,I2859,I532777,I532803,);
nand I_31171 (I532811,I532803,I197403);
not I_31172 (I532828,I532811);
DFFARX1 I_31173 (I197400,I2859,I532777,I532854,);
not I_31174 (I532862,I532854);
nor I_31175 (I532879,I197406,I197400);
not I_31176 (I532896,I532879);
DFFARX1 I_31177 (I532896,I2859,I532777,I532763,);
or I_31178 (I532927,I197409,I197406);
DFFARX1 I_31179 (I532927,I2859,I532777,I532766,);
not I_31180 (I532958,I197415);
nor I_31181 (I532975,I532958,I197427);
nor I_31182 (I532992,I532975,I197400);
nor I_31183 (I533009,I197427,I197412);
nor I_31184 (I533026,I532862,I533009);
nor I_31185 (I532751,I532828,I533026);
not I_31186 (I533057,I533009);
nand I_31187 (I532754,I533057,I532811);
nand I_31188 (I532748,I533057,I532879);
nor I_31189 (I532745,I533009,I532992);
nor I_31190 (I533116,I197418,I197409);
not I_31191 (I533133,I533116);
DFFARX1 I_31192 (I533116,I2859,I532777,I533159,);
not I_31193 (I532769,I533159);
nor I_31194 (I533181,I197418,I197424);
DFFARX1 I_31195 (I533181,I2859,I532777,I533207,);
and I_31196 (I533215,I533207,I197406);
nor I_31197 (I533232,I533215,I533133);
DFFARX1 I_31198 (I533232,I2859,I532777,I532760,);
nor I_31199 (I533263,I533207,I532992);
DFFARX1 I_31200 (I533263,I2859,I532777,I532742,);
nor I_31201 (I532757,I533207,I532896);
not I_31202 (I533338,I2866);
DFFARX1 I_31203 (I2428,I2859,I533338,I533364,);
nand I_31204 (I533372,I533364,I2724);
not I_31205 (I533389,I533372);
DFFARX1 I_31206 (I2140,I2859,I533338,I533415,);
not I_31207 (I533423,I533415);
nor I_31208 (I533440,I1580,I2820);
not I_31209 (I533457,I533440);
DFFARX1 I_31210 (I533457,I2859,I533338,I533324,);
or I_31211 (I533488,I1404,I1580);
DFFARX1 I_31212 (I533488,I2859,I533338,I533327,);
not I_31213 (I533519,I2828);
nor I_31214 (I533536,I533519,I2748);
nor I_31215 (I533553,I533536,I2820);
nor I_31216 (I533570,I2748,I2532);
nor I_31217 (I533587,I533423,I533570);
nor I_31218 (I533312,I533389,I533587);
not I_31219 (I533618,I533570);
nand I_31220 (I533315,I533618,I533372);
nand I_31221 (I533309,I533618,I533440);
nor I_31222 (I533306,I533570,I533553);
nor I_31223 (I533677,I2372,I1404);
not I_31224 (I533694,I533677);
DFFARX1 I_31225 (I533677,I2859,I533338,I533720,);
not I_31226 (I533330,I533720);
nor I_31227 (I533742,I2372,I1364);
DFFARX1 I_31228 (I533742,I2859,I533338,I533768,);
and I_31229 (I533776,I533768,I1580);
nor I_31230 (I533793,I533776,I533694);
DFFARX1 I_31231 (I533793,I2859,I533338,I533321,);
nor I_31232 (I533824,I533768,I533553);
DFFARX1 I_31233 (I533824,I2859,I533338,I533303,);
nor I_31234 (I533318,I533768,I533457);
not I_31235 (I533899,I2866);
DFFARX1 I_31236 (I330717,I2859,I533899,I533925,);
nand I_31237 (I533933,I533925,I330735);
not I_31238 (I533950,I533933);
DFFARX1 I_31239 (I330714,I2859,I533899,I533976,);
not I_31240 (I533984,I533976);
nor I_31241 (I534001,I330729,I330723);
not I_31242 (I534018,I534001);
DFFARX1 I_31243 (I534018,I2859,I533899,I533885,);
or I_31244 (I534049,I330720,I330729);
DFFARX1 I_31245 (I534049,I2859,I533899,I533888,);
not I_31246 (I534080,I330720);
nor I_31247 (I534097,I534080,I330726);
nor I_31248 (I534114,I534097,I330723);
nor I_31249 (I534131,I330726,I330714);
nor I_31250 (I534148,I533984,I534131);
nor I_31251 (I533873,I533950,I534148);
not I_31252 (I534179,I534131);
nand I_31253 (I533876,I534179,I533933);
nand I_31254 (I533870,I534179,I534001);
nor I_31255 (I533867,I534131,I534114);
nor I_31256 (I534238,I330717,I330720);
not I_31257 (I534255,I534238);
DFFARX1 I_31258 (I534238,I2859,I533899,I534281,);
not I_31259 (I533891,I534281);
nor I_31260 (I534303,I330717,I330732);
DFFARX1 I_31261 (I534303,I2859,I533899,I534329,);
and I_31262 (I534337,I534329,I330729);
nor I_31263 (I534354,I534337,I534255);
DFFARX1 I_31264 (I534354,I2859,I533899,I533882,);
nor I_31265 (I534385,I534329,I534114);
DFFARX1 I_31266 (I534385,I2859,I533899,I533864,);
nor I_31267 (I533879,I534329,I534018);
not I_31268 (I534460,I2866);
DFFARX1 I_31269 (I324399,I2859,I534460,I534486,);
DFFARX1 I_31270 (I324396,I2859,I534460,I534503,);
not I_31271 (I534511,I534503);
nor I_31272 (I534428,I534486,I534511);
DFFARX1 I_31273 (I534511,I2859,I534460,I534443,);
nor I_31274 (I534556,I324411,I324393);
and I_31275 (I534573,I534556,I324390);
nor I_31276 (I534590,I534573,I324411);
not I_31277 (I534607,I324411);
and I_31278 (I534624,I534607,I324396);
nand I_31279 (I534641,I534624,I324408);
nor I_31280 (I534658,I534607,I534641);
DFFARX1 I_31281 (I534658,I2859,I534460,I534425,);
not I_31282 (I534689,I534641);
nand I_31283 (I534706,I534511,I534689);
nand I_31284 (I534437,I534573,I534689);
DFFARX1 I_31285 (I534607,I2859,I534460,I534452,);
not I_31286 (I534751,I324402);
nor I_31287 (I534768,I534751,I324396);
nor I_31288 (I534785,I534768,I534590);
DFFARX1 I_31289 (I534785,I2859,I534460,I534449,);
not I_31290 (I534816,I534768);
DFFARX1 I_31291 (I534816,I2859,I534460,I534842,);
not I_31292 (I534850,I534842);
nor I_31293 (I534446,I534850,I534768);
nor I_31294 (I534881,I534751,I324390);
and I_31295 (I534898,I534881,I324405);
or I_31296 (I534915,I534898,I324393);
DFFARX1 I_31297 (I534915,I2859,I534460,I534941,);
not I_31298 (I534949,I534941);
nand I_31299 (I534966,I534949,I534689);
not I_31300 (I534440,I534966);
nand I_31301 (I534434,I534966,I534706);
nand I_31302 (I534431,I534949,I534573);
not I_31303 (I535055,I2866);
DFFARX1 I_31304 (I335993,I2859,I535055,I535081,);
DFFARX1 I_31305 (I335990,I2859,I535055,I535098,);
not I_31306 (I535106,I535098);
nor I_31307 (I535023,I535081,I535106);
DFFARX1 I_31308 (I535106,I2859,I535055,I535038,);
nor I_31309 (I535151,I336005,I335987);
and I_31310 (I535168,I535151,I335984);
nor I_31311 (I535185,I535168,I336005);
not I_31312 (I535202,I336005);
and I_31313 (I535219,I535202,I335990);
nand I_31314 (I535236,I535219,I336002);
nor I_31315 (I535253,I535202,I535236);
DFFARX1 I_31316 (I535253,I2859,I535055,I535020,);
not I_31317 (I535284,I535236);
nand I_31318 (I535301,I535106,I535284);
nand I_31319 (I535032,I535168,I535284);
DFFARX1 I_31320 (I535202,I2859,I535055,I535047,);
not I_31321 (I535346,I335996);
nor I_31322 (I535363,I535346,I335990);
nor I_31323 (I535380,I535363,I535185);
DFFARX1 I_31324 (I535380,I2859,I535055,I535044,);
not I_31325 (I535411,I535363);
DFFARX1 I_31326 (I535411,I2859,I535055,I535437,);
not I_31327 (I535445,I535437);
nor I_31328 (I535041,I535445,I535363);
nor I_31329 (I535476,I535346,I335984);
and I_31330 (I535493,I535476,I335999);
or I_31331 (I535510,I535493,I335987);
DFFARX1 I_31332 (I535510,I2859,I535055,I535536,);
not I_31333 (I535544,I535536);
nand I_31334 (I535561,I535544,I535284);
not I_31335 (I535035,I535561);
nand I_31336 (I535029,I535561,I535301);
nand I_31337 (I535026,I535544,I535168);
not I_31338 (I535650,I2866);
DFFARX1 I_31339 (I91167,I2859,I535650,I535676,);
DFFARX1 I_31340 (I91170,I2859,I535650,I535693,);
not I_31341 (I535701,I535693);
nor I_31342 (I535618,I535676,I535701);
DFFARX1 I_31343 (I535701,I2859,I535650,I535633,);
nor I_31344 (I535746,I91176,I91170);
and I_31345 (I535763,I535746,I91173);
nor I_31346 (I535780,I535763,I91176);
not I_31347 (I535797,I91176);
and I_31348 (I535814,I535797,I91167);
nand I_31349 (I535831,I535814,I91185);
nor I_31350 (I535848,I535797,I535831);
DFFARX1 I_31351 (I535848,I2859,I535650,I535615,);
not I_31352 (I535879,I535831);
nand I_31353 (I535896,I535701,I535879);
nand I_31354 (I535627,I535763,I535879);
DFFARX1 I_31355 (I535797,I2859,I535650,I535642,);
not I_31356 (I535941,I91179);
nor I_31357 (I535958,I535941,I91167);
nor I_31358 (I535975,I535958,I535780);
DFFARX1 I_31359 (I535975,I2859,I535650,I535639,);
not I_31360 (I536006,I535958);
DFFARX1 I_31361 (I536006,I2859,I535650,I536032,);
not I_31362 (I536040,I536032);
nor I_31363 (I535636,I536040,I535958);
nor I_31364 (I536071,I535941,I91182);
and I_31365 (I536088,I536071,I91188);
or I_31366 (I536105,I536088,I91191);
DFFARX1 I_31367 (I536105,I2859,I535650,I536131,);
not I_31368 (I536139,I536131);
nand I_31369 (I536156,I536139,I535879);
not I_31370 (I535630,I536156);
nand I_31371 (I535624,I536156,I535896);
nand I_31372 (I535621,I536139,I535763);
not I_31373 (I536245,I2866);
DFFARX1 I_31374 (I72127,I2859,I536245,I536271,);
DFFARX1 I_31375 (I72130,I2859,I536245,I536288,);
not I_31376 (I536296,I536288);
nor I_31377 (I536213,I536271,I536296);
DFFARX1 I_31378 (I536296,I2859,I536245,I536228,);
nor I_31379 (I536341,I72136,I72130);
and I_31380 (I536358,I536341,I72133);
nor I_31381 (I536375,I536358,I72136);
not I_31382 (I536392,I72136);
and I_31383 (I536409,I536392,I72127);
nand I_31384 (I536426,I536409,I72145);
nor I_31385 (I536443,I536392,I536426);
DFFARX1 I_31386 (I536443,I2859,I536245,I536210,);
not I_31387 (I536474,I536426);
nand I_31388 (I536491,I536296,I536474);
nand I_31389 (I536222,I536358,I536474);
DFFARX1 I_31390 (I536392,I2859,I536245,I536237,);
not I_31391 (I536536,I72139);
nor I_31392 (I536553,I536536,I72127);
nor I_31393 (I536570,I536553,I536375);
DFFARX1 I_31394 (I536570,I2859,I536245,I536234,);
not I_31395 (I536601,I536553);
DFFARX1 I_31396 (I536601,I2859,I536245,I536627,);
not I_31397 (I536635,I536627);
nor I_31398 (I536231,I536635,I536553);
nor I_31399 (I536666,I536536,I72142);
and I_31400 (I536683,I536666,I72148);
or I_31401 (I536700,I536683,I72151);
DFFARX1 I_31402 (I536700,I2859,I536245,I536726,);
not I_31403 (I536734,I536726);
nand I_31404 (I536751,I536734,I536474);
not I_31405 (I536225,I536751);
nand I_31406 (I536219,I536751,I536491);
nand I_31407 (I536216,I536734,I536358);
not I_31408 (I536840,I2866);
DFFARX1 I_31409 (I165848,I2859,I536840,I536866,);
DFFARX1 I_31410 (I165854,I2859,I536840,I536883,);
not I_31411 (I536891,I536883);
nor I_31412 (I536808,I536866,I536891);
DFFARX1 I_31413 (I536891,I2859,I536840,I536823,);
nor I_31414 (I536936,I165863,I165848);
and I_31415 (I536953,I536936,I165875);
nor I_31416 (I536970,I536953,I165863);
not I_31417 (I536987,I165863);
and I_31418 (I537004,I536987,I165851);
nand I_31419 (I537021,I537004,I165872);
nor I_31420 (I537038,I536987,I537021);
DFFARX1 I_31421 (I537038,I2859,I536840,I536805,);
not I_31422 (I537069,I537021);
nand I_31423 (I537086,I536891,I537069);
nand I_31424 (I536817,I536953,I537069);
DFFARX1 I_31425 (I536987,I2859,I536840,I536832,);
not I_31426 (I537131,I165860);
nor I_31427 (I537148,I537131,I165851);
nor I_31428 (I537165,I537148,I536970);
DFFARX1 I_31429 (I537165,I2859,I536840,I536829,);
not I_31430 (I537196,I537148);
DFFARX1 I_31431 (I537196,I2859,I536840,I537222,);
not I_31432 (I537230,I537222);
nor I_31433 (I536826,I537230,I537148);
nor I_31434 (I537261,I537131,I165857);
and I_31435 (I537278,I537261,I165869);
or I_31436 (I537295,I537278,I165866);
DFFARX1 I_31437 (I537295,I2859,I536840,I537321,);
not I_31438 (I537329,I537321);
nand I_31439 (I537346,I537329,I537069);
not I_31440 (I536820,I537346);
nand I_31441 (I536814,I537346,I537086);
nand I_31442 (I536811,I537329,I536953);
not I_31443 (I537435,I2866);
DFFARX1 I_31444 (I25891,I2859,I537435,I537461,);
DFFARX1 I_31445 (I25879,I2859,I537435,I537478,);
not I_31446 (I537486,I537478);
nor I_31447 (I537403,I537461,I537486);
DFFARX1 I_31448 (I537486,I2859,I537435,I537418,);
nor I_31449 (I537531,I25870,I25894);
and I_31450 (I537548,I537531,I25873);
nor I_31451 (I537565,I537548,I25870);
not I_31452 (I537582,I25870);
and I_31453 (I537599,I537582,I25876);
nand I_31454 (I537616,I537599,I25888);
nor I_31455 (I537633,I537582,I537616);
DFFARX1 I_31456 (I537633,I2859,I537435,I537400,);
not I_31457 (I537664,I537616);
nand I_31458 (I537681,I537486,I537664);
nand I_31459 (I537412,I537548,I537664);
DFFARX1 I_31460 (I537582,I2859,I537435,I537427,);
not I_31461 (I537726,I25870);
nor I_31462 (I537743,I537726,I25876);
nor I_31463 (I537760,I537743,I537565);
DFFARX1 I_31464 (I537760,I2859,I537435,I537424,);
not I_31465 (I537791,I537743);
DFFARX1 I_31466 (I537791,I2859,I537435,I537817,);
not I_31467 (I537825,I537817);
nor I_31468 (I537421,I537825,I537743);
nor I_31469 (I537856,I537726,I25873);
and I_31470 (I537873,I537856,I25882);
or I_31471 (I537890,I537873,I25885);
DFFARX1 I_31472 (I537890,I2859,I537435,I537916,);
not I_31473 (I537924,I537916);
nand I_31474 (I537941,I537924,I537664);
not I_31475 (I537415,I537941);
nand I_31476 (I537409,I537941,I537681);
nand I_31477 (I537406,I537924,I537548);
not I_31478 (I538030,I2866);
DFFARX1 I_31479 (I274737,I2859,I538030,I538056,);
DFFARX1 I_31480 (I274719,I2859,I538030,I538073,);
not I_31481 (I538081,I538073);
nor I_31482 (I537998,I538056,I538081);
DFFARX1 I_31483 (I538081,I2859,I538030,I538013,);
nor I_31484 (I538126,I274725,I274728);
and I_31485 (I538143,I538126,I274716);
nor I_31486 (I538160,I538143,I274725);
not I_31487 (I538177,I274725);
and I_31488 (I538194,I538177,I274734);
nand I_31489 (I538211,I538194,I274722);
nor I_31490 (I538228,I538177,I538211);
DFFARX1 I_31491 (I538228,I2859,I538030,I537995,);
not I_31492 (I538259,I538211);
nand I_31493 (I538276,I538081,I538259);
nand I_31494 (I538007,I538143,I538259);
DFFARX1 I_31495 (I538177,I2859,I538030,I538022,);
not I_31496 (I538321,I274719);
nor I_31497 (I538338,I538321,I274734);
nor I_31498 (I538355,I538338,I538160);
DFFARX1 I_31499 (I538355,I2859,I538030,I538019,);
not I_31500 (I538386,I538338);
DFFARX1 I_31501 (I538386,I2859,I538030,I538412,);
not I_31502 (I538420,I538412);
nor I_31503 (I538016,I538420,I538338);
nor I_31504 (I538451,I538321,I274731);
and I_31505 (I538468,I538451,I274740);
or I_31506 (I538485,I538468,I274716);
DFFARX1 I_31507 (I538485,I2859,I538030,I538511,);
not I_31508 (I538519,I538511);
nand I_31509 (I538536,I538519,I538259);
not I_31510 (I538010,I538536);
nand I_31511 (I538004,I538536,I538276);
nand I_31512 (I538001,I538519,I538143);
not I_31513 (I538625,I2866);
DFFARX1 I_31514 (I402511,I2859,I538625,I538651,);
DFFARX1 I_31515 (I402529,I2859,I538625,I538668,);
not I_31516 (I538676,I538668);
nor I_31517 (I538593,I538651,I538676);
DFFARX1 I_31518 (I538676,I2859,I538625,I538608,);
nor I_31519 (I538721,I402508,I402520);
and I_31520 (I538738,I538721,I402505);
nor I_31521 (I538755,I538738,I402508);
not I_31522 (I538772,I402508);
and I_31523 (I538789,I538772,I402514);
nand I_31524 (I538806,I538789,I402526);
nor I_31525 (I538823,I538772,I538806);
DFFARX1 I_31526 (I538823,I2859,I538625,I538590,);
not I_31527 (I538854,I538806);
nand I_31528 (I538871,I538676,I538854);
nand I_31529 (I538602,I538738,I538854);
DFFARX1 I_31530 (I538772,I2859,I538625,I538617,);
not I_31531 (I538916,I402517);
nor I_31532 (I538933,I538916,I402514);
nor I_31533 (I538950,I538933,I538755);
DFFARX1 I_31534 (I538950,I2859,I538625,I538614,);
not I_31535 (I538981,I538933);
DFFARX1 I_31536 (I538981,I2859,I538625,I539007,);
not I_31537 (I539015,I539007);
nor I_31538 (I538611,I539015,I538933);
nor I_31539 (I539046,I538916,I402505);
and I_31540 (I539063,I539046,I402532);
or I_31541 (I539080,I539063,I402523);
DFFARX1 I_31542 (I539080,I2859,I538625,I539106,);
not I_31543 (I539114,I539106);
nand I_31544 (I539131,I539114,I538854);
not I_31545 (I538605,I539131);
nand I_31546 (I538599,I539131,I538871);
nand I_31547 (I538596,I539114,I538738);
not I_31548 (I539220,I2866);
DFFARX1 I_31549 (I437231,I2859,I539220,I539246,);
DFFARX1 I_31550 (I437222,I2859,I539220,I539263,);
not I_31551 (I539271,I539263);
nor I_31552 (I539188,I539246,I539271);
DFFARX1 I_31553 (I539271,I2859,I539220,I539203,);
nor I_31554 (I539316,I437228,I437237);
and I_31555 (I539333,I539316,I437240);
nor I_31556 (I539350,I539333,I437228);
not I_31557 (I539367,I437228);
and I_31558 (I539384,I539367,I437219);
nand I_31559 (I539401,I539384,I437225);
nor I_31560 (I539418,I539367,I539401);
DFFARX1 I_31561 (I539418,I2859,I539220,I539185,);
not I_31562 (I539449,I539401);
nand I_31563 (I539466,I539271,I539449);
nand I_31564 (I539197,I539333,I539449);
DFFARX1 I_31565 (I539367,I2859,I539220,I539212,);
not I_31566 (I539511,I437234);
nor I_31567 (I539528,I539511,I437219);
nor I_31568 (I539545,I539528,I539350);
DFFARX1 I_31569 (I539545,I2859,I539220,I539209,);
not I_31570 (I539576,I539528);
DFFARX1 I_31571 (I539576,I2859,I539220,I539602,);
not I_31572 (I539610,I539602);
nor I_31573 (I539206,I539610,I539528);
nor I_31574 (I539641,I539511,I437219);
and I_31575 (I539658,I539641,I437222);
or I_31576 (I539675,I539658,I437225);
DFFARX1 I_31577 (I539675,I2859,I539220,I539701,);
not I_31578 (I539709,I539701);
nand I_31579 (I539726,I539709,I539449);
not I_31580 (I539200,I539726);
nand I_31581 (I539194,I539726,I539466);
nand I_31582 (I539191,I539709,I539333);
not I_31583 (I539815,I2866);
DFFARX1 I_31584 (I62012,I2859,I539815,I539841,);
DFFARX1 I_31585 (I62015,I2859,I539815,I539858,);
not I_31586 (I539866,I539858);
nor I_31587 (I539783,I539841,I539866);
DFFARX1 I_31588 (I539866,I2859,I539815,I539798,);
nor I_31589 (I539911,I62021,I62015);
and I_31590 (I539928,I539911,I62018);
nor I_31591 (I539945,I539928,I62021);
not I_31592 (I539962,I62021);
and I_31593 (I539979,I539962,I62012);
nand I_31594 (I539996,I539979,I62030);
nor I_31595 (I540013,I539962,I539996);
DFFARX1 I_31596 (I540013,I2859,I539815,I539780,);
not I_31597 (I540044,I539996);
nand I_31598 (I540061,I539866,I540044);
nand I_31599 (I539792,I539928,I540044);
DFFARX1 I_31600 (I539962,I2859,I539815,I539807,);
not I_31601 (I540106,I62024);
nor I_31602 (I540123,I540106,I62012);
nor I_31603 (I540140,I540123,I539945);
DFFARX1 I_31604 (I540140,I2859,I539815,I539804,);
not I_31605 (I540171,I540123);
DFFARX1 I_31606 (I540171,I2859,I539815,I540197,);
not I_31607 (I540205,I540197);
nor I_31608 (I539801,I540205,I540123);
nor I_31609 (I540236,I540106,I62027);
and I_31610 (I540253,I540236,I62033);
or I_31611 (I540270,I540253,I62036);
DFFARX1 I_31612 (I540270,I2859,I539815,I540296,);
not I_31613 (I540304,I540296);
nand I_31614 (I540321,I540304,I540044);
not I_31615 (I539795,I540321);
nand I_31616 (I539789,I540321,I540061);
nand I_31617 (I539786,I540304,I539928);
not I_31618 (I540410,I2866);
DFFARX1 I_31619 (I124593,I2859,I540410,I540436,);
DFFARX1 I_31620 (I124587,I2859,I540410,I540453,);
not I_31621 (I540461,I540453);
nor I_31622 (I540378,I540436,I540461);
DFFARX1 I_31623 (I540461,I2859,I540410,I540393,);
nor I_31624 (I540506,I124575,I124596);
and I_31625 (I540523,I540506,I124590);
nor I_31626 (I540540,I540523,I124575);
not I_31627 (I540557,I124575);
and I_31628 (I540574,I540557,I124572);
nand I_31629 (I540591,I540574,I124584);
nor I_31630 (I540608,I540557,I540591);
DFFARX1 I_31631 (I540608,I2859,I540410,I540375,);
not I_31632 (I540639,I540591);
nand I_31633 (I540656,I540461,I540639);
nand I_31634 (I540387,I540523,I540639);
DFFARX1 I_31635 (I540557,I2859,I540410,I540402,);
not I_31636 (I540701,I124599);
nor I_31637 (I540718,I540701,I124572);
nor I_31638 (I540735,I540718,I540540);
DFFARX1 I_31639 (I540735,I2859,I540410,I540399,);
not I_31640 (I540766,I540718);
DFFARX1 I_31641 (I540766,I2859,I540410,I540792,);
not I_31642 (I540800,I540792);
nor I_31643 (I540396,I540800,I540718);
nor I_31644 (I540831,I540701,I124581);
and I_31645 (I540848,I540831,I124578);
or I_31646 (I540865,I540848,I124572);
DFFARX1 I_31647 (I540865,I2859,I540410,I540891,);
not I_31648 (I540899,I540891);
nand I_31649 (I540916,I540899,I540639);
not I_31650 (I540390,I540916);
nand I_31651 (I540384,I540916,I540656);
nand I_31652 (I540381,I540899,I540523);
not I_31653 (I541005,I2866);
DFFARX1 I_31654 (I289765,I2859,I541005,I541031,);
DFFARX1 I_31655 (I289747,I2859,I541005,I541048,);
not I_31656 (I541056,I541048);
nor I_31657 (I540973,I541031,I541056);
DFFARX1 I_31658 (I541056,I2859,I541005,I540988,);
nor I_31659 (I541101,I289753,I289756);
and I_31660 (I541118,I541101,I289744);
nor I_31661 (I541135,I541118,I289753);
not I_31662 (I541152,I289753);
and I_31663 (I541169,I541152,I289762);
nand I_31664 (I541186,I541169,I289750);
nor I_31665 (I541203,I541152,I541186);
DFFARX1 I_31666 (I541203,I2859,I541005,I540970,);
not I_31667 (I541234,I541186);
nand I_31668 (I541251,I541056,I541234);
nand I_31669 (I540982,I541118,I541234);
DFFARX1 I_31670 (I541152,I2859,I541005,I540997,);
not I_31671 (I541296,I289747);
nor I_31672 (I541313,I541296,I289762);
nor I_31673 (I541330,I541313,I541135);
DFFARX1 I_31674 (I541330,I2859,I541005,I540994,);
not I_31675 (I541361,I541313);
DFFARX1 I_31676 (I541361,I2859,I541005,I541387,);
not I_31677 (I541395,I541387);
nor I_31678 (I540991,I541395,I541313);
nor I_31679 (I541426,I541296,I289759);
and I_31680 (I541443,I541426,I289768);
or I_31681 (I541460,I541443,I289744);
DFFARX1 I_31682 (I541460,I2859,I541005,I541486,);
not I_31683 (I541494,I541486);
nand I_31684 (I541511,I541494,I541234);
not I_31685 (I540985,I541511);
nand I_31686 (I540979,I541511,I541251);
nand I_31687 (I540976,I541494,I541118);
not I_31688 (I541600,I2866);
DFFARX1 I_31689 (I236589,I2859,I541600,I541626,);
DFFARX1 I_31690 (I236583,I2859,I541600,I541643,);
not I_31691 (I541651,I541643);
nor I_31692 (I541568,I541626,I541651);
DFFARX1 I_31693 (I541651,I2859,I541600,I541583,);
nor I_31694 (I541696,I236580,I236571);
and I_31695 (I541713,I541696,I236568);
nor I_31696 (I541730,I541713,I236580);
not I_31697 (I541747,I236580);
and I_31698 (I541764,I541747,I236574);
nand I_31699 (I541781,I541764,I236586);
nor I_31700 (I541798,I541747,I541781);
DFFARX1 I_31701 (I541798,I2859,I541600,I541565,);
not I_31702 (I541829,I541781);
nand I_31703 (I541846,I541651,I541829);
nand I_31704 (I541577,I541713,I541829);
DFFARX1 I_31705 (I541747,I2859,I541600,I541592,);
not I_31706 (I541891,I236592);
nor I_31707 (I541908,I541891,I236574);
nor I_31708 (I541925,I541908,I541730);
DFFARX1 I_31709 (I541925,I2859,I541600,I541589,);
not I_31710 (I541956,I541908);
DFFARX1 I_31711 (I541956,I2859,I541600,I541982,);
not I_31712 (I541990,I541982);
nor I_31713 (I541586,I541990,I541908);
nor I_31714 (I542021,I541891,I236571);
and I_31715 (I542038,I542021,I236577);
or I_31716 (I542055,I542038,I236568);
DFFARX1 I_31717 (I542055,I2859,I541600,I542081,);
not I_31718 (I542089,I542081);
nand I_31719 (I542106,I542089,I541829);
not I_31720 (I541580,I542106);
nand I_31721 (I541574,I542106,I541846);
nand I_31722 (I541571,I542089,I541713);
not I_31723 (I542195,I2866);
DFFARX1 I_31724 (I332304,I2859,I542195,I542221,);
DFFARX1 I_31725 (I332301,I2859,I542195,I542238,);
not I_31726 (I542246,I542238);
nor I_31727 (I542163,I542221,I542246);
DFFARX1 I_31728 (I542246,I2859,I542195,I542178,);
nor I_31729 (I542291,I332316,I332298);
and I_31730 (I542308,I542291,I332295);
nor I_31731 (I542325,I542308,I332316);
not I_31732 (I542342,I332316);
and I_31733 (I542359,I542342,I332301);
nand I_31734 (I542376,I542359,I332313);
nor I_31735 (I542393,I542342,I542376);
DFFARX1 I_31736 (I542393,I2859,I542195,I542160,);
not I_31737 (I542424,I542376);
nand I_31738 (I542441,I542246,I542424);
nand I_31739 (I542172,I542308,I542424);
DFFARX1 I_31740 (I542342,I2859,I542195,I542187,);
not I_31741 (I542486,I332307);
nor I_31742 (I542503,I542486,I332301);
nor I_31743 (I542520,I542503,I542325);
DFFARX1 I_31744 (I542520,I2859,I542195,I542184,);
not I_31745 (I542551,I542503);
DFFARX1 I_31746 (I542551,I2859,I542195,I542577,);
not I_31747 (I542585,I542577);
nor I_31748 (I542181,I542585,I542503);
nor I_31749 (I542616,I542486,I332295);
and I_31750 (I542633,I542616,I332310);
or I_31751 (I542650,I542633,I332298);
DFFARX1 I_31752 (I542650,I2859,I542195,I542676,);
not I_31753 (I542684,I542676);
nand I_31754 (I542701,I542684,I542424);
not I_31755 (I542175,I542701);
nand I_31756 (I542169,I542701,I542441);
nand I_31757 (I542166,I542684,I542308);
not I_31758 (I542790,I2866);
DFFARX1 I_31759 (I172920,I2859,I542790,I542816,);
DFFARX1 I_31760 (I172926,I2859,I542790,I542833,);
not I_31761 (I542841,I542833);
nor I_31762 (I542758,I542816,I542841);
DFFARX1 I_31763 (I542841,I2859,I542790,I542773,);
nor I_31764 (I542886,I172935,I172920);
and I_31765 (I542903,I542886,I172947);
nor I_31766 (I542920,I542903,I172935);
not I_31767 (I542937,I172935);
and I_31768 (I542954,I542937,I172923);
nand I_31769 (I542971,I542954,I172944);
nor I_31770 (I542988,I542937,I542971);
DFFARX1 I_31771 (I542988,I2859,I542790,I542755,);
not I_31772 (I543019,I542971);
nand I_31773 (I543036,I542841,I543019);
nand I_31774 (I542767,I542903,I543019);
DFFARX1 I_31775 (I542937,I2859,I542790,I542782,);
not I_31776 (I543081,I172932);
nor I_31777 (I543098,I543081,I172923);
nor I_31778 (I543115,I543098,I542920);
DFFARX1 I_31779 (I543115,I2859,I542790,I542779,);
not I_31780 (I543146,I543098);
DFFARX1 I_31781 (I543146,I2859,I542790,I543172,);
not I_31782 (I543180,I543172);
nor I_31783 (I542776,I543180,I543098);
nor I_31784 (I543211,I543081,I172929);
and I_31785 (I543228,I543211,I172941);
or I_31786 (I543245,I543228,I172938);
DFFARX1 I_31787 (I543245,I2859,I542790,I543271,);
not I_31788 (I543279,I543271);
nand I_31789 (I543296,I543279,I543019);
not I_31790 (I542770,I543296);
nand I_31791 (I542764,I543296,I543036);
nand I_31792 (I542761,I543279,I542903);
not I_31793 (I543385,I2866);
DFFARX1 I_31794 (I110802,I2859,I543385,I543411,);
DFFARX1 I_31795 (I110805,I2859,I543385,I543428,);
not I_31796 (I543436,I543428);
nor I_31797 (I543353,I543411,I543436);
DFFARX1 I_31798 (I543436,I2859,I543385,I543368,);
nor I_31799 (I543481,I110811,I110805);
and I_31800 (I543498,I543481,I110808);
nor I_31801 (I543515,I543498,I110811);
not I_31802 (I543532,I110811);
and I_31803 (I543549,I543532,I110802);
nand I_31804 (I543566,I543549,I110820);
nor I_31805 (I543583,I543532,I543566);
DFFARX1 I_31806 (I543583,I2859,I543385,I543350,);
not I_31807 (I543614,I543566);
nand I_31808 (I543631,I543436,I543614);
nand I_31809 (I543362,I543498,I543614);
DFFARX1 I_31810 (I543532,I2859,I543385,I543377,);
not I_31811 (I543676,I110814);
nor I_31812 (I543693,I543676,I110802);
nor I_31813 (I543710,I543693,I543515);
DFFARX1 I_31814 (I543710,I2859,I543385,I543374,);
not I_31815 (I543741,I543693);
DFFARX1 I_31816 (I543741,I2859,I543385,I543767,);
not I_31817 (I543775,I543767);
nor I_31818 (I543371,I543775,I543693);
nor I_31819 (I543806,I543676,I110817);
and I_31820 (I543823,I543806,I110823);
or I_31821 (I543840,I543823,I110826);
DFFARX1 I_31822 (I543840,I2859,I543385,I543866,);
not I_31823 (I543874,I543866);
nand I_31824 (I543891,I543874,I543614);
not I_31825 (I543365,I543891);
nand I_31826 (I543359,I543891,I543631);
nand I_31827 (I543356,I543874,I543498);
not I_31828 (I543980,I2866);
DFFARX1 I_31829 (I268379,I2859,I543980,I544006,);
DFFARX1 I_31830 (I268361,I2859,I543980,I544023,);
not I_31831 (I544031,I544023);
nor I_31832 (I543948,I544006,I544031);
DFFARX1 I_31833 (I544031,I2859,I543980,I543963,);
nor I_31834 (I544076,I268367,I268370);
and I_31835 (I544093,I544076,I268358);
nor I_31836 (I544110,I544093,I268367);
not I_31837 (I544127,I268367);
and I_31838 (I544144,I544127,I268376);
nand I_31839 (I544161,I544144,I268364);
nor I_31840 (I544178,I544127,I544161);
DFFARX1 I_31841 (I544178,I2859,I543980,I543945,);
not I_31842 (I544209,I544161);
nand I_31843 (I544226,I544031,I544209);
nand I_31844 (I543957,I544093,I544209);
DFFARX1 I_31845 (I544127,I2859,I543980,I543972,);
not I_31846 (I544271,I268361);
nor I_31847 (I544288,I544271,I268376);
nor I_31848 (I544305,I544288,I544110);
DFFARX1 I_31849 (I544305,I2859,I543980,I543969,);
not I_31850 (I544336,I544288);
DFFARX1 I_31851 (I544336,I2859,I543980,I544362,);
not I_31852 (I544370,I544362);
nor I_31853 (I543966,I544370,I544288);
nor I_31854 (I544401,I544271,I268373);
and I_31855 (I544418,I544401,I268382);
or I_31856 (I544435,I544418,I268358);
DFFARX1 I_31857 (I544435,I2859,I543980,I544461,);
not I_31858 (I544469,I544461);
nand I_31859 (I544486,I544469,I544209);
not I_31860 (I543960,I544486);
nand I_31861 (I543954,I544486,I544226);
nand I_31862 (I543951,I544469,I544093);
not I_31863 (I544575,I2866);
DFFARX1 I_31864 (I440061,I2859,I544575,I544601,);
DFFARX1 I_31865 (I440073,I2859,I544575,I544618,);
not I_31866 (I544626,I544618);
nor I_31867 (I544543,I544601,I544626);
DFFARX1 I_31868 (I544626,I2859,I544575,I544558,);
nor I_31869 (I544671,I440070,I440064);
and I_31870 (I544688,I544671,I440058);
nor I_31871 (I544705,I544688,I440070);
not I_31872 (I544722,I440070);
and I_31873 (I544739,I544722,I440067);
nand I_31874 (I544756,I544739,I440058);
nor I_31875 (I544773,I544722,I544756);
DFFARX1 I_31876 (I544773,I2859,I544575,I544540,);
not I_31877 (I544804,I544756);
nand I_31878 (I544821,I544626,I544804);
nand I_31879 (I544552,I544688,I544804);
DFFARX1 I_31880 (I544722,I2859,I544575,I544567,);
not I_31881 (I544866,I440082);
nor I_31882 (I544883,I544866,I440067);
nor I_31883 (I544900,I544883,I544705);
DFFARX1 I_31884 (I544900,I2859,I544575,I544564,);
not I_31885 (I544931,I544883);
DFFARX1 I_31886 (I544931,I2859,I544575,I544957,);
not I_31887 (I544965,I544957);
nor I_31888 (I544561,I544965,I544883);
nor I_31889 (I544996,I544866,I440076);
and I_31890 (I545013,I544996,I440079);
or I_31891 (I545030,I545013,I440061);
DFFARX1 I_31892 (I545030,I2859,I544575,I545056,);
not I_31893 (I545064,I545056);
nand I_31894 (I545081,I545064,I544804);
not I_31895 (I544555,I545081);
nand I_31896 (I544549,I545081,I544821);
nand I_31897 (I544546,I545064,I544688);
not I_31898 (I545170,I2866);
DFFARX1 I_31899 (I482255,I2859,I545170,I545196,);
DFFARX1 I_31900 (I482267,I2859,I545170,I545213,);
not I_31901 (I545221,I545213);
nor I_31902 (I545138,I545196,I545221);
DFFARX1 I_31903 (I545221,I2859,I545170,I545153,);
nor I_31904 (I545266,I482264,I482258);
and I_31905 (I545283,I545266,I482252);
nor I_31906 (I545300,I545283,I482264);
not I_31907 (I545317,I482264);
and I_31908 (I545334,I545317,I482261);
nand I_31909 (I545351,I545334,I482252);
nor I_31910 (I545368,I545317,I545351);
DFFARX1 I_31911 (I545368,I2859,I545170,I545135,);
not I_31912 (I545399,I545351);
nand I_31913 (I545416,I545221,I545399);
nand I_31914 (I545147,I545283,I545399);
DFFARX1 I_31915 (I545317,I2859,I545170,I545162,);
not I_31916 (I545461,I482276);
nor I_31917 (I545478,I545461,I482261);
nor I_31918 (I545495,I545478,I545300);
DFFARX1 I_31919 (I545495,I2859,I545170,I545159,);
not I_31920 (I545526,I545478);
DFFARX1 I_31921 (I545526,I2859,I545170,I545552,);
not I_31922 (I545560,I545552);
nor I_31923 (I545156,I545560,I545478);
nor I_31924 (I545591,I545461,I482270);
and I_31925 (I545608,I545591,I482273);
or I_31926 (I545625,I545608,I482255);
DFFARX1 I_31927 (I545625,I2859,I545170,I545651,);
not I_31928 (I545659,I545651);
nand I_31929 (I545676,I545659,I545399);
not I_31930 (I545150,I545676);
nand I_31931 (I545144,I545676,I545416);
nand I_31932 (I545141,I545659,I545283);
not I_31933 (I545765,I2866);
DFFARX1 I_31934 (I490925,I2859,I545765,I545791,);
DFFARX1 I_31935 (I490937,I2859,I545765,I545808,);
not I_31936 (I545816,I545808);
nor I_31937 (I545733,I545791,I545816);
DFFARX1 I_31938 (I545816,I2859,I545765,I545748,);
nor I_31939 (I545861,I490934,I490928);
and I_31940 (I545878,I545861,I490922);
nor I_31941 (I545895,I545878,I490934);
not I_31942 (I545912,I490934);
and I_31943 (I545929,I545912,I490931);
nand I_31944 (I545946,I545929,I490922);
nor I_31945 (I545963,I545912,I545946);
DFFARX1 I_31946 (I545963,I2859,I545765,I545730,);
not I_31947 (I545994,I545946);
nand I_31948 (I546011,I545816,I545994);
nand I_31949 (I545742,I545878,I545994);
DFFARX1 I_31950 (I545912,I2859,I545765,I545757,);
not I_31951 (I546056,I490946);
nor I_31952 (I546073,I546056,I490931);
nor I_31953 (I546090,I546073,I545895);
DFFARX1 I_31954 (I546090,I2859,I545765,I545754,);
not I_31955 (I546121,I546073);
DFFARX1 I_31956 (I546121,I2859,I545765,I546147,);
not I_31957 (I546155,I546147);
nor I_31958 (I545751,I546155,I546073);
nor I_31959 (I546186,I546056,I490940);
and I_31960 (I546203,I546186,I490943);
or I_31961 (I546220,I546203,I490925);
DFFARX1 I_31962 (I546220,I2859,I545765,I546246,);
not I_31963 (I546254,I546246);
nand I_31964 (I546271,I546254,I545994);
not I_31965 (I545745,I546271);
nand I_31966 (I545739,I546271,I546011);
nand I_31967 (I545736,I546254,I545878);
not I_31968 (I546360,I2866);
DFFARX1 I_31969 (I283985,I2859,I546360,I546386,);
DFFARX1 I_31970 (I283967,I2859,I546360,I546403,);
not I_31971 (I546411,I546403);
nor I_31972 (I546328,I546386,I546411);
DFFARX1 I_31973 (I546411,I2859,I546360,I546343,);
nor I_31974 (I546456,I283973,I283976);
and I_31975 (I546473,I546456,I283964);
nor I_31976 (I546490,I546473,I283973);
not I_31977 (I546507,I283973);
and I_31978 (I546524,I546507,I283982);
nand I_31979 (I546541,I546524,I283970);
nor I_31980 (I546558,I546507,I546541);
DFFARX1 I_31981 (I546558,I2859,I546360,I546325,);
not I_31982 (I546589,I546541);
nand I_31983 (I546606,I546411,I546589);
nand I_31984 (I546337,I546473,I546589);
DFFARX1 I_31985 (I546507,I2859,I546360,I546352,);
not I_31986 (I546651,I283967);
nor I_31987 (I546668,I546651,I283982);
nor I_31988 (I546685,I546668,I546490);
DFFARX1 I_31989 (I546685,I2859,I546360,I546349,);
not I_31990 (I546716,I546668);
DFFARX1 I_31991 (I546716,I2859,I546360,I546742,);
not I_31992 (I546750,I546742);
nor I_31993 (I546346,I546750,I546668);
nor I_31994 (I546781,I546651,I283979);
and I_31995 (I546798,I546781,I283988);
or I_31996 (I546815,I546798,I283964);
DFFARX1 I_31997 (I546815,I2859,I546360,I546841,);
not I_31998 (I546849,I546841);
nand I_31999 (I546866,I546849,I546589);
not I_32000 (I546340,I546866);
nand I_32001 (I546334,I546866,I546606);
nand I_32002 (I546331,I546849,I546473);
not I_32003 (I546955,I2866);
DFFARX1 I_32004 (I290921,I2859,I546955,I546981,);
DFFARX1 I_32005 (I290903,I2859,I546955,I546998,);
not I_32006 (I547006,I546998);
nor I_32007 (I546923,I546981,I547006);
DFFARX1 I_32008 (I547006,I2859,I546955,I546938,);
nor I_32009 (I547051,I290909,I290912);
and I_32010 (I547068,I547051,I290900);
nor I_32011 (I547085,I547068,I290909);
not I_32012 (I547102,I290909);
and I_32013 (I547119,I547102,I290918);
nand I_32014 (I547136,I547119,I290906);
nor I_32015 (I547153,I547102,I547136);
DFFARX1 I_32016 (I547153,I2859,I546955,I546920,);
not I_32017 (I547184,I547136);
nand I_32018 (I547201,I547006,I547184);
nand I_32019 (I546932,I547068,I547184);
DFFARX1 I_32020 (I547102,I2859,I546955,I546947,);
not I_32021 (I547246,I290903);
nor I_32022 (I547263,I547246,I290918);
nor I_32023 (I547280,I547263,I547085);
DFFARX1 I_32024 (I547280,I2859,I546955,I546944,);
not I_32025 (I547311,I547263);
DFFARX1 I_32026 (I547311,I2859,I546955,I547337,);
not I_32027 (I547345,I547337);
nor I_32028 (I546941,I547345,I547263);
nor I_32029 (I547376,I547246,I290915);
and I_32030 (I547393,I547376,I290924);
or I_32031 (I547410,I547393,I290900);
DFFARX1 I_32032 (I547410,I2859,I546955,I547436,);
not I_32033 (I547444,I547436);
nand I_32034 (I547461,I547444,I547184);
not I_32035 (I546935,I547461);
nand I_32036 (I546929,I547461,I547201);
nand I_32037 (I546926,I547444,I547068);
not I_32038 (I547550,I2866);
DFFARX1 I_32039 (I31688,I2859,I547550,I547576,);
DFFARX1 I_32040 (I31676,I2859,I547550,I547593,);
not I_32041 (I547601,I547593);
nor I_32042 (I547518,I547576,I547601);
DFFARX1 I_32043 (I547601,I2859,I547550,I547533,);
nor I_32044 (I547646,I31667,I31691);
and I_32045 (I547663,I547646,I31670);
nor I_32046 (I547680,I547663,I31667);
not I_32047 (I547697,I31667);
and I_32048 (I547714,I547697,I31673);
nand I_32049 (I547731,I547714,I31685);
nor I_32050 (I547748,I547697,I547731);
DFFARX1 I_32051 (I547748,I2859,I547550,I547515,);
not I_32052 (I547779,I547731);
nand I_32053 (I547796,I547601,I547779);
nand I_32054 (I547527,I547663,I547779);
DFFARX1 I_32055 (I547697,I2859,I547550,I547542,);
not I_32056 (I547841,I31667);
nor I_32057 (I547858,I547841,I31673);
nor I_32058 (I547875,I547858,I547680);
DFFARX1 I_32059 (I547875,I2859,I547550,I547539,);
not I_32060 (I547906,I547858);
DFFARX1 I_32061 (I547906,I2859,I547550,I547932,);
not I_32062 (I547940,I547932);
nor I_32063 (I547536,I547940,I547858);
nor I_32064 (I547971,I547841,I31670);
and I_32065 (I547988,I547971,I31679);
or I_32066 (I548005,I547988,I31682);
DFFARX1 I_32067 (I548005,I2859,I547550,I548031,);
not I_32068 (I548039,I548031);
nand I_32069 (I548056,I548039,I547779);
not I_32070 (I547530,I548056);
nand I_32071 (I547524,I548056,I547796);
nand I_32072 (I547521,I548039,I547663);
not I_32073 (I548145,I2866);
DFFARX1 I_32074 (I266067,I2859,I548145,I548171,);
DFFARX1 I_32075 (I266049,I2859,I548145,I548188,);
not I_32076 (I548196,I548188);
nor I_32077 (I548113,I548171,I548196);
DFFARX1 I_32078 (I548196,I2859,I548145,I548128,);
nor I_32079 (I548241,I266055,I266058);
and I_32080 (I548258,I548241,I266046);
nor I_32081 (I548275,I548258,I266055);
not I_32082 (I548292,I266055);
and I_32083 (I548309,I548292,I266064);
nand I_32084 (I548326,I548309,I266052);
nor I_32085 (I548343,I548292,I548326);
DFFARX1 I_32086 (I548343,I2859,I548145,I548110,);
not I_32087 (I548374,I548326);
nand I_32088 (I548391,I548196,I548374);
nand I_32089 (I548122,I548258,I548374);
DFFARX1 I_32090 (I548292,I2859,I548145,I548137,);
not I_32091 (I548436,I266049);
nor I_32092 (I548453,I548436,I266064);
nor I_32093 (I548470,I548453,I548275);
DFFARX1 I_32094 (I548470,I2859,I548145,I548134,);
not I_32095 (I548501,I548453);
DFFARX1 I_32096 (I548501,I2859,I548145,I548527,);
not I_32097 (I548535,I548527);
nor I_32098 (I548131,I548535,I548453);
nor I_32099 (I548566,I548436,I266061);
and I_32100 (I548583,I548566,I266070);
or I_32101 (I548600,I548583,I266046);
DFFARX1 I_32102 (I548600,I2859,I548145,I548626,);
not I_32103 (I548634,I548626);
nand I_32104 (I548651,I548634,I548374);
not I_32105 (I548125,I548651);
nand I_32106 (I548119,I548651,I548391);
nand I_32107 (I548116,I548634,I548258);
not I_32108 (I548740,I2866);
DFFARX1 I_32109 (I424889,I2859,I548740,I548766,);
DFFARX1 I_32110 (I424880,I2859,I548740,I548783,);
not I_32111 (I548791,I548783);
nor I_32112 (I548708,I548766,I548791);
DFFARX1 I_32113 (I548791,I2859,I548740,I548723,);
nor I_32114 (I548836,I424886,I424895);
and I_32115 (I548853,I548836,I424898);
nor I_32116 (I548870,I548853,I424886);
not I_32117 (I548887,I424886);
and I_32118 (I548904,I548887,I424877);
nand I_32119 (I548921,I548904,I424883);
nor I_32120 (I548938,I548887,I548921);
DFFARX1 I_32121 (I548938,I2859,I548740,I548705,);
not I_32122 (I548969,I548921);
nand I_32123 (I548986,I548791,I548969);
nand I_32124 (I548717,I548853,I548969);
DFFARX1 I_32125 (I548887,I2859,I548740,I548732,);
not I_32126 (I549031,I424892);
nor I_32127 (I549048,I549031,I424877);
nor I_32128 (I549065,I549048,I548870);
DFFARX1 I_32129 (I549065,I2859,I548740,I548729,);
not I_32130 (I549096,I549048);
DFFARX1 I_32131 (I549096,I2859,I548740,I549122,);
not I_32132 (I549130,I549122);
nor I_32133 (I548726,I549130,I549048);
nor I_32134 (I549161,I549031,I424877);
and I_32135 (I549178,I549161,I424880);
or I_32136 (I549195,I549178,I424883);
DFFARX1 I_32137 (I549195,I2859,I548740,I549221,);
not I_32138 (I549229,I549221);
nand I_32139 (I549246,I549229,I548969);
not I_32140 (I548720,I549246);
nand I_32141 (I548714,I549246,I548986);
nand I_32142 (I548711,I549229,I548853);
not I_32143 (I549335,I2866);
DFFARX1 I_32144 (I20094,I2859,I549335,I549361,);
DFFARX1 I_32145 (I20082,I2859,I549335,I549378,);
not I_32146 (I549386,I549378);
nor I_32147 (I549303,I549361,I549386);
DFFARX1 I_32148 (I549386,I2859,I549335,I549318,);
nor I_32149 (I549431,I20073,I20097);
and I_32150 (I549448,I549431,I20076);
nor I_32151 (I549465,I549448,I20073);
not I_32152 (I549482,I20073);
and I_32153 (I549499,I549482,I20079);
nand I_32154 (I549516,I549499,I20091);
nor I_32155 (I549533,I549482,I549516);
DFFARX1 I_32156 (I549533,I2859,I549335,I549300,);
not I_32157 (I549564,I549516);
nand I_32158 (I549581,I549386,I549564);
nand I_32159 (I549312,I549448,I549564);
DFFARX1 I_32160 (I549482,I2859,I549335,I549327,);
not I_32161 (I549626,I20073);
nor I_32162 (I549643,I549626,I20079);
nor I_32163 (I549660,I549643,I549465);
DFFARX1 I_32164 (I549660,I2859,I549335,I549324,);
not I_32165 (I549691,I549643);
DFFARX1 I_32166 (I549691,I2859,I549335,I549717,);
not I_32167 (I549725,I549717);
nor I_32168 (I549321,I549725,I549643);
nor I_32169 (I549756,I549626,I20076);
and I_32170 (I549773,I549756,I20085);
or I_32171 (I549790,I549773,I20088);
DFFARX1 I_32172 (I549790,I2859,I549335,I549816,);
not I_32173 (I549824,I549816);
nand I_32174 (I549841,I549824,I549564);
not I_32175 (I549315,I549841);
nand I_32176 (I549309,I549841,I549581);
nand I_32177 (I549306,I549824,I549448);
not I_32178 (I549930,I2866);
DFFARX1 I_32179 (I117215,I2859,I549930,I549956,);
DFFARX1 I_32180 (I117209,I2859,I549930,I549973,);
not I_32181 (I549981,I549973);
nor I_32182 (I549898,I549956,I549981);
DFFARX1 I_32183 (I549981,I2859,I549930,I549913,);
nor I_32184 (I550026,I117197,I117218);
and I_32185 (I550043,I550026,I117212);
nor I_32186 (I550060,I550043,I117197);
not I_32187 (I550077,I117197);
and I_32188 (I550094,I550077,I117194);
nand I_32189 (I550111,I550094,I117206);
nor I_32190 (I550128,I550077,I550111);
DFFARX1 I_32191 (I550128,I2859,I549930,I549895,);
not I_32192 (I550159,I550111);
nand I_32193 (I550176,I549981,I550159);
nand I_32194 (I549907,I550043,I550159);
DFFARX1 I_32195 (I550077,I2859,I549930,I549922,);
not I_32196 (I550221,I117221);
nor I_32197 (I550238,I550221,I117194);
nor I_32198 (I550255,I550238,I550060);
DFFARX1 I_32199 (I550255,I2859,I549930,I549919,);
not I_32200 (I550286,I550238);
DFFARX1 I_32201 (I550286,I2859,I549930,I550312,);
not I_32202 (I550320,I550312);
nor I_32203 (I549916,I550320,I550238);
nor I_32204 (I550351,I550221,I117203);
and I_32205 (I550368,I550351,I117200);
or I_32206 (I550385,I550368,I117194);
DFFARX1 I_32207 (I550385,I2859,I549930,I550411,);
not I_32208 (I550419,I550411);
nand I_32209 (I550436,I550419,I550159);
not I_32210 (I549910,I550436);
nand I_32211 (I549904,I550436,I550176);
nand I_32212 (I549901,I550419,I550043);
not I_32213 (I550525,I2866);
DFFARX1 I_32214 (I337047,I2859,I550525,I550551,);
DFFARX1 I_32215 (I337044,I2859,I550525,I550568,);
not I_32216 (I550576,I550568);
nor I_32217 (I550493,I550551,I550576);
DFFARX1 I_32218 (I550576,I2859,I550525,I550508,);
nor I_32219 (I550621,I337059,I337041);
and I_32220 (I550638,I550621,I337038);
nor I_32221 (I550655,I550638,I337059);
not I_32222 (I550672,I337059);
and I_32223 (I550689,I550672,I337044);
nand I_32224 (I550706,I550689,I337056);
nor I_32225 (I550723,I550672,I550706);
DFFARX1 I_32226 (I550723,I2859,I550525,I550490,);
not I_32227 (I550754,I550706);
nand I_32228 (I550771,I550576,I550754);
nand I_32229 (I550502,I550638,I550754);
DFFARX1 I_32230 (I550672,I2859,I550525,I550517,);
not I_32231 (I550816,I337050);
nor I_32232 (I550833,I550816,I337044);
nor I_32233 (I550850,I550833,I550655);
DFFARX1 I_32234 (I550850,I2859,I550525,I550514,);
not I_32235 (I550881,I550833);
DFFARX1 I_32236 (I550881,I2859,I550525,I550907,);
not I_32237 (I550915,I550907);
nor I_32238 (I550511,I550915,I550833);
nor I_32239 (I550946,I550816,I337038);
and I_32240 (I550963,I550946,I337053);
or I_32241 (I550980,I550963,I337041);
DFFARX1 I_32242 (I550980,I2859,I550525,I551006,);
not I_32243 (I551014,I551006);
nand I_32244 (I551031,I551014,I550754);
not I_32245 (I550505,I551031);
nand I_32246 (I550499,I551031,I550771);
nand I_32247 (I550496,I551014,I550638);
not I_32248 (I551120,I2866);
DFFARX1 I_32249 (I524702,I2859,I551120,I551146,);
DFFARX1 I_32250 (I524693,I2859,I551120,I551163,);
not I_32251 (I551171,I551163);
nor I_32252 (I551088,I551146,I551171);
DFFARX1 I_32253 (I551171,I2859,I551120,I551103,);
nor I_32254 (I551216,I524684,I524699);
and I_32255 (I551233,I551216,I524687);
nor I_32256 (I551250,I551233,I524684);
not I_32257 (I551267,I524684);
and I_32258 (I551284,I551267,I524690);
nand I_32259 (I551301,I551284,I524708);
nor I_32260 (I551318,I551267,I551301);
DFFARX1 I_32261 (I551318,I2859,I551120,I551085,);
not I_32262 (I551349,I551301);
nand I_32263 (I551366,I551171,I551349);
nand I_32264 (I551097,I551233,I551349);
DFFARX1 I_32265 (I551267,I2859,I551120,I551112,);
not I_32266 (I551411,I524684);
nor I_32267 (I551428,I551411,I524690);
nor I_32268 (I551445,I551428,I551250);
DFFARX1 I_32269 (I551445,I2859,I551120,I551109,);
not I_32270 (I551476,I551428);
DFFARX1 I_32271 (I551476,I2859,I551120,I551502,);
not I_32272 (I551510,I551502);
nor I_32273 (I551106,I551510,I551428);
nor I_32274 (I551541,I551411,I524687);
and I_32275 (I551558,I551541,I524696);
or I_32276 (I551575,I551558,I524705);
DFFARX1 I_32277 (I551575,I2859,I551120,I551601,);
not I_32278 (I551609,I551601);
nand I_32279 (I551626,I551609,I551349);
not I_32280 (I551100,I551626);
nand I_32281 (I551094,I551626,I551366);
nand I_32282 (I551091,I551609,I551233);
not I_32283 (I551715,I2866);
DFFARX1 I_32284 (I533330,I2859,I551715,I551741,);
DFFARX1 I_32285 (I533315,I2859,I551715,I551758,);
not I_32286 (I551766,I551758);
nor I_32287 (I551683,I551741,I551766);
DFFARX1 I_32288 (I551766,I2859,I551715,I551698,);
nor I_32289 (I551811,I533312,I533321);
and I_32290 (I551828,I551811,I533327);
nor I_32291 (I551845,I551828,I533312);
not I_32292 (I551862,I533312);
and I_32293 (I551879,I551862,I533309);
nand I_32294 (I551896,I551879,I533303);
nor I_32295 (I551913,I551862,I551896);
DFFARX1 I_32296 (I551913,I2859,I551715,I551680,);
not I_32297 (I551944,I551896);
nand I_32298 (I551961,I551766,I551944);
nand I_32299 (I551692,I551828,I551944);
DFFARX1 I_32300 (I551862,I2859,I551715,I551707,);
not I_32301 (I552006,I533303);
nor I_32302 (I552023,I552006,I533309);
nor I_32303 (I552040,I552023,I551845);
DFFARX1 I_32304 (I552040,I2859,I551715,I551704,);
not I_32305 (I552071,I552023);
DFFARX1 I_32306 (I552071,I2859,I551715,I552097,);
not I_32307 (I552105,I552097);
nor I_32308 (I551701,I552105,I552023);
nor I_32309 (I552136,I552006,I533318);
and I_32310 (I552153,I552136,I533324);
or I_32311 (I552170,I552153,I533306);
DFFARX1 I_32312 (I552170,I2859,I551715,I552196,);
not I_32313 (I552204,I552196);
nand I_32314 (I552221,I552204,I551944);
not I_32315 (I551695,I552221);
nand I_32316 (I551689,I552221,I551961);
nand I_32317 (I551686,I552204,I551828);
not I_32318 (I552310,I2866);
DFFARX1 I_32319 (I477631,I2859,I552310,I552336,);
DFFARX1 I_32320 (I477643,I2859,I552310,I552353,);
not I_32321 (I552361,I552353);
nor I_32322 (I552278,I552336,I552361);
DFFARX1 I_32323 (I552361,I2859,I552310,I552293,);
nor I_32324 (I552406,I477640,I477634);
and I_32325 (I552423,I552406,I477628);
nor I_32326 (I552440,I552423,I477640);
not I_32327 (I552457,I477640);
and I_32328 (I552474,I552457,I477637);
nand I_32329 (I552491,I552474,I477628);
nor I_32330 (I552508,I552457,I552491);
DFFARX1 I_32331 (I552508,I2859,I552310,I552275,);
not I_32332 (I552539,I552491);
nand I_32333 (I552556,I552361,I552539);
nand I_32334 (I552287,I552423,I552539);
DFFARX1 I_32335 (I552457,I2859,I552310,I552302,);
not I_32336 (I552601,I477652);
nor I_32337 (I552618,I552601,I477637);
nor I_32338 (I552635,I552618,I552440);
DFFARX1 I_32339 (I552635,I2859,I552310,I552299,);
not I_32340 (I552666,I552618);
DFFARX1 I_32341 (I552666,I2859,I552310,I552692,);
not I_32342 (I552700,I552692);
nor I_32343 (I552296,I552700,I552618);
nor I_32344 (I552731,I552601,I477646);
and I_32345 (I552748,I552731,I477649);
or I_32346 (I552765,I552748,I477631);
DFFARX1 I_32347 (I552765,I2859,I552310,I552791,);
not I_32348 (I552799,I552791);
nand I_32349 (I552816,I552799,I552539);
not I_32350 (I552290,I552816);
nand I_32351 (I552284,I552816,I552556);
nand I_32352 (I552281,I552799,I552423);
not I_32353 (I552905,I2866);
DFFARX1 I_32354 (I57252,I2859,I552905,I552931,);
DFFARX1 I_32355 (I57255,I2859,I552905,I552948,);
not I_32356 (I552956,I552948);
nor I_32357 (I552873,I552931,I552956);
DFFARX1 I_32358 (I552956,I2859,I552905,I552888,);
nor I_32359 (I553001,I57261,I57255);
and I_32360 (I553018,I553001,I57258);
nor I_32361 (I553035,I553018,I57261);
not I_32362 (I553052,I57261);
and I_32363 (I553069,I553052,I57252);
nand I_32364 (I553086,I553069,I57270);
nor I_32365 (I553103,I553052,I553086);
DFFARX1 I_32366 (I553103,I2859,I552905,I552870,);
not I_32367 (I553134,I553086);
nand I_32368 (I553151,I552956,I553134);
nand I_32369 (I552882,I553018,I553134);
DFFARX1 I_32370 (I553052,I2859,I552905,I552897,);
not I_32371 (I553196,I57264);
nor I_32372 (I553213,I553196,I57252);
nor I_32373 (I553230,I553213,I553035);
DFFARX1 I_32374 (I553230,I2859,I552905,I552894,);
not I_32375 (I553261,I553213);
DFFARX1 I_32376 (I553261,I2859,I552905,I553287,);
not I_32377 (I553295,I553287);
nor I_32378 (I552891,I553295,I553213);
nor I_32379 (I553326,I553196,I57267);
and I_32380 (I553343,I553326,I57273);
or I_32381 (I553360,I553343,I57276);
DFFARX1 I_32382 (I553360,I2859,I552905,I553386,);
not I_32383 (I553394,I553386);
nand I_32384 (I553411,I553394,I553134);
not I_32385 (I552885,I553411);
nand I_32386 (I552879,I553411,I553151);
nand I_32387 (I552876,I553394,I553018);
not I_32388 (I553500,I2866);
DFFARX1 I_32389 (I245259,I2859,I553500,I553526,);
DFFARX1 I_32390 (I245253,I2859,I553500,I553543,);
not I_32391 (I553551,I553543);
nor I_32392 (I553468,I553526,I553551);
DFFARX1 I_32393 (I553551,I2859,I553500,I553483,);
nor I_32394 (I553596,I245250,I245241);
and I_32395 (I553613,I553596,I245238);
nor I_32396 (I553630,I553613,I245250);
not I_32397 (I553647,I245250);
and I_32398 (I553664,I553647,I245244);
nand I_32399 (I553681,I553664,I245256);
nor I_32400 (I553698,I553647,I553681);
DFFARX1 I_32401 (I553698,I2859,I553500,I553465,);
not I_32402 (I553729,I553681);
nand I_32403 (I553746,I553551,I553729);
nand I_32404 (I553477,I553613,I553729);
DFFARX1 I_32405 (I553647,I2859,I553500,I553492,);
not I_32406 (I553791,I245262);
nor I_32407 (I553808,I553791,I245244);
nor I_32408 (I553825,I553808,I553630);
DFFARX1 I_32409 (I553825,I2859,I553500,I553489,);
not I_32410 (I553856,I553808);
DFFARX1 I_32411 (I553856,I2859,I553500,I553882,);
not I_32412 (I553890,I553882);
nor I_32413 (I553486,I553890,I553808);
nor I_32414 (I553921,I553791,I245241);
and I_32415 (I553938,I553921,I245247);
or I_32416 (I553955,I553938,I245238);
DFFARX1 I_32417 (I553955,I2859,I553500,I553981,);
not I_32418 (I553989,I553981);
nand I_32419 (I554006,I553989,I553729);
not I_32420 (I553480,I554006);
nand I_32421 (I553474,I554006,I553746);
nand I_32422 (I553471,I553989,I553613);
not I_32423 (I554095,I2866);
DFFARX1 I_32424 (I417035,I2859,I554095,I554121,);
DFFARX1 I_32425 (I417026,I2859,I554095,I554138,);
not I_32426 (I554146,I554138);
nor I_32427 (I554063,I554121,I554146);
DFFARX1 I_32428 (I554146,I2859,I554095,I554078,);
nor I_32429 (I554191,I417032,I417041);
and I_32430 (I554208,I554191,I417044);
nor I_32431 (I554225,I554208,I417032);
not I_32432 (I554242,I417032);
and I_32433 (I554259,I554242,I417023);
nand I_32434 (I554276,I554259,I417029);
nor I_32435 (I554293,I554242,I554276);
DFFARX1 I_32436 (I554293,I2859,I554095,I554060,);
not I_32437 (I554324,I554276);
nand I_32438 (I554341,I554146,I554324);
nand I_32439 (I554072,I554208,I554324);
DFFARX1 I_32440 (I554242,I2859,I554095,I554087,);
not I_32441 (I554386,I417038);
nor I_32442 (I554403,I554386,I417023);
nor I_32443 (I554420,I554403,I554225);
DFFARX1 I_32444 (I554420,I2859,I554095,I554084,);
not I_32445 (I554451,I554403);
DFFARX1 I_32446 (I554451,I2859,I554095,I554477,);
not I_32447 (I554485,I554477);
nor I_32448 (I554081,I554485,I554403);
nor I_32449 (I554516,I554386,I417023);
and I_32450 (I554533,I554516,I417026);
or I_32451 (I554550,I554533,I417029);
DFFARX1 I_32452 (I554550,I2859,I554095,I554576,);
not I_32453 (I554584,I554576);
nand I_32454 (I554601,I554584,I554324);
not I_32455 (I554075,I554601);
nand I_32456 (I554069,I554601,I554341);
nand I_32457 (I554066,I554584,I554208);
not I_32458 (I554690,I2866);
DFFARX1 I_32459 (I176184,I2859,I554690,I554716,);
DFFARX1 I_32460 (I176190,I2859,I554690,I554733,);
not I_32461 (I554741,I554733);
nor I_32462 (I554658,I554716,I554741);
DFFARX1 I_32463 (I554741,I2859,I554690,I554673,);
nor I_32464 (I554786,I176199,I176184);
and I_32465 (I554803,I554786,I176211);
nor I_32466 (I554820,I554803,I176199);
not I_32467 (I554837,I176199);
and I_32468 (I554854,I554837,I176187);
nand I_32469 (I554871,I554854,I176208);
nor I_32470 (I554888,I554837,I554871);
DFFARX1 I_32471 (I554888,I2859,I554690,I554655,);
not I_32472 (I554919,I554871);
nand I_32473 (I554936,I554741,I554919);
nand I_32474 (I554667,I554803,I554919);
DFFARX1 I_32475 (I554837,I2859,I554690,I554682,);
not I_32476 (I554981,I176196);
nor I_32477 (I554998,I554981,I176187);
nor I_32478 (I555015,I554998,I554820);
DFFARX1 I_32479 (I555015,I2859,I554690,I554679,);
not I_32480 (I555046,I554998);
DFFARX1 I_32481 (I555046,I2859,I554690,I555072,);
not I_32482 (I555080,I555072);
nor I_32483 (I554676,I555080,I554998);
nor I_32484 (I555111,I554981,I176193);
and I_32485 (I555128,I555111,I176205);
or I_32486 (I555145,I555128,I176202);
DFFARX1 I_32487 (I555145,I2859,I554690,I555171,);
not I_32488 (I555179,I555171);
nand I_32489 (I555196,I555179,I554919);
not I_32490 (I554670,I555196);
nand I_32491 (I554664,I555196,I554936);
nand I_32492 (I554661,I555179,I554803);
not I_32493 (I555285,I2866);
DFFARX1 I_32494 (I385069,I2859,I555285,I555311,);
DFFARX1 I_32495 (I385087,I2859,I555285,I555328,);
not I_32496 (I555336,I555328);
nor I_32497 (I555253,I555311,I555336);
DFFARX1 I_32498 (I555336,I2859,I555285,I555268,);
nor I_32499 (I555381,I385066,I385078);
and I_32500 (I555398,I555381,I385063);
nor I_32501 (I555415,I555398,I385066);
not I_32502 (I555432,I385066);
and I_32503 (I555449,I555432,I385072);
nand I_32504 (I555466,I555449,I385084);
nor I_32505 (I555483,I555432,I555466);
DFFARX1 I_32506 (I555483,I2859,I555285,I555250,);
not I_32507 (I555514,I555466);
nand I_32508 (I555531,I555336,I555514);
nand I_32509 (I555262,I555398,I555514);
DFFARX1 I_32510 (I555432,I2859,I555285,I555277,);
not I_32511 (I555576,I385075);
nor I_32512 (I555593,I555576,I385072);
nor I_32513 (I555610,I555593,I555415);
DFFARX1 I_32514 (I555610,I2859,I555285,I555274,);
not I_32515 (I555641,I555593);
DFFARX1 I_32516 (I555641,I2859,I555285,I555667,);
not I_32517 (I555675,I555667);
nor I_32518 (I555271,I555675,I555593);
nor I_32519 (I555706,I555576,I385063);
and I_32520 (I555723,I555706,I385090);
or I_32521 (I555740,I555723,I385081);
DFFARX1 I_32522 (I555740,I2859,I555285,I555766,);
not I_32523 (I555774,I555766);
nand I_32524 (I555791,I555774,I555514);
not I_32525 (I555265,I555791);
nand I_32526 (I555259,I555791,I555531);
nand I_32527 (I555256,I555774,I555398);
not I_32528 (I555880,I2866);
DFFARX1 I_32529 (I197944,I2859,I555880,I555906,);
DFFARX1 I_32530 (I197950,I2859,I555880,I555923,);
not I_32531 (I555931,I555923);
nor I_32532 (I555848,I555906,I555931);
DFFARX1 I_32533 (I555931,I2859,I555880,I555863,);
nor I_32534 (I555976,I197959,I197944);
and I_32535 (I555993,I555976,I197971);
nor I_32536 (I556010,I555993,I197959);
not I_32537 (I556027,I197959);
and I_32538 (I556044,I556027,I197947);
nand I_32539 (I556061,I556044,I197968);
nor I_32540 (I556078,I556027,I556061);
DFFARX1 I_32541 (I556078,I2859,I555880,I555845,);
not I_32542 (I556109,I556061);
nand I_32543 (I556126,I555931,I556109);
nand I_32544 (I555857,I555993,I556109);
DFFARX1 I_32545 (I556027,I2859,I555880,I555872,);
not I_32546 (I556171,I197956);
nor I_32547 (I556188,I556171,I197947);
nor I_32548 (I556205,I556188,I556010);
DFFARX1 I_32549 (I556205,I2859,I555880,I555869,);
not I_32550 (I556236,I556188);
DFFARX1 I_32551 (I556236,I2859,I555880,I556262,);
not I_32552 (I556270,I556262);
nor I_32553 (I555866,I556270,I556188);
nor I_32554 (I556301,I556171,I197953);
and I_32555 (I556318,I556301,I197965);
or I_32556 (I556335,I556318,I197962);
DFFARX1 I_32557 (I556335,I2859,I555880,I556361,);
not I_32558 (I556369,I556361);
nand I_32559 (I556386,I556369,I556109);
not I_32560 (I555860,I556386);
nand I_32561 (I555854,I556386,I556126);
nand I_32562 (I555851,I556369,I555993);
not I_32563 (I556475,I2866);
DFFARX1 I_32564 (I223295,I2859,I556475,I556501,);
DFFARX1 I_32565 (I223289,I2859,I556475,I556518,);
not I_32566 (I556526,I556518);
nor I_32567 (I556443,I556501,I556526);
DFFARX1 I_32568 (I556526,I2859,I556475,I556458,);
nor I_32569 (I556571,I223286,I223277);
and I_32570 (I556588,I556571,I223274);
nor I_32571 (I556605,I556588,I223286);
not I_32572 (I556622,I223286);
and I_32573 (I556639,I556622,I223280);
nand I_32574 (I556656,I556639,I223292);
nor I_32575 (I556673,I556622,I556656);
DFFARX1 I_32576 (I556673,I2859,I556475,I556440,);
not I_32577 (I556704,I556656);
nand I_32578 (I556721,I556526,I556704);
nand I_32579 (I556452,I556588,I556704);
DFFARX1 I_32580 (I556622,I2859,I556475,I556467,);
not I_32581 (I556766,I223298);
nor I_32582 (I556783,I556766,I223280);
nor I_32583 (I556800,I556783,I556605);
DFFARX1 I_32584 (I556800,I2859,I556475,I556464,);
not I_32585 (I556831,I556783);
DFFARX1 I_32586 (I556831,I2859,I556475,I556857,);
not I_32587 (I556865,I556857);
nor I_32588 (I556461,I556865,I556783);
nor I_32589 (I556896,I556766,I223277);
and I_32590 (I556913,I556896,I223283);
or I_32591 (I556930,I556913,I223274);
DFFARX1 I_32592 (I556930,I2859,I556475,I556956,);
not I_32593 (I556964,I556956);
nand I_32594 (I556981,I556964,I556704);
not I_32595 (I556455,I556981);
nand I_32596 (I556449,I556981,I556721);
nand I_32597 (I556446,I556964,I556588);
not I_32598 (I557070,I2866);
DFFARX1 I_32599 (I194136,I2859,I557070,I557096,);
DFFARX1 I_32600 (I194142,I2859,I557070,I557113,);
not I_32601 (I557121,I557113);
nor I_32602 (I557038,I557096,I557121);
DFFARX1 I_32603 (I557121,I2859,I557070,I557053,);
nor I_32604 (I557166,I194151,I194136);
and I_32605 (I557183,I557166,I194163);
nor I_32606 (I557200,I557183,I194151);
not I_32607 (I557217,I194151);
and I_32608 (I557234,I557217,I194139);
nand I_32609 (I557251,I557234,I194160);
nor I_32610 (I557268,I557217,I557251);
DFFARX1 I_32611 (I557268,I2859,I557070,I557035,);
not I_32612 (I557299,I557251);
nand I_32613 (I557316,I557121,I557299);
nand I_32614 (I557047,I557183,I557299);
DFFARX1 I_32615 (I557217,I2859,I557070,I557062,);
not I_32616 (I557361,I194148);
nor I_32617 (I557378,I557361,I194139);
nor I_32618 (I557395,I557378,I557200);
DFFARX1 I_32619 (I557395,I2859,I557070,I557059,);
not I_32620 (I557426,I557378);
DFFARX1 I_32621 (I557426,I2859,I557070,I557452,);
not I_32622 (I557460,I557452);
nor I_32623 (I557056,I557460,I557378);
nor I_32624 (I557491,I557361,I194145);
and I_32625 (I557508,I557491,I194157);
or I_32626 (I557525,I557508,I194154);
DFFARX1 I_32627 (I557525,I2859,I557070,I557551,);
not I_32628 (I557559,I557551);
nand I_32629 (I557576,I557559,I557299);
not I_32630 (I557050,I557576);
nand I_32631 (I557044,I557576,I557316);
nand I_32632 (I557041,I557559,I557183);
not I_32633 (I557665,I2866);
DFFARX1 I_32634 (I523546,I2859,I557665,I557691,);
DFFARX1 I_32635 (I523537,I2859,I557665,I557708,);
not I_32636 (I557716,I557708);
nor I_32637 (I557633,I557691,I557716);
DFFARX1 I_32638 (I557716,I2859,I557665,I557648,);
nor I_32639 (I557761,I523528,I523543);
and I_32640 (I557778,I557761,I523531);
nor I_32641 (I557795,I557778,I523528);
not I_32642 (I557812,I523528);
and I_32643 (I557829,I557812,I523534);
nand I_32644 (I557846,I557829,I523552);
nor I_32645 (I557863,I557812,I557846);
DFFARX1 I_32646 (I557863,I2859,I557665,I557630,);
not I_32647 (I557894,I557846);
nand I_32648 (I557911,I557716,I557894);
nand I_32649 (I557642,I557778,I557894);
DFFARX1 I_32650 (I557812,I2859,I557665,I557657,);
not I_32651 (I557956,I523528);
nor I_32652 (I557973,I557956,I523534);
nor I_32653 (I557990,I557973,I557795);
DFFARX1 I_32654 (I557990,I2859,I557665,I557654,);
not I_32655 (I558021,I557973);
DFFARX1 I_32656 (I558021,I2859,I557665,I558047,);
not I_32657 (I558055,I558047);
nor I_32658 (I557651,I558055,I557973);
nor I_32659 (I558086,I557956,I523531);
and I_32660 (I558103,I558086,I523540);
or I_32661 (I558120,I558103,I523549);
DFFARX1 I_32662 (I558120,I2859,I557665,I558146,);
not I_32663 (I558154,I558146);
nand I_32664 (I558171,I558154,I557894);
not I_32665 (I557645,I558171);
nand I_32666 (I557639,I558171,I557911);
nand I_32667 (I557636,I558154,I557778);
not I_32668 (I558260,I2866);
DFFARX1 I_32669 (I361289,I2859,I558260,I558286,);
DFFARX1 I_32670 (I361286,I2859,I558260,I558303,);
not I_32671 (I558311,I558303);
nor I_32672 (I558228,I558286,I558311);
DFFARX1 I_32673 (I558311,I2859,I558260,I558243,);
nor I_32674 (I558356,I361301,I361283);
and I_32675 (I558373,I558356,I361280);
nor I_32676 (I558390,I558373,I361301);
not I_32677 (I558407,I361301);
and I_32678 (I558424,I558407,I361286);
nand I_32679 (I558441,I558424,I361298);
nor I_32680 (I558458,I558407,I558441);
DFFARX1 I_32681 (I558458,I2859,I558260,I558225,);
not I_32682 (I558489,I558441);
nand I_32683 (I558506,I558311,I558489);
nand I_32684 (I558237,I558373,I558489);
DFFARX1 I_32685 (I558407,I2859,I558260,I558252,);
not I_32686 (I558551,I361292);
nor I_32687 (I558568,I558551,I361286);
nor I_32688 (I558585,I558568,I558390);
DFFARX1 I_32689 (I558585,I2859,I558260,I558249,);
not I_32690 (I558616,I558568);
DFFARX1 I_32691 (I558616,I2859,I558260,I558642,);
not I_32692 (I558650,I558642);
nor I_32693 (I558246,I558650,I558568);
nor I_32694 (I558681,I558551,I361280);
and I_32695 (I558698,I558681,I361295);
or I_32696 (I558715,I558698,I361283);
DFFARX1 I_32697 (I558715,I2859,I558260,I558741,);
not I_32698 (I558749,I558741);
nand I_32699 (I558766,I558749,I558489);
not I_32700 (I558240,I558766);
nand I_32701 (I558234,I558766,I558506);
nand I_32702 (I558231,I558749,I558373);
not I_32703 (I558855,I2866);
DFFARX1 I_32704 (I191416,I2859,I558855,I558881,);
DFFARX1 I_32705 (I191422,I2859,I558855,I558898,);
not I_32706 (I558906,I558898);
nor I_32707 (I558823,I558881,I558906);
DFFARX1 I_32708 (I558906,I2859,I558855,I558838,);
nor I_32709 (I558951,I191431,I191416);
and I_32710 (I558968,I558951,I191443);
nor I_32711 (I558985,I558968,I191431);
not I_32712 (I559002,I191431);
and I_32713 (I559019,I559002,I191419);
nand I_32714 (I559036,I559019,I191440);
nor I_32715 (I559053,I559002,I559036);
DFFARX1 I_32716 (I559053,I2859,I558855,I558820,);
not I_32717 (I559084,I559036);
nand I_32718 (I559101,I558906,I559084);
nand I_32719 (I558832,I558968,I559084);
DFFARX1 I_32720 (I559002,I2859,I558855,I558847,);
not I_32721 (I559146,I191428);
nor I_32722 (I559163,I559146,I191419);
nor I_32723 (I559180,I559163,I558985);
DFFARX1 I_32724 (I559180,I2859,I558855,I558844,);
not I_32725 (I559211,I559163);
DFFARX1 I_32726 (I559211,I2859,I558855,I559237,);
not I_32727 (I559245,I559237);
nor I_32728 (I558841,I559245,I559163);
nor I_32729 (I559276,I559146,I191425);
and I_32730 (I559293,I559276,I191437);
or I_32731 (I559310,I559293,I191434);
DFFARX1 I_32732 (I559310,I2859,I558855,I559336,);
not I_32733 (I559344,I559336);
nand I_32734 (I559361,I559344,I559084);
not I_32735 (I558835,I559361);
nand I_32736 (I558829,I559361,I559101);
nand I_32737 (I558826,I559344,I558968);
not I_32738 (I559450,I2866);
DFFARX1 I_32739 (I123539,I2859,I559450,I559476,);
DFFARX1 I_32740 (I123533,I2859,I559450,I559493,);
not I_32741 (I559501,I559493);
nor I_32742 (I559418,I559476,I559501);
DFFARX1 I_32743 (I559501,I2859,I559450,I559433,);
nor I_32744 (I559546,I123521,I123542);
and I_32745 (I559563,I559546,I123536);
nor I_32746 (I559580,I559563,I123521);
not I_32747 (I559597,I123521);
and I_32748 (I559614,I559597,I123518);
nand I_32749 (I559631,I559614,I123530);
nor I_32750 (I559648,I559597,I559631);
DFFARX1 I_32751 (I559648,I2859,I559450,I559415,);
not I_32752 (I559679,I559631);
nand I_32753 (I559696,I559501,I559679);
nand I_32754 (I559427,I559563,I559679);
DFFARX1 I_32755 (I559597,I2859,I559450,I559442,);
not I_32756 (I559741,I123545);
nor I_32757 (I559758,I559741,I123518);
nor I_32758 (I559775,I559758,I559580);
DFFARX1 I_32759 (I559775,I2859,I559450,I559439,);
not I_32760 (I559806,I559758);
DFFARX1 I_32761 (I559806,I2859,I559450,I559832,);
not I_32762 (I559840,I559832);
nor I_32763 (I559436,I559840,I559758);
nor I_32764 (I559871,I559741,I123527);
and I_32765 (I559888,I559871,I123524);
or I_32766 (I559905,I559888,I123518);
DFFARX1 I_32767 (I559905,I2859,I559450,I559931,);
not I_32768 (I559939,I559931);
nand I_32769 (I559956,I559939,I559679);
not I_32770 (I559430,I559956);
nand I_32771 (I559424,I559956,I559696);
nand I_32772 (I559421,I559939,I559563);
not I_32773 (I560045,I2866);
DFFARX1 I_32774 (I126701,I2859,I560045,I560071,);
DFFARX1 I_32775 (I126695,I2859,I560045,I560088,);
not I_32776 (I560096,I560088);
nor I_32777 (I560013,I560071,I560096);
DFFARX1 I_32778 (I560096,I2859,I560045,I560028,);
nor I_32779 (I560141,I126683,I126704);
and I_32780 (I560158,I560141,I126698);
nor I_32781 (I560175,I560158,I126683);
not I_32782 (I560192,I126683);
and I_32783 (I560209,I560192,I126680);
nand I_32784 (I560226,I560209,I126692);
nor I_32785 (I560243,I560192,I560226);
DFFARX1 I_32786 (I560243,I2859,I560045,I560010,);
not I_32787 (I560274,I560226);
nand I_32788 (I560291,I560096,I560274);
nand I_32789 (I560022,I560158,I560274);
DFFARX1 I_32790 (I560192,I2859,I560045,I560037,);
not I_32791 (I560336,I126707);
nor I_32792 (I560353,I560336,I126680);
nor I_32793 (I560370,I560353,I560175);
DFFARX1 I_32794 (I560370,I2859,I560045,I560034,);
not I_32795 (I560401,I560353);
DFFARX1 I_32796 (I560401,I2859,I560045,I560427,);
not I_32797 (I560435,I560427);
nor I_32798 (I560031,I560435,I560353);
nor I_32799 (I560466,I560336,I126689);
and I_32800 (I560483,I560466,I126686);
or I_32801 (I560500,I560483,I126680);
DFFARX1 I_32802 (I560500,I2859,I560045,I560526,);
not I_32803 (I560534,I560526);
nand I_32804 (I560551,I560534,I560274);
not I_32805 (I560025,I560551);
nand I_32806 (I560019,I560551,I560291);
nand I_32807 (I560016,I560534,I560158);
not I_32808 (I560640,I2866);
DFFARX1 I_32809 (I371503,I2859,I560640,I560666,);
DFFARX1 I_32810 (I371521,I2859,I560640,I560683,);
not I_32811 (I560691,I560683);
nor I_32812 (I560608,I560666,I560691);
DFFARX1 I_32813 (I560691,I2859,I560640,I560623,);
nor I_32814 (I560736,I371500,I371512);
and I_32815 (I560753,I560736,I371497);
nor I_32816 (I560770,I560753,I371500);
not I_32817 (I560787,I371500);
and I_32818 (I560804,I560787,I371506);
nand I_32819 (I560821,I560804,I371518);
nor I_32820 (I560838,I560787,I560821);
DFFARX1 I_32821 (I560838,I2859,I560640,I560605,);
not I_32822 (I560869,I560821);
nand I_32823 (I560886,I560691,I560869);
nand I_32824 (I560617,I560753,I560869);
DFFARX1 I_32825 (I560787,I2859,I560640,I560632,);
not I_32826 (I560931,I371509);
nor I_32827 (I560948,I560931,I371506);
nor I_32828 (I560965,I560948,I560770);
DFFARX1 I_32829 (I560965,I2859,I560640,I560629,);
not I_32830 (I560996,I560948);
DFFARX1 I_32831 (I560996,I2859,I560640,I561022,);
not I_32832 (I561030,I561022);
nor I_32833 (I560626,I561030,I560948);
nor I_32834 (I561061,I560931,I371497);
and I_32835 (I561078,I561061,I371524);
or I_32836 (I561095,I561078,I371515);
DFFARX1 I_32837 (I561095,I2859,I560640,I561121,);
not I_32838 (I561129,I561121);
nand I_32839 (I561146,I561129,I560869);
not I_32840 (I560620,I561146);
nand I_32841 (I560614,I561146,I560886);
nand I_32842 (I560611,I561129,I560753);
not I_32843 (I561235,I2866);
DFFARX1 I_32844 (I103067,I2859,I561235,I561261,);
DFFARX1 I_32845 (I103070,I2859,I561235,I561278,);
not I_32846 (I561286,I561278);
nor I_32847 (I561203,I561261,I561286);
DFFARX1 I_32848 (I561286,I2859,I561235,I561218,);
nor I_32849 (I561331,I103076,I103070);
and I_32850 (I561348,I561331,I103073);
nor I_32851 (I561365,I561348,I103076);
not I_32852 (I561382,I103076);
and I_32853 (I561399,I561382,I103067);
nand I_32854 (I561416,I561399,I103085);
nor I_32855 (I561433,I561382,I561416);
DFFARX1 I_32856 (I561433,I2859,I561235,I561200,);
not I_32857 (I561464,I561416);
nand I_32858 (I561481,I561286,I561464);
nand I_32859 (I561212,I561348,I561464);
DFFARX1 I_32860 (I561382,I2859,I561235,I561227,);
not I_32861 (I561526,I103079);
nor I_32862 (I561543,I561526,I103067);
nor I_32863 (I561560,I561543,I561365);
DFFARX1 I_32864 (I561560,I2859,I561235,I561224,);
not I_32865 (I561591,I561543);
DFFARX1 I_32866 (I561591,I2859,I561235,I561617,);
not I_32867 (I561625,I561617);
nor I_32868 (I561221,I561625,I561543);
nor I_32869 (I561656,I561526,I103082);
and I_32870 (I561673,I561656,I103088);
or I_32871 (I561690,I561673,I103091);
DFFARX1 I_32872 (I561690,I2859,I561235,I561716,);
not I_32873 (I561724,I561716);
nand I_32874 (I561741,I561724,I561464);
not I_32875 (I561215,I561741);
nand I_32876 (I561209,I561741,I561481);
nand I_32877 (I561206,I561724,I561348);
not I_32878 (I561830,I2866);
DFFARX1 I_32879 (I134606,I2859,I561830,I561856,);
DFFARX1 I_32880 (I134600,I2859,I561830,I561873,);
not I_32881 (I561881,I561873);
nor I_32882 (I561798,I561856,I561881);
DFFARX1 I_32883 (I561881,I2859,I561830,I561813,);
nor I_32884 (I561926,I134588,I134609);
and I_32885 (I561943,I561926,I134603);
nor I_32886 (I561960,I561943,I134588);
not I_32887 (I561977,I134588);
and I_32888 (I561994,I561977,I134585);
nand I_32889 (I562011,I561994,I134597);
nor I_32890 (I562028,I561977,I562011);
DFFARX1 I_32891 (I562028,I2859,I561830,I561795,);
not I_32892 (I562059,I562011);
nand I_32893 (I562076,I561881,I562059);
nand I_32894 (I561807,I561943,I562059);
DFFARX1 I_32895 (I561977,I2859,I561830,I561822,);
not I_32896 (I562121,I134612);
nor I_32897 (I562138,I562121,I134585);
nor I_32898 (I562155,I562138,I561960);
DFFARX1 I_32899 (I562155,I2859,I561830,I561819,);
not I_32900 (I562186,I562138);
DFFARX1 I_32901 (I562186,I2859,I561830,I562212,);
not I_32902 (I562220,I562212);
nor I_32903 (I561816,I562220,I562138);
nor I_32904 (I562251,I562121,I134594);
and I_32905 (I562268,I562251,I134591);
or I_32906 (I562285,I562268,I134585);
DFFARX1 I_32907 (I562285,I2859,I561830,I562311,);
not I_32908 (I562319,I562311);
nand I_32909 (I562336,I562319,I562059);
not I_32910 (I561810,I562336);
nand I_32911 (I561804,I562336,I562076);
nand I_32912 (I561801,I562319,I561943);
not I_32913 (I562425,I2866);
DFFARX1 I_32914 (I237745,I2859,I562425,I562451,);
DFFARX1 I_32915 (I237739,I2859,I562425,I562468,);
not I_32916 (I562476,I562468);
nor I_32917 (I562393,I562451,I562476);
DFFARX1 I_32918 (I562476,I2859,I562425,I562408,);
nor I_32919 (I562521,I237736,I237727);
and I_32920 (I562538,I562521,I237724);
nor I_32921 (I562555,I562538,I237736);
not I_32922 (I562572,I237736);
and I_32923 (I562589,I562572,I237730);
nand I_32924 (I562606,I562589,I237742);
nor I_32925 (I562623,I562572,I562606);
DFFARX1 I_32926 (I562623,I2859,I562425,I562390,);
not I_32927 (I562654,I562606);
nand I_32928 (I562671,I562476,I562654);
nand I_32929 (I562402,I562538,I562654);
DFFARX1 I_32930 (I562572,I2859,I562425,I562417,);
not I_32931 (I562716,I237748);
nor I_32932 (I562733,I562716,I237730);
nor I_32933 (I562750,I562733,I562555);
DFFARX1 I_32934 (I562750,I2859,I562425,I562414,);
not I_32935 (I562781,I562733);
DFFARX1 I_32936 (I562781,I2859,I562425,I562807,);
not I_32937 (I562815,I562807);
nor I_32938 (I562411,I562815,I562733);
nor I_32939 (I562846,I562716,I237727);
and I_32940 (I562863,I562846,I237733);
or I_32941 (I562880,I562863,I237724);
DFFARX1 I_32942 (I562880,I2859,I562425,I562906,);
not I_32943 (I562914,I562906);
nand I_32944 (I562931,I562914,I562654);
not I_32945 (I562405,I562931);
nand I_32946 (I562399,I562931,I562671);
nand I_32947 (I562396,I562914,I562538);
not I_32948 (I563020,I2866);
DFFARX1 I_32949 (I6389,I2859,I563020,I563046,);
DFFARX1 I_32950 (I6371,I2859,I563020,I563063,);
not I_32951 (I563071,I563063);
nor I_32952 (I562988,I563046,I563071);
DFFARX1 I_32953 (I563071,I2859,I563020,I563003,);
nor I_32954 (I563116,I6371,I6386);
and I_32955 (I563133,I563116,I6380);
nor I_32956 (I563150,I563133,I6371);
not I_32957 (I563167,I6371);
and I_32958 (I563184,I563167,I6374);
nand I_32959 (I563201,I563184,I6377);
nor I_32960 (I563218,I563167,I563201);
DFFARX1 I_32961 (I563218,I2859,I563020,I562985,);
not I_32962 (I563249,I563201);
nand I_32963 (I563266,I563071,I563249);
nand I_32964 (I562997,I563133,I563249);
DFFARX1 I_32965 (I563167,I2859,I563020,I563012,);
not I_32966 (I563311,I6383);
nor I_32967 (I563328,I563311,I6374);
nor I_32968 (I563345,I563328,I563150);
DFFARX1 I_32969 (I563345,I2859,I563020,I563009,);
not I_32970 (I563376,I563328);
DFFARX1 I_32971 (I563376,I2859,I563020,I563402,);
not I_32972 (I563410,I563402);
nor I_32973 (I563006,I563410,I563328);
nor I_32974 (I563441,I563311,I6395);
and I_32975 (I563458,I563441,I6392);
or I_32976 (I563475,I563458,I6374);
DFFARX1 I_32977 (I563475,I2859,I563020,I563501,);
not I_32978 (I563509,I563501);
nand I_32979 (I563526,I563509,I563249);
not I_32980 (I563000,I563526);
nand I_32981 (I562994,I563526,I563266);
nand I_32982 (I562991,I563509,I563133);
not I_32983 (I563615,I2866);
DFFARX1 I_32984 (I437792,I2859,I563615,I563641,);
DFFARX1 I_32985 (I437783,I2859,I563615,I563658,);
not I_32986 (I563666,I563658);
nor I_32987 (I563583,I563641,I563666);
DFFARX1 I_32988 (I563666,I2859,I563615,I563598,);
nor I_32989 (I563711,I437789,I437798);
and I_32990 (I563728,I563711,I437801);
nor I_32991 (I563745,I563728,I437789);
not I_32992 (I563762,I437789);
and I_32993 (I563779,I563762,I437780);
nand I_32994 (I563796,I563779,I437786);
nor I_32995 (I563813,I563762,I563796);
DFFARX1 I_32996 (I563813,I2859,I563615,I563580,);
not I_32997 (I563844,I563796);
nand I_32998 (I563861,I563666,I563844);
nand I_32999 (I563592,I563728,I563844);
DFFARX1 I_33000 (I563762,I2859,I563615,I563607,);
not I_33001 (I563906,I437795);
nor I_33002 (I563923,I563906,I437780);
nor I_33003 (I563940,I563923,I563745);
DFFARX1 I_33004 (I563940,I2859,I563615,I563604,);
not I_33005 (I563971,I563923);
DFFARX1 I_33006 (I563971,I2859,I563615,I563997,);
not I_33007 (I564005,I563997);
nor I_33008 (I563601,I564005,I563923);
nor I_33009 (I564036,I563906,I437780);
and I_33010 (I564053,I564036,I437783);
or I_33011 (I564070,I564053,I437786);
DFFARX1 I_33012 (I564070,I2859,I563615,I564096,);
not I_33013 (I564104,I564096);
nand I_33014 (I564121,I564104,I563844);
not I_33015 (I563595,I564121);
nand I_33016 (I563589,I564121,I563861);
nand I_33017 (I563586,I564104,I563728);
not I_33018 (I564210,I2866);
DFFARX1 I_33019 (I73317,I2859,I564210,I564236,);
DFFARX1 I_33020 (I73320,I2859,I564210,I564253,);
not I_33021 (I564261,I564253);
nor I_33022 (I564178,I564236,I564261);
DFFARX1 I_33023 (I564261,I2859,I564210,I564193,);
nor I_33024 (I564306,I73326,I73320);
and I_33025 (I564323,I564306,I73323);
nor I_33026 (I564340,I564323,I73326);
not I_33027 (I564357,I73326);
and I_33028 (I564374,I564357,I73317);
nand I_33029 (I564391,I564374,I73335);
nor I_33030 (I564408,I564357,I564391);
DFFARX1 I_33031 (I564408,I2859,I564210,I564175,);
not I_33032 (I564439,I564391);
nand I_33033 (I564456,I564261,I564439);
nand I_33034 (I564187,I564323,I564439);
DFFARX1 I_33035 (I564357,I2859,I564210,I564202,);
not I_33036 (I564501,I73329);
nor I_33037 (I564518,I564501,I73317);
nor I_33038 (I564535,I564518,I564340);
DFFARX1 I_33039 (I564535,I2859,I564210,I564199,);
not I_33040 (I564566,I564518);
DFFARX1 I_33041 (I564566,I2859,I564210,I564592,);
not I_33042 (I564600,I564592);
nor I_33043 (I564196,I564600,I564518);
nor I_33044 (I564631,I564501,I73332);
and I_33045 (I564648,I564631,I73338);
or I_33046 (I564665,I564648,I73341);
DFFARX1 I_33047 (I564665,I2859,I564210,I564691,);
not I_33048 (I564699,I564691);
nand I_33049 (I564716,I564699,I564439);
not I_33050 (I564190,I564716);
nand I_33051 (I564184,I564716,I564456);
nand I_33052 (I564181,I564699,I564323);
not I_33053 (I564805,I2866);
DFFARX1 I_33054 (I59037,I2859,I564805,I564831,);
DFFARX1 I_33055 (I59040,I2859,I564805,I564848,);
not I_33056 (I564856,I564848);
nor I_33057 (I564773,I564831,I564856);
DFFARX1 I_33058 (I564856,I2859,I564805,I564788,);
nor I_33059 (I564901,I59046,I59040);
and I_33060 (I564918,I564901,I59043);
nor I_33061 (I564935,I564918,I59046);
not I_33062 (I564952,I59046);
and I_33063 (I564969,I564952,I59037);
nand I_33064 (I564986,I564969,I59055);
nor I_33065 (I565003,I564952,I564986);
DFFARX1 I_33066 (I565003,I2859,I564805,I564770,);
not I_33067 (I565034,I564986);
nand I_33068 (I565051,I564856,I565034);
nand I_33069 (I564782,I564918,I565034);
DFFARX1 I_33070 (I564952,I2859,I564805,I564797,);
not I_33071 (I565096,I59049);
nor I_33072 (I565113,I565096,I59037);
nor I_33073 (I565130,I565113,I564935);
DFFARX1 I_33074 (I565130,I2859,I564805,I564794,);
not I_33075 (I565161,I565113);
DFFARX1 I_33076 (I565161,I2859,I564805,I565187,);
not I_33077 (I565195,I565187);
nor I_33078 (I564791,I565195,I565113);
nor I_33079 (I565226,I565096,I59052);
and I_33080 (I565243,I565226,I59058);
or I_33081 (I565260,I565243,I59061);
DFFARX1 I_33082 (I565260,I2859,I564805,I565286,);
not I_33083 (I565294,I565286);
nand I_33084 (I565311,I565294,I565034);
not I_33085 (I564785,I565311);
nand I_33086 (I564779,I565311,I565051);
nand I_33087 (I564776,I565294,I564918);
not I_33088 (I565400,I2866);
DFFARX1 I_33089 (I56062,I2859,I565400,I565426,);
DFFARX1 I_33090 (I56065,I2859,I565400,I565443,);
not I_33091 (I565451,I565443);
nor I_33092 (I565368,I565426,I565451);
DFFARX1 I_33093 (I565451,I2859,I565400,I565383,);
nor I_33094 (I565496,I56071,I56065);
and I_33095 (I565513,I565496,I56068);
nor I_33096 (I565530,I565513,I56071);
not I_33097 (I565547,I56071);
and I_33098 (I565564,I565547,I56062);
nand I_33099 (I565581,I565564,I56080);
nor I_33100 (I565598,I565547,I565581);
DFFARX1 I_33101 (I565598,I2859,I565400,I565365,);
not I_33102 (I565629,I565581);
nand I_33103 (I565646,I565451,I565629);
nand I_33104 (I565377,I565513,I565629);
DFFARX1 I_33105 (I565547,I2859,I565400,I565392,);
not I_33106 (I565691,I56074);
nor I_33107 (I565708,I565691,I56062);
nor I_33108 (I565725,I565708,I565530);
DFFARX1 I_33109 (I565725,I2859,I565400,I565389,);
not I_33110 (I565756,I565708);
DFFARX1 I_33111 (I565756,I2859,I565400,I565782,);
not I_33112 (I565790,I565782);
nor I_33113 (I565386,I565790,I565708);
nor I_33114 (I565821,I565691,I56077);
and I_33115 (I565838,I565821,I56083);
or I_33116 (I565855,I565838,I56086);
DFFARX1 I_33117 (I565855,I2859,I565400,I565881,);
not I_33118 (I565889,I565881);
nand I_33119 (I565906,I565889,I565629);
not I_33120 (I565380,I565906);
nand I_33121 (I565374,I565906,I565646);
nand I_33122 (I565371,I565889,I565513);
not I_33123 (I565995,I2866);
DFFARX1 I_33124 (I107232,I2859,I565995,I566021,);
DFFARX1 I_33125 (I107235,I2859,I565995,I566038,);
not I_33126 (I566046,I566038);
nor I_33127 (I565963,I566021,I566046);
DFFARX1 I_33128 (I566046,I2859,I565995,I565978,);
nor I_33129 (I566091,I107241,I107235);
and I_33130 (I566108,I566091,I107238);
nor I_33131 (I566125,I566108,I107241);
not I_33132 (I566142,I107241);
and I_33133 (I566159,I566142,I107232);
nand I_33134 (I566176,I566159,I107250);
nor I_33135 (I566193,I566142,I566176);
DFFARX1 I_33136 (I566193,I2859,I565995,I565960,);
not I_33137 (I566224,I566176);
nand I_33138 (I566241,I566046,I566224);
nand I_33139 (I565972,I566108,I566224);
DFFARX1 I_33140 (I566142,I2859,I565995,I565987,);
not I_33141 (I566286,I107244);
nor I_33142 (I566303,I566286,I107232);
nor I_33143 (I566320,I566303,I566125);
DFFARX1 I_33144 (I566320,I2859,I565995,I565984,);
not I_33145 (I566351,I566303);
DFFARX1 I_33146 (I566351,I2859,I565995,I566377,);
not I_33147 (I566385,I566377);
nor I_33148 (I565981,I566385,I566303);
nor I_33149 (I566416,I566286,I107247);
and I_33150 (I566433,I566416,I107253);
or I_33151 (I566450,I566433,I107256);
DFFARX1 I_33152 (I566450,I2859,I565995,I566476,);
not I_33153 (I566484,I566476);
nand I_33154 (I566501,I566484,I566224);
not I_33155 (I565975,I566501);
nand I_33156 (I565969,I566501,I566241);
nand I_33157 (I565966,I566484,I566108);
not I_33158 (I566590,I2866);
DFFARX1 I_33159 (I421523,I2859,I566590,I566616,);
DFFARX1 I_33160 (I421514,I2859,I566590,I566633,);
not I_33161 (I566641,I566633);
nor I_33162 (I566558,I566616,I566641);
DFFARX1 I_33163 (I566641,I2859,I566590,I566573,);
nor I_33164 (I566686,I421520,I421529);
and I_33165 (I566703,I566686,I421532);
nor I_33166 (I566720,I566703,I421520);
not I_33167 (I566737,I421520);
and I_33168 (I566754,I566737,I421511);
nand I_33169 (I566771,I566754,I421517);
nor I_33170 (I566788,I566737,I566771);
DFFARX1 I_33171 (I566788,I2859,I566590,I566555,);
not I_33172 (I566819,I566771);
nand I_33173 (I566836,I566641,I566819);
nand I_33174 (I566567,I566703,I566819);
DFFARX1 I_33175 (I566737,I2859,I566590,I566582,);
not I_33176 (I566881,I421526);
nor I_33177 (I566898,I566881,I421511);
nor I_33178 (I566915,I566898,I566720);
DFFARX1 I_33179 (I566915,I2859,I566590,I566579,);
not I_33180 (I566946,I566898);
DFFARX1 I_33181 (I566946,I2859,I566590,I566972,);
not I_33182 (I566980,I566972);
nor I_33183 (I566576,I566980,I566898);
nor I_33184 (I567011,I566881,I421511);
and I_33185 (I567028,I567011,I421514);
or I_33186 (I567045,I567028,I421517);
DFFARX1 I_33187 (I567045,I2859,I566590,I567071,);
not I_33188 (I567079,I567071);
nand I_33189 (I567096,I567079,I566819);
not I_33190 (I566570,I567096);
nand I_33191 (I566564,I567096,I566836);
nand I_33192 (I566561,I567079,I566703);
not I_33193 (I567185,I2866);
DFFARX1 I_33194 (I137241,I2859,I567185,I567211,);
DFFARX1 I_33195 (I137235,I2859,I567185,I567228,);
not I_33196 (I567236,I567228);
nor I_33197 (I567153,I567211,I567236);
DFFARX1 I_33198 (I567236,I2859,I567185,I567168,);
nor I_33199 (I567281,I137223,I137244);
and I_33200 (I567298,I567281,I137238);
nor I_33201 (I567315,I567298,I137223);
not I_33202 (I567332,I137223);
and I_33203 (I567349,I567332,I137220);
nand I_33204 (I567366,I567349,I137232);
nor I_33205 (I567383,I567332,I567366);
DFFARX1 I_33206 (I567383,I2859,I567185,I567150,);
not I_33207 (I567414,I567366);
nand I_33208 (I567431,I567236,I567414);
nand I_33209 (I567162,I567298,I567414);
DFFARX1 I_33210 (I567332,I2859,I567185,I567177,);
not I_33211 (I567476,I137247);
nor I_33212 (I567493,I567476,I137220);
nor I_33213 (I567510,I567493,I567315);
DFFARX1 I_33214 (I567510,I2859,I567185,I567174,);
not I_33215 (I567541,I567493);
DFFARX1 I_33216 (I567541,I2859,I567185,I567567,);
not I_33217 (I567575,I567567);
nor I_33218 (I567171,I567575,I567493);
nor I_33219 (I567606,I567476,I137229);
and I_33220 (I567623,I567606,I137226);
or I_33221 (I567640,I567623,I137220);
DFFARX1 I_33222 (I567640,I2859,I567185,I567666,);
not I_33223 (I567674,I567666);
nand I_33224 (I567691,I567674,I567414);
not I_33225 (I567165,I567691);
nand I_33226 (I567159,I567691,I567431);
nand I_33227 (I567156,I567674,I567298);
not I_33228 (I567780,I2866);
DFFARX1 I_33229 (I1500,I2859,I567780,I567806,);
DFFARX1 I_33230 (I2412,I2859,I567780,I567823,);
not I_33231 (I567831,I567823);
nor I_33232 (I567748,I567806,I567831);
DFFARX1 I_33233 (I567831,I2859,I567780,I567763,);
nor I_33234 (I567876,I1916,I1852);
and I_33235 (I567893,I567876,I2196);
nor I_33236 (I567910,I567893,I1916);
not I_33237 (I567927,I1916);
and I_33238 (I567944,I567927,I2628);
nand I_33239 (I567961,I567944,I2164);
nor I_33240 (I567978,I567927,I567961);
DFFARX1 I_33241 (I567978,I2859,I567780,I567745,);
not I_33242 (I568009,I567961);
nand I_33243 (I568026,I567831,I568009);
nand I_33244 (I567757,I567893,I568009);
DFFARX1 I_33245 (I567927,I2859,I567780,I567772,);
not I_33246 (I568071,I2380);
nor I_33247 (I568088,I568071,I2628);
nor I_33248 (I568105,I568088,I567910);
DFFARX1 I_33249 (I568105,I2859,I567780,I567769,);
not I_33250 (I568136,I568088);
DFFARX1 I_33251 (I568136,I2859,I567780,I568162,);
not I_33252 (I568170,I568162);
nor I_33253 (I567766,I568170,I568088);
nor I_33254 (I568201,I568071,I1380);
and I_33255 (I568218,I568201,I1844);
or I_33256 (I568235,I568218,I1980);
DFFARX1 I_33257 (I568235,I2859,I567780,I568261,);
not I_33258 (I568269,I568261);
nand I_33259 (I568286,I568269,I568009);
not I_33260 (I567760,I568286);
nand I_33261 (I567754,I568286,I568026);
nand I_33262 (I567751,I568269,I567893);
not I_33263 (I568375,I2866);
DFFARX1 I_33264 (I520656,I2859,I568375,I568401,);
DFFARX1 I_33265 (I520647,I2859,I568375,I568418,);
not I_33266 (I568426,I568418);
nor I_33267 (I568343,I568401,I568426);
DFFARX1 I_33268 (I568426,I2859,I568375,I568358,);
nor I_33269 (I568471,I520638,I520653);
and I_33270 (I568488,I568471,I520641);
nor I_33271 (I568505,I568488,I520638);
not I_33272 (I568522,I520638);
and I_33273 (I568539,I568522,I520644);
nand I_33274 (I568556,I568539,I520662);
nor I_33275 (I568573,I568522,I568556);
DFFARX1 I_33276 (I568573,I2859,I568375,I568340,);
not I_33277 (I568604,I568556);
nand I_33278 (I568621,I568426,I568604);
nand I_33279 (I568352,I568488,I568604);
DFFARX1 I_33280 (I568522,I2859,I568375,I568367,);
not I_33281 (I568666,I520638);
nor I_33282 (I568683,I568666,I520644);
nor I_33283 (I568700,I568683,I568505);
DFFARX1 I_33284 (I568700,I2859,I568375,I568364,);
not I_33285 (I568731,I568683);
DFFARX1 I_33286 (I568731,I2859,I568375,I568757,);
not I_33287 (I568765,I568757);
nor I_33288 (I568361,I568765,I568683);
nor I_33289 (I568796,I568666,I520641);
and I_33290 (I568813,I568796,I520650);
or I_33291 (I568830,I568813,I520659);
DFFARX1 I_33292 (I568830,I2859,I568375,I568856,);
not I_33293 (I568864,I568856);
nand I_33294 (I568881,I568864,I568604);
not I_33295 (I568355,I568881);
nand I_33296 (I568349,I568881,I568621);
nand I_33297 (I568346,I568864,I568488);
not I_33298 (I568970,I2866);
DFFARX1 I_33299 (I287453,I2859,I568970,I568996,);
DFFARX1 I_33300 (I287435,I2859,I568970,I569013,);
not I_33301 (I569021,I569013);
nor I_33302 (I568938,I568996,I569021);
DFFARX1 I_33303 (I569021,I2859,I568970,I568953,);
nor I_33304 (I569066,I287441,I287444);
and I_33305 (I569083,I569066,I287432);
nor I_33306 (I569100,I569083,I287441);
not I_33307 (I569117,I287441);
and I_33308 (I569134,I569117,I287450);
nand I_33309 (I569151,I569134,I287438);
nor I_33310 (I569168,I569117,I569151);
DFFARX1 I_33311 (I569168,I2859,I568970,I568935,);
not I_33312 (I569199,I569151);
nand I_33313 (I569216,I569021,I569199);
nand I_33314 (I568947,I569083,I569199);
DFFARX1 I_33315 (I569117,I2859,I568970,I568962,);
not I_33316 (I569261,I287435);
nor I_33317 (I569278,I569261,I287450);
nor I_33318 (I569295,I569278,I569100);
DFFARX1 I_33319 (I569295,I2859,I568970,I568959,);
not I_33320 (I569326,I569278);
DFFARX1 I_33321 (I569326,I2859,I568970,I569352,);
not I_33322 (I569360,I569352);
nor I_33323 (I568956,I569360,I569278);
nor I_33324 (I569391,I569261,I287447);
and I_33325 (I569408,I569391,I287456);
or I_33326 (I569425,I569408,I287432);
DFFARX1 I_33327 (I569425,I2859,I568970,I569451,);
not I_33328 (I569459,I569451);
nand I_33329 (I569476,I569459,I569199);
not I_33330 (I568950,I569476);
nand I_33331 (I568944,I569476,I569216);
nand I_33332 (I568941,I569459,I569083);
not I_33333 (I569565,I2866);
DFFARX1 I_33334 (I107827,I2859,I569565,I569591,);
DFFARX1 I_33335 (I107830,I2859,I569565,I569608,);
not I_33336 (I569616,I569608);
nor I_33337 (I569533,I569591,I569616);
DFFARX1 I_33338 (I569616,I2859,I569565,I569548,);
nor I_33339 (I569661,I107836,I107830);
and I_33340 (I569678,I569661,I107833);
nor I_33341 (I569695,I569678,I107836);
not I_33342 (I569712,I107836);
and I_33343 (I569729,I569712,I107827);
nand I_33344 (I569746,I569729,I107845);
nor I_33345 (I569763,I569712,I569746);
DFFARX1 I_33346 (I569763,I2859,I569565,I569530,);
not I_33347 (I569794,I569746);
nand I_33348 (I569811,I569616,I569794);
nand I_33349 (I569542,I569678,I569794);
DFFARX1 I_33350 (I569712,I2859,I569565,I569557,);
not I_33351 (I569856,I107839);
nor I_33352 (I569873,I569856,I107827);
nor I_33353 (I569890,I569873,I569695);
DFFARX1 I_33354 (I569890,I2859,I569565,I569554,);
not I_33355 (I569921,I569873);
DFFARX1 I_33356 (I569921,I2859,I569565,I569947,);
not I_33357 (I569955,I569947);
nor I_33358 (I569551,I569955,I569873);
nor I_33359 (I569986,I569856,I107842);
and I_33360 (I570003,I569986,I107848);
or I_33361 (I570020,I570003,I107851);
DFFARX1 I_33362 (I570020,I2859,I569565,I570046,);
not I_33363 (I570054,I570046);
nand I_33364 (I570071,I570054,I569794);
not I_33365 (I569545,I570071);
nand I_33366 (I569539,I570071,I569811);
nand I_33367 (I569536,I570054,I569678);
not I_33368 (I570160,I2866);
DFFARX1 I_33369 (I24310,I2859,I570160,I570186,);
DFFARX1 I_33370 (I24298,I2859,I570160,I570203,);
not I_33371 (I570211,I570203);
nor I_33372 (I570128,I570186,I570211);
DFFARX1 I_33373 (I570211,I2859,I570160,I570143,);
nor I_33374 (I570256,I24289,I24313);
and I_33375 (I570273,I570256,I24292);
nor I_33376 (I570290,I570273,I24289);
not I_33377 (I570307,I24289);
and I_33378 (I570324,I570307,I24295);
nand I_33379 (I570341,I570324,I24307);
nor I_33380 (I570358,I570307,I570341);
DFFARX1 I_33381 (I570358,I2859,I570160,I570125,);
not I_33382 (I570389,I570341);
nand I_33383 (I570406,I570211,I570389);
nand I_33384 (I570137,I570273,I570389);
DFFARX1 I_33385 (I570307,I2859,I570160,I570152,);
not I_33386 (I570451,I24289);
nor I_33387 (I570468,I570451,I24295);
nor I_33388 (I570485,I570468,I570290);
DFFARX1 I_33389 (I570485,I2859,I570160,I570149,);
not I_33390 (I570516,I570468);
DFFARX1 I_33391 (I570516,I2859,I570160,I570542,);
not I_33392 (I570550,I570542);
nor I_33393 (I570146,I570550,I570468);
nor I_33394 (I570581,I570451,I24292);
and I_33395 (I570598,I570581,I24301);
or I_33396 (I570615,I570598,I24304);
DFFARX1 I_33397 (I570615,I2859,I570160,I570641,);
not I_33398 (I570649,I570641);
nand I_33399 (I570666,I570649,I570389);
not I_33400 (I570140,I570666);
nand I_33401 (I570134,I570666,I570406);
nand I_33402 (I570131,I570649,I570273);
not I_33403 (I570755,I2866);
DFFARX1 I_33404 (I244681,I2859,I570755,I570781,);
DFFARX1 I_33405 (I244675,I2859,I570755,I570798,);
not I_33406 (I570806,I570798);
nor I_33407 (I570723,I570781,I570806);
DFFARX1 I_33408 (I570806,I2859,I570755,I570738,);
nor I_33409 (I570851,I244672,I244663);
and I_33410 (I570868,I570851,I244660);
nor I_33411 (I570885,I570868,I244672);
not I_33412 (I570902,I244672);
and I_33413 (I570919,I570902,I244666);
nand I_33414 (I570936,I570919,I244678);
nor I_33415 (I570953,I570902,I570936);
DFFARX1 I_33416 (I570953,I2859,I570755,I570720,);
not I_33417 (I570984,I570936);
nand I_33418 (I571001,I570806,I570984);
nand I_33419 (I570732,I570868,I570984);
DFFARX1 I_33420 (I570902,I2859,I570755,I570747,);
not I_33421 (I571046,I244684);
nor I_33422 (I571063,I571046,I244666);
nor I_33423 (I571080,I571063,I570885);
DFFARX1 I_33424 (I571080,I2859,I570755,I570744,);
not I_33425 (I571111,I571063);
DFFARX1 I_33426 (I571111,I2859,I570755,I571137,);
not I_33427 (I571145,I571137);
nor I_33428 (I570741,I571145,I571063);
nor I_33429 (I571176,I571046,I244663);
and I_33430 (I571193,I571176,I244669);
or I_33431 (I571210,I571193,I244660);
DFFARX1 I_33432 (I571210,I2859,I570755,I571236,);
not I_33433 (I571244,I571236);
nand I_33434 (I571261,I571244,I570984);
not I_33435 (I570735,I571261);
nand I_33436 (I570729,I571261,I571001);
nand I_33437 (I570726,I571244,I570868);
not I_33438 (I571350,I2866);
DFFARX1 I_33439 (I504114,I2859,I571350,I571376,);
DFFARX1 I_33440 (I504117,I2859,I571350,I571393,);
not I_33441 (I571401,I571393);
nor I_33442 (I571318,I571376,I571401);
DFFARX1 I_33443 (I571401,I2859,I571350,I571333,);
nor I_33444 (I571446,I504117,I504132);
and I_33445 (I571463,I571446,I504126);
nor I_33446 (I571480,I571463,I504117);
not I_33447 (I571497,I504117);
and I_33448 (I571514,I571497,I504135);
nand I_33449 (I571531,I571514,I504123);
nor I_33450 (I571548,I571497,I571531);
DFFARX1 I_33451 (I571548,I2859,I571350,I571315,);
not I_33452 (I571579,I571531);
nand I_33453 (I571596,I571401,I571579);
nand I_33454 (I571327,I571463,I571579);
DFFARX1 I_33455 (I571497,I2859,I571350,I571342,);
not I_33456 (I571641,I504129);
nor I_33457 (I571658,I571641,I504135);
nor I_33458 (I571675,I571658,I571480);
DFFARX1 I_33459 (I571675,I2859,I571350,I571339,);
not I_33460 (I571706,I571658);
DFFARX1 I_33461 (I571706,I2859,I571350,I571732,);
not I_33462 (I571740,I571732);
nor I_33463 (I571336,I571740,I571658);
nor I_33464 (I571771,I571641,I504114);
and I_33465 (I571788,I571771,I504138);
or I_33466 (I571805,I571788,I504120);
DFFARX1 I_33467 (I571805,I2859,I571350,I571831,);
not I_33468 (I571839,I571831);
nand I_33469 (I571856,I571839,I571579);
not I_33470 (I571330,I571856);
nand I_33471 (I571324,I571856,I571596);
nand I_33472 (I571321,I571839,I571463);
not I_33473 (I571945,I2866);
DFFARX1 I_33474 (I66177,I2859,I571945,I571971,);
DFFARX1 I_33475 (I66180,I2859,I571945,I571988,);
not I_33476 (I571996,I571988);
nor I_33477 (I571913,I571971,I571996);
DFFARX1 I_33478 (I571996,I2859,I571945,I571928,);
nor I_33479 (I572041,I66186,I66180);
and I_33480 (I572058,I572041,I66183);
nor I_33481 (I572075,I572058,I66186);
not I_33482 (I572092,I66186);
and I_33483 (I572109,I572092,I66177);
nand I_33484 (I572126,I572109,I66195);
nor I_33485 (I572143,I572092,I572126);
DFFARX1 I_33486 (I572143,I2859,I571945,I571910,);
not I_33487 (I572174,I572126);
nand I_33488 (I572191,I571996,I572174);
nand I_33489 (I571922,I572058,I572174);
DFFARX1 I_33490 (I572092,I2859,I571945,I571937,);
not I_33491 (I572236,I66189);
nor I_33492 (I572253,I572236,I66177);
nor I_33493 (I572270,I572253,I572075);
DFFARX1 I_33494 (I572270,I2859,I571945,I571934,);
not I_33495 (I572301,I572253);
DFFARX1 I_33496 (I572301,I2859,I571945,I572327,);
not I_33497 (I572335,I572327);
nor I_33498 (I571931,I572335,I572253);
nor I_33499 (I572366,I572236,I66192);
and I_33500 (I572383,I572366,I66198);
or I_33501 (I572400,I572383,I66201);
DFFARX1 I_33502 (I572400,I2859,I571945,I572426,);
not I_33503 (I572434,I572426);
nand I_33504 (I572451,I572434,I572174);
not I_33505 (I571925,I572451);
nand I_33506 (I571919,I572451,I572191);
nand I_33507 (I571916,I572434,I572058);
not I_33508 (I572540,I2866);
DFFARX1 I_33509 (I200120,I2859,I572540,I572566,);
DFFARX1 I_33510 (I200123,I2859,I572540,I572583,);
not I_33511 (I572591,I572583);
nor I_33512 (I572508,I572566,I572591);
DFFARX1 I_33513 (I572591,I2859,I572540,I572523,);
nor I_33514 (I572636,I200126,I200144);
and I_33515 (I572653,I572636,I200129);
nor I_33516 (I572670,I572653,I200126);
not I_33517 (I572687,I200126);
and I_33518 (I572704,I572687,I200138);
nand I_33519 (I572721,I572704,I200141);
nor I_33520 (I572738,I572687,I572721);
DFFARX1 I_33521 (I572738,I2859,I572540,I572505,);
not I_33522 (I572769,I572721);
nand I_33523 (I572786,I572591,I572769);
nand I_33524 (I572517,I572653,I572769);
DFFARX1 I_33525 (I572687,I2859,I572540,I572532,);
not I_33526 (I572831,I200132);
nor I_33527 (I572848,I572831,I200138);
nor I_33528 (I572865,I572848,I572670);
DFFARX1 I_33529 (I572865,I2859,I572540,I572529,);
not I_33530 (I572896,I572848);
DFFARX1 I_33531 (I572896,I2859,I572540,I572922,);
not I_33532 (I572930,I572922);
nor I_33533 (I572526,I572930,I572848);
nor I_33534 (I572961,I572831,I200120);
and I_33535 (I572978,I572961,I200135);
or I_33536 (I572995,I572978,I200123);
DFFARX1 I_33537 (I572995,I2859,I572540,I573021,);
not I_33538 (I573029,I573021);
nand I_33539 (I573046,I573029,I572769);
not I_33540 (I572520,I573046);
nand I_33541 (I572514,I573046,I572786);
nand I_33542 (I572511,I573029,I572653);
not I_33543 (I573135,I2866);
DFFARX1 I_33544 (I203095,I2859,I573135,I573161,);
DFFARX1 I_33545 (I203098,I2859,I573135,I573178,);
not I_33546 (I573186,I573178);
nor I_33547 (I573103,I573161,I573186);
DFFARX1 I_33548 (I573186,I2859,I573135,I573118,);
nor I_33549 (I573231,I203101,I203119);
and I_33550 (I573248,I573231,I203104);
nor I_33551 (I573265,I573248,I203101);
not I_33552 (I573282,I203101);
and I_33553 (I573299,I573282,I203113);
nand I_33554 (I573316,I573299,I203116);
nor I_33555 (I573333,I573282,I573316);
DFFARX1 I_33556 (I573333,I2859,I573135,I573100,);
not I_33557 (I573364,I573316);
nand I_33558 (I573381,I573186,I573364);
nand I_33559 (I573112,I573248,I573364);
DFFARX1 I_33560 (I573282,I2859,I573135,I573127,);
not I_33561 (I573426,I203107);
nor I_33562 (I573443,I573426,I203113);
nor I_33563 (I573460,I573443,I573265);
DFFARX1 I_33564 (I573460,I2859,I573135,I573124,);
not I_33565 (I573491,I573443);
DFFARX1 I_33566 (I573491,I2859,I573135,I573517,);
not I_33567 (I573525,I573517);
nor I_33568 (I573121,I573525,I573443);
nor I_33569 (I573556,I573426,I203095);
and I_33570 (I573573,I573556,I203110);
or I_33571 (I573590,I573573,I203098);
DFFARX1 I_33572 (I573590,I2859,I573135,I573616,);
not I_33573 (I573624,I573616);
nand I_33574 (I573641,I573624,I573364);
not I_33575 (I573115,I573641);
nand I_33576 (I573109,I573641,I573381);
nand I_33577 (I573106,I573624,I573248);
not I_33578 (I573730,I2866);
DFFARX1 I_33579 (I171832,I2859,I573730,I573756,);
DFFARX1 I_33580 (I171838,I2859,I573730,I573773,);
not I_33581 (I573781,I573773);
nor I_33582 (I573698,I573756,I573781);
DFFARX1 I_33583 (I573781,I2859,I573730,I573713,);
nor I_33584 (I573826,I171847,I171832);
and I_33585 (I573843,I573826,I171859);
nor I_33586 (I573860,I573843,I171847);
not I_33587 (I573877,I171847);
and I_33588 (I573894,I573877,I171835);
nand I_33589 (I573911,I573894,I171856);
nor I_33590 (I573928,I573877,I573911);
DFFARX1 I_33591 (I573928,I2859,I573730,I573695,);
not I_33592 (I573959,I573911);
nand I_33593 (I573976,I573781,I573959);
nand I_33594 (I573707,I573843,I573959);
DFFARX1 I_33595 (I573877,I2859,I573730,I573722,);
not I_33596 (I574021,I171844);
nor I_33597 (I574038,I574021,I171835);
nor I_33598 (I574055,I574038,I573860);
DFFARX1 I_33599 (I574055,I2859,I573730,I573719,);
not I_33600 (I574086,I574038);
DFFARX1 I_33601 (I574086,I2859,I573730,I574112,);
not I_33602 (I574120,I574112);
nor I_33603 (I573716,I574120,I574038);
nor I_33604 (I574151,I574021,I171841);
and I_33605 (I574168,I574151,I171853);
or I_33606 (I574185,I574168,I171850);
DFFARX1 I_33607 (I574185,I2859,I573730,I574211,);
not I_33608 (I574219,I574211);
nand I_33609 (I574236,I574219,I573959);
not I_33610 (I573710,I574236);
nand I_33611 (I573704,I574236,I573976);
nand I_33612 (I573701,I574219,I573843);
endmodule


