module test_I3211(I1902,I1294,I3447,I1301,I3211);
input I1902,I1294,I3447,I1301;
output I3211;
wire I3263,I3464,I3512,I3481,I2962,I2583,I2575,I2569,I3246,I2566,I2945,I3543,I2832;
not I_0(I3263,I2569);
or I_1(I3464,I3447,I2575);
DFFARX1 I_2(I3481,I1294,I3246,,,I3512,);
DFFARX1 I_3(I3464,I1294,I3246,,,I3481,);
and I_4(I3211,I3543,I3512);
nor I_5(I2962,I2945);
not I_6(I2583,I1301);
DFFARX1 I_7(I1294,I2583,,,I2575,);
nand I_8(I2569,I2832,I2962);
not I_9(I3246,I1301);
not I_10(I2566,I2945);
DFFARX1 I_11(I1902,I1294,I2583,,,I2945,);
nand I_12(I3543,I3263,I2566);
DFFARX1 I_13(I1294,I2583,,,I2832,);
endmodule


