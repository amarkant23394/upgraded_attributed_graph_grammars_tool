module test_I3263(I2798,I1917,I2651,I1902,I1294,I1301,I3263);
input I2798,I1917,I2651,I1902,I1294,I1301;
output I3263;
wire I2815,I2668,I1914,I2583,I2569,I2962,I2945,I2832;
not I_0(I3263,I2569);
or I_1(I2815,I2798,I1917);
nand I_2(I2668,I2651,I1914);
DFFARX1 I_3(I1294,,,I1914,);
not I_4(I2583,I1301);
nand I_5(I2569,I2832,I2962);
nor I_6(I2962,I2945,I2668);
DFFARX1 I_7(I1902,I1294,I2583,,,I2945,);
DFFARX1 I_8(I2815,I1294,I2583,,,I2832,);
endmodule


