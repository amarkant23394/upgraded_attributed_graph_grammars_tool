module test_I2311(I1287,I1231,I2311);
input I1287,I1231;
output I2311;
wire I2294;
nor I_0(I2294,I1287,I1231);
not I_1(I2311,I2294);
endmodule


