module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_8_r_10,n11_10,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_8_r_10,n11_10,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
nor I_40(N1371_0_r_10,n37_10,n38_10);
nor I_41(N1508_0_r_10,n37_10,n58_10);
nand I_42(N6147_2_r_10,n39_10,n40_10);
not I_43(N6147_3_r_10,n39_10);
nor I_44(N1372_4_r_10,n46_10,n49_10);
nor I_45(N1508_4_r_10,n51_10,n52_10);
nor I_46(N1507_6_r_10,n49_10,n60_10);
nor I_47(N1508_6_r_10,n49_10,n50_10);
nor I_48(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_49(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_50(N6147_9_r_10,n36_10,n37_10);
nor I_51(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_52(I_BUFF_1_9_r_10,n48_10);
nor I_53(N3_8_r_10,n44_10,n47_10);
not I_54(n11_10,blif_reset_net_8_r_10);
not I_55(n35_10,n49_10);
nor I_56(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_57(n37_10,N1508_10_r_8);
not I_58(n38_10,n46_10);
nand I_59(n39_10,n43_10,n44_10);
nand I_60(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_61(n41_10,n42_10,N1508_10_r_8);
not I_62(n42_10,n44_10);
nor I_63(n43_10,n45_10,N1508_10_r_8);
nand I_64(n44_10,n54_10,N1508_6_r_8);
nor I_65(n45_10,n59_10,G199_8_r_8);
nand I_66(n46_10,n61_10,n_42_8_r_8);
nor I_67(n47_10,n46_10,n48_10);
nand I_68(n48_10,n62_10,n63_10);
nand I_69(n49_10,n56_10,N1508_1_r_8);
not I_70(n50_10,n45_10);
nor I_71(n51_10,n42_10,n53_10);
not I_72(n52_10,N1372_4_r_10);
nor I_73(n53_10,n48_10,n50_10);
and I_74(n54_10,n55_10,G199_8_r_8);
nand I_75(n55_10,n56_10,n57_10);
nand I_76(n56_10,N1507_6_r_8,N6147_9_r_8);
not I_77(n57_10,N1508_1_r_8);
nor I_78(n58_10,n35_10,n45_10);
nor I_79(n59_10,N1371_0_r_8,N1508_1_r_8);
nor I_80(n60_10,n37_10,n46_10);
or I_81(n61_10,N1371_0_r_8,N1508_1_r_8);
nor I_82(n62_10,N6147_9_r_8,N6134_9_r_8);
or I_83(n63_10,n64_10,N1507_6_r_8);
nor I_84(n64_10,N1508_6_r_8,n_42_8_r_8);
endmodule


