module test_I2827(I1407,I1351,I2827);
input I1407,I1351;
output I2827;
wire I2776;
not I_0(I2776,I1407);
nor I_1(I2827,I2776,I1351);
endmodule


