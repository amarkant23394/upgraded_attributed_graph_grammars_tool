module test_I15143(I10647,I10961,I1470,I15143);
input I10647,I10961,I1470;
output I15143;
wire I12913,I12930,I12718,I10615,I10639,I12599,I11201,I12964,I12882,I12848,I10609;
DFFARX1 I_0(I1470,,,I12913,);
and I_1(I12930,I12913,I10609);
nor I_2(I12718,I10615,I10639);
DFFARX1 I_3(I10961,I1470,I10647,,,I10615,);
DFFARX1 I_4(I11201,I1470,I10647,,,I10639,);
nand I_5(I12599,I12718,I12964);
not I_6(I15143,I12599);
and I_7(I11201,I10961);
nor I_8(I12964,I12930,I12882);
not I_9(I12882,I12848);
DFFARX1 I_10(I1470,,,I12848,);
DFFARX1 I_11(I1470,I10647,,,I10609,);
endmodule


