module test_I8998(I6924,I5642,I5368,I5070,I8998);
input I6924,I5642,I5368,I5070;
output I8998;
wire I7026,I7057,I6975,I6881,I6992,I5097;
not I_0(I7026,I5070);
not I_1(I7057,I7026);
nor I_2(I6975,I6924,I5070);
nand I_3(I6881,I6992,I7057);
nand I_4(I6992,I6975,I5097);
not I_5(I8998,I6881);
nand I_6(I5097,I5642,I5368);
endmodule


