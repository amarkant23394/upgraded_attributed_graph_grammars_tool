module test_final(IN_1_0_l_5,IN_2_0_l_5,IN_3_0_l_5,IN_4_0_l_5,IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0);
input IN_1_0_l_5,IN_2_0_l_5,IN_3_0_l_5,IN_4_0_l_5,IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0;
wire N1371_0_r_5,N1508_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1507_6_r_5,N1508_6_r_5,n_431_5_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,N1508_0_r_0,n_102_5_r_0,N3_8_l_0,n5_0,n40_0,n4_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0;
nor I_0(N1371_0_r_5,n28_5,n39_5);
not I_1(N1508_0_r_5,n39_5);
nor I_2(N6147_2_r_5,n28_5,n37_5);
nand I_3(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_4(n_431_5_r_5,blif_clk_net_5_r_0,n5_0,G78_5_r_5,);
nand I_5(n_576_5_r_5,n26_5,n27_5);
not I_6(n_102_5_r_5,n28_5);
nand I_7(n_547_5_r_5,n31_5,n32_5);
nor I_8(N1507_6_r_5,n30_5,n32_5);
nor I_9(N1508_6_r_5,n39_5,n41_5);
nand I_10(n_431_5_r_5,n34_5,n35_5);
nor I_11(n26_5,n29_5,n30_5);
nor I_12(n27_5,IN_2_0_l_5,n28_5);
nor I_13(n28_5,n29_5,n44_5);
not I_14(n29_5,IN_1_0_l_5);
nand I_15(n30_5,N1508_0_r_5,n43_5);
nor I_16(n31_5,n28_5,n33_5);
nor I_17(n32_5,IN_3_1_l_5,n40_5);
nor I_18(n33_5,IN_2_0_l_5,n29_5);
or I_19(n34_5,IN_2_0_l_5,n29_5);
nand I_20(n35_5,n32_5,n36_5);
not I_21(n36_5,n30_5);
nor I_22(n37_5,N1507_6_r_5,n38_5);
and I_23(n38_5,n39_5,n40_5);
nand I_24(n39_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_25(n40_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_26(n41_5,n28_5,n42_5);
or I_27(n42_5,n32_5,n36_5);
or I_28(n43_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_29(n44_5,IN_3_0_l_5,IN_4_0_l_5);
nor I_30(N1371_0_r_0,n24_0,n25_0);
not I_31(N1508_0_r_0,n25_0);
nor I_32(N6147_2_r_0,n28_0,n29_0);
nand I_33(n_429_or_0_5_r_0,n4_0,n25_0);
DFFARX1 I_34(n4_0,blif_clk_net_5_r_0,n5_0,G78_5_r_0,);
nand I_35(n_576_5_r_0,n23_0,n24_0);
not I_36(n_102_5_r_0,n40_0);
nand I_37(n_547_5_r_0,n26_0,n27_0);
nor I_38(N1507_6_r_0,n_102_5_r_0,n37_0);
nor I_39(N1508_6_r_0,n25_0,n33_0);
and I_40(N3_8_l_0,n32_0,n_429_or_0_5_r_5);
not I_41(n5_0,blif_reset_net_5_r_0);
DFFARX1 I_42(N3_8_l_0,blif_clk_net_5_r_0,n5_0,n40_0,);
not I_43(n4_0,n31_0);
nor I_44(n23_0,n40_0,n25_0);
and I_45(n24_0,n4_0,n39_0);
nand I_46(n25_0,G78_5_r_5,n_576_5_r_5);
nor I_47(n26_0,n40_0,n24_0);
nor I_48(n27_0,N1508_6_r_5,N6147_2_r_5);
nor I_49(n28_0,n25_0,N6147_2_r_5);
nand I_50(n29_0,n_102_5_r_0,n30_0);
nand I_51(n30_0,n27_0,n31_0);
nand I_52(n31_0,n_102_5_r_5,n_547_5_r_5);
nand I_53(n32_0,N1371_0_r_5,N6147_2_r_5);
nand I_54(n33_0,n34_0,n35_0);
nand I_55(n34_0,n_102_5_r_0,n36_0);
not I_56(n35_0,N6147_2_r_5);
not I_57(n36_0,n27_0);
nor I_58(n37_0,n36_0,n38_0);
nand I_59(n38_0,N1508_0_r_0,n35_0);
or I_60(n39_0,n_429_or_0_5_r_5,N1371_0_r_5);
endmodule


