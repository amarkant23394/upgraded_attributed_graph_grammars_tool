module test_I6843(I2742,I4017,I1477,I1470,I6843);
input I2742,I4017,I1477,I1470;
output I6843;
wire I6781,I3975,I3966,I3954,I6826,I6442,I6329,I6493,I4068,I4308,I4034,I4130,I3957,I2724,I3983;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
nor I_1(I3975,I4308,I4034);
or I_2(I3966,I4068,I4034);
not I_3(I3954,I4068);
nand I_4(I6826,I6781,I6442);
nor I_5(I6442,I3975,I3954);
not I_6(I6329,I1477);
DFFARX1 I_7(I3966,I1470,I6329,,,I6493,);
and I_8(I6843,I6493,I6826);
nor I_9(I4068,I2742,I2724);
DFFARX1 I_10(I1470,I3983,,,I4308,);
DFFARX1 I_11(I4017,I1470,I3983,,,I4034,);
nor I_12(I4130,I4068);
nand I_13(I3957,I4308,I4130);
DFFARX1 I_14(I1470,,,I2724,);
not I_15(I3983,I1477);
endmodule


