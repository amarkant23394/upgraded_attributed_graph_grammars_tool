module test_I1483(I1383,I1477,I1470,I1483);
input I1383,I1477,I1470;
output I1483;
wire I1518,I1880;
not I_0(I1518,I1477);
DFFARX1 I_1(I1383,I1470,I1518,,,I1880,);
DFFARX1 I_2(I1880,I1470,I1518,,,I1483,);
endmodule


