module test_I8862(I1477,I8862);
input I1477;
output I8862;
wire ;
not I_0(I8862,I1477);
endmodule


