module test_I1307(I1215,I1294,I1301,I1307);
input I1215,I1294,I1301;
output I1307;
wire I1873,I1342,I1780;
DFFARX1 I_0(I1780,I1294,I1342,,,I1873,);
not I_1(I1342,I1301);
and I_2(I1307,I1780,I1873);
DFFARX1 I_3(I1215,I1294,I1342,,,I1780,);
endmodule


