module test_final(IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5,N3_2_l_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_5,blif_clk_net_1_r_8,n8_8,G42_1_r_5,);
nor I_1(n_572_1_r_5,n21_5,n22_5);
nand I_2(n_573_1_r_5,n13_5,n16_5);
nor I_3(n_549_1_r_5,n21_5,n17_5);
nand I_4(n_569_1_r_5,n13_5,n15_5);
nor I_5(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_6(G199_2_l_5,blif_clk_net_1_r_8,n8_8,ACVQN2_3_r_5,);
nor I_7(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_8(n_42_2_l_5,blif_clk_net_1_r_8,n8_8,ACVQN1_5_r_5,);
not I_9(P6_5_r_5,P6_5_r_internal_5);
and I_10(N3_2_l_5,IN_6_2_l_5,n19_5);
DFFARX1 I_11(N3_2_l_5,blif_clk_net_1_r_8,n8_8,G199_2_l_5,);
DFFARX1 I_12(IN_1_3_l_5,blif_clk_net_1_r_8,n8_8,ACVQN2_3_l_5,);
not I_13(n13_5,ACVQN2_3_l_5);
DFFARX1 I_14(IN_2_3_l_5,blif_clk_net_1_r_8,n8_8,ACVQN1_3_l_5,);
and I_15(N1_4_l_5,IN_6_4_l_5,n20_5);
DFFARX1 I_16(N1_4_l_5,blif_clk_net_1_r_8,n8_8,n21_5,);
not I_17(n15_5,n21_5);
DFFARX1 I_18(IN_3_4_l_5,blif_clk_net_1_r_8,n8_8,n22_5,);
nor I_19(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_20(ACVQN2_3_l_5,blif_clk_net_1_r_8,n8_8,n11_internal_5,);
not I_21(n11_5,n11_internal_5);
nor I_22(n_42_2_l_5,IN_1_2_l_5,IN_3_2_l_5);
not I_23(n1_5,n18_5);
DFFARX1 I_24(n1_5,blif_clk_net_1_r_8,n8_8,P6_5_r_internal_5,);
not I_25(n16_5,n_42_2_l_5);
nor I_26(n17_5,n22_5,n18_5);
nand I_27(n18_5,IN_4_3_l_5,ACVQN1_3_l_5);
nand I_28(n19_5,IN_2_2_l_5,IN_3_2_l_5);
nand I_29(n20_5,IN_1_4_l_5,IN_2_4_l_5);
DFFARX1 I_30(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_31(n_572_1_r_8,n39_8,n23_8);
and I_32(n_549_1_r_8,n38_8,n23_8);
nand I_33(n_569_1_r_8,n38_8,n24_8);
nor I_34(n_452_1_r_8,n25_8,n26_8);
nor I_35(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_36(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_37(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_38(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_39(n_431_0_l_8,n29_8,n_569_1_r_5);
not I_40(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_41(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_42(n19_8,G78_0_l_8);
DFFARX1 I_43(n_573_1_r_5,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_44(n22_8,n39_8);
DFFARX1 I_45(n_266_and_0_3_r_5,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_46(n4_1_r_8,G78_0_l_8,n33_8);
nor I_47(N3_2_r_8,n22_8,n35_8);
nor I_48(N1_4_r_8,n27_8,n37_8);
nand I_49(n23_8,n32_8,G42_1_r_5);
not I_50(n24_8,n23_8);
nand I_51(n25_8,n36_8,n_572_1_r_5);
nand I_52(n26_8,n27_8,n28_8);
nor I_53(n27_8,n31_8,n_549_1_r_5);
not I_54(n28_8,P6_5_r_5);
and I_55(n29_8,n30_8,ACVQN2_3_r_5);
nor I_56(n30_8,n31_8,n_452_1_r_5);
not I_57(n31_8,G42_1_r_5);
and I_58(n32_8,n28_8,n_549_1_r_5);
nand I_59(n33_8,n28_8,n34_8);
not I_60(n34_8,n25_8);
nor I_61(n35_8,n34_8,P6_5_r_5);
not I_62(n36_8,ACVQN1_5_r_5);
nor I_63(n37_8,n19_8,n38_8);
endmodule


