module test_I16232(I1477,I1470,I14356,I14605,I16232);
input I1477,I1470,I14356,I14605;
output I16232;
wire I14338,I16356,I16339,I16240,I16661,I14347,I14353,I16678,I14808,I16644,I14370;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
DFFARX1 I_1(I14356,I1470,I16240,,,I16356,);
nor I_2(I16339,I14353,I14338);
DFFARX1 I_3(I16678,I1470,I16240,,,I16232,);
not I_4(I16240,I1477);
nand I_5(I16661,I16644,I16356);
DFFARX1 I_6(I1470,I14370,,,I14347,);
not I_7(I14353,I14808);
and I_8(I16678,I16339,I16661);
DFFARX1 I_9(I1470,I14370,,,I14808,);
DFFARX1 I_10(I14347,I1470,I16240,,,I16644,);
not I_11(I14370,I1477);
endmodule


