module test_I7535(I6826,I1477,I1470,I6705,I7535);
input I6826,I1477,I1470,I6705;
output I7535;
wire I6297,I6300,I7946,I7714,I7881,I7570,I6329,I7587,I6843,I6493,I6291;
DFFARX1 I_0(I6843,I1470,I6329,,,I6297,);
DFFARX1 I_1(I1470,I6329,,,I6300,);
DFFARX1 I_2(I7881,I1470,I7570,,,I7946,);
not I_3(I7714,I6297);
nand I_4(I7881,I7587,I6291);
not I_5(I7570,I1477);
not I_6(I6329,I1477);
not I_7(I7587,I6300);
and I_8(I7535,I7714,I7946);
and I_9(I6843,I6493,I6826);
DFFARX1 I_10(I1470,I6329,,,I6493,);
DFFARX1 I_11(I6705,I1470,I6329,,,I6291,);
endmodule


