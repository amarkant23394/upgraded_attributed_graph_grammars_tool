module test_I2651(I1316,I2406,I1294,I1301,I2651);
input I1316,I2406,I1294,I1301;
output I2651;
wire I2600,I1911,I2005,I1937,I2022,I2039,I1908,I2070,I1310,I2488;
not I_0(I2600,I1911);
nand I_1(I1911,I2070,I2488);
nor I_2(I2005,I1310);
nor I_3(I2651,I2600,I1908);
not I_4(I1937,I1301);
nand I_5(I2022,I2005,I1316);
DFFARX1 I_6(I2022,I1294,I1937,,,I2039,);
not I_7(I1908,I2039);
not I_8(I2070,I1310);
DFFARX1 I_9(I1294,,,I1310,);
not I_10(I2488,I2406);
endmodule


