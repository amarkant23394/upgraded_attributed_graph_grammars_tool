module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_8_r_6,n9_6,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_6,n30_6,n33_6);
nor I_37(N1508_0_r_6,n33_6,n44_6);
not I_38(N1372_1_r_6,n41_6);
nor I_39(N1508_1_r_6,n40_6,n41_6);
nor I_40(N1507_6_r_6,n39_6,n45_6);
nor I_41(N1508_6_r_6,n37_6,n38_6);
nor I_42(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_43(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_44(N6147_9_r_6,n32_6,n33_6);
nor I_45(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_46(I_BUFF_1_9_r_6,n37_6);
not I_47(N1372_10_r_6,n43_6);
nor I_48(N1508_10_r_6,n42_6,n43_6);
nor I_49(N3_8_r_6,n36_6,N1507_6_r_3);
not I_50(n9_6,blif_reset_net_8_r_6);
nor I_51(n30_6,n53_6,N1372_1_r_3);
not I_52(n31_6,n36_6);
nor I_53(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_54(n33_6,N1507_6_r_3);
not I_55(n34_6,n35_6);
nand I_56(n35_6,n49_6,G42_7_r_3);
nand I_57(n36_6,n51_6,N6134_9_r_3);
nand I_58(n37_6,n54_6,n_452_7_r_3);
or I_59(n38_6,n35_6,n39_6);
nor I_60(n39_6,n40_6,n45_6);
and I_61(n40_6,n46_6,n47_6);
nand I_62(n41_6,n30_6,n31_6);
nor I_63(n42_6,n34_6,n40_6);
nand I_64(n43_6,n30_6,N1507_6_r_3);
nor I_65(n44_6,n31_6,n40_6);
nor I_66(n45_6,n35_6,n36_6);
nor I_67(n46_6,N1372_1_r_3,N1508_1_r_3);
or I_68(n47_6,n48_6,N1508_6_r_3);
nor I_69(n48_6,n_569_7_r_3,N1508_6_r_3);
and I_70(n49_6,n50_6,G42_7_r_3);
nand I_71(n50_6,n51_6,n52_6);
nand I_72(n51_6,N1508_1_r_3,N1507_6_r_3);
not I_73(n52_6,N6134_9_r_3);
nor I_74(n53_6,n_573_7_r_3,n_549_7_r_3);
or I_75(n54_6,n_573_7_r_3,n_549_7_r_3);
endmodule


