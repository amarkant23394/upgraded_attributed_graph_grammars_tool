module test_I4263(I1477,I1359,I2776,I1415,I1447,I1431,I1470,I4263);
input I1477,I1359,I2776,I1415,I1447,I1431,I1470;
output I4263;
wire I2733,I3107,I3076,I2980,I3983,I3200,I3310,I2745,I3217,I3293,I2759,I2844,I2827,I4246;
nand I_0(I2733,I3217,I3107);
nor I_1(I3107,I3076,I2844);
DFFARX1 I_2(I1447,I1470,I2759,,,I3076,);
nand I_3(I2980,I2776,I1415);
not I_4(I3983,I1477);
DFFARX1 I_5(I1431,I1470,I2759,,,I3200,);
and I_6(I4263,I4246,I2733);
and I_7(I3310,I2844,I3293);
nor I_8(I2745,I2980,I3310);
not I_9(I3217,I3200);
not I_10(I3293,I3217);
not I_11(I2759,I1477);
nand I_12(I2844,I2827,I1359);
nor I_13(I2827,I2776);
DFFARX1 I_14(I2745,I1470,I3983,,,I4246,);
endmodule


