module test_final(G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11,n_431_0_l_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_11,blif_clk_net_1_r_3,n9_3,G42_1_r_11,);
nor I_1(n_572_1_r_11,n29_11,n30_11);
nand I_2(n_573_1_r_11,n26_11,n28_11);
nor I_3(n_549_1_r_11,n27_11,n32_11);
nand I_4(n_569_1_r_11,n45_11,n28_11);
nor I_5(n_452_1_r_11,n43_11,n44_11);
nor I_6(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_7(N3_2_r_11,blif_clk_net_1_r_3,n9_3,G199_2_r_11,);
DFFARX1 I_8(n24_11,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_11,);
nor I_9(n_266_and_0_3_r_11,n20_11,n37_11);
or I_10(n_431_0_l_11,IN_8_0_l_11,n33_11);
DFFARX1 I_11(n_431_0_l_11,blif_clk_net_1_r_3,n9_3,n43_11,);
not I_12(n26_11,n43_11);
DFFARX1 I_13(IN_2_5_l_11,blif_clk_net_1_r_3,n9_3,n44_11,);
DFFARX1 I_14(IN_1_5_l_11,blif_clk_net_1_r_3,n9_3,n45_11,);
not I_15(n27_11,n45_11);
nor I_16(n4_1_r_11,n44_11,n25_11);
nor I_17(N3_2_r_11,n45_11,n40_11);
nand I_18(n24_11,IN_11_0_l_11,n39_11);
nand I_19(n25_11,IN_7_0_l_11,n38_11);
DFFARX1 I_20(n25_11,blif_clk_net_1_r_3,n9_3,n20_internal_11,);
not I_21(n20_11,n20_internal_11);
not I_22(n28_11,n25_11);
not I_23(n29_11,G1_0_l_11);
nand I_24(n30_11,n26_11,n31_11);
not I_25(n31_11,IN_5_0_l_11);
and I_26(n32_11,n26_11,n44_11);
and I_27(n33_11,IN_2_0_l_11,n34_11);
nor I_28(n34_11,IN_4_0_l_11,n29_11);
not I_29(n35_11,G2_0_l_11);
nand I_30(n36_11,G1_0_l_11,n31_11);
nor I_31(n37_11,IN_5_0_l_11,n29_11);
nor I_32(n38_11,G2_0_l_11,n31_11);
nor I_33(n39_11,G2_0_l_11,IN_10_0_l_11);
nor I_34(n40_11,G2_0_l_11,n41_11);
nor I_35(n41_11,IN_10_0_l_11,n42_11);
not I_36(n42_11,IN_11_0_l_11);
DFFARX1 I_37(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_38(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_39(n_573_1_r_3,n26_3,n27_3);
nor I_40(n_549_1_r_3,n40_3,n32_3);
nand I_41(n_569_1_r_3,n27_3,n31_3);
and I_42(n_452_1_r_3,n26_3,ACVQN2_3_r_11);
nor I_43(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_44(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_45(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_46(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_47(n4_1_l_3,G42_1_r_11,ACVQN2_3_r_11);
not I_48(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_49(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_50(n22_3,G42_1_l_3);
DFFARX1 I_51(n_569_1_r_11,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_52(n_452_1_r_11,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_53(n25_3,n25_internal_3);
nor I_54(n4_1_r_3,n40_3,n36_3);
nor I_55(N3_2_r_3,n26_3,n37_3);
nor I_56(n_572_1_l_3,n_573_1_r_11,n_549_1_r_11);
DFFARX1 I_57(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_58(n26_3,n_572_1_r_11,G199_2_r_11);
not I_59(n27_3,n_42_2_r_11);
nor I_60(n28_3,n29_3,n_42_2_r_11);
nor I_61(n29_3,n30_3,n_549_1_r_11);
not I_62(n30_3,n_266_and_0_3_r_11);
nor I_63(n31_3,n40_3,n_572_1_r_11);
nor I_64(n32_3,n25_3,n33_3);
nand I_65(n33_3,n22_3,G42_1_r_11);
or I_66(n34_3,n_572_1_r_11,n_42_2_r_11);
nand I_67(n35_3,ACVQN1_3_r_3,G42_1_r_11);
nor I_68(n36_3,G199_2_r_11,ACVQN2_3_r_11);
nor I_69(n37_3,n38_3,n39_3);
not I_70(n38_3,n_572_1_l_3);
nand I_71(n39_3,n27_3,n30_3);
endmodule


