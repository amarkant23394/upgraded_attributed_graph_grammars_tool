module test_I11751(I1477,I9049,I9083,I8947,I6896,I1470,I11751);
input I1477,I9049,I9083,I8947,I6896,I1470;
output I11751;
wire I9320,I8845,I8836,I9179,I8839,I11344,I9337,I9303,I9210,I8862,I8848,I9413,I11672,I11361,I9066,I11310;
not I_0(I9320,I9303);
or I_1(I8845,I9179,I9066);
nand I_2(I8836,I9320,I9210);
DFFARX1 I_3(I6896,I1470,I8862,,,I9179,);
DFFARX1 I_4(I9337,I1470,I8862,,,I8839,);
nor I_5(I11344,I8848,I8839);
nor I_6(I9337,I9320);
DFFARX1 I_7(I1470,I8862,,,I9303,);
nor I_8(I9210,I9179,I8947);
not I_9(I8862,I1477);
nor I_10(I8848,I9083,I9413);
and I_11(I9413,I8947);
DFFARX1 I_12(I8836,I1470,I11310,,,I11672,);
nand I_13(I11361,I11344,I8845);
DFFARX1 I_14(I9049,I1470,I8862,,,I9066,);
not I_15(I11310,I1477);
nand I_16(I11751,I11672,I11361);
endmodule


