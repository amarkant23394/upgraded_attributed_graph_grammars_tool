module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_8_r_6,n9_6,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N1371_0_r_6,n30_6,n33_6);
nor I_42(N1508_0_r_6,n33_6,n44_6);
not I_43(N1372_1_r_6,n41_6);
nor I_44(N1508_1_r_6,n40_6,n41_6);
nor I_45(N1507_6_r_6,n39_6,n45_6);
nor I_46(N1508_6_r_6,n37_6,n38_6);
nor I_47(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_48(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_49(N6147_9_r_6,n32_6,n33_6);
nor I_50(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_51(I_BUFF_1_9_r_6,n37_6);
not I_52(N1372_10_r_6,n43_6);
nor I_53(N1508_10_r_6,n42_6,n43_6);
nor I_54(N3_8_r_6,n36_6,N1508_0_r_1);
not I_55(n9_6,blif_reset_net_8_r_6);
nor I_56(n30_6,n53_6,n_572_7_r_1);
not I_57(n31_6,n36_6);
nor I_58(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_59(n33_6,N1508_0_r_1);
not I_60(n34_6,n35_6);
nand I_61(n35_6,n49_6,G42_7_r_1);
nand I_62(n36_6,n51_6,n_549_7_r_1);
nand I_63(n37_6,n54_6,G42_7_r_1);
or I_64(n38_6,n35_6,n39_6);
nor I_65(n39_6,n40_6,n45_6);
and I_66(n40_6,n46_6,n47_6);
nand I_67(n41_6,n30_6,n31_6);
nor I_68(n42_6,n34_6,n40_6);
nand I_69(n43_6,n30_6,N1508_0_r_1);
nor I_70(n44_6,n31_6,n40_6);
nor I_71(n45_6,n35_6,n36_6);
nor I_72(n46_6,n_572_7_r_1,N1507_6_r_1);
or I_73(n47_6,n48_6,N1508_6_r_1);
nor I_74(n48_6,N1507_6_r_1,n_569_7_r_1);
and I_75(n49_6,n50_6,n_573_7_r_1);
nand I_76(n50_6,n51_6,n52_6);
nand I_77(n51_6,N1508_6_r_1,N6134_9_r_1);
not I_78(n52_6,n_549_7_r_1);
nor I_79(n53_6,N6147_9_r_1,N1508_0_r_1);
or I_80(n54_6,N6147_9_r_1,N1508_0_r_1);
endmodule


