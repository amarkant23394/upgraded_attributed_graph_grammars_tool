module test_final(IN_1_2_l_2,IN_2_2_l_2,G1_3_l_2,G2_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_5_3_l_2,IN_7_3_l_2,IN_8_3_l_2,IN_10_3_l_2,IN_11_3_l_2,blif_clk_net_1_r_5,blif_reset_net_1_r_5,G199_1_r_5,G214_1_r_5,ACVQN1_2_r_5,P6_2_r_5,n_429_or_0_3_r_5,G78_3_r_5,n_576_3_r_5,n_102_3_r_5,n_547_3_r_5,n_42_5_r_5,G199_5_r_5);
input IN_1_2_l_2,IN_2_2_l_2,G1_3_l_2,G2_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_5_3_l_2,IN_7_3_l_2,IN_8_3_l_2,IN_10_3_l_2,IN_11_3_l_2,blif_clk_net_1_r_5,blif_reset_net_1_r_5;
output G199_1_r_5,G214_1_r_5,ACVQN1_2_r_5,P6_2_r_5,n_429_or_0_3_r_5,G78_3_r_5,n_576_3_r_5,n_102_3_r_5,n_547_3_r_5,n_42_5_r_5,G199_5_r_5;
wire ACVQN2_0_r_2,n_266_and_0_0_r_2,G199_1_r_2,G214_1_r_2,n_429_or_0_3_r_2,G78_3_r_2,n_576_3_r_2,n_102_3_r_2,n_547_3_r_2,n_42_5_r_2,G199_5_r_2,ACVQN1_2_l_2,P6_2_l_2,P6_internal_2_l_2,n_429_or_0_3_l_2,n12_3_l_2,n_431_3_l_2,G78_3_l_2,n_576_3_l_2,n11_3_l_2,n_102_3_l_2,n_547_3_l_2,n13_3_l_2,n14_3_l_2,n15_3_l_2,n16_3_l_2,ACVQN1_0_r_2,N1_1_r_2,n3_1_r_2,n12_3_r_2,n_431_3_r_2,n11_3_r_2,n13_3_r_2,n14_3_r_2,n15_3_r_2,n16_3_r_2,N3_5_r_2,n3_5_r_2,n1_1_r_5,ACVQN1_2_l_5,P6_2_l_5,P6_internal_2_l_5,n_429_or_0_3_l_5,n12_3_l_5,n_431_3_l_5,G78_3_l_5,n_576_3_l_5,n11_3_l_5,n_102_3_l_5,n_547_3_l_5,n13_3_l_5,n14_3_l_5,n15_3_l_5,n16_3_l_5,N1_1_r_5,n3_1_r_5,P6_internal_2_r_5,n12_3_r_5,n_431_3_r_5,n11_3_r_5,n13_3_r_5,n14_3_r_5,n15_3_r_5,n16_3_r_5,N3_5_r_5,n3_5_r_5;
DFFARX1 I_0(P6_2_l_2,blif_clk_net_1_r_5,n1_1_r_5,ACVQN2_0_r_2,);
and I_1(n_266_and_0_0_r_2,n_102_3_l_2,ACVQN1_0_r_2);
DFFARX1 I_2(N1_1_r_2,blif_clk_net_1_r_5,n1_1_r_5,G199_1_r_2,);
DFFARX1 I_3(n_547_3_l_2,blif_clk_net_1_r_5,n1_1_r_5,G214_1_r_2,);
nand I_4(n_429_or_0_3_r_2,ACVQN1_2_l_2,n12_3_r_2);
DFFARX1 I_5(n_431_3_r_2,blif_clk_net_1_r_5,n1_1_r_5,G78_3_r_2,);
nand I_6(n_576_3_r_2,ACVQN1_2_l_2,n11_3_r_2);
not I_7(n_102_3_r_2,G78_3_l_2);
nand I_8(n_547_3_r_2,n_102_3_l_2,n13_3_r_2);
nor I_9(n_42_5_r_2,ACVQN1_2_l_2,P6_2_l_2);
DFFARX1 I_10(N3_5_r_2,blif_clk_net_1_r_5,n1_1_r_5,G199_5_r_2,);
DFFARX1 I_11(IN_2_2_l_2,blif_clk_net_1_r_5,n1_1_r_5,ACVQN1_2_l_2,);
not I_12(P6_2_l_2,P6_internal_2_l_2);
DFFARX1 I_13(IN_1_2_l_2,blif_clk_net_1_r_5,n1_1_r_5,P6_internal_2_l_2,);
nand I_14(n_429_or_0_3_l_2,G1_3_l_2,n12_3_l_2);
not I_15(n12_3_l_2,IN_5_3_l_2);
or I_16(n_431_3_l_2,IN_8_3_l_2,n14_3_l_2);
DFFARX1 I_17(n_431_3_l_2,blif_clk_net_1_r_5,n1_1_r_5,G78_3_l_2,);
nand I_18(n_576_3_l_2,IN_7_3_l_2,n11_3_l_2);
nor I_19(n11_3_l_2,G2_3_l_2,n12_3_l_2);
not I_20(n_102_3_l_2,G2_3_l_2);
nand I_21(n_547_3_l_2,IN_11_3_l_2,n13_3_l_2);
nor I_22(n13_3_l_2,G2_3_l_2,IN_10_3_l_2);
and I_23(n14_3_l_2,IN_2_3_l_2,n15_3_l_2);
nor I_24(n15_3_l_2,IN_4_3_l_2,n16_3_l_2);
not I_25(n16_3_l_2,G1_3_l_2);
DFFARX1 I_26(G78_3_l_2,blif_clk_net_1_r_5,n1_1_r_5,ACVQN1_0_r_2,);
and I_27(N1_1_r_2,G78_3_l_2,n3_1_r_2);
nand I_28(n3_1_r_2,n_576_3_l_2,n_547_3_l_2);
not I_29(n12_3_r_2,n_429_or_0_3_l_2);
or I_30(n_431_3_r_2,n_429_or_0_3_l_2,n14_3_r_2);
nor I_31(n11_3_r_2,G78_3_l_2,n12_3_r_2);
nor I_32(n13_3_r_2,G78_3_l_2,n_576_3_l_2);
and I_33(n14_3_r_2,n_576_3_l_2,n15_3_r_2);
nor I_34(n15_3_r_2,P6_2_l_2,n16_3_r_2);
not I_35(n16_3_r_2,ACVQN1_2_l_2);
and I_36(N3_5_r_2,n_102_3_l_2,n3_5_r_2);
nand I_37(n3_5_r_2,ACVQN1_2_l_2,n_429_or_0_3_l_2);
DFFARX1 I_38(N1_1_r_5,blif_clk_net_1_r_5,n1_1_r_5,G199_1_r_5,);
DFFARX1 I_39(ACVQN1_2_l_5,blif_clk_net_1_r_5,n1_1_r_5,G214_1_r_5,);
DFFARX1 I_40(n_429_or_0_3_l_5,blif_clk_net_1_r_5,n1_1_r_5,ACVQN1_2_r_5,);
not I_41(P6_2_r_5,P6_internal_2_r_5);
nand I_42(n_429_or_0_3_r_5,n_576_3_l_5,n12_3_r_5);
DFFARX1 I_43(n_431_3_r_5,blif_clk_net_1_r_5,n1_1_r_5,G78_3_r_5,);
nand I_44(n_576_3_r_5,P6_2_l_5,n11_3_r_5);
not I_45(n_102_3_r_5,ACVQN1_2_l_5);
nand I_46(n_547_3_r_5,G78_3_l_5,n13_3_r_5);
nor I_47(n_42_5_r_5,n_576_3_l_5,n_102_3_l_5);
DFFARX1 I_48(N3_5_r_5,blif_clk_net_1_r_5,n1_1_r_5,G199_5_r_5,);
not I_49(n1_1_r_5,blif_reset_net_1_r_5);
DFFARX1 I_50(G214_1_r_2,blif_clk_net_1_r_5,n1_1_r_5,ACVQN1_2_l_5,);
not I_51(P6_2_l_5,P6_internal_2_l_5);
DFFARX1 I_52(G199_5_r_2,blif_clk_net_1_r_5,n1_1_r_5,P6_internal_2_l_5,);
nand I_53(n_429_or_0_3_l_5,n12_3_l_5,n_576_3_r_2);
not I_54(n12_3_l_5,G78_3_r_2);
or I_55(n_431_3_l_5,n14_3_l_5,n_547_3_r_2);
DFFARX1 I_56(n_431_3_l_5,blif_clk_net_1_r_5,n1_1_r_5,G78_3_l_5,);
nand I_57(n_576_3_l_5,n11_3_l_5,n_266_and_0_0_r_2);
nor I_58(n11_3_l_5,n12_3_l_5,n_102_3_r_2);
not I_59(n_102_3_l_5,n_102_3_r_2);
nand I_60(n_547_3_l_5,n13_3_l_5,ACVQN2_0_r_2);
nor I_61(n13_3_l_5,n_102_3_r_2,n_42_5_r_2);
and I_62(n14_3_l_5,n15_3_l_5,G199_1_r_2);
nor I_63(n15_3_l_5,n16_3_l_5,n_429_or_0_3_r_2);
not I_64(n16_3_l_5,n_576_3_r_2);
and I_65(N1_1_r_5,n_102_3_l_5,n3_1_r_5);
nand I_66(n3_1_r_5,ACVQN1_2_l_5,n_547_3_l_5);
DFFARX1 I_67(G78_3_l_5,blif_clk_net_1_r_5,n1_1_r_5,P6_internal_2_r_5,);
not I_68(n12_3_r_5,n_102_3_l_5);
or I_69(n_431_3_r_5,P6_2_l_5,n14_3_r_5);
nor I_70(n11_3_r_5,ACVQN1_2_l_5,n12_3_r_5);
nor I_71(n13_3_r_5,ACVQN1_2_l_5,n_576_3_l_5);
and I_72(n14_3_r_5,n_429_or_0_3_l_5,n15_3_r_5);
nor I_73(n15_3_r_5,G78_3_l_5,n16_3_r_5);
not I_74(n16_3_r_5,n_576_3_l_5);
and I_75(N3_5_r_5,n_429_or_0_3_l_5,n3_5_r_5);
nand I_76(n3_5_r_5,P6_2_l_5,n_576_3_l_5);
endmodule


