module test_I6011(I1477,I1470,I6011);
input I1477,I1470;
output I6011;
wire I4917,I5994,I2143,I4544,I4506,I4512,I4521,I4869,I4674,I2149,I2155,I4742,I4807,I4824,I4790,I4773;
nor I_0(I4917,I4869,I4674);
nand I_1(I5994,I4512,I4506);
DFFARX1 I_2(I1470,,,I2143,);
not I_3(I4544,I1477);
and I_4(I6011,I5994,I4521);
nand I_5(I4506,I4869,I4773);
nand I_6(I4512,I4824,I4790);
DFFARX1 I_7(I4917,I1470,I4544,,,I4521,);
DFFARX1 I_8(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_9(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_10(I1470,,,I2149,);
DFFARX1 I_11(I1470,,,I2155,);
DFFARX1 I_12(I1470,I4544,,,I4742,);
DFFARX1 I_13(I1470,I4544,,,I4807,);
and I_14(I4824,I4807,I2143);
nor I_15(I4790,I4674,I4773);
not I_16(I4773,I4742);
endmodule


