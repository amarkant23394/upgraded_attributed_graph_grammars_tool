module test_I12605(I10633,I1477,I12814,I10618,I9477,I9465,I1470,I12605);
input I10633,I1477,I12814,I10618,I9477,I9465,I1470;
output I12605;
wire I10647,I11105,I12930,I12947,I12831,I12848,I10715,I13023,I10766,I10636,I10732,I12619,I12913,I10609;
not I_0(I10647,I1477);
and I_1(I11105,I10766);
and I_2(I12930,I12913,I10609);
nor I_3(I12947,I12930,I12848);
and I_4(I12831,I12814,I10618);
DFFARX1 I_5(I12831,I1470,I12619,,,I12848,);
nor I_6(I10715,I9477);
DFFARX1 I_7(I10636,I1470,I12619,,,I13023,);
not I_8(I10766,I9477);
nor I_9(I10636,I10732,I10766);
nand I_10(I10732,I10715,I9465);
not I_11(I12619,I1477);
DFFARX1 I_12(I10633,I1470,I12619,,,I12913,);
nand I_13(I12605,I13023,I12947);
DFFARX1 I_14(I11105,I1470,I10647,,,I10609,);
endmodule


