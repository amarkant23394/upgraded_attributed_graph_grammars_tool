module test_I13740(I1477,I1470,I11990,I13740);
input I1477,I1470,I11990;
output I13740;
wire I12270,I12239,I14162,I10014,I11938,I12208,I13775,I11973;
nand I_0(I12270,I11990,I10014);
DFFARX1 I_1(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_2(I11938,I1470,I13775,,,I14162,);
DFFARX1 I_3(I1470,,,I10014,);
and I_4(I11938,I12270,I12239);
DFFARX1 I_5(I1470,I11973,,,I12208,);
not I_6(I13775,I1477);
DFFARX1 I_7(I14162,I1470,I13775,,,I13740,);
not I_8(I11973,I1477);
endmodule


