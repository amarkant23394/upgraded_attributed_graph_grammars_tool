module test_I12930(I10879,I9477,I10698,I1477,I1470,I10732,I12930);
input I10879,I9477,I10698,I1477,I1470,I10732;
output I12930;
wire I12619,I10647,I11105,I12913,I10633,I10766,I10896,I11009,I11088,I11026,I10609;
not I_0(I12619,I1477);
not I_1(I10647,I1477);
and I_2(I11105,I10766,I11088);
DFFARX1 I_3(I10633,I1470,I12619,,,I12913,);
and I_4(I12930,I12913,I10609);
nand I_5(I10633,I10896,I11026);
not I_6(I10766,I9477);
DFFARX1 I_7(I10879,I1470,I10647,,,I10896,);
DFFARX1 I_8(I1470,I10647,,,I11009,);
nand I_9(I11088,I11009,I10698);
nor I_10(I11026,I11009,I10732);
DFFARX1 I_11(I11105,I1470,I10647,,,I10609,);
endmodule


