module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_5_r_7,n6_7,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_5_r_7,n6_7,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_5_r_7,n6_7,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_5_r_7,n6_7,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
nor I_43(N1371_0_r_7,n53_7,n52_7);
nor I_44(N1508_0_r_7,n51_7,n52_7);
nand I_45(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_46(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_47(n_576_5_r_7,n31_7,n32_7);
nor I_48(n_102_5_r_7,N1508_4_r_9,G78_5_r_9);
nand I_49(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_50(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_51(n_572_7_r_7,n54_7,n33_7);
nand I_52(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_53(n_549_7_r_7,n53_7,n36_7);
nand I_54(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_55(n_452_7_r_7,n_547_5_r_9,N6147_9_r_9);
nor I_56(n4_7_l_7,n_576_5_r_9,N6134_9_r_9);
not I_57(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_58(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_59(n30_7,n53_7);
and I_60(N3_8_l_7,n50_7,N1508_4_r_9);
DFFARX1 I_61(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_62(n_431_5_r_7,n40_7,n41_7);
nor I_63(n4_7_r_7,n54_7,n49_7);
and I_64(n31_7,n_102_5_r_7,n39_7);
not I_65(n32_7,n_576_5_r_9);
nor I_66(n33_7,n34_7,n_576_5_r_9);
and I_67(n34_7,n35_7,N1372_4_r_9);
not I_68(n35_7,G199_8_r_9);
nor I_69(n36_7,n37_7,n_576_5_r_9);
or I_70(n37_7,n54_7,N1508_4_r_9);
or I_71(n38_7,n_42_8_r_9,N1372_4_r_9);
nor I_72(n39_7,n_452_7_r_7,G78_5_r_9);
nand I_73(n40_7,n46_7,n47_7);
nand I_74(n41_7,n42_7,n43_7);
nor I_75(n42_7,n44_7,n45_7);
nor I_76(n43_7,n_42_8_r_9,N1372_4_r_9);
nor I_77(n44_7,G199_8_r_9,N6147_2_r_9);
nor I_78(n45_7,G78_5_r_9,n_576_5_r_9);
nand I_79(n46_7,n35_7,N1372_4_r_9);
not I_80(n47_7,n_576_5_r_9);
or I_81(n48_7,n_452_7_r_7,G78_5_r_9);
not I_82(n49_7,n_452_7_r_7);
nand I_83(n50_7,N6147_2_r_9,n_42_8_r_9);
and I_84(n51_7,n_452_7_r_7,n45_7);
not I_85(n52_7,n44_7);
endmodule


