module test_I10633(I1477,I10664,I10845,I9477,I9576,I1470,I10633);
input I1477,I10664,I10845,I9477,I9576,I1470;
output I10633;
wire I10879,I10647,I11009,I11026,I10715,I9638,I10862,I9816,I10896,I9453,I10732,I9491,I9468,I9462,I9465,I9864;
or I_0(I10879,I10862,I9462);
not I_1(I10647,I1477);
nand I_2(I10633,I10896,I11026);
DFFARX1 I_3(I9468,I1470,I10647,,,I11009,);
nor I_4(I11026,I11009,I10732);
nor I_5(I10715,I10664,I9477);
nor I_6(I9638,I9576);
and I_7(I10862,I10845,I9453);
DFFARX1 I_8(I1470,I9491,,,I9816,);
DFFARX1 I_9(I10879,I1470,I10647,,,I10896,);
nand I_10(I9453,I9816);
nand I_11(I10732,I10715,I9465);
not I_12(I9491,I1477);
DFFARX1 I_13(I9864,I1470,I9491,,,I9468,);
not I_14(I9462,I9576);
nand I_15(I9465,I9816,I9638);
nor I_16(I9864,I9816);
endmodule


