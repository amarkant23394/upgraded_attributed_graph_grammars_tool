module test_I6309(I2742,I4017,I1477,I1470,I6309);
input I2742,I4017,I1477,I1470;
output I6309;
wire I3975,I3966,I3954,I6442,I6329,I6493,I4068,I4308,I4034,I6459,I2724,I3983;
nor I_0(I3975,I4308,I4034);
or I_1(I3966,I4068,I4034);
not I_2(I3954,I4068);
nand I_3(I6309,I6493,I6459);
nor I_4(I6442,I3975,I3954);
not I_5(I6329,I1477);
DFFARX1 I_6(I3966,I1470,I6329,,,I6493,);
nor I_7(I4068,I2742,I2724);
DFFARX1 I_8(I1470,I3983,,,I4308,);
DFFARX1 I_9(I4017,I1470,I3983,,,I4034,);
not I_10(I6459,I6442);
DFFARX1 I_11(I1470,,,I2724,);
not I_12(I3983,I1477);
endmodule


