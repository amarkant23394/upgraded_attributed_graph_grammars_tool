module test_I11184(I1477,I9771,I8193,I9576,I1470,I11184);
input I1477,I9771,I8193,I9576,I1470;
output I11184;
wire I10647,I10664,I9474,I9471,I10715,I9542,I9638,I11167,I9816,I11150,I10732,I9491,I9477,I9833,I9465,I9621;
not I_0(I10647,I1477);
not I_1(I10664,I9471);
or I_2(I9474,I9576,I9542);
nor I_3(I9471,I9542);
nor I_4(I10715,I10664,I9477);
DFFARX1 I_5(I1470,I9491,,,I9542,);
nor I_6(I9638,I9621,I9576);
nand I_7(I11184,I11167,I10732);
not I_8(I11167,I11150);
DFFARX1 I_9(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_10(I9474,I1470,I10647,,,I11150,);
nand I_11(I10732,I10715,I9465);
not I_12(I9491,I1477);
nor I_13(I9477,I9771,I9833);
and I_14(I9833,I9816);
nand I_15(I9465,I9816,I9638);
DFFARX1 I_16(I1470,I9491,,,I9621,);
endmodule


