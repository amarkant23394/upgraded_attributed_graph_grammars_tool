module test_I10715(I9491,I8216,I8753,I1470,I9525,I8193,I9672,I10715);
input I9491,I8216,I8753,I1470,I9525,I8193,I9672;
output I10715;
wire I9477,I8187,I9542,I10664,I9754,I9816,I9559,I9771,I8178,I9833,I9689,I9471;
nor I_0(I9477,I9771,I9833);
nor I_1(I10715,I10664,I9477);
DFFARX1 I_2(I1470,I8216,,,I8187,);
DFFARX1 I_3(I9525,I1470,I9491,,,I9542,);
not I_4(I10664,I9471);
DFFARX1 I_5(I8187,I1470,I9491,,,I9754,);
DFFARX1 I_6(I8193,I1470,I9491,,,I9816,);
not I_7(I9559,I9542);
and I_8(I9771,I9754,I8178);
DFFARX1 I_9(I8753,I1470,I8216,,,I8178,);
and I_10(I9833,I9816,I9559);
DFFARX1 I_11(I9672,I1470,I9491,,,I9689,);
nor I_12(I9471,I9689,I9542);
endmodule


