module test_I6705(I1477,I2745,I3217,I1470,I6705);
input I1477,I2745,I3217,I1470;
output I6705;
wire I2733,I3107,I3076,I4435,I3972,I3983,I2742,I3155,I6329,I4068,I4263,I2724,I6688,I2963,I4452,I2759,I3948,I4246;
nand I_0(I2733,I3217,I3107);
nor I_1(I3107,I3076);
DFFARX1 I_2(I1470,I2759,,,I3076,);
and I_3(I6705,I6688,I3972);
and I_4(I4435,I4068);
or I_5(I3972,I4263,I4068);
not I_6(I3983,I1477);
or I_7(I2742,I3076,I2963);
or I_8(I3155,I3076);
not I_9(I6329,I1477);
nor I_10(I4068,I2742,I2724);
and I_11(I4263,I4246,I2733);
DFFARX1 I_12(I3155,I1470,I2759,,,I2724,);
DFFARX1 I_13(I3948,I1470,I6329,,,I6688,);
DFFARX1 I_14(I1470,I2759,,,I2963,);
or I_15(I4452,I4263,I4435);
not I_16(I2759,I1477);
DFFARX1 I_17(I4452,I1470,I3983,,,I3948,);
DFFARX1 I_18(I2745,I1470,I3983,,,I4246,);
endmodule


