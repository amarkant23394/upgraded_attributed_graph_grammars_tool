module test_I11057(I1477,I9771,I1470,I11057);
input I1477,I9771,I1470;
output I11057;
wire I9477,I10647,I9833,I9491,I10797,I9816,I10766,I9468,I11009,I9621,I9864;
nor I_0(I9477,I9771,I9833);
not I_1(I10647,I1477);
and I_2(I9833,I9816);
not I_3(I9491,I1477);
not I_4(I10797,I10766);
nor I_5(I11057,I11009,I10797);
DFFARX1 I_6(I1470,I9491,,,I9816,);
not I_7(I10766,I9477);
DFFARX1 I_8(I9864,I1470,I9491,,,I9468,);
DFFARX1 I_9(I9468,I1470,I10647,,,I11009,);
DFFARX1 I_10(I1470,I9491,,,I9621,);
nor I_11(I9864,I9816,I9621);
endmodule


