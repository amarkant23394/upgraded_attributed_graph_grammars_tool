module test_I8736(I4629,I1477,I1470,I8736);
input I4629,I1477,I1470;
output I8736;
wire I8216,I5864,I5751,I4595,I4536,I4515,I4527,I5881,I5915,I5731;
not I_0(I8216,I1477);
nor I_1(I5864,I4536,I4515);
not I_2(I5751,I1477);
DFFARX1 I_3(I1470,,,I4595,);
nor I_4(I4536,I4595);
not I_5(I4515,I4629);
or I_6(I4527,I4629,I4595);
not I_7(I5881,I5864);
DFFARX1 I_8(I4527,I1470,I5751,,,I5915,);
nand I_9(I5731,I5915,I5881);
DFFARX1 I_10(I5731,I1470,I8216,,,I8736,);
endmodule


