module test_I4578(I1477,I1231,I1303,I1375,I1287,I2441,I1470,I4578);
input I1477,I1231,I1303,I1375,I1287,I2441,I1470;
output I4578;
wire I2311,I2540,I4561,I2458,I2152,I2345,I2161,I2173,I2181,I2509,I2557,I2294,I2232;
not I_0(I2311,I2294);
DFFARX1 I_1(I1470,I2181,,,I2540,);
nand I_2(I4561,I2152,I2173);
DFFARX1 I_3(I2441,I1470,I2181,,,I2458,);
DFFARX1 I_4(I2458,I1470,I2181,,,I2152,);
and I_5(I4578,I4561,I2161);
DFFARX1 I_6(I1375,I1470,I2181,,,I2345,);
nand I_7(I2161,I2345,I2311);
nand I_8(I2173,I2557,I2509);
not I_9(I2181,I1477);
nor I_10(I2509,I2458,I2232);
and I_11(I2557,I2540,I1303);
nor I_12(I2294,I1287,I1231);
DFFARX1 I_13(I1470,I2181,,,I2232,);
endmodule


