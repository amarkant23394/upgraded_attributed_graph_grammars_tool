module test_I17384(I15582,I17628,I1477,I1470,I17384);
input I15582,I17628,I1477,I1470;
output I17384;
wire I17413,I17645,I17696,I17662;
not I_0(I17413,I1477);
or I_1(I17645,I17628,I15582);
DFFARX1 I_2(I17662,I1470,I17413,,,I17696,);
DFFARX1 I_3(I17645,I1470,I17413,,,I17662,);
not I_4(I17384,I17696);
endmodule


