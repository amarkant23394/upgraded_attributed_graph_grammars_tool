module test_c6288_7_355(IN_1,IN_2,IN_3,IN_4,IN_5,N6150,N6147,N6134);
input IN_1,IN_2,IN_3,IN_4,IN_5;
output N6150,N6147,N6134;
wire N6145,N6141,N6146,N6124;
nor I_0(N6145,N6141,IN_1);
nor I_1(N6150,N6145,N6146);
not I_2(N6141,IN_2);
not I_3(N6146,N6141);
nor I_4(N6147,N6141,N6124);
nor I_5(N6124,IN_3,IN_4);
nor I_6(N6134,N6124,IN_5);
endmodule


