module test_I6329(I1477,I6329);
input I1477;
output I6329;
wire ;
not I_0(I6329,I1477);
endmodule


