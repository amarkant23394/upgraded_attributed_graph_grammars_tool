module test_I6300(I3951,I3945,I1477,I1470,I4356,I6300);
input I3951,I3945,I1477,I1470,I4356;
output I6300;
wire I6606,I3960,I6589,I6329,I6572,I3983;
DFFARX1 I_0(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_1(I4356,I1470,I3983,,,I3960,);
and I_2(I6589,I6572,I3960);
not I_3(I6329,I1477);
nand I_4(I6572,I3951,I3945);
DFFARX1 I_5(I6606,I1470,I6329,,,I6300,);
not I_6(I3983,I1477);
endmodule


