module test_final(G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7,n_431_0_l_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_7,blif_clk_net_1_r_8,n8_8,G42_1_r_7,);
nor I_1(n_572_1_r_7,n30_7,n31_7);
nand I_2(n_573_1_r_7,IN_7_0_l_7,n28_7);
nor I_3(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_4(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_5(N1_4_r_7,blif_clk_net_1_r_8,n8_8,G199_4_r_7,);
DFFARX1 I_6(n26_7,blif_clk_net_1_r_8,n8_8,G214_4_r_7,);
DFFARX1 I_7(n5_7,blif_clk_net_1_r_8,n8_8,ACVQN1_5_r_7,);
not I_8(P6_5_r_7,P6_5_r_internal_7);
or I_9(n_431_0_l_7,IN_8_0_l_7,n36_7);
DFFARX1 I_10(n_431_0_l_7,blif_clk_net_1_r_8,n8_8,n43_7,);
not I_11(n27_7,n43_7);
DFFARX1 I_12(IN_2_5_l_7,blif_clk_net_1_r_8,n8_8,ACVQN1_5_l_7,);
DFFARX1 I_13(IN_1_5_l_7,blif_clk_net_1_r_8,n8_8,n44_7,);
nor I_14(n4_1_r_7,n30_7,n38_7);
nor I_15(N1_4_r_7,n27_7,n40_7);
nand I_16(n26_7,IN_11_0_l_7,n39_7);
not I_17(n5_7,G2_0_l_7);
DFFARX1 I_18(ACVQN1_5_l_7,blif_clk_net_1_r_8,n8_8,P6_5_r_internal_7,);
nor I_19(n28_7,n26_7,n29_7);
not I_20(n29_7,IN_5_0_l_7);
not I_21(n30_7,G1_0_l_7);
nand I_22(n31_7,n27_7,n29_7);
nor I_23(n32_7,ACVQN1_5_l_7,n34_7);
nor I_24(n33_7,G2_0_l_7,n29_7);
not I_25(n34_7,IN_7_0_l_7);
nor I_26(n35_7,n43_7,n44_7);
and I_27(n36_7,IN_2_0_l_7,n37_7);
nor I_28(n37_7,IN_4_0_l_7,n30_7);
nand I_29(n38_7,G2_0_l_7,n29_7);
nor I_30(n39_7,G2_0_l_7,IN_10_0_l_7);
nor I_31(n40_7,n44_7,n41_7);
nor I_32(n41_7,n34_7,n42_7);
nand I_33(n42_7,IN_5_0_l_7,n5_7);
DFFARX1 I_34(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_35(n_572_1_r_8,n39_8,n23_8);
and I_36(n_549_1_r_8,n38_8,n23_8);
nand I_37(n_569_1_r_8,n38_8,n24_8);
nor I_38(n_452_1_r_8,n25_8,n26_8);
nor I_39(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_40(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_41(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_42(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_43(n_431_0_l_8,n29_8,P6_5_r_7);
not I_44(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_45(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_46(n19_8,G78_0_l_8);
DFFARX1 I_47(n_572_1_r_7,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_48(n22_8,n39_8);
DFFARX1 I_49(G199_4_r_7,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_50(n4_1_r_8,G78_0_l_8,n33_8);
nor I_51(N3_2_r_8,n22_8,n35_8);
nor I_52(N1_4_r_8,n27_8,n37_8);
nand I_53(n23_8,n32_8,G42_1_r_7);
not I_54(n24_8,n23_8);
nand I_55(n25_8,n36_8,n_569_1_r_7);
nand I_56(n26_8,n27_8,n28_8);
nor I_57(n27_8,n31_8,n_549_1_r_7);
not I_58(n28_8,G214_4_r_7);
and I_59(n29_8,n30_8,G42_1_r_7);
nor I_60(n30_8,n31_8,n_572_1_r_7);
not I_61(n31_8,n_573_1_r_7);
and I_62(n32_8,n28_8,n_549_1_r_7);
nand I_63(n33_8,n28_8,n34_8);
not I_64(n34_8,n25_8);
nor I_65(n35_8,n34_8,G214_4_r_7);
not I_66(n36_8,ACVQN1_5_r_7);
nor I_67(n37_8,n19_8,n38_8);
endmodule


