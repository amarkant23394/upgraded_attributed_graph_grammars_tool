module test_I5249(I1518,I3388,I1504,I3487,I1489,I2103,I1470,I3538,I5249);
input I1518,I3388,I1504,I3487,I1489,I2103,I1470,I3538;
output I5249;
wire I3846,I3504,I3521,I3380,I1495,I3555,I3747;
nor I_0(I3846,I3747,I3555);
and I_1(I3504,I3487,I1489);
nor I_2(I3521,I3504,I1495);
nand I_3(I3380,I3521,I3846);
DFFARX1 I_4(I2103,I1470,I1518,,,I1495,);
DFFARX1 I_5(I3538,I1470,I3388,,,I3555,);
not I_6(I5249,I3380);
DFFARX1 I_7(I1504,I1470,I3388,,,I3747,);
endmodule


