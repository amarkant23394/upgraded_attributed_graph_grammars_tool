module test_I6442(I1477,I2810,I1470,I6442);
input I1477,I2810,I1470;
output I6442;
wire I3076,I3983,I2742,I3954,I3155,I4068,I2724,I3975,I4000,I2963,I4308,I4034,I2730,I2759,I4017,I3124,I2727;
nor I_0(I6442,I3975,I3954);
DFFARX1 I_1(I1470,I2759,,,I3076,);
not I_2(I3983,I1477);
or I_3(I2742,I3076,I2963);
not I_4(I3954,I4068);
or I_5(I3155,I3076);
nor I_6(I4068,I2742,I2724);
DFFARX1 I_7(I3155,I1470,I2759,,,I2724,);
nor I_8(I3975,I4308,I4034);
nand I_9(I4000,I2724);
DFFARX1 I_10(I1470,I2759,,,I2963,);
DFFARX1 I_11(I2727,I1470,I3983,,,I4308,);
DFFARX1 I_12(I4017,I1470,I3983,,,I4034,);
not I_13(I2730,I3076);
not I_14(I2759,I1477);
and I_15(I4017,I4000,I2730);
nor I_16(I3124,I3076);
nand I_17(I2727,I2810,I3124);
endmodule


