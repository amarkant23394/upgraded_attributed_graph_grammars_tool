module test_I7427(I1477,I1470,I7427);
input I1477,I1470;
output I7427;
wire I5594,I6907,I7410,I5512,I5082,I5105;
DFFARX1 I_0(I5512,I1470,I5105,,,I5594,);
not I_1(I7427,I7410);
not I_2(I6907,I1477);
DFFARX1 I_3(I5082,I1470,I6907,,,I7410,);
DFFARX1 I_4(I1470,I5105,,,I5512,);
not I_5(I5082,I5594);
not I_6(I5105,I1477);
endmodule


