module test_final(G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11,n_431_0_l_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_11,blif_clk_net_1_r_9,n5_9,G42_1_r_11,);
nor I_1(n_572_1_r_11,n29_11,n30_11);
nand I_2(n_573_1_r_11,n26_11,n28_11);
nor I_3(n_549_1_r_11,n27_11,n32_11);
nand I_4(n_569_1_r_11,n45_11,n28_11);
nor I_5(n_452_1_r_11,n43_11,n44_11);
nor I_6(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_7(N3_2_r_11,blif_clk_net_1_r_9,n5_9,G199_2_r_11,);
DFFARX1 I_8(n24_11,blif_clk_net_1_r_9,n5_9,ACVQN2_3_r_11,);
nor I_9(n_266_and_0_3_r_11,n20_11,n37_11);
or I_10(n_431_0_l_11,IN_8_0_l_11,n33_11);
DFFARX1 I_11(n_431_0_l_11,blif_clk_net_1_r_9,n5_9,n43_11,);
not I_12(n26_11,n43_11);
DFFARX1 I_13(IN_2_5_l_11,blif_clk_net_1_r_9,n5_9,n44_11,);
DFFARX1 I_14(IN_1_5_l_11,blif_clk_net_1_r_9,n5_9,n45_11,);
not I_15(n27_11,n45_11);
nor I_16(n4_1_r_11,n44_11,n25_11);
nor I_17(N3_2_r_11,n45_11,n40_11);
nand I_18(n24_11,IN_11_0_l_11,n39_11);
nand I_19(n25_11,IN_7_0_l_11,n38_11);
DFFARX1 I_20(n25_11,blif_clk_net_1_r_9,n5_9,n20_internal_11,);
not I_21(n20_11,n20_internal_11);
not I_22(n28_11,n25_11);
not I_23(n29_11,G1_0_l_11);
nand I_24(n30_11,n26_11,n31_11);
not I_25(n31_11,IN_5_0_l_11);
and I_26(n32_11,n26_11,n44_11);
and I_27(n33_11,IN_2_0_l_11,n34_11);
nor I_28(n34_11,IN_4_0_l_11,n29_11);
not I_29(n35_11,G2_0_l_11);
nand I_30(n36_11,G1_0_l_11,n31_11);
nor I_31(n37_11,IN_5_0_l_11,n29_11);
nor I_32(n38_11,G2_0_l_11,n31_11);
nor I_33(n39_11,G2_0_l_11,IN_10_0_l_11);
nor I_34(n40_11,G2_0_l_11,n41_11);
nor I_35(n41_11,IN_10_0_l_11,n42_11);
not I_36(n42_11,IN_11_0_l_11);
DFFARX1 I_37(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_38(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_39(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_40(n_549_1_r_9,n17_9,n18_9);
or I_41(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_42(n_452_1_r_9,n26_9,n25_9);
nor I_43(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_44(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_45(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_46(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_47(N3_2_l_9,n22_9,G199_2_r_11);
not I_48(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_49(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_50(n16_9,n27_9);
DFFARX1 I_51(G42_1_r_11,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_52(n15_9,n26_9);
DFFARX1 I_53(n_572_1_r_11,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_54(n29_9,n29_internal_9);
and I_55(N1_4_l_9,n24_9,n_266_and_0_3_r_11);
DFFARX1 I_56(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_57(ACVQN2_3_r_11,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_58(n28_9,n28_internal_9);
nor I_59(n4_1_r_9,n27_9,n26_9);
nor I_60(N3_2_r_9,n15_9,n21_9);
nor I_61(N1_4_r_9,n16_9,n21_9);
nor I_62(n_42_2_l_9,n_573_1_r_11,n_549_1_r_11);
not I_63(n17_9,n_452_1_r_9);
nand I_64(n18_9,n27_9,n15_9);
nor I_65(n19_9,n29_9,n20_9);
not I_66(n20_9,n_569_1_r_11);
and I_67(n21_9,n23_9,n_569_1_r_11);
nand I_68(n22_9,n_549_1_r_11,n_42_2_r_11);
nor I_69(n23_9,n29_9,n28_9);
nand I_70(n24_9,G42_1_r_11,n_452_1_r_11);
endmodule


