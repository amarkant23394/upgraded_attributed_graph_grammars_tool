module test_I6878(I7122,I5085,I1477,I1470,I6878);
input I7122,I5085,I1477,I1470;
output I6878;
wire I7190,I7156,I6907,I7139;
DFFARX1 I_0(I7156,I1470,I6907,,,I7190,);
DFFARX1 I_1(I7139,I1470,I6907,,,I7156,);
not I_2(I6907,I1477);
or I_3(I7139,I7122,I5085);
not I_4(I6878,I7190);
endmodule


