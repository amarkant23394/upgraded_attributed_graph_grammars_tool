module test_I4807(I1477,I1470,I2198,I1271,I4807);
input I1477,I1470,I2198,I1271;
output I4807;
wire I2181,I4544,I2170,I2232,I2215;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
not I_2(I2170,I2232);
DFFARX1 I_3(I2215,I1470,I2181,,,I2232,);
DFFARX1 I_4(I2170,I1470,I4544,,,I4807,);
and I_5(I2215,I2198,I1271);
endmodule


