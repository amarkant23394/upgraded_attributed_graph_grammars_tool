module test_I2492(I1231,I1327,I1477,I1470,I2424,I1375,I1287,I2492);
input I1231,I1327,I1477,I1470,I2424,I1375,I1287;
output I2492;
wire I2362,I2441,I2475,I2181,I2294,I2458,I2345;
and I_0(I2492,I2294,I2475);
not I_1(I2362,I2345);
and I_2(I2441,I2424,I1327);
nor I_3(I2475,I2458,I2362);
not I_4(I2181,I1477);
nor I_5(I2294,I1287,I1231);
DFFARX1 I_6(I2441,I1470,I2181,,,I2458,);
DFFARX1 I_7(I1375,I1470,I2181,,,I2345,);
endmodule


