module test_I8124(I7652,I1477,I1470,I6459,I6318,I6705,I6657,I8124);
input I7652,I1477,I1470,I6459,I6318,I6705,I6657;
output I8124;
wire I8107,I6321,I8090,I8011,I7570,I6309,I6493,I8028,I7994,I7977,I7669;
not I_0(I8107,I8090);
nand I_1(I6321,I6705,I6657);
DFFARX1 I_2(I6309,I1470,I7570,,,I8090,);
nor I_3(I8011,I7669,I7994);
not I_4(I7570,I1477);
nand I_5(I6309,I6493,I6459);
DFFARX1 I_6(I1470,,,I6493,);
and I_7(I8028,I7977,I8011);
not I_8(I7994,I7977);
or I_9(I8124,I8107,I8028);
DFFARX1 I_10(I6321,I1470,I7570,,,I7977,);
nand I_11(I7669,I7652,I6318);
endmodule


