module test_I11361(I9320,I9032,I1477,I8913,I6992,I7026,I8947,I1470,I8879,I11361);
input I9320,I9032,I1477,I8913,I6992,I7026,I8947,I1470,I8879;
output I11361;
wire I8845,I9179,I8839,I11344,I9337,I9396,I9049,I8862,I6881,I8848,I9083,I9413,I6896,I9066,I6869;
or I_0(I8845,I9179,I9066);
DFFARX1 I_1(I6896,I1470,I8862,,,I9179,);
DFFARX1 I_2(I9337,I1470,I8862,,,I8839,);
nor I_3(I11344,I8848,I8839);
nor I_4(I9337,I9320,I8913);
not I_5(I9396,I9320);
or I_6(I9049,I9032,I6869);
not I_7(I8862,I1477);
nand I_8(I6881,I6992);
nor I_9(I8848,I9083,I9413);
nand I_10(I9083,I8879,I6881);
and I_11(I9413,I8947,I9396);
nor I_12(I6896,I6992,I7026);
nand I_13(I11361,I11344,I8845);
DFFARX1 I_14(I9049,I1470,I8862,,,I9066,);
DFFARX1 I_15(I1470,,,I6869,);
endmodule


