module test_final(IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_reset_net_0_r_1,blif_clk_net_0_r_1,ACVQN2_0_r_1,n_266_and_0_0_r_1,G199_1_r_1,G214_1_r_1,ACVQN1_2_r_1,P6_2_r_1,n_429_or_0_3_r_1,G78_3_r_1,n_576_3_r_1,n_102_3_r_1,n_547_3_r_1);
input IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_reset_net_0_r_1,blif_clk_net_0_r_1;
output ACVQN2_0_r_1,n_266_and_0_0_r_1,G199_1_r_1,G214_1_r_1,ACVQN1_2_r_1,P6_2_r_1,n_429_or_0_3_r_1,G78_3_r_1,n_576_3_r_1,n_102_3_r_1,n_547_3_r_1;
wire ACVQN2_0_r_8,n_266_and_0_0_r_8,ACVQN1_2_r_8,P6_2_r_8,n_429_or_0_3_r_8,G78_3_r_8,n_576_3_r_8,n_102_3_r_8,n_547_3_r_8,n_42_5_r_8,G199_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8,ACVQN1_0_l_8,N1_1_l_8,G199_1_l_8,G214_1_l_8,n3_1_l_8,n_42_5_l_8,N3_5_l_8,G199_5_l_8,n3_5_l_8,ACVQN1_0_r_8,P6_internal_2_r_8,n12_3_r_8,n_431_3_r_8,n11_3_r_8,n13_3_r_8,n14_3_r_8,n15_3_r_8,n16_3_r_8,N3_5_r_8,n3_5_r_8,n1_0_r_1,ACVQN1_2_l_1,P6_2_l_1,P6_internal_2_l_1,n_429_or_0_3_l_1,n12_3_l_1,n_431_3_l_1,G78_3_l_1,n_576_3_l_1,n11_3_l_1,n_102_3_l_1,n_547_3_l_1,n13_3_l_1,n14_3_l_1,n15_3_l_1,n16_3_l_1,ACVQN1_0_r_1,N1_1_r_1,n3_1_r_1,P6_internal_2_r_1,n12_3_r_1,n_431_3_r_1,n11_3_r_1,n13_3_r_1,n14_3_r_1,n15_3_r_1,n16_3_r_1;
DFFARX1 I_0(n_266_and_0_0_l_8,blif_clk_net_0_r_1,n1_0_r_1,ACVQN2_0_r_8,);
and I_1(n_266_and_0_0_r_8,G199_5_l_8,ACVQN1_0_r_8);
DFFARX1 I_2(G199_5_l_8,blif_clk_net_0_r_1,n1_0_r_1,ACVQN1_2_r_8,);
not I_3(P6_2_r_8,P6_internal_2_r_8);
nand I_4(n_429_or_0_3_r_8,G199_5_l_8,n12_3_r_8);
DFFARX1 I_5(n_431_3_r_8,blif_clk_net_0_r_1,n1_0_r_1,G78_3_r_8,);
nand I_6(n_576_3_r_8,n_42_5_l_8,n11_3_r_8);
not I_7(n_102_3_r_8,n_266_and_0_0_l_8);
nand I_8(n_547_3_r_8,ACVQN2_0_l_8,n13_3_r_8);
nor I_9(n_42_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8);
DFFARX1 I_10(N3_5_r_8,blif_clk_net_0_r_1,n1_0_r_1,G199_5_r_8,);
DFFARX1 I_11(IN_1_0_l_8,blif_clk_net_0_r_1,n1_0_r_1,ACVQN2_0_l_8,);
and I_12(n_266_and_0_0_l_8,IN_4_0_l_8,ACVQN1_0_l_8);
DFFARX1 I_13(IN_2_0_l_8,blif_clk_net_0_r_1,n1_0_r_1,ACVQN1_0_l_8,);
and I_14(N1_1_l_8,IN_6_1_l_8,n3_1_l_8);
DFFARX1 I_15(N1_1_l_8,blif_clk_net_0_r_1,n1_0_r_1,G199_1_l_8,);
DFFARX1 I_16(IN_3_1_l_8,blif_clk_net_0_r_1,n1_0_r_1,G214_1_l_8,);
nand I_17(n3_1_l_8,IN_1_1_l_8,IN_2_1_l_8);
nor I_18(n_42_5_l_8,IN_1_5_l_8,IN_3_5_l_8);
and I_19(N3_5_l_8,IN_6_5_l_8,n3_5_l_8);
DFFARX1 I_20(N3_5_l_8,blif_clk_net_0_r_1,n1_0_r_1,G199_5_l_8,);
nand I_21(n3_5_l_8,IN_2_5_l_8,IN_3_5_l_8);
DFFARX1 I_22(G214_1_l_8,blif_clk_net_0_r_1,n1_0_r_1,ACVQN1_0_r_8,);
DFFARX1 I_23(G214_1_l_8,blif_clk_net_0_r_1,n1_0_r_1,P6_internal_2_r_8,);
not I_24(n12_3_r_8,G199_1_l_8);
or I_25(n_431_3_r_8,n_42_5_l_8,n14_3_r_8);
nor I_26(n11_3_r_8,n_266_and_0_0_l_8,n12_3_r_8);
nor I_27(n13_3_r_8,n_266_and_0_0_l_8,G199_1_l_8);
and I_28(n14_3_r_8,ACVQN2_0_l_8,n15_3_r_8);
nor I_29(n15_3_r_8,G199_1_l_8,n16_3_r_8);
not I_30(n16_3_r_8,G199_5_l_8);
and I_31(N3_5_r_8,n_42_5_l_8,n3_5_r_8);
nand I_32(n3_5_r_8,ACVQN2_0_l_8,G214_1_l_8);
DFFARX1 I_33(P6_2_l_1,blif_clk_net_0_r_1,n1_0_r_1,ACVQN2_0_r_1,);
and I_34(n_266_and_0_0_r_1,n_102_3_l_1,ACVQN1_0_r_1);
DFFARX1 I_35(N1_1_r_1,blif_clk_net_0_r_1,n1_0_r_1,G199_1_r_1,);
DFFARX1 I_36(n_576_3_l_1,blif_clk_net_0_r_1,n1_0_r_1,G214_1_r_1,);
DFFARX1 I_37(n_547_3_l_1,blif_clk_net_0_r_1,n1_0_r_1,ACVQN1_2_r_1,);
not I_38(P6_2_r_1,P6_internal_2_r_1);
nand I_39(n_429_or_0_3_r_1,ACVQN1_2_l_1,n12_3_r_1);
DFFARX1 I_40(n_431_3_r_1,blif_clk_net_0_r_1,n1_0_r_1,G78_3_r_1,);
nand I_41(n_576_3_r_1,n_547_3_l_1,n11_3_r_1);
not I_42(n_102_3_r_1,n_576_3_l_1);
nand I_43(n_547_3_r_1,P6_2_l_1,n13_3_r_1);
not I_44(n1_0_r_1,blif_reset_net_0_r_1);
DFFARX1 I_45(n_102_3_r_8,blif_clk_net_0_r_1,n1_0_r_1,ACVQN1_2_l_1,);
not I_46(P6_2_l_1,P6_internal_2_l_1);
DFFARX1 I_47(n_547_3_r_8,blif_clk_net_0_r_1,n1_0_r_1,P6_internal_2_l_1,);
nand I_48(n_429_or_0_3_l_1,n12_3_l_1,n_576_3_r_8);
not I_49(n12_3_l_1,G78_3_r_8);
or I_50(n_431_3_l_1,n14_3_l_1,n_42_5_r_8);
DFFARX1 I_51(n_431_3_l_1,blif_clk_net_0_r_1,n1_0_r_1,G78_3_l_1,);
nand I_52(n_576_3_l_1,n11_3_l_1,ACVQN1_2_r_8);
nor I_53(n11_3_l_1,n12_3_l_1,n_266_and_0_0_r_8);
not I_54(n_102_3_l_1,n_266_and_0_0_r_8);
nand I_55(n_547_3_l_1,n13_3_l_1,ACVQN2_0_r_8);
nor I_56(n13_3_l_1,n_266_and_0_0_r_8,P6_2_r_8);
and I_57(n14_3_l_1,n15_3_l_1,n_429_or_0_3_r_8);
nor I_58(n15_3_l_1,n16_3_l_1,G199_5_r_8);
not I_59(n16_3_l_1,n_576_3_r_8);
DFFARX1 I_60(n_429_or_0_3_l_1,blif_clk_net_0_r_1,n1_0_r_1,ACVQN1_0_r_1,);
and I_61(N1_1_r_1,n_429_or_0_3_l_1,n3_1_r_1);
nand I_62(n3_1_r_1,n_429_or_0_3_l_1,G78_3_l_1);
DFFARX1 I_63(ACVQN1_2_l_1,blif_clk_net_0_r_1,n1_0_r_1,P6_internal_2_r_1,);
not I_64(n12_3_r_1,n_102_3_l_1);
or I_65(n_431_3_r_1,P6_2_l_1,n14_3_r_1);
nor I_66(n11_3_r_1,G78_3_l_1,n12_3_r_1);
nor I_67(n13_3_r_1,G78_3_l_1,n_576_3_l_1);
and I_68(n14_3_r_1,ACVQN1_2_l_1,n15_3_r_1);
nor I_69(n15_3_r_1,n_576_3_l_1,n16_3_r_1);
not I_70(n16_3_r_1,ACVQN1_2_l_1);
endmodule


