module test_I2844(I1407,I1351,I1359,I2844);
input I1407,I1351,I1359;
output I2844;
wire I2776,I2827;
nand I_0(I2844,I2827,I1359);
not I_1(I2776,I1407);
nor I_2(I2827,I2776,I1351);
endmodule


