module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_3_r_10,blif_reset_net_3_r_10,n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10);
input IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_3_r_10,blif_reset_net_3_r_10;
output n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10;
wire ACVQN2_0_r_14,n_266_and_0_0_r_14,G199_1_r_14,G214_1_r_14,ACVQN1_2_r_14,P6_2_r_14,n_429_or_0_3_r_14,G78_3_r_14,n_576_3_r_14,n_102_3_r_14,n_547_3_r_14,ACVQN2_0_l_14,n_266_and_0_0_l_14,ACVQN1_0_l_14,N1_1_l_14,G199_1_l_14,G214_1_l_14,n3_1_l_14,n_42_5_l_14,N3_5_l_14,G199_5_l_14,n3_5_l_14,ACVQN1_0_r_14,N1_1_r_14,n3_1_r_14,P6_internal_2_r_14,n12_3_r_14,n_431_3_r_14,n11_3_r_14,n13_3_r_14,n14_3_r_14,n15_3_r_14,n16_3_r_14,n2_3_r_10,ACVQN2_0_l_10,n_266_and_0_0_l_10,ACVQN1_0_l_10,n4_4_l_10,G42_4_l_10,n_87_4_l_10,n_572_4_l_10,n_573_4_l_10,n_549_4_l_10,n7_4_l_10,n_569_4_l_10,n_452_4_l_10,n12_3_r_10,n_431_3_r_10,n11_3_r_10,n13_3_r_10,n14_3_r_10,n15_3_r_10,n16_3_r_10,n4_4_r_10,n_87_4_r_10,n7_4_r_10;
DFFARX1 I_0(n_266_and_0_0_l_14,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_r_14,);
and I_1(n_266_and_0_0_r_14,G199_5_l_14,ACVQN1_0_r_14);
DFFARX1 I_2(N1_1_r_14,blif_clk_net_3_r_10,n2_3_r_10,G199_1_r_14,);
DFFARX1 I_3(G199_1_l_14,blif_clk_net_3_r_10,n2_3_r_10,G214_1_r_14,);
DFFARX1 I_4(ACVQN2_0_l_14,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_2_r_14,);
not I_5(P6_2_r_14,P6_internal_2_r_14);
nand I_6(n_429_or_0_3_r_14,G214_1_l_14,n12_3_r_14);
DFFARX1 I_7(n_431_3_r_14,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_14,);
nand I_8(n_576_3_r_14,ACVQN2_0_l_14,n11_3_r_14);
not I_9(n_102_3_r_14,G199_5_l_14);
nand I_10(n_547_3_r_14,n_266_and_0_0_l_14,n13_3_r_14);
DFFARX1 I_11(IN_1_0_l_14,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_14,);
and I_12(n_266_and_0_0_l_14,IN_4_0_l_14,ACVQN1_0_l_14);
DFFARX1 I_13(IN_2_0_l_14,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_14,);
and I_14(N1_1_l_14,IN_6_1_l_14,n3_1_l_14);
DFFARX1 I_15(N1_1_l_14,blif_clk_net_3_r_10,n2_3_r_10,G199_1_l_14,);
DFFARX1 I_16(IN_3_1_l_14,blif_clk_net_3_r_10,n2_3_r_10,G214_1_l_14,);
nand I_17(n3_1_l_14,IN_1_1_l_14,IN_2_1_l_14);
nor I_18(n_42_5_l_14,IN_1_5_l_14,IN_3_5_l_14);
and I_19(N3_5_l_14,IN_6_5_l_14,n3_5_l_14);
DFFARX1 I_20(N3_5_l_14,blif_clk_net_3_r_10,n2_3_r_10,G199_5_l_14,);
nand I_21(n3_5_l_14,IN_2_5_l_14,IN_3_5_l_14);
DFFARX1 I_22(G214_1_l_14,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_r_14,);
and I_23(N1_1_r_14,G214_1_l_14,n3_1_r_14);
nand I_24(n3_1_r_14,ACVQN2_0_l_14,n_42_5_l_14);
DFFARX1 I_25(G199_5_l_14,blif_clk_net_3_r_10,n2_3_r_10,P6_internal_2_r_14,);
not I_26(n12_3_r_14,n_42_5_l_14);
or I_27(n_431_3_r_14,n_266_and_0_0_l_14,n14_3_r_14);
nor I_28(n11_3_r_14,G199_5_l_14,n12_3_r_14);
nor I_29(n13_3_r_14,G199_1_l_14,G199_5_l_14);
and I_30(n14_3_r_14,n_42_5_l_14,n15_3_r_14);
nor I_31(n15_3_r_14,G199_1_l_14,n16_3_r_14);
not I_32(n16_3_r_14,G214_1_l_14);
nand I_33(n_429_or_0_3_r_10,n_266_and_0_0_l_10,n12_3_r_10);
DFFARX1 I_34(n_431_3_r_10,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_10,);
nand I_35(n_576_3_r_10,ACVQN2_0_l_10,n11_3_r_10);
not I_36(n_102_3_r_10,G42_4_l_10);
nand I_37(n_547_3_r_10,n_569_4_l_10,n13_3_r_10);
DFFARX1 I_38(n4_4_r_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_10,);
nor I_39(n_572_4_r_10,ACVQN2_0_l_10,n_573_4_l_10);
or I_40(n_573_4_r_10,n_569_4_l_10,n_452_4_l_10);
nor I_41(n_549_4_r_10,n_572_4_l_10,n7_4_r_10);
or I_42(n_569_4_r_10,n_572_4_l_10,n_569_4_l_10);
nor I_43(n_452_4_r_10,n_266_and_0_0_l_10,n_452_4_l_10);
not I_44(n2_3_r_10,blif_reset_net_3_r_10);
DFFARX1 I_45(n_547_3_r_14,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_10,);
and I_46(n_266_and_0_0_l_10,ACVQN1_0_l_10,n_576_3_r_14);
DFFARX1 I_47(P6_2_r_14,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_10,);
nor I_48(n4_4_l_10,G78_3_r_14,n_102_3_r_14);
DFFARX1 I_49(n4_4_l_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_l_10,);
not I_50(n_87_4_l_10,G214_1_r_14);
nor I_51(n_572_4_l_10,G199_1_r_14,G214_1_r_14);
or I_52(n_573_4_l_10,ACVQN1_2_r_14,n_429_or_0_3_r_14);
nor I_53(n_549_4_l_10,n7_4_l_10,n_266_and_0_0_r_14);
and I_54(n7_4_l_10,n_87_4_l_10,ACVQN2_0_r_14);
or I_55(n_569_4_l_10,n_266_and_0_0_r_14,ACVQN1_2_r_14);
nor I_56(n_452_4_l_10,n_429_or_0_3_r_14,G78_3_r_14);
not I_57(n12_3_r_10,n_549_4_l_10);
or I_58(n_431_3_r_10,n_572_4_l_10,n14_3_r_10);
nor I_59(n11_3_r_10,G42_4_l_10,n12_3_r_10);
nor I_60(n13_3_r_10,G42_4_l_10,n_549_4_l_10);
and I_61(n14_3_r_10,ACVQN2_0_l_10,n15_3_r_10);
nor I_62(n15_3_r_10,n_573_4_l_10,n16_3_r_10);
not I_63(n16_3_r_10,n_266_and_0_0_l_10);
nor I_64(n4_4_r_10,n_266_and_0_0_l_10,G42_4_l_10);
not I_65(n_87_4_r_10,ACVQN2_0_l_10);
and I_66(n7_4_r_10,n_452_4_l_10,n_87_4_r_10);
endmodule


