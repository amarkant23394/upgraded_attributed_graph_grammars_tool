module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_5_r_11,n9_11,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
not I_44(N1372_1_r_11,n53_11);
nor I_45(N1508_1_r_11,n39_11,n53_11);
nor I_46(N6147_2_r_11,n48_11,n49_11);
nor I_47(N6147_3_r_11,n44_11,n45_11);
nand I_48(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_49(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_50(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_51(n_102_5_r_11,n39_11);
nand I_52(n_547_5_r_11,n36_11,n37_11);
nor I_53(N1507_6_r_11,n52_11,n57_11);
nor I_54(N1508_6_r_11,n46_11,n51_11);
nor I_55(N1372_10_r_11,n43_11,n47_11);
nor I_56(N1508_10_r_11,n55_11,n56_11);
nand I_57(n_431_5_r_11,n40_11,n41_11);
not I_58(n9_11,blif_reset_net_5_r_11);
nor I_59(n36_11,n38_11,n39_11);
not I_60(n37_11,n40_11);
nor I_61(n38_11,n60_11,N6147_3_r_10);
nor I_62(n39_11,n54_11,N6147_3_r_10);
nand I_63(n40_11,N6147_2_r_10,n_42_8_r_10);
nand I_64(n41_11,n_102_5_r_11,n42_11);
and I_65(n42_11,n58_11,N6147_9_r_10);
not I_66(n43_11,n44_11);
nor I_67(n44_11,n40_11,G199_8_r_10);
nand I_68(n45_11,n46_11,n47_11);
not I_69(n46_11,n38_11);
nand I_70(n47_11,n59_11,n62_11);
and I_71(n48_11,n37_11,n47_11);
or I_72(n49_11,n44_11,n50_11);
nor I_73(n50_11,n60_11,n61_11);
or I_74(n51_11,n_102_5_r_11,n52_11);
nor I_75(n52_11,n42_11,n57_11);
nand I_76(n53_11,n37_11,n50_11);
or I_77(n54_11,N1371_0_r_10,N1508_6_r_10);
nor I_78(n55_11,n38_11,n42_11);
not I_79(n56_11,N1372_10_r_11);
and I_80(n57_11,n38_11,n50_11);
and I_81(n58_11,n59_11,N6134_9_r_10);
or I_82(n59_11,n63_11,N1508_0_r_10);
not I_83(n60_11,N6147_2_r_10);
nor I_84(n61_11,N1508_0_r_10,N1508_4_r_10);
nand I_85(n62_11,N1507_6_r_10,N1371_0_r_10);
and I_86(n63_11,N1507_6_r_10,N1371_0_r_10);
endmodule


