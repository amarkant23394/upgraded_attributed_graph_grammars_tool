module test_I3969(I2810,I1431,I4017,I1447,I2844,I2980,I1470_clk,I1477_rst,I3969);
input I2810,I1431,I4017,I1447,I2844,I2980,I1470_clk,I1477_rst;
output I3969;
wire I4325,I4034,I3310,I3983_rst,I3124,I3076,I3217,I3107,I4308,I4246,I3200,I2759_rst,I2727,I2745,I4263,I4051,I2733;
and I_0(I4325,I4308,I4051);
DFFARX1 I_1 (I4017,I1470_clk,I3983_rst,I4034);
and I_2(I3310,I2844);
not I_3(I3983_rst,I1477_rst);
nor I_4(I3969,I4263,I4325);
nor I_5(I3124,I3076);
DFFARX1 I_6 (I1447,I1470_clk,I2759_rst,I3076);
not I_7(I3217,I3200);
nor I_8(I3107,I3076,I2844);
DFFARX1 I_9 (I2727,I1470_clk,I3983_rst,I4308);
DFFARX1 I_10 (I2745,I1470_clk,I3983_rst,I4246);
DFFARX1 I_11 (I1431,I1470_clk,I2759_rst,I3200);
not I_12(I2759_rst,I1477_rst);
nand I_13(I2727,I2810,I3124);
nor I_14(I2745,I2980,I3310);
and I_15(I4263,I4246,I2733);
not I_16(I4051,I4034);
nand I_17(I2733,I3217,I3107);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule