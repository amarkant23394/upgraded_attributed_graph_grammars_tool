module test_I14982(I12865,I1477,I1470,I14982);
input I12865,I1477,I1470;
output I14982;
wire I12619,I13023,I12718,I10615,I12596,I13119,I13102,I10639;
not I_0(I12619,I1477);
DFFARX1 I_1(I1470,I12619,,,I13023,);
nor I_2(I12718,I10615,I10639);
not I_3(I14982,I12596);
DFFARX1 I_4(I1470,,,I10615,);
DFFARX1 I_5(I13119,I1470,I12619,,,I12596,);
or I_6(I13119,I12718,I13102);
and I_7(I13102,I13023,I12865);
DFFARX1 I_8(I1470,,,I10639,);
endmodule


