module test_I2617(I1410,I1322,I1294,I1639,I1301,I2617);
input I1410,I1322,I1294,I1639,I1301;
output I2617;
wire I1316,I1342,I2005,I2313,I1937,I2022,I2039,I1908,I2234,I1331,I1509,I1304,I1954,I1926;
nand I_0(I1316,I1509);
not I_1(I1342,I1301);
nor I_2(I2005,I1954);
DFFARX1 I_3(I1331,I1294,I1937,,,I2313,);
not I_4(I1937,I1301);
nand I_5(I2022,I2005,I1316);
DFFARX1 I_6(I2022,I1294,I1937,,,I2039,);
not I_7(I1908,I2039);
nand I_8(I2234,I1954,I1304);
nor I_9(I2617,I1908,I1926);
nor I_10(I1331,I1639,I1410);
DFFARX1 I_11(I1294,I1342,,,I1509,);
DFFARX1 I_12(I1509,I1294,I1342,,,I1304,);
not I_13(I1954,I1322);
nor I_14(I1926,I2313,I2234);
endmodule


