module test_final(IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_5_r,blif_reset_net_5_r,N6147_2_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_5_r,blif_reset_net_5_r;
output N6147_2_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N6147_2_l,n5_2_l,n6_2_l,N6138_2_l,n7_2_l,N1372_4_l,N1508_4_l,n6_4_l,n7_4_l,n8_4_l,N6150_9_l,N6147_9_l,N6134_9_l,n3_9_l,I_BUFF_1_9_l,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n6_4_r,n7_4_r,n8_4_r,n_431_5_r,n2_5_r,n11_5_r,n12_5_r,n13_5_r,n14_5_r,n15_5_r,n16_5_r,N3_8_r,n3_8_r,N6150_9_r,n3_9_r;
nor I_0(N6147_2_l,n5_2_l,n6_2_l);
nor I_1(n5_2_l,IN_5_2_l,n7_2_l);
not I_2(n6_2_l,N6138_2_l);
nor I_3(N6138_2_l,IN_1_2_l,IN_2_2_l);
nor I_4(n7_2_l,IN_3_2_l,IN_4_2_l);
not I_5(N1372_4_l,n7_4_l);
nor I_6(N1508_4_l,n6_4_l,n7_4_l);
nor I_7(n6_4_l,IN_5_4_l,n8_4_l);
nand I_8(n7_4_l,IN_1_4_l,IN_2_4_l);
and I_9(n8_4_l,IN_3_4_l,IN_4_4_l);
not I_10(N6150_9_l,IN_2_9_l);
nor I_11(N6147_9_l,N6150_9_l,n3_9_l);
nor I_12(N6134_9_l,IN_5_9_l,n3_9_l);
nor I_13(n3_9_l,IN_3_9_l,IN_4_9_l);
buf I_14(I_BUFF_1_9_l,IN_1_9_l);
nor I_15(N6147_2_r,n5_2_r,n6_2_r);
nor I_16(n5_2_r,n7_2_r,N1372_4_l);
not I_17(n6_2_r,N6138_2_r);
nor I_18(N6138_2_r,I_BUFF_1_9_l,N6147_2_l);
nor I_19(n7_2_r,N6147_2_l,N1508_4_l);
not I_20(N1372_4_r,n7_4_r);
nor I_21(N1508_4_r,n6_4_r,n7_4_r);
nor I_22(n6_4_r,n8_4_r,N1372_4_l);
nand I_23(n7_4_r,N6134_9_l,I_BUFF_1_9_l);
and I_24(n8_4_r,N6147_2_l,N6134_9_l);
nand I_25(n_429_or_0_5_r,n12_5_r,N1508_4_l);
DFFARX1 I_26(n_431_5_r,blif_clk_net_5_r,n2_5_r,G78_5_r,);
nand I_27(n_576_5_r,n11_5_r,N1508_4_l);
not I_28(n_102_5_r,N6134_9_l);
nand I_29(n_547_5_r,n13_5_r,I_BUFF_1_9_l);
or I_30(n_431_5_r,n14_5_r,N6147_9_l);
not I_31(n2_5_r,blif_reset_net_5_r);
nor I_32(n11_5_r,n12_5_r,N6134_9_l);
not I_33(n12_5_r,N6147_9_l);
nor I_34(n13_5_r,N6134_9_l,N6147_2_l);
and I_35(n14_5_r,n15_5_r,N6147_9_l);
nor I_36(n15_5_r,n16_5_r,N6147_9_l);
not I_37(n16_5_r,N1508_4_l);
nor I_38(n_42_8_r,N1508_4_l,N1372_4_l);
DFFARX1 I_39(N3_8_r,blif_clk_net_5_r,n2_5_r,G199_8_r,);
and I_40(N3_8_r,n3_8_r,N1508_4_l);
nand I_41(n3_8_r,N1508_4_l,N6134_9_l);
not I_42(N6150_9_r,N1372_4_l);
nor I_43(N6147_9_r,N6150_9_r,n3_9_r);
nor I_44(N6134_9_r,n3_9_r,N6134_9_l);
nor I_45(n3_9_r,N6147_9_l,N6147_2_l);
buf I_46(I_BUFF_1_9_r,N1372_4_l);
endmodule


