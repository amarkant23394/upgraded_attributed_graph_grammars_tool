module test_I9525(I8753,I1477,I8674,I8377,I8250,I5737,I8233,I1470,I9525);
input I8753,I1477,I8674,I8377,I8250,I5737,I8233,I1470;
output I9525;
wire I8527,I8202,I8496,I9508,I8770,I8216,I8561,I8184,I8462,I8267,I8199,I5713,I8544;
nand I_0(I8527,I8233,I5713);
nand I_1(I8202,I8267,I8496);
nor I_2(I8496,I8462,I8377);
and I_3(I9525,I9508,I8184);
nand I_4(I9508,I8199,I8202);
or I_5(I8770,I8753,I8674);
not I_6(I8216,I1477);
and I_7(I8561,I8527,I8544);
DFFARX1 I_8(I8561,I1470,I8216,,,I8184,);
DFFARX1 I_9(I1470,I8216,,,I8462,);
nand I_10(I8267,I8250,I5737);
DFFARX1 I_11(I8770,I1470,I8216,,,I8199,);
DFFARX1 I_12(I1470,,,I5713,);
nand I_13(I8544,I8527,I8462);
endmodule


