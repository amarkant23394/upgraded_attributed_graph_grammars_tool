module test_I8830(I1477,I6992,I7026,I1470,I8830);
input I1477,I6992,I7026,I1470;
output I8830;
wire I7190,I6893,I6878,I9179,I6907,I8896,I8913,I8981,I7269,I8862,I7286,I6896,I7156,I6872,I9227,I8964;
DFFARX1 I_0(I7156,I1470,I6907,,,I7190,);
nand I_1(I8830,I8913,I9227);
nand I_2(I6893,I7156,I7286);
not I_3(I6878,I7190);
DFFARX1 I_4(I6896,I1470,I8862,,,I9179,);
not I_5(I6907,I1477);
nor I_6(I8896,I6893,I6872);
nand I_7(I8913,I8896,I6878);
not I_8(I8981,I8964);
DFFARX1 I_9(I1470,I6907,,,I7269,);
not I_10(I8862,I1477);
nor I_11(I7286,I7269,I6992);
nor I_12(I6896,I6992,I7026);
DFFARX1 I_13(I1470,I6907,,,I7156,);
DFFARX1 I_14(I7269,I1470,I6907,,,I6872,);
nor I_15(I9227,I9179,I8981);
not I_16(I8964,I6893);
endmodule


