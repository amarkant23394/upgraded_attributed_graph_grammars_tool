module test_I1331(I1223,I1255,I1294,I1239,I1207,I1301,I1331);
input I1223,I1255,I1294,I1239,I1207,I1301;
output I1331;
wire I1410,I1622,I1342,I1639;
nor I_0(I1410,I1223,I1239);
DFFARX1 I_1(I1255,I1294,I1342,,,I1622,);
not I_2(I1342,I1301);
nor I_3(I1331,I1639,I1410);
and I_4(I1639,I1622,I1207);
endmodule


