module test_I4530(I1477,I1470,I1303,I4578,I2695,I4530);
input I1477,I1470,I1303,I4578,I2695;
output I4530;
wire I2540,I2143,I2181,I4544,I2170,I2557,I4869,I4886,I2149,I4595,I2232,I4807,I4824,I4612;
DFFARX1 I_0(I1470,I2181,,,I2540,);
DFFARX1 I_1(I2557,I1470,I2181,,,I2143,);
not I_2(I2181,I1477);
not I_3(I4544,I1477);
not I_4(I2170,I2232);
and I_5(I2557,I2540,I1303);
DFFARX1 I_6(I2149,I1470,I4544,,,I4869,);
and I_7(I4886,I4869,I4612);
DFFARX1 I_8(I2695,I1470,I2181,,,I2149,);
DFFARX1 I_9(I4578,I1470,I4544,,,I4595,);
DFFARX1 I_10(I1470,I2181,,,I2232,);
DFFARX1 I_11(I2170,I1470,I4544,,,I4807,);
and I_12(I4824,I4807,I2143);
nor I_13(I4530,I4824,I4886);
not I_14(I4612,I4595);
endmodule


