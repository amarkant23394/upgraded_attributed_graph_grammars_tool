module test_I6411(I3954,I1477,I1470,I3969,I6411);
input I3954,I1477,I1470,I3969;
output I6411;
wire I3963,I6346,I6363,I6380,I6329,I4181,I4034;
nor I_0(I3963,I4181,I4034);
nand I_1(I6346,I3969,I3954);
and I_2(I6363,I6346,I3963);
DFFARX1 I_3(I6363,I1470,I6329,,,I6380,);
not I_4(I6329,I1477);
DFFARX1 I_5(I1470,,,I4181,);
DFFARX1 I_6(I6380,I1470,I6329,,,I6411,);
DFFARX1 I_7(I1470,,,I4034,);
endmodule


