module test_I2634(I2022,I1294,I1331,I1954,I1988,I1301,I2634);
input I2022,I1294,I1331,I1954,I1988,I1301;
output I2634;
wire I2268,I1304,I2313,I2251,I1937,I2039,I1908,I2234,I2617,I2070,I1929,I1310,I1926;
and I_0(I2268,I2070,I2251);
DFFARX1 I_1(I1294,,,I1304,);
DFFARX1 I_2(I1331,I1294,I1937,,,I2313,);
nand I_3(I2251,I2234,I1988);
not I_4(I1937,I1301);
DFFARX1 I_5(I2022,I1294,I1937,,,I2039,);
not I_6(I1908,I2039);
nand I_7(I2234,I1954,I1304);
nand I_8(I2634,I2617,I1929);
nor I_9(I2617,I1908,I1926);
not I_10(I2070,I1310);
DFFARX1 I_11(I2268,I1294,I1937,,,I1929,);
DFFARX1 I_12(I1294,,,I1310,);
nor I_13(I1926,I2313,I2234);
endmodule


