module test_I2764(I1937,I1331,I1294,I1954,I1687,I2764);
input I1937,I1331,I1294,I1954,I1687;
output I2764;
wire I1316,I2344,I2005,I2313,I1971,I2022,I1923,I1988,I1509,I1334,I1310;
not I_0(I2764,I1923);
nand I_1(I1316,I1509,I1687);
nor I_2(I2344,I2313,I1988);
nor I_3(I2005,I1954,I1310);
DFFARX1 I_4(I1331,I1294,I1937,,,I2313,);
nor I_5(I1971,I1310);
nand I_6(I2022,I2005,I1316);
nand I_7(I1923,I2022,I2344);
nand I_8(I1988,I1971,I1334);
DFFARX1 I_9(I1294,,,I1509,);
DFFARX1 I_10(I1294,,,I1334,);
DFFARX1 I_11(I1294,,,I1310,);
endmodule


