module test_I2945(I1322,I1294,I2155,I1301,I2945);
input I1322,I1294,I2155,I1301;
output I2945;
wire I2172,I2583,I1902,I2203,I2234,I1937,I1342,I1954,I1509,I1304;
DFFARX1 I_0(I2155,I1294,I1937,,,I2172,);
not I_1(I2583,I1301);
and I_2(I1902,I2234,I2203);
DFFARX1 I_3(I2172,I1294,I1937,,,I2203,);
nand I_4(I2234,I1954,I1304);
not I_5(I1937,I1301);
not I_6(I1342,I1301);
not I_7(I1954,I1322);
DFFARX1 I_8(I1294,I1342,,,I1509,);
DFFARX1 I_9(I1509,I1294,I1342,,,I1304,);
DFFARX1 I_10(I1902,I1294,I2583,,,I2945,);
endmodule


