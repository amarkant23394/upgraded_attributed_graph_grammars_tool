module test_I9542(I8770,I8527,I8267,I8496,I1477,I1470,I9542);
input I8770,I8527,I8267,I8496,I1477,I1470;
output I9542;
wire I9508,I8202,I8216,I8199,I8544,I8184,I8561,I9525,I9491;
nand I_0(I9508,I8199,I8202);
DFFARX1 I_1(I9525,I1470,I9491,,,I9542,);
nand I_2(I8202,I8267,I8496);
not I_3(I8216,I1477);
DFFARX1 I_4(I8770,I1470,I8216,,,I8199,);
nand I_5(I8544,I8527);
DFFARX1 I_6(I8561,I1470,I8216,,,I8184,);
and I_7(I8561,I8527,I8544);
and I_8(I9525,I9508,I8184);
not I_9(I9491,I1477);
endmodule


