module test_final(IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_2,n_572_1_r_2,n_573_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2,N3_2_l_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n4_1_r_2,blif_clk_net_1_r_1,n5_1,G42_1_r_2,);
nor I_1(n_572_1_r_2,n26_2,n18_2);
nand I_2(n_573_1_r_2,n17_2,n19_2);
nor I_3(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_4(n_569_1_r_2,n13_2,n19_2);
not I_5(n_452_1_r_2,n_573_1_r_2);
nor I_6(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_7(N3_2_r_2,blif_clk_net_1_r_1,n5_1,G199_2_r_2,);
DFFARX1 I_8(ACVQN2_3_l_2,blif_clk_net_1_r_1,n5_1,ACVQN1_5_r_2,);
not I_9(P6_5_r_2,P6_5_r_internal_2);
and I_10(N3_2_l_2,IN_6_2_l_2,n24_2);
DFFARX1 I_11(N3_2_l_2,blif_clk_net_1_r_1,n5_1,G199_2_l_2,);
not I_12(n13_2,G199_2_l_2);
DFFARX1 I_13(IN_1_3_l_2,blif_clk_net_1_r_1,n5_1,ACVQN2_3_l_2,);
DFFARX1 I_14(IN_2_3_l_2,blif_clk_net_1_r_1,n5_1,n16_2,);
and I_15(N1_4_l_2,IN_6_4_l_2,n25_2);
DFFARX1 I_16(N1_4_l_2,blif_clk_net_1_r_1,n5_1,n26_2,);
DFFARX1 I_17(IN_3_4_l_2,blif_clk_net_1_r_1,n5_1,n17_internal_2,);
not I_18(n17_2,n17_internal_2);
nor I_19(n4_1_r_2,n26_2,n22_2);
nor I_20(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_21(G199_2_l_2,blif_clk_net_1_r_1,n5_1,P6_5_r_internal_2,);
nor I_22(n18_2,IN_1_2_l_2,IN_3_2_l_2);
nand I_23(n19_2,IN_4_3_l_2,n16_2);
nor I_24(n20_2,n26_2,n21_2);
not I_25(n21_2,n18_2);
and I_26(n22_2,IN_4_3_l_2,n16_2);
nor I_27(n23_2,n13_2,n21_2);
nand I_28(n24_2,IN_2_2_l_2,IN_3_2_l_2);
nand I_29(n25_2,IN_1_4_l_2,IN_2_4_l_2);
DFFARX1 I_30(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_31(n_572_1_r_1,n26_1,n19_1);
nand I_32(n_573_1_r_1,n16_1,n18_1);
nor I_33(n_549_1_r_1,n20_1,n21_1);
nor I_34(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_35(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_36(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_37(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_38(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_39(N3_2_l_1,n23_1,n_452_1_r_2);
not I_40(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_41(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_42(n17_1,n26_1);
DFFARX1 I_43(G199_2_r_2,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_44(n16_1,n16_internal_1);
DFFARX1 I_45(n_42_2_r_2,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_46(N1_4_l_1,n25_1,n_569_1_r_2);
DFFARX1 I_47(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_48(G42_1_r_2,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_49(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_50(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_51(n14_1,n14_internal_1);
nor I_52(N1_4_r_1,n17_1,n24_1);
nand I_53(n18_1,ACVQN1_3_l_1,n_572_1_r_2);
nor I_54(n19_1,G42_1_r_2,n_549_1_r_2);
not I_55(n20_1,n18_1);
nor I_56(n21_1,n26_1,n22_1);
not I_57(n22_1,n19_1);
nand I_58(n23_1,G42_1_r_2,n_572_1_r_2);
nor I_59(n24_1,n18_1,n22_1);
nand I_60(n25_1,ACVQN1_5_r_2,P6_5_r_2);
endmodule


