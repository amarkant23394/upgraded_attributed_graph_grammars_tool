module test_I15582(I1477,I14066,I1470,I15582);
input I1477,I14066,I1470;
output I15582;
wire I14083,I13746,I13775,I15611,I15928;
not I_0(I15582,I15928);
DFFARX1 I_1(I14066,I1470,I13775,,,I14083,);
not I_2(I13746,I14083);
not I_3(I13775,I1477);
not I_4(I15611,I1477);
DFFARX1 I_5(I13746,I1470,I15611,,,I15928,);
endmodule


