module test_I2897(I1294,I1331,I1954,I2406,I1687,I1937,I2897);
input I1294,I1331,I1954,I2406,I1687,I1937;
output I2897;
wire I1911,I2005,I2313,I2022,I1316,I2600,I1971,I1334,I1310,I2488,I2344,I2070,I1923,I1988,I1509;
nand I_0(I1911,I2070,I2488);
nor I_1(I2005,I1954,I1310);
DFFARX1 I_2(I1331,I1294,I1937,,,I2313,);
nand I_3(I2022,I2005,I1316);
nand I_4(I1316,I1509,I1687);
nand I_5(I2897,I2600,I1923);
not I_6(I2600,I1911);
nor I_7(I1971,I1310);
DFFARX1 I_8(I1294,,,I1334,);
DFFARX1 I_9(I1294,,,I1310,);
not I_10(I2488,I2406);
nor I_11(I2344,I2313,I1988);
not I_12(I2070,I1310);
nand I_13(I1923,I2022,I2344);
nand I_14(I1988,I1971,I1334);
DFFARX1 I_15(I1294,,,I1509,);
endmodule


