module test_I4356(I2878,I1447,I1477,I1470,I2793,I1335,I4356);
input I2878,I1447,I1477,I1470,I2793,I1335;
output I4356;
wire I2810,I3217,I2759,I3124,I2727,I3200,I4113,I3076,I4308,I2751,I3983;
nand I_0(I2810,I2793,I1335);
not I_1(I3217,I3200);
not I_2(I2759,I1477);
nor I_3(I3124,I3076,I2878);
nand I_4(I2727,I2810,I3124);
DFFARX1 I_5(I1470,I2759,,,I3200,);
DFFARX1 I_6(I2751,I1470,I3983,,,I4113,);
DFFARX1 I_7(I1447,I1470,I2759,,,I3076,);
DFFARX1 I_8(I2727,I1470,I3983,,,I4308,);
nor I_9(I4356,I4308,I4113);
nor I_10(I2751,I3076,I3217);
not I_11(I3983,I1477);
endmodule


