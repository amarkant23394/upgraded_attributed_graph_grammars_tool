module test_I7587(I1477,I6572,I1470,I7587);
input I1477,I6572,I1470;
output I7587;
wire I6606,I3960,I6589,I6329,I6300;
DFFARX1 I_0(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_1(I1470,,,I3960,);
and I_2(I6589,I6572,I3960);
not I_3(I6329,I1477);
not I_4(I7587,I6300);
DFFARX1 I_5(I6606,I1470,I6329,,,I6300,);
endmodule


