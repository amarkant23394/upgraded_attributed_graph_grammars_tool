module test_I5073(I1477,I5334,I3589,I1470,I5073);
input I1477,I5334,I3589,I1470;
output I5073;
wire I5416,I5450,I3388,I5351,I3350,I5433,I5122,I3356,I5105;
nand I_0(I5416,I5122,I3356);
and I_1(I5450,I5416,I5433);
not I_2(I3388,I1477);
DFFARX1 I_3(I5334,I1470,I5105,,,I5351,);
DFFARX1 I_4(I5450,I1470,I5105,,,I5073,);
DFFARX1 I_5(I1470,I3388,,,I3350,);
nand I_6(I5433,I5416,I5351);
not I_7(I5122,I3350);
DFFARX1 I_8(I3589,I1470,I3388,,,I3356,);
not I_9(I5105,I1477);
endmodule


