module test_I14939(I1477,I1470,I14939);
input I1477,I1470;
output I14939;
wire I12619,I12670,I15016,I12584,I14999,I12590,I12930,I12783,I12752,I12913,I14965,I12581,I10609;
not I_0(I12619,I1477);
DFFARX1 I_1(I1470,I12619,,,I12670,);
nand I_2(I15016,I14999,I12581);
and I_3(I12584,I12670,I12783);
nor I_4(I14999,I12584,I12590);
not I_5(I12590,I12752);
and I_6(I12930,I12913,I10609);
DFFARX1 I_7(I1470,I12619,,,I12783,);
DFFARX1 I_8(I1470,I12619,,,I12752,);
DFFARX1 I_9(I1470,I12619,,,I12913,);
DFFARX1 I_10(I15016,I1470,I14965,,,I14939,);
not I_11(I14965,I1477);
DFFARX1 I_12(I12930,I1470,I12619,,,I12581,);
DFFARX1 I_13(I1470,,,I10609,);
endmodule


