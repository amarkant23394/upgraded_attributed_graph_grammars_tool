module test_final(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470,I1477,I16208,I16211,I16205,I16214,I16220,I16223,I16202,I16232,I16229,I16217,I16226,I16801,I16804,I16786,I16807,I16798,I16789,I16780,I16810,I16795,I16792,I16783,I17402,I17387,I17384,I17381,I17399,I17396,I17375,I17378,I17405,I17390,I17393);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1470,I1477;
output I16208,I16211,I16205,I16214,I16220,I16223,I16202,I16232,I16229,I16217,I16226,I16801,I16804,I16786,I16807,I16798,I16789,I16780,I16810,I16795,I16792,I16783,I17402,I17387,I17384,I17381,I17399,I17396,I17375,I17378,I17405,I17390,I17393;
wire I1518,I1535,I1552,I1569,I1586,I1603,I1620,I1637,I1507,I1668,I1492,I1699,I1716,I1733,I1750,I1767,I1784,I1801,I1489,I1832,I1849,I1486,I1880,I1897,I1504,I1928,I1501,I1959,I1976,I1480,I1483,I2021,I2038,I2055,I2072,I1510,I2103,I1495,I1498,I2181,I2198,I2215,I2232,I2170,I2263,I2158,I2294,I2311,I2328,I2345,I2362,I2161,I2393,I2146,I2424,I2441,I2458,I2475,I2492,I2509,I2152,I2540,I2557,I2574,I2164,I2173,I2143,I2633,I2167,I2155,I2678,I2695,I2149,I2759,I2776,I2793,I2810,I2827,I2844,I2861,I2878,I2895,I2912,I2929,I2946,I2963,I2980,I2748,I3011,I3028,I3045,I2721,I3076,I2742,I3107,I3124,I2727,I3155,I2724,I2730,I3200,I3217,I3234,I2736,I2751,I2739,I3293,I3310,I2745,I2733,I3388,I3405,I3422,I3362,I3453,I3470,I3487,I3504,I3521,I3538,I3555,I3572,I3589,I3356,I3620,I3637,I3353,I3668,I3685,I3702,I3365,I3350,I3747,I3764,I3781,I3798,I3815,I3371,I3846,I3380,I3877,I3374,I3377,I3368,I3359,I3983,I4000,I4017,I4034,I4051,I4068,I3966,I3954,I4113,I4130,I4147,I4164,I4181,I3963,I4212,I4229,I4246,I4263,I3972,I3951,I4308,I4325,I3969,I4356,I3960,I3975,I4401,I4418,I4435,I4452,I3948,I3957,I3945,I4544,I4561,I4578,I4595,I4612,I4629,I4527,I4515,I4674,I4691,I4708,I4725,I4742,I4524,I4773,I4790,I4807,I4824,I4533,I4512,I4869,I4886,I4530,I4917,I4521,I4536,I4962,I4979,I4996,I5013,I4509,I4518,I4506,I5105,I5122,I5139,I5156,I5079,I5187,I5204,I5094,I5076,I5249,I5266,I5283,I5300,I5317,I5334,I5351,I5368,I5385,I5091,I5416,I5433,I5450,I5073,I5481,I5070,I5512,I5529,I5546,I5563,I5085,I5594,I5082,I5625,I5642,I5659,I5088,I5097,I5067,I5751,I5768,I5785,I5802,I5740,I5833,I5728,I5864,I5881,I5898,I5915,I5932,I5731,I5963,I5716,I5994,I6011,I6028,I6045,I6062,I6079,I5722,I6110,I6127,I6144,I5734,I5743,I5713,I6203,I5737,I5725,I6248,I6265,I5719,I6329,I6346,I6363,I6380,I6318,I6411,I6306,I6442,I6459,I6476,I6493,I6510,I6309,I6541,I6294,I6572,I6589,I6606,I6623,I6640,I6657,I6300,I6688,I6705,I6722,I6312,I6321,I6291,I6781,I6315,I6303,I6826,I6843,I6297,I6907,I6924,I6941,I6958,I6975,I6992,I7009,I7026,I6896,I7057,I6881,I7088,I7105,I7122,I7139,I7156,I7173,I7190,I6878,I7221,I7238,I6875,I7269,I7286,I6893,I7317,I6890,I7348,I7365,I6869,I6872,I7410,I7427,I7444,I7461,I6899,I7492,I6884,I6887,I7570,I7587,I7604,I7621,I7544,I7652,I7669,I7559,I7541,I7714,I7731,I7748,I7765,I7782,I7799,I7816,I7833,I7850,I7556,I7881,I7898,I7915,I7538,I7946,I7535,I7977,I7994,I8011,I8028,I7550,I8059,I7547,I8090,I8107,I8124,I7553,I7562,I7532,I8216,I8233,I8250,I8267,I8190,I8298,I8315,I8205,I8187,I8360,I8377,I8394,I8411,I8428,I8445,I8462,I8479,I8496,I8202,I8527,I8544,I8561,I8184,I8592,I8181,I8623,I8640,I8657,I8674,I8196,I8705,I8193,I8736,I8753,I8770,I8199,I8208,I8178,I8862,I8879,I8896,I8913,I8930,I8947,I8964,I8981,I8998,I9015,I9032,I9049,I9066,I9083,I8851,I9114,I9131,I9148,I8824,I9179,I8845,I9210,I9227,I8830,I9258,I8827,I8833,I9303,I9320,I9337,I8839,I8854,I8842,I9396,I9413,I8848,I8836,I9491,I9508,I9525,I9542,I9559,I9576,I9474,I9462,I9621,I9638,I9655,I9672,I9689,I9471,I9720,I9737,I9754,I9771,I9480,I9459,I9816,I9833,I9477,I9864,I9468,I9483,I9909,I9926,I9943,I9960,I9456,I9465,I9453,I10052,I10069,I10086,I10103,I10120,I10137,I10154,I10023,I10185,I10202,I10219,I10236,I10253,I10270,I10287,I10020,I10014,I10332,I10349,I10366,I10041,I10397,I10414,I10032,I10026,I10459,I10029,I10490,I10507,I10044,I10538,I10038,I10035,I10583,I10017,I10647,I10664,I10681,I10698,I10715,I10732,I10749,I10766,I10636,I10797,I10621,I10828,I10845,I10862,I10879,I10896,I10913,I10930,I10618,I10961,I10978,I10615,I11009,I11026,I10633,I11057,I10630,I11088,I11105,I10609,I10612,I11150,I11167,I11184,I11201,I10639,I11232,I10624,I10627,I11310,I11327,I11344,I11361,I11378,I11395,I11412,I11429,I11299,I11460,I11284,I11491,I11508,I11525,I11542,I11559,I11576,I11593,I11281,I11624,I11641,I11278,I11672,I11689,I11296,I11720,I11293,I11751,I11768,I11272,I11275,I11813,I11830,I11847,I11864,I11302,I11895,I11287,I11290,I11973,I11990,I12007,I12024,I12041,I12058,I12075,I11944,I12106,I12123,I12140,I12157,I12174,I12191,I12208,I11941,I12239,I11935,I12270,I12287,I12304,I11965,I11938,I12349,I11962,I12380,I11959,I11956,I12425,I12442,I12459,I12476,I12493,I11950,I12524,I12541,I11953,I11947,I12619,I12636,I12653,I12670,I12687,I12587,I12718,I12735,I12752,I12590,I12783,I12584,I12814,I12831,I12848,I12865,I12882,I12593,I12913,I12930,I12947,I12964,I12599,I12602,I12581,I13023,I13040,I13057,I12611,I12608,I13102,I13119,I12596,I12605,I13197,I13214,I13231,I13248,I13265,I13165,I13296,I13313,I13330,I13168,I13361,I13162,I13392,I13409,I13426,I13443,I13460,I13171,I13491,I13508,I13525,I13542,I13177,I13180,I13159,I13601,I13618,I13635,I13189,I13186,I13680,I13697,I13174,I13183,I13775,I13792,I13809,I13826,I13843,I13860,I13758,I13891,I13908,I13925,I13761,I13743,I13970,I13987,I14004,I13764,I13755,I14049,I14066,I14083,I13746,I14114,I14131,I13737,I14162,I14179,I14196,I13767,I14227,I14244,I14261,I14278,I13752,I13749,I13740,I14370,I14387,I14404,I14421,I14438,I14455,I14472,I14341,I14503,I14520,I14537,I14554,I14571,I14588,I14605,I14338,I14332,I14650,I14667,I14684,I14359,I14715,I14732,I14350,I14344,I14777,I14347,I14808,I14825,I14362,I14856,I14356,I14353,I14901,I14335,I14965,I14982,I14999,I15016,I14939,I15047,I15064,I14954,I14936,I15109,I15126,I15143,I15160,I15177,I15194,I15211,I15228,I15245,I14951,I15276,I15293,I15310,I14933,I15341,I14930,I15372,I15389,I15406,I15423,I14945,I15454,I14942,I15485,I15502,I15519,I14948,I14957,I14927,I15611,I15628,I15645,I15662,I15679,I15696,I15713,I15730,I15747,I15764,I15781,I15798,I15815,I15832,I15600,I15863,I15880,I15897,I15573,I15928,I15594,I15959,I15976,I15579,I16007,I15576,I15582,I16052,I16069,I16086,I15588,I15603,I15591,I16145,I16162,I15597,I15585,I16240,I16257,I16274,I16291,I16308,I16339,I16356,I16373,I16404,I16435,I16452,I16469,I16486,I16503,I16534,I16551,I16568,I16585,I16644,I16661,I16678,I16723,I16740,I16818,I16835,I16852,I16869,I16886,I16903,I16934,I16951,I16968,I17013,I17030,I17047,I17092,I17109,I17126,I17157,I17174,I17205,I17222,I17239,I17270,I17287,I17304,I17321,I17413,I17430,I17447,I17464,I17481,I17498,I17515,I17532,I17563,I17594,I17611,I17628,I17645,I17662,I17679,I17696,I17727,I17744,I17775,I17792,I17823,I17854,I17871,I17916,I17933,I17950,I17967,I17998;
DFFARX1 I_0(I16291,I1470,I16240,,,I16208,);
not I_1(I16211,I16373);
and I_2(I16205,I16291,I16404);
nand I_3(I16214,I16291,I16503);
nand I_4(I16220,I16339,I16585);
not I_5(I16223,I16551);
DFFARX1 I_6(I16551,I1470,I16240,,,I16202,);
DFFARX1 I_7(I16678,I1470,I16240,,,I16232,);
nor I_8(I16229,I16644,I16551);
DFFARX1 I_9(I16740,I1470,I16240,,,I16217,);
nand I_10(I16226,I16644,I16568);
not I_11(I16801,I16886);
nand I_12(I16804,I16934,I16903);
DFFARX1 I_13(I16934,I1470,I16818,,,I16786,);
nor I_14(I16807,I17047,I16869);
nand I_15(I16798,I17047,I16968);
not I_16(I16789,I17126);
DFFARX1 I_17(I17174,I1470,I16818,,,I16780,);
DFFARX1 I_18(I17239,I1470,I16818,,,I16810,);
DFFARX1 I_19(I17321,I1470,I16818,,,I16795,);
nand I_20(I16792,I17205,I16951);
DFFARX1 I_21(I17205,I1470,I16818,,,I16783,);
nor I_22(I17402,I17498,I17532);
nand I_23(I17387,I17498,I17563);
not I_24(I17384,I17696);
DFFARX1 I_25(I17727,I1470,I17413,,,I17381,);
nand I_26(I17399,I17662,I17792);
not I_27(I17396,I17775);
DFFARX1 I_28(I17871,I1470,I17413,,,I17375,);
DFFARX1 I_29(I17775,I1470,I17413,,,I17378,);
DFFARX1 I_30(I17967,I1470,I17413,,,I17405,);
DFFARX1 I_31(I17998,I1470,I17413,,,I17390,);
nand I_32(I17393,I17933,I17823);
not I_33(I1518,I1477);
not I_34(I1535,I1455);
nor I_35(I1552,I1215,I1399);
nand I_36(I1569,I1552,I1463);
nor I_37(I1586,I1535,I1215);
nand I_38(I1603,I1586,I1423);
not I_39(I1620,I1603);
not I_40(I1637,I1215);
nor I_41(I1507,I1603,I1637);
not I_42(I1668,I1637);
nand I_43(I1492,I1603,I1668);
not I_44(I1699,I1207);
nor I_45(I1716,I1699,I1367);
and I_46(I1733,I1716,I1439);
or I_47(I1750,I1733,I1279);
DFFARX1 I_48(I1750,I1470,I1518,,,I1767,);
nor I_49(I1784,I1767,I1620);
DFFARX1 I_50(I1767,I1470,I1518,,,I1801,);
not I_51(I1489,I1801);
nand I_52(I1832,I1535,I1207);
and I_53(I1849,I1832,I1784);
DFFARX1 I_54(I1832,I1470,I1518,,,I1486,);
DFFARX1 I_55(I1383,I1470,I1518,,,I1880,);
nor I_56(I1897,I1880,I1603);
nand I_57(I1504,I1767,I1897);
nor I_58(I1928,I1880,I1668);
not I_59(I1501,I1880);
nand I_60(I1959,I1880,I1569);
and I_61(I1976,I1637,I1959);
DFFARX1 I_62(I1976,I1470,I1518,,,I1480,);
DFFARX1 I_63(I1880,I1470,I1518,,,I1483,);
DFFARX1 I_64(I1295,I1470,I1518,,,I2021,);
not I_65(I2038,I2021);
nand I_66(I2055,I2038,I1603);
and I_67(I2072,I1832,I2055);
DFFARX1 I_68(I2072,I1470,I1518,,,I1510,);
or I_69(I2103,I2038,I1849);
DFFARX1 I_70(I2103,I1470,I1518,,,I1495,);
nand I_71(I1498,I2038,I1928);
not I_72(I2181,I1477);
nand I_73(I2198,I1343,I1231);
and I_74(I2215,I2198,I1271);
DFFARX1 I_75(I2215,I1470,I2181,,,I2232,);
not I_76(I2170,I2232);
DFFARX1 I_77(I2232,I1470,I2181,,,I2263,);
not I_78(I2158,I2263);
nor I_79(I2294,I1287,I1231);
not I_80(I2311,I2294);
nor I_81(I2328,I2232,I2311);
DFFARX1 I_82(I1375,I1470,I2181,,,I2345,);
not I_83(I2362,I2345);
nand I_84(I2161,I2345,I2311);
DFFARX1 I_85(I2345,I1470,I2181,,,I2393,);
and I_86(I2146,I2232,I2393);
nand I_87(I2424,I1223,I1255);
and I_88(I2441,I2424,I1327);
DFFARX1 I_89(I2441,I1470,I2181,,,I2458,);
nor I_90(I2475,I2458,I2362);
and I_91(I2492,I2294,I2475);
nor I_92(I2509,I2458,I2232);
DFFARX1 I_93(I2458,I1470,I2181,,,I2152,);
DFFARX1 I_94(I1247,I1470,I2181,,,I2540,);
and I_95(I2557,I2540,I1303);
or I_96(I2574,I2557,I2492);
DFFARX1 I_97(I2574,I1470,I2181,,,I2164,);
nand I_98(I2173,I2557,I2509);
DFFARX1 I_99(I2557,I1470,I2181,,,I2143,);
DFFARX1 I_100(I1239,I1470,I2181,,,I2633,);
nand I_101(I2167,I2633,I2328);
DFFARX1 I_102(I2633,I1470,I2181,,,I2155,);
nand I_103(I2678,I2633,I2294);
and I_104(I2695,I2345,I2678);
DFFARX1 I_105(I2695,I1470,I2181,,,I2149,);
not I_106(I2759,I1477);
not I_107(I2776,I1407);
nor I_108(I2793,I1351,I1319);
nand I_109(I2810,I2793,I1335);
nor I_110(I2827,I2776,I1351);
nand I_111(I2844,I2827,I1359);
not I_112(I2861,I1351);
not I_113(I2878,I2861);
not I_114(I2895,I1415);
nor I_115(I2912,I2895,I1311);
and I_116(I2929,I2912,I1391);
or I_117(I2946,I2929,I1263);
DFFARX1 I_118(I2946,I1470,I2759,,,I2963,);
nand I_119(I2980,I2776,I1415);
or I_120(I2748,I2980,I2963);
not I_121(I3011,I2980);
nor I_122(I3028,I2963,I3011);
and I_123(I3045,I2861,I3028);
nand I_124(I2721,I2980,I2878);
DFFARX1 I_125(I1447,I1470,I2759,,,I3076,);
or I_126(I2742,I3076,I2963);
nor I_127(I3107,I3076,I2844);
nor I_128(I3124,I3076,I2878);
nand I_129(I2727,I2810,I3124);
or I_130(I3155,I3076,I3045);
DFFARX1 I_131(I3155,I1470,I2759,,,I2724,);
not I_132(I2730,I3076);
DFFARX1 I_133(I1431,I1470,I2759,,,I3200,);
not I_134(I3217,I3200);
nor I_135(I3234,I3217,I2810);
DFFARX1 I_136(I3234,I1470,I2759,,,I2736,);
nor I_137(I2751,I3076,I3217);
nor I_138(I2739,I3217,I2980);
not I_139(I3293,I3217);
and I_140(I3310,I2844,I3293);
nor I_141(I2745,I2980,I3310);
nand I_142(I2733,I3217,I3107);
not I_143(I3388,I1477);
or I_144(I3405,I1480,I1495);
or I_145(I3422,I1483,I1480);
DFFARX1 I_146(I3422,I1470,I3388,,,I3362,);
nor I_147(I3453,I1486,I1501);
not I_148(I3470,I3453);
not I_149(I3487,I1486);
and I_150(I3504,I3487,I1489);
nor I_151(I3521,I3504,I1495);
nor I_152(I3538,I1492,I1510);
DFFARX1 I_153(I3538,I1470,I3388,,,I3555,);
nand I_154(I3572,I3555,I3405);
and I_155(I3589,I3521,I3572);
DFFARX1 I_156(I3589,I1470,I3388,,,I3356,);
nor I_157(I3620,I1492,I1483);
DFFARX1 I_158(I3620,I1470,I3388,,,I3637,);
and I_159(I3353,I3453,I3637);
DFFARX1 I_160(I1507,I1470,I3388,,,I3668,);
and I_161(I3685,I3668,I1498);
DFFARX1 I_162(I3685,I1470,I3388,,,I3702,);
not I_163(I3365,I3702);
DFFARX1 I_164(I3685,I1470,I3388,,,I3350,);
DFFARX1 I_165(I1504,I1470,I3388,,,I3747,);
not I_166(I3764,I3747);
nor I_167(I3781,I3422,I3764);
and I_168(I3798,I3685,I3781);
or I_169(I3815,I3405,I3798);
DFFARX1 I_170(I3815,I1470,I3388,,,I3371,);
nor I_171(I3846,I3747,I3555);
nand I_172(I3380,I3521,I3846);
nor I_173(I3877,I3747,I3470);
nand I_174(I3374,I3620,I3877);
not I_175(I3377,I3747);
nand I_176(I3368,I3747,I3470);
DFFARX1 I_177(I3747,I1470,I3388,,,I3359,);
not I_178(I3983,I1477);
nand I_179(I4000,I2721,I2724);
and I_180(I4017,I4000,I2730);
DFFARX1 I_181(I4017,I1470,I3983,,,I4034,);
not I_182(I4051,I4034);
nor I_183(I4068,I2742,I2724);
or I_184(I3966,I4068,I4034);
not I_185(I3954,I4068);
DFFARX1 I_186(I2751,I1470,I3983,,,I4113,);
nor I_187(I4130,I4113,I4068);
nand I_188(I4147,I2739,I2736);
and I_189(I4164,I4147,I2748);
DFFARX1 I_190(I4164,I1470,I3983,,,I4181,);
nor I_191(I3963,I4181,I4034);
not I_192(I4212,I4181);
nor I_193(I4229,I4113,I4212);
DFFARX1 I_194(I2745,I1470,I3983,,,I4246,);
and I_195(I4263,I4246,I2733);
or I_196(I3972,I4263,I4068);
nand I_197(I3951,I4263,I4229);
DFFARX1 I_198(I2727,I1470,I3983,,,I4308,);
and I_199(I4325,I4308,I4051);
nor I_200(I3969,I4263,I4325);
nor I_201(I4356,I4308,I4113);
DFFARX1 I_202(I4356,I1470,I3983,,,I3960,);
nor I_203(I3975,I4308,I4034);
not I_204(I4401,I4308);
nor I_205(I4418,I4181,I4401);
and I_206(I4435,I4068,I4418);
or I_207(I4452,I4263,I4435);
DFFARX1 I_208(I4452,I1470,I3983,,,I3948,);
nand I_209(I3957,I4308,I4130);
nand I_210(I3945,I4308,I4212);
not I_211(I4544,I1477);
nand I_212(I4561,I2152,I2173);
and I_213(I4578,I4561,I2161);
DFFARX1 I_214(I4578,I1470,I4544,,,I4595,);
not I_215(I4612,I4595);
nor I_216(I4629,I2167,I2173);
or I_217(I4527,I4629,I4595);
not I_218(I4515,I4629);
DFFARX1 I_219(I2155,I1470,I4544,,,I4674,);
nor I_220(I4691,I4674,I4629);
nand I_221(I4708,I2146,I2164);
and I_222(I4725,I4708,I2158);
DFFARX1 I_223(I4725,I1470,I4544,,,I4742,);
nor I_224(I4524,I4742,I4595);
not I_225(I4773,I4742);
nor I_226(I4790,I4674,I4773);
DFFARX1 I_227(I2170,I1470,I4544,,,I4807,);
and I_228(I4824,I4807,I2143);
or I_229(I4533,I4824,I4629);
nand I_230(I4512,I4824,I4790);
DFFARX1 I_231(I2149,I1470,I4544,,,I4869,);
and I_232(I4886,I4869,I4612);
nor I_233(I4530,I4824,I4886);
nor I_234(I4917,I4869,I4674);
DFFARX1 I_235(I4917,I1470,I4544,,,I4521,);
nor I_236(I4536,I4869,I4595);
not I_237(I4962,I4869);
nor I_238(I4979,I4742,I4962);
and I_239(I4996,I4629,I4979);
or I_240(I5013,I4824,I4996);
DFFARX1 I_241(I5013,I1470,I4544,,,I4509,);
nand I_242(I4518,I4869,I4691);
nand I_243(I4506,I4869,I4773);
not I_244(I5105,I1477);
not I_245(I5122,I3350);
nor I_246(I5139,I3380,I3359);
nand I_247(I5156,I5139,I3371);
DFFARX1 I_248(I5156,I1470,I5105,,,I5079,);
nor I_249(I5187,I5122,I3380);
nand I_250(I5204,I5187,I3353);
not I_251(I5094,I5204);
DFFARX1 I_252(I5204,I1470,I5105,,,I5076,);
not I_253(I5249,I3380);
not I_254(I5266,I5249);
not I_255(I5283,I3356);
nor I_256(I5300,I5283,I3374);
and I_257(I5317,I5300,I3365);
or I_258(I5334,I5317,I3362);
DFFARX1 I_259(I5334,I1470,I5105,,,I5351,);
nor I_260(I5368,I5351,I5204);
nor I_261(I5385,I5351,I5266);
nand I_262(I5091,I5156,I5385);
nand I_263(I5416,I5122,I3356);
nand I_264(I5433,I5416,I5351);
and I_265(I5450,I5416,I5433);
DFFARX1 I_266(I5450,I1470,I5105,,,I5073,);
DFFARX1 I_267(I5416,I1470,I5105,,,I5481,);
and I_268(I5070,I5249,I5481);
DFFARX1 I_269(I3368,I1470,I5105,,,I5512,);
not I_270(I5529,I5512);
nor I_271(I5546,I5204,I5529);
and I_272(I5563,I5512,I5546);
nand I_273(I5085,I5512,I5266);
DFFARX1 I_274(I5512,I1470,I5105,,,I5594,);
not I_275(I5082,I5594);
DFFARX1 I_276(I3377,I1470,I5105,,,I5625,);
not I_277(I5642,I5625);
or I_278(I5659,I5642,I5563);
DFFARX1 I_279(I5659,I1470,I5105,,,I5088,);
nand I_280(I5097,I5642,I5368);
DFFARX1 I_281(I5642,I1470,I5105,,,I5067,);
not I_282(I5751,I1477);
nand I_283(I5768,I4530,I4515);
and I_284(I5785,I5768,I4524);
DFFARX1 I_285(I5785,I1470,I5751,,,I5802,);
not I_286(I5740,I5802);
DFFARX1 I_287(I5802,I1470,I5751,,,I5833,);
not I_288(I5728,I5833);
nor I_289(I5864,I4536,I4515);
not I_290(I5881,I5864);
nor I_291(I5898,I5802,I5881);
DFFARX1 I_292(I4527,I1470,I5751,,,I5915,);
not I_293(I5932,I5915);
nand I_294(I5731,I5915,I5881);
DFFARX1 I_295(I5915,I1470,I5751,,,I5963,);
and I_296(I5716,I5802,I5963);
nand I_297(I5994,I4512,I4506);
and I_298(I6011,I5994,I4521);
DFFARX1 I_299(I6011,I1470,I5751,,,I6028,);
nor I_300(I6045,I6028,I5932);
and I_301(I6062,I5864,I6045);
nor I_302(I6079,I6028,I5802);
DFFARX1 I_303(I6028,I1470,I5751,,,I5722,);
DFFARX1 I_304(I4509,I1470,I5751,,,I6110,);
and I_305(I6127,I6110,I4533);
or I_306(I6144,I6127,I6062);
DFFARX1 I_307(I6144,I1470,I5751,,,I5734,);
nand I_308(I5743,I6127,I6079);
DFFARX1 I_309(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_310(I4518,I1470,I5751,,,I6203,);
nand I_311(I5737,I6203,I5898);
DFFARX1 I_312(I6203,I1470,I5751,,,I5725,);
nand I_313(I6248,I6203,I5864);
and I_314(I6265,I5915,I6248);
DFFARX1 I_315(I6265,I1470,I5751,,,I5719,);
not I_316(I6329,I1477);
nand I_317(I6346,I3969,I3954);
and I_318(I6363,I6346,I3963);
DFFARX1 I_319(I6363,I1470,I6329,,,I6380,);
not I_320(I6318,I6380);
DFFARX1 I_321(I6380,I1470,I6329,,,I6411,);
not I_322(I6306,I6411);
nor I_323(I6442,I3975,I3954);
not I_324(I6459,I6442);
nor I_325(I6476,I6380,I6459);
DFFARX1 I_326(I3966,I1470,I6329,,,I6493,);
not I_327(I6510,I6493);
nand I_328(I6309,I6493,I6459);
DFFARX1 I_329(I6493,I1470,I6329,,,I6541,);
and I_330(I6294,I6380,I6541);
nand I_331(I6572,I3951,I3945);
and I_332(I6589,I6572,I3960);
DFFARX1 I_333(I6589,I1470,I6329,,,I6606,);
nor I_334(I6623,I6606,I6510);
and I_335(I6640,I6442,I6623);
nor I_336(I6657,I6606,I6380);
DFFARX1 I_337(I6606,I1470,I6329,,,I6300,);
DFFARX1 I_338(I3948,I1470,I6329,,,I6688,);
and I_339(I6705,I6688,I3972);
or I_340(I6722,I6705,I6640);
DFFARX1 I_341(I6722,I1470,I6329,,,I6312,);
nand I_342(I6321,I6705,I6657);
DFFARX1 I_343(I6705,I1470,I6329,,,I6291,);
DFFARX1 I_344(I3957,I1470,I6329,,,I6781,);
nand I_345(I6315,I6781,I6476);
DFFARX1 I_346(I6781,I1470,I6329,,,I6303,);
nand I_347(I6826,I6781,I6442);
and I_348(I6843,I6493,I6826);
DFFARX1 I_349(I6843,I1470,I6329,,,I6297,);
not I_350(I6907,I1477);
not I_351(I6924,I5073);
nor I_352(I6941,I5070,I5094);
nand I_353(I6958,I6941,I5091);
nor I_354(I6975,I6924,I5070);
nand I_355(I6992,I6975,I5097);
not I_356(I7009,I6992);
not I_357(I7026,I5070);
nor I_358(I6896,I6992,I7026);
not I_359(I7057,I7026);
nand I_360(I6881,I6992,I7057);
not I_361(I7088,I5088);
nor I_362(I7105,I7088,I5079);
and I_363(I7122,I7105,I5076);
or I_364(I7139,I7122,I5085);
DFFARX1 I_365(I7139,I1470,I6907,,,I7156,);
nor I_366(I7173,I7156,I7009);
DFFARX1 I_367(I7156,I1470,I6907,,,I7190,);
not I_368(I6878,I7190);
nand I_369(I7221,I6924,I5088);
and I_370(I7238,I7221,I7173);
DFFARX1 I_371(I7221,I1470,I6907,,,I6875,);
DFFARX1 I_372(I5067,I1470,I6907,,,I7269,);
nor I_373(I7286,I7269,I6992);
nand I_374(I6893,I7156,I7286);
nor I_375(I7317,I7269,I7057);
not I_376(I6890,I7269);
nand I_377(I7348,I7269,I6958);
and I_378(I7365,I7026,I7348);
DFFARX1 I_379(I7365,I1470,I6907,,,I6869,);
DFFARX1 I_380(I7269,I1470,I6907,,,I6872,);
DFFARX1 I_381(I5082,I1470,I6907,,,I7410,);
not I_382(I7427,I7410);
nand I_383(I7444,I7427,I6992);
and I_384(I7461,I7221,I7444);
DFFARX1 I_385(I7461,I1470,I6907,,,I6899,);
or I_386(I7492,I7427,I7238);
DFFARX1 I_387(I7492,I1470,I6907,,,I6884,);
nand I_388(I6887,I7427,I7317);
not I_389(I7570,I1477);
not I_390(I7587,I6300);
nor I_391(I7604,I6297,I6294);
nand I_392(I7621,I7604,I6315);
DFFARX1 I_393(I7621,I1470,I7570,,,I7544,);
nor I_394(I7652,I7587,I6297);
nand I_395(I7669,I7652,I6318);
not I_396(I7559,I7669);
DFFARX1 I_397(I7669,I1470,I7570,,,I7541,);
not I_398(I7714,I6297);
not I_399(I7731,I7714);
not I_400(I7748,I6291);
nor I_401(I7765,I7748,I6303);
and I_402(I7782,I7765,I6312);
or I_403(I7799,I7782,I6306);
DFFARX1 I_404(I7799,I1470,I7570,,,I7816,);
nor I_405(I7833,I7816,I7669);
nor I_406(I7850,I7816,I7731);
nand I_407(I7556,I7621,I7850);
nand I_408(I7881,I7587,I6291);
nand I_409(I7898,I7881,I7816);
and I_410(I7915,I7881,I7898);
DFFARX1 I_411(I7915,I1470,I7570,,,I7538,);
DFFARX1 I_412(I7881,I1470,I7570,,,I7946,);
and I_413(I7535,I7714,I7946);
DFFARX1 I_414(I6321,I1470,I7570,,,I7977,);
not I_415(I7994,I7977);
nor I_416(I8011,I7669,I7994);
and I_417(I8028,I7977,I8011);
nand I_418(I7550,I7977,I7731);
DFFARX1 I_419(I7977,I1470,I7570,,,I8059,);
not I_420(I7547,I8059);
DFFARX1 I_421(I6309,I1470,I7570,,,I8090,);
not I_422(I8107,I8090);
or I_423(I8124,I8107,I8028);
DFFARX1 I_424(I8124,I1470,I7570,,,I7553,);
nand I_425(I7562,I8107,I7833);
DFFARX1 I_426(I8107,I1470,I7570,,,I7532,);
not I_427(I8216,I1477);
not I_428(I8233,I5722);
nor I_429(I8250,I5719,I5716);
nand I_430(I8267,I8250,I5737);
DFFARX1 I_431(I8267,I1470,I8216,,,I8190,);
nor I_432(I8298,I8233,I5719);
nand I_433(I8315,I8298,I5740);
not I_434(I8205,I8315);
DFFARX1 I_435(I8315,I1470,I8216,,,I8187,);
not I_436(I8360,I5719);
not I_437(I8377,I8360);
not I_438(I8394,I5713);
nor I_439(I8411,I8394,I5725);
and I_440(I8428,I8411,I5734);
or I_441(I8445,I8428,I5728);
DFFARX1 I_442(I8445,I1470,I8216,,,I8462,);
nor I_443(I8479,I8462,I8315);
nor I_444(I8496,I8462,I8377);
nand I_445(I8202,I8267,I8496);
nand I_446(I8527,I8233,I5713);
nand I_447(I8544,I8527,I8462);
and I_448(I8561,I8527,I8544);
DFFARX1 I_449(I8561,I1470,I8216,,,I8184,);
DFFARX1 I_450(I8527,I1470,I8216,,,I8592,);
and I_451(I8181,I8360,I8592);
DFFARX1 I_452(I5743,I1470,I8216,,,I8623,);
not I_453(I8640,I8623);
nor I_454(I8657,I8315,I8640);
and I_455(I8674,I8623,I8657);
nand I_456(I8196,I8623,I8377);
DFFARX1 I_457(I8623,I1470,I8216,,,I8705,);
not I_458(I8193,I8705);
DFFARX1 I_459(I5731,I1470,I8216,,,I8736,);
not I_460(I8753,I8736);
or I_461(I8770,I8753,I8674);
DFFARX1 I_462(I8770,I1470,I8216,,,I8199,);
nand I_463(I8208,I8753,I8479);
DFFARX1 I_464(I8753,I1470,I8216,,,I8178,);
not I_465(I8862,I1477);
not I_466(I8879,I6887);
nor I_467(I8896,I6893,I6872);
nand I_468(I8913,I8896,I6878);
nor I_469(I8930,I8879,I6893);
nand I_470(I8947,I8930,I6884);
not I_471(I8964,I6893);
not I_472(I8981,I8964);
not I_473(I8998,I6881);
nor I_474(I9015,I8998,I6899);
and I_475(I9032,I9015,I6890);
or I_476(I9049,I9032,I6869);
DFFARX1 I_477(I9049,I1470,I8862,,,I9066,);
nand I_478(I9083,I8879,I6881);
or I_479(I8851,I9083,I9066);
not I_480(I9114,I9083);
nor I_481(I9131,I9066,I9114);
and I_482(I9148,I8964,I9131);
nand I_483(I8824,I9083,I8981);
DFFARX1 I_484(I6896,I1470,I8862,,,I9179,);
or I_485(I8845,I9179,I9066);
nor I_486(I9210,I9179,I8947);
nor I_487(I9227,I9179,I8981);
nand I_488(I8830,I8913,I9227);
or I_489(I9258,I9179,I9148);
DFFARX1 I_490(I9258,I1470,I8862,,,I8827,);
not I_491(I8833,I9179);
DFFARX1 I_492(I6875,I1470,I8862,,,I9303,);
not I_493(I9320,I9303);
nor I_494(I9337,I9320,I8913);
DFFARX1 I_495(I9337,I1470,I8862,,,I8839,);
nor I_496(I8854,I9179,I9320);
nor I_497(I8842,I9320,I9083);
not I_498(I9396,I9320);
and I_499(I9413,I8947,I9396);
nor I_500(I8848,I9083,I9413);
nand I_501(I8836,I9320,I9210);
not I_502(I9491,I1477);
nand I_503(I9508,I8199,I8202);
and I_504(I9525,I9508,I8184);
DFFARX1 I_505(I9525,I1470,I9491,,,I9542,);
not I_506(I9559,I9542);
nor I_507(I9576,I8181,I8202);
or I_508(I9474,I9576,I9542);
not I_509(I9462,I9576);
DFFARX1 I_510(I8205,I1470,I9491,,,I9621,);
nor I_511(I9638,I9621,I9576);
nand I_512(I9655,I8190,I8196);
and I_513(I9672,I9655,I8208);
DFFARX1 I_514(I9672,I1470,I9491,,,I9689,);
nor I_515(I9471,I9689,I9542);
not I_516(I9720,I9689);
nor I_517(I9737,I9621,I9720);
DFFARX1 I_518(I8187,I1470,I9491,,,I9754,);
and I_519(I9771,I9754,I8178);
or I_520(I9480,I9771,I9576);
nand I_521(I9459,I9771,I9737);
DFFARX1 I_522(I8193,I1470,I9491,,,I9816,);
and I_523(I9833,I9816,I9559);
nor I_524(I9477,I9771,I9833);
nor I_525(I9864,I9816,I9621);
DFFARX1 I_526(I9864,I1470,I9491,,,I9468,);
nor I_527(I9483,I9816,I9542);
not I_528(I9909,I9816);
nor I_529(I9926,I9689,I9909);
and I_530(I9943,I9576,I9926);
or I_531(I9960,I9771,I9943);
DFFARX1 I_532(I9960,I1470,I9491,,,I9456,);
nand I_533(I9465,I9816,I9638);
nand I_534(I9453,I9816,I9720);
not I_535(I10052,I1477);
nand I_536(I10069,I7559,I7535);
and I_537(I10086,I10069,I7544);
DFFARX1 I_538(I10086,I1470,I10052,,,I10103,);
nor I_539(I10120,I7538,I7535);
DFFARX1 I_540(I7553,I1470,I10052,,,I10137,);
nand I_541(I10154,I10137,I10120);
DFFARX1 I_542(I10137,I1470,I10052,,,I10023,);
nand I_543(I10185,I7547,I7562);
and I_544(I10202,I10185,I7541);
DFFARX1 I_545(I10202,I1470,I10052,,,I10219,);
not I_546(I10236,I10219);
nor I_547(I10253,I10103,I10236);
and I_548(I10270,I10120,I10253);
and I_549(I10287,I10219,I10154);
DFFARX1 I_550(I10287,I1470,I10052,,,I10020,);
DFFARX1 I_551(I10219,I1470,I10052,,,I10014,);
DFFARX1 I_552(I7532,I1470,I10052,,,I10332,);
and I_553(I10349,I10332,I7550);
nand I_554(I10366,I10349,I10219);
nor I_555(I10041,I10349,I10120);
not I_556(I10397,I10349);
nor I_557(I10414,I10103,I10397);
nand I_558(I10032,I10137,I10414);
nand I_559(I10026,I10219,I10397);
or I_560(I10459,I10349,I10270);
DFFARX1 I_561(I10459,I1470,I10052,,,I10029,);
DFFARX1 I_562(I7556,I1470,I10052,,,I10490,);
and I_563(I10507,I10490,I10366);
DFFARX1 I_564(I10507,I1470,I10052,,,I10044,);
nor I_565(I10538,I10490,I10103);
nand I_566(I10038,I10349,I10538);
not I_567(I10035,I10490);
DFFARX1 I_568(I10490,I1470,I10052,,,I10583,);
and I_569(I10017,I10490,I10583);
not I_570(I10647,I1477);
not I_571(I10664,I9471);
nor I_572(I10681,I9477,I9480);
nand I_573(I10698,I10681,I9456);
nor I_574(I10715,I10664,I9477);
nand I_575(I10732,I10715,I9465);
not I_576(I10749,I10732);
not I_577(I10766,I9477);
nor I_578(I10636,I10732,I10766);
not I_579(I10797,I10766);
nand I_580(I10621,I10732,I10797);
not I_581(I10828,I9459);
nor I_582(I10845,I10828,I9483);
and I_583(I10862,I10845,I9453);
or I_584(I10879,I10862,I9462);
DFFARX1 I_585(I10879,I1470,I10647,,,I10896,);
nor I_586(I10913,I10896,I10749);
DFFARX1 I_587(I10896,I1470,I10647,,,I10930,);
not I_588(I10618,I10930);
nand I_589(I10961,I10664,I9459);
and I_590(I10978,I10961,I10913);
DFFARX1 I_591(I10961,I1470,I10647,,,I10615,);
DFFARX1 I_592(I9468,I1470,I10647,,,I11009,);
nor I_593(I11026,I11009,I10732);
nand I_594(I10633,I10896,I11026);
nor I_595(I11057,I11009,I10797);
not I_596(I10630,I11009);
nand I_597(I11088,I11009,I10698);
and I_598(I11105,I10766,I11088);
DFFARX1 I_599(I11105,I1470,I10647,,,I10609,);
DFFARX1 I_600(I11009,I1470,I10647,,,I10612,);
DFFARX1 I_601(I9474,I1470,I10647,,,I11150,);
not I_602(I11167,I11150);
nand I_603(I11184,I11167,I10732);
and I_604(I11201,I10961,I11184);
DFFARX1 I_605(I11201,I1470,I10647,,,I10639,);
or I_606(I11232,I11167,I10978);
DFFARX1 I_607(I11232,I1470,I10647,,,I10624,);
nand I_608(I10627,I11167,I11057);
not I_609(I11310,I1477);
not I_610(I11327,I8830);
nor I_611(I11344,I8848,I8839);
nand I_612(I11361,I11344,I8845);
nor I_613(I11378,I11327,I8848);
nand I_614(I11395,I11378,I8851);
not I_615(I11412,I11395);
not I_616(I11429,I8848);
nor I_617(I11299,I11395,I11429);
not I_618(I11460,I11429);
nand I_619(I11284,I11395,I11460);
not I_620(I11491,I8827);
nor I_621(I11508,I11491,I8842);
and I_622(I11525,I11508,I8824);
or I_623(I11542,I11525,I8833);
DFFARX1 I_624(I11542,I1470,I11310,,,I11559,);
nor I_625(I11576,I11559,I11412);
DFFARX1 I_626(I11559,I1470,I11310,,,I11593,);
not I_627(I11281,I11593);
nand I_628(I11624,I11327,I8827);
and I_629(I11641,I11624,I11576);
DFFARX1 I_630(I11624,I1470,I11310,,,I11278,);
DFFARX1 I_631(I8836,I1470,I11310,,,I11672,);
nor I_632(I11689,I11672,I11395);
nand I_633(I11296,I11559,I11689);
nor I_634(I11720,I11672,I11460);
not I_635(I11293,I11672);
nand I_636(I11751,I11672,I11361);
and I_637(I11768,I11429,I11751);
DFFARX1 I_638(I11768,I1470,I11310,,,I11272,);
DFFARX1 I_639(I11672,I1470,I11310,,,I11275,);
DFFARX1 I_640(I8854,I1470,I11310,,,I11813,);
not I_641(I11830,I11813);
nand I_642(I11847,I11830,I11395);
and I_643(I11864,I11624,I11847);
DFFARX1 I_644(I11864,I1470,I11310,,,I11302,);
or I_645(I11895,I11830,I11641);
DFFARX1 I_646(I11895,I1470,I11310,,,I11287,);
nand I_647(I11290,I11830,I11720);
not I_648(I11973,I1477);
not I_649(I11990,I10032);
nor I_650(I12007,I10020,I10029);
nand I_651(I12024,I12007,I10044);
nor I_652(I12041,I11990,I10020);
nand I_653(I12058,I12041,I10026);
DFFARX1 I_654(I12058,I1470,I11973,,,I12075,);
not I_655(I11944,I12075);
not I_656(I12106,I10020);
not I_657(I12123,I12106);
not I_658(I12140,I10014);
nor I_659(I12157,I12140,I10035);
and I_660(I12174,I12157,I10017);
or I_661(I12191,I12174,I10023);
DFFARX1 I_662(I12191,I1470,I11973,,,I12208,);
DFFARX1 I_663(I12208,I1470,I11973,,,I11941,);
DFFARX1 I_664(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_665(I12208,I1470,I11973,,,I11935,);
nand I_666(I12270,I11990,I10014);
nand I_667(I12287,I12270,I12024);
and I_668(I12304,I12106,I12287);
DFFARX1 I_669(I12304,I1470,I11973,,,I11965,);
and I_670(I11938,I12270,I12239);
DFFARX1 I_671(I10041,I1470,I11973,,,I12349,);
nor I_672(I11962,I12349,I12270);
nor I_673(I12380,I12349,I12024);
nand I_674(I11959,I12058,I12380);
not I_675(I11956,I12349);
DFFARX1 I_676(I10038,I1470,I11973,,,I12425,);
not I_677(I12442,I12425);
nor I_678(I12459,I12442,I12123);
and I_679(I12476,I12349,I12459);
or I_680(I12493,I12270,I12476);
DFFARX1 I_681(I12493,I1470,I11973,,,I11950,);
not I_682(I12524,I12442);
nor I_683(I12541,I12349,I12524);
nand I_684(I11953,I12442,I12541);
nand I_685(I11947,I12106,I12524);
not I_686(I12619,I1477);
nand I_687(I12636,I10612,I10639);
and I_688(I12653,I12636,I10627);
DFFARX1 I_689(I12653,I1470,I12619,,,I12670,);
not I_690(I12687,I12670);
DFFARX1 I_691(I12670,I1470,I12619,,,I12587,);
nor I_692(I12718,I10615,I10639);
DFFARX1 I_693(I10630,I1470,I12619,,,I12735,);
DFFARX1 I_694(I12735,I1470,I12619,,,I12752,);
not I_695(I12590,I12752);
DFFARX1 I_696(I12735,I1470,I12619,,,I12783,);
and I_697(I12584,I12670,I12783);
nand I_698(I12814,I10624,I10621);
and I_699(I12831,I12814,I10618);
DFFARX1 I_700(I12831,I1470,I12619,,,I12848,);
nor I_701(I12865,I12848,I12687);
not I_702(I12882,I12848);
nand I_703(I12593,I12670,I12882);
DFFARX1 I_704(I10633,I1470,I12619,,,I12913,);
and I_705(I12930,I12913,I10609);
nor I_706(I12947,I12930,I12848);
nor I_707(I12964,I12930,I12882);
nand I_708(I12599,I12718,I12964);
not I_709(I12602,I12930);
DFFARX1 I_710(I12930,I1470,I12619,,,I12581,);
DFFARX1 I_711(I10636,I1470,I12619,,,I13023,);
nand I_712(I13040,I13023,I12735);
and I_713(I13057,I12718,I13040);
DFFARX1 I_714(I13057,I1470,I12619,,,I12611,);
nor I_715(I12608,I13023,I12930);
and I_716(I13102,I13023,I12865);
or I_717(I13119,I12718,I13102);
DFFARX1 I_718(I13119,I1470,I12619,,,I12596,);
nand I_719(I12605,I13023,I12947);
not I_720(I13197,I1477);
nand I_721(I13214,I11275,I11302);
and I_722(I13231,I13214,I11290);
DFFARX1 I_723(I13231,I1470,I13197,,,I13248,);
not I_724(I13265,I13248);
DFFARX1 I_725(I13248,I1470,I13197,,,I13165,);
nor I_726(I13296,I11278,I11302);
DFFARX1 I_727(I11293,I1470,I13197,,,I13313,);
DFFARX1 I_728(I13313,I1470,I13197,,,I13330,);
not I_729(I13168,I13330);
DFFARX1 I_730(I13313,I1470,I13197,,,I13361,);
and I_731(I13162,I13248,I13361);
nand I_732(I13392,I11287,I11284);
and I_733(I13409,I13392,I11281);
DFFARX1 I_734(I13409,I1470,I13197,,,I13426,);
nor I_735(I13443,I13426,I13265);
not I_736(I13460,I13426);
nand I_737(I13171,I13248,I13460);
DFFARX1 I_738(I11296,I1470,I13197,,,I13491,);
and I_739(I13508,I13491,I11272);
nor I_740(I13525,I13508,I13426);
nor I_741(I13542,I13508,I13460);
nand I_742(I13177,I13296,I13542);
not I_743(I13180,I13508);
DFFARX1 I_744(I13508,I1470,I13197,,,I13159,);
DFFARX1 I_745(I11299,I1470,I13197,,,I13601,);
nand I_746(I13618,I13601,I13313);
and I_747(I13635,I13296,I13618);
DFFARX1 I_748(I13635,I1470,I13197,,,I13189,);
nor I_749(I13186,I13601,I13508);
and I_750(I13680,I13601,I13443);
or I_751(I13697,I13296,I13680);
DFFARX1 I_752(I13697,I1470,I13197,,,I13174,);
nand I_753(I13183,I13601,I13525);
not I_754(I13775,I1477);
nand I_755(I13792,I11953,I11965);
and I_756(I13809,I13792,I11947);
DFFARX1 I_757(I13809,I1470,I13775,,,I13826,);
nor I_758(I13843,I11959,I11965);
nor I_759(I13860,I13843,I13826);
not I_760(I13758,I13843);
DFFARX1 I_761(I11944,I1470,I13775,,,I13891,);
not I_762(I13908,I13891);
nor I_763(I13925,I13843,I13908);
nand I_764(I13761,I13891,I13860);
DFFARX1 I_765(I13891,I1470,I13775,,,I13743,);
nand I_766(I13970,I11935,I11950);
and I_767(I13987,I13970,I11941);
DFFARX1 I_768(I13987,I1470,I13775,,,I14004,);
nor I_769(I13764,I14004,I13826);
nand I_770(I13755,I14004,I13925);
DFFARX1 I_771(I11962,I1470,I13775,,,I14049,);
and I_772(I14066,I14049,I11956);
DFFARX1 I_773(I14066,I1470,I13775,,,I14083,);
not I_774(I13746,I14083);
nand I_775(I14114,I14066,I14004);
and I_776(I14131,I13826,I14114);
DFFARX1 I_777(I14131,I1470,I13775,,,I13737,);
DFFARX1 I_778(I11938,I1470,I13775,,,I14162,);
nand I_779(I14179,I14162,I13826);
and I_780(I14196,I14004,I14179);
DFFARX1 I_781(I14196,I1470,I13775,,,I13767,);
not I_782(I14227,I14162);
nor I_783(I14244,I13843,I14227);
and I_784(I14261,I14162,I14244);
or I_785(I14278,I14066,I14261);
DFFARX1 I_786(I14278,I1470,I13775,,,I13752,);
nand I_787(I13749,I14162,I13908);
DFFARX1 I_788(I14162,I1470,I13775,,,I13740,);
not I_789(I14370,I1477);
nand I_790(I14387,I13171,I13186);
and I_791(I14404,I14387,I13183);
DFFARX1 I_792(I14404,I1470,I14370,,,I14421,);
nor I_793(I14438,I13159,I13186);
DFFARX1 I_794(I13177,I1470,I14370,,,I14455,);
nand I_795(I14472,I14455,I14438);
DFFARX1 I_796(I14455,I1470,I14370,,,I14341,);
nand I_797(I14503,I13180,I13168);
and I_798(I14520,I14503,I13174);
DFFARX1 I_799(I14520,I1470,I14370,,,I14537,);
not I_800(I14554,I14537);
nor I_801(I14571,I14421,I14554);
and I_802(I14588,I14438,I14571);
and I_803(I14605,I14537,I14472);
DFFARX1 I_804(I14605,I1470,I14370,,,I14338,);
DFFARX1 I_805(I14537,I1470,I14370,,,I14332,);
DFFARX1 I_806(I13165,I1470,I14370,,,I14650,);
and I_807(I14667,I14650,I13189);
nand I_808(I14684,I14667,I14537);
nor I_809(I14359,I14667,I14438);
not I_810(I14715,I14667);
nor I_811(I14732,I14421,I14715);
nand I_812(I14350,I14455,I14732);
nand I_813(I14344,I14537,I14715);
or I_814(I14777,I14667,I14588);
DFFARX1 I_815(I14777,I1470,I14370,,,I14347,);
DFFARX1 I_816(I13162,I1470,I14370,,,I14808,);
and I_817(I14825,I14808,I14684);
DFFARX1 I_818(I14825,I1470,I14370,,,I14362,);
nor I_819(I14856,I14808,I14421);
nand I_820(I14356,I14667,I14856);
not I_821(I14353,I14808);
DFFARX1 I_822(I14808,I1470,I14370,,,I14901,);
and I_823(I14335,I14808,I14901);
not I_824(I14965,I1477);
not I_825(I14982,I12596);
nor I_826(I14999,I12584,I12590);
nand I_827(I15016,I14999,I12581);
DFFARX1 I_828(I15016,I1470,I14965,,,I14939,);
nor I_829(I15047,I14982,I12584);
nand I_830(I15064,I15047,I12587);
not I_831(I14954,I15064);
DFFARX1 I_832(I15064,I1470,I14965,,,I14936,);
not I_833(I15109,I12584);
not I_834(I15126,I15109);
not I_835(I15143,I12599);
nor I_836(I15160,I15143,I12611);
and I_837(I15177,I15160,I12593);
or I_838(I15194,I15177,I12608);
DFFARX1 I_839(I15194,I1470,I14965,,,I15211,);
nor I_840(I15228,I15211,I15064);
nor I_841(I15245,I15211,I15126);
nand I_842(I14951,I15016,I15245);
nand I_843(I15276,I14982,I12599);
nand I_844(I15293,I15276,I15211);
and I_845(I15310,I15276,I15293);
DFFARX1 I_846(I15310,I1470,I14965,,,I14933,);
DFFARX1 I_847(I15276,I1470,I14965,,,I15341,);
and I_848(I14930,I15109,I15341);
DFFARX1 I_849(I12602,I1470,I14965,,,I15372,);
not I_850(I15389,I15372);
nor I_851(I15406,I15064,I15389);
and I_852(I15423,I15372,I15406);
nand I_853(I14945,I15372,I15126);
DFFARX1 I_854(I15372,I1470,I14965,,,I15454,);
not I_855(I14942,I15454);
DFFARX1 I_856(I12605,I1470,I14965,,,I15485,);
not I_857(I15502,I15485);
or I_858(I15519,I15502,I15423);
DFFARX1 I_859(I15519,I1470,I14965,,,I14948,);
nand I_860(I14957,I15502,I15228);
DFFARX1 I_861(I15502,I1470,I14965,,,I14927,);
not I_862(I15611,I1477);
not I_863(I15628,I13743);
nor I_864(I15645,I13761,I13740);
nand I_865(I15662,I15645,I13764);
nor I_866(I15679,I15628,I13761);
nand I_867(I15696,I15679,I13758);
not I_868(I15713,I13761);
not I_869(I15730,I15713);
not I_870(I15747,I13749);
nor I_871(I15764,I15747,I13737);
and I_872(I15781,I15764,I13755);
or I_873(I15798,I15781,I13767);
DFFARX1 I_874(I15798,I1470,I15611,,,I15815,);
nand I_875(I15832,I15628,I13749);
or I_876(I15600,I15832,I15815);
not I_877(I15863,I15832);
nor I_878(I15880,I15815,I15863);
and I_879(I15897,I15713,I15880);
nand I_880(I15573,I15832,I15730);
DFFARX1 I_881(I13746,I1470,I15611,,,I15928,);
or I_882(I15594,I15928,I15815);
nor I_883(I15959,I15928,I15696);
nor I_884(I15976,I15928,I15730);
nand I_885(I15579,I15662,I15976);
or I_886(I16007,I15928,I15897);
DFFARX1 I_887(I16007,I1470,I15611,,,I15576,);
not I_888(I15582,I15928);
DFFARX1 I_889(I13752,I1470,I15611,,,I16052,);
not I_890(I16069,I16052);
nor I_891(I16086,I16069,I15662);
DFFARX1 I_892(I16086,I1470,I15611,,,I15588,);
nor I_893(I15603,I15928,I16069);
nor I_894(I15591,I16069,I15832);
not I_895(I16145,I16069);
and I_896(I16162,I15696,I16145);
nor I_897(I15597,I15832,I16162);
nand I_898(I15585,I16069,I15959);
not I_899(I16240,I1477);
nand I_900(I16257,I14341,I14338);
and I_901(I16274,I16257,I14332);
DFFARX1 I_902(I16274,I1470,I16240,,,I16291,);
not I_903(I16308,I16291);
nor I_904(I16339,I14353,I14338);
DFFARX1 I_905(I14356,I1470,I16240,,,I16356,);
DFFARX1 I_906(I16356,I1470,I16240,,,I16373,);
DFFARX1 I_907(I16356,I1470,I16240,,,I16404,);
nand I_908(I16435,I14359,I14350);
and I_909(I16452,I16435,I14362);
DFFARX1 I_910(I16452,I1470,I16240,,,I16469,);
nor I_911(I16486,I16469,I16308);
not I_912(I16503,I16469);
DFFARX1 I_913(I14335,I1470,I16240,,,I16534,);
and I_914(I16551,I16534,I14344);
nor I_915(I16568,I16551,I16469);
nor I_916(I16585,I16551,I16503);
DFFARX1 I_917(I14347,I1470,I16240,,,I16644,);
nand I_918(I16661,I16644,I16356);
and I_919(I16678,I16339,I16661);
and I_920(I16723,I16644,I16486);
or I_921(I16740,I16339,I16723);
not I_922(I16818,I1477);
nand I_923(I16835,I14936,I14948);
and I_924(I16852,I16835,I14957);
DFFARX1 I_925(I16852,I1470,I16818,,,I16869,);
nor I_926(I16886,I14951,I14948);
nor I_927(I16903,I16886,I16869);
DFFARX1 I_928(I14945,I1470,I16818,,,I16934,);
not I_929(I16951,I16934);
nor I_930(I16968,I16886,I16951);
nand I_931(I17013,I14942,I14939);
and I_932(I17030,I17013,I14930);
DFFARX1 I_933(I17030,I1470,I16818,,,I17047,);
DFFARX1 I_934(I14954,I1470,I16818,,,I17092,);
and I_935(I17109,I17092,I14933);
DFFARX1 I_936(I17109,I1470,I16818,,,I17126,);
nand I_937(I17157,I17109,I17047);
and I_938(I17174,I16869,I17157);
DFFARX1 I_939(I14927,I1470,I16818,,,I17205,);
nand I_940(I17222,I17205,I16869);
and I_941(I17239,I17047,I17222);
not I_942(I17270,I17205);
nor I_943(I17287,I16886,I17270);
and I_944(I17304,I17205,I17287);
or I_945(I17321,I17109,I17304);
not I_946(I17413,I1477);
not I_947(I17430,I15579);
nor I_948(I17447,I15597,I15588);
nand I_949(I17464,I17447,I15594);
nor I_950(I17481,I17430,I15597);
nand I_951(I17498,I17481,I15600);
not I_952(I17515,I17498);
not I_953(I17532,I15597);
not I_954(I17563,I17532);
not I_955(I17594,I15576);
nor I_956(I17611,I17594,I15591);
and I_957(I17628,I17611,I15573);
or I_958(I17645,I17628,I15582);
DFFARX1 I_959(I17645,I1470,I17413,,,I17662,);
nor I_960(I17679,I17662,I17515);
DFFARX1 I_961(I17662,I1470,I17413,,,I17696,);
nand I_962(I17727,I17430,I15576);
and I_963(I17744,I17727,I17679);
DFFARX1 I_964(I15585,I1470,I17413,,,I17775,);
nor I_965(I17792,I17775,I17498);
nor I_966(I17823,I17775,I17563);
nand I_967(I17854,I17775,I17464);
and I_968(I17871,I17532,I17854);
DFFARX1 I_969(I15603,I1470,I17413,,,I17916,);
not I_970(I17933,I17916);
nand I_971(I17950,I17933,I17498);
and I_972(I17967,I17727,I17950);
or I_973(I17998,I17933,I17744);
endmodule


