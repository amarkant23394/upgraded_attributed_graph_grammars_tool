module test_I15579(I1477,I13987,I13809,I1470,I15579);
input I1477,I13987,I13809,I1470;
output I15579;
wire I15645,I14004,I15730,I13860,I13746,I15662,I13891,I14083,I13775,I15611,I15928,I13761,I15713,I13740,I13764,I13826,I14162,I15976;
nor I_0(I15645,I13761,I13740);
DFFARX1 I_1(I13987,I1470,I13775,,,I14004,);
not I_2(I15730,I15713);
nor I_3(I13860,I13826);
not I_4(I13746,I14083);
nand I_5(I15662,I15645,I13764);
DFFARX1 I_6(I1470,I13775,,,I13891,);
DFFARX1 I_7(I1470,I13775,,,I14083,);
nand I_8(I15579,I15662,I15976);
not I_9(I13775,I1477);
not I_10(I15611,I1477);
DFFARX1 I_11(I13746,I1470,I15611,,,I15928,);
nand I_12(I13761,I13891,I13860);
not I_13(I15713,I13761);
DFFARX1 I_14(I14162,I1470,I13775,,,I13740,);
nor I_15(I13764,I14004,I13826);
DFFARX1 I_16(I13809,I1470,I13775,,,I13826,);
DFFARX1 I_17(I1470,I13775,,,I14162,);
nor I_18(I15976,I15928,I15730);
endmodule


