module test_I9754(I8233,I1477,I1470,I9754);
input I8233,I1477,I1470;
output I9754;
wire I8187,I8216,I5802,I8298,I5719,I5740,I8315,I9491;
DFFARX1 I_0(I8315,I1470,I8216,,,I8187,);
not I_1(I8216,I1477);
DFFARX1 I_2(I8187,I1470,I9491,,,I9754,);
DFFARX1 I_3(I1470,,,I5802,);
nor I_4(I8298,I8233,I5719);
DFFARX1 I_5(I1470,,,I5719,);
not I_6(I5740,I5802);
nand I_7(I8315,I8298,I5740);
not I_8(I9491,I1477);
endmodule


