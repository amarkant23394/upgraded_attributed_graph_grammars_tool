module test_final(IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_reset_net_0_r_4,blif_clk_net_0_r_4,ACVQN2_0_r_4,n_266_and_0_0_r_4,ACVQN1_2_r_4,P6_2_r_4,n_429_or_0_3_r_4,G78_3_r_4,n_576_3_r_4,n_102_3_r_4,n_547_3_r_4,n_42_5_r_4,G199_5_r_4);
input IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_reset_net_0_r_4,blif_clk_net_0_r_4;
output ACVQN2_0_r_4,n_266_and_0_0_r_4,ACVQN1_2_r_4,P6_2_r_4,n_429_or_0_3_r_4,G78_3_r_4,n_576_3_r_4,n_102_3_r_4,n_547_3_r_4,n_42_5_r_4,G199_5_r_4;
wire ACVQN2_0_r_8,n_266_and_0_0_r_8,ACVQN1_2_r_8,P6_2_r_8,n_429_or_0_3_r_8,G78_3_r_8,n_576_3_r_8,n_102_3_r_8,n_547_3_r_8,n_42_5_r_8,G199_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8,ACVQN1_0_l_8,N1_1_l_8,G199_1_l_8,G214_1_l_8,n3_1_l_8,n_42_5_l_8,N3_5_l_8,G199_5_l_8,n3_5_l_8,ACVQN1_0_r_8,P6_internal_2_r_8,n12_3_r_8,n_431_3_r_8,n11_3_r_8,n13_3_r_8,n14_3_r_8,n15_3_r_8,n16_3_r_8,N3_5_r_8,n3_5_r_8,n1_0_r_4,ACVQN2_0_l_4,n_266_and_0_0_l_4,ACVQN1_0_l_4,n4_4_l_4,G42_4_l_4,n_87_4_l_4,n_572_4_l_4,n_573_4_l_4,n_549_4_l_4,n7_4_l_4,n_569_4_l_4,n_452_4_l_4,ACVQN1_0_r_4,P6_internal_2_r_4,n12_3_r_4,n_431_3_r_4,n11_3_r_4,n13_3_r_4,n14_3_r_4,n15_3_r_4,n16_3_r_4,N3_5_r_4,n3_5_r_4;
DFFARX1 I_0(n_266_and_0_0_l_8,blif_clk_net_0_r_4,n1_0_r_4,ACVQN2_0_r_8,);
and I_1(n_266_and_0_0_r_8,G199_5_l_8,ACVQN1_0_r_8);
DFFARX1 I_2(G199_5_l_8,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_2_r_8,);
not I_3(P6_2_r_8,P6_internal_2_r_8);
nand I_4(n_429_or_0_3_r_8,G199_5_l_8,n12_3_r_8);
DFFARX1 I_5(n_431_3_r_8,blif_clk_net_0_r_4,n1_0_r_4,G78_3_r_8,);
nand I_6(n_576_3_r_8,n_42_5_l_8,n11_3_r_8);
not I_7(n_102_3_r_8,n_266_and_0_0_l_8);
nand I_8(n_547_3_r_8,ACVQN2_0_l_8,n13_3_r_8);
nor I_9(n_42_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8);
DFFARX1 I_10(N3_5_r_8,blif_clk_net_0_r_4,n1_0_r_4,G199_5_r_8,);
DFFARX1 I_11(IN_1_0_l_8,blif_clk_net_0_r_4,n1_0_r_4,ACVQN2_0_l_8,);
and I_12(n_266_and_0_0_l_8,IN_4_0_l_8,ACVQN1_0_l_8);
DFFARX1 I_13(IN_2_0_l_8,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_0_l_8,);
and I_14(N1_1_l_8,IN_6_1_l_8,n3_1_l_8);
DFFARX1 I_15(N1_1_l_8,blif_clk_net_0_r_4,n1_0_r_4,G199_1_l_8,);
DFFARX1 I_16(IN_3_1_l_8,blif_clk_net_0_r_4,n1_0_r_4,G214_1_l_8,);
nand I_17(n3_1_l_8,IN_1_1_l_8,IN_2_1_l_8);
nor I_18(n_42_5_l_8,IN_1_5_l_8,IN_3_5_l_8);
and I_19(N3_5_l_8,IN_6_5_l_8,n3_5_l_8);
DFFARX1 I_20(N3_5_l_8,blif_clk_net_0_r_4,n1_0_r_4,G199_5_l_8,);
nand I_21(n3_5_l_8,IN_2_5_l_8,IN_3_5_l_8);
DFFARX1 I_22(G214_1_l_8,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_0_r_8,);
DFFARX1 I_23(G214_1_l_8,blif_clk_net_0_r_4,n1_0_r_4,P6_internal_2_r_8,);
not I_24(n12_3_r_8,G199_1_l_8);
or I_25(n_431_3_r_8,n_42_5_l_8,n14_3_r_8);
nor I_26(n11_3_r_8,n_266_and_0_0_l_8,n12_3_r_8);
nor I_27(n13_3_r_8,n_266_and_0_0_l_8,G199_1_l_8);
and I_28(n14_3_r_8,ACVQN2_0_l_8,n15_3_r_8);
nor I_29(n15_3_r_8,G199_1_l_8,n16_3_r_8);
not I_30(n16_3_r_8,G199_5_l_8);
and I_31(N3_5_r_8,n_42_5_l_8,n3_5_r_8);
nand I_32(n3_5_r_8,ACVQN2_0_l_8,G214_1_l_8);
DFFARX1 I_33(n_569_4_l_4,blif_clk_net_0_r_4,n1_0_r_4,ACVQN2_0_r_4,);
and I_34(n_266_and_0_0_r_4,ACVQN2_0_l_4,ACVQN1_0_r_4);
DFFARX1 I_35(n_266_and_0_0_l_4,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_2_r_4,);
not I_36(P6_2_r_4,P6_internal_2_r_4);
nand I_37(n_429_or_0_3_r_4,G42_4_l_4,n12_3_r_4);
DFFARX1 I_38(n_431_3_r_4,blif_clk_net_0_r_4,n1_0_r_4,G78_3_r_4,);
nand I_39(n_576_3_r_4,n_573_4_l_4,n11_3_r_4);
not I_40(n_102_3_r_4,n_569_4_l_4);
nand I_41(n_547_3_r_4,ACVQN2_0_l_4,n13_3_r_4);
nor I_42(n_42_5_r_4,G42_4_l_4,n_549_4_l_4);
DFFARX1 I_43(N3_5_r_4,blif_clk_net_0_r_4,n1_0_r_4,G199_5_r_4,);
not I_44(n1_0_r_4,blif_reset_net_0_r_4);
DFFARX1 I_45(n_266_and_0_0_r_8,blif_clk_net_0_r_4,n1_0_r_4,ACVQN2_0_l_4,);
and I_46(n_266_and_0_0_l_4,ACVQN1_0_l_4,n_576_3_r_8);
DFFARX1 I_47(n_42_5_r_8,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_0_l_4,);
nor I_48(n4_4_l_4,ACVQN1_2_r_8,n_547_3_r_8);
DFFARX1 I_49(n4_4_l_4,blif_clk_net_0_r_4,n1_0_r_4,G42_4_l_4,);
not I_50(n_87_4_l_4,G78_3_r_8);
nor I_51(n_572_4_l_4,n_429_or_0_3_r_8,G78_3_r_8);
or I_52(n_573_4_l_4,ACVQN2_0_r_8,P6_2_r_8);
nor I_53(n_549_4_l_4,n7_4_l_4,G199_5_r_8);
and I_54(n7_4_l_4,n_87_4_l_4,n_102_3_r_8);
or I_55(n_569_4_l_4,ACVQN2_0_r_8,G199_5_r_8);
nor I_56(n_452_4_l_4,ACVQN1_2_r_8,P6_2_r_8);
DFFARX1 I_57(n_549_4_l_4,blif_clk_net_0_r_4,n1_0_r_4,ACVQN1_0_r_4,);
DFFARX1 I_58(ACVQN2_0_l_4,blif_clk_net_0_r_4,n1_0_r_4,P6_internal_2_r_4,);
not I_59(n12_3_r_4,n_266_and_0_0_l_4);
or I_60(n_431_3_r_4,n_572_4_l_4,n14_3_r_4);
nor I_61(n11_3_r_4,n_569_4_l_4,n12_3_r_4);
nor I_62(n13_3_r_4,n_572_4_l_4,n_569_4_l_4);
and I_63(n14_3_r_4,n_452_4_l_4,n15_3_r_4);
nor I_64(n15_3_r_4,n_266_and_0_0_l_4,n16_3_r_4);
not I_65(n16_3_r_4,G42_4_l_4);
and I_66(N3_5_r_4,n_573_4_l_4,n3_5_r_4);
nand I_67(n3_5_r_4,n_549_4_l_4,n_452_4_l_4);
endmodule


