module Benchmark_testing10000(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2703,I2711,I2719,I2727,I2735,I2743,I2751,I2759,I2767,I2775,I2783,I2791,I2799,I2807,I2815,I2823,I2831,I2839,I2847,I2855,I2863,I2871,I2879,I2887,I2895,I2903,I2911,I2919,I2927,I2935,I2943,I2951,I2959,I2966,I2973,I114083,I114077,I114074,I114086,I114071,I114092,I114101,I114095,I114098,I114089,I114080,I115883,I115868,I115865,I115862,I115880,I115877,I115856,I115859,I115886,I115871,I115874,I117209,I117194,I117191,I117188,I117206,I117203,I117182,I117185,I117212,I117197,I117200,I121013,I121016,I121010,I121019,I121025,I121028,I121007,I121037,I121034,I121022,I121031,I121591,I121594,I121588,I121597,I121603,I121606,I121585,I121615,I121612,I121600,I121609,I122768,I122753,I122750,I122762,I122756,I122771,I122741,I122759,I122765,I122744,I122747,I129273,I129261,I129270,I129279,I129258,I129276,I129267,I129282,I129255,I129264,I129252,I132916,I132931,I132928,I132913,I132910,I132937,I132925,I132919,I132934,I132922,I132907,I134177,I134171,I134168,I134180,I134165,I134186,I134195,I134189,I134192,I134183,I134174,I134787,I134772,I134769,I134766,I134784,I134781,I134760,I134763,I134790,I134775,I134778,I141853,I141856,I141838,I141859,I141850,I141841,I141832,I141862,I141847,I141844,I141835,I142436,I142433,I142427,I142454,I142445,I142439,I142442,I142457,I142451,I142448,I142430,I143621,I143609,I143618,I143627,I143606,I143624,I143615,I143630,I143603,I143612,I143600,I145295,I145310,I145292,I145307,I145289,I145286,I145301,I145298,I145304,I145313,I145283,I145941,I145956,I145938,I145953,I145935,I145932,I145947,I145944,I145950,I145959,I145929,I146587,I146581,I146578,I146590,I146575,I146596,I146605,I146599,I146602,I146593,I146584,I149084,I149057,I149078,I149063,I149060,I149066,I149072,I149087,I149075,I149081,I149069,I149713,I149701,I149704,I149689,I149695,I149707,I149716,I149686,I149710,I149698,I149692,I150285,I150273,I150282,I150291,I150270,I150288,I150279,I150294,I150267,I150276,I150264,I150852,I150837,I150834,I150831,I150849,I150846,I150825,I150828,I150855,I150840,I150843);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2703,I2711,I2719,I2727,I2735,I2743,I2751,I2759,I2767,I2775,I2783,I2791,I2799,I2807,I2815,I2823,I2831,I2839,I2847,I2855,I2863,I2871,I2879,I2887,I2895,I2903,I2911,I2919,I2927,I2935,I2943,I2951,I2959,I2966,I2973;
output I114083,I114077,I114074,I114086,I114071,I114092,I114101,I114095,I114098,I114089,I114080,I115883,I115868,I115865,I115862,I115880,I115877,I115856,I115859,I115886,I115871,I115874,I117209,I117194,I117191,I117188,I117206,I117203,I117182,I117185,I117212,I117197,I117200,I121013,I121016,I121010,I121019,I121025,I121028,I121007,I121037,I121034,I121022,I121031,I121591,I121594,I121588,I121597,I121603,I121606,I121585,I121615,I121612,I121600,I121609,I122768,I122753,I122750,I122762,I122756,I122771,I122741,I122759,I122765,I122744,I122747,I129273,I129261,I129270,I129279,I129258,I129276,I129267,I129282,I129255,I129264,I129252,I132916,I132931,I132928,I132913,I132910,I132937,I132925,I132919,I132934,I132922,I132907,I134177,I134171,I134168,I134180,I134165,I134186,I134195,I134189,I134192,I134183,I134174,I134787,I134772,I134769,I134766,I134784,I134781,I134760,I134763,I134790,I134775,I134778,I141853,I141856,I141838,I141859,I141850,I141841,I141832,I141862,I141847,I141844,I141835,I142436,I142433,I142427,I142454,I142445,I142439,I142442,I142457,I142451,I142448,I142430,I143621,I143609,I143618,I143627,I143606,I143624,I143615,I143630,I143603,I143612,I143600,I145295,I145310,I145292,I145307,I145289,I145286,I145301,I145298,I145304,I145313,I145283,I145941,I145956,I145938,I145953,I145935,I145932,I145947,I145944,I145950,I145959,I145929,I146587,I146581,I146578,I146590,I146575,I146596,I146605,I146599,I146602,I146593,I146584,I149084,I149057,I149078,I149063,I149060,I149066,I149072,I149087,I149075,I149081,I149069,I149713,I149701,I149704,I149689,I149695,I149707,I149716,I149686,I149710,I149698,I149692,I150285,I150273,I150282,I150291,I150270,I150288,I150279,I150294,I150267,I150276,I150264,I150852,I150837,I150834,I150831,I150849,I150846,I150825,I150828,I150855,I150840,I150843;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2703,I2711,I2719,I2727,I2735,I2743,I2751,I2759,I2767,I2775,I2783,I2791,I2799,I2807,I2815,I2823,I2831,I2839,I2847,I2855,I2863,I2871,I2879,I2887,I2895,I2903,I2911,I2919,I2927,I2935,I2943,I2951,I2959,I2966,I2973,I3014,I3031,I3048,I3065,I3082,I3099,I2997,I2985,I3144,I3161,I3178,I3195,I3212,I2994,I3243,I3260,I3277,I3294,I3003,I2982,I3339,I3356,I3000,I3387,I2991,I3006,I3432,I3449,I3466,I3483,I2979,I2988,I2976,I3575,I3592,I3609,I3626,I3643,I3660,I3558,I3546,I3705,I3722,I3739,I3756,I3773,I3555,I3804,I3821,I3838,I3855,I3564,I3543,I3900,I3917,I3561,I3948,I3552,I3567,I3993,I4010,I4027,I4044,I3540,I3549,I3537,I4136,I4153,I4170,I4187,I4204,I4221,I4119,I4107,I4266,I4283,I4300,I4317,I4334,I4116,I4365,I4382,I4399,I4416,I4125,I4104,I4461,I4478,I4122,I4509,I4113,I4128,I4554,I4571,I4588,I4605,I4101,I4110,I4098,I4697,I4714,I4731,I4748,I4671,I4779,I4796,I4686,I4668,I4841,I4858,I4875,I4892,I4909,I4926,I4943,I4960,I4977,I4683,I5008,I5025,I5042,I4665,I5073,I4662,I5104,I5121,I5138,I5155,I4677,I5186,I4674,I5217,I5234,I5251,I4680,I4689,I4659,I5343,I5360,I5377,I5394,I5317,I5425,I5442,I5332,I5314,I5487,I5504,I5521,I5538,I5555,I5572,I5589,I5606,I5623,I5329,I5654,I5671,I5688,I5311,I5719,I5308,I5750,I5767,I5784,I5801,I5323,I5832,I5320,I5863,I5880,I5897,I5326,I5335,I5305,I5989,I6006,I6023,I6040,I5960,I6071,I6088,I6105,I6122,I6139,I6156,I6173,I6190,I6207,I6224,I5975,I5972,I6269,I5957,I6300,I5954,I6331,I6348,I6365,I6382,I6399,I6416,I5981,I6447,I5969,I5963,I6492,I6509,I5978,I6540,I6557,I6574,I5966,I5951,I6652,I6669,I6635,I6614,I6714,I6731,I6748,I6765,I6782,I6799,I6816,I6833,I6850,I6641,I6881,I6898,I6915,I6932,I6644,I6963,I6980,I6997,I7014,I7031,I6629,I7062,I7079,I6632,I6626,I6620,I7138,I6638,I7169,I6623,I6617,I7247,I7264,I7281,I7298,I7315,I7332,I7349,I7366,I7236,I7397,I7221,I7428,I7445,I7462,I7479,I7496,I7513,I7530,I7218,I7561,I7578,I7215,I7609,I7626,I7233,I7657,I7230,I7688,I7705,I7209,I7212,I7750,I7767,I7784,I7801,I7239,I7832,I7224,I7227,I7910,I7927,I7944,I7961,I7978,I7995,I8012,I8029,I7899,I8060,I7884,I8091,I8108,I8125,I8142,I8159,I8176,I8193,I7881,I8224,I8241,I7878,I8272,I8289,I7896,I8320,I7893,I8351,I8368,I7872,I7875,I8413,I8430,I8447,I8464,I7902,I8495,I7887,I7890,I8573,I8590,I8607,I8624,I8641,I8658,I8675,I8692,I8562,I8723,I8547,I8754,I8771,I8788,I8805,I8822,I8839,I8856,I8544,I8887,I8904,I8541,I8935,I8952,I8559,I8983,I8556,I9014,I9031,I8535,I8538,I9076,I9093,I9110,I9127,I8565,I9158,I8550,I8553,I9236,I9253,I9270,I9287,I9304,I9321,I9338,I9355,I9225,I9386,I9210,I9417,I9434,I9451,I9468,I9485,I9502,I9519,I9207,I9550,I9567,I9204,I9598,I9615,I9222,I9646,I9219,I9677,I9694,I9198,I9201,I9739,I9756,I9773,I9790,I9228,I9821,I9213,I9216,I9899,I9916,I9933,I9950,I9967,I9984,I10001,I9870,I10032,I10049,I10066,I10083,I10100,I10117,I10134,I9867,I10165,I9861,I10196,I10213,I10230,I9891,I9864,I10275,I9888,I10306,I9885,I9882,I10351,I10368,I10385,I10402,I10419,I9876,I10450,I10467,I9879,I9873,I10545,I10562,I10579,I10596,I10613,I10630,I10647,I10516,I10678,I10695,I10712,I10729,I10746,I10763,I10780,I10513,I10811,I10507,I10842,I10859,I10876,I10537,I10510,I10921,I10534,I10952,I10531,I10528,I10997,I11014,I11031,I11048,I11065,I10522,I11096,I11113,I10525,I10519,I11191,I11208,I11225,I11242,I11259,I11276,I11293,I11162,I11324,I11341,I11358,I11375,I11392,I11409,I11426,I11159,I11457,I11153,I11488,I11505,I11522,I11183,I11156,I11567,I11180,I11598,I11177,I11174,I11643,I11660,I11677,I11694,I11711,I11168,I11742,I11759,I11171,I11165,I11837,I11854,I11871,I11888,I11905,I11799,I11936,I11953,I11970,I11987,I12004,I12021,I11808,I12052,I11802,I12083,I12100,I12117,I12134,I11829,I11826,I12179,I12196,I12213,I11823,I12244,I11820,I11811,I12289,I12306,I12323,I11814,I11817,I12368,I12385,I11805,I12449,I12466,I12483,I12500,I12517,I12417,I12548,I12565,I12582,I12420,I12613,I12414,I12644,I12661,I12678,I12695,I12712,I12423,I12743,I12760,I12777,I12794,I12429,I12432,I12411,I12853,I12870,I12887,I12441,I12438,I12932,I12949,I12426,I12435,I13027,I13044,I13061,I13078,I13095,I13112,I13129,I12998,I13160,I13177,I13194,I13211,I13228,I13245,I13262,I12995,I12989,I13307,I13324,I13341,I13016,I13372,I13389,I13007,I13001,I13434,I13004,I13465,I13482,I13019,I13513,I13013,I13010,I13558,I12992,I13622,I13639,I13656,I13673,I13690,I13707,I13724,I13741,I13758,I13775,I13792,I13809,I13826,I13843,I13611,I13874,I13891,I13908,I13584,I13939,I13605,I13970,I13987,I13590,I14018,I13587,I13593,I14063,I14080,I14097,I13599,I13614,I13602,I14156,I14173,I13608,I13596,I14251,I14268,I14285,I14302,I14240,I14333,I14228,I14364,I14381,I14398,I14415,I14432,I14231,I14463,I14216,I14494,I14511,I14528,I14545,I14562,I14579,I14222,I14610,I14627,I14644,I14234,I14243,I14213,I14703,I14237,I14225,I14748,I14765,I14219,I14829,I14846,I14863,I14880,I14818,I14911,I14806,I14942,I14959,I14976,I14993,I15010,I14809,I15041,I14794,I15072,I15089,I15106,I15123,I15140,I15157,I14800,I15188,I15205,I15222,I14812,I14821,I14791,I15281,I14815,I14803,I15326,I15343,I14797,I15407,I15424,I15441,I15458,I15475,I15492,I15390,I15378,I15537,I15554,I15571,I15588,I15605,I15387,I15636,I15653,I15670,I15687,I15396,I15375,I15732,I15749,I15393,I15780,I15384,I15399,I15825,I15842,I15859,I15876,I15372,I15381,I15369,I15968,I15985,I16002,I16019,I16036,I16053,I15951,I15939,I16098,I16115,I16132,I16149,I16166,I15948,I16197,I16214,I16231,I16248,I15957,I15936,I16293,I16310,I15954,I16341,I15945,I15960,I16386,I16403,I16420,I16437,I15933,I15942,I15930,I16529,I16546,I16563,I16580,I16597,I16614,I16512,I16500,I16659,I16676,I16693,I16710,I16727,I16509,I16758,I16775,I16792,I16809,I16518,I16497,I16854,I16871,I16515,I16902,I16506,I16521,I16947,I16964,I16981,I16998,I16494,I16503,I16491,I17090,I17107,I17124,I17141,I17064,I17172,I17189,I17079,I17061,I17234,I17251,I17268,I17285,I17302,I17319,I17336,I17353,I17370,I17076,I17401,I17418,I17435,I17058,I17466,I17055,I17497,I17514,I17531,I17548,I17070,I17579,I17067,I17610,I17627,I17644,I17073,I17082,I17052,I17736,I17753,I17770,I17787,I17710,I17818,I17835,I17725,I17707,I17880,I17897,I17914,I17931,I17948,I17965,I17982,I17999,I18016,I17722,I18047,I18064,I18081,I17704,I18112,I17701,I18143,I18160,I18177,I18194,I17716,I18225,I17713,I18256,I18273,I18290,I17719,I17728,I17698,I18382,I18399,I18416,I18433,I18356,I18464,I18481,I18371,I18353,I18526,I18543,I18560,I18577,I18594,I18611,I18628,I18645,I18662,I18368,I18693,I18710,I18727,I18350,I18758,I18347,I18789,I18806,I18823,I18840,I18362,I18871,I18359,I18902,I18919,I18936,I18365,I18374,I18344,I19028,I19045,I19062,I19079,I18999,I19110,I19127,I19144,I19161,I19178,I19195,I19212,I19229,I19246,I19263,I19014,I19011,I19308,I18996,I19339,I18993,I19370,I19387,I19404,I19421,I19438,I19455,I19020,I19486,I19008,I19002,I19531,I19548,I19017,I19579,I19596,I19613,I19005,I18990,I19691,I19708,I19725,I19665,I19756,I19773,I19790,I19807,I19824,I19841,I19858,I19875,I19892,I19659,I19923,I19940,I19656,I19971,I19988,I20005,I19668,I19653,I20050,I20067,I20084,I20101,I20118,I19674,I20149,I19683,I20180,I19677,I19680,I19671,I19662,I20286,I20303,I20320,I20337,I20354,I20371,I20388,I20405,I20275,I20436,I20260,I20467,I20484,I20501,I20518,I20535,I20552,I20569,I20257,I20600,I20617,I20254,I20648,I20665,I20272,I20696,I20269,I20727,I20744,I20248,I20251,I20789,I20806,I20823,I20840,I20278,I20871,I20263,I20266,I20949,I20966,I20983,I21000,I21017,I21034,I21051,I21068,I20938,I21099,I20923,I21130,I21147,I21164,I21181,I21198,I21215,I21232,I20920,I21263,I21280,I20917,I21311,I21328,I20935,I21359,I20932,I21390,I21407,I20911,I20914,I21452,I21469,I21486,I21503,I20941,I21534,I20926,I20929,I21612,I21629,I21646,I21663,I21680,I21697,I21714,I21731,I21601,I21762,I21586,I21793,I21810,I21827,I21844,I21861,I21878,I21895,I21583,I21926,I21943,I21580,I21974,I21991,I21598,I22022,I21595,I22053,I22070,I21574,I21577,I22115,I22132,I22149,I22166,I21604,I22197,I21589,I21592,I22275,I22292,I22309,I22326,I22343,I22360,I22377,I22394,I22264,I22425,I22249,I22456,I22473,I22490,I22507,I22524,I22541,I22558,I22246,I22589,I22606,I22243,I22637,I22654,I22261,I22685,I22258,I22716,I22733,I22237,I22240,I22778,I22795,I22812,I22829,I22267,I22860,I22252,I22255,I22938,I22955,I22972,I22989,I23006,I23023,I23040,I23057,I22927,I23088,I22912,I23119,I23136,I23153,I23170,I23187,I23204,I23221,I22909,I23252,I23269,I22906,I23300,I23317,I22924,I23348,I22921,I23379,I23396,I22900,I22903,I23441,I23458,I23475,I23492,I22930,I23523,I22915,I22918,I23601,I23618,I23635,I23652,I23669,I23686,I23703,I23720,I23590,I23751,I23575,I23782,I23799,I23816,I23833,I23850,I23867,I23884,I23572,I23915,I23932,I23569,I23963,I23980,I23587,I24011,I23584,I24042,I24059,I23563,I23566,I24104,I24121,I24138,I24155,I23593,I24186,I23578,I23581,I24264,I24281,I24298,I24315,I24332,I24349,I24366,I24235,I24397,I24414,I24431,I24448,I24465,I24482,I24499,I24232,I24530,I24226,I24561,I24578,I24595,I24256,I24229,I24640,I24253,I24671,I24250,I24247,I24716,I24733,I24750,I24767,I24784,I24241,I24815,I24832,I24244,I24238,I24910,I24927,I24944,I24961,I24978,I24878,I25009,I25026,I25043,I24881,I25074,I24875,I25105,I25122,I25139,I25156,I25173,I24884,I25204,I25221,I25238,I25255,I24890,I24893,I24872,I25314,I25331,I25348,I24902,I24899,I25393,I25410,I24887,I24896,I25488,I25505,I25522,I25539,I25556,I25456,I25587,I25604,I25621,I25459,I25652,I25453,I25683,I25700,I25717,I25734,I25751,I25462,I25782,I25799,I25816,I25833,I25468,I25471,I25450,I25892,I25909,I25926,I25480,I25477,I25971,I25988,I25465,I25474,I26066,I26083,I26100,I26117,I26134,I26034,I26165,I26182,I26199,I26037,I26230,I26031,I26261,I26278,I26295,I26312,I26329,I26040,I26360,I26377,I26394,I26411,I26046,I26049,I26028,I26470,I26487,I26504,I26058,I26055,I26549,I26566,I26043,I26052,I26644,I26661,I26678,I26695,I26712,I26612,I26743,I26760,I26777,I26615,I26808,I26609,I26839,I26856,I26873,I26890,I26907,I26618,I26938,I26955,I26972,I26989,I26624,I26627,I26606,I27048,I27065,I27082,I26636,I26633,I27127,I27144,I26621,I26630,I27222,I27239,I27256,I27273,I27290,I27190,I27321,I27338,I27355,I27193,I27386,I27187,I27417,I27434,I27451,I27468,I27485,I27196,I27516,I27533,I27550,I27567,I27202,I27205,I27184,I27626,I27643,I27660,I27214,I27211,I27705,I27722,I27199,I27208,I27800,I27817,I27834,I27851,I27868,I27768,I27899,I27916,I27933,I27950,I27967,I27984,I28001,I28018,I27774,I27765,I28063,I28080,I27789,I28111,I28128,I27777,I28159,I28176,I27783,I28207,I27771,I28238,I27762,I28269,I28286,I27792,I28317,I27786,I28348,I27780,I28412,I28429,I28446,I28463,I28401,I28494,I28511,I28528,I28545,I28562,I28579,I28596,I28386,I28627,I28383,I28658,I28395,I28689,I28706,I28723,I28389,I28404,I28768,I28785,I28374,I28816,I28392,I28847,I28864,I28398,I28895,I28912,I28377,I28380,I28990,I29007,I29024,I29041,I28979,I29072,I29089,I29106,I29123,I29140,I29157,I29174,I28964,I29205,I28961,I29236,I28973,I29267,I29284,I29301,I28967,I28982,I29346,I29363,I28952,I29394,I28970,I29425,I29442,I28976,I29473,I29490,I28955,I28958,I29568,I29585,I29602,I29619,I29636,I29653,I29551,I29684,I29701,I29718,I29554,I29536,I29763,I29780,I29797,I29557,I29548,I29842,I29859,I29876,I29539,I29907,I29924,I29530,I29955,I29972,I29989,I29560,I30020,I30037,I30054,I30071,I29545,I29542,I29533,I30163,I30180,I30197,I30214,I30231,I30248,I30146,I30279,I30296,I30313,I30149,I30131,I30358,I30375,I30392,I30152,I30143,I30437,I30454,I30471,I30134,I30502,I30519,I30125,I30550,I30567,I30584,I30155,I30615,I30632,I30649,I30666,I30140,I30137,I30128,I30758,I30775,I30792,I30809,I30826,I30843,I30741,I30874,I30891,I30908,I30744,I30726,I30953,I30970,I30987,I30747,I30738,I31032,I31049,I31066,I30729,I31097,I31114,I30720,I31145,I31162,I31179,I30750,I31210,I31227,I31244,I31261,I30735,I30732,I30723,I31353,I31370,I31387,I31404,I31421,I31438,I31336,I31469,I31486,I31503,I31339,I31321,I31548,I31565,I31582,I31342,I31333,I31627,I31644,I31661,I31324,I31692,I31709,I31315,I31740,I31757,I31774,I31345,I31805,I31822,I31839,I31856,I31330,I31327,I31318,I31948,I31965,I31982,I31999,I32016,I32033,I31931,I32064,I32081,I32098,I31934,I31916,I32143,I32160,I32177,I31937,I31928,I32222,I32239,I32256,I31919,I32287,I32304,I31910,I32335,I32352,I32369,I31940,I32400,I32417,I32434,I32451,I31925,I31922,I31913,I32543,I32560,I32577,I32594,I32611,I32628,I32645,I32514,I32676,I32693,I32710,I32727,I32744,I32761,I32778,I32511,I32505,I32823,I32840,I32857,I32532,I32888,I32905,I32523,I32517,I32950,I32520,I32981,I32998,I32535,I33029,I32529,I32526,I33074,I32508,I33138,I33155,I33172,I33189,I33206,I33223,I33240,I33257,I33274,I33291,I33308,I33325,I33342,I33359,I33127,I33390,I33407,I33424,I33100,I33455,I33121,I33486,I33503,I33106,I33534,I33103,I33109,I33579,I33596,I33613,I33115,I33130,I33118,I33672,I33689,I33124,I33112,I33767,I33784,I33801,I33818,I33835,I33852,I33869,I33886,I33903,I33920,I33937,I33954,I33971,I33988,I33756,I34019,I34036,I34053,I33729,I34084,I33750,I34115,I34132,I33735,I34163,I33732,I33738,I34208,I34225,I34242,I33744,I33759,I33747,I34301,I34318,I33753,I33741,I34396,I34413,I34430,I34447,I34464,I34481,I34498,I34515,I34532,I34549,I34566,I34583,I34600,I34617,I34385,I34648,I34665,I34682,I34358,I34713,I34379,I34744,I34761,I34364,I34792,I34361,I34367,I34837,I34854,I34871,I34373,I34388,I34376,I34930,I34947,I34382,I34370,I35025,I35042,I35059,I35076,I35093,I35110,I35127,I35144,I35161,I35178,I35195,I35212,I35229,I35246,I35014,I35277,I35294,I35311,I34987,I35342,I35008,I35373,I35390,I34993,I35421,I34990,I34996,I35466,I35483,I35500,I35002,I35017,I35005,I35559,I35576,I35011,I34999,I35654,I35671,I35688,I35705,I35722,I35739,I35756,I35773,I35790,I35807,I35824,I35841,I35858,I35875,I35643,I35906,I35923,I35940,I35616,I35971,I35637,I36002,I36019,I35622,I36050,I35619,I35625,I36095,I36112,I36129,I35631,I35646,I35634,I36188,I36205,I35640,I35628,I36283,I36300,I36317,I36334,I36272,I36365,I36260,I36396,I36413,I36430,I36447,I36464,I36263,I36495,I36248,I36526,I36543,I36560,I36577,I36594,I36611,I36254,I36642,I36659,I36676,I36266,I36275,I36245,I36735,I36269,I36257,I36780,I36797,I36251,I36861,I36878,I36895,I36912,I36835,I36943,I36960,I36850,I36832,I37005,I37022,I37039,I37056,I37073,I37090,I37107,I37124,I37141,I36847,I37172,I37189,I37206,I36829,I37237,I36826,I37268,I37285,I37302,I37319,I36841,I37350,I36838,I37381,I37398,I37415,I36844,I36853,I36823,I37507,I37524,I37541,I37558,I37478,I37589,I37606,I37623,I37640,I37657,I37674,I37691,I37708,I37725,I37742,I37493,I37490,I37787,I37475,I37818,I37472,I37849,I37866,I37883,I37900,I37917,I37934,I37499,I37965,I37487,I37481,I38010,I38027,I37496,I38058,I38075,I38092,I37484,I37469,I38170,I38187,I38204,I38221,I38141,I38252,I38269,I38286,I38303,I38320,I38337,I38354,I38371,I38388,I38405,I38156,I38153,I38450,I38138,I38481,I38135,I38512,I38529,I38546,I38563,I38580,I38597,I38162,I38628,I38150,I38144,I38673,I38690,I38159,I38721,I38738,I38755,I38147,I38132,I38833,I38850,I38867,I38807,I38898,I38915,I38932,I38949,I38966,I38983,I39000,I39017,I39034,I38801,I39065,I39082,I38798,I39113,I39130,I39147,I38810,I38795,I39192,I39209,I39226,I39243,I39260,I38816,I39291,I38825,I39322,I38819,I38822,I38813,I38804,I39428,I39445,I39411,I39390,I39490,I39507,I39524,I39541,I39558,I39575,I39592,I39609,I39626,I39417,I39657,I39674,I39691,I39708,I39420,I39739,I39756,I39773,I39790,I39807,I39405,I39838,I39855,I39408,I39402,I39396,I39914,I39414,I39945,I39399,I39393,I40023,I40040,I40006,I39985,I40085,I40102,I40119,I40136,I40153,I40170,I40187,I40204,I40221,I40012,I40252,I40269,I40286,I40303,I40015,I40334,I40351,I40368,I40385,I40402,I40000,I40433,I40450,I40003,I39997,I39991,I40509,I40009,I40540,I39994,I39988,I40618,I40635,I40601,I40580,I40680,I40697,I40714,I40731,I40748,I40765,I40782,I40799,I40816,I40607,I40847,I40864,I40881,I40898,I40610,I40929,I40946,I40963,I40980,I40997,I40595,I41028,I41045,I40598,I40592,I40586,I41104,I40604,I41135,I40589,I40583,I41213,I41230,I41247,I41264,I41281,I41298,I41315,I41332,I41202,I41363,I41187,I41394,I41411,I41428,I41445,I41462,I41479,I41496,I41184,I41527,I41544,I41181,I41575,I41592,I41199,I41623,I41196,I41654,I41671,I41175,I41178,I41716,I41733,I41750,I41767,I41205,I41798,I41190,I41193,I41876,I41893,I41910,I41927,I41944,I41961,I41978,I41995,I41865,I42026,I41850,I42057,I42074,I42091,I42108,I42125,I42142,I42159,I41847,I42190,I42207,I41844,I42238,I42255,I41862,I42286,I41859,I42317,I42334,I41838,I41841,I42379,I42396,I42413,I42430,I41868,I42461,I41853,I41856,I42539,I42556,I42573,I42590,I42607,I42624,I42641,I42658,I42528,I42689,I42513,I42720,I42737,I42754,I42771,I42788,I42805,I42822,I42510,I42853,I42870,I42507,I42901,I42918,I42525,I42949,I42522,I42980,I42997,I42501,I42504,I43042,I43059,I43076,I43093,I42531,I43124,I42516,I42519,I43202,I43219,I43236,I43253,I43270,I43287,I43304,I43321,I43191,I43352,I43176,I43383,I43400,I43417,I43434,I43451,I43468,I43485,I43173,I43516,I43533,I43170,I43564,I43581,I43188,I43612,I43185,I43643,I43660,I43164,I43167,I43705,I43722,I43739,I43756,I43194,I43787,I43179,I43182,I43865,I43882,I43899,I43916,I43933,I43950,I43967,I43984,I43854,I44015,I43839,I44046,I44063,I44080,I44097,I44114,I44131,I44148,I43836,I44179,I44196,I43833,I44227,I44244,I43851,I44275,I43848,I44306,I44323,I43827,I43830,I44368,I44385,I44402,I44419,I43857,I44450,I43842,I43845,I44528,I44545,I44562,I44579,I44596,I44613,I44630,I44647,I44517,I44678,I44502,I44709,I44726,I44743,I44760,I44777,I44794,I44811,I44499,I44842,I44859,I44496,I44890,I44907,I44514,I44938,I44511,I44969,I44986,I44490,I44493,I45031,I45048,I45065,I45082,I44520,I45113,I44505,I44508,I45191,I45208,I45225,I45242,I45259,I45276,I45293,I45310,I45180,I45341,I45165,I45372,I45389,I45406,I45423,I45440,I45457,I45474,I45162,I45505,I45522,I45159,I45553,I45570,I45177,I45601,I45174,I45632,I45649,I45153,I45156,I45694,I45711,I45728,I45745,I45183,I45776,I45168,I45171,I45854,I45871,I45888,I45905,I45922,I45939,I45956,I45825,I45987,I46004,I46021,I46038,I46055,I46072,I46089,I45822,I46120,I45816,I46151,I46168,I46185,I45846,I45819,I46230,I45843,I46261,I45840,I45837,I46306,I46323,I46340,I46357,I46374,I45831,I46405,I46422,I45834,I45828,I46500,I46517,I46534,I46551,I46568,I46585,I46602,I46471,I46633,I46650,I46667,I46684,I46701,I46718,I46735,I46468,I46766,I46462,I46797,I46814,I46831,I46492,I46465,I46876,I46489,I46907,I46486,I46483,I46952,I46969,I46986,I47003,I47020,I46477,I47051,I47068,I46480,I46474,I47146,I47163,I47180,I47197,I47214,I47231,I47248,I47117,I47279,I47296,I47313,I47330,I47347,I47364,I47381,I47114,I47412,I47108,I47443,I47460,I47477,I47138,I47111,I47522,I47135,I47553,I47132,I47129,I47598,I47615,I47632,I47649,I47666,I47123,I47697,I47714,I47126,I47120,I47792,I47809,I47826,I47843,I47860,I47877,I47894,I47763,I47925,I47942,I47959,I47976,I47993,I48010,I48027,I47760,I48058,I47754,I48089,I48106,I48123,I47784,I47757,I48168,I47781,I48199,I47778,I47775,I48244,I48261,I48278,I48295,I48312,I47769,I48343,I48360,I47772,I47766,I48438,I48455,I48472,I48489,I48506,I48523,I48540,I48409,I48571,I48588,I48605,I48622,I48639,I48656,I48673,I48406,I48704,I48400,I48735,I48752,I48769,I48430,I48403,I48814,I48427,I48845,I48424,I48421,I48890,I48907,I48924,I48941,I48958,I48415,I48989,I49006,I48418,I48412,I49084,I49101,I49118,I49135,I49152,I49046,I49183,I49200,I49217,I49234,I49251,I49268,I49055,I49299,I49049,I49330,I49347,I49364,I49381,I49076,I49073,I49426,I49443,I49460,I49070,I49491,I49067,I49058,I49536,I49553,I49570,I49061,I49064,I49615,I49632,I49052,I49696,I49713,I49730,I49747,I49764,I49658,I49795,I49812,I49829,I49846,I49863,I49880,I49667,I49911,I49661,I49942,I49959,I49976,I49993,I49688,I49685,I50038,I50055,I50072,I49682,I50103,I49679,I49670,I50148,I50165,I50182,I49673,I49676,I50227,I50244,I49664,I50308,I50325,I50342,I50359,I50376,I50276,I50407,I50424,I50441,I50279,I50472,I50273,I50503,I50520,I50537,I50554,I50571,I50282,I50602,I50619,I50636,I50653,I50288,I50291,I50270,I50712,I50729,I50746,I50300,I50297,I50791,I50808,I50285,I50294,I50886,I50903,I50920,I50937,I50954,I50854,I50985,I51002,I51019,I50857,I51050,I50851,I51081,I51098,I51115,I51132,I51149,I50860,I51180,I51197,I51214,I51231,I50866,I50869,I50848,I51290,I51307,I51324,I50878,I50875,I51369,I51386,I50863,I50872,I51464,I51481,I51498,I51515,I51532,I51432,I51563,I51580,I51597,I51435,I51628,I51429,I51659,I51676,I51693,I51710,I51727,I51438,I51758,I51775,I51792,I51809,I51444,I51447,I51426,I51868,I51885,I51902,I51456,I51453,I51947,I51964,I51441,I51450,I52042,I52059,I52076,I52093,I52110,I52010,I52141,I52158,I52175,I52013,I52206,I52007,I52237,I52254,I52271,I52288,I52305,I52016,I52336,I52353,I52370,I52387,I52022,I52025,I52004,I52446,I52463,I52480,I52034,I52031,I52525,I52542,I52019,I52028,I52620,I52637,I52654,I52671,I52688,I52588,I52719,I52736,I52753,I52591,I52784,I52585,I52815,I52832,I52849,I52866,I52883,I52594,I52914,I52931,I52948,I52965,I52600,I52603,I52582,I53024,I53041,I53058,I52612,I52609,I53103,I53120,I52597,I52606,I53198,I53215,I53232,I53249,I53266,I53166,I53297,I53314,I53331,I53169,I53362,I53163,I53393,I53410,I53427,I53444,I53461,I53172,I53492,I53509,I53526,I53543,I53178,I53181,I53160,I53602,I53619,I53636,I53190,I53187,I53681,I53698,I53175,I53184,I53776,I53793,I53810,I53827,I53844,I53861,I53759,I53892,I53909,I53926,I53762,I53744,I53971,I53988,I54005,I53765,I53756,I54050,I54067,I54084,I53747,I54115,I54132,I53738,I54163,I54180,I54197,I53768,I54228,I54245,I54262,I54279,I53753,I53750,I53741,I54371,I54388,I54405,I54422,I54439,I54456,I54354,I54487,I54504,I54521,I54357,I54339,I54566,I54583,I54600,I54360,I54351,I54645,I54662,I54679,I54342,I54710,I54727,I54333,I54758,I54775,I54792,I54363,I54823,I54840,I54857,I54874,I54348,I54345,I54336,I54966,I54983,I55000,I55017,I55034,I55051,I54949,I55082,I55099,I55116,I54952,I54934,I55161,I55178,I55195,I54955,I54946,I55240,I55257,I55274,I54937,I55305,I55322,I54928,I55353,I55370,I55387,I54958,I55418,I55435,I55452,I55469,I54943,I54940,I54931,I55561,I55578,I55595,I55612,I55629,I55646,I55544,I55677,I55694,I55711,I55547,I55529,I55756,I55773,I55790,I55550,I55541,I55835,I55852,I55869,I55532,I55900,I55917,I55523,I55948,I55965,I55982,I55553,I56013,I56030,I56047,I56064,I55538,I55535,I55526,I56156,I56173,I56190,I56207,I56224,I56241,I56139,I56272,I56289,I56306,I56142,I56124,I56351,I56368,I56385,I56145,I56136,I56430,I56447,I56464,I56127,I56495,I56512,I56118,I56543,I56560,I56577,I56148,I56608,I56625,I56642,I56659,I56133,I56130,I56121,I56751,I56768,I56785,I56802,I56819,I56836,I56853,I56722,I56884,I56901,I56918,I56935,I56952,I56969,I56986,I56719,I56713,I57031,I57048,I57065,I56740,I57096,I57113,I56731,I56725,I57158,I56728,I57189,I57206,I56743,I57237,I56737,I56734,I57282,I56716,I57346,I57363,I57380,I57397,I57414,I57431,I57448,I57317,I57479,I57496,I57513,I57530,I57547,I57564,I57581,I57314,I57308,I57626,I57643,I57660,I57335,I57691,I57708,I57326,I57320,I57753,I57323,I57784,I57801,I57338,I57832,I57332,I57329,I57877,I57311,I57941,I57958,I57975,I57992,I58009,I58026,I58043,I57912,I58074,I58091,I58108,I58125,I58142,I58159,I58176,I57909,I57903,I58221,I58238,I58255,I57930,I58286,I58303,I57921,I57915,I58348,I57918,I58379,I58396,I57933,I58427,I57927,I57924,I58472,I57906,I58536,I58553,I58570,I58587,I58604,I58621,I58638,I58655,I58672,I58689,I58706,I58723,I58740,I58757,I58525,I58788,I58805,I58822,I58498,I58853,I58519,I58884,I58901,I58504,I58932,I58501,I58507,I58977,I58994,I59011,I58513,I58528,I58516,I59070,I59087,I58522,I58510,I59165,I59182,I59199,I59216,I59233,I59250,I59267,I59284,I59301,I59318,I59335,I59352,I59369,I59386,I59154,I59417,I59434,I59451,I59127,I59482,I59148,I59513,I59530,I59133,I59561,I59130,I59136,I59606,I59623,I59640,I59142,I59157,I59145,I59699,I59716,I59151,I59139,I59794,I59811,I59828,I59845,I59862,I59879,I59896,I59913,I59930,I59947,I59964,I59981,I59998,I60015,I59783,I60046,I60063,I60080,I59756,I60111,I59777,I60142,I60159,I59762,I60190,I59759,I59765,I60235,I60252,I60269,I59771,I59786,I59774,I60328,I60345,I59780,I59768,I60423,I60440,I60457,I60474,I60491,I60508,I60406,I60394,I60553,I60570,I60587,I60604,I60621,I60403,I60652,I60669,I60686,I60703,I60412,I60391,I60748,I60765,I60409,I60796,I60400,I60415,I60841,I60858,I60875,I60892,I60388,I60397,I60385,I60984,I61001,I61018,I61035,I60958,I61066,I61083,I60973,I60955,I61128,I61145,I61162,I61179,I61196,I61213,I61230,I61247,I61264,I60970,I61295,I61312,I61329,I60952,I61360,I60949,I61391,I61408,I61425,I61442,I60964,I61473,I60961,I61504,I61521,I61538,I60967,I60976,I60946,I61630,I61647,I61664,I61681,I61604,I61712,I61729,I61619,I61601,I61774,I61791,I61808,I61825,I61842,I61859,I61876,I61893,I61910,I61616,I61941,I61958,I61975,I61598,I62006,I61595,I62037,I62054,I62071,I62088,I61610,I62119,I61607,I62150,I62167,I62184,I61613,I61622,I61592,I62276,I62293,I62310,I62327,I62250,I62358,I62375,I62265,I62247,I62420,I62437,I62454,I62471,I62488,I62505,I62522,I62539,I62556,I62262,I62587,I62604,I62621,I62244,I62652,I62241,I62683,I62700,I62717,I62734,I62256,I62765,I62253,I62796,I62813,I62830,I62259,I62268,I62238,I62922,I62939,I62956,I62973,I62896,I63004,I63021,I62911,I62893,I63066,I63083,I63100,I63117,I63134,I63151,I63168,I63185,I63202,I62908,I63233,I63250,I63267,I62890,I63298,I62887,I63329,I63346,I63363,I63380,I62902,I63411,I62899,I63442,I63459,I63476,I62905,I62914,I62884,I63568,I63585,I63602,I63619,I63542,I63650,I63667,I63557,I63539,I63712,I63729,I63746,I63763,I63780,I63797,I63814,I63831,I63848,I63554,I63879,I63896,I63913,I63536,I63944,I63533,I63975,I63992,I64009,I64026,I63548,I64057,I63545,I64088,I64105,I64122,I63551,I63560,I63530,I64214,I64231,I64248,I64265,I64188,I64296,I64313,I64203,I64185,I64358,I64375,I64392,I64409,I64426,I64443,I64460,I64477,I64494,I64200,I64525,I64542,I64559,I64182,I64590,I64179,I64621,I64638,I64655,I64672,I64194,I64703,I64191,I64734,I64751,I64768,I64197,I64206,I64176,I64860,I64877,I64894,I64911,I64834,I64942,I64959,I64849,I64831,I65004,I65021,I65038,I65055,I65072,I65089,I65106,I65123,I65140,I64846,I65171,I65188,I65205,I64828,I65236,I64825,I65267,I65284,I65301,I65318,I64840,I65349,I64837,I65380,I65397,I65414,I64843,I64852,I64822,I65506,I65523,I65540,I65557,I65480,I65588,I65605,I65495,I65477,I65650,I65667,I65684,I65701,I65718,I65735,I65752,I65769,I65786,I65492,I65817,I65834,I65851,I65474,I65882,I65471,I65913,I65930,I65947,I65964,I65486,I65995,I65483,I66026,I66043,I66060,I65489,I65498,I65468,I66152,I66169,I66186,I66203,I66123,I66234,I66251,I66268,I66285,I66302,I66319,I66336,I66353,I66370,I66387,I66138,I66135,I66432,I66120,I66463,I66117,I66494,I66511,I66528,I66545,I66562,I66579,I66144,I66610,I66132,I66126,I66655,I66672,I66141,I66703,I66720,I66737,I66129,I66114,I66815,I66832,I66849,I66866,I66786,I66897,I66914,I66931,I66948,I66965,I66982,I66999,I67016,I67033,I67050,I66801,I66798,I67095,I66783,I67126,I66780,I67157,I67174,I67191,I67208,I67225,I67242,I66807,I67273,I66795,I66789,I67318,I67335,I66804,I67366,I67383,I67400,I66792,I66777,I67478,I67495,I67512,I67452,I67543,I67560,I67577,I67594,I67611,I67628,I67645,I67662,I67679,I67446,I67710,I67727,I67443,I67758,I67775,I67792,I67455,I67440,I67837,I67854,I67871,I67888,I67905,I67461,I67936,I67470,I67967,I67464,I67467,I67458,I67449,I68073,I68090,I68107,I68047,I68138,I68155,I68172,I68189,I68206,I68223,I68240,I68257,I68274,I68041,I68305,I68322,I68038,I68353,I68370,I68387,I68050,I68035,I68432,I68449,I68466,I68483,I68500,I68056,I68531,I68065,I68562,I68059,I68062,I68053,I68044,I68668,I68685,I68702,I68719,I68736,I68753,I68770,I68787,I68657,I68818,I68642,I68849,I68866,I68883,I68900,I68917,I68934,I68951,I68639,I68982,I68999,I68636,I69030,I69047,I68654,I69078,I68651,I69109,I69126,I68630,I68633,I69171,I69188,I69205,I69222,I68660,I69253,I68645,I68648,I69331,I69348,I69365,I69382,I69399,I69416,I69433,I69450,I69320,I69481,I69305,I69512,I69529,I69546,I69563,I69580,I69597,I69614,I69302,I69645,I69662,I69299,I69693,I69710,I69317,I69741,I69314,I69772,I69789,I69293,I69296,I69834,I69851,I69868,I69885,I69323,I69916,I69308,I69311,I69994,I70011,I70028,I70045,I70062,I70079,I70096,I70113,I69983,I70144,I69968,I70175,I70192,I70209,I70226,I70243,I70260,I70277,I69965,I70308,I70325,I69962,I70356,I70373,I69980,I70404,I69977,I70435,I70452,I69956,I69959,I70497,I70514,I70531,I70548,I69986,I70579,I69971,I69974,I70657,I70674,I70691,I70708,I70725,I70742,I70759,I70776,I70646,I70807,I70631,I70838,I70855,I70872,I70889,I70906,I70923,I70940,I70628,I70971,I70988,I70625,I71019,I71036,I70643,I71067,I70640,I71098,I71115,I70619,I70622,I71160,I71177,I71194,I71211,I70649,I71242,I70634,I70637,I71320,I71337,I71354,I71371,I71388,I71405,I71422,I71439,I71309,I71470,I71294,I71501,I71518,I71535,I71552,I71569,I71586,I71603,I71291,I71634,I71651,I71288,I71682,I71699,I71306,I71730,I71303,I71761,I71778,I71282,I71285,I71823,I71840,I71857,I71874,I71312,I71905,I71297,I71300,I71983,I72000,I72017,I72034,I72051,I72068,I72085,I72102,I71972,I72133,I71957,I72164,I72181,I72198,I72215,I72232,I72249,I72266,I71954,I72297,I72314,I71951,I72345,I72362,I71969,I72393,I71966,I72424,I72441,I71945,I71948,I72486,I72503,I72520,I72537,I71975,I72568,I71960,I71963,I72646,I72663,I72680,I72697,I72714,I72731,I72748,I72765,I72635,I72796,I72620,I72827,I72844,I72861,I72878,I72895,I72912,I72929,I72617,I72960,I72977,I72614,I73008,I73025,I72632,I73056,I72629,I73087,I73104,I72608,I72611,I73149,I73166,I73183,I73200,I72638,I73231,I72623,I72626,I73309,I73326,I73343,I73360,I73377,I73394,I73411,I73280,I73442,I73459,I73476,I73493,I73510,I73527,I73544,I73277,I73575,I73271,I73606,I73623,I73640,I73301,I73274,I73685,I73298,I73716,I73295,I73292,I73761,I73778,I73795,I73812,I73829,I73286,I73860,I73877,I73289,I73283,I73955,I73972,I73989,I74006,I74023,I74040,I74057,I73926,I74088,I74105,I74122,I74139,I74156,I74173,I74190,I73923,I74221,I73917,I74252,I74269,I74286,I73947,I73920,I74331,I73944,I74362,I73941,I73938,I74407,I74424,I74441,I74458,I74475,I73932,I74506,I74523,I73935,I73929,I74601,I74618,I74635,I74652,I74669,I74686,I74703,I74572,I74734,I74751,I74768,I74785,I74802,I74819,I74836,I74569,I74867,I74563,I74898,I74915,I74932,I74593,I74566,I74977,I74590,I75008,I74587,I74584,I75053,I75070,I75087,I75104,I75121,I74578,I75152,I75169,I74581,I74575,I75247,I75264,I75281,I75298,I75315,I75332,I75349,I75218,I75380,I75397,I75414,I75431,I75448,I75465,I75482,I75215,I75513,I75209,I75544,I75561,I75578,I75239,I75212,I75623,I75236,I75654,I75233,I75230,I75699,I75716,I75733,I75750,I75767,I75224,I75798,I75815,I75227,I75221,I75893,I75910,I75927,I75944,I75961,I75978,I75995,I75864,I76026,I76043,I76060,I76077,I76094,I76111,I76128,I75861,I76159,I75855,I76190,I76207,I76224,I75885,I75858,I76269,I75882,I76300,I75879,I75876,I76345,I76362,I76379,I76396,I76413,I75870,I76444,I76461,I75873,I75867,I76539,I76556,I76573,I76590,I76607,I76507,I76638,I76655,I76672,I76510,I76703,I76504,I76734,I76751,I76768,I76785,I76802,I76513,I76833,I76850,I76867,I76884,I76519,I76522,I76501,I76943,I76960,I76977,I76531,I76528,I77022,I77039,I76516,I76525,I77117,I77134,I77151,I77168,I77185,I77085,I77216,I77233,I77250,I77088,I77281,I77082,I77312,I77329,I77346,I77363,I77380,I77091,I77411,I77428,I77445,I77462,I77097,I77100,I77079,I77521,I77538,I77555,I77109,I77106,I77600,I77617,I77094,I77103,I77695,I77712,I77729,I77746,I77763,I77663,I77794,I77811,I77828,I77666,I77859,I77660,I77890,I77907,I77924,I77941,I77958,I77669,I77989,I78006,I78023,I78040,I77675,I77678,I77657,I78099,I78116,I78133,I77687,I77684,I78178,I78195,I77672,I77681,I78273,I78290,I78307,I78324,I78341,I78358,I78256,I78389,I78406,I78423,I78259,I78241,I78468,I78485,I78502,I78262,I78253,I78547,I78564,I78581,I78244,I78612,I78629,I78235,I78660,I78677,I78694,I78265,I78725,I78742,I78759,I78776,I78250,I78247,I78238,I78868,I78885,I78902,I78919,I78936,I78953,I78851,I78984,I79001,I79018,I78854,I78836,I79063,I79080,I79097,I78857,I78848,I79142,I79159,I79176,I78839,I79207,I79224,I78830,I79255,I79272,I79289,I78860,I79320,I79337,I79354,I79371,I78845,I78842,I78833,I79463,I79480,I79497,I79514,I79531,I79548,I79446,I79579,I79596,I79613,I79449,I79431,I79658,I79675,I79692,I79452,I79443,I79737,I79754,I79771,I79434,I79802,I79819,I79425,I79850,I79867,I79884,I79455,I79915,I79932,I79949,I79966,I79440,I79437,I79428,I80058,I80075,I80092,I80109,I80126,I80143,I80041,I80174,I80191,I80208,I80044,I80026,I80253,I80270,I80287,I80047,I80038,I80332,I80349,I80366,I80029,I80397,I80414,I80020,I80445,I80462,I80479,I80050,I80510,I80527,I80544,I80561,I80035,I80032,I80023,I80653,I80670,I80687,I80704,I80721,I80738,I80755,I80624,I80786,I80803,I80820,I80837,I80854,I80871,I80888,I80621,I80615,I80933,I80950,I80967,I80642,I80998,I81015,I80633,I80627,I81060,I80630,I81091,I81108,I80645,I81139,I80639,I80636,I81184,I80618,I81248,I81265,I81282,I81299,I81316,I81333,I81350,I81219,I81381,I81398,I81415,I81432,I81449,I81466,I81483,I81216,I81210,I81528,I81545,I81562,I81237,I81593,I81610,I81228,I81222,I81655,I81225,I81686,I81703,I81240,I81734,I81234,I81231,I81779,I81213,I81843,I81860,I81877,I81894,I81911,I81928,I81945,I81814,I81976,I81993,I82010,I82027,I82044,I82061,I82078,I81811,I81805,I82123,I82140,I82157,I81832,I82188,I82205,I81823,I81817,I82250,I81820,I82281,I82298,I81835,I82329,I81829,I81826,I82374,I81808,I82438,I82455,I82472,I82489,I82506,I82523,I82540,I82409,I82571,I82588,I82605,I82622,I82639,I82656,I82673,I82406,I82400,I82718,I82735,I82752,I82427,I82783,I82800,I82418,I82412,I82845,I82415,I82876,I82893,I82430,I82924,I82424,I82421,I82969,I82403,I83033,I83050,I83067,I83084,I83101,I83118,I83135,I83152,I83169,I83186,I83203,I83220,I83237,I83254,I83022,I83285,I83302,I83319,I82995,I83350,I83016,I83381,I83398,I83001,I83429,I82998,I83004,I83474,I83491,I83508,I83010,I83025,I83013,I83567,I83584,I83019,I83007,I83662,I83679,I83696,I83713,I83730,I83747,I83764,I83781,I83798,I83815,I83832,I83849,I83866,I83883,I83651,I83914,I83931,I83948,I83624,I83979,I83645,I84010,I84027,I83630,I84058,I83627,I83633,I84103,I84120,I84137,I83639,I83654,I83642,I84196,I84213,I83648,I83636,I84291,I84308,I84325,I84342,I84359,I84376,I84393,I84410,I84427,I84444,I84461,I84478,I84495,I84512,I84280,I84543,I84560,I84577,I84253,I84608,I84274,I84639,I84656,I84259,I84687,I84256,I84262,I84732,I84749,I84766,I84268,I84283,I84271,I84825,I84842,I84277,I84265,I84920,I84937,I84954,I84971,I84988,I85005,I85022,I85039,I85056,I85073,I85090,I85107,I85124,I85141,I84909,I85172,I85189,I85206,I84882,I85237,I84903,I85268,I85285,I84888,I85316,I84885,I84891,I85361,I85378,I85395,I84897,I84912,I84900,I85454,I85471,I84906,I84894,I85549,I85566,I85583,I85600,I85538,I85631,I85526,I85662,I85679,I85696,I85713,I85730,I85529,I85761,I85514,I85792,I85809,I85826,I85843,I85860,I85877,I85520,I85908,I85925,I85942,I85532,I85541,I85511,I86001,I85535,I85523,I86046,I86063,I85517,I86127,I86144,I86161,I86178,I86195,I86212,I86110,I86098,I86257,I86274,I86291,I86308,I86325,I86107,I86356,I86373,I86390,I86407,I86116,I86095,I86452,I86469,I86113,I86500,I86104,I86119,I86545,I86562,I86579,I86596,I86092,I86101,I86089,I86688,I86705,I86722,I86739,I86756,I86773,I86671,I86659,I86818,I86835,I86852,I86869,I86886,I86668,I86917,I86934,I86951,I86968,I86677,I86656,I87013,I87030,I86674,I87061,I86665,I86680,I87106,I87123,I87140,I87157,I86653,I86662,I86650,I87249,I87266,I87283,I87300,I87317,I87334,I87232,I87220,I87379,I87396,I87413,I87430,I87447,I87229,I87478,I87495,I87512,I87529,I87238,I87217,I87574,I87591,I87235,I87622,I87226,I87241,I87667,I87684,I87701,I87718,I87214,I87223,I87211,I87810,I87827,I87844,I87861,I87784,I87892,I87909,I87799,I87781,I87954,I87971,I87988,I88005,I88022,I88039,I88056,I88073,I88090,I87796,I88121,I88138,I88155,I87778,I88186,I87775,I88217,I88234,I88251,I88268,I87790,I88299,I87787,I88330,I88347,I88364,I87793,I87802,I87772,I88456,I88473,I88490,I88507,I88430,I88538,I88555,I88445,I88427,I88600,I88617,I88634,I88651,I88668,I88685,I88702,I88719,I88736,I88442,I88767,I88784,I88801,I88424,I88832,I88421,I88863,I88880,I88897,I88914,I88436,I88945,I88433,I88976,I88993,I89010,I88439,I88448,I88418,I89102,I89119,I89136,I89153,I89076,I89184,I89201,I89091,I89073,I89246,I89263,I89280,I89297,I89314,I89331,I89348,I89365,I89382,I89088,I89413,I89430,I89447,I89070,I89478,I89067,I89509,I89526,I89543,I89560,I89082,I89591,I89079,I89622,I89639,I89656,I89085,I89094,I89064,I89748,I89765,I89782,I89799,I89722,I89830,I89847,I89737,I89719,I89892,I89909,I89926,I89943,I89960,I89977,I89994,I90011,I90028,I89734,I90059,I90076,I90093,I89716,I90124,I89713,I90155,I90172,I90189,I90206,I89728,I90237,I89725,I90268,I90285,I90302,I89731,I89740,I89710,I90394,I90411,I90428,I90445,I90365,I90476,I90493,I90510,I90527,I90544,I90561,I90578,I90595,I90612,I90629,I90380,I90377,I90674,I90362,I90705,I90359,I90736,I90753,I90770,I90787,I90804,I90821,I90386,I90852,I90374,I90368,I90897,I90914,I90383,I90945,I90962,I90979,I90371,I90356,I91057,I91074,I91091,I91108,I91028,I91139,I91156,I91173,I91190,I91207,I91224,I91241,I91258,I91275,I91292,I91043,I91040,I91337,I91025,I91368,I91022,I91399,I91416,I91433,I91450,I91467,I91484,I91049,I91515,I91037,I91031,I91560,I91577,I91046,I91608,I91625,I91642,I91034,I91019,I91720,I91737,I91754,I91771,I91691,I91802,I91819,I91836,I91853,I91870,I91887,I91904,I91921,I91938,I91955,I91706,I91703,I92000,I91688,I92031,I91685,I92062,I92079,I92096,I92113,I92130,I92147,I91712,I92178,I91700,I91694,I92223,I92240,I91709,I92271,I92288,I92305,I91697,I91682,I92383,I92400,I92417,I92357,I92448,I92465,I92482,I92499,I92516,I92533,I92550,I92567,I92584,I92351,I92615,I92632,I92348,I92663,I92680,I92697,I92360,I92345,I92742,I92759,I92776,I92793,I92810,I92366,I92841,I92375,I92872,I92369,I92372,I92363,I92354,I92978,I92995,I93012,I93029,I93046,I93063,I93080,I93097,I92967,I93128,I92952,I93159,I93176,I93193,I93210,I93227,I93244,I93261,I92949,I93292,I93309,I92946,I93340,I93357,I92964,I93388,I92961,I93419,I93436,I92940,I92943,I93481,I93498,I93515,I93532,I92970,I93563,I92955,I92958,I93641,I93658,I93675,I93692,I93709,I93726,I93743,I93760,I93630,I93791,I93615,I93822,I93839,I93856,I93873,I93890,I93907,I93924,I93612,I93955,I93972,I93609,I94003,I94020,I93627,I94051,I93624,I94082,I94099,I93603,I93606,I94144,I94161,I94178,I94195,I93633,I94226,I93618,I93621,I94304,I94321,I94338,I94355,I94372,I94389,I94406,I94275,I94437,I94454,I94471,I94488,I94505,I94522,I94539,I94272,I94570,I94266,I94601,I94618,I94635,I94296,I94269,I94680,I94293,I94711,I94290,I94287,I94756,I94773,I94790,I94807,I94824,I94281,I94855,I94872,I94284,I94278,I94950,I94967,I94984,I95001,I95018,I95035,I95052,I94921,I95083,I95100,I95117,I95134,I95151,I95168,I95185,I94918,I95216,I94912,I95247,I95264,I95281,I94942,I94915,I95326,I94939,I95357,I94936,I94933,I95402,I95419,I95436,I95453,I95470,I94927,I95501,I95518,I94930,I94924,I95596,I95613,I95630,I95647,I95664,I95681,I95698,I95567,I95729,I95746,I95763,I95780,I95797,I95814,I95831,I95564,I95862,I95558,I95893,I95910,I95927,I95588,I95561,I95972,I95585,I96003,I95582,I95579,I96048,I96065,I96082,I96099,I96116,I95573,I96147,I96164,I95576,I95570,I96242,I96259,I96276,I96293,I96310,I96327,I96344,I96213,I96375,I96392,I96409,I96426,I96443,I96460,I96477,I96210,I96508,I96204,I96539,I96556,I96573,I96234,I96207,I96618,I96231,I96649,I96228,I96225,I96694,I96711,I96728,I96745,I96762,I96219,I96793,I96810,I96222,I96216,I96888,I96905,I96922,I96939,I96956,I96973,I96990,I96859,I97021,I97038,I97055,I97072,I97089,I97106,I97123,I96856,I97154,I96850,I97185,I97202,I97219,I96880,I96853,I97264,I96877,I97295,I96874,I96871,I97340,I97357,I97374,I97391,I97408,I96865,I97439,I97456,I96868,I96862,I97534,I97551,I97568,I97585,I97602,I97502,I97633,I97650,I97667,I97505,I97698,I97499,I97729,I97746,I97763,I97780,I97797,I97508,I97828,I97845,I97862,I97879,I97514,I97517,I97496,I97938,I97955,I97972,I97526,I97523,I98017,I98034,I97511,I97520,I98112,I98129,I98146,I98163,I98180,I98080,I98211,I98228,I98245,I98083,I98276,I98077,I98307,I98324,I98341,I98358,I98375,I98086,I98406,I98423,I98440,I98457,I98092,I98095,I98074,I98516,I98533,I98550,I98104,I98101,I98595,I98612,I98089,I98098,I98690,I98707,I98724,I98741,I98758,I98658,I98789,I98806,I98823,I98840,I98857,I98874,I98891,I98908,I98664,I98655,I98953,I98970,I98679,I99001,I99018,I98667,I99049,I99066,I98673,I99097,I98661,I99128,I98652,I99159,I99176,I98682,I99207,I98676,I99238,I98670,I99302,I99319,I99336,I99353,I99291,I99384,I99401,I99418,I99435,I99452,I99469,I99486,I99276,I99517,I99273,I99548,I99285,I99579,I99596,I99613,I99279,I99294,I99658,I99675,I99264,I99706,I99282,I99737,I99754,I99288,I99785,I99802,I99267,I99270,I99880,I99897,I99914,I99931,I99948,I99965,I99863,I99996,I100013,I100030,I99866,I99848,I100075,I100092,I100109,I99869,I99860,I100154,I100171,I100188,I99851,I100219,I100236,I99842,I100267,I100284,I100301,I99872,I100332,I100349,I100366,I100383,I99857,I99854,I99845,I100475,I100492,I100509,I100526,I100543,I100560,I100458,I100591,I100608,I100625,I100461,I100443,I100670,I100687,I100704,I100464,I100455,I100749,I100766,I100783,I100446,I100814,I100831,I100437,I100862,I100879,I100896,I100467,I100927,I100944,I100961,I100978,I100452,I100449,I100440,I101070,I101087,I101104,I101121,I101138,I101155,I101053,I101186,I101203,I101220,I101056,I101038,I101265,I101282,I101299,I101059,I101050,I101344,I101361,I101378,I101041,I101409,I101426,I101032,I101457,I101474,I101491,I101062,I101522,I101539,I101556,I101573,I101047,I101044,I101035,I101665,I101682,I101699,I101716,I101733,I101750,I101648,I101781,I101798,I101815,I101651,I101633,I101860,I101877,I101894,I101654,I101645,I101939,I101956,I101973,I101636,I102004,I102021,I101627,I102052,I102069,I102086,I101657,I102117,I102134,I102151,I102168,I101642,I101639,I101630,I102260,I102277,I102294,I102311,I102328,I102345,I102243,I102376,I102393,I102410,I102246,I102228,I102455,I102472,I102489,I102249,I102240,I102534,I102551,I102568,I102231,I102599,I102616,I102222,I102647,I102664,I102681,I102252,I102712,I102729,I102746,I102763,I102237,I102234,I102225,I102855,I102872,I102889,I102906,I102923,I102940,I102957,I102826,I102988,I103005,I103022,I103039,I103056,I103073,I103090,I102823,I102817,I103135,I103152,I103169,I102844,I103200,I103217,I102835,I102829,I103262,I102832,I103293,I103310,I102847,I103341,I102841,I102838,I103386,I102820,I103450,I103467,I103484,I103501,I103518,I103535,I103552,I103421,I103583,I103600,I103617,I103634,I103651,I103668,I103685,I103418,I103412,I103730,I103747,I103764,I103439,I103795,I103812,I103430,I103424,I103857,I103427,I103888,I103905,I103442,I103936,I103436,I103433,I103981,I103415,I104045,I104062,I104079,I104096,I104113,I104130,I104147,I104164,I104181,I104198,I104215,I104232,I104249,I104266,I104034,I104297,I104314,I104331,I104007,I104362,I104028,I104393,I104410,I104013,I104441,I104010,I104016,I104486,I104503,I104520,I104022,I104037,I104025,I104579,I104596,I104031,I104019,I104674,I104691,I104708,I104725,I104742,I104759,I104776,I104793,I104810,I104827,I104844,I104861,I104878,I104895,I104663,I104926,I104943,I104960,I104636,I104991,I104657,I105022,I105039,I104642,I105070,I104639,I104645,I105115,I105132,I105149,I104651,I104666,I104654,I105208,I105225,I104660,I104648,I105303,I105320,I105337,I105354,I105371,I105388,I105405,I105422,I105439,I105456,I105473,I105490,I105507,I105524,I105292,I105555,I105572,I105589,I105265,I105620,I105286,I105651,I105668,I105271,I105699,I105268,I105274,I105744,I105761,I105778,I105280,I105295,I105283,I105837,I105854,I105289,I105277,I105932,I105949,I105966,I105983,I106000,I106017,I106034,I106051,I106068,I106085,I106102,I106119,I106136,I106153,I105921,I106184,I106201,I106218,I105894,I106249,I105915,I106280,I106297,I105900,I106328,I105897,I105903,I106373,I106390,I106407,I105909,I105924,I105912,I106466,I106483,I105918,I105906,I106561,I106578,I106595,I106612,I106550,I106643,I106538,I106674,I106691,I106708,I106725,I106742,I106541,I106773,I106526,I106804,I106821,I106838,I106855,I106872,I106889,I106532,I106920,I106937,I106954,I106544,I106553,I106523,I107013,I106547,I106535,I107058,I107075,I106529,I107139,I107156,I107173,I107190,I107128,I107221,I107116,I107252,I107269,I107286,I107303,I107320,I107119,I107351,I107104,I107382,I107399,I107416,I107433,I107450,I107467,I107110,I107498,I107515,I107532,I107122,I107131,I107101,I107591,I107125,I107113,I107636,I107653,I107107,I107717,I107734,I107751,I107768,I107706,I107799,I107694,I107830,I107847,I107864,I107881,I107898,I107697,I107929,I107682,I107960,I107977,I107994,I108011,I108028,I108045,I107688,I108076,I108093,I108110,I107700,I107709,I107679,I108169,I107703,I107691,I108214,I108231,I107685,I108295,I108312,I108329,I108346,I108363,I108380,I108278,I108266,I108425,I108442,I108459,I108476,I108493,I108275,I108524,I108541,I108558,I108575,I108284,I108263,I108620,I108637,I108281,I108668,I108272,I108287,I108713,I108730,I108747,I108764,I108260,I108269,I108257,I108856,I108873,I108890,I108907,I108830,I108938,I108955,I108845,I108827,I109000,I109017,I109034,I109051,I109068,I109085,I109102,I109119,I109136,I108842,I109167,I109184,I109201,I108824,I109232,I108821,I109263,I109280,I109297,I109314,I108836,I109345,I108833,I109376,I109393,I109410,I108839,I108848,I108818,I109502,I109519,I109536,I109553,I109476,I109584,I109601,I109491,I109473,I109646,I109663,I109680,I109697,I109714,I109731,I109748,I109765,I109782,I109488,I109813,I109830,I109847,I109470,I109878,I109467,I109909,I109926,I109943,I109960,I109482,I109991,I109479,I110022,I110039,I110056,I109485,I109494,I109464,I110148,I110165,I110182,I110199,I110122,I110230,I110247,I110137,I110119,I110292,I110309,I110326,I110343,I110360,I110377,I110394,I110411,I110428,I110134,I110459,I110476,I110493,I110116,I110524,I110113,I110555,I110572,I110589,I110606,I110128,I110637,I110125,I110668,I110685,I110702,I110131,I110140,I110110,I110794,I110811,I110828,I110845,I110765,I110876,I110893,I110910,I110927,I110944,I110961,I110978,I110995,I111012,I111029,I110780,I110777,I111074,I110762,I111105,I110759,I111136,I111153,I111170,I111187,I111204,I111221,I110786,I111252,I110774,I110768,I111297,I111314,I110783,I111345,I111362,I111379,I110771,I110756,I111457,I111474,I111491,I111508,I111428,I111539,I111556,I111573,I111590,I111607,I111624,I111641,I111658,I111675,I111692,I111443,I111440,I111737,I111425,I111768,I111422,I111799,I111816,I111833,I111850,I111867,I111884,I111449,I111915,I111437,I111431,I111960,I111977,I111446,I112008,I112025,I112042,I111434,I111419,I112120,I112137,I112154,I112171,I112091,I112202,I112219,I112236,I112253,I112270,I112287,I112304,I112321,I112338,I112355,I112106,I112103,I112400,I112088,I112431,I112085,I112462,I112479,I112496,I112513,I112530,I112547,I112112,I112578,I112100,I112094,I112623,I112640,I112109,I112671,I112688,I112705,I112097,I112082,I112783,I112800,I112817,I112834,I112754,I112865,I112882,I112899,I112916,I112933,I112950,I112967,I112984,I113001,I113018,I112769,I112766,I113063,I112751,I113094,I112748,I113125,I113142,I113159,I113176,I113193,I113210,I112775,I113241,I112763,I112757,I113286,I113303,I112772,I113334,I113351,I113368,I112760,I112745,I113446,I113463,I113480,I113497,I113417,I113528,I113545,I113562,I113579,I113596,I113613,I113630,I113647,I113664,I113681,I113432,I113429,I113726,I113414,I113757,I113411,I113788,I113805,I113822,I113839,I113856,I113873,I113438,I113904,I113426,I113420,I113949,I113966,I113435,I113997,I114014,I114031,I113423,I113408,I114109,I114126,I114143,I114174,I114191,I114208,I114225,I114242,I114259,I114276,I114293,I114310,I114341,I114358,I114389,I114406,I114423,I114468,I114485,I114502,I114519,I114536,I114567,I114598,I114704,I114721,I114687,I114666,I114766,I114783,I114800,I114817,I114834,I114851,I114868,I114885,I114902,I114693,I114933,I114950,I114967,I114984,I114696,I115015,I115032,I115049,I115066,I115083,I114681,I115114,I115131,I114684,I114678,I114672,I115190,I114690,I115221,I114675,I114669,I115299,I115316,I115282,I115261,I115361,I115378,I115395,I115412,I115429,I115446,I115463,I115480,I115497,I115288,I115528,I115545,I115562,I115579,I115291,I115610,I115627,I115644,I115661,I115678,I115276,I115709,I115726,I115279,I115273,I115267,I115785,I115285,I115816,I115270,I115264,I115894,I115911,I115928,I115945,I115962,I115979,I115996,I116013,I116044,I116075,I116092,I116109,I116126,I116143,I116160,I116177,I116208,I116225,I116256,I116273,I116304,I116335,I116352,I116397,I116414,I116431,I116448,I116479,I116557,I116574,I116591,I116608,I116625,I116642,I116659,I116676,I116546,I116707,I116531,I116738,I116755,I116772,I116789,I116806,I116823,I116840,I116528,I116871,I116888,I116525,I116919,I116936,I116543,I116967,I116540,I116998,I117015,I116519,I116522,I117060,I117077,I117094,I117111,I116549,I117142,I116534,I116537,I117220,I117237,I117254,I117271,I117288,I117305,I117322,I117339,I117370,I117401,I117418,I117435,I117452,I117469,I117486,I117503,I117534,I117551,I117582,I117599,I117630,I117661,I117678,I117723,I117740,I117757,I117774,I117805,I117883,I117900,I117917,I117934,I117951,I117968,I117985,I118002,I117872,I118033,I117857,I118064,I118081,I118098,I118115,I118132,I118149,I118166,I117854,I118197,I118214,I117851,I118245,I118262,I117869,I118293,I117866,I118324,I118341,I117845,I117848,I118386,I118403,I118420,I118437,I117875,I118468,I117860,I117863,I118546,I118563,I118580,I118597,I118614,I118631,I118648,I118665,I118535,I118696,I118520,I118727,I118744,I118761,I118778,I118795,I118812,I118829,I118517,I118860,I118877,I118514,I118908,I118925,I118532,I118956,I118529,I118987,I119004,I118508,I118511,I119049,I119066,I119083,I119100,I118538,I119131,I118523,I118526,I119209,I119226,I119243,I119260,I119277,I119294,I119311,I119180,I119342,I119359,I119376,I119393,I119410,I119427,I119444,I119177,I119475,I119171,I119506,I119523,I119540,I119201,I119174,I119585,I119198,I119616,I119195,I119192,I119661,I119678,I119695,I119712,I119729,I119186,I119760,I119777,I119189,I119183,I119855,I119872,I119889,I119906,I119923,I119817,I119954,I119971,I119988,I120005,I120022,I120039,I119826,I120070,I119820,I120101,I120118,I120135,I120152,I119847,I119844,I120197,I120214,I120231,I119841,I120262,I119838,I119829,I120307,I120324,I120341,I119832,I119835,I120386,I120403,I119823,I120467,I120484,I120501,I120518,I120535,I120435,I120566,I120583,I120600,I120438,I120631,I120432,I120662,I120679,I120696,I120713,I120730,I120441,I120761,I120778,I120795,I120812,I120447,I120450,I120429,I120871,I120888,I120905,I120459,I120456,I120950,I120967,I120444,I120453,I121045,I121062,I121079,I121096,I121113,I121144,I121161,I121178,I121209,I121240,I121257,I121274,I121291,I121308,I121339,I121356,I121373,I121390,I121449,I121466,I121483,I121528,I121545,I121623,I121640,I121657,I121674,I121691,I121722,I121739,I121756,I121787,I121818,I121835,I121852,I121869,I121886,I121917,I121934,I121951,I121968,I122027,I122044,I122061,I122106,I122123,I122201,I122218,I122235,I122252,I122269,I122169,I122300,I122317,I122334,I122172,I122365,I122166,I122396,I122413,I122430,I122447,I122464,I122175,I122495,I122512,I122529,I122546,I122181,I122184,I122163,I122605,I122622,I122639,I122193,I122190,I122684,I122701,I122178,I122187,I122779,I122796,I122813,I122830,I122861,I122878,I122895,I122912,I122929,I122946,I122963,I122994,I123025,I123056,I123073,I123090,I123135,I123152,I123183,I123214,I123231,I123262,I123279,I123357,I123374,I123391,I123408,I123425,I123442,I123340,I123473,I123490,I123507,I123343,I123325,I123552,I123569,I123586,I123346,I123337,I123631,I123648,I123665,I123328,I123696,I123713,I123319,I123744,I123761,I123778,I123349,I123809,I123826,I123843,I123860,I123334,I123331,I123322,I123952,I123969,I123986,I124003,I124020,I124037,I123935,I124068,I124085,I124102,I123938,I123920,I124147,I124164,I124181,I123941,I123932,I124226,I124243,I124260,I123923,I124291,I124308,I123914,I124339,I124356,I124373,I123944,I124404,I124421,I124438,I124455,I123929,I123926,I123917,I124547,I124564,I124581,I124598,I124615,I124632,I124530,I124663,I124680,I124697,I124533,I124515,I124742,I124759,I124776,I124536,I124527,I124821,I124838,I124855,I124518,I124886,I124903,I124509,I124934,I124951,I124968,I124539,I124999,I125016,I125033,I125050,I124524,I124521,I124512,I125142,I125159,I125176,I125193,I125210,I125227,I125244,I125113,I125275,I125292,I125309,I125326,I125343,I125360,I125377,I125110,I125104,I125422,I125439,I125456,I125131,I125487,I125504,I125122,I125116,I125549,I125119,I125580,I125597,I125134,I125628,I125128,I125125,I125673,I125107,I125737,I125754,I125771,I125788,I125805,I125822,I125839,I125708,I125870,I125887,I125904,I125921,I125938,I125955,I125972,I125705,I125699,I126017,I126034,I126051,I125726,I126082,I126099,I125717,I125711,I126144,I125714,I126175,I126192,I125729,I126223,I125723,I125720,I126268,I125702,I126332,I126349,I126366,I126383,I126400,I126417,I126434,I126303,I126465,I126482,I126499,I126516,I126533,I126550,I126567,I126300,I126294,I126612,I126629,I126646,I126321,I126677,I126694,I126312,I126306,I126739,I126309,I126770,I126787,I126324,I126818,I126318,I126315,I126863,I126297,I126927,I126944,I126961,I126978,I126995,I127012,I127029,I127046,I127063,I127080,I127097,I127114,I127131,I127148,I126916,I127179,I127196,I127213,I126889,I127244,I126910,I127275,I127292,I126895,I127323,I126892,I126898,I127368,I127385,I127402,I126904,I126919,I126907,I127461,I127478,I126913,I126901,I127556,I127573,I127590,I127607,I127545,I127638,I127533,I127669,I127686,I127703,I127720,I127737,I127536,I127768,I127521,I127799,I127816,I127833,I127850,I127867,I127884,I127527,I127915,I127932,I127949,I127539,I127548,I127518,I128008,I127542,I127530,I128053,I128070,I127524,I128134,I128151,I128168,I128185,I128123,I128216,I128111,I128247,I128264,I128281,I128298,I128315,I128114,I128346,I128099,I128377,I128394,I128411,I128428,I128445,I128462,I128105,I128493,I128510,I128527,I128117,I128126,I128096,I128586,I128120,I128108,I128631,I128648,I128102,I128712,I128729,I128746,I128763,I128701,I128794,I128689,I128825,I128842,I128859,I128876,I128893,I128692,I128924,I128677,I128955,I128972,I128989,I129006,I129023,I129040,I128683,I129071,I129088,I129105,I128695,I128704,I128674,I129164,I128698,I128686,I129209,I129226,I128680,I129290,I129307,I129324,I129341,I129358,I129375,I129420,I129437,I129454,I129471,I129488,I129519,I129536,I129553,I129570,I129615,I129632,I129663,I129708,I129725,I129742,I129759,I129851,I129868,I129885,I129902,I129919,I129936,I129834,I129822,I129981,I129998,I130015,I130032,I130049,I129831,I130080,I130097,I130114,I130131,I129840,I129819,I130176,I130193,I129837,I130224,I129828,I129843,I130269,I130286,I130303,I130320,I129816,I129825,I129813,I130412,I130429,I130446,I130463,I130480,I130497,I130395,I130383,I130542,I130559,I130576,I130593,I130610,I130392,I130641,I130658,I130675,I130692,I130401,I130380,I130737,I130754,I130398,I130785,I130389,I130404,I130830,I130847,I130864,I130881,I130377,I130386,I130374,I130973,I130990,I131007,I131024,I130947,I131055,I131072,I130962,I130944,I131117,I131134,I131151,I131168,I131185,I131202,I131219,I131236,I131253,I130959,I131284,I131301,I131318,I130941,I131349,I130938,I131380,I131397,I131414,I131431,I130953,I131462,I130950,I131493,I131510,I131527,I130956,I130965,I130935,I131619,I131636,I131653,I131670,I131590,I131701,I131718,I131735,I131752,I131769,I131786,I131803,I131820,I131837,I131854,I131605,I131602,I131899,I131587,I131930,I131584,I131961,I131978,I131995,I132012,I132029,I132046,I131611,I132077,I131599,I131593,I132122,I132139,I131608,I132170,I132187,I132204,I131596,I131581,I132282,I132299,I132316,I132333,I132253,I132364,I132381,I132398,I132415,I132432,I132449,I132466,I132483,I132500,I132517,I132268,I132265,I132562,I132250,I132593,I132247,I132624,I132641,I132658,I132675,I132692,I132709,I132274,I132740,I132262,I132256,I132785,I132802,I132271,I132833,I132850,I132867,I132259,I132244,I132945,I132962,I132979,I132996,I133027,I133044,I133061,I133078,I133095,I133112,I133129,I133146,I133163,I133180,I133225,I133256,I133287,I133304,I133321,I133338,I133355,I133372,I133403,I133448,I133465,I133496,I133513,I133530,I133608,I133625,I133642,I133582,I133673,I133690,I133707,I133724,I133741,I133758,I133775,I133792,I133809,I133576,I133840,I133857,I133573,I133888,I133905,I133922,I133585,I133570,I133967,I133984,I134001,I134018,I134035,I133591,I134066,I133600,I134097,I133594,I133597,I133588,I133579,I134203,I134220,I134237,I134268,I134285,I134302,I134319,I134336,I134353,I134370,I134387,I134404,I134435,I134452,I134483,I134500,I134517,I134562,I134579,I134596,I134613,I134630,I134661,I134692,I134798,I134815,I134832,I134849,I134866,I134883,I134900,I134917,I134948,I134979,I134996,I135013,I135030,I135047,I135064,I135081,I135112,I135129,I135160,I135177,I135208,I135239,I135256,I135301,I135318,I135335,I135352,I135383,I135461,I135478,I135495,I135512,I135529,I135546,I135563,I135580,I135450,I135611,I135435,I135642,I135659,I135676,I135693,I135710,I135727,I135744,I135432,I135775,I135792,I135429,I135823,I135840,I135447,I135871,I135444,I135902,I135919,I135423,I135426,I135964,I135981,I135998,I136015,I135453,I136046,I135438,I135441,I136124,I136141,I136158,I136175,I136192,I136209,I136226,I136243,I136113,I136274,I136098,I136305,I136322,I136339,I136356,I136373,I136390,I136407,I136095,I136438,I136455,I136092,I136486,I136503,I136110,I136534,I136107,I136565,I136582,I136086,I136089,I136627,I136644,I136661,I136678,I136116,I136709,I136101,I136104,I136787,I136804,I136821,I136838,I136855,I136872,I136889,I136906,I136776,I136937,I136761,I136968,I136985,I137002,I137019,I137036,I137053,I137070,I136758,I137101,I137118,I136755,I137149,I137166,I136773,I137197,I136770,I137228,I137245,I136749,I136752,I137290,I137307,I137324,I137341,I136779,I137372,I136764,I136767,I137450,I137467,I137484,I137501,I137518,I137535,I137552,I137569,I137439,I137600,I137424,I137631,I137648,I137665,I137682,I137699,I137716,I137733,I137421,I137764,I137781,I137418,I137812,I137829,I137436,I137860,I137433,I137891,I137908,I137412,I137415,I137953,I137970,I137987,I138004,I137442,I138035,I137427,I137430,I138113,I138130,I138147,I138164,I138181,I138198,I138215,I138232,I138102,I138263,I138087,I138294,I138311,I138328,I138345,I138362,I138379,I138396,I138084,I138427,I138444,I138081,I138475,I138492,I138099,I138523,I138096,I138554,I138571,I138075,I138078,I138616,I138633,I138650,I138667,I138105,I138698,I138090,I138093,I138776,I138793,I138810,I138827,I138844,I138861,I138878,I138747,I138909,I138926,I138943,I138960,I138977,I138994,I139011,I138744,I139042,I138738,I139073,I139090,I139107,I138768,I138741,I139152,I138765,I139183,I138762,I138759,I139228,I139245,I139262,I139279,I139296,I138753,I139327,I139344,I138756,I138750,I139422,I139439,I139456,I139473,I139490,I139507,I139524,I139393,I139555,I139572,I139589,I139606,I139623,I139640,I139657,I139390,I139688,I139384,I139719,I139736,I139753,I139414,I139387,I139798,I139411,I139829,I139408,I139405,I139874,I139891,I139908,I139925,I139942,I139399,I139973,I139990,I139402,I139396,I140068,I140085,I140102,I140119,I140136,I140153,I140170,I140039,I140201,I140218,I140235,I140252,I140269,I140286,I140303,I140036,I140334,I140030,I140365,I140382,I140399,I140060,I140033,I140444,I140057,I140475,I140054,I140051,I140520,I140537,I140554,I140571,I140588,I140045,I140619,I140636,I140048,I140042,I140714,I140731,I140748,I140765,I140782,I140682,I140813,I140830,I140847,I140685,I140878,I140679,I140909,I140926,I140943,I140960,I140977,I140688,I141008,I141025,I141042,I141059,I140694,I140697,I140676,I141118,I141135,I141152,I140706,I140703,I141197,I141214,I140691,I140700,I141292,I141309,I141326,I141343,I141360,I141260,I141391,I141408,I141425,I141263,I141456,I141257,I141487,I141504,I141521,I141538,I141555,I141266,I141586,I141603,I141620,I141637,I141272,I141275,I141254,I141696,I141713,I141730,I141284,I141281,I141775,I141792,I141269,I141278,I141870,I141887,I141904,I141921,I141938,I141955,I141986,I142003,I142020,I142065,I142082,I142099,I142144,I142161,I142178,I142209,I142226,I142257,I142274,I142291,I142322,I142339,I142356,I142373,I142465,I142482,I142499,I142516,I142533,I142550,I142567,I142598,I142615,I142632,I142649,I142666,I142683,I142700,I142745,I142762,I142779,I142810,I142827,I142872,I142903,I142920,I142951,I142996,I143060,I143077,I143094,I143111,I143049,I143142,I143037,I143173,I143190,I143207,I143224,I143241,I143040,I143272,I143025,I143303,I143320,I143337,I143354,I143371,I143388,I143031,I143419,I143436,I143453,I143043,I143052,I143022,I143512,I143046,I143034,I143557,I143574,I143028,I143638,I143655,I143672,I143689,I143706,I143723,I143768,I143785,I143802,I143819,I143836,I143867,I143884,I143901,I143918,I143963,I143980,I144011,I144056,I144073,I144090,I144107,I144199,I144216,I144233,I144250,I144267,I144284,I144182,I144170,I144329,I144346,I144363,I144380,I144397,I144179,I144428,I144445,I144462,I144479,I144188,I144167,I144524,I144541,I144185,I144572,I144176,I144191,I144617,I144634,I144651,I144668,I144164,I144173,I144161,I144760,I144777,I144794,I144811,I144828,I144845,I144743,I144731,I144890,I144907,I144924,I144941,I144958,I144740,I144989,I145006,I145023,I145040,I144749,I144728,I145085,I145102,I144746,I145133,I144737,I144752,I145178,I145195,I145212,I145229,I144725,I144734,I144722,I145321,I145338,I145355,I145372,I145403,I145420,I145465,I145482,I145499,I145516,I145533,I145550,I145567,I145584,I145601,I145632,I145649,I145666,I145697,I145728,I145745,I145762,I145779,I145810,I145841,I145858,I145875,I145967,I145984,I146001,I146018,I146049,I146066,I146111,I146128,I146145,I146162,I146179,I146196,I146213,I146230,I146247,I146278,I146295,I146312,I146343,I146374,I146391,I146408,I146425,I146456,I146487,I146504,I146521,I146613,I146630,I146647,I146678,I146695,I146712,I146729,I146746,I146763,I146780,I146797,I146814,I146845,I146862,I146893,I146910,I146927,I146972,I146989,I147006,I147023,I147040,I147071,I147102,I147208,I147225,I147242,I147259,I147276,I147293,I147310,I147327,I147197,I147358,I147182,I147389,I147406,I147423,I147440,I147457,I147474,I147491,I147179,I147522,I147539,I147176,I147570,I147587,I147194,I147618,I147191,I147649,I147666,I147170,I147173,I147711,I147728,I147745,I147762,I147200,I147793,I147185,I147188,I147871,I147888,I147905,I147922,I147939,I147956,I147973,I147842,I148004,I148021,I148038,I148055,I148072,I148089,I148106,I147839,I148137,I147833,I148168,I148185,I148202,I147863,I147836,I148247,I147860,I148278,I147857,I147854,I148323,I148340,I148357,I148374,I148391,I147848,I148422,I148439,I147851,I147845,I148517,I148534,I148551,I148568,I148585,I148485,I148616,I148633,I148650,I148488,I148681,I148482,I148712,I148729,I148746,I148763,I148780,I148491,I148811,I148828,I148845,I148862,I148497,I148500,I148479,I148921,I148938,I148955,I148509,I148506,I149000,I149017,I148494,I148503,I149095,I149112,I149129,I149146,I149163,I149180,I149197,I149214,I149231,I149248,I149265,I149282,I149299,I149316,I149347,I149364,I149381,I149412,I149443,I149460,I149491,I149536,I149553,I149570,I149629,I149646,I149724,I149741,I149758,I149775,I149806,I149837,I149854,I149871,I149888,I149905,I149936,I149967,I149984,I150001,I150018,I150035,I150052,I150083,I150100,I150117,I150176,I150221,I150238,I150302,I150319,I150336,I150353,I150370,I150387,I150432,I150449,I150466,I150483,I150500,I150531,I150548,I150565,I150582,I150627,I150644,I150675,I150720,I150737,I150754,I150771,I150863,I150880,I150897,I150914,I150931,I150948,I150965,I150982,I151013,I151044,I151061,I151078,I151095,I151112,I151129,I151146,I151177,I151194,I151225,I151242,I151273,I151304,I151321,I151366,I151383,I151400,I151417,I151448;
not I_0 (I3014,I2973);
nand I_1 (I3031,I1847,I2799);
and I_2 (I3048,I3031,I1447);
DFFARX1 I_3 (I3065,I3048,I2966,I3014,);
not I_4 (I3082,I3065);
nor I_5 (I3099,I2111,I2799);
or I_6 (I2997,I3099,I3065);
not I_7 (I2985,I3099);
DFFARX1 I_8 (I3144,I1375,I2966,I3014,);
nor I_9 (I3161,I3144,I3099);
nand I_10 (I3178,I1367,I1991);
and I_11 (I3195,I3178,I1663);
DFFARX1 I_12 (I3212,I3195,I2966,I3014,);
nor I_13 (I2994,I3212,I3065);
not I_14 (I3243,I3212);
nor I_15 (I3260,I3144,I3243);
DFFARX1 I_16 (I3277,I1575,I2966,I3014,);
and I_17 (I3294,I3277,I2943);
or I_18 (I3003,I3294,I3099);
nand I_19 (I2982,I3294,I3260);
DFFARX1 I_20 (I3339,I2079,I2966,I3014,);
and I_21 (I3356,I3339,I3082);
nor I_22 (I3000,I3294,I3356);
nor I_23 (I3387,I3339,I3144);
DFFARX1 I_24 (I2991,I3387,I2966,I3014,);
nor I_25 (I3006,I3339,I3065);
not I_26 (I3432,I3339);
nor I_27 (I3449,I3212,I3432);
and I_28 (I3466,I3099,I3449);
or I_29 (I3483,I3294,I3466);
DFFARX1 I_30 (I2979,I3483,I2966,I3014,);
nand I_31 (I2988,I3339,I3161);
nand I_32 (I2976,I3339,I3243);
not I_33 (I3575,I2973);
nand I_34 (I3592,I1927,I2599);
and I_35 (I3609,I3592,I1879);
DFFARX1 I_36 (I3626,I3609,I2966,I3575,);
not I_37 (I3643,I3626);
nor I_38 (I3660,I2583,I2599);
or I_39 (I3558,I3660,I3626);
not I_40 (I3546,I3660);
DFFARX1 I_41 (I3705,I2127,I2966,I3575,);
nor I_42 (I3722,I3705,I3660);
nand I_43 (I3739,I2687,I2119);
and I_44 (I3756,I3739,I1623);
DFFARX1 I_45 (I3773,I3756,I2966,I3575,);
nor I_46 (I3555,I3773,I3626);
not I_47 (I3804,I3773);
nor I_48 (I3821,I3705,I3804);
DFFARX1 I_49 (I3838,I2463,I2966,I3575,);
and I_50 (I3855,I3838,I2199);
or I_51 (I3564,I3855,I3660);
nand I_52 (I3543,I3855,I3821);
DFFARX1 I_53 (I3900,I2143,I2966,I3575,);
and I_54 (I3917,I3900,I3643);
nor I_55 (I3561,I3855,I3917);
nor I_56 (I3948,I3900,I3705);
DFFARX1 I_57 (I3552,I3948,I2966,I3575,);
nor I_58 (I3567,I3900,I3626);
not I_59 (I3993,I3900);
nor I_60 (I4010,I3773,I3993);
and I_61 (I4027,I3660,I4010);
or I_62 (I4044,I3855,I4027);
DFFARX1 I_63 (I3540,I4044,I2966,I3575,);
nand I_64 (I3549,I3900,I3722);
nand I_65 (I3537,I3900,I3804);
not I_66 (I4136,I2973);
nand I_67 (I4153,I2887,I1951);
and I_68 (I4170,I4153,I2207);
DFFARX1 I_69 (I4187,I4170,I2966,I4136,);
not I_70 (I4204,I4187);
nor I_71 (I4221,I2055,I1951);
or I_72 (I4119,I4221,I4187);
not I_73 (I4107,I4221);
DFFARX1 I_74 (I4266,I1271,I2966,I4136,);
nor I_75 (I4283,I4266,I4221);
nand I_76 (I4300,I2623,I2431);
and I_77 (I4317,I4300,I2719);
DFFARX1 I_78 (I4334,I4317,I2966,I4136,);
nor I_79 (I4116,I4334,I4187);
not I_80 (I4365,I4334);
nor I_81 (I4382,I4266,I4365);
DFFARX1 I_82 (I4399,I2479,I2966,I4136,);
and I_83 (I4416,I4399,I2727);
or I_84 (I4125,I4416,I4221);
nand I_85 (I4104,I4416,I4382);
DFFARX1 I_86 (I4461,I1911,I2966,I4136,);
and I_87 (I4478,I4461,I4204);
nor I_88 (I4122,I4416,I4478);
nor I_89 (I4509,I4461,I4266);
DFFARX1 I_90 (I4113,I4509,I2966,I4136,);
nor I_91 (I4128,I4461,I4187);
not I_92 (I4554,I4461);
nor I_93 (I4571,I4334,I4554);
and I_94 (I4588,I4221,I4571);
or I_95 (I4605,I4416,I4588);
DFFARX1 I_96 (I4101,I4605,I2966,I4136,);
nand I_97 (I4110,I4461,I4283);
nand I_98 (I4098,I4461,I4365);
not I_99 (I4697,I2973);
not I_100 (I4714,I2359);
nor I_101 (I4731,I1407,I2575);
nand I_102 (I4748,I4731,I2487);
DFFARX1 I_103 (I4671,I4748,I2966,I4697,);
nor I_104 (I4779,I4714,I1407);
nand I_105 (I4796,I4779,I1535);
not I_106 (I4686,I4796);
DFFARX1 I_107 (I4668,I4796,I2966,I4697,);
not I_108 (I4841,I1407);
not I_109 (I4858,I4841);
not I_110 (I4875,I2927);
nor I_111 (I4892,I4875,I1783);
and I_112 (I4909,I4892,I1759);
or I_113 (I4926,I4909,I2679);
DFFARX1 I_114 (I4943,I4926,I2966,I4697,);
nor I_115 (I4960,I4943,I4796);
nor I_116 (I4977,I4943,I4858);
nand I_117 (I4683,I4748,I4977);
nand I_118 (I5008,I4714,I2927);
nand I_119 (I5025,I5008,I4943);
and I_120 (I5042,I5008,I5025);
DFFARX1 I_121 (I4665,I5042,I2966,I4697,);
DFFARX1 I_122 (I5073,I5008,I2966,I4697,);
and I_123 (I4662,I4841,I5073);
DFFARX1 I_124 (I5104,I2471,I2966,I4697,);
not I_125 (I5121,I5104);
nor I_126 (I5138,I4796,I5121);
and I_127 (I5155,I5104,I5138);
nand I_128 (I4677,I5104,I4858);
DFFARX1 I_129 (I5186,I5104,I2966,I4697,);
not I_130 (I4674,I5186);
DFFARX1 I_131 (I5217,I2255,I2966,I4697,);
not I_132 (I5234,I5217);
or I_133 (I5251,I5234,I5155);
DFFARX1 I_134 (I4680,I5251,I2966,I4697,);
nand I_135 (I4689,I5234,I4960);
DFFARX1 I_136 (I4659,I5234,I2966,I4697,);
not I_137 (I5343,I2973);
not I_138 (I5360,I2175);
nor I_139 (I5377,I2423,I2071);
nand I_140 (I5394,I5377,I1263);
DFFARX1 I_141 (I5317,I5394,I2966,I5343,);
nor I_142 (I5425,I5360,I2423);
nand I_143 (I5442,I5425,I2407);
not I_144 (I5332,I5442);
DFFARX1 I_145 (I5314,I5442,I2966,I5343,);
not I_146 (I5487,I2423);
not I_147 (I5504,I5487);
not I_148 (I5521,I1431);
nor I_149 (I5538,I5521,I2063);
and I_150 (I5555,I5538,I2863);
or I_151 (I5572,I5555,I2783);
DFFARX1 I_152 (I5589,I5572,I2966,I5343,);
nor I_153 (I5606,I5589,I5442);
nor I_154 (I5623,I5589,I5504);
nand I_155 (I5329,I5394,I5623);
nand I_156 (I5654,I5360,I1431);
nand I_157 (I5671,I5654,I5589);
and I_158 (I5688,I5654,I5671);
DFFARX1 I_159 (I5311,I5688,I2966,I5343,);
DFFARX1 I_160 (I5719,I5654,I2966,I5343,);
and I_161 (I5308,I5487,I5719);
DFFARX1 I_162 (I5750,I2895,I2966,I5343,);
not I_163 (I5767,I5750);
nor I_164 (I5784,I5442,I5767);
and I_165 (I5801,I5750,I5784);
nand I_166 (I5323,I5750,I5504);
DFFARX1 I_167 (I5832,I5750,I2966,I5343,);
not I_168 (I5320,I5832);
DFFARX1 I_169 (I5863,I1719,I2966,I5343,);
not I_170 (I5880,I5863);
or I_171 (I5897,I5880,I5801);
DFFARX1 I_172 (I5326,I5897,I2966,I5343,);
nand I_173 (I5335,I5880,I5606);
DFFARX1 I_174 (I5305,I5880,I2966,I5343,);
not I_175 (I5989,I2973);
not I_176 (I6006,I1607);
nor I_177 (I6023,I1359,I1871);
nand I_178 (I6040,I6023,I1727);
DFFARX1 I_179 (I5960,I6040,I2966,I5989,);
nor I_180 (I6071,I6006,I1359);
nand I_181 (I6088,I6071,I2263);
nand I_182 (I6105,I6088,I6040);
not I_183 (I6122,I1359);
not I_184 (I6139,I2543);
nor I_185 (I6156,I6139,I1943);
and I_186 (I6173,I6156,I2039);
or I_187 (I6190,I6173,I1775);
DFFARX1 I_188 (I6207,I6190,I2966,I5989,);
nor I_189 (I6224,I6207,I6088);
nand I_190 (I5975,I6122,I6224);
not I_191 (I5972,I6207);
and I_192 (I6269,I6207,I6105);
DFFARX1 I_193 (I5957,I6269,I2966,I5989,);
DFFARX1 I_194 (I6300,I6207,I2966,I5989,);
and I_195 (I5954,I6122,I6300);
nand I_196 (I6331,I6006,I2543);
not I_197 (I6348,I6331);
nor I_198 (I6365,I6207,I6348);
DFFARX1 I_199 (I6382,I2271,I2966,I5989,);
nand I_200 (I6399,I6382,I6331);
and I_201 (I6416,I6122,I6399);
DFFARX1 I_202 (I5981,I6416,I2966,I5989,);
not I_203 (I6447,I6382);
nand I_204 (I5969,I6382,I6365);
nand I_205 (I5963,I6382,I6348);
DFFARX1 I_206 (I6492,I1415,I2966,I5989,);
not I_207 (I6509,I6492);
nor I_208 (I5978,I6382,I6509);
nor I_209 (I6540,I6509,I6447);
and I_210 (I6557,I6088,I6540);
or I_211 (I6574,I6331,I6557);
DFFARX1 I_212 (I5966,I6574,I2966,I5989,);
DFFARX1 I_213 (I5951,I6509,I2966,I5989,);
not I_214 (I6652,I2973);
or I_215 (I6669,I1807,I1543);
not I_216 (I6635,I6669);
DFFARX1 I_217 (I6614,I6669,I2966,I6652,);
or I_218 (I6714,I2375,I1807);
nor I_219 (I6731,I1591,I1711);
nor I_220 (I6748,I6731,I6669);
not I_221 (I6765,I1591);
and I_222 (I6782,I6765,I2751);
nor I_223 (I6799,I6782,I1543);
DFFARX1 I_224 (I6816,I6799,I2966,I6652,);
nor I_225 (I6833,I1503,I1479);
DFFARX1 I_226 (I6850,I6833,I2966,I6652,);
nor I_227 (I6641,I6850,I6799);
not I_228 (I6881,I6850);
nor I_229 (I6898,I1503,I2375);
nand I_230 (I6915,I6799,I6898);
and I_231 (I6932,I6714,I6915);
DFFARX1 I_232 (I6644,I6932,I2966,I6652,);
DFFARX1 I_233 (I6963,I2855,I2966,I6652,);
and I_234 (I6980,I6963,I1439);
nor I_235 (I6997,I6980,I6881);
and I_236 (I7014,I6898,I6997);
or I_237 (I7031,I6731,I7014);
DFFARX1 I_238 (I6629,I7031,I2966,I6652,);
not I_239 (I7062,I6980);
nor I_240 (I7079,I6669,I7062);
nand I_241 (I6632,I6714,I7079);
nand I_242 (I6626,I6850,I7062);
DFFARX1 I_243 (I6620,I6980,I2966,I6652,);
DFFARX1 I_244 (I7138,I1735,I2966,I6652,);
nand I_245 (I6638,I7138,I6748);
DFFARX1 I_246 (I7169,I7138,I2966,I6652,);
not I_247 (I6623,I7169);
and I_248 (I6617,I7138,I6816);
not I_249 (I7247,I2973);
not I_250 (I7264,I2959);
nor I_251 (I7281,I1935,I2247);
nand I_252 (I7298,I7281,I2439);
nor I_253 (I7315,I7264,I1935);
nand I_254 (I7332,I7315,I2815);
not I_255 (I7349,I7332);
not I_256 (I7366,I1935);
nor I_257 (I7236,I7332,I7366);
not I_258 (I7397,I7366);
nand I_259 (I7221,I7332,I7397);
not I_260 (I7428,I2335);
nor I_261 (I7445,I7428,I1743);
and I_262 (I7462,I7445,I1255);
or I_263 (I7479,I7462,I2831);
DFFARX1 I_264 (I7496,I7479,I2966,I7247,);
nor I_265 (I7513,I7496,I7349);
DFFARX1 I_266 (I7530,I7496,I2966,I7247,);
not I_267 (I7218,I7530);
nand I_268 (I7561,I7264,I2335);
and I_269 (I7578,I7561,I7513);
DFFARX1 I_270 (I7215,I7561,I2966,I7247,);
DFFARX1 I_271 (I7609,I2343,I2966,I7247,);
nor I_272 (I7626,I7609,I7332);
nand I_273 (I7233,I7496,I7626);
nor I_274 (I7657,I7609,I7397);
not I_275 (I7230,I7609);
nand I_276 (I7688,I7609,I7298);
and I_277 (I7705,I7366,I7688);
DFFARX1 I_278 (I7209,I7705,I2966,I7247,);
DFFARX1 I_279 (I7212,I7609,I2966,I7247,);
DFFARX1 I_280 (I7750,I2511,I2966,I7247,);
not I_281 (I7767,I7750);
nand I_282 (I7784,I7767,I7332);
and I_283 (I7801,I7561,I7784);
DFFARX1 I_284 (I7239,I7801,I2966,I7247,);
or I_285 (I7832,I7767,I7578);
DFFARX1 I_286 (I7224,I7832,I2966,I7247,);
nand I_287 (I7227,I7767,I7657);
not I_288 (I7910,I2973);
not I_289 (I7927,I1855);
nor I_290 (I7944,I1799,I1559);
nand I_291 (I7961,I7944,I2695);
nor I_292 (I7978,I7927,I1799);
nand I_293 (I7995,I7978,I1687);
not I_294 (I8012,I7995);
not I_295 (I8029,I1799);
nor I_296 (I7899,I7995,I8029);
not I_297 (I8060,I8029);
nand I_298 (I7884,I7995,I8060);
not I_299 (I8091,I1703);
nor I_300 (I8108,I8091,I2527);
and I_301 (I8125,I8108,I1207);
or I_302 (I8142,I8125,I2295);
DFFARX1 I_303 (I8159,I8142,I2966,I7910,);
nor I_304 (I8176,I8159,I8012);
DFFARX1 I_305 (I8193,I8159,I2966,I7910,);
not I_306 (I7881,I8193);
nand I_307 (I8224,I7927,I1703);
and I_308 (I8241,I8224,I8176);
DFFARX1 I_309 (I7878,I8224,I2966,I7910,);
DFFARX1 I_310 (I8272,I2911,I2966,I7910,);
nor I_311 (I8289,I8272,I7995);
nand I_312 (I7896,I8159,I8289);
nor I_313 (I8320,I8272,I8060);
not I_314 (I7893,I8272);
nand I_315 (I8351,I8272,I7961);
and I_316 (I8368,I8029,I8351);
DFFARX1 I_317 (I7872,I8368,I2966,I7910,);
DFFARX1 I_318 (I7875,I8272,I2966,I7910,);
DFFARX1 I_319 (I8413,I2351,I2966,I7910,);
not I_320 (I8430,I8413);
nand I_321 (I8447,I8430,I7995);
and I_322 (I8464,I8224,I8447);
DFFARX1 I_323 (I7902,I8464,I2966,I7910,);
or I_324 (I8495,I8430,I8241);
DFFARX1 I_325 (I7887,I8495,I2966,I7910,);
nand I_326 (I7890,I8430,I8320);
not I_327 (I8573,I2973);
not I_328 (I8590,I1351);
nor I_329 (I8607,I1471,I2807);
nand I_330 (I8624,I8607,I1455);
nor I_331 (I8641,I8590,I1471);
nand I_332 (I8658,I8641,I1831);
not I_333 (I8675,I8658);
not I_334 (I8692,I1471);
nor I_335 (I8562,I8658,I8692);
not I_336 (I8723,I8692);
nand I_337 (I8547,I8658,I8723);
not I_338 (I8754,I1303);
nor I_339 (I8771,I8754,I2663);
and I_340 (I8788,I8771,I2759);
or I_341 (I8805,I8788,I1919);
DFFARX1 I_342 (I8822,I8805,I2966,I8573,);
nor I_343 (I8839,I8822,I8675);
DFFARX1 I_344 (I8856,I8822,I2966,I8573,);
not I_345 (I8544,I8856);
nand I_346 (I8887,I8590,I1303);
and I_347 (I8904,I8887,I8839);
DFFARX1 I_348 (I8541,I8887,I2966,I8573,);
DFFARX1 I_349 (I8935,I2015,I2966,I8573,);
nor I_350 (I8952,I8935,I8658);
nand I_351 (I8559,I8822,I8952);
nor I_352 (I8983,I8935,I8723);
not I_353 (I8556,I8935);
nand I_354 (I9014,I8935,I8624);
and I_355 (I9031,I8692,I9014);
DFFARX1 I_356 (I8535,I9031,I2966,I8573,);
DFFARX1 I_357 (I8538,I8935,I2966,I8573,);
DFFARX1 I_358 (I9076,I1423,I2966,I8573,);
not I_359 (I9093,I9076);
nand I_360 (I9110,I9093,I8658);
and I_361 (I9127,I8887,I9110);
DFFARX1 I_362 (I8565,I9127,I2966,I8573,);
or I_363 (I9158,I9093,I8904);
DFFARX1 I_364 (I8550,I9158,I2966,I8573,);
nand I_365 (I8553,I9093,I8983);
not I_366 (I9236,I2973);
not I_367 (I9253,I2231);
nor I_368 (I9270,I2903,I1655);
nand I_369 (I9287,I9270,I2191);
nor I_370 (I9304,I9253,I2903);
nand I_371 (I9321,I9304,I2655);
not I_372 (I9338,I9321);
not I_373 (I9355,I2903);
nor I_374 (I9225,I9321,I9355);
not I_375 (I9386,I9355);
nand I_376 (I9210,I9321,I9386);
not I_377 (I9417,I1343);
nor I_378 (I9434,I9417,I2607);
and I_379 (I9451,I9434,I2775);
or I_380 (I9468,I9451,I2503);
DFFARX1 I_381 (I9485,I9468,I2966,I9236,);
nor I_382 (I9502,I9485,I9338);
DFFARX1 I_383 (I9519,I9485,I2966,I9236,);
not I_384 (I9207,I9519);
nand I_385 (I9550,I9253,I1343);
and I_386 (I9567,I9550,I9502);
DFFARX1 I_387 (I9204,I9550,I2966,I9236,);
DFFARX1 I_388 (I9598,I2303,I2966,I9236,);
nor I_389 (I9615,I9598,I9321);
nand I_390 (I9222,I9485,I9615);
nor I_391 (I9646,I9598,I9386);
not I_392 (I9219,I9598);
nand I_393 (I9677,I9598,I9287);
and I_394 (I9694,I9355,I9677);
DFFARX1 I_395 (I9198,I9694,I2966,I9236,);
DFFARX1 I_396 (I9201,I9598,I2966,I9236,);
DFFARX1 I_397 (I9739,I2167,I2966,I9236,);
not I_398 (I9756,I9739);
nand I_399 (I9773,I9756,I9321);
and I_400 (I9790,I9550,I9773);
DFFARX1 I_401 (I9228,I9790,I2966,I9236,);
or I_402 (I9821,I9756,I9567);
DFFARX1 I_403 (I9213,I9821,I2966,I9236,);
nand I_404 (I9216,I9756,I9646);
not I_405 (I9899,I2973);
not I_406 (I9916,I1751);
nor I_407 (I9933,I2047,I2287);
nand I_408 (I9950,I9933,I2951);
nor I_409 (I9967,I9916,I2047);
nand I_410 (I9984,I9967,I1679);
DFFARX1 I_411 (I10001,I9984,I2966,I9899,);
not I_412 (I9870,I10001);
not I_413 (I10032,I2047);
not I_414 (I10049,I10032);
not I_415 (I10066,I2711);
nor I_416 (I10083,I10066,I2455);
and I_417 (I10100,I10083,I2767);
or I_418 (I10117,I10100,I2239);
DFFARX1 I_419 (I10134,I10117,I2966,I9899,);
DFFARX1 I_420 (I9867,I10134,I2966,I9899,);
DFFARX1 I_421 (I10165,I10134,I2966,I9899,);
DFFARX1 I_422 (I9861,I10134,I2966,I9899,);
nand I_423 (I10196,I9916,I2711);
nand I_424 (I10213,I10196,I9950);
and I_425 (I10230,I10032,I10213);
DFFARX1 I_426 (I9891,I10230,I2966,I9899,);
and I_427 (I9864,I10196,I10165);
DFFARX1 I_428 (I10275,I1887,I2966,I9899,);
nor I_429 (I9888,I10275,I10196);
nor I_430 (I10306,I10275,I9950);
nand I_431 (I9885,I9984,I10306);
not I_432 (I9882,I10275);
DFFARX1 I_433 (I10351,I1999,I2966,I9899,);
not I_434 (I10368,I10351);
nor I_435 (I10385,I10368,I10049);
and I_436 (I10402,I10275,I10385);
or I_437 (I10419,I10196,I10402);
DFFARX1 I_438 (I9876,I10419,I2966,I9899,);
not I_439 (I10450,I10368);
nor I_440 (I10467,I10275,I10450);
nand I_441 (I9879,I10368,I10467);
nand I_442 (I9873,I10032,I10450);
not I_443 (I10545,I2973);
not I_444 (I10562,I2383);
nor I_445 (I10579,I2703,I1311);
nand I_446 (I10596,I10579,I1639);
nor I_447 (I10613,I10562,I2703);
nand I_448 (I10630,I10613,I1599);
DFFARX1 I_449 (I10647,I10630,I2966,I10545,);
not I_450 (I10516,I10647);
not I_451 (I10678,I2703);
not I_452 (I10695,I10678);
not I_453 (I10712,I1583);
nor I_454 (I10729,I10712,I2319);
and I_455 (I10746,I10729,I1519);
or I_456 (I10763,I10746,I1239);
DFFARX1 I_457 (I10780,I10763,I2966,I10545,);
DFFARX1 I_458 (I10513,I10780,I2966,I10545,);
DFFARX1 I_459 (I10811,I10780,I2966,I10545,);
DFFARX1 I_460 (I10507,I10780,I2966,I10545,);
nand I_461 (I10842,I10562,I1583);
nand I_462 (I10859,I10842,I10596);
and I_463 (I10876,I10678,I10859);
DFFARX1 I_464 (I10537,I10876,I2966,I10545,);
and I_465 (I10510,I10842,I10811);
DFFARX1 I_466 (I10921,I2095,I2966,I10545,);
nor I_467 (I10534,I10921,I10842);
nor I_468 (I10952,I10921,I10596);
nand I_469 (I10531,I10630,I10952);
not I_470 (I10528,I10921);
DFFARX1 I_471 (I10997,I1695,I2966,I10545,);
not I_472 (I11014,I10997);
nor I_473 (I11031,I11014,I10695);
and I_474 (I11048,I10921,I11031);
or I_475 (I11065,I10842,I11048);
DFFARX1 I_476 (I10522,I11065,I2966,I10545,);
not I_477 (I11096,I11014);
nor I_478 (I11113,I10921,I11096);
nand I_479 (I10525,I11014,I11113);
nand I_480 (I10519,I10678,I11096);
not I_481 (I11191,I2973);
not I_482 (I11208,I2639);
nor I_483 (I11225,I2743,I2023);
nand I_484 (I11242,I11225,I2311);
nor I_485 (I11259,I11208,I2743);
nand I_486 (I11276,I11259,I1903);
DFFARX1 I_487 (I11293,I11276,I2966,I11191,);
not I_488 (I11162,I11293);
not I_489 (I11324,I2743);
not I_490 (I11341,I11324);
not I_491 (I11358,I2879);
nor I_492 (I11375,I11358,I1527);
and I_493 (I11392,I11375,I1895);
or I_494 (I11409,I11392,I2631);
DFFARX1 I_495 (I11426,I11409,I2966,I11191,);
DFFARX1 I_496 (I11159,I11426,I2966,I11191,);
DFFARX1 I_497 (I11457,I11426,I2966,I11191,);
DFFARX1 I_498 (I11153,I11426,I2966,I11191,);
nand I_499 (I11488,I11208,I2879);
nand I_500 (I11505,I11488,I11242);
and I_501 (I11522,I11324,I11505);
DFFARX1 I_502 (I11183,I11522,I2966,I11191,);
and I_503 (I11156,I11488,I11457);
DFFARX1 I_504 (I11567,I1767,I2966,I11191,);
nor I_505 (I11180,I11567,I11488);
nor I_506 (I11598,I11567,I11242);
nand I_507 (I11177,I11276,I11598);
not I_508 (I11174,I11567);
DFFARX1 I_509 (I11643,I1615,I2966,I11191,);
not I_510 (I11660,I11643);
nor I_511 (I11677,I11660,I11341);
and I_512 (I11694,I11567,I11677);
or I_513 (I11711,I11488,I11694);
DFFARX1 I_514 (I11168,I11711,I2966,I11191,);
not I_515 (I11742,I11660);
nor I_516 (I11759,I11567,I11742);
nand I_517 (I11171,I11660,I11759);
nand I_518 (I11165,I11324,I11742);
not I_519 (I11837,I2973);
or I_520 (I11854,I2791,I1967);
or I_521 (I11871,I2399,I2791);
nor I_522 (I11888,I1463,I2135);
DFFARX1 I_523 (I11905,I11888,I2966,I11837,);
DFFARX1 I_524 (I11799,I11888,I2966,I11837,);
not I_525 (I11936,I1463);
and I_526 (I11953,I11936,I2495);
nor I_527 (I11970,I11953,I1967);
nor I_528 (I11987,I1631,I1327);
DFFARX1 I_529 (I12004,I11987,I2966,I11837,);
not I_530 (I12021,I12004);
DFFARX1 I_531 (I11808,I12004,I2966,I11837,);
nor I_532 (I12052,I1631,I2399);
and I_533 (I11802,I12052,I11905);
DFFARX1 I_534 (I12083,I1295,I2966,I11837,);
and I_535 (I12100,I12083,I1391);
nand I_536 (I12117,I12100,I11871);
and I_537 (I12134,I12004,I12117);
DFFARX1 I_538 (I11829,I12134,I2966,I11837,);
nor I_539 (I11826,I12100,I11970);
not I_540 (I12179,I12100);
nor I_541 (I12196,I11854,I12179);
nor I_542 (I12213,I12100,I12052);
nand I_543 (I11823,I11871,I12213);
nor I_544 (I12244,I12100,I12021);
not I_545 (I11820,I12100);
nand I_546 (I11811,I12100,I12021);
DFFARX1 I_547 (I12289,I2671,I2966,I11837,);
and I_548 (I12306,I12289,I12196);
or I_549 (I12323,I11854,I12306);
DFFARX1 I_550 (I11814,I12323,I2966,I11837,);
nand I_551 (I11817,I12289,I12244);
nand I_552 (I12368,I12289,I11970);
and I_553 (I12385,I11888,I12368);
DFFARX1 I_554 (I11805,I12385,I2966,I11837,);
not I_555 (I12449,I2973);
nand I_556 (I12466,I2823,I1863);
and I_557 (I12483,I12466,I2559);
DFFARX1 I_558 (I12500,I12483,I2966,I12449,);
not I_559 (I12517,I12500);
DFFARX1 I_560 (I12417,I12500,I2966,I12449,);
nor I_561 (I12548,I1791,I1863);
DFFARX1 I_562 (I12565,I1319,I2966,I12449,);
DFFARX1 I_563 (I12582,I12565,I2966,I12449,);
not I_564 (I12420,I12582);
DFFARX1 I_565 (I12613,I12565,I2966,I12449,);
and I_566 (I12414,I12500,I12613);
nand I_567 (I12644,I2847,I1959);
and I_568 (I12661,I12644,I2535);
DFFARX1 I_569 (I12678,I12661,I2966,I12449,);
nor I_570 (I12695,I12678,I12517);
not I_571 (I12712,I12678);
nand I_572 (I12423,I12500,I12712);
DFFARX1 I_573 (I12743,I2215,I2966,I12449,);
and I_574 (I12760,I12743,I2591);
nor I_575 (I12777,I12760,I12678);
nor I_576 (I12794,I12760,I12712);
nand I_577 (I12429,I12548,I12794);
not I_578 (I12432,I12760);
DFFARX1 I_579 (I12411,I12760,I2966,I12449,);
DFFARX1 I_580 (I12853,I1975,I2966,I12449,);
nand I_581 (I12870,I12853,I12565);
and I_582 (I12887,I12548,I12870);
DFFARX1 I_583 (I12441,I12887,I2966,I12449,);
nor I_584 (I12438,I12853,I12760);
and I_585 (I12932,I12853,I12695);
or I_586 (I12949,I12548,I12932);
DFFARX1 I_587 (I12426,I12949,I2966,I12449,);
nand I_588 (I12435,I12853,I12777);
not I_589 (I13027,I2973);
nand I_590 (I13044,I1551,I1495);
and I_591 (I13061,I13044,I2447);
DFFARX1 I_592 (I13078,I13061,I2966,I13027,);
nor I_593 (I13095,I1279,I1495);
DFFARX1 I_594 (I13112,I2151,I2966,I13027,);
nand I_595 (I13129,I13112,I13095);
DFFARX1 I_596 (I12998,I13112,I2966,I13027,);
nand I_597 (I13160,I1823,I1215);
and I_598 (I13177,I13160,I2103);
DFFARX1 I_599 (I13194,I13177,I2966,I13027,);
not I_600 (I13211,I13194);
nor I_601 (I13228,I13078,I13211);
and I_602 (I13245,I13095,I13228);
and I_603 (I13262,I13194,I13129);
DFFARX1 I_604 (I12995,I13262,I2966,I13027,);
DFFARX1 I_605 (I12989,I13194,I2966,I13027,);
DFFARX1 I_606 (I13307,I2159,I2966,I13027,);
and I_607 (I13324,I13307,I1983);
nand I_608 (I13341,I13324,I13194);
nor I_609 (I13016,I13324,I13095);
not I_610 (I13372,I13324);
nor I_611 (I13389,I13078,I13372);
nand I_612 (I13007,I13112,I13389);
nand I_613 (I13001,I13194,I13372);
or I_614 (I13434,I13324,I13245);
DFFARX1 I_615 (I13004,I13434,I2966,I13027,);
DFFARX1 I_616 (I13465,I1335,I2966,I13027,);
and I_617 (I13482,I13465,I13341);
DFFARX1 I_618 (I13019,I13482,I2966,I13027,);
nor I_619 (I13513,I13465,I13078);
nand I_620 (I13013,I13324,I13513);
not I_621 (I13010,I13465);
DFFARX1 I_622 (I13558,I13465,I2966,I13027,);
and I_623 (I12992,I13465,I13558);
not I_624 (I13622,I2973);
not I_625 (I13639,I2391);
nor I_626 (I13656,I1815,I2007);
nand I_627 (I13673,I13656,I1287);
nor I_628 (I13690,I13639,I1815);
nand I_629 (I13707,I13690,I2839);
not I_630 (I13724,I1815);
not I_631 (I13741,I13724);
not I_632 (I13758,I2567);
nor I_633 (I13775,I13758,I1487);
and I_634 (I13792,I13775,I1399);
or I_635 (I13809,I13792,I1671);
DFFARX1 I_636 (I13826,I13809,I2966,I13622,);
nand I_637 (I13843,I13639,I2567);
or I_638 (I13611,I13843,I13826);
not I_639 (I13874,I13843);
nor I_640 (I13891,I13826,I13874);
and I_641 (I13908,I13724,I13891);
nand I_642 (I13584,I13843,I13741);
DFFARX1 I_643 (I13939,I1247,I2966,I13622,);
or I_644 (I13605,I13939,I13826);
nor I_645 (I13970,I13939,I13707);
nor I_646 (I13987,I13939,I13741);
nand I_647 (I13590,I13673,I13987);
or I_648 (I14018,I13939,I13908);
DFFARX1 I_649 (I13587,I14018,I2966,I13622,);
not I_650 (I13593,I13939);
DFFARX1 I_651 (I14063,I2871,I2966,I13622,);
not I_652 (I14080,I14063);
nor I_653 (I14097,I14080,I13673);
DFFARX1 I_654 (I13599,I14097,I2966,I13622,);
nor I_655 (I13614,I13939,I14080);
nor I_656 (I13602,I14080,I13843);
not I_657 (I14156,I14080);
and I_658 (I14173,I13707,I14156);
nor I_659 (I13608,I13843,I14173);
nand I_660 (I13596,I14080,I13970);
not I_661 (I14251,I2973);
nand I_662 (I14268,I2519,I2031);
and I_663 (I14285,I14268,I1383);
DFFARX1 I_664 (I14302,I14285,I2966,I14251,);
not I_665 (I14240,I14302);
DFFARX1 I_666 (I14333,I14302,I2966,I14251,);
not I_667 (I14228,I14333);
nor I_668 (I14364,I1511,I2031);
not I_669 (I14381,I14364);
nor I_670 (I14398,I14302,I14381);
DFFARX1 I_671 (I14415,I2647,I2966,I14251,);
not I_672 (I14432,I14415);
nand I_673 (I14231,I14415,I14381);
DFFARX1 I_674 (I14463,I14415,I2966,I14251,);
and I_675 (I14216,I14302,I14463);
nand I_676 (I14494,I2087,I2183);
and I_677 (I14511,I14494,I1839);
DFFARX1 I_678 (I14528,I14511,I2966,I14251,);
nor I_679 (I14545,I14528,I14432);
and I_680 (I14562,I14364,I14545);
nor I_681 (I14579,I14528,I14302);
DFFARX1 I_682 (I14222,I14528,I2966,I14251,);
DFFARX1 I_683 (I14610,I1231,I2966,I14251,);
and I_684 (I14627,I14610,I1647);
or I_685 (I14644,I14627,I14562);
DFFARX1 I_686 (I14234,I14644,I2966,I14251,);
nand I_687 (I14243,I14627,I14579);
DFFARX1 I_688 (I14213,I14627,I2966,I14251,);
DFFARX1 I_689 (I14703,I1223,I2966,I14251,);
nand I_690 (I14237,I14703,I14398);
DFFARX1 I_691 (I14225,I14703,I2966,I14251,);
nand I_692 (I14748,I14703,I14364);
and I_693 (I14765,I14415,I14748);
DFFARX1 I_694 (I14219,I14765,I2966,I14251,);
not I_695 (I14829,I2973);
nand I_696 (I14846,I2279,I2615);
and I_697 (I14863,I14846,I2551);
DFFARX1 I_698 (I14880,I14863,I2966,I14829,);
not I_699 (I14818,I14880);
DFFARX1 I_700 (I14911,I14880,I2966,I14829,);
not I_701 (I14806,I14911);
nor I_702 (I14942,I2327,I2615);
not I_703 (I14959,I14942);
nor I_704 (I14976,I14880,I14959);
DFFARX1 I_705 (I14993,I2367,I2966,I14829,);
not I_706 (I15010,I14993);
nand I_707 (I14809,I14993,I14959);
DFFARX1 I_708 (I15041,I14993,I2966,I14829,);
and I_709 (I14794,I14880,I15041);
nand I_710 (I15072,I2919,I2935);
and I_711 (I15089,I15072,I2223);
DFFARX1 I_712 (I15106,I15089,I2966,I14829,);
nor I_713 (I15123,I15106,I15010);
and I_714 (I15140,I14942,I15123);
nor I_715 (I15157,I15106,I14880);
DFFARX1 I_716 (I14800,I15106,I2966,I14829,);
DFFARX1 I_717 (I15188,I1567,I2966,I14829,);
and I_718 (I15205,I15188,I2415);
or I_719 (I15222,I15205,I15140);
DFFARX1 I_720 (I14812,I15222,I2966,I14829,);
nand I_721 (I14821,I15205,I15157);
DFFARX1 I_722 (I14791,I15205,I2966,I14829,);
DFFARX1 I_723 (I15281,I2735,I2966,I14829,);
nand I_724 (I14815,I15281,I14976);
DFFARX1 I_725 (I14803,I15281,I2966,I14829,);
nand I_726 (I15326,I15281,I14942);
and I_727 (I15343,I14993,I15326);
DFFARX1 I_728 (I14797,I15343,I2966,I14829,);
not I_729 (I15407,I2973);
nand I_730 (I15424,I13584,I13587);
and I_731 (I15441,I15424,I13593);
DFFARX1 I_732 (I15458,I15441,I2966,I15407,);
not I_733 (I15475,I15458);
nor I_734 (I15492,I13605,I13587);
or I_735 (I15390,I15492,I15458);
not I_736 (I15378,I15492);
DFFARX1 I_737 (I15537,I13614,I2966,I15407,);
nor I_738 (I15554,I15537,I15492);
nand I_739 (I15571,I13602,I13599);
and I_740 (I15588,I15571,I13611);
DFFARX1 I_741 (I15605,I15588,I2966,I15407,);
nor I_742 (I15387,I15605,I15458);
not I_743 (I15636,I15605);
nor I_744 (I15653,I15537,I15636);
DFFARX1 I_745 (I15670,I13608,I2966,I15407,);
and I_746 (I15687,I15670,I13596);
or I_747 (I15396,I15687,I15492);
nand I_748 (I15375,I15687,I15653);
DFFARX1 I_749 (I15732,I13590,I2966,I15407,);
and I_750 (I15749,I15732,I15475);
nor I_751 (I15393,I15687,I15749);
nor I_752 (I15780,I15732,I15537);
DFFARX1 I_753 (I15384,I15780,I2966,I15407,);
nor I_754 (I15399,I15732,I15458);
not I_755 (I15825,I15732);
nor I_756 (I15842,I15605,I15825);
and I_757 (I15859,I15492,I15842);
or I_758 (I15876,I15687,I15859);
DFFARX1 I_759 (I15372,I15876,I2966,I15407,);
nand I_760 (I15381,I15732,I15554);
nand I_761 (I15369,I15732,I15636);
not I_762 (I15968,I2973);
nand I_763 (I15985,I9891,I9882);
and I_764 (I16002,I15985,I9885);
DFFARX1 I_765 (I16019,I16002,I2966,I15968,);
not I_766 (I16036,I16019);
nor I_767 (I16053,I9861,I9882);
or I_768 (I15951,I16053,I16019);
not I_769 (I15939,I16053);
DFFARX1 I_770 (I16098,I9876,I2966,I15968,);
nor I_771 (I16115,I16098,I16053);
nand I_772 (I16132,I9864,I9879);
and I_773 (I16149,I16132,I9873);
DFFARX1 I_774 (I16166,I16149,I2966,I15968,);
nor I_775 (I15948,I16166,I16019);
not I_776 (I16197,I16166);
nor I_777 (I16214,I16098,I16197);
DFFARX1 I_778 (I16231,I9888,I2966,I15968,);
and I_779 (I16248,I16231,I9867);
or I_780 (I15957,I16248,I16053);
nand I_781 (I15936,I16248,I16214);
DFFARX1 I_782 (I16293,I9870,I2966,I15968,);
and I_783 (I16310,I16293,I16036);
nor I_784 (I15954,I16248,I16310);
nor I_785 (I16341,I16293,I16098);
DFFARX1 I_786 (I15945,I16341,I2966,I15968,);
nor I_787 (I15960,I16293,I16019);
not I_788 (I16386,I16293);
nor I_789 (I16403,I16166,I16386);
and I_790 (I16420,I16053,I16403);
or I_791 (I16437,I16248,I16420);
DFFARX1 I_792 (I15933,I16437,I2966,I15968,);
nand I_793 (I15942,I16293,I16115);
nand I_794 (I15930,I16293,I16197);
not I_795 (I16529,I2973);
nand I_796 (I16546,I5326,I5329);
and I_797 (I16563,I16546,I5311);
DFFARX1 I_798 (I16580,I16563,I2966,I16529,);
not I_799 (I16597,I16580);
nor I_800 (I16614,I5308,I5329);
or I_801 (I16512,I16614,I16580);
not I_802 (I16500,I16614);
DFFARX1 I_803 (I16659,I5332,I2966,I16529,);
nor I_804 (I16676,I16659,I16614);
nand I_805 (I16693,I5317,I5323);
and I_806 (I16710,I16693,I5335);
DFFARX1 I_807 (I16727,I16710,I2966,I16529,);
nor I_808 (I16509,I16727,I16580);
not I_809 (I16758,I16727);
nor I_810 (I16775,I16659,I16758);
DFFARX1 I_811 (I16792,I5314,I2966,I16529,);
and I_812 (I16809,I16792,I5305);
or I_813 (I16518,I16809,I16614);
nand I_814 (I16497,I16809,I16775);
DFFARX1 I_815 (I16854,I5320,I2966,I16529,);
and I_816 (I16871,I16854,I16597);
nor I_817 (I16515,I16809,I16871);
nor I_818 (I16902,I16854,I16659);
DFFARX1 I_819 (I16506,I16902,I2966,I16529,);
nor I_820 (I16521,I16854,I16580);
not I_821 (I16947,I16854);
nor I_822 (I16964,I16727,I16947);
and I_823 (I16981,I16614,I16964);
or I_824 (I16998,I16809,I16981);
DFFARX1 I_825 (I16494,I16998,I2966,I16529,);
nand I_826 (I16503,I16854,I16676);
nand I_827 (I16491,I16854,I16758);
not I_828 (I17090,I2973);
not I_829 (I17107,I5969);
nor I_830 (I17124,I5957,I5963);
nand I_831 (I17141,I17124,I5972);
DFFARX1 I_832 (I17064,I17141,I2966,I17090,);
nor I_833 (I17172,I17107,I5957);
nand I_834 (I17189,I17172,I5960);
not I_835 (I17079,I17189);
DFFARX1 I_836 (I17061,I17189,I2966,I17090,);
not I_837 (I17234,I5957);
not I_838 (I17251,I17234);
not I_839 (I17268,I5981);
nor I_840 (I17285,I17268,I5954);
and I_841 (I17302,I17285,I5975);
or I_842 (I17319,I17302,I5966);
DFFARX1 I_843 (I17336,I17319,I2966,I17090,);
nor I_844 (I17353,I17336,I17189);
nor I_845 (I17370,I17336,I17251);
nand I_846 (I17076,I17141,I17370);
nand I_847 (I17401,I17107,I5981);
nand I_848 (I17418,I17401,I17336);
and I_849 (I17435,I17401,I17418);
DFFARX1 I_850 (I17058,I17435,I2966,I17090,);
DFFARX1 I_851 (I17466,I17401,I2966,I17090,);
and I_852 (I17055,I17234,I17466);
DFFARX1 I_853 (I17497,I5951,I2966,I17090,);
not I_854 (I17514,I17497);
nor I_855 (I17531,I17189,I17514);
and I_856 (I17548,I17497,I17531);
nand I_857 (I17070,I17497,I17251);
DFFARX1 I_858 (I17579,I17497,I2966,I17090,);
not I_859 (I17067,I17579);
DFFARX1 I_860 (I17610,I5978,I2966,I17090,);
not I_861 (I17627,I17610);
or I_862 (I17644,I17627,I17548);
DFFARX1 I_863 (I17073,I17644,I2966,I17090,);
nand I_864 (I17082,I17627,I17353);
DFFARX1 I_865 (I17052,I17627,I2966,I17090,);
not I_866 (I17736,I2973);
not I_867 (I17753,I8553);
nor I_868 (I17770,I8550,I8538);
nand I_869 (I17787,I17770,I8541);
DFFARX1 I_870 (I17710,I17787,I2966,I17736,);
nor I_871 (I17818,I17753,I8550);
nand I_872 (I17835,I17818,I8547);
not I_873 (I17725,I17835);
DFFARX1 I_874 (I17707,I17835,I2966,I17736,);
not I_875 (I17880,I8550);
not I_876 (I17897,I17880);
not I_877 (I17914,I8559);
nor I_878 (I17931,I17914,I8535);
and I_879 (I17948,I17931,I8556);
or I_880 (I17965,I17948,I8544);
DFFARX1 I_881 (I17982,I17965,I2966,I17736,);
nor I_882 (I17999,I17982,I17835);
nor I_883 (I18016,I17982,I17897);
nand I_884 (I17722,I17787,I18016);
nand I_885 (I18047,I17753,I8559);
nand I_886 (I18064,I18047,I17982);
and I_887 (I18081,I18047,I18064);
DFFARX1 I_888 (I17704,I18081,I2966,I17736,);
DFFARX1 I_889 (I18112,I18047,I2966,I17736,);
and I_890 (I17701,I17880,I18112);
DFFARX1 I_891 (I18143,I8565,I2966,I17736,);
not I_892 (I18160,I18143);
nor I_893 (I18177,I17835,I18160);
and I_894 (I18194,I18143,I18177);
nand I_895 (I17716,I18143,I17897);
DFFARX1 I_896 (I18225,I18143,I2966,I17736,);
not I_897 (I17713,I18225);
DFFARX1 I_898 (I18256,I8562,I2966,I17736,);
not I_899 (I18273,I18256);
or I_900 (I18290,I18273,I18194);
DFFARX1 I_901 (I17719,I18290,I2966,I17736,);
nand I_902 (I17728,I18273,I17999);
DFFARX1 I_903 (I17698,I18273,I2966,I17736,);
not I_904 (I18382,I2973);
not I_905 (I18399,I9216);
nor I_906 (I18416,I9213,I9201);
nand I_907 (I18433,I18416,I9204);
DFFARX1 I_908 (I18356,I18433,I2966,I18382,);
nor I_909 (I18464,I18399,I9213);
nand I_910 (I18481,I18464,I9210);
not I_911 (I18371,I18481);
DFFARX1 I_912 (I18353,I18481,I2966,I18382,);
not I_913 (I18526,I9213);
not I_914 (I18543,I18526);
not I_915 (I18560,I9222);
nor I_916 (I18577,I18560,I9198);
and I_917 (I18594,I18577,I9219);
or I_918 (I18611,I18594,I9207);
DFFARX1 I_919 (I18628,I18611,I2966,I18382,);
nor I_920 (I18645,I18628,I18481);
nor I_921 (I18662,I18628,I18543);
nand I_922 (I18368,I18433,I18662);
nand I_923 (I18693,I18399,I9222);
nand I_924 (I18710,I18693,I18628);
and I_925 (I18727,I18693,I18710);
DFFARX1 I_926 (I18350,I18727,I2966,I18382,);
DFFARX1 I_927 (I18758,I18693,I2966,I18382,);
and I_928 (I18347,I18526,I18758);
DFFARX1 I_929 (I18789,I9228,I2966,I18382,);
not I_930 (I18806,I18789);
nor I_931 (I18823,I18481,I18806);
and I_932 (I18840,I18789,I18823);
nand I_933 (I18362,I18789,I18543);
DFFARX1 I_934 (I18871,I18789,I2966,I18382,);
not I_935 (I18359,I18871);
DFFARX1 I_936 (I18902,I9225,I2966,I18382,);
not I_937 (I18919,I18902);
or I_938 (I18936,I18919,I18840);
DFFARX1 I_939 (I18365,I18936,I2966,I18382,);
nand I_940 (I18374,I18919,I18645);
DFFARX1 I_941 (I18344,I18919,I2966,I18382,);
not I_942 (I19028,I2973);
not I_943 (I19045,I17713);
nor I_944 (I19062,I17701,I17725);
nand I_945 (I19079,I19062,I17710);
DFFARX1 I_946 (I18999,I19079,I2966,I19028,);
nor I_947 (I19110,I19045,I17701);
nand I_948 (I19127,I19110,I17728);
nand I_949 (I19144,I19127,I19079);
not I_950 (I19161,I17701);
not I_951 (I19178,I17698);
nor I_952 (I19195,I19178,I17707);
and I_953 (I19212,I19195,I17722);
or I_954 (I19229,I19212,I17704);
DFFARX1 I_955 (I19246,I19229,I2966,I19028,);
nor I_956 (I19263,I19246,I19127);
nand I_957 (I19014,I19161,I19263);
not I_958 (I19011,I19246);
and I_959 (I19308,I19246,I19144);
DFFARX1 I_960 (I18996,I19308,I2966,I19028,);
DFFARX1 I_961 (I19339,I19246,I2966,I19028,);
and I_962 (I18993,I19161,I19339);
nand I_963 (I19370,I19045,I17698);
not I_964 (I19387,I19370);
nor I_965 (I19404,I19246,I19387);
DFFARX1 I_966 (I19421,I17719,I2966,I19028,);
nand I_967 (I19438,I19421,I19370);
and I_968 (I19455,I19161,I19438);
DFFARX1 I_969 (I19020,I19455,I2966,I19028,);
not I_970 (I19486,I19421);
nand I_971 (I19008,I19421,I19404);
nand I_972 (I19002,I19421,I19387);
DFFARX1 I_973 (I19531,I17716,I2966,I19028,);
not I_974 (I19548,I19531);
nor I_975 (I19017,I19421,I19548);
nor I_976 (I19579,I19548,I19486);
and I_977 (I19596,I19127,I19579);
or I_978 (I19613,I19370,I19596);
DFFARX1 I_979 (I19005,I19613,I2966,I19028,);
DFFARX1 I_980 (I18990,I19548,I2966,I19028,);
not I_981 (I19691,I2973);
or I_982 (I19708,I7872,I7887);
or I_983 (I19725,I7875,I7872);
DFFARX1 I_984 (I19665,I19725,I2966,I19691,);
nor I_985 (I19756,I7878,I7893);
not I_986 (I19773,I19756);
not I_987 (I19790,I7878);
and I_988 (I19807,I19790,I7881);
nor I_989 (I19824,I19807,I7887);
nor I_990 (I19841,I7884,I7902);
DFFARX1 I_991 (I19858,I19841,I2966,I19691,);
nand I_992 (I19875,I19858,I19708);
and I_993 (I19892,I19824,I19875);
DFFARX1 I_994 (I19659,I19892,I2966,I19691,);
nor I_995 (I19923,I7884,I7875);
DFFARX1 I_996 (I19940,I19923,I2966,I19691,);
and I_997 (I19656,I19756,I19940);
DFFARX1 I_998 (I19971,I7899,I2966,I19691,);
and I_999 (I19988,I19971,I7890);
DFFARX1 I_1000 (I20005,I19988,I2966,I19691,);
not I_1001 (I19668,I20005);
DFFARX1 I_1002 (I19653,I19988,I2966,I19691,);
DFFARX1 I_1003 (I20050,I7896,I2966,I19691,);
not I_1004 (I20067,I20050);
nor I_1005 (I20084,I19725,I20067);
and I_1006 (I20101,I19988,I20084);
or I_1007 (I20118,I19708,I20101);
DFFARX1 I_1008 (I19674,I20118,I2966,I19691,);
nor I_1009 (I20149,I20050,I19858);
nand I_1010 (I19683,I19824,I20149);
nor I_1011 (I20180,I20050,I19773);
nand I_1012 (I19677,I19923,I20180);
not I_1013 (I19680,I20050);
nand I_1014 (I19671,I20050,I19773);
DFFARX1 I_1015 (I19662,I20050,I2966,I19691,);
not I_1016 (I20286,I2973);
not I_1017 (I20303,I2994);
nor I_1018 (I20320,I3000,I3003);
nand I_1019 (I20337,I20320,I2979);
nor I_1020 (I20354,I20303,I3000);
nand I_1021 (I20371,I20354,I2988);
not I_1022 (I20388,I20371);
not I_1023 (I20405,I3000);
nor I_1024 (I20275,I20371,I20405);
not I_1025 (I20436,I20405);
nand I_1026 (I20260,I20371,I20436);
not I_1027 (I20467,I2982);
nor I_1028 (I20484,I20467,I3006);
and I_1029 (I20501,I20484,I2976);
or I_1030 (I20518,I20501,I2985);
DFFARX1 I_1031 (I20535,I20518,I2966,I20286,);
nor I_1032 (I20552,I20535,I20388);
DFFARX1 I_1033 (I20569,I20535,I2966,I20286,);
not I_1034 (I20257,I20569);
nand I_1035 (I20600,I20303,I2982);
and I_1036 (I20617,I20600,I20552);
DFFARX1 I_1037 (I20254,I20600,I2966,I20286,);
DFFARX1 I_1038 (I20648,I2991,I2966,I20286,);
nor I_1039 (I20665,I20648,I20371);
nand I_1040 (I20272,I20535,I20665);
nor I_1041 (I20696,I20648,I20436);
not I_1042 (I20269,I20648);
nand I_1043 (I20727,I20648,I20337);
and I_1044 (I20744,I20405,I20727);
DFFARX1 I_1045 (I20248,I20744,I2966,I20286,);
DFFARX1 I_1046 (I20251,I20648,I2966,I20286,);
DFFARX1 I_1047 (I20789,I2997,I2966,I20286,);
not I_1048 (I20806,I20789);
nand I_1049 (I20823,I20806,I20371);
and I_1050 (I20840,I20600,I20823);
DFFARX1 I_1051 (I20278,I20840,I2966,I20286,);
or I_1052 (I20871,I20806,I20617);
DFFARX1 I_1053 (I20263,I20871,I2966,I20286,);
nand I_1054 (I20266,I20806,I20696);
not I_1055 (I20949,I2973);
not I_1056 (I20966,I19671);
nor I_1057 (I20983,I19665,I19656);
nand I_1058 (I21000,I20983,I19668);
nor I_1059 (I21017,I20966,I19665);
nand I_1060 (I21034,I21017,I19683);
not I_1061 (I21051,I21034);
not I_1062 (I21068,I19665);
nor I_1063 (I20938,I21034,I21068);
not I_1064 (I21099,I21068);
nand I_1065 (I20923,I21034,I21099);
not I_1066 (I21130,I19659);
nor I_1067 (I21147,I21130,I19653);
and I_1068 (I21164,I21147,I19680);
or I_1069 (I21181,I21164,I19677);
DFFARX1 I_1070 (I21198,I21181,I2966,I20949,);
nor I_1071 (I21215,I21198,I21051);
DFFARX1 I_1072 (I21232,I21198,I2966,I20949,);
not I_1073 (I20920,I21232);
nand I_1074 (I21263,I20966,I19659);
and I_1075 (I21280,I21263,I21215);
DFFARX1 I_1076 (I20917,I21263,I2966,I20949,);
DFFARX1 I_1077 (I21311,I19674,I2966,I20949,);
nor I_1078 (I21328,I21311,I21034);
nand I_1079 (I20935,I21198,I21328);
nor I_1080 (I21359,I21311,I21099);
not I_1081 (I20932,I21311);
nand I_1082 (I21390,I21311,I21000);
and I_1083 (I21407,I21068,I21390);
DFFARX1 I_1084 (I20911,I21407,I2966,I20949,);
DFFARX1 I_1085 (I20914,I21311,I2966,I20949,);
DFFARX1 I_1086 (I21452,I19662,I2966,I20949,);
not I_1087 (I21469,I21452);
nand I_1088 (I21486,I21469,I21034);
and I_1089 (I21503,I21263,I21486);
DFFARX1 I_1090 (I20941,I21503,I2966,I20949,);
or I_1091 (I21534,I21469,I21280);
DFFARX1 I_1092 (I20926,I21534,I2966,I20949,);
nand I_1093 (I20929,I21469,I21359);
not I_1094 (I21612,I2973);
not I_1095 (I21629,I11805);
nor I_1096 (I21646,I11808,I11814);
nand I_1097 (I21663,I21646,I11820);
nor I_1098 (I21680,I21629,I11808);
nand I_1099 (I21697,I21680,I11799);
not I_1100 (I21714,I21697);
not I_1101 (I21731,I11808);
nor I_1102 (I21601,I21697,I21731);
not I_1103 (I21762,I21731);
nand I_1104 (I21586,I21697,I21762);
not I_1105 (I21793,I11811);
nor I_1106 (I21810,I21793,I11826);
and I_1107 (I21827,I21810,I11829);
or I_1108 (I21844,I21827,I11802);
DFFARX1 I_1109 (I21861,I21844,I2966,I21612,);
nor I_1110 (I21878,I21861,I21714);
DFFARX1 I_1111 (I21895,I21861,I2966,I21612,);
not I_1112 (I21583,I21895);
nand I_1113 (I21926,I21629,I11811);
and I_1114 (I21943,I21926,I21878);
DFFARX1 I_1115 (I21580,I21926,I2966,I21612,);
DFFARX1 I_1116 (I21974,I11823,I2966,I21612,);
nor I_1117 (I21991,I21974,I21697);
nand I_1118 (I21598,I21861,I21991);
nor I_1119 (I22022,I21974,I21762);
not I_1120 (I21595,I21974);
nand I_1121 (I22053,I21974,I21663);
and I_1122 (I22070,I21731,I22053);
DFFARX1 I_1123 (I21574,I22070,I2966,I21612,);
DFFARX1 I_1124 (I21577,I21974,I2966,I21612,);
DFFARX1 I_1125 (I22115,I11817,I2966,I21612,);
not I_1126 (I22132,I22115);
nand I_1127 (I22149,I22132,I21697);
and I_1128 (I22166,I21926,I22149);
DFFARX1 I_1129 (I21604,I22166,I2966,I21612,);
or I_1130 (I22197,I22132,I21943);
DFFARX1 I_1131 (I21589,I22197,I2966,I21612,);
nand I_1132 (I21592,I22132,I22022);
not I_1133 (I22275,I2973);
not I_1134 (I22292,I4665);
nor I_1135 (I22309,I4662,I4686);
nand I_1136 (I22326,I22309,I4683);
nor I_1137 (I22343,I22292,I4662);
nand I_1138 (I22360,I22343,I4689);
not I_1139 (I22377,I22360);
not I_1140 (I22394,I4662);
nor I_1141 (I22264,I22360,I22394);
not I_1142 (I22425,I22394);
nand I_1143 (I22249,I22360,I22425);
not I_1144 (I22456,I4680);
nor I_1145 (I22473,I22456,I4671);
and I_1146 (I22490,I22473,I4668);
or I_1147 (I22507,I22490,I4677);
DFFARX1 I_1148 (I22524,I22507,I2966,I22275,);
nor I_1149 (I22541,I22524,I22377);
DFFARX1 I_1150 (I22558,I22524,I2966,I22275,);
not I_1151 (I22246,I22558);
nand I_1152 (I22589,I22292,I4680);
and I_1153 (I22606,I22589,I22541);
DFFARX1 I_1154 (I22243,I22589,I2966,I22275,);
DFFARX1 I_1155 (I22637,I4659,I2966,I22275,);
nor I_1156 (I22654,I22637,I22360);
nand I_1157 (I22261,I22524,I22654);
nor I_1158 (I22685,I22637,I22425);
not I_1159 (I22258,I22637);
nand I_1160 (I22716,I22637,I22326);
and I_1161 (I22733,I22394,I22716);
DFFARX1 I_1162 (I22237,I22733,I2966,I22275,);
DFFARX1 I_1163 (I22240,I22637,I2966,I22275,);
DFFARX1 I_1164 (I22778,I4674,I2966,I22275,);
not I_1165 (I22795,I22778);
nand I_1166 (I22812,I22795,I22360);
and I_1167 (I22829,I22589,I22812);
DFFARX1 I_1168 (I22267,I22829,I2966,I22275,);
or I_1169 (I22860,I22795,I22606);
DFFARX1 I_1170 (I22252,I22860,I2966,I22275,);
nand I_1171 (I22255,I22795,I22685);
not I_1172 (I22938,I2973);
not I_1173 (I22955,I3555);
nor I_1174 (I22972,I3561,I3564);
nand I_1175 (I22989,I22972,I3540);
nor I_1176 (I23006,I22955,I3561);
nand I_1177 (I23023,I23006,I3549);
not I_1178 (I23040,I23023);
not I_1179 (I23057,I3561);
nor I_1180 (I22927,I23023,I23057);
not I_1181 (I23088,I23057);
nand I_1182 (I22912,I23023,I23088);
not I_1183 (I23119,I3543);
nor I_1184 (I23136,I23119,I3567);
and I_1185 (I23153,I23136,I3537);
or I_1186 (I23170,I23153,I3546);
DFFARX1 I_1187 (I23187,I23170,I2966,I22938,);
nor I_1188 (I23204,I23187,I23040);
DFFARX1 I_1189 (I23221,I23187,I2966,I22938,);
not I_1190 (I22909,I23221);
nand I_1191 (I23252,I22955,I3543);
and I_1192 (I23269,I23252,I23204);
DFFARX1 I_1193 (I22906,I23252,I2966,I22938,);
DFFARX1 I_1194 (I23300,I3552,I2966,I22938,);
nor I_1195 (I23317,I23300,I23023);
nand I_1196 (I22924,I23187,I23317);
nor I_1197 (I23348,I23300,I23088);
not I_1198 (I22921,I23300);
nand I_1199 (I23379,I23300,I22989);
and I_1200 (I23396,I23057,I23379);
DFFARX1 I_1201 (I22900,I23396,I2966,I22938,);
DFFARX1 I_1202 (I22903,I23300,I2966,I22938,);
DFFARX1 I_1203 (I23441,I3558,I2966,I22938,);
not I_1204 (I23458,I23441);
nand I_1205 (I23475,I23458,I23023);
and I_1206 (I23492,I23252,I23475);
DFFARX1 I_1207 (I22930,I23492,I2966,I22938,);
or I_1208 (I23523,I23458,I23269);
DFFARX1 I_1209 (I22915,I23523,I2966,I22938,);
nand I_1210 (I22918,I23458,I23348);
not I_1211 (I23601,I2973);
not I_1212 (I23618,I10519);
nor I_1213 (I23635,I10516,I10534);
nand I_1214 (I23652,I23635,I10537);
nor I_1215 (I23669,I23618,I10516);
nand I_1216 (I23686,I23669,I10522);
not I_1217 (I23703,I23686);
not I_1218 (I23720,I10516);
nor I_1219 (I23590,I23686,I23720);
not I_1220 (I23751,I23720);
nand I_1221 (I23575,I23686,I23751);
not I_1222 (I23782,I10531);
nor I_1223 (I23799,I23782,I10513);
and I_1224 (I23816,I23799,I10507);
or I_1225 (I23833,I23816,I10525);
DFFARX1 I_1226 (I23850,I23833,I2966,I23601,);
nor I_1227 (I23867,I23850,I23703);
DFFARX1 I_1228 (I23884,I23850,I2966,I23601,);
not I_1229 (I23572,I23884);
nand I_1230 (I23915,I23618,I10531);
and I_1231 (I23932,I23915,I23867);
DFFARX1 I_1232 (I23569,I23915,I2966,I23601,);
DFFARX1 I_1233 (I23963,I10510,I2966,I23601,);
nor I_1234 (I23980,I23963,I23686);
nand I_1235 (I23587,I23850,I23980);
nor I_1236 (I24011,I23963,I23751);
not I_1237 (I23584,I23963);
nand I_1238 (I24042,I23963,I23652);
and I_1239 (I24059,I23720,I24042);
DFFARX1 I_1240 (I23563,I24059,I2966,I23601,);
DFFARX1 I_1241 (I23566,I23963,I2966,I23601,);
DFFARX1 I_1242 (I24104,I10528,I2966,I23601,);
not I_1243 (I24121,I24104);
nand I_1244 (I24138,I24121,I23686);
and I_1245 (I24155,I23915,I24138);
DFFARX1 I_1246 (I23593,I24155,I2966,I23601,);
or I_1247 (I24186,I24121,I23932);
DFFARX1 I_1248 (I23578,I24186,I2966,I23601,);
nand I_1249 (I23581,I24121,I24011);
not I_1250 (I24264,I2973);
not I_1251 (I24281,I20272);
nor I_1252 (I24298,I20251,I20263);
nand I_1253 (I24315,I24298,I20266);
nor I_1254 (I24332,I24281,I20251);
nand I_1255 (I24349,I24332,I20248);
DFFARX1 I_1256 (I24366,I24349,I2966,I24264,);
not I_1257 (I24235,I24366);
not I_1258 (I24397,I20251);
not I_1259 (I24414,I24397);
not I_1260 (I24431,I20269);
nor I_1261 (I24448,I24431,I20260);
and I_1262 (I24465,I24448,I20254);
or I_1263 (I24482,I24465,I20278);
DFFARX1 I_1264 (I24499,I24482,I2966,I24264,);
DFFARX1 I_1265 (I24232,I24499,I2966,I24264,);
DFFARX1 I_1266 (I24530,I24499,I2966,I24264,);
DFFARX1 I_1267 (I24226,I24499,I2966,I24264,);
nand I_1268 (I24561,I24281,I20269);
nand I_1269 (I24578,I24561,I24315);
and I_1270 (I24595,I24397,I24578);
DFFARX1 I_1271 (I24256,I24595,I2966,I24264,);
and I_1272 (I24229,I24561,I24530);
DFFARX1 I_1273 (I24640,I20275,I2966,I24264,);
nor I_1274 (I24253,I24640,I24561);
nor I_1275 (I24671,I24640,I24315);
nand I_1276 (I24250,I24349,I24671);
not I_1277 (I24247,I24640);
DFFARX1 I_1278 (I24716,I20257,I2966,I24264,);
not I_1279 (I24733,I24716);
nor I_1280 (I24750,I24733,I24414);
and I_1281 (I24767,I24640,I24750);
or I_1282 (I24784,I24561,I24767);
DFFARX1 I_1283 (I24241,I24784,I2966,I24264,);
not I_1284 (I24815,I24733);
nor I_1285 (I24832,I24640,I24815);
nand I_1286 (I24244,I24733,I24832);
nand I_1287 (I24238,I24397,I24815);
not I_1288 (I24910,I2973);
nand I_1289 (I24927,I4113,I4128);
and I_1290 (I24944,I24927,I4116);
DFFARX1 I_1291 (I24961,I24944,I2966,I24910,);
not I_1292 (I24978,I24961);
DFFARX1 I_1293 (I24878,I24961,I2966,I24910,);
nor I_1294 (I25009,I4125,I4128);
DFFARX1 I_1295 (I25026,I4110,I2966,I24910,);
DFFARX1 I_1296 (I25043,I25026,I2966,I24910,);
not I_1297 (I24881,I25043);
DFFARX1 I_1298 (I25074,I25026,I2966,I24910,);
and I_1299 (I24875,I24961,I25074);
nand I_1300 (I25105,I4101,I4098);
and I_1301 (I25122,I25105,I4104);
DFFARX1 I_1302 (I25139,I25122,I2966,I24910,);
nor I_1303 (I25156,I25139,I24978);
not I_1304 (I25173,I25139);
nand I_1305 (I24884,I24961,I25173);
DFFARX1 I_1306 (I25204,I4107,I2966,I24910,);
and I_1307 (I25221,I25204,I4119);
nor I_1308 (I25238,I25221,I25139);
nor I_1309 (I25255,I25221,I25173);
nand I_1310 (I24890,I25009,I25255);
not I_1311 (I24893,I25221);
DFFARX1 I_1312 (I24872,I25221,I2966,I24910,);
DFFARX1 I_1313 (I25314,I4122,I2966,I24910,);
nand I_1314 (I25331,I25314,I25026);
and I_1315 (I25348,I25009,I25331);
DFFARX1 I_1316 (I24902,I25348,I2966,I24910,);
nor I_1317 (I24899,I25314,I25221);
and I_1318 (I25393,I25314,I25156);
or I_1319 (I25410,I25009,I25393);
DFFARX1 I_1320 (I24887,I25410,I2966,I24910,);
nand I_1321 (I24896,I25314,I25238);
not I_1322 (I25488,I2973);
nand I_1323 (I25505,I16506,I16521);
and I_1324 (I25522,I25505,I16509);
DFFARX1 I_1325 (I25539,I25522,I2966,I25488,);
not I_1326 (I25556,I25539);
DFFARX1 I_1327 (I25456,I25539,I2966,I25488,);
nor I_1328 (I25587,I16518,I16521);
DFFARX1 I_1329 (I25604,I16503,I2966,I25488,);
DFFARX1 I_1330 (I25621,I25604,I2966,I25488,);
not I_1331 (I25459,I25621);
DFFARX1 I_1332 (I25652,I25604,I2966,I25488,);
and I_1333 (I25453,I25539,I25652);
nand I_1334 (I25683,I16494,I16491);
and I_1335 (I25700,I25683,I16497);
DFFARX1 I_1336 (I25717,I25700,I2966,I25488,);
nor I_1337 (I25734,I25717,I25556);
not I_1338 (I25751,I25717);
nand I_1339 (I25462,I25539,I25751);
DFFARX1 I_1340 (I25782,I16500,I2966,I25488,);
and I_1341 (I25799,I25782,I16512);
nor I_1342 (I25816,I25799,I25717);
nor I_1343 (I25833,I25799,I25751);
nand I_1344 (I25468,I25587,I25833);
not I_1345 (I25471,I25799);
DFFARX1 I_1346 (I25450,I25799,I2966,I25488,);
DFFARX1 I_1347 (I25892,I16515,I2966,I25488,);
nand I_1348 (I25909,I25892,I25604);
and I_1349 (I25926,I25587,I25909);
DFFARX1 I_1350 (I25480,I25926,I2966,I25488,);
nor I_1351 (I25477,I25892,I25799);
and I_1352 (I25971,I25892,I25734);
or I_1353 (I25988,I25587,I25971);
DFFARX1 I_1354 (I25465,I25988,I2966,I25488,);
nand I_1355 (I25474,I25892,I25816);
not I_1356 (I26066,I2973);
nand I_1357 (I26083,I17073,I17055);
and I_1358 (I26100,I26083,I17067);
DFFARX1 I_1359 (I26117,I26100,I2966,I26066,);
not I_1360 (I26134,I26117);
DFFARX1 I_1361 (I26034,I26117,I2966,I26066,);
nor I_1362 (I26165,I17070,I17055);
DFFARX1 I_1363 (I26182,I17079,I2966,I26066,);
DFFARX1 I_1364 (I26199,I26182,I2966,I26066,);
not I_1365 (I26037,I26199);
DFFARX1 I_1366 (I26230,I26182,I2966,I26066,);
and I_1367 (I26031,I26117,I26230);
nand I_1368 (I26261,I17058,I17082);
and I_1369 (I26278,I26261,I17061);
DFFARX1 I_1370 (I26295,I26278,I2966,I26066,);
nor I_1371 (I26312,I26295,I26134);
not I_1372 (I26329,I26295);
nand I_1373 (I26040,I26117,I26329);
DFFARX1 I_1374 (I26360,I17064,I2966,I26066,);
and I_1375 (I26377,I26360,I17076);
nor I_1376 (I26394,I26377,I26295);
nor I_1377 (I26411,I26377,I26329);
nand I_1378 (I26046,I26165,I26411);
not I_1379 (I26049,I26377);
DFFARX1 I_1380 (I26028,I26377,I2966,I26066,);
DFFARX1 I_1381 (I26470,I17052,I2966,I26066,);
nand I_1382 (I26487,I26470,I26182);
and I_1383 (I26504,I26165,I26487);
DFFARX1 I_1384 (I26058,I26504,I2966,I26066,);
nor I_1385 (I26055,I26470,I26377);
and I_1386 (I26549,I26470,I26312);
or I_1387 (I26566,I26165,I26549);
DFFARX1 I_1388 (I26043,I26566,I2966,I26066,);
nand I_1389 (I26052,I26470,I26394);
not I_1390 (I26644,I2973);
nand I_1391 (I26661,I18365,I18347);
and I_1392 (I26678,I26661,I18359);
DFFARX1 I_1393 (I26695,I26678,I2966,I26644,);
not I_1394 (I26712,I26695);
DFFARX1 I_1395 (I26612,I26695,I2966,I26644,);
nor I_1396 (I26743,I18362,I18347);
DFFARX1 I_1397 (I26760,I18371,I2966,I26644,);
DFFARX1 I_1398 (I26777,I26760,I2966,I26644,);
not I_1399 (I26615,I26777);
DFFARX1 I_1400 (I26808,I26760,I2966,I26644,);
and I_1401 (I26609,I26695,I26808);
nand I_1402 (I26839,I18350,I18374);
and I_1403 (I26856,I26839,I18353);
DFFARX1 I_1404 (I26873,I26856,I2966,I26644,);
nor I_1405 (I26890,I26873,I26712);
not I_1406 (I26907,I26873);
nand I_1407 (I26618,I26695,I26907);
DFFARX1 I_1408 (I26938,I18356,I2966,I26644,);
and I_1409 (I26955,I26938,I18368);
nor I_1410 (I26972,I26955,I26873);
nor I_1411 (I26989,I26955,I26907);
nand I_1412 (I26624,I26743,I26989);
not I_1413 (I26627,I26955);
DFFARX1 I_1414 (I26606,I26955,I2966,I26644,);
DFFARX1 I_1415 (I27048,I18344,I2966,I26644,);
nand I_1416 (I27065,I27048,I26760);
and I_1417 (I27082,I26743,I27065);
DFFARX1 I_1418 (I26636,I27082,I2966,I26644,);
nor I_1419 (I26633,I27048,I26955);
and I_1420 (I27127,I27048,I26890);
or I_1421 (I27144,I26743,I27127);
DFFARX1 I_1422 (I26621,I27144,I2966,I26644,);
nand I_1423 (I26630,I27048,I26972);
not I_1424 (I27222,I2973);
nand I_1425 (I27239,I6614,I6617);
and I_1426 (I27256,I27239,I6623);
DFFARX1 I_1427 (I27273,I27256,I2966,I27222,);
not I_1428 (I27290,I27273);
DFFARX1 I_1429 (I27190,I27273,I2966,I27222,);
nor I_1430 (I27321,I6635,I6617);
DFFARX1 I_1431 (I27338,I6626,I2966,I27222,);
DFFARX1 I_1432 (I27355,I27338,I2966,I27222,);
not I_1433 (I27193,I27355);
DFFARX1 I_1434 (I27386,I27338,I2966,I27222,);
and I_1435 (I27187,I27273,I27386);
nand I_1436 (I27417,I6632,I6629);
and I_1437 (I27434,I27417,I6641);
DFFARX1 I_1438 (I27451,I27434,I2966,I27222,);
nor I_1439 (I27468,I27451,I27290);
not I_1440 (I27485,I27451);
nand I_1441 (I27196,I27273,I27485);
DFFARX1 I_1442 (I27516,I6638,I2966,I27222,);
and I_1443 (I27533,I27516,I6644);
nor I_1444 (I27550,I27533,I27451);
nor I_1445 (I27567,I27533,I27485);
nand I_1446 (I27202,I27321,I27567);
not I_1447 (I27205,I27533);
DFFARX1 I_1448 (I27184,I27533,I2966,I27222,);
DFFARX1 I_1449 (I27626,I6620,I2966,I27222,);
nand I_1450 (I27643,I27626,I27338);
and I_1451 (I27660,I27321,I27643);
DFFARX1 I_1452 (I27214,I27660,I2966,I27222,);
nor I_1453 (I27211,I27626,I27533);
and I_1454 (I27705,I27626,I27468);
or I_1455 (I27722,I27321,I27705);
DFFARX1 I_1456 (I27199,I27722,I2966,I27222,);
nand I_1457 (I27208,I27626,I27550);
not I_1458 (I27800,I2973);
or I_1459 (I27817,I26624,I26615);
or I_1460 (I27834,I26612,I26624);
nor I_1461 (I27851,I26618,I26609);
not I_1462 (I27868,I27851);
DFFARX1 I_1463 (I27768,I27851,I2966,I27800,);
nand I_1464 (I27899,I27851,I27817);
not I_1465 (I27916,I26618);
and I_1466 (I27933,I27916,I26621);
nor I_1467 (I27950,I27933,I26615);
nor I_1468 (I27967,I26636,I26627);
DFFARX1 I_1469 (I27984,I27967,I2966,I27800,);
nor I_1470 (I28001,I27984,I27868);
not I_1471 (I28018,I27984);
nand I_1472 (I27774,I27851,I28018);
DFFARX1 I_1473 (I27765,I27984,I2966,I27800,);
nor I_1474 (I28063,I26636,I26612);
nand I_1475 (I28080,I27834,I28063);
nor I_1476 (I27789,I27817,I28063);
and I_1477 (I28111,I28063,I28001);
or I_1478 (I28128,I27950,I28111);
DFFARX1 I_1479 (I27777,I28128,I2966,I27800,);
DFFARX1 I_1480 (I28159,I26630,I2966,I27800,);
and I_1481 (I28176,I28159,I26633);
not I_1482 (I27783,I28176);
DFFARX1 I_1483 (I28207,I28176,I2966,I27800,);
not I_1484 (I27771,I28207);
and I_1485 (I28238,I28176,I27899);
DFFARX1 I_1486 (I27762,I28238,I2966,I27800,);
DFFARX1 I_1487 (I28269,I26606,I2966,I27800,);
and I_1488 (I28286,I28269,I28080);
DFFARX1 I_1489 (I27792,I28286,I2966,I27800,);
nor I_1490 (I28317,I28269,I28176);
nand I_1491 (I27786,I27950,I28317);
nor I_1492 (I28348,I28269,I28018);
nand I_1493 (I27780,I27834,I28348);
not I_1494 (I28412,I2973);
or I_1495 (I28429,I24256,I24241);
or I_1496 (I28446,I24250,I24256);
nor I_1497 (I28463,I24244,I24232);
or I_1498 (I28401,I28463,I28429);
not I_1499 (I28494,I24244);
and I_1500 (I28511,I28494,I24253);
nor I_1501 (I28528,I28511,I24241);
not I_1502 (I28545,I28528);
nor I_1503 (I28562,I24238,I24229);
DFFARX1 I_1504 (I28579,I28562,I2966,I28412,);
nor I_1505 (I28596,I28579,I28528);
nand I_1506 (I28386,I28429,I28596);
nor I_1507 (I28627,I28579,I28545);
not I_1508 (I28383,I28579);
nor I_1509 (I28658,I24238,I24250);
or I_1510 (I28395,I28429,I28658);
DFFARX1 I_1511 (I28689,I24247,I2966,I28412,);
and I_1512 (I28706,I28689,I24226);
nor I_1513 (I28723,I28706,I28579);
DFFARX1 I_1514 (I28389,I28723,I2966,I28412,);
nor I_1515 (I28404,I28706,I28658);
not I_1516 (I28768,I28706);
nor I_1517 (I28785,I28446,I28768);
nand I_1518 (I28374,I28706,I28545);
DFFARX1 I_1519 (I28816,I24235,I2966,I28412,);
nor I_1520 (I28392,I28816,I28446);
not I_1521 (I28847,I28816);
and I_1522 (I28864,I28658,I28847);
nor I_1523 (I28398,I28463,I28864);
and I_1524 (I28895,I28816,I28785);
or I_1525 (I28912,I28463,I28895);
DFFARX1 I_1526 (I28377,I28912,I2966,I28412,);
nand I_1527 (I28380,I28816,I28627);
not I_1528 (I28990,I2973);
or I_1529 (I29007,I12441,I12414);
or I_1530 (I29024,I12411,I12441);
nor I_1531 (I29041,I12423,I12435);
or I_1532 (I28979,I29041,I29007);
not I_1533 (I29072,I12423);
and I_1534 (I29089,I29072,I12429);
nor I_1535 (I29106,I29089,I12414);
not I_1536 (I29123,I29106);
nor I_1537 (I29140,I12417,I12438);
DFFARX1 I_1538 (I29157,I29140,I2966,I28990,);
nor I_1539 (I29174,I29157,I29106);
nand I_1540 (I28964,I29007,I29174);
nor I_1541 (I29205,I29157,I29123);
not I_1542 (I28961,I29157);
nor I_1543 (I29236,I12417,I12411);
or I_1544 (I28973,I29007,I29236);
DFFARX1 I_1545 (I29267,I12432,I2966,I28990,);
and I_1546 (I29284,I29267,I12420);
nor I_1547 (I29301,I29284,I29157);
DFFARX1 I_1548 (I28967,I29301,I2966,I28990,);
nor I_1549 (I28982,I29284,I29236);
not I_1550 (I29346,I29284);
nor I_1551 (I29363,I29024,I29346);
nand I_1552 (I28952,I29284,I29123);
DFFARX1 I_1553 (I29394,I12426,I2966,I28990,);
nor I_1554 (I28970,I29394,I29024);
not I_1555 (I29425,I29394);
and I_1556 (I29442,I29236,I29425);
nor I_1557 (I28976,I29041,I29442);
and I_1558 (I29473,I29394,I29363);
or I_1559 (I29490,I29041,I29473);
DFFARX1 I_1560 (I28955,I29490,I2966,I28990,);
nand I_1561 (I28958,I29394,I29205);
not I_1562 (I29568,I2973);
nand I_1563 (I29585,I15372,I15378);
and I_1564 (I29602,I29585,I15375);
DFFARX1 I_1565 (I29619,I29602,I2966,I29568,);
nor I_1566 (I29636,I15399,I15378);
nor I_1567 (I29653,I29636,I29619);
not I_1568 (I29551,I29636);
DFFARX1 I_1569 (I29684,I15390,I2966,I29568,);
not I_1570 (I29701,I29684);
nor I_1571 (I29718,I29636,I29701);
nand I_1572 (I29554,I29684,I29653);
DFFARX1 I_1573 (I29536,I29684,I2966,I29568,);
nand I_1574 (I29763,I15393,I15396);
and I_1575 (I29780,I29763,I15369);
DFFARX1 I_1576 (I29797,I29780,I2966,I29568,);
nor I_1577 (I29557,I29797,I29619);
nand I_1578 (I29548,I29797,I29718);
DFFARX1 I_1579 (I29842,I15387,I2966,I29568,);
and I_1580 (I29859,I29842,I15381);
DFFARX1 I_1581 (I29876,I29859,I2966,I29568,);
not I_1582 (I29539,I29876);
nand I_1583 (I29907,I29859,I29797);
and I_1584 (I29924,I29619,I29907);
DFFARX1 I_1585 (I29530,I29924,I2966,I29568,);
DFFARX1 I_1586 (I29955,I15384,I2966,I29568,);
nand I_1587 (I29972,I29955,I29619);
and I_1588 (I29989,I29797,I29972);
DFFARX1 I_1589 (I29560,I29989,I2966,I29568,);
not I_1590 (I30020,I29955);
nor I_1591 (I30037,I29636,I30020);
and I_1592 (I30054,I29955,I30037);
or I_1593 (I30071,I29859,I30054);
DFFARX1 I_1594 (I29545,I30071,I2966,I29568,);
nand I_1595 (I29542,I29955,I29701);
DFFARX1 I_1596 (I29533,I29955,I2966,I29568,);
not I_1597 (I30163,I2973);
nand I_1598 (I30180,I13004,I12995);
and I_1599 (I30197,I30180,I13013);
DFFARX1 I_1600 (I30214,I30197,I2966,I30163,);
nor I_1601 (I30231,I12992,I12995);
nor I_1602 (I30248,I30231,I30214);
not I_1603 (I30146,I30231);
DFFARX1 I_1604 (I30279,I13001,I2966,I30163,);
not I_1605 (I30296,I30279);
nor I_1606 (I30313,I30231,I30296);
nand I_1607 (I30149,I30279,I30248);
DFFARX1 I_1608 (I30131,I30279,I2966,I30163,);
nand I_1609 (I30358,I13016,I12998);
and I_1610 (I30375,I30358,I13019);
DFFARX1 I_1611 (I30392,I30375,I2966,I30163,);
nor I_1612 (I30152,I30392,I30214);
nand I_1613 (I30143,I30392,I30313);
DFFARX1 I_1614 (I30437,I13007,I2966,I30163,);
and I_1615 (I30454,I30437,I12989);
DFFARX1 I_1616 (I30471,I30454,I2966,I30163,);
not I_1617 (I30134,I30471);
nand I_1618 (I30502,I30454,I30392);
and I_1619 (I30519,I30214,I30502);
DFFARX1 I_1620 (I30125,I30519,I2966,I30163,);
DFFARX1 I_1621 (I30550,I13010,I2966,I30163,);
nand I_1622 (I30567,I30550,I30214);
and I_1623 (I30584,I30392,I30567);
DFFARX1 I_1624 (I30155,I30584,I2966,I30163,);
not I_1625 (I30615,I30550);
nor I_1626 (I30632,I30231,I30615);
and I_1627 (I30649,I30550,I30632);
or I_1628 (I30666,I30454,I30649);
DFFARX1 I_1629 (I30140,I30666,I2966,I30163,);
nand I_1630 (I30137,I30550,I30296);
DFFARX1 I_1631 (I30128,I30550,I2966,I30163,);
not I_1632 (I30758,I2973);
nand I_1633 (I30775,I19008,I19020);
and I_1634 (I30792,I30775,I18999);
DFFARX1 I_1635 (I30809,I30792,I2966,I30758,);
nor I_1636 (I30826,I18990,I19020);
nor I_1637 (I30843,I30826,I30809);
not I_1638 (I30741,I30826);
DFFARX1 I_1639 (I30874,I19002,I2966,I30758,);
not I_1640 (I30891,I30874);
nor I_1641 (I30908,I30826,I30891);
nand I_1642 (I30744,I30874,I30843);
DFFARX1 I_1643 (I30726,I30874,I2966,I30758,);
nand I_1644 (I30953,I19017,I19005);
and I_1645 (I30970,I30953,I18993);
DFFARX1 I_1646 (I30987,I30970,I2966,I30758,);
nor I_1647 (I30747,I30987,I30809);
nand I_1648 (I30738,I30987,I30908);
DFFARX1 I_1649 (I31032,I19011,I2966,I30758,);
and I_1650 (I31049,I31032,I18996);
DFFARX1 I_1651 (I31066,I31049,I2966,I30758,);
not I_1652 (I30729,I31066);
nand I_1653 (I31097,I31049,I30987);
and I_1654 (I31114,I30809,I31097);
DFFARX1 I_1655 (I30720,I31114,I2966,I30758,);
DFFARX1 I_1656 (I31145,I19014,I2966,I30758,);
nand I_1657 (I31162,I31145,I30809);
and I_1658 (I31179,I30987,I31162);
DFFARX1 I_1659 (I30750,I31179,I2966,I30758,);
not I_1660 (I31210,I31145);
nor I_1661 (I31227,I30826,I31210);
and I_1662 (I31244,I31145,I31227);
or I_1663 (I31261,I31049,I31244);
DFFARX1 I_1664 (I30735,I31261,I2966,I30758,);
nand I_1665 (I30732,I31145,I30891);
DFFARX1 I_1666 (I30723,I31145,I2966,I30758,);
not I_1667 (I31353,I2973);
nand I_1668 (I31370,I15933,I15939);
and I_1669 (I31387,I31370,I15936);
DFFARX1 I_1670 (I31404,I31387,I2966,I31353,);
nor I_1671 (I31421,I15960,I15939);
nor I_1672 (I31438,I31421,I31404);
not I_1673 (I31336,I31421);
DFFARX1 I_1674 (I31469,I15951,I2966,I31353,);
not I_1675 (I31486,I31469);
nor I_1676 (I31503,I31421,I31486);
nand I_1677 (I31339,I31469,I31438);
DFFARX1 I_1678 (I31321,I31469,I2966,I31353,);
nand I_1679 (I31548,I15954,I15957);
and I_1680 (I31565,I31548,I15930);
DFFARX1 I_1681 (I31582,I31565,I2966,I31353,);
nor I_1682 (I31342,I31582,I31404);
nand I_1683 (I31333,I31582,I31503);
DFFARX1 I_1684 (I31627,I15948,I2966,I31353,);
and I_1685 (I31644,I31627,I15942);
DFFARX1 I_1686 (I31661,I31644,I2966,I31353,);
not I_1687 (I31324,I31661);
nand I_1688 (I31692,I31644,I31582);
and I_1689 (I31709,I31404,I31692);
DFFARX1 I_1690 (I31315,I31709,I2966,I31353,);
DFFARX1 I_1691 (I31740,I15945,I2966,I31353,);
nand I_1692 (I31757,I31740,I31404);
and I_1693 (I31774,I31582,I31757);
DFFARX1 I_1694 (I31345,I31774,I2966,I31353,);
not I_1695 (I31805,I31740);
nor I_1696 (I31822,I31421,I31805);
and I_1697 (I31839,I31740,I31822);
or I_1698 (I31856,I31644,I31839);
DFFARX1 I_1699 (I31330,I31856,I2966,I31353,);
nand I_1700 (I31327,I31740,I31486);
DFFARX1 I_1701 (I31318,I31740,I2966,I31353,);
not I_1702 (I31948,I2973);
nand I_1703 (I31965,I7227,I7233);
and I_1704 (I31982,I31965,I7215);
DFFARX1 I_1705 (I31999,I31982,I2966,I31948,);
nor I_1706 (I32016,I7209,I7233);
nor I_1707 (I32033,I32016,I31999);
not I_1708 (I31931,I32016);
DFFARX1 I_1709 (I32064,I7239,I2966,I31948,);
not I_1710 (I32081,I32064);
nor I_1711 (I32098,I32016,I32081);
nand I_1712 (I31934,I32064,I32033);
DFFARX1 I_1713 (I31916,I32064,I2966,I31948,);
nand I_1714 (I32143,I7230,I7221);
and I_1715 (I32160,I32143,I7224);
DFFARX1 I_1716 (I32177,I32160,I2966,I31948,);
nor I_1717 (I31937,I32177,I31999);
nand I_1718 (I31928,I32177,I32098);
DFFARX1 I_1719 (I32222,I7236,I2966,I31948,);
and I_1720 (I32239,I32222,I7212);
DFFARX1 I_1721 (I32256,I32239,I2966,I31948,);
not I_1722 (I31919,I32256);
nand I_1723 (I32287,I32239,I32177);
and I_1724 (I32304,I31999,I32287);
DFFARX1 I_1725 (I31910,I32304,I2966,I31948,);
DFFARX1 I_1726 (I32335,I7218,I2966,I31948,);
nand I_1727 (I32352,I32335,I31999);
and I_1728 (I32369,I32177,I32352);
DFFARX1 I_1729 (I31940,I32369,I2966,I31948,);
not I_1730 (I32400,I32335);
nor I_1731 (I32417,I32016,I32400);
and I_1732 (I32434,I32335,I32417);
or I_1733 (I32451,I32239,I32434);
DFFARX1 I_1734 (I31925,I32451,I2966,I31948,);
nand I_1735 (I31922,I32335,I32081);
DFFARX1 I_1736 (I31913,I32335,I2966,I31948,);
not I_1737 (I32543,I2973);
nand I_1738 (I32560,I22267,I22237);
and I_1739 (I32577,I32560,I22255);
DFFARX1 I_1740 (I32594,I32577,I2966,I32543,);
nor I_1741 (I32611,I22249,I22237);
DFFARX1 I_1742 (I32628,I22246,I2966,I32543,);
nand I_1743 (I32645,I32628,I32611);
DFFARX1 I_1744 (I32514,I32628,I2966,I32543,);
nand I_1745 (I32676,I22240,I22243);
and I_1746 (I32693,I32676,I22261);
DFFARX1 I_1747 (I32710,I32693,I2966,I32543,);
not I_1748 (I32727,I32710);
nor I_1749 (I32744,I32594,I32727);
and I_1750 (I32761,I32611,I32744);
and I_1751 (I32778,I32710,I32645);
DFFARX1 I_1752 (I32511,I32778,I2966,I32543,);
DFFARX1 I_1753 (I32505,I32710,I2966,I32543,);
DFFARX1 I_1754 (I32823,I22264,I2966,I32543,);
and I_1755 (I32840,I32823,I22258);
nand I_1756 (I32857,I32840,I32710);
nor I_1757 (I32532,I32840,I32611);
not I_1758 (I32888,I32840);
nor I_1759 (I32905,I32594,I32888);
nand I_1760 (I32523,I32628,I32905);
nand I_1761 (I32517,I32710,I32888);
or I_1762 (I32950,I32840,I32761);
DFFARX1 I_1763 (I32520,I32950,I2966,I32543,);
DFFARX1 I_1764 (I32981,I22252,I2966,I32543,);
and I_1765 (I32998,I32981,I32857);
DFFARX1 I_1766 (I32535,I32998,I2966,I32543,);
nor I_1767 (I33029,I32981,I32594);
nand I_1768 (I32529,I32840,I33029);
not I_1769 (I32526,I32981);
DFFARX1 I_1770 (I33074,I32981,I2966,I32543,);
and I_1771 (I32508,I32981,I33074);
not I_1772 (I33138,I2973);
not I_1773 (I33155,I27774);
nor I_1774 (I33172,I27765,I27792);
nand I_1775 (I33189,I33172,I27762);
nor I_1776 (I33206,I33155,I27765);
nand I_1777 (I33223,I33206,I27786);
not I_1778 (I33240,I27765);
not I_1779 (I33257,I33240);
not I_1780 (I33274,I27771);
nor I_1781 (I33291,I33274,I27789);
and I_1782 (I33308,I33291,I27780);
or I_1783 (I33325,I33308,I27777);
DFFARX1 I_1784 (I33342,I33325,I2966,I33138,);
nand I_1785 (I33359,I33155,I27771);
or I_1786 (I33127,I33359,I33342);
not I_1787 (I33390,I33359);
nor I_1788 (I33407,I33342,I33390);
and I_1789 (I33424,I33240,I33407);
nand I_1790 (I33100,I33359,I33257);
DFFARX1 I_1791 (I33455,I27768,I2966,I33138,);
or I_1792 (I33121,I33455,I33342);
nor I_1793 (I33486,I33455,I33223);
nor I_1794 (I33503,I33455,I33257);
nand I_1795 (I33106,I33189,I33503);
or I_1796 (I33534,I33455,I33424);
DFFARX1 I_1797 (I33103,I33534,I2966,I33138,);
not I_1798 (I33109,I33455);
DFFARX1 I_1799 (I33579,I27783,I2966,I33138,);
not I_1800 (I33596,I33579);
nor I_1801 (I33613,I33596,I33189);
DFFARX1 I_1802 (I33115,I33613,I2966,I33138,);
nor I_1803 (I33130,I33455,I33596);
nor I_1804 (I33118,I33596,I33359);
not I_1805 (I33672,I33596);
and I_1806 (I33689,I33223,I33672);
nor I_1807 (I33124,I33359,I33689);
nand I_1808 (I33112,I33596,I33486);
not I_1809 (I33767,I2973);
not I_1810 (I33784,I11171);
nor I_1811 (I33801,I11180,I11183);
nand I_1812 (I33818,I33801,I11168);
nor I_1813 (I33835,I33784,I11180);
nand I_1814 (I33852,I33835,I11165);
not I_1815 (I33869,I11180);
not I_1816 (I33886,I33869);
not I_1817 (I33903,I11153);
nor I_1818 (I33920,I33903,I11159);
and I_1819 (I33937,I33920,I11156);
or I_1820 (I33954,I33937,I11177);
DFFARX1 I_1821 (I33971,I33954,I2966,I33767,);
nand I_1822 (I33988,I33784,I11153);
or I_1823 (I33756,I33988,I33971);
not I_1824 (I34019,I33988);
nor I_1825 (I34036,I33971,I34019);
and I_1826 (I34053,I33869,I34036);
nand I_1827 (I33729,I33988,I33886);
DFFARX1 I_1828 (I34084,I11162,I2966,I33767,);
or I_1829 (I33750,I34084,I33971);
nor I_1830 (I34115,I34084,I33852);
nor I_1831 (I34132,I34084,I33886);
nand I_1832 (I33735,I33818,I34132);
or I_1833 (I34163,I34084,I34053);
DFFARX1 I_1834 (I33732,I34163,I2966,I33767,);
not I_1835 (I33738,I34084);
DFFARX1 I_1836 (I34208,I11174,I2966,I33767,);
not I_1837 (I34225,I34208);
nor I_1838 (I34242,I34225,I33818);
DFFARX1 I_1839 (I33744,I34242,I2966,I33767,);
nor I_1840 (I33759,I34084,I34225);
nor I_1841 (I33747,I34225,I33988);
not I_1842 (I34301,I34225);
and I_1843 (I34318,I33852,I34301);
nor I_1844 (I33753,I33988,I34318);
nand I_1845 (I33741,I34225,I34115);
not I_1846 (I34396,I2973);
not I_1847 (I34413,I14797);
nor I_1848 (I34430,I14821,I14806);
nand I_1849 (I34447,I34430,I14791);
nor I_1850 (I34464,I34413,I14821);
nand I_1851 (I34481,I34464,I14818);
not I_1852 (I34498,I14821);
not I_1853 (I34515,I34498);
not I_1854 (I34532,I14800);
nor I_1855 (I34549,I34532,I14794);
and I_1856 (I34566,I34549,I14815);
or I_1857 (I34583,I34566,I14803);
DFFARX1 I_1858 (I34600,I34583,I2966,I34396,);
nand I_1859 (I34617,I34413,I14800);
or I_1860 (I34385,I34617,I34600);
not I_1861 (I34648,I34617);
nor I_1862 (I34665,I34600,I34648);
and I_1863 (I34682,I34498,I34665);
nand I_1864 (I34358,I34617,I34515);
DFFARX1 I_1865 (I34713,I14812,I2966,I34396,);
or I_1866 (I34379,I34713,I34600);
nor I_1867 (I34744,I34713,I34481);
nor I_1868 (I34761,I34713,I34515);
nand I_1869 (I34364,I34447,I34761);
or I_1870 (I34792,I34713,I34682);
DFFARX1 I_1871 (I34361,I34792,I2966,I34396,);
not I_1872 (I34367,I34713);
DFFARX1 I_1873 (I34837,I14809,I2966,I34396,);
not I_1874 (I34854,I34837);
nor I_1875 (I34871,I34854,I34447);
DFFARX1 I_1876 (I34373,I34871,I2966,I34396,);
nor I_1877 (I34388,I34713,I34854);
nor I_1878 (I34376,I34854,I34617);
not I_1879 (I34930,I34854);
and I_1880 (I34947,I34481,I34930);
nor I_1881 (I34382,I34617,I34947);
nand I_1882 (I34370,I34854,I34744);
not I_1883 (I35025,I2973);
not I_1884 (I35042,I26058);
nor I_1885 (I35059,I26031,I26049);
nand I_1886 (I35076,I35059,I26034);
nor I_1887 (I35093,I35042,I26031);
nand I_1888 (I35110,I35093,I26052);
not I_1889 (I35127,I26031);
not I_1890 (I35144,I35127);
not I_1891 (I35161,I26028);
nor I_1892 (I35178,I35161,I26055);
and I_1893 (I35195,I35178,I26046);
or I_1894 (I35212,I35195,I26037);
DFFARX1 I_1895 (I35229,I35212,I2966,I35025,);
nand I_1896 (I35246,I35042,I26028);
or I_1897 (I35014,I35246,I35229);
not I_1898 (I35277,I35246);
nor I_1899 (I35294,I35229,I35277);
and I_1900 (I35311,I35127,I35294);
nand I_1901 (I34987,I35246,I35144);
DFFARX1 I_1902 (I35342,I26040,I2966,I35025,);
or I_1903 (I35008,I35342,I35229);
nor I_1904 (I35373,I35342,I35110);
nor I_1905 (I35390,I35342,I35144);
nand I_1906 (I34993,I35076,I35390);
or I_1907 (I35421,I35342,I35311);
DFFARX1 I_1908 (I34990,I35421,I2966,I35025,);
not I_1909 (I34996,I35342);
DFFARX1 I_1910 (I35466,I26043,I2966,I35025,);
not I_1911 (I35483,I35466);
nor I_1912 (I35500,I35483,I35076);
DFFARX1 I_1913 (I35002,I35500,I2966,I35025,);
nor I_1914 (I35017,I35342,I35483);
nor I_1915 (I35005,I35483,I35246);
not I_1916 (I35559,I35483);
and I_1917 (I35576,I35110,I35559);
nor I_1918 (I35011,I35246,I35576);
nand I_1919 (I34999,I35483,I35373);
not I_1920 (I35654,I2973);
not I_1921 (I35671,I14219);
nor I_1922 (I35688,I14243,I14228);
nand I_1923 (I35705,I35688,I14213);
nor I_1924 (I35722,I35671,I14243);
nand I_1925 (I35739,I35722,I14240);
not I_1926 (I35756,I14243);
not I_1927 (I35773,I35756);
not I_1928 (I35790,I14222);
nor I_1929 (I35807,I35790,I14216);
and I_1930 (I35824,I35807,I14237);
or I_1931 (I35841,I35824,I14225);
DFFARX1 I_1932 (I35858,I35841,I2966,I35654,);
nand I_1933 (I35875,I35671,I14222);
or I_1934 (I35643,I35875,I35858);
not I_1935 (I35906,I35875);
nor I_1936 (I35923,I35858,I35906);
and I_1937 (I35940,I35756,I35923);
nand I_1938 (I35616,I35875,I35773);
DFFARX1 I_1939 (I35971,I14234,I2966,I35654,);
or I_1940 (I35637,I35971,I35858);
nor I_1941 (I36002,I35971,I35739);
nor I_1942 (I36019,I35971,I35773);
nand I_1943 (I35622,I35705,I36019);
or I_1944 (I36050,I35971,I35940);
DFFARX1 I_1945 (I35619,I36050,I2966,I35654,);
not I_1946 (I35625,I35971);
DFFARX1 I_1947 (I36095,I14231,I2966,I35654,);
not I_1948 (I36112,I36095);
nor I_1949 (I36129,I36112,I35705);
DFFARX1 I_1950 (I35631,I36129,I2966,I35654,);
nor I_1951 (I35646,I35971,I36112);
nor I_1952 (I35634,I36112,I35875);
not I_1953 (I36188,I36112);
and I_1954 (I36205,I35739,I36188);
nor I_1955 (I35640,I35875,I36205);
nand I_1956 (I35628,I36112,I36002);
not I_1957 (I36283,I2973);
nand I_1958 (I36300,I23572,I23569);
and I_1959 (I36317,I36300,I23593);
DFFARX1 I_1960 (I36334,I36317,I2966,I36283,);
not I_1961 (I36272,I36334);
DFFARX1 I_1962 (I36365,I36334,I2966,I36283,);
not I_1963 (I36260,I36365);
nor I_1964 (I36396,I23575,I23569);
not I_1965 (I36413,I36396);
nor I_1966 (I36430,I36334,I36413);
DFFARX1 I_1967 (I36447,I23590,I2966,I36283,);
not I_1968 (I36464,I36447);
nand I_1969 (I36263,I36447,I36413);
DFFARX1 I_1970 (I36495,I36447,I2966,I36283,);
and I_1971 (I36248,I36334,I36495);
nand I_1972 (I36526,I23578,I23563);
and I_1973 (I36543,I36526,I23581);
DFFARX1 I_1974 (I36560,I36543,I2966,I36283,);
nor I_1975 (I36577,I36560,I36464);
and I_1976 (I36594,I36396,I36577);
nor I_1977 (I36611,I36560,I36334);
DFFARX1 I_1978 (I36254,I36560,I2966,I36283,);
DFFARX1 I_1979 (I36642,I23584,I2966,I36283,);
and I_1980 (I36659,I36642,I23587);
or I_1981 (I36676,I36659,I36594);
DFFARX1 I_1982 (I36266,I36676,I2966,I36283,);
nand I_1983 (I36275,I36659,I36611);
DFFARX1 I_1984 (I36245,I36659,I2966,I36283,);
DFFARX1 I_1985 (I36735,I23566,I2966,I36283,);
nand I_1986 (I36269,I36735,I36430);
DFFARX1 I_1987 (I36257,I36735,I2966,I36283,);
nand I_1988 (I36780,I36735,I36396);
and I_1989 (I36797,I36447,I36780);
DFFARX1 I_1990 (I36251,I36797,I2966,I36283,);
not I_1991 (I36861,I2973);
not I_1992 (I36878,I22918);
nor I_1993 (I36895,I22915,I22903);
nand I_1994 (I36912,I36895,I22906);
DFFARX1 I_1995 (I36835,I36912,I2966,I36861,);
nor I_1996 (I36943,I36878,I22915);
nand I_1997 (I36960,I36943,I22912);
not I_1998 (I36850,I36960);
DFFARX1 I_1999 (I36832,I36960,I2966,I36861,);
not I_2000 (I37005,I22915);
not I_2001 (I37022,I37005);
not I_2002 (I37039,I22924);
nor I_2003 (I37056,I37039,I22900);
and I_2004 (I37073,I37056,I22921);
or I_2005 (I37090,I37073,I22909);
DFFARX1 I_2006 (I37107,I37090,I2966,I36861,);
nor I_2007 (I37124,I37107,I36960);
nor I_2008 (I37141,I37107,I37022);
nand I_2009 (I36847,I36912,I37141);
nand I_2010 (I37172,I36878,I22924);
nand I_2011 (I37189,I37172,I37107);
and I_2012 (I37206,I37172,I37189);
DFFARX1 I_2013 (I36829,I37206,I2966,I36861,);
DFFARX1 I_2014 (I37237,I37172,I2966,I36861,);
and I_2015 (I36826,I37005,I37237);
DFFARX1 I_2016 (I37268,I22930,I2966,I36861,);
not I_2017 (I37285,I37268);
nor I_2018 (I37302,I36960,I37285);
and I_2019 (I37319,I37268,I37302);
nand I_2020 (I36841,I37268,I37022);
DFFARX1 I_2021 (I37350,I37268,I2966,I36861,);
not I_2022 (I36838,I37350);
DFFARX1 I_2023 (I37381,I22927,I2966,I36861,);
not I_2024 (I37398,I37381);
or I_2025 (I37415,I37398,I37319);
DFFARX1 I_2026 (I36844,I37415,I2966,I36861,);
nand I_2027 (I36853,I37398,I37124);
DFFARX1 I_2028 (I36823,I37398,I2966,I36861,);
not I_2029 (I37507,I2973);
not I_2030 (I37524,I20911);
nor I_2031 (I37541,I20920,I20932);
nand I_2032 (I37558,I37541,I20923);
DFFARX1 I_2033 (I37478,I37558,I2966,I37507,);
nor I_2034 (I37589,I37524,I20920);
nand I_2035 (I37606,I37589,I20935);
nand I_2036 (I37623,I37606,I37558);
not I_2037 (I37640,I20920);
not I_2038 (I37657,I20941);
nor I_2039 (I37674,I37657,I20917);
and I_2040 (I37691,I37674,I20926);
or I_2041 (I37708,I37691,I20914);
DFFARX1 I_2042 (I37725,I37708,I2966,I37507,);
nor I_2043 (I37742,I37725,I37606);
nand I_2044 (I37493,I37640,I37742);
not I_2045 (I37490,I37725);
and I_2046 (I37787,I37725,I37623);
DFFARX1 I_2047 (I37475,I37787,I2966,I37507,);
DFFARX1 I_2048 (I37818,I37725,I2966,I37507,);
and I_2049 (I37472,I37640,I37818);
nand I_2050 (I37849,I37524,I20941);
not I_2051 (I37866,I37849);
nor I_2052 (I37883,I37725,I37866);
DFFARX1 I_2053 (I37900,I20938,I2966,I37507,);
nand I_2054 (I37917,I37900,I37849);
and I_2055 (I37934,I37640,I37917);
DFFARX1 I_2056 (I37499,I37934,I2966,I37507,);
not I_2057 (I37965,I37900);
nand I_2058 (I37487,I37900,I37883);
nand I_2059 (I37481,I37900,I37866);
DFFARX1 I_2060 (I38010,I20929,I2966,I37507,);
not I_2061 (I38027,I38010);
nor I_2062 (I37496,I37900,I38027);
nor I_2063 (I38058,I38027,I37965);
and I_2064 (I38075,I37606,I38058);
or I_2065 (I38092,I37849,I38075);
DFFARX1 I_2066 (I37484,I38092,I2966,I37507,);
DFFARX1 I_2067 (I37469,I38027,I2966,I37507,);
not I_2068 (I38170,I2973);
not I_2069 (I38187,I30735);
nor I_2070 (I38204,I30747,I30750);
nand I_2071 (I38221,I38204,I30738);
DFFARX1 I_2072 (I38141,I38221,I2966,I38170,);
nor I_2073 (I38252,I38187,I30747);
nand I_2074 (I38269,I38252,I30723);
nand I_2075 (I38286,I38269,I38221);
not I_2076 (I38303,I30747);
not I_2077 (I38320,I30726);
nor I_2078 (I38337,I38320,I30729);
and I_2079 (I38354,I38337,I30732);
or I_2080 (I38371,I38354,I30741);
DFFARX1 I_2081 (I38388,I38371,I2966,I38170,);
nor I_2082 (I38405,I38388,I38269);
nand I_2083 (I38156,I38303,I38405);
not I_2084 (I38153,I38388);
and I_2085 (I38450,I38388,I38286);
DFFARX1 I_2086 (I38138,I38450,I2966,I38170,);
DFFARX1 I_2087 (I38481,I38388,I2966,I38170,);
and I_2088 (I38135,I38303,I38481);
nand I_2089 (I38512,I38187,I30726);
not I_2090 (I38529,I38512);
nor I_2091 (I38546,I38388,I38529);
DFFARX1 I_2092 (I38563,I30744,I2966,I38170,);
nand I_2093 (I38580,I38563,I38512);
and I_2094 (I38597,I38303,I38580);
DFFARX1 I_2095 (I38162,I38597,I2966,I38170,);
not I_2096 (I38628,I38563);
nand I_2097 (I38150,I38563,I38546);
nand I_2098 (I38144,I38563,I38529);
DFFARX1 I_2099 (I38673,I30720,I2966,I38170,);
not I_2100 (I38690,I38673);
nor I_2101 (I38159,I38563,I38690);
nor I_2102 (I38721,I38690,I38628);
and I_2103 (I38738,I38269,I38721);
or I_2104 (I38755,I38512,I38738);
DFFARX1 I_2105 (I38147,I38755,I2966,I38170,);
DFFARX1 I_2106 (I38132,I38690,I2966,I38170,);
not I_2107 (I38833,I2973);
or I_2108 (I38850,I36245,I36263);
or I_2109 (I38867,I36248,I36245);
DFFARX1 I_2110 (I38807,I38867,I2966,I38833,);
nor I_2111 (I38898,I36257,I36260);
not I_2112 (I38915,I38898);
not I_2113 (I38932,I36257);
and I_2114 (I38949,I38932,I36266);
nor I_2115 (I38966,I38949,I36263);
nor I_2116 (I38983,I36272,I36251);
DFFARX1 I_2117 (I39000,I38983,I2966,I38833,);
nand I_2118 (I39017,I39000,I38850);
and I_2119 (I39034,I38966,I39017);
DFFARX1 I_2120 (I38801,I39034,I2966,I38833,);
nor I_2121 (I39065,I36272,I36248);
DFFARX1 I_2122 (I39082,I39065,I2966,I38833,);
and I_2123 (I38798,I38898,I39082);
DFFARX1 I_2124 (I39113,I36275,I2966,I38833,);
and I_2125 (I39130,I39113,I36269);
DFFARX1 I_2126 (I39147,I39130,I2966,I38833,);
not I_2127 (I38810,I39147);
DFFARX1 I_2128 (I38795,I39130,I2966,I38833,);
DFFARX1 I_2129 (I39192,I36254,I2966,I38833,);
not I_2130 (I39209,I39192);
nor I_2131 (I39226,I38867,I39209);
and I_2132 (I39243,I39130,I39226);
or I_2133 (I39260,I38850,I39243);
DFFARX1 I_2134 (I38816,I39260,I2966,I38833,);
nor I_2135 (I39291,I39192,I39000);
nand I_2136 (I38825,I38966,I39291);
nor I_2137 (I39322,I39192,I38915);
nand I_2138 (I38819,I39065,I39322);
not I_2139 (I38822,I39192);
nand I_2140 (I38813,I39192,I38915);
DFFARX1 I_2141 (I38804,I39192,I2966,I38833,);
not I_2142 (I39428,I2973);
or I_2143 (I39445,I30131,I30143);
not I_2144 (I39411,I39445);
DFFARX1 I_2145 (I39390,I39445,I2966,I39428,);
or I_2146 (I39490,I30155,I30131);
nor I_2147 (I39507,I30149,I30134);
nor I_2148 (I39524,I39507,I39445);
not I_2149 (I39541,I30149);
and I_2150 (I39558,I39541,I30146);
nor I_2151 (I39575,I39558,I30143);
DFFARX1 I_2152 (I39592,I39575,I2966,I39428,);
nor I_2153 (I39609,I30140,I30137);
DFFARX1 I_2154 (I39626,I39609,I2966,I39428,);
nor I_2155 (I39417,I39626,I39575);
not I_2156 (I39657,I39626);
nor I_2157 (I39674,I30140,I30155);
nand I_2158 (I39691,I39575,I39674);
and I_2159 (I39708,I39490,I39691);
DFFARX1 I_2160 (I39420,I39708,I2966,I39428,);
DFFARX1 I_2161 (I39739,I30152,I2966,I39428,);
and I_2162 (I39756,I39739,I30125);
nor I_2163 (I39773,I39756,I39657);
and I_2164 (I39790,I39674,I39773);
or I_2165 (I39807,I39507,I39790);
DFFARX1 I_2166 (I39405,I39807,I2966,I39428,);
not I_2167 (I39838,I39756);
nor I_2168 (I39855,I39445,I39838);
nand I_2169 (I39408,I39490,I39855);
nand I_2170 (I39402,I39626,I39838);
DFFARX1 I_2171 (I39396,I39756,I2966,I39428,);
DFFARX1 I_2172 (I39914,I30128,I2966,I39428,);
nand I_2173 (I39414,I39914,I39524);
DFFARX1 I_2174 (I39945,I39914,I2966,I39428,);
not I_2175 (I39399,I39945);
and I_2176 (I39393,I39914,I39592);
not I_2177 (I40023,I2973);
or I_2178 (I40040,I21589,I21577);
not I_2179 (I40006,I40040);
DFFARX1 I_2180 (I39985,I40040,I2966,I40023,);
or I_2181 (I40085,I21574,I21589);
nor I_2182 (I40102,I21604,I21595);
nor I_2183 (I40119,I40102,I40040);
not I_2184 (I40136,I21604);
and I_2185 (I40153,I40136,I21583);
nor I_2186 (I40170,I40153,I21577);
DFFARX1 I_2187 (I40187,I40170,I2966,I40023,);
nor I_2188 (I40204,I21586,I21580);
DFFARX1 I_2189 (I40221,I40204,I2966,I40023,);
nor I_2190 (I40012,I40221,I40170);
not I_2191 (I40252,I40221);
nor I_2192 (I40269,I21586,I21574);
nand I_2193 (I40286,I40170,I40269);
and I_2194 (I40303,I40085,I40286);
DFFARX1 I_2195 (I40015,I40303,I2966,I40023,);
DFFARX1 I_2196 (I40334,I21601,I2966,I40023,);
and I_2197 (I40351,I40334,I21598);
nor I_2198 (I40368,I40351,I40252);
and I_2199 (I40385,I40269,I40368);
or I_2200 (I40402,I40102,I40385);
DFFARX1 I_2201 (I40000,I40402,I2966,I40023,);
not I_2202 (I40433,I40351);
nor I_2203 (I40450,I40040,I40433);
nand I_2204 (I40003,I40085,I40450);
nand I_2205 (I39997,I40221,I40433);
DFFARX1 I_2206 (I39991,I40351,I2966,I40023,);
DFFARX1 I_2207 (I40509,I21592,I2966,I40023,);
nand I_2208 (I40009,I40509,I40119);
DFFARX1 I_2209 (I40540,I40509,I2966,I40023,);
not I_2210 (I39994,I40540);
and I_2211 (I39988,I40509,I40187);
not I_2212 (I40618,I2973);
or I_2213 (I40635,I31916,I31928);
not I_2214 (I40601,I40635);
DFFARX1 I_2215 (I40580,I40635,I2966,I40618,);
or I_2216 (I40680,I31940,I31916);
nor I_2217 (I40697,I31934,I31919);
nor I_2218 (I40714,I40697,I40635);
not I_2219 (I40731,I31934);
and I_2220 (I40748,I40731,I31931);
nor I_2221 (I40765,I40748,I31928);
DFFARX1 I_2222 (I40782,I40765,I2966,I40618,);
nor I_2223 (I40799,I31925,I31922);
DFFARX1 I_2224 (I40816,I40799,I2966,I40618,);
nor I_2225 (I40607,I40816,I40765);
not I_2226 (I40847,I40816);
nor I_2227 (I40864,I31925,I31940);
nand I_2228 (I40881,I40765,I40864);
and I_2229 (I40898,I40680,I40881);
DFFARX1 I_2230 (I40610,I40898,I2966,I40618,);
DFFARX1 I_2231 (I40929,I31937,I2966,I40618,);
and I_2232 (I40946,I40929,I31910);
nor I_2233 (I40963,I40946,I40847);
and I_2234 (I40980,I40864,I40963);
or I_2235 (I40997,I40697,I40980);
DFFARX1 I_2236 (I40595,I40997,I2966,I40618,);
not I_2237 (I41028,I40946);
nor I_2238 (I41045,I40635,I41028);
nand I_2239 (I40598,I40680,I41045);
nand I_2240 (I40592,I40816,I41028);
DFFARX1 I_2241 (I40586,I40946,I2966,I40618,);
DFFARX1 I_2242 (I41104,I31913,I2966,I40618,);
nand I_2243 (I40604,I41104,I40714);
DFFARX1 I_2244 (I41135,I41104,I2966,I40618,);
not I_2245 (I40589,I41135);
and I_2246 (I40583,I41104,I40782);
not I_2247 (I41213,I2973);
not I_2248 (I41230,I29548);
nor I_2249 (I41247,I29557,I29539);
nand I_2250 (I41264,I41247,I29560);
nor I_2251 (I41281,I41230,I29557);
nand I_2252 (I41298,I41281,I29551);
not I_2253 (I41315,I41298);
not I_2254 (I41332,I29557);
nor I_2255 (I41202,I41298,I41332);
not I_2256 (I41363,I41332);
nand I_2257 (I41187,I41298,I41363);
not I_2258 (I41394,I29545);
nor I_2259 (I41411,I41394,I29536);
and I_2260 (I41428,I41411,I29533);
or I_2261 (I41445,I41428,I29530);
DFFARX1 I_2262 (I41462,I41445,I2966,I41213,);
nor I_2263 (I41479,I41462,I41315);
DFFARX1 I_2264 (I41496,I41462,I2966,I41213,);
not I_2265 (I41184,I41496);
nand I_2266 (I41527,I41230,I29545);
and I_2267 (I41544,I41527,I41479);
DFFARX1 I_2268 (I41181,I41527,I2966,I41213,);
DFFARX1 I_2269 (I41575,I29554,I2966,I41213,);
nor I_2270 (I41592,I41575,I41298);
nand I_2271 (I41199,I41462,I41592);
nor I_2272 (I41623,I41575,I41363);
not I_2273 (I41196,I41575);
nand I_2274 (I41654,I41575,I41264);
and I_2275 (I41671,I41332,I41654);
DFFARX1 I_2276 (I41175,I41671,I2966,I41213,);
DFFARX1 I_2277 (I41178,I41575,I2966,I41213,);
DFFARX1 I_2278 (I41716,I29542,I2966,I41213,);
not I_2279 (I41733,I41716);
nand I_2280 (I41750,I41733,I41298);
and I_2281 (I41767,I41527,I41750);
DFFARX1 I_2282 (I41205,I41767,I2966,I41213,);
or I_2283 (I41798,I41733,I41544);
DFFARX1 I_2284 (I41190,I41798,I2966,I41213,);
nand I_2285 (I41193,I41733,I41623);
not I_2286 (I41876,I2973);
not I_2287 (I41893,I28377);
nor I_2288 (I41910,I28398,I28404);
nand I_2289 (I41927,I41910,I28392);
nor I_2290 (I41944,I41893,I28398);
nand I_2291 (I41961,I41944,I28374);
not I_2292 (I41978,I41961);
not I_2293 (I41995,I28398);
nor I_2294 (I41865,I41961,I41995);
not I_2295 (I42026,I41995);
nand I_2296 (I41850,I41961,I42026);
not I_2297 (I42057,I28380);
nor I_2298 (I42074,I42057,I28401);
and I_2299 (I42091,I42074,I28389);
or I_2300 (I42108,I42091,I28395);
DFFARX1 I_2301 (I42125,I42108,I2966,I41876,);
nor I_2302 (I42142,I42125,I41978);
DFFARX1 I_2303 (I42159,I42125,I2966,I41876,);
not I_2304 (I41847,I42159);
nand I_2305 (I42190,I41893,I28380);
and I_2306 (I42207,I42190,I42142);
DFFARX1 I_2307 (I41844,I42190,I2966,I41876,);
DFFARX1 I_2308 (I42238,I28386,I2966,I41876,);
nor I_2309 (I42255,I42238,I41961);
nand I_2310 (I41862,I42125,I42255);
nor I_2311 (I42286,I42238,I42026);
not I_2312 (I41859,I42238);
nand I_2313 (I42317,I42238,I41927);
and I_2314 (I42334,I41995,I42317);
DFFARX1 I_2315 (I41838,I42334,I2966,I41876,);
DFFARX1 I_2316 (I41841,I42238,I2966,I41876,);
DFFARX1 I_2317 (I42379,I28383,I2966,I41876,);
not I_2318 (I42396,I42379);
nand I_2319 (I42413,I42396,I41961);
and I_2320 (I42430,I42190,I42413);
DFFARX1 I_2321 (I41868,I42430,I2966,I41876,);
or I_2322 (I42461,I42396,I42207);
DFFARX1 I_2323 (I41853,I42461,I2966,I41876,);
nand I_2324 (I41856,I42396,I42286);
not I_2325 (I42539,I2973);
not I_2326 (I42556,I37472);
nor I_2327 (I42573,I37478,I37484);
nand I_2328 (I42590,I42573,I37487);
nor I_2329 (I42607,I42556,I37478);
nand I_2330 (I42624,I42607,I37469);
not I_2331 (I42641,I42624);
not I_2332 (I42658,I37478);
nor I_2333 (I42528,I42624,I42658);
not I_2334 (I42689,I42658);
nand I_2335 (I42513,I42624,I42689);
not I_2336 (I42720,I37481);
nor I_2337 (I42737,I42720,I37475);
and I_2338 (I42754,I42737,I37490);
or I_2339 (I42771,I42754,I37496);
DFFARX1 I_2340 (I42788,I42771,I2966,I42539,);
nor I_2341 (I42805,I42788,I42641);
DFFARX1 I_2342 (I42822,I42788,I2966,I42539,);
not I_2343 (I42510,I42822);
nand I_2344 (I42853,I42556,I37481);
and I_2345 (I42870,I42853,I42805);
DFFARX1 I_2346 (I42507,I42853,I2966,I42539,);
DFFARX1 I_2347 (I42901,I37493,I2966,I42539,);
nor I_2348 (I42918,I42901,I42624);
nand I_2349 (I42525,I42788,I42918);
nor I_2350 (I42949,I42901,I42689);
not I_2351 (I42522,I42901);
nand I_2352 (I42980,I42901,I42590);
and I_2353 (I42997,I42658,I42980);
DFFARX1 I_2354 (I42501,I42997,I2966,I42539,);
DFFARX1 I_2355 (I42504,I42901,I2966,I42539,);
DFFARX1 I_2356 (I43042,I37499,I2966,I42539,);
not I_2357 (I43059,I43042);
nand I_2358 (I43076,I43059,I42624);
and I_2359 (I43093,I42853,I43076);
DFFARX1 I_2360 (I42531,I43093,I2966,I42539,);
or I_2361 (I43124,I43059,I42870);
DFFARX1 I_2362 (I42516,I43124,I2966,I42539,);
nand I_2363 (I42519,I43059,I42949);
not I_2364 (I43202,I2973);
not I_2365 (I43219,I32523);
nor I_2366 (I43236,I32520,I32511);
nand I_2367 (I43253,I43236,I32514);
nor I_2368 (I43270,I43219,I32520);
nand I_2369 (I43287,I43270,I32508);
not I_2370 (I43304,I43287);
not I_2371 (I43321,I32520);
nor I_2372 (I43191,I43287,I43321);
not I_2373 (I43352,I43321);
nand I_2374 (I43176,I43287,I43352);
not I_2375 (I43383,I32529);
nor I_2376 (I43400,I43383,I32532);
and I_2377 (I43417,I43400,I32517);
or I_2378 (I43434,I43417,I32505);
DFFARX1 I_2379 (I43451,I43434,I2966,I43202,);
nor I_2380 (I43468,I43451,I43304);
DFFARX1 I_2381 (I43485,I43451,I2966,I43202,);
not I_2382 (I43173,I43485);
nand I_2383 (I43516,I43219,I32529);
and I_2384 (I43533,I43516,I43468);
DFFARX1 I_2385 (I43170,I43516,I2966,I43202,);
DFFARX1 I_2386 (I43564,I32526,I2966,I43202,);
nor I_2387 (I43581,I43564,I43287);
nand I_2388 (I43188,I43451,I43581);
nor I_2389 (I43612,I43564,I43352);
not I_2390 (I43185,I43564);
nand I_2391 (I43643,I43564,I43253);
and I_2392 (I43660,I43321,I43643);
DFFARX1 I_2393 (I43164,I43660,I2966,I43202,);
DFFARX1 I_2394 (I43167,I43564,I2966,I43202,);
DFFARX1 I_2395 (I43705,I32535,I2966,I43202,);
not I_2396 (I43722,I43705);
nand I_2397 (I43739,I43722,I43287);
and I_2398 (I43756,I43516,I43739);
DFFARX1 I_2399 (I43194,I43756,I2966,I43202,);
or I_2400 (I43787,I43722,I43533);
DFFARX1 I_2401 (I43179,I43787,I2966,I43202,);
nand I_2402 (I43182,I43722,I43612);
not I_2403 (I43865,I2973);
not I_2404 (I43882,I25465);
nor I_2405 (I43899,I25477,I25459);
nand I_2406 (I43916,I43899,I25480);
nor I_2407 (I43933,I43882,I25477);
nand I_2408 (I43950,I43933,I25471);
not I_2409 (I43967,I43950);
not I_2410 (I43984,I25477);
nor I_2411 (I43854,I43950,I43984);
not I_2412 (I44015,I43984);
nand I_2413 (I43839,I43950,I44015);
not I_2414 (I44046,I25462);
nor I_2415 (I44063,I44046,I25456);
and I_2416 (I44080,I44063,I25468);
or I_2417 (I44097,I44080,I25453);
DFFARX1 I_2418 (I44114,I44097,I2966,I43865,);
nor I_2419 (I44131,I44114,I43967);
DFFARX1 I_2420 (I44148,I44114,I2966,I43865,);
not I_2421 (I43836,I44148);
nand I_2422 (I44179,I43882,I25462);
and I_2423 (I44196,I44179,I44131);
DFFARX1 I_2424 (I43833,I44179,I2966,I43865,);
DFFARX1 I_2425 (I44227,I25450,I2966,I43865,);
nor I_2426 (I44244,I44227,I43950);
nand I_2427 (I43851,I44114,I44244);
nor I_2428 (I44275,I44227,I44015);
not I_2429 (I43848,I44227);
nand I_2430 (I44306,I44227,I43916);
and I_2431 (I44323,I43984,I44306);
DFFARX1 I_2432 (I43827,I44323,I2966,I43865,);
DFFARX1 I_2433 (I43830,I44227,I2966,I43865,);
DFFARX1 I_2434 (I44368,I25474,I2966,I43865,);
not I_2435 (I44385,I44368);
nand I_2436 (I44402,I44385,I43950);
and I_2437 (I44419,I44179,I44402);
DFFARX1 I_2438 (I43857,I44419,I2966,I43865,);
or I_2439 (I44450,I44385,I44196);
DFFARX1 I_2440 (I43842,I44450,I2966,I43865,);
nand I_2441 (I43845,I44385,I44275);
not I_2442 (I44528,I2973);
not I_2443 (I44545,I28955);
nor I_2444 (I44562,I28976,I28982);
nand I_2445 (I44579,I44562,I28970);
nor I_2446 (I44596,I44545,I28976);
nand I_2447 (I44613,I44596,I28952);
not I_2448 (I44630,I44613);
not I_2449 (I44647,I28976);
nor I_2450 (I44517,I44613,I44647);
not I_2451 (I44678,I44647);
nand I_2452 (I44502,I44613,I44678);
not I_2453 (I44709,I28958);
nor I_2454 (I44726,I44709,I28979);
and I_2455 (I44743,I44726,I28967);
or I_2456 (I44760,I44743,I28973);
DFFARX1 I_2457 (I44777,I44760,I2966,I44528,);
nor I_2458 (I44794,I44777,I44630);
DFFARX1 I_2459 (I44811,I44777,I2966,I44528,);
not I_2460 (I44499,I44811);
nand I_2461 (I44842,I44545,I28958);
and I_2462 (I44859,I44842,I44794);
DFFARX1 I_2463 (I44496,I44842,I2966,I44528,);
DFFARX1 I_2464 (I44890,I28964,I2966,I44528,);
nor I_2465 (I44907,I44890,I44613);
nand I_2466 (I44514,I44777,I44907);
nor I_2467 (I44938,I44890,I44678);
not I_2468 (I44511,I44890);
nand I_2469 (I44969,I44890,I44579);
and I_2470 (I44986,I44647,I44969);
DFFARX1 I_2471 (I44490,I44986,I2966,I44528,);
DFFARX1 I_2472 (I44493,I44890,I2966,I44528,);
DFFARX1 I_2473 (I45031,I28961,I2966,I44528,);
not I_2474 (I45048,I45031);
nand I_2475 (I45065,I45048,I44613);
and I_2476 (I45082,I44842,I45065);
DFFARX1 I_2477 (I44520,I45082,I2966,I44528,);
or I_2478 (I45113,I45048,I44859);
DFFARX1 I_2479 (I44505,I45113,I2966,I44528,);
nand I_2480 (I44508,I45048,I44938);
not I_2481 (I45191,I2973);
not I_2482 (I45208,I33106);
nor I_2483 (I45225,I33124,I33115);
nand I_2484 (I45242,I45225,I33121);
nor I_2485 (I45259,I45208,I33124);
nand I_2486 (I45276,I45259,I33127);
not I_2487 (I45293,I45276);
not I_2488 (I45310,I33124);
nor I_2489 (I45180,I45276,I45310);
not I_2490 (I45341,I45310);
nand I_2491 (I45165,I45276,I45341);
not I_2492 (I45372,I33103);
nor I_2493 (I45389,I45372,I33118);
and I_2494 (I45406,I45389,I33100);
or I_2495 (I45423,I45406,I33109);
DFFARX1 I_2496 (I45440,I45423,I2966,I45191,);
nor I_2497 (I45457,I45440,I45293);
DFFARX1 I_2498 (I45474,I45440,I2966,I45191,);
not I_2499 (I45162,I45474);
nand I_2500 (I45505,I45208,I33103);
and I_2501 (I45522,I45505,I45457);
DFFARX1 I_2502 (I45159,I45505,I2966,I45191,);
DFFARX1 I_2503 (I45553,I33112,I2966,I45191,);
nor I_2504 (I45570,I45553,I45276);
nand I_2505 (I45177,I45440,I45570);
nor I_2506 (I45601,I45553,I45341);
not I_2507 (I45174,I45553);
nand I_2508 (I45632,I45553,I45242);
and I_2509 (I45649,I45310,I45632);
DFFARX1 I_2510 (I45153,I45649,I2966,I45191,);
DFFARX1 I_2511 (I45156,I45553,I2966,I45191,);
DFFARX1 I_2512 (I45694,I33130,I2966,I45191,);
not I_2513 (I45711,I45694);
nand I_2514 (I45728,I45711,I45276);
and I_2515 (I45745,I45505,I45728);
DFFARX1 I_2516 (I45183,I45745,I2966,I45191,);
or I_2517 (I45776,I45711,I45522);
DFFARX1 I_2518 (I45168,I45776,I2966,I45191,);
nand I_2519 (I45171,I45711,I45601);
not I_2520 (I45854,I2973);
not I_2521 (I45871,I43851);
nor I_2522 (I45888,I43830,I43842);
nand I_2523 (I45905,I45888,I43845);
nor I_2524 (I45922,I45871,I43830);
nand I_2525 (I45939,I45922,I43827);
DFFARX1 I_2526 (I45956,I45939,I2966,I45854,);
not I_2527 (I45825,I45956);
not I_2528 (I45987,I43830);
not I_2529 (I46004,I45987);
not I_2530 (I46021,I43848);
nor I_2531 (I46038,I46021,I43839);
and I_2532 (I46055,I46038,I43833);
or I_2533 (I46072,I46055,I43857);
DFFARX1 I_2534 (I46089,I46072,I2966,I45854,);
DFFARX1 I_2535 (I45822,I46089,I2966,I45854,);
DFFARX1 I_2536 (I46120,I46089,I2966,I45854,);
DFFARX1 I_2537 (I45816,I46089,I2966,I45854,);
nand I_2538 (I46151,I45871,I43848);
nand I_2539 (I46168,I46151,I45905);
and I_2540 (I46185,I45987,I46168);
DFFARX1 I_2541 (I45846,I46185,I2966,I45854,);
and I_2542 (I45819,I46151,I46120);
DFFARX1 I_2543 (I46230,I43854,I2966,I45854,);
nor I_2544 (I45843,I46230,I46151);
nor I_2545 (I46261,I46230,I45905);
nand I_2546 (I45840,I45939,I46261);
not I_2547 (I45837,I46230);
DFFARX1 I_2548 (I46306,I43836,I2966,I45854,);
not I_2549 (I46323,I46306);
nor I_2550 (I46340,I46323,I46004);
and I_2551 (I46357,I46230,I46340);
or I_2552 (I46374,I46151,I46357);
DFFARX1 I_2553 (I45831,I46374,I2966,I45854,);
not I_2554 (I46405,I46323);
nor I_2555 (I46422,I46230,I46405);
nand I_2556 (I45834,I46323,I46422);
nand I_2557 (I45828,I45987,I46405);
not I_2558 (I46500,I2973);
not I_2559 (I46517,I31324);
nor I_2560 (I46534,I31336,I31330);
nand I_2561 (I46551,I46534,I31315);
nor I_2562 (I46568,I46517,I31336);
nand I_2563 (I46585,I46568,I31342);
DFFARX1 I_2564 (I46602,I46585,I2966,I46500,);
not I_2565 (I46471,I46602);
not I_2566 (I46633,I31336);
not I_2567 (I46650,I46633);
not I_2568 (I46667,I31339);
nor I_2569 (I46684,I46667,I31321);
and I_2570 (I46701,I46684,I31318);
or I_2571 (I46718,I46701,I31345);
DFFARX1 I_2572 (I46735,I46718,I2966,I46500,);
DFFARX1 I_2573 (I46468,I46735,I2966,I46500,);
DFFARX1 I_2574 (I46766,I46735,I2966,I46500,);
DFFARX1 I_2575 (I46462,I46735,I2966,I46500,);
nand I_2576 (I46797,I46517,I31339);
nand I_2577 (I46814,I46797,I46551);
and I_2578 (I46831,I46633,I46814);
DFFARX1 I_2579 (I46492,I46831,I2966,I46500,);
and I_2580 (I46465,I46797,I46766);
DFFARX1 I_2581 (I46876,I31333,I2966,I46500,);
nor I_2582 (I46489,I46876,I46797);
nor I_2583 (I46907,I46876,I46551);
nand I_2584 (I46486,I46585,I46907);
not I_2585 (I46483,I46876);
DFFARX1 I_2586 (I46952,I31327,I2966,I46500,);
not I_2587 (I46969,I46952);
nor I_2588 (I46986,I46969,I46650);
and I_2589 (I47003,I46876,I46986);
or I_2590 (I47020,I46797,I47003);
DFFARX1 I_2591 (I46477,I47020,I2966,I46500,);
not I_2592 (I47051,I46969);
nor I_2593 (I47068,I46876,I47051);
nand I_2594 (I46480,I46969,I47068);
nand I_2595 (I46474,I46633,I47051);
not I_2596 (I47146,I2973);
not I_2597 (I47163,I39405);
nor I_2598 (I47180,I39393,I39396);
nand I_2599 (I47197,I47180,I39420);
nor I_2600 (I47214,I47163,I39393);
nand I_2601 (I47231,I47214,I39402);
DFFARX1 I_2602 (I47248,I47231,I2966,I47146,);
not I_2603 (I47117,I47248);
not I_2604 (I47279,I39393);
not I_2605 (I47296,I47279);
not I_2606 (I47313,I39399);
nor I_2607 (I47330,I47313,I39414);
and I_2608 (I47347,I47330,I39390);
or I_2609 (I47364,I47347,I39417);
DFFARX1 I_2610 (I47381,I47364,I2966,I47146,);
DFFARX1 I_2611 (I47114,I47381,I2966,I47146,);
DFFARX1 I_2612 (I47412,I47381,I2966,I47146,);
DFFARX1 I_2613 (I47108,I47381,I2966,I47146,);
nand I_2614 (I47443,I47163,I39399);
nand I_2615 (I47460,I47443,I47197);
and I_2616 (I47477,I47279,I47460);
DFFARX1 I_2617 (I47138,I47477,I2966,I47146,);
and I_2618 (I47111,I47443,I47412);
DFFARX1 I_2619 (I47522,I39408,I2966,I47146,);
nor I_2620 (I47135,I47522,I47443);
nor I_2621 (I47553,I47522,I47197);
nand I_2622 (I47132,I47231,I47553);
not I_2623 (I47129,I47522);
DFFARX1 I_2624 (I47598,I39411,I2966,I47146,);
not I_2625 (I47615,I47598);
nor I_2626 (I47632,I47615,I47296);
and I_2627 (I47649,I47522,I47632);
or I_2628 (I47666,I47443,I47649);
DFFARX1 I_2629 (I47123,I47666,I2966,I47146,);
not I_2630 (I47697,I47615);
nor I_2631 (I47714,I47522,I47697);
nand I_2632 (I47126,I47615,I47714);
nand I_2633 (I47120,I47279,I47697);
not I_2634 (I47792,I2973);
not I_2635 (I47809,I24887);
nor I_2636 (I47826,I24890,I24872);
nand I_2637 (I47843,I47826,I24899);
nor I_2638 (I47860,I47809,I24890);
nand I_2639 (I47877,I47860,I24878);
DFFARX1 I_2640 (I47894,I47877,I2966,I47792,);
not I_2641 (I47763,I47894);
not I_2642 (I47925,I24890);
not I_2643 (I47942,I47925);
not I_2644 (I47959,I24884);
nor I_2645 (I47976,I47959,I24896);
and I_2646 (I47993,I47976,I24902);
or I_2647 (I48010,I47993,I24881);
DFFARX1 I_2648 (I48027,I48010,I2966,I47792,);
DFFARX1 I_2649 (I47760,I48027,I2966,I47792,);
DFFARX1 I_2650 (I48058,I48027,I2966,I47792,);
DFFARX1 I_2651 (I47754,I48027,I2966,I47792,);
nand I_2652 (I48089,I47809,I24884);
nand I_2653 (I48106,I48089,I47843);
and I_2654 (I48123,I47925,I48106);
DFFARX1 I_2655 (I47784,I48123,I2966,I47792,);
and I_2656 (I47757,I48089,I48058);
DFFARX1 I_2657 (I48168,I24893,I2966,I47792,);
nor I_2658 (I47781,I48168,I48089);
nor I_2659 (I48199,I48168,I47843);
nand I_2660 (I47778,I47877,I48199);
not I_2661 (I47775,I48168);
DFFARX1 I_2662 (I48244,I24875,I2966,I47792,);
not I_2663 (I48261,I48244);
nor I_2664 (I48278,I48261,I47942);
and I_2665 (I48295,I48168,I48278);
or I_2666 (I48312,I48089,I48295);
DFFARX1 I_2667 (I47769,I48312,I2966,I47792,);
not I_2668 (I48343,I48261);
nor I_2669 (I48360,I48168,I48343);
nand I_2670 (I47772,I48261,I48360);
nand I_2671 (I47766,I47925,I48343);
not I_2672 (I48438,I2973);
not I_2673 (I48455,I27199);
nor I_2674 (I48472,I27202,I27184);
nand I_2675 (I48489,I48472,I27211);
nor I_2676 (I48506,I48455,I27202);
nand I_2677 (I48523,I48506,I27190);
DFFARX1 I_2678 (I48540,I48523,I2966,I48438,);
not I_2679 (I48409,I48540);
not I_2680 (I48571,I27202);
not I_2681 (I48588,I48571);
not I_2682 (I48605,I27196);
nor I_2683 (I48622,I48605,I27208);
and I_2684 (I48639,I48622,I27214);
or I_2685 (I48656,I48639,I27193);
DFFARX1 I_2686 (I48673,I48656,I2966,I48438,);
DFFARX1 I_2687 (I48406,I48673,I2966,I48438,);
DFFARX1 I_2688 (I48704,I48673,I2966,I48438,);
DFFARX1 I_2689 (I48400,I48673,I2966,I48438,);
nand I_2690 (I48735,I48455,I27196);
nand I_2691 (I48752,I48735,I48489);
and I_2692 (I48769,I48571,I48752);
DFFARX1 I_2693 (I48430,I48769,I2966,I48438,);
and I_2694 (I48403,I48735,I48704);
DFFARX1 I_2695 (I48814,I27205,I2966,I48438,);
nor I_2696 (I48427,I48814,I48735);
nor I_2697 (I48845,I48814,I48489);
nand I_2698 (I48424,I48523,I48845);
not I_2699 (I48421,I48814);
DFFARX1 I_2700 (I48890,I27187,I2966,I48438,);
not I_2701 (I48907,I48890);
nor I_2702 (I48924,I48907,I48588);
and I_2703 (I48941,I48814,I48924);
or I_2704 (I48958,I48735,I48941);
DFFARX1 I_2705 (I48415,I48958,I2966,I48438,);
not I_2706 (I48989,I48907);
nor I_2707 (I49006,I48814,I48989);
nand I_2708 (I48418,I48907,I49006);
nand I_2709 (I48412,I48571,I48989);
not I_2710 (I49084,I2973);
or I_2711 (I49101,I44502,I44490);
or I_2712 (I49118,I44499,I44502);
nor I_2713 (I49135,I44493,I44514);
DFFARX1 I_2714 (I49152,I49135,I2966,I49084,);
DFFARX1 I_2715 (I49046,I49135,I2966,I49084,);
not I_2716 (I49183,I44493);
and I_2717 (I49200,I49183,I44508);
nor I_2718 (I49217,I49200,I44490);
nor I_2719 (I49234,I44505,I44520);
DFFARX1 I_2720 (I49251,I49234,I2966,I49084,);
not I_2721 (I49268,I49251);
DFFARX1 I_2722 (I49055,I49251,I2966,I49084,);
nor I_2723 (I49299,I44505,I44499);
and I_2724 (I49049,I49299,I49152);
DFFARX1 I_2725 (I49330,I44517,I2966,I49084,);
and I_2726 (I49347,I49330,I44496);
nand I_2727 (I49364,I49347,I49118);
and I_2728 (I49381,I49251,I49364);
DFFARX1 I_2729 (I49076,I49381,I2966,I49084,);
nor I_2730 (I49073,I49347,I49217);
not I_2731 (I49426,I49347);
nor I_2732 (I49443,I49101,I49426);
nor I_2733 (I49460,I49347,I49299);
nand I_2734 (I49070,I49118,I49460);
nor I_2735 (I49491,I49347,I49268);
not I_2736 (I49067,I49347);
nand I_2737 (I49058,I49347,I49268);
DFFARX1 I_2738 (I49536,I44511,I2966,I49084,);
and I_2739 (I49553,I49536,I49443);
or I_2740 (I49570,I49101,I49553);
DFFARX1 I_2741 (I49061,I49570,I2966,I49084,);
nand I_2742 (I49064,I49536,I49491);
nand I_2743 (I49615,I49536,I49217);
and I_2744 (I49632,I49135,I49615);
DFFARX1 I_2745 (I49052,I49632,I2966,I49084,);
not I_2746 (I49696,I2973);
or I_2747 (I49713,I40601,I40610);
or I_2748 (I49730,I40595,I40601);
nor I_2749 (I49747,I40589,I40583);
DFFARX1 I_2750 (I49764,I49747,I2966,I49696,);
DFFARX1 I_2751 (I49658,I49747,I2966,I49696,);
not I_2752 (I49795,I40589);
and I_2753 (I49812,I49795,I40580);
nor I_2754 (I49829,I49812,I40610);
nor I_2755 (I49846,I40607,I40604);
DFFARX1 I_2756 (I49863,I49846,I2966,I49696,);
not I_2757 (I49880,I49863);
DFFARX1 I_2758 (I49667,I49863,I2966,I49696,);
nor I_2759 (I49911,I40607,I40595);
and I_2760 (I49661,I49911,I49764);
DFFARX1 I_2761 (I49942,I40586,I2966,I49696,);
and I_2762 (I49959,I49942,I40592);
nand I_2763 (I49976,I49959,I49730);
and I_2764 (I49993,I49863,I49976);
DFFARX1 I_2765 (I49688,I49993,I2966,I49696,);
nor I_2766 (I49685,I49959,I49829);
not I_2767 (I50038,I49959);
nor I_2768 (I50055,I49713,I50038);
nor I_2769 (I50072,I49959,I49911);
nand I_2770 (I49682,I49730,I50072);
nor I_2771 (I50103,I49959,I49880);
not I_2772 (I49679,I49959);
nand I_2773 (I49670,I49959,I49880);
DFFARX1 I_2774 (I50148,I40598,I2966,I49696,);
and I_2775 (I50165,I50148,I50055);
or I_2776 (I50182,I49713,I50165);
DFFARX1 I_2777 (I49673,I50182,I2966,I49696,);
nand I_2778 (I49676,I50148,I50103);
nand I_2779 (I50227,I50148,I49829);
and I_2780 (I50244,I49747,I50227);
DFFARX1 I_2781 (I49664,I50244,I2966,I49696,);
not I_2782 (I50308,I2973);
nand I_2783 (I50325,I39985,I39988);
and I_2784 (I50342,I50325,I39994);
DFFARX1 I_2785 (I50359,I50342,I2966,I50308,);
not I_2786 (I50376,I50359);
DFFARX1 I_2787 (I50276,I50359,I2966,I50308,);
nor I_2788 (I50407,I40006,I39988);
DFFARX1 I_2789 (I50424,I39997,I2966,I50308,);
DFFARX1 I_2790 (I50441,I50424,I2966,I50308,);
not I_2791 (I50279,I50441);
DFFARX1 I_2792 (I50472,I50424,I2966,I50308,);
and I_2793 (I50273,I50359,I50472);
nand I_2794 (I50503,I40003,I40000);
and I_2795 (I50520,I50503,I40012);
DFFARX1 I_2796 (I50537,I50520,I2966,I50308,);
nor I_2797 (I50554,I50537,I50376);
not I_2798 (I50571,I50537);
nand I_2799 (I50282,I50359,I50571);
DFFARX1 I_2800 (I50602,I40009,I2966,I50308,);
and I_2801 (I50619,I50602,I40015);
nor I_2802 (I50636,I50619,I50537);
nor I_2803 (I50653,I50619,I50571);
nand I_2804 (I50288,I50407,I50653);
not I_2805 (I50291,I50619);
DFFARX1 I_2806 (I50270,I50619,I2966,I50308,);
DFFARX1 I_2807 (I50712,I39991,I2966,I50308,);
nand I_2808 (I50729,I50712,I50424);
and I_2809 (I50746,I50407,I50729);
DFFARX1 I_2810 (I50300,I50746,I2966,I50308,);
nor I_2811 (I50297,I50712,I50619);
and I_2812 (I50791,I50712,I50554);
or I_2813 (I50808,I50407,I50791);
DFFARX1 I_2814 (I50285,I50808,I2966,I50308,);
nand I_2815 (I50294,I50712,I50636);
not I_2816 (I50886,I2973);
nand I_2817 (I50903,I38159,I38138);
and I_2818 (I50920,I50903,I38135);
DFFARX1 I_2819 (I50937,I50920,I2966,I50886,);
not I_2820 (I50954,I50937);
DFFARX1 I_2821 (I50854,I50937,I2966,I50886,);
nor I_2822 (I50985,I38144,I38138);
DFFARX1 I_2823 (I51002,I38132,I2966,I50886,);
DFFARX1 I_2824 (I51019,I51002,I2966,I50886,);
not I_2825 (I50857,I51019);
DFFARX1 I_2826 (I51050,I51002,I2966,I50886,);
and I_2827 (I50851,I50937,I51050);
nand I_2828 (I51081,I38162,I38153);
and I_2829 (I51098,I51081,I38150);
DFFARX1 I_2830 (I51115,I51098,I2966,I50886,);
nor I_2831 (I51132,I51115,I50954);
not I_2832 (I51149,I51115);
nand I_2833 (I50860,I50937,I51149);
DFFARX1 I_2834 (I51180,I38147,I2966,I50886,);
and I_2835 (I51197,I51180,I38156);
nor I_2836 (I51214,I51197,I51115);
nor I_2837 (I51231,I51197,I51149);
nand I_2838 (I50866,I50985,I51231);
not I_2839 (I50869,I51197);
DFFARX1 I_2840 (I50848,I51197,I2966,I50886,);
DFFARX1 I_2841 (I51290,I38141,I2966,I50886,);
nand I_2842 (I51307,I51290,I51002);
and I_2843 (I51324,I50985,I51307);
DFFARX1 I_2844 (I50878,I51324,I2966,I50886,);
nor I_2845 (I50875,I51290,I51197);
and I_2846 (I51369,I51290,I51132);
or I_2847 (I51386,I50985,I51369);
DFFARX1 I_2848 (I50863,I51386,I2966,I50886,);
nand I_2849 (I50872,I51290,I51214);
not I_2850 (I51464,I2973);
nand I_2851 (I51481,I43167,I43194);
and I_2852 (I51498,I51481,I43182);
DFFARX1 I_2853 (I51515,I51498,I2966,I51464,);
not I_2854 (I51532,I51515);
DFFARX1 I_2855 (I51432,I51515,I2966,I51464,);
nor I_2856 (I51563,I43170,I43194);
DFFARX1 I_2857 (I51580,I43185,I2966,I51464,);
DFFARX1 I_2858 (I51597,I51580,I2966,I51464,);
not I_2859 (I51435,I51597);
DFFARX1 I_2860 (I51628,I51580,I2966,I51464,);
and I_2861 (I51429,I51515,I51628);
nand I_2862 (I51659,I43179,I43176);
and I_2863 (I51676,I51659,I43173);
DFFARX1 I_2864 (I51693,I51676,I2966,I51464,);
nor I_2865 (I51710,I51693,I51532);
not I_2866 (I51727,I51693);
nand I_2867 (I51438,I51515,I51727);
DFFARX1 I_2868 (I51758,I43188,I2966,I51464,);
and I_2869 (I51775,I51758,I43164);
nor I_2870 (I51792,I51775,I51693);
nor I_2871 (I51809,I51775,I51727);
nand I_2872 (I51444,I51563,I51809);
not I_2873 (I51447,I51775);
DFFARX1 I_2874 (I51426,I51775,I2966,I51464,);
DFFARX1 I_2875 (I51868,I43191,I2966,I51464,);
nand I_2876 (I51885,I51868,I51580);
and I_2877 (I51902,I51563,I51885);
DFFARX1 I_2878 (I51456,I51902,I2966,I51464,);
nor I_2879 (I51453,I51868,I51775);
and I_2880 (I51947,I51868,I51710);
or I_2881 (I51964,I51563,I51947);
DFFARX1 I_2882 (I51441,I51964,I2966,I51464,);
nand I_2883 (I51450,I51868,I51792);
not I_2884 (I52042,I2973);
nand I_2885 (I52059,I45831,I45828);
and I_2886 (I52076,I52059,I45840);
DFFARX1 I_2887 (I52093,I52076,I2966,I52042,);
not I_2888 (I52110,I52093);
DFFARX1 I_2889 (I52010,I52093,I2966,I52042,);
nor I_2890 (I52141,I45837,I45828);
DFFARX1 I_2891 (I52158,I45843,I2966,I52042,);
DFFARX1 I_2892 (I52175,I52158,I2966,I52042,);
not I_2893 (I52013,I52175);
DFFARX1 I_2894 (I52206,I52158,I2966,I52042,);
and I_2895 (I52007,I52093,I52206);
nand I_2896 (I52237,I45819,I45822);
and I_2897 (I52254,I52237,I45846);
DFFARX1 I_2898 (I52271,I52254,I2966,I52042,);
nor I_2899 (I52288,I52271,I52110);
not I_2900 (I52305,I52271);
nand I_2901 (I52016,I52093,I52305);
DFFARX1 I_2902 (I52336,I45825,I2966,I52042,);
and I_2903 (I52353,I52336,I45816);
nor I_2904 (I52370,I52353,I52271);
nor I_2905 (I52387,I52353,I52305);
nand I_2906 (I52022,I52141,I52387);
not I_2907 (I52025,I52353);
DFFARX1 I_2908 (I52004,I52353,I2966,I52042,);
DFFARX1 I_2909 (I52446,I45834,I2966,I52042,);
nand I_2910 (I52463,I52446,I52158);
and I_2911 (I52480,I52141,I52463);
DFFARX1 I_2912 (I52034,I52480,I2966,I52042,);
nor I_2913 (I52031,I52446,I52353);
and I_2914 (I52525,I52446,I52288);
or I_2915 (I52542,I52141,I52525);
DFFARX1 I_2916 (I52019,I52542,I2966,I52042,);
nand I_2917 (I52028,I52446,I52370);
not I_2918 (I52620,I2973);
nand I_2919 (I52637,I34376,I34379);
and I_2920 (I52654,I52637,I34385);
DFFARX1 I_2921 (I52671,I52654,I2966,I52620,);
not I_2922 (I52688,I52671);
DFFARX1 I_2923 (I52588,I52671,I2966,I52620,);
nor I_2924 (I52719,I34382,I34379);
DFFARX1 I_2925 (I52736,I34361,I2966,I52620,);
DFFARX1 I_2926 (I52753,I52736,I2966,I52620,);
not I_2927 (I52591,I52753);
DFFARX1 I_2928 (I52784,I52736,I2966,I52620,);
and I_2929 (I52585,I52671,I52784);
nand I_2930 (I52815,I34358,I34373);
and I_2931 (I52832,I52815,I34370);
DFFARX1 I_2932 (I52849,I52832,I2966,I52620,);
nor I_2933 (I52866,I52849,I52688);
not I_2934 (I52883,I52849);
nand I_2935 (I52594,I52671,I52883);
DFFARX1 I_2936 (I52914,I34388,I2966,I52620,);
and I_2937 (I52931,I52914,I34367);
nor I_2938 (I52948,I52931,I52849);
nor I_2939 (I52965,I52931,I52883);
nand I_2940 (I52600,I52719,I52965);
not I_2941 (I52603,I52931);
DFFARX1 I_2942 (I52582,I52931,I2966,I52620,);
DFFARX1 I_2943 (I53024,I34364,I2966,I52620,);
nand I_2944 (I53041,I53024,I52736);
and I_2945 (I53058,I52719,I53041);
DFFARX1 I_2946 (I52612,I53058,I2966,I52620,);
nor I_2947 (I52609,I53024,I52931);
and I_2948 (I53103,I53024,I52866);
or I_2949 (I53120,I52719,I53103);
DFFARX1 I_2950 (I52597,I53120,I2966,I52620,);
nand I_2951 (I52606,I53024,I52948);
not I_2952 (I53198,I2973);
nand I_2953 (I53215,I47123,I47120);
and I_2954 (I53232,I53215,I47132);
DFFARX1 I_2955 (I53249,I53232,I2966,I53198,);
not I_2956 (I53266,I53249);
DFFARX1 I_2957 (I53166,I53249,I2966,I53198,);
nor I_2958 (I53297,I47129,I47120);
DFFARX1 I_2959 (I53314,I47135,I2966,I53198,);
DFFARX1 I_2960 (I53331,I53314,I2966,I53198,);
not I_2961 (I53169,I53331);
DFFARX1 I_2962 (I53362,I53314,I2966,I53198,);
and I_2963 (I53163,I53249,I53362);
nand I_2964 (I53393,I47111,I47114);
and I_2965 (I53410,I53393,I47138);
DFFARX1 I_2966 (I53427,I53410,I2966,I53198,);
nor I_2967 (I53444,I53427,I53266);
not I_2968 (I53461,I53427);
nand I_2969 (I53172,I53249,I53461);
DFFARX1 I_2970 (I53492,I47117,I2966,I53198,);
and I_2971 (I53509,I53492,I47108);
nor I_2972 (I53526,I53509,I53427);
nor I_2973 (I53543,I53509,I53461);
nand I_2974 (I53178,I53297,I53543);
not I_2975 (I53181,I53509);
DFFARX1 I_2976 (I53160,I53509,I2966,I53198,);
DFFARX1 I_2977 (I53602,I47126,I2966,I53198,);
nand I_2978 (I53619,I53602,I53314);
and I_2979 (I53636,I53297,I53619);
DFFARX1 I_2980 (I53190,I53636,I2966,I53198,);
nor I_2981 (I53187,I53602,I53509);
and I_2982 (I53681,I53602,I53444);
or I_2983 (I53698,I53297,I53681);
DFFARX1 I_2984 (I53175,I53698,I2966,I53198,);
nand I_2985 (I53184,I53602,I53526);
not I_2986 (I53776,I2973);
nand I_2987 (I53793,I35634,I35625);
and I_2988 (I53810,I53793,I35643);
DFFARX1 I_2989 (I53827,I53810,I2966,I53776,);
nor I_2990 (I53844,I35640,I35625);
nor I_2991 (I53861,I53844,I53827);
not I_2992 (I53759,I53844);
DFFARX1 I_2993 (I53892,I35622,I2966,I53776,);
not I_2994 (I53909,I53892);
nor I_2995 (I53926,I53844,I53909);
nand I_2996 (I53762,I53892,I53861);
DFFARX1 I_2997 (I53744,I53892,I2966,I53776,);
nand I_2998 (I53971,I35631,I35646);
and I_2999 (I53988,I53971,I35637);
DFFARX1 I_3000 (I54005,I53988,I2966,I53776,);
nor I_3001 (I53765,I54005,I53827);
nand I_3002 (I53756,I54005,I53926);
DFFARX1 I_3003 (I54050,I35619,I2966,I53776,);
and I_3004 (I54067,I54050,I35628);
DFFARX1 I_3005 (I54084,I54067,I2966,I53776,);
not I_3006 (I53747,I54084);
nand I_3007 (I54115,I54067,I54005);
and I_3008 (I54132,I53827,I54115);
DFFARX1 I_3009 (I53738,I54132,I2966,I53776,);
DFFARX1 I_3010 (I54163,I35616,I2966,I53776,);
nand I_3011 (I54180,I54163,I53827);
and I_3012 (I54197,I54005,I54180);
DFFARX1 I_3013 (I53768,I54197,I2966,I53776,);
not I_3014 (I54228,I54163);
nor I_3015 (I54245,I53844,I54228);
and I_3016 (I54262,I54163,I54245);
or I_3017 (I54279,I54067,I54262);
DFFARX1 I_3018 (I53753,I54279,I2966,I53776,);
nand I_3019 (I53750,I54163,I53909);
DFFARX1 I_3020 (I53741,I54163,I2966,I53776,);
not I_3021 (I54371,I2973);
nand I_3022 (I54388,I33747,I33738);
and I_3023 (I54405,I54388,I33756);
DFFARX1 I_3024 (I54422,I54405,I2966,I54371,);
nor I_3025 (I54439,I33753,I33738);
nor I_3026 (I54456,I54439,I54422);
not I_3027 (I54354,I54439);
DFFARX1 I_3028 (I54487,I33735,I2966,I54371,);
not I_3029 (I54504,I54487);
nor I_3030 (I54521,I54439,I54504);
nand I_3031 (I54357,I54487,I54456);
DFFARX1 I_3032 (I54339,I54487,I2966,I54371,);
nand I_3033 (I54566,I33744,I33759);
and I_3034 (I54583,I54566,I33750);
DFFARX1 I_3035 (I54600,I54583,I2966,I54371,);
nor I_3036 (I54360,I54600,I54422);
nand I_3037 (I54351,I54600,I54521);
DFFARX1 I_3038 (I54645,I33732,I2966,I54371,);
and I_3039 (I54662,I54645,I33741);
DFFARX1 I_3040 (I54679,I54662,I2966,I54371,);
not I_3041 (I54342,I54679);
nand I_3042 (I54710,I54662,I54600);
and I_3043 (I54727,I54422,I54710);
DFFARX1 I_3044 (I54333,I54727,I2966,I54371,);
DFFARX1 I_3045 (I54758,I33729,I2966,I54371,);
nand I_3046 (I54775,I54758,I54422);
and I_3047 (I54792,I54600,I54775);
DFFARX1 I_3048 (I54363,I54792,I2966,I54371,);
not I_3049 (I54823,I54758);
nor I_3050 (I54840,I54439,I54823);
and I_3051 (I54857,I54758,I54840);
or I_3052 (I54874,I54662,I54857);
DFFARX1 I_3053 (I54348,I54874,I2966,I54371,);
nand I_3054 (I54345,I54758,I54504);
DFFARX1 I_3055 (I54336,I54758,I2966,I54371,);
not I_3056 (I54966,I2973);
nand I_3057 (I54983,I53187,I53190);
and I_3058 (I55000,I54983,I53184);
DFFARX1 I_3059 (I55017,I55000,I2966,I54966,);
nor I_3060 (I55034,I53181,I53190);
nor I_3061 (I55051,I55034,I55017);
not I_3062 (I54949,I55034);
DFFARX1 I_3063 (I55082,I53163,I2966,I54966,);
not I_3064 (I55099,I55082);
nor I_3065 (I55116,I55034,I55099);
nand I_3066 (I54952,I55082,I55051);
DFFARX1 I_3067 (I54934,I55082,I2966,I54966,);
nand I_3068 (I55161,I53172,I53169);
and I_3069 (I55178,I55161,I53178);
DFFARX1 I_3070 (I55195,I55178,I2966,I54966,);
nor I_3071 (I54955,I55195,I55017);
nand I_3072 (I54946,I55195,I55116);
DFFARX1 I_3073 (I55240,I53160,I2966,I54966,);
and I_3074 (I55257,I55240,I53175);
DFFARX1 I_3075 (I55274,I55257,I2966,I54966,);
not I_3076 (I54937,I55274);
nand I_3077 (I55305,I55257,I55195);
and I_3078 (I55322,I55017,I55305);
DFFARX1 I_3079 (I54928,I55322,I2966,I54966,);
DFFARX1 I_3080 (I55353,I53166,I2966,I54966,);
nand I_3081 (I55370,I55353,I55017);
and I_3082 (I55387,I55195,I55370);
DFFARX1 I_3083 (I54958,I55387,I2966,I54966,);
not I_3084 (I55418,I55353);
nor I_3085 (I55435,I55034,I55418);
and I_3086 (I55452,I55353,I55435);
or I_3087 (I55469,I55257,I55452);
DFFARX1 I_3088 (I54943,I55469,I2966,I54966,);
nand I_3089 (I54940,I55353,I55099);
DFFARX1 I_3090 (I54931,I55353,I2966,I54966,);
not I_3091 (I55561,I2973);
nand I_3092 (I55578,I35005,I34996);
and I_3093 (I55595,I55578,I35014);
DFFARX1 I_3094 (I55612,I55595,I2966,I55561,);
nor I_3095 (I55629,I35011,I34996);
nor I_3096 (I55646,I55629,I55612);
not I_3097 (I55544,I55629);
DFFARX1 I_3098 (I55677,I34993,I2966,I55561,);
not I_3099 (I55694,I55677);
nor I_3100 (I55711,I55629,I55694);
nand I_3101 (I55547,I55677,I55646);
DFFARX1 I_3102 (I55529,I55677,I2966,I55561,);
nand I_3103 (I55756,I35002,I35017);
and I_3104 (I55773,I55756,I35008);
DFFARX1 I_3105 (I55790,I55773,I2966,I55561,);
nor I_3106 (I55550,I55790,I55612);
nand I_3107 (I55541,I55790,I55711);
DFFARX1 I_3108 (I55835,I34990,I2966,I55561,);
and I_3109 (I55852,I55835,I34999);
DFFARX1 I_3110 (I55869,I55852,I2966,I55561,);
not I_3111 (I55532,I55869);
nand I_3112 (I55900,I55852,I55790);
and I_3113 (I55917,I55612,I55900);
DFFARX1 I_3114 (I55523,I55917,I2966,I55561,);
DFFARX1 I_3115 (I55948,I34987,I2966,I55561,);
nand I_3116 (I55965,I55948,I55612);
and I_3117 (I55982,I55790,I55965);
DFFARX1 I_3118 (I55553,I55982,I2966,I55561,);
not I_3119 (I56013,I55948);
nor I_3120 (I56030,I55629,I56013);
and I_3121 (I56047,I55948,I56030);
or I_3122 (I56064,I55852,I56047);
DFFARX1 I_3123 (I55538,I56064,I2966,I55561,);
nand I_3124 (I55535,I55948,I55694);
DFFARX1 I_3125 (I55526,I55948,I2966,I55561,);
not I_3126 (I56156,I2973);
nand I_3127 (I56173,I47772,I47784);
and I_3128 (I56190,I56173,I47766);
DFFARX1 I_3129 (I56207,I56190,I2966,I56156,);
nor I_3130 (I56224,I47778,I47784);
nor I_3131 (I56241,I56224,I56207);
not I_3132 (I56139,I56224);
DFFARX1 I_3133 (I56272,I47763,I2966,I56156,);
not I_3134 (I56289,I56272);
nor I_3135 (I56306,I56224,I56289);
nand I_3136 (I56142,I56272,I56241);
DFFARX1 I_3137 (I56124,I56272,I2966,I56156,);
nand I_3138 (I56351,I47754,I47769);
and I_3139 (I56368,I56351,I47760);
DFFARX1 I_3140 (I56385,I56368,I2966,I56156,);
nor I_3141 (I56145,I56385,I56207);
nand I_3142 (I56136,I56385,I56306);
DFFARX1 I_3143 (I56430,I47781,I2966,I56156,);
and I_3144 (I56447,I56430,I47775);
DFFARX1 I_3145 (I56464,I56447,I2966,I56156,);
not I_3146 (I56127,I56464);
nand I_3147 (I56495,I56447,I56385);
and I_3148 (I56512,I56207,I56495);
DFFARX1 I_3149 (I56118,I56512,I2966,I56156,);
DFFARX1 I_3150 (I56543,I47757,I2966,I56156,);
nand I_3151 (I56560,I56543,I56207);
and I_3152 (I56577,I56385,I56560);
DFFARX1 I_3153 (I56148,I56577,I2966,I56156,);
not I_3154 (I56608,I56543);
nor I_3155 (I56625,I56224,I56608);
and I_3156 (I56642,I56543,I56625);
or I_3157 (I56659,I56447,I56642);
DFFARX1 I_3158 (I56133,I56659,I2966,I56156,);
nand I_3159 (I56130,I56543,I56289);
DFFARX1 I_3160 (I56121,I56543,I2966,I56156,);
not I_3161 (I56751,I2973);
nand I_3162 (I56768,I45183,I45153);
and I_3163 (I56785,I56768,I45171);
DFFARX1 I_3164 (I56802,I56785,I2966,I56751,);
nor I_3165 (I56819,I45165,I45153);
DFFARX1 I_3166 (I56836,I45162,I2966,I56751,);
nand I_3167 (I56853,I56836,I56819);
DFFARX1 I_3168 (I56722,I56836,I2966,I56751,);
nand I_3169 (I56884,I45156,I45159);
and I_3170 (I56901,I56884,I45177);
DFFARX1 I_3171 (I56918,I56901,I2966,I56751,);
not I_3172 (I56935,I56918);
nor I_3173 (I56952,I56802,I56935);
and I_3174 (I56969,I56819,I56952);
and I_3175 (I56986,I56918,I56853);
DFFARX1 I_3176 (I56719,I56986,I2966,I56751,);
DFFARX1 I_3177 (I56713,I56918,I2966,I56751,);
DFFARX1 I_3178 (I57031,I45180,I2966,I56751,);
and I_3179 (I57048,I57031,I45174);
nand I_3180 (I57065,I57048,I56918);
nor I_3181 (I56740,I57048,I56819);
not I_3182 (I57096,I57048);
nor I_3183 (I57113,I56802,I57096);
nand I_3184 (I56731,I56836,I57113);
nand I_3185 (I56725,I56918,I57096);
or I_3186 (I57158,I57048,I56969);
DFFARX1 I_3187 (I56728,I57158,I2966,I56751,);
DFFARX1 I_3188 (I57189,I45168,I2966,I56751,);
and I_3189 (I57206,I57189,I57065);
DFFARX1 I_3190 (I56743,I57206,I2966,I56751,);
nor I_3191 (I57237,I57189,I56802);
nand I_3192 (I56737,I57048,I57237);
not I_3193 (I56734,I57189);
DFFARX1 I_3194 (I57282,I57189,I2966,I56751,);
and I_3195 (I56716,I57189,I57282);
not I_3196 (I57346,I2973);
nand I_3197 (I57363,I41868,I41838);
and I_3198 (I57380,I57363,I41856);
DFFARX1 I_3199 (I57397,I57380,I2966,I57346,);
nor I_3200 (I57414,I41850,I41838);
DFFARX1 I_3201 (I57431,I41847,I2966,I57346,);
nand I_3202 (I57448,I57431,I57414);
DFFARX1 I_3203 (I57317,I57431,I2966,I57346,);
nand I_3204 (I57479,I41841,I41844);
and I_3205 (I57496,I57479,I41862);
DFFARX1 I_3206 (I57513,I57496,I2966,I57346,);
not I_3207 (I57530,I57513);
nor I_3208 (I57547,I57397,I57530);
and I_3209 (I57564,I57414,I57547);
and I_3210 (I57581,I57513,I57448);
DFFARX1 I_3211 (I57314,I57581,I2966,I57346,);
DFFARX1 I_3212 (I57308,I57513,I2966,I57346,);
DFFARX1 I_3213 (I57626,I41865,I2966,I57346,);
and I_3214 (I57643,I57626,I41859);
nand I_3215 (I57660,I57643,I57513);
nor I_3216 (I57335,I57643,I57414);
not I_3217 (I57691,I57643);
nor I_3218 (I57708,I57397,I57691);
nand I_3219 (I57326,I57431,I57708);
nand I_3220 (I57320,I57513,I57691);
or I_3221 (I57753,I57643,I57564);
DFFARX1 I_3222 (I57323,I57753,I2966,I57346,);
DFFARX1 I_3223 (I57784,I41853,I2966,I57346,);
and I_3224 (I57801,I57784,I57660);
DFFARX1 I_3225 (I57338,I57801,I2966,I57346,);
nor I_3226 (I57832,I57784,I57397);
nand I_3227 (I57332,I57643,I57832);
not I_3228 (I57329,I57784);
DFFARX1 I_3229 (I57877,I57784,I2966,I57346,);
and I_3230 (I57311,I57784,I57877);
not I_3231 (I57941,I2973);
nand I_3232 (I57958,I54348,I54333);
and I_3233 (I57975,I57958,I54339);
DFFARX1 I_3234 (I57992,I57975,I2966,I57941,);
nor I_3235 (I58009,I54342,I54333);
DFFARX1 I_3236 (I58026,I54354,I2966,I57941,);
nand I_3237 (I58043,I58026,I58009);
DFFARX1 I_3238 (I57912,I58026,I2966,I57941,);
nand I_3239 (I58074,I54345,I54336);
and I_3240 (I58091,I58074,I54363);
DFFARX1 I_3241 (I58108,I58091,I2966,I57941,);
not I_3242 (I58125,I58108);
nor I_3243 (I58142,I57992,I58125);
and I_3244 (I58159,I58009,I58142);
and I_3245 (I58176,I58108,I58043);
DFFARX1 I_3246 (I57909,I58176,I2966,I57941,);
DFFARX1 I_3247 (I57903,I58108,I2966,I57941,);
DFFARX1 I_3248 (I58221,I54351,I2966,I57941,);
and I_3249 (I58238,I58221,I54357);
nand I_3250 (I58255,I58238,I58108);
nor I_3251 (I57930,I58238,I58009);
not I_3252 (I58286,I58238);
nor I_3253 (I58303,I57992,I58286);
nand I_3254 (I57921,I58026,I58303);
nand I_3255 (I57915,I58108,I58286);
or I_3256 (I58348,I58238,I58159);
DFFARX1 I_3257 (I57918,I58348,I2966,I57941,);
DFFARX1 I_3258 (I58379,I54360,I2966,I57941,);
and I_3259 (I58396,I58379,I58255);
DFFARX1 I_3260 (I57933,I58396,I2966,I57941,);
nor I_3261 (I58427,I58379,I57992);
nand I_3262 (I57927,I58238,I58427);
not I_3263 (I57924,I58379);
DFFARX1 I_3264 (I58472,I58379,I2966,I57941,);
and I_3265 (I57906,I58379,I58472);
not I_3266 (I58536,I2973);
not I_3267 (I58553,I54934);
nor I_3268 (I58570,I54952,I54931);
nand I_3269 (I58587,I58570,I54955);
nor I_3270 (I58604,I58553,I54952);
nand I_3271 (I58621,I58604,I54949);
not I_3272 (I58638,I54952);
not I_3273 (I58655,I58638);
not I_3274 (I58672,I54940);
nor I_3275 (I58689,I58672,I54928);
and I_3276 (I58706,I58689,I54946);
or I_3277 (I58723,I58706,I54958);
DFFARX1 I_3278 (I58740,I58723,I2966,I58536,);
nand I_3279 (I58757,I58553,I54940);
or I_3280 (I58525,I58757,I58740);
not I_3281 (I58788,I58757);
nor I_3282 (I58805,I58740,I58788);
and I_3283 (I58822,I58638,I58805);
nand I_3284 (I58498,I58757,I58655);
DFFARX1 I_3285 (I58853,I54937,I2966,I58536,);
or I_3286 (I58519,I58853,I58740);
nor I_3287 (I58884,I58853,I58621);
nor I_3288 (I58901,I58853,I58655);
nand I_3289 (I58504,I58587,I58901);
or I_3290 (I58932,I58853,I58822);
DFFARX1 I_3291 (I58501,I58932,I2966,I58536,);
not I_3292 (I58507,I58853);
DFFARX1 I_3293 (I58977,I54943,I2966,I58536,);
not I_3294 (I58994,I58977);
nor I_3295 (I59011,I58994,I58587);
DFFARX1 I_3296 (I58513,I59011,I2966,I58536,);
nor I_3297 (I58528,I58853,I58994);
nor I_3298 (I58516,I58994,I58757);
not I_3299 (I59070,I58994);
and I_3300 (I59087,I58621,I59070);
nor I_3301 (I58522,I58757,I59087);
nand I_3302 (I58510,I58994,I58884);
not I_3303 (I59165,I2973);
not I_3304 (I59182,I55529);
nor I_3305 (I59199,I55547,I55526);
nand I_3306 (I59216,I59199,I55550);
nor I_3307 (I59233,I59182,I55547);
nand I_3308 (I59250,I59233,I55544);
not I_3309 (I59267,I55547);
not I_3310 (I59284,I59267);
not I_3311 (I59301,I55535);
nor I_3312 (I59318,I59301,I55523);
and I_3313 (I59335,I59318,I55541);
or I_3314 (I59352,I59335,I55553);
DFFARX1 I_3315 (I59369,I59352,I2966,I59165,);
nand I_3316 (I59386,I59182,I55535);
or I_3317 (I59154,I59386,I59369);
not I_3318 (I59417,I59386);
nor I_3319 (I59434,I59369,I59417);
and I_3320 (I59451,I59267,I59434);
nand I_3321 (I59127,I59386,I59284);
DFFARX1 I_3322 (I59482,I55532,I2966,I59165,);
or I_3323 (I59148,I59482,I59369);
nor I_3324 (I59513,I59482,I59250);
nor I_3325 (I59530,I59482,I59284);
nand I_3326 (I59133,I59216,I59530);
or I_3327 (I59561,I59482,I59451);
DFFARX1 I_3328 (I59130,I59561,I2966,I59165,);
not I_3329 (I59136,I59482);
DFFARX1 I_3330 (I59606,I55538,I2966,I59165,);
not I_3331 (I59623,I59606);
nor I_3332 (I59640,I59623,I59216);
DFFARX1 I_3333 (I59142,I59640,I2966,I59165,);
nor I_3334 (I59157,I59482,I59623);
nor I_3335 (I59145,I59623,I59386);
not I_3336 (I59699,I59623);
and I_3337 (I59716,I59250,I59699);
nor I_3338 (I59151,I59386,I59716);
nand I_3339 (I59139,I59623,I59513);
not I_3340 (I59794,I2973);
not I_3341 (I59811,I42519);
nor I_3342 (I59828,I42525,I42504);
nand I_3343 (I59845,I59828,I42510);
nor I_3344 (I59862,I59811,I42525);
nand I_3345 (I59879,I59862,I42516);
not I_3346 (I59896,I42525);
not I_3347 (I59913,I59896);
not I_3348 (I59930,I42513);
nor I_3349 (I59947,I59930,I42531);
and I_3350 (I59964,I59947,I42522);
or I_3351 (I59981,I59964,I42501);
DFFARX1 I_3352 (I59998,I59981,I2966,I59794,);
nand I_3353 (I60015,I59811,I42513);
or I_3354 (I59783,I60015,I59998);
not I_3355 (I60046,I60015);
nor I_3356 (I60063,I59998,I60046);
and I_3357 (I60080,I59896,I60063);
nand I_3358 (I59756,I60015,I59913);
DFFARX1 I_3359 (I60111,I42528,I2966,I59794,);
or I_3360 (I59777,I60111,I59998);
nor I_3361 (I60142,I60111,I59879);
nor I_3362 (I60159,I60111,I59913);
nand I_3363 (I59762,I59845,I60159);
or I_3364 (I60190,I60111,I60080);
DFFARX1 I_3365 (I59759,I60190,I2966,I59794,);
not I_3366 (I59765,I60111);
DFFARX1 I_3367 (I60235,I42507,I2966,I59794,);
not I_3368 (I60252,I60235);
nor I_3369 (I60269,I60252,I59845);
DFFARX1 I_3370 (I59771,I60269,I2966,I59794,);
nor I_3371 (I59786,I60111,I60252);
nor I_3372 (I59774,I60252,I60015);
not I_3373 (I60328,I60252);
and I_3374 (I60345,I59879,I60328);
nor I_3375 (I59780,I60015,I60345);
nand I_3376 (I59768,I60252,I60142);
not I_3377 (I60423,I2973);
nand I_3378 (I60440,I36844,I36847);
and I_3379 (I60457,I60440,I36829);
DFFARX1 I_3380 (I60474,I60457,I2966,I60423,);
not I_3381 (I60491,I60474);
nor I_3382 (I60508,I36826,I36847);
or I_3383 (I60406,I60508,I60474);
not I_3384 (I60394,I60508);
DFFARX1 I_3385 (I60553,I36850,I2966,I60423,);
nor I_3386 (I60570,I60553,I60508);
nand I_3387 (I60587,I36835,I36841);
and I_3388 (I60604,I60587,I36853);
DFFARX1 I_3389 (I60621,I60604,I2966,I60423,);
nor I_3390 (I60403,I60621,I60474);
not I_3391 (I60652,I60621);
nor I_3392 (I60669,I60553,I60652);
DFFARX1 I_3393 (I60686,I36832,I2966,I60423,);
and I_3394 (I60703,I60686,I36823);
or I_3395 (I60412,I60703,I60508);
nand I_3396 (I60391,I60703,I60669);
DFFARX1 I_3397 (I60748,I36838,I2966,I60423,);
and I_3398 (I60765,I60748,I60491);
nor I_3399 (I60409,I60703,I60765);
nor I_3400 (I60796,I60748,I60553);
DFFARX1 I_3401 (I60400,I60796,I2966,I60423,);
nor I_3402 (I60415,I60748,I60474);
not I_3403 (I60841,I60748);
nor I_3404 (I60858,I60621,I60841);
and I_3405 (I60875,I60508,I60858);
or I_3406 (I60892,I60703,I60875);
DFFARX1 I_3407 (I60388,I60892,I2966,I60423,);
nand I_3408 (I60397,I60748,I60570);
nand I_3409 (I60385,I60748,I60652);
not I_3410 (I60984,I2973);
not I_3411 (I61001,I57918);
nor I_3412 (I61018,I57903,I57930);
nand I_3413 (I61035,I61018,I57906);
DFFARX1 I_3414 (I60958,I61035,I2966,I60984,);
nor I_3415 (I61066,I61001,I57903);
nand I_3416 (I61083,I61066,I57921);
not I_3417 (I60973,I61083);
DFFARX1 I_3418 (I60955,I61083,I2966,I60984,);
not I_3419 (I61128,I57903);
not I_3420 (I61145,I61128);
not I_3421 (I61162,I57933);
nor I_3422 (I61179,I61162,I57915);
and I_3423 (I61196,I61179,I57924);
or I_3424 (I61213,I61196,I57909);
DFFARX1 I_3425 (I61230,I61213,I2966,I60984,);
nor I_3426 (I61247,I61230,I61083);
nor I_3427 (I61264,I61230,I61145);
nand I_3428 (I60970,I61035,I61264);
nand I_3429 (I61295,I61001,I57933);
nand I_3430 (I61312,I61295,I61230);
and I_3431 (I61329,I61295,I61312);
DFFARX1 I_3432 (I60952,I61329,I2966,I60984,);
DFFARX1 I_3433 (I61360,I61295,I2966,I60984,);
and I_3434 (I60949,I61128,I61360);
DFFARX1 I_3435 (I61391,I57912,I2966,I60984,);
not I_3436 (I61408,I61391);
nor I_3437 (I61425,I61083,I61408);
and I_3438 (I61442,I61391,I61425);
nand I_3439 (I60964,I61391,I61145);
DFFARX1 I_3440 (I61473,I61391,I2966,I60984,);
not I_3441 (I60961,I61473);
DFFARX1 I_3442 (I61504,I57927,I2966,I60984,);
not I_3443 (I61521,I61504);
or I_3444 (I61538,I61521,I61442);
DFFARX1 I_3445 (I60967,I61538,I2966,I60984,);
nand I_3446 (I60976,I61521,I61247);
DFFARX1 I_3447 (I60946,I61521,I2966,I60984,);
not I_3448 (I61630,I2973);
not I_3449 (I61647,I41193);
nor I_3450 (I61664,I41190,I41178);
nand I_3451 (I61681,I61664,I41181);
DFFARX1 I_3452 (I61604,I61681,I2966,I61630,);
nor I_3453 (I61712,I61647,I41190);
nand I_3454 (I61729,I61712,I41187);
not I_3455 (I61619,I61729);
DFFARX1 I_3456 (I61601,I61729,I2966,I61630,);
not I_3457 (I61774,I41190);
not I_3458 (I61791,I61774);
not I_3459 (I61808,I41199);
nor I_3460 (I61825,I61808,I41175);
and I_3461 (I61842,I61825,I41196);
or I_3462 (I61859,I61842,I41184);
DFFARX1 I_3463 (I61876,I61859,I2966,I61630,);
nor I_3464 (I61893,I61876,I61729);
nor I_3465 (I61910,I61876,I61791);
nand I_3466 (I61616,I61681,I61910);
nand I_3467 (I61941,I61647,I41199);
nand I_3468 (I61958,I61941,I61876);
and I_3469 (I61975,I61941,I61958);
DFFARX1 I_3470 (I61598,I61975,I2966,I61630,);
DFFARX1 I_3471 (I62006,I61941,I2966,I61630,);
and I_3472 (I61595,I61774,I62006);
DFFARX1 I_3473 (I62037,I41205,I2966,I61630,);
not I_3474 (I62054,I62037);
nor I_3475 (I62071,I61729,I62054);
and I_3476 (I62088,I62037,I62071);
nand I_3477 (I61610,I62037,I61791);
DFFARX1 I_3478 (I62119,I62037,I2966,I61630,);
not I_3479 (I61607,I62119);
DFFARX1 I_3480 (I62150,I41202,I2966,I61630,);
not I_3481 (I62167,I62150);
or I_3482 (I62184,I62167,I62088);
DFFARX1 I_3483 (I61613,I62184,I2966,I61630,);
nand I_3484 (I61622,I62167,I61893);
DFFARX1 I_3485 (I61592,I62167,I2966,I61630,);
not I_3486 (I62276,I2973);
not I_3487 (I62293,I56145);
nor I_3488 (I62310,I56121,I56127);
nand I_3489 (I62327,I62310,I56130);
DFFARX1 I_3490 (I62250,I62327,I2966,I62276,);
nor I_3491 (I62358,I62293,I56121);
nand I_3492 (I62375,I62358,I56139);
not I_3493 (I62265,I62375);
DFFARX1 I_3494 (I62247,I62375,I2966,I62276,);
not I_3495 (I62420,I56121);
not I_3496 (I62437,I62420);
not I_3497 (I62454,I56118);
nor I_3498 (I62471,I62454,I56133);
and I_3499 (I62488,I62471,I56124);
or I_3500 (I62505,I62488,I56136);
DFFARX1 I_3501 (I62522,I62505,I2966,I62276,);
nor I_3502 (I62539,I62522,I62375);
nor I_3503 (I62556,I62522,I62437);
nand I_3504 (I62262,I62327,I62556);
nand I_3505 (I62587,I62293,I56118);
nand I_3506 (I62604,I62587,I62522);
and I_3507 (I62621,I62587,I62604);
DFFARX1 I_3508 (I62244,I62621,I2966,I62276,);
DFFARX1 I_3509 (I62652,I62587,I2966,I62276,);
and I_3510 (I62241,I62420,I62652);
DFFARX1 I_3511 (I62683,I56148,I2966,I62276,);
not I_3512 (I62700,I62683);
nor I_3513 (I62717,I62375,I62700);
and I_3514 (I62734,I62683,I62717);
nand I_3515 (I62256,I62683,I62437);
DFFARX1 I_3516 (I62765,I62683,I2966,I62276,);
not I_3517 (I62253,I62765);
DFFARX1 I_3518 (I62796,I56142,I2966,I62276,);
not I_3519 (I62813,I62796);
or I_3520 (I62830,I62813,I62734);
DFFARX1 I_3521 (I62259,I62830,I2966,I62276,);
nand I_3522 (I62268,I62813,I62539);
DFFARX1 I_3523 (I62238,I62813,I2966,I62276,);
not I_3524 (I62922,I2973);
not I_3525 (I62939,I48418);
nor I_3526 (I62956,I48430,I48412);
nand I_3527 (I62973,I62956,I48427);
DFFARX1 I_3528 (I62896,I62973,I2966,I62922,);
nor I_3529 (I63004,I62939,I48430);
nand I_3530 (I63021,I63004,I48415);
not I_3531 (I62911,I63021);
DFFARX1 I_3532 (I62893,I63021,I2966,I62922,);
not I_3533 (I63066,I48430);
not I_3534 (I63083,I63066);
not I_3535 (I63100,I48424);
nor I_3536 (I63117,I63100,I48403);
and I_3537 (I63134,I63117,I48406);
or I_3538 (I63151,I63134,I48409);
DFFARX1 I_3539 (I63168,I63151,I2966,I62922,);
nor I_3540 (I63185,I63168,I63021);
nor I_3541 (I63202,I63168,I63083);
nand I_3542 (I62908,I62973,I63202);
nand I_3543 (I63233,I62939,I48424);
nand I_3544 (I63250,I63233,I63168);
and I_3545 (I63267,I63233,I63250);
DFFARX1 I_3546 (I62890,I63267,I2966,I62922,);
DFFARX1 I_3547 (I63298,I63233,I2966,I62922,);
and I_3548 (I62887,I63066,I63298);
DFFARX1 I_3549 (I63329,I48400,I2966,I62922,);
not I_3550 (I63346,I63329);
nor I_3551 (I63363,I63021,I63346);
and I_3552 (I63380,I63329,I63363);
nand I_3553 (I62902,I63329,I63083);
DFFARX1 I_3554 (I63411,I63329,I2966,I62922,);
not I_3555 (I62899,I63411);
DFFARX1 I_3556 (I63442,I48421,I2966,I62922,);
not I_3557 (I63459,I63442);
or I_3558 (I63476,I63459,I63380);
DFFARX1 I_3559 (I62905,I63476,I2966,I62922,);
nand I_3560 (I62914,I63459,I63185);
DFFARX1 I_3561 (I62884,I63459,I2966,I62922,);
not I_3562 (I63568,I2973);
not I_3563 (I63585,I58498);
nor I_3564 (I63602,I58513,I58528);
nand I_3565 (I63619,I63602,I58516);
DFFARX1 I_3566 (I63542,I63619,I2966,I63568,);
nor I_3567 (I63650,I63585,I58513);
nand I_3568 (I63667,I63650,I58519);
not I_3569 (I63557,I63667);
DFFARX1 I_3570 (I63539,I63667,I2966,I63568,);
not I_3571 (I63712,I58513);
not I_3572 (I63729,I63712);
not I_3573 (I63746,I58525);
nor I_3574 (I63763,I63746,I58522);
and I_3575 (I63780,I63763,I58501);
or I_3576 (I63797,I63780,I58510);
DFFARX1 I_3577 (I63814,I63797,I2966,I63568,);
nor I_3578 (I63831,I63814,I63667);
nor I_3579 (I63848,I63814,I63729);
nand I_3580 (I63554,I63619,I63848);
nand I_3581 (I63879,I63585,I58525);
nand I_3582 (I63896,I63879,I63814);
and I_3583 (I63913,I63879,I63896);
DFFARX1 I_3584 (I63536,I63913,I2966,I63568,);
DFFARX1 I_3585 (I63944,I63879,I2966,I63568,);
and I_3586 (I63533,I63712,I63944);
DFFARX1 I_3587 (I63975,I58507,I2966,I63568,);
not I_3588 (I63992,I63975);
nor I_3589 (I64009,I63667,I63992);
and I_3590 (I64026,I63975,I64009);
nand I_3591 (I63548,I63975,I63729);
DFFARX1 I_3592 (I64057,I63975,I2966,I63568,);
not I_3593 (I63545,I64057);
DFFARX1 I_3594 (I64088,I58504,I2966,I63568,);
not I_3595 (I64105,I64088);
or I_3596 (I64122,I64105,I64026);
DFFARX1 I_3597 (I63551,I64122,I2966,I63568,);
nand I_3598 (I63560,I64105,I63831);
DFFARX1 I_3599 (I63530,I64105,I2966,I63568,);
not I_3600 (I64214,I2973);
not I_3601 (I64231,I38795);
nor I_3602 (I64248,I38825,I38804);
nand I_3603 (I64265,I64248,I38816);
DFFARX1 I_3604 (I64188,I64265,I2966,I64214,);
nor I_3605 (I64296,I64231,I38825);
nand I_3606 (I64313,I64296,I38798);
not I_3607 (I64203,I64313);
DFFARX1 I_3608 (I64185,I64313,I2966,I64214,);
not I_3609 (I64358,I38825);
not I_3610 (I64375,I64358);
not I_3611 (I64392,I38801);
nor I_3612 (I64409,I64392,I38819);
and I_3613 (I64426,I64409,I38810);
or I_3614 (I64443,I64426,I38807);
DFFARX1 I_3615 (I64460,I64443,I2966,I64214,);
nor I_3616 (I64477,I64460,I64313);
nor I_3617 (I64494,I64460,I64375);
nand I_3618 (I64200,I64265,I64494);
nand I_3619 (I64525,I64231,I38801);
nand I_3620 (I64542,I64525,I64460);
and I_3621 (I64559,I64525,I64542);
DFFARX1 I_3622 (I64182,I64559,I2966,I64214,);
DFFARX1 I_3623 (I64590,I64525,I2966,I64214,);
and I_3624 (I64179,I64358,I64590);
DFFARX1 I_3625 (I64621,I38813,I2966,I64214,);
not I_3626 (I64638,I64621);
nor I_3627 (I64655,I64313,I64638);
and I_3628 (I64672,I64621,I64655);
nand I_3629 (I64194,I64621,I64375);
DFFARX1 I_3630 (I64703,I64621,I2966,I64214,);
not I_3631 (I64191,I64703);
DFFARX1 I_3632 (I64734,I38822,I2966,I64214,);
not I_3633 (I64751,I64734);
or I_3634 (I64768,I64751,I64672);
DFFARX1 I_3635 (I64197,I64768,I2966,I64214,);
nand I_3636 (I64206,I64751,I64477);
DFFARX1 I_3637 (I64176,I64751,I2966,I64214,);
not I_3638 (I64860,I2973);
not I_3639 (I64877,I52019);
nor I_3640 (I64894,I52007,I52013);
nand I_3641 (I64911,I64894,I52004);
DFFARX1 I_3642 (I64834,I64911,I2966,I64860,);
nor I_3643 (I64942,I64877,I52007);
nand I_3644 (I64959,I64942,I52010);
not I_3645 (I64849,I64959);
DFFARX1 I_3646 (I64831,I64959,I2966,I64860,);
not I_3647 (I65004,I52007);
not I_3648 (I65021,I65004);
not I_3649 (I65038,I52022);
nor I_3650 (I65055,I65038,I52034);
and I_3651 (I65072,I65055,I52016);
or I_3652 (I65089,I65072,I52031);
DFFARX1 I_3653 (I65106,I65089,I2966,I64860,);
nor I_3654 (I65123,I65106,I64959);
nor I_3655 (I65140,I65106,I65021);
nand I_3656 (I64846,I64911,I65140);
nand I_3657 (I65171,I64877,I52022);
nand I_3658 (I65188,I65171,I65106);
and I_3659 (I65205,I65171,I65188);
DFFARX1 I_3660 (I64828,I65205,I2966,I64860,);
DFFARX1 I_3661 (I65236,I65171,I2966,I64860,);
and I_3662 (I64825,I65004,I65236);
DFFARX1 I_3663 (I65267,I52025,I2966,I64860,);
not I_3664 (I65284,I65267);
nor I_3665 (I65301,I64959,I65284);
and I_3666 (I65318,I65267,I65301);
nand I_3667 (I64840,I65267,I65021);
DFFARX1 I_3668 (I65349,I65267,I2966,I64860,);
not I_3669 (I64837,I65349);
DFFARX1 I_3670 (I65380,I52028,I2966,I64860,);
not I_3671 (I65397,I65380);
or I_3672 (I65414,I65397,I65318);
DFFARX1 I_3673 (I64843,I65414,I2966,I64860,);
nand I_3674 (I64852,I65397,I65123);
DFFARX1 I_3675 (I64822,I65397,I2966,I64860,);
not I_3676 (I65506,I2973);
not I_3677 (I65523,I49064);
nor I_3678 (I65540,I49046,I49061);
nand I_3679 (I65557,I65540,I49070);
DFFARX1 I_3680 (I65480,I65557,I2966,I65506,);
nor I_3681 (I65588,I65523,I49046);
nand I_3682 (I65605,I65588,I49073);
not I_3683 (I65495,I65605);
DFFARX1 I_3684 (I65477,I65605,I2966,I65506,);
not I_3685 (I65650,I49046);
not I_3686 (I65667,I65650);
not I_3687 (I65684,I49076);
nor I_3688 (I65701,I65684,I49052);
and I_3689 (I65718,I65701,I49055);
or I_3690 (I65735,I65718,I49049);
DFFARX1 I_3691 (I65752,I65735,I2966,I65506,);
nor I_3692 (I65769,I65752,I65605);
nor I_3693 (I65786,I65752,I65667);
nand I_3694 (I65492,I65557,I65786);
nand I_3695 (I65817,I65523,I49076);
nand I_3696 (I65834,I65817,I65752);
and I_3697 (I65851,I65817,I65834);
DFFARX1 I_3698 (I65474,I65851,I2966,I65506,);
DFFARX1 I_3699 (I65882,I65817,I2966,I65506,);
and I_3700 (I65471,I65650,I65882);
DFFARX1 I_3701 (I65913,I49058,I2966,I65506,);
not I_3702 (I65930,I65913);
nor I_3703 (I65947,I65605,I65930);
and I_3704 (I65964,I65913,I65947);
nand I_3705 (I65486,I65913,I65667);
DFFARX1 I_3706 (I65995,I65913,I2966,I65506,);
not I_3707 (I65483,I65995);
DFFARX1 I_3708 (I66026,I49067,I2966,I65506,);
not I_3709 (I66043,I66026);
or I_3710 (I66060,I66043,I65964);
DFFARX1 I_3711 (I65489,I66060,I2966,I65506,);
nand I_3712 (I65498,I66043,I65769);
DFFARX1 I_3713 (I65468,I66043,I2966,I65506,);
not I_3714 (I66152,I2973);
not I_3715 (I66169,I52582);
nor I_3716 (I66186,I52588,I52585);
nand I_3717 (I66203,I66186,I52603);
DFFARX1 I_3718 (I66123,I66203,I2966,I66152,);
nor I_3719 (I66234,I66169,I52588);
nand I_3720 (I66251,I66234,I52612);
nand I_3721 (I66268,I66251,I66203);
not I_3722 (I66285,I52588);
not I_3723 (I66302,I52606);
nor I_3724 (I66319,I66302,I52597);
and I_3725 (I66336,I66319,I52600);
or I_3726 (I66353,I66336,I52591);
DFFARX1 I_3727 (I66370,I66353,I2966,I66152,);
nor I_3728 (I66387,I66370,I66251);
nand I_3729 (I66138,I66285,I66387);
not I_3730 (I66135,I66370);
and I_3731 (I66432,I66370,I66268);
DFFARX1 I_3732 (I66120,I66432,I2966,I66152,);
DFFARX1 I_3733 (I66463,I66370,I2966,I66152,);
and I_3734 (I66117,I66285,I66463);
nand I_3735 (I66494,I66169,I52606);
not I_3736 (I66511,I66494);
nor I_3737 (I66528,I66370,I66511);
DFFARX1 I_3738 (I66545,I52609,I2966,I66152,);
nand I_3739 (I66562,I66545,I66494);
and I_3740 (I66579,I66285,I66562);
DFFARX1 I_3741 (I66144,I66579,I2966,I66152,);
not I_3742 (I66610,I66545);
nand I_3743 (I66132,I66545,I66528);
nand I_3744 (I66126,I66545,I66511);
DFFARX1 I_3745 (I66655,I52594,I2966,I66152,);
not I_3746 (I66672,I66655);
nor I_3747 (I66141,I66545,I66672);
nor I_3748 (I66703,I66672,I66610);
and I_3749 (I66720,I66251,I66703);
or I_3750 (I66737,I66494,I66720);
DFFARX1 I_3751 (I66129,I66737,I2966,I66152,);
DFFARX1 I_3752 (I66114,I66672,I2966,I66152,);
not I_3753 (I66815,I2973);
not I_3754 (I66832,I50848);
nor I_3755 (I66849,I50854,I50851);
nand I_3756 (I66866,I66849,I50869);
DFFARX1 I_3757 (I66786,I66866,I2966,I66815,);
nor I_3758 (I66897,I66832,I50854);
nand I_3759 (I66914,I66897,I50878);
nand I_3760 (I66931,I66914,I66866);
not I_3761 (I66948,I50854);
not I_3762 (I66965,I50872);
nor I_3763 (I66982,I66965,I50863);
and I_3764 (I66999,I66982,I50866);
or I_3765 (I67016,I66999,I50857);
DFFARX1 I_3766 (I67033,I67016,I2966,I66815,);
nor I_3767 (I67050,I67033,I66914);
nand I_3768 (I66801,I66948,I67050);
not I_3769 (I66798,I67033);
and I_3770 (I67095,I67033,I66931);
DFFARX1 I_3771 (I66783,I67095,I2966,I66815,);
DFFARX1 I_3772 (I67126,I67033,I2966,I66815,);
and I_3773 (I66780,I66948,I67126);
nand I_3774 (I67157,I66832,I50872);
not I_3775 (I67174,I67157);
nor I_3776 (I67191,I67033,I67174);
DFFARX1 I_3777 (I67208,I50875,I2966,I66815,);
nand I_3778 (I67225,I67208,I67157);
and I_3779 (I67242,I66948,I67225);
DFFARX1 I_3780 (I66807,I67242,I2966,I66815,);
not I_3781 (I67273,I67208);
nand I_3782 (I66795,I67208,I67191);
nand I_3783 (I66789,I67208,I67174);
DFFARX1 I_3784 (I67318,I50860,I2966,I66815,);
not I_3785 (I67335,I67318);
nor I_3786 (I66804,I67208,I67335);
nor I_3787 (I67366,I67335,I67273);
and I_3788 (I67383,I66914,I67366);
or I_3789 (I67400,I67157,I67383);
DFFARX1 I_3790 (I66792,I67400,I2966,I66815,);
DFFARX1 I_3791 (I66777,I67335,I2966,I66815,);
not I_3792 (I67478,I2973);
or I_3793 (I67495,I60967,I60961);
or I_3794 (I67512,I60955,I60967);
DFFARX1 I_3795 (I67452,I67512,I2966,I67478,);
nor I_3796 (I67543,I60973,I60964);
not I_3797 (I67560,I67543);
not I_3798 (I67577,I60973);
and I_3799 (I67594,I67577,I60970);
nor I_3800 (I67611,I67594,I60961);
nor I_3801 (I67628,I60946,I60952);
DFFARX1 I_3802 (I67645,I67628,I2966,I67478,);
nand I_3803 (I67662,I67645,I67495);
and I_3804 (I67679,I67611,I67662);
DFFARX1 I_3805 (I67446,I67679,I2966,I67478,);
nor I_3806 (I67710,I60946,I60955);
DFFARX1 I_3807 (I67727,I67710,I2966,I67478,);
and I_3808 (I67443,I67543,I67727);
DFFARX1 I_3809 (I67758,I60958,I2966,I67478,);
and I_3810 (I67775,I67758,I60976);
DFFARX1 I_3811 (I67792,I67775,I2966,I67478,);
not I_3812 (I67455,I67792);
DFFARX1 I_3813 (I67440,I67775,I2966,I67478,);
DFFARX1 I_3814 (I67837,I60949,I2966,I67478,);
not I_3815 (I67854,I67837);
nor I_3816 (I67871,I67512,I67854);
and I_3817 (I67888,I67775,I67871);
or I_3818 (I67905,I67495,I67888);
DFFARX1 I_3819 (I67461,I67905,I2966,I67478,);
nor I_3820 (I67936,I67837,I67645);
nand I_3821 (I67470,I67611,I67936);
nor I_3822 (I67967,I67837,I67560);
nand I_3823 (I67464,I67710,I67967);
not I_3824 (I67467,I67837);
nand I_3825 (I67458,I67837,I67560);
DFFARX1 I_3826 (I67449,I67837,I2966,I67478,);
not I_3827 (I68073,I2973);
or I_3828 (I68090,I66807,I66792);
or I_3829 (I68107,I66789,I66807);
DFFARX1 I_3830 (I68047,I68107,I2966,I68073,);
nor I_3831 (I68138,I66777,I66786);
not I_3832 (I68155,I68138);
not I_3833 (I68172,I66777);
and I_3834 (I68189,I68172,I66801);
nor I_3835 (I68206,I68189,I66792);
nor I_3836 (I68223,I66780,I66795);
DFFARX1 I_3837 (I68240,I68223,I2966,I68073,);
nand I_3838 (I68257,I68240,I68090);
and I_3839 (I68274,I68206,I68257);
DFFARX1 I_3840 (I68041,I68274,I2966,I68073,);
nor I_3841 (I68305,I66780,I66789);
DFFARX1 I_3842 (I68322,I68305,I2966,I68073,);
and I_3843 (I68038,I68138,I68322);
DFFARX1 I_3844 (I68353,I66783,I2966,I68073,);
and I_3845 (I68370,I68353,I66804);
DFFARX1 I_3846 (I68387,I68370,I2966,I68073,);
not I_3847 (I68050,I68387);
DFFARX1 I_3848 (I68035,I68370,I2966,I68073,);
DFFARX1 I_3849 (I68432,I66798,I2966,I68073,);
not I_3850 (I68449,I68432);
nor I_3851 (I68466,I68107,I68449);
and I_3852 (I68483,I68370,I68466);
or I_3853 (I68500,I68090,I68483);
DFFARX1 I_3854 (I68056,I68500,I2966,I68073,);
nor I_3855 (I68531,I68432,I68240);
nand I_3856 (I68065,I68206,I68531);
nor I_3857 (I68562,I68432,I68155);
nand I_3858 (I68059,I68305,I68562);
not I_3859 (I68062,I68432);
nand I_3860 (I68053,I68432,I68155);
DFFARX1 I_3861 (I68044,I68432,I2966,I68073,);
not I_3862 (I68668,I2973);
not I_3863 (I68685,I56731);
nor I_3864 (I68702,I56728,I56719);
nand I_3865 (I68719,I68702,I56722);
nor I_3866 (I68736,I68685,I56728);
nand I_3867 (I68753,I68736,I56716);
not I_3868 (I68770,I68753);
not I_3869 (I68787,I56728);
nor I_3870 (I68657,I68753,I68787);
not I_3871 (I68818,I68787);
nand I_3872 (I68642,I68753,I68818);
not I_3873 (I68849,I56737);
nor I_3874 (I68866,I68849,I56740);
and I_3875 (I68883,I68866,I56725);
or I_3876 (I68900,I68883,I56713);
DFFARX1 I_3877 (I68917,I68900,I2966,I68668,);
nor I_3878 (I68934,I68917,I68770);
DFFARX1 I_3879 (I68951,I68917,I2966,I68668,);
not I_3880 (I68639,I68951);
nand I_3881 (I68982,I68685,I56737);
and I_3882 (I68999,I68982,I68934);
DFFARX1 I_3883 (I68636,I68982,I2966,I68668,);
DFFARX1 I_3884 (I69030,I56734,I2966,I68668,);
nor I_3885 (I69047,I69030,I68753);
nand I_3886 (I68654,I68917,I69047);
nor I_3887 (I69078,I69030,I68818);
not I_3888 (I68651,I69030);
nand I_3889 (I69109,I69030,I68719);
and I_3890 (I69126,I68787,I69109);
DFFARX1 I_3891 (I68630,I69126,I2966,I68668,);
DFFARX1 I_3892 (I68633,I69030,I2966,I68668,);
DFFARX1 I_3893 (I69171,I56743,I2966,I68668,);
not I_3894 (I69188,I69171);
nand I_3895 (I69205,I69188,I68753);
and I_3896 (I69222,I68982,I69205);
DFFARX1 I_3897 (I68660,I69222,I2966,I68668,);
or I_3898 (I69253,I69188,I68999);
DFFARX1 I_3899 (I68645,I69253,I2966,I68668,);
nand I_3900 (I68648,I69188,I69078);
not I_3901 (I69331,I2973);
not I_3902 (I69348,I59762);
nor I_3903 (I69365,I59780,I59771);
nand I_3904 (I69382,I69365,I59777);
nor I_3905 (I69399,I69348,I59780);
nand I_3906 (I69416,I69399,I59783);
not I_3907 (I69433,I69416);
not I_3908 (I69450,I59780);
nor I_3909 (I69320,I69416,I69450);
not I_3910 (I69481,I69450);
nand I_3911 (I69305,I69416,I69481);
not I_3912 (I69512,I59759);
nor I_3913 (I69529,I69512,I59774);
and I_3914 (I69546,I69529,I59756);
or I_3915 (I69563,I69546,I59765);
DFFARX1 I_3916 (I69580,I69563,I2966,I69331,);
nor I_3917 (I69597,I69580,I69433);
DFFARX1 I_3918 (I69614,I69580,I2966,I69331,);
not I_3919 (I69302,I69614);
nand I_3920 (I69645,I69348,I59759);
and I_3921 (I69662,I69645,I69597);
DFFARX1 I_3922 (I69299,I69645,I2966,I69331,);
DFFARX1 I_3923 (I69693,I59768,I2966,I69331,);
nor I_3924 (I69710,I69693,I69416);
nand I_3925 (I69317,I69580,I69710);
nor I_3926 (I69741,I69693,I69481);
not I_3927 (I69314,I69693);
nand I_3928 (I69772,I69693,I69382);
and I_3929 (I69789,I69450,I69772);
DFFARX1 I_3930 (I69293,I69789,I2966,I69331,);
DFFARX1 I_3931 (I69296,I69693,I2966,I69331,);
DFFARX1 I_3932 (I69834,I59786,I2966,I69331,);
not I_3933 (I69851,I69834);
nand I_3934 (I69868,I69851,I69416);
and I_3935 (I69885,I69645,I69868);
DFFARX1 I_3936 (I69323,I69885,I2966,I69331,);
or I_3937 (I69916,I69851,I69662);
DFFARX1 I_3938 (I69308,I69916,I2966,I69331,);
nand I_3939 (I69311,I69851,I69741);
not I_3940 (I69994,I2973);
not I_3941 (I70011,I60403);
nor I_3942 (I70028,I60409,I60412);
nand I_3943 (I70045,I70028,I60388);
nor I_3944 (I70062,I70011,I60409);
nand I_3945 (I70079,I70062,I60397);
not I_3946 (I70096,I70079);
not I_3947 (I70113,I60409);
nor I_3948 (I69983,I70079,I70113);
not I_3949 (I70144,I70113);
nand I_3950 (I69968,I70079,I70144);
not I_3951 (I70175,I60391);
nor I_3952 (I70192,I70175,I60415);
and I_3953 (I70209,I70192,I60385);
or I_3954 (I70226,I70209,I60394);
DFFARX1 I_3955 (I70243,I70226,I2966,I69994,);
nor I_3956 (I70260,I70243,I70096);
DFFARX1 I_3957 (I70277,I70243,I2966,I69994,);
not I_3958 (I69965,I70277);
nand I_3959 (I70308,I70011,I60391);
and I_3960 (I70325,I70308,I70260);
DFFARX1 I_3961 (I69962,I70308,I2966,I69994,);
DFFARX1 I_3962 (I70356,I60400,I2966,I69994,);
nor I_3963 (I70373,I70356,I70079);
nand I_3964 (I69980,I70243,I70373);
nor I_3965 (I70404,I70356,I70144);
not I_3966 (I69977,I70356);
nand I_3967 (I70435,I70356,I70045);
and I_3968 (I70452,I70113,I70435);
DFFARX1 I_3969 (I69956,I70452,I2966,I69994,);
DFFARX1 I_3970 (I69959,I70356,I2966,I69994,);
DFFARX1 I_3971 (I70497,I60406,I2966,I69994,);
not I_3972 (I70514,I70497);
nand I_3973 (I70531,I70514,I70079);
and I_3974 (I70548,I70308,I70531);
DFFARX1 I_3975 (I69986,I70548,I2966,I69994,);
or I_3976 (I70579,I70514,I70325);
DFFARX1 I_3977 (I69971,I70579,I2966,I69994,);
nand I_3978 (I69974,I70514,I70404);
not I_3979 (I70657,I2973);
not I_3980 (I70674,I46474);
nor I_3981 (I70691,I46471,I46489);
nand I_3982 (I70708,I70691,I46492);
nor I_3983 (I70725,I70674,I46471);
nand I_3984 (I70742,I70725,I46477);
not I_3985 (I70759,I70742);
not I_3986 (I70776,I46471);
nor I_3987 (I70646,I70742,I70776);
not I_3988 (I70807,I70776);
nand I_3989 (I70631,I70742,I70807);
not I_3990 (I70838,I46486);
nor I_3991 (I70855,I70838,I46468);
and I_3992 (I70872,I70855,I46462);
or I_3993 (I70889,I70872,I46480);
DFFARX1 I_3994 (I70906,I70889,I2966,I70657,);
nor I_3995 (I70923,I70906,I70759);
DFFARX1 I_3996 (I70940,I70906,I2966,I70657,);
not I_3997 (I70628,I70940);
nand I_3998 (I70971,I70674,I46486);
and I_3999 (I70988,I70971,I70923);
DFFARX1 I_4000 (I70625,I70971,I2966,I70657,);
DFFARX1 I_4001 (I71019,I46465,I2966,I70657,);
nor I_4002 (I71036,I71019,I70742);
nand I_4003 (I70643,I70906,I71036);
nor I_4004 (I71067,I71019,I70807);
not I_4005 (I70640,I71019);
nand I_4006 (I71098,I71019,I70708);
and I_4007 (I71115,I70776,I71098);
DFFARX1 I_4008 (I70619,I71115,I2966,I70657,);
DFFARX1 I_4009 (I70622,I71019,I2966,I70657,);
DFFARX1 I_4010 (I71160,I46483,I2966,I70657,);
not I_4011 (I71177,I71160);
nand I_4012 (I71194,I71177,I70742);
and I_4013 (I71211,I70971,I71194);
DFFARX1 I_4014 (I70649,I71211,I2966,I70657,);
or I_4015 (I71242,I71177,I70988);
DFFARX1 I_4016 (I70634,I71242,I2966,I70657,);
nand I_4017 (I70637,I71177,I71067);
not I_4018 (I71320,I2973);
not I_4019 (I71337,I50285);
nor I_4020 (I71354,I50297,I50279);
nand I_4021 (I71371,I71354,I50300);
nor I_4022 (I71388,I71337,I50297);
nand I_4023 (I71405,I71388,I50291);
not I_4024 (I71422,I71405);
not I_4025 (I71439,I50297);
nor I_4026 (I71309,I71405,I71439);
not I_4027 (I71470,I71439);
nand I_4028 (I71294,I71405,I71470);
not I_4029 (I71501,I50282);
nor I_4030 (I71518,I71501,I50276);
and I_4031 (I71535,I71518,I50288);
or I_4032 (I71552,I71535,I50273);
DFFARX1 I_4033 (I71569,I71552,I2966,I71320,);
nor I_4034 (I71586,I71569,I71422);
DFFARX1 I_4035 (I71603,I71569,I2966,I71320,);
not I_4036 (I71291,I71603);
nand I_4037 (I71634,I71337,I50282);
and I_4038 (I71651,I71634,I71586);
DFFARX1 I_4039 (I71288,I71634,I2966,I71320,);
DFFARX1 I_4040 (I71682,I50270,I2966,I71320,);
nor I_4041 (I71699,I71682,I71405);
nand I_4042 (I71306,I71569,I71699);
nor I_4043 (I71730,I71682,I71470);
not I_4044 (I71303,I71682);
nand I_4045 (I71761,I71682,I71371);
and I_4046 (I71778,I71439,I71761);
DFFARX1 I_4047 (I71282,I71778,I2966,I71320,);
DFFARX1 I_4048 (I71285,I71682,I2966,I71320,);
DFFARX1 I_4049 (I71823,I50294,I2966,I71320,);
not I_4050 (I71840,I71823);
nand I_4051 (I71857,I71840,I71405);
and I_4052 (I71874,I71634,I71857);
DFFARX1 I_4053 (I71312,I71874,I2966,I71320,);
or I_4054 (I71905,I71840,I71651);
DFFARX1 I_4055 (I71297,I71905,I2966,I71320,);
nand I_4056 (I71300,I71840,I71730);
not I_4057 (I71983,I2973);
not I_4058 (I72000,I51441);
nor I_4059 (I72017,I51453,I51435);
nand I_4060 (I72034,I72017,I51456);
nor I_4061 (I72051,I72000,I51453);
nand I_4062 (I72068,I72051,I51447);
not I_4063 (I72085,I72068);
not I_4064 (I72102,I51453);
nor I_4065 (I71972,I72068,I72102);
not I_4066 (I72133,I72102);
nand I_4067 (I71957,I72068,I72133);
not I_4068 (I72164,I51438);
nor I_4069 (I72181,I72164,I51432);
and I_4070 (I72198,I72181,I51444);
or I_4071 (I72215,I72198,I51429);
DFFARX1 I_4072 (I72232,I72215,I2966,I71983,);
nor I_4073 (I72249,I72232,I72085);
DFFARX1 I_4074 (I72266,I72232,I2966,I71983,);
not I_4075 (I71954,I72266);
nand I_4076 (I72297,I72000,I51438);
and I_4077 (I72314,I72297,I72249);
DFFARX1 I_4078 (I71951,I72297,I2966,I71983,);
DFFARX1 I_4079 (I72345,I51426,I2966,I71983,);
nor I_4080 (I72362,I72345,I72068);
nand I_4081 (I71969,I72232,I72362);
nor I_4082 (I72393,I72345,I72133);
not I_4083 (I71966,I72345);
nand I_4084 (I72424,I72345,I72034);
and I_4085 (I72441,I72102,I72424);
DFFARX1 I_4086 (I71945,I72441,I2966,I71983,);
DFFARX1 I_4087 (I71948,I72345,I2966,I71983,);
DFFARX1 I_4088 (I72486,I51450,I2966,I71983,);
not I_4089 (I72503,I72486);
nand I_4090 (I72520,I72503,I72068);
and I_4091 (I72537,I72297,I72520);
DFFARX1 I_4092 (I71975,I72537,I2966,I71983,);
or I_4093 (I72568,I72503,I72314);
DFFARX1 I_4094 (I71960,I72568,I2966,I71983,);
nand I_4095 (I71963,I72503,I72393);
not I_4096 (I72646,I2973);
not I_4097 (I72663,I65474);
nor I_4098 (I72680,I65471,I65495);
nand I_4099 (I72697,I72680,I65492);
nor I_4100 (I72714,I72663,I65471);
nand I_4101 (I72731,I72714,I65498);
not I_4102 (I72748,I72731);
not I_4103 (I72765,I65471);
nor I_4104 (I72635,I72731,I72765);
not I_4105 (I72796,I72765);
nand I_4106 (I72620,I72731,I72796);
not I_4107 (I72827,I65489);
nor I_4108 (I72844,I72827,I65480);
and I_4109 (I72861,I72844,I65477);
or I_4110 (I72878,I72861,I65486);
DFFARX1 I_4111 (I72895,I72878,I2966,I72646,);
nor I_4112 (I72912,I72895,I72748);
DFFARX1 I_4113 (I72929,I72895,I2966,I72646,);
not I_4114 (I72617,I72929);
nand I_4115 (I72960,I72663,I65489);
and I_4116 (I72977,I72960,I72912);
DFFARX1 I_4117 (I72614,I72960,I2966,I72646,);
DFFARX1 I_4118 (I73008,I65468,I2966,I72646,);
nor I_4119 (I73025,I73008,I72731);
nand I_4120 (I72632,I72895,I73025);
nor I_4121 (I73056,I73008,I72796);
not I_4122 (I72629,I73008);
nand I_4123 (I73087,I73008,I72697);
and I_4124 (I73104,I72765,I73087);
DFFARX1 I_4125 (I72608,I73104,I2966,I72646,);
DFFARX1 I_4126 (I72611,I73008,I2966,I72646,);
DFFARX1 I_4127 (I73149,I65483,I2966,I72646,);
not I_4128 (I73166,I73149);
nand I_4129 (I73183,I73166,I72731);
and I_4130 (I73200,I72960,I73183);
DFFARX1 I_4131 (I72638,I73200,I2966,I72646,);
or I_4132 (I73231,I73166,I72977);
DFFARX1 I_4133 (I72623,I73231,I2966,I72646,);
nand I_4134 (I72626,I73166,I73056);
not I_4135 (I73309,I2973);
not I_4136 (I73326,I49676);
nor I_4137 (I73343,I49685,I49670);
nand I_4138 (I73360,I73343,I49658);
nor I_4139 (I73377,I73326,I49685);
nand I_4140 (I73394,I73377,I49661);
DFFARX1 I_4141 (I73411,I73394,I2966,I73309,);
not I_4142 (I73280,I73411);
not I_4143 (I73442,I49685);
not I_4144 (I73459,I73442);
not I_4145 (I73476,I49673);
nor I_4146 (I73493,I73476,I49667);
and I_4147 (I73510,I73493,I49664);
or I_4148 (I73527,I73510,I49679);
DFFARX1 I_4149 (I73544,I73527,I2966,I73309,);
DFFARX1 I_4150 (I73277,I73544,I2966,I73309,);
DFFARX1 I_4151 (I73575,I73544,I2966,I73309,);
DFFARX1 I_4152 (I73271,I73544,I2966,I73309,);
nand I_4153 (I73606,I73326,I49673);
nand I_4154 (I73623,I73606,I73360);
and I_4155 (I73640,I73442,I73623);
DFFARX1 I_4156 (I73301,I73640,I2966,I73309,);
and I_4157 (I73274,I73606,I73575);
DFFARX1 I_4158 (I73685,I49688,I2966,I73309,);
nor I_4159 (I73298,I73685,I73606);
nor I_4160 (I73716,I73685,I73360);
nand I_4161 (I73295,I73394,I73716);
not I_4162 (I73292,I73685);
DFFARX1 I_4163 (I73761,I49682,I2966,I73309,);
not I_4164 (I73778,I73761);
nor I_4165 (I73795,I73778,I73459);
and I_4166 (I73812,I73685,I73795);
or I_4167 (I73829,I73606,I73812);
DFFARX1 I_4168 (I73286,I73829,I2966,I73309,);
not I_4169 (I73860,I73778);
nor I_4170 (I73877,I73685,I73860);
nand I_4171 (I73289,I73778,I73877);
nand I_4172 (I73283,I73442,I73860);
not I_4173 (I73955,I2973);
not I_4174 (I73972,I62905);
nor I_4175 (I73989,I62896,I62887);
nand I_4176 (I74006,I73989,I62902);
nor I_4177 (I74023,I73972,I62896);
nand I_4178 (I74040,I74023,I62899);
DFFARX1 I_4179 (I74057,I74040,I2966,I73955,);
not I_4180 (I73926,I74057);
not I_4181 (I74088,I62896);
not I_4182 (I74105,I74088);
not I_4183 (I74122,I62908);
nor I_4184 (I74139,I74122,I62893);
and I_4185 (I74156,I74139,I62911);
or I_4186 (I74173,I74156,I62884);
DFFARX1 I_4187 (I74190,I74173,I2966,I73955,);
DFFARX1 I_4188 (I73923,I74190,I2966,I73955,);
DFFARX1 I_4189 (I74221,I74190,I2966,I73955,);
DFFARX1 I_4190 (I73917,I74190,I2966,I73955,);
nand I_4191 (I74252,I73972,I62908);
nand I_4192 (I74269,I74252,I74006);
and I_4193 (I74286,I74088,I74269);
DFFARX1 I_4194 (I73947,I74286,I2966,I73955,);
and I_4195 (I73920,I74252,I74221);
DFFARX1 I_4196 (I74331,I62914,I2966,I73955,);
nor I_4197 (I73944,I74331,I74252);
nor I_4198 (I74362,I74331,I74006);
nand I_4199 (I73941,I74040,I74362);
not I_4200 (I73938,I74331);
DFFARX1 I_4201 (I74407,I62890,I2966,I73955,);
not I_4202 (I74424,I74407);
nor I_4203 (I74441,I74424,I74105);
and I_4204 (I74458,I74331,I74441);
or I_4205 (I74475,I74252,I74458);
DFFARX1 I_4206 (I73932,I74475,I2966,I73955,);
not I_4207 (I74506,I74424);
nor I_4208 (I74523,I74331,I74506);
nand I_4209 (I73935,I74424,I74523);
nand I_4210 (I73929,I74088,I74506);
not I_4211 (I74601,I2973);
not I_4212 (I74618,I53747);
nor I_4213 (I74635,I53759,I53753);
nand I_4214 (I74652,I74635,I53738);
nor I_4215 (I74669,I74618,I53759);
nand I_4216 (I74686,I74669,I53765);
DFFARX1 I_4217 (I74703,I74686,I2966,I74601,);
not I_4218 (I74572,I74703);
not I_4219 (I74734,I53759);
not I_4220 (I74751,I74734);
not I_4221 (I74768,I53762);
nor I_4222 (I74785,I74768,I53744);
and I_4223 (I74802,I74785,I53741);
or I_4224 (I74819,I74802,I53768);
DFFARX1 I_4225 (I74836,I74819,I2966,I74601,);
DFFARX1 I_4226 (I74569,I74836,I2966,I74601,);
DFFARX1 I_4227 (I74867,I74836,I2966,I74601,);
DFFARX1 I_4228 (I74563,I74836,I2966,I74601,);
nand I_4229 (I74898,I74618,I53762);
nand I_4230 (I74915,I74898,I74652);
and I_4231 (I74932,I74734,I74915);
DFFARX1 I_4232 (I74593,I74932,I2966,I74601,);
and I_4233 (I74566,I74898,I74867);
DFFARX1 I_4234 (I74977,I53756,I2966,I74601,);
nor I_4235 (I74590,I74977,I74898);
nor I_4236 (I75008,I74977,I74652);
nand I_4237 (I74587,I74686,I75008);
not I_4238 (I74584,I74977);
DFFARX1 I_4239 (I75053,I53750,I2966,I74601,);
not I_4240 (I75070,I75053);
nor I_4241 (I75087,I75070,I74751);
and I_4242 (I75104,I74977,I75087);
or I_4243 (I75121,I74898,I75104);
DFFARX1 I_4244 (I74578,I75121,I2966,I74601,);
not I_4245 (I75152,I75070);
nor I_4246 (I75169,I74977,I75152);
nand I_4247 (I74581,I75070,I75169);
nand I_4248 (I74575,I74734,I75152);
not I_4249 (I75247,I2973);
not I_4250 (I75264,I72632);
nor I_4251 (I75281,I72611,I72623);
nand I_4252 (I75298,I75281,I72626);
nor I_4253 (I75315,I75264,I72611);
nand I_4254 (I75332,I75315,I72608);
DFFARX1 I_4255 (I75349,I75332,I2966,I75247,);
not I_4256 (I75218,I75349);
not I_4257 (I75380,I72611);
not I_4258 (I75397,I75380);
not I_4259 (I75414,I72629);
nor I_4260 (I75431,I75414,I72620);
and I_4261 (I75448,I75431,I72614);
or I_4262 (I75465,I75448,I72638);
DFFARX1 I_4263 (I75482,I75465,I2966,I75247,);
DFFARX1 I_4264 (I75215,I75482,I2966,I75247,);
DFFARX1 I_4265 (I75513,I75482,I2966,I75247,);
DFFARX1 I_4266 (I75209,I75482,I2966,I75247,);
nand I_4267 (I75544,I75264,I72629);
nand I_4268 (I75561,I75544,I75298);
and I_4269 (I75578,I75380,I75561);
DFFARX1 I_4270 (I75239,I75578,I2966,I75247,);
and I_4271 (I75212,I75544,I75513);
DFFARX1 I_4272 (I75623,I72635,I2966,I75247,);
nor I_4273 (I75236,I75623,I75544);
nor I_4274 (I75654,I75623,I75298);
nand I_4275 (I75233,I75332,I75654);
not I_4276 (I75230,I75623);
DFFARX1 I_4277 (I75699,I72617,I2966,I75247,);
not I_4278 (I75716,I75699);
nor I_4279 (I75733,I75716,I75397);
and I_4280 (I75750,I75623,I75733);
or I_4281 (I75767,I75544,I75750);
DFFARX1 I_4282 (I75224,I75767,I2966,I75247,);
not I_4283 (I75798,I75716);
nor I_4284 (I75815,I75623,I75798);
nand I_4285 (I75227,I75716,I75815);
nand I_4286 (I75221,I75380,I75798);
not I_4287 (I75893,I2973);
not I_4288 (I75910,I64197);
nor I_4289 (I75927,I64188,I64179);
nand I_4290 (I75944,I75927,I64194);
nor I_4291 (I75961,I75910,I64188);
nand I_4292 (I75978,I75961,I64191);
DFFARX1 I_4293 (I75995,I75978,I2966,I75893,);
not I_4294 (I75864,I75995);
not I_4295 (I76026,I64188);
not I_4296 (I76043,I76026);
not I_4297 (I76060,I64200);
nor I_4298 (I76077,I76060,I64185);
and I_4299 (I76094,I76077,I64203);
or I_4300 (I76111,I76094,I64176);
DFFARX1 I_4301 (I76128,I76111,I2966,I75893,);
DFFARX1 I_4302 (I75861,I76128,I2966,I75893,);
DFFARX1 I_4303 (I76159,I76128,I2966,I75893,);
DFFARX1 I_4304 (I75855,I76128,I2966,I75893,);
nand I_4305 (I76190,I75910,I64200);
nand I_4306 (I76207,I76190,I75944);
and I_4307 (I76224,I76026,I76207);
DFFARX1 I_4308 (I75885,I76224,I2966,I75893,);
and I_4309 (I75858,I76190,I76159);
DFFARX1 I_4310 (I76269,I64206,I2966,I75893,);
nor I_4311 (I75882,I76269,I76190);
nor I_4312 (I76300,I76269,I75944);
nand I_4313 (I75879,I75978,I76300);
not I_4314 (I75876,I76269);
DFFARX1 I_4315 (I76345,I64182,I2966,I75893,);
not I_4316 (I76362,I76345);
nor I_4317 (I76379,I76362,I76043);
and I_4318 (I76396,I76269,I76379);
or I_4319 (I76413,I76190,I76396);
DFFARX1 I_4320 (I75870,I76413,I2966,I75893,);
not I_4321 (I76444,I76362);
nor I_4322 (I76461,I76269,I76444);
nand I_4323 (I75873,I76362,I76461);
nand I_4324 (I75867,I76026,I76444);
not I_4325 (I76539,I2973);
nand I_4326 (I76556,I70622,I70649);
and I_4327 (I76573,I76556,I70637);
DFFARX1 I_4328 (I76590,I76573,I2966,I76539,);
not I_4329 (I76607,I76590);
DFFARX1 I_4330 (I76507,I76590,I2966,I76539,);
nor I_4331 (I76638,I70625,I70649);
DFFARX1 I_4332 (I76655,I70640,I2966,I76539,);
DFFARX1 I_4333 (I76672,I76655,I2966,I76539,);
not I_4334 (I76510,I76672);
DFFARX1 I_4335 (I76703,I76655,I2966,I76539,);
and I_4336 (I76504,I76590,I76703);
nand I_4337 (I76734,I70634,I70631);
and I_4338 (I76751,I76734,I70628);
DFFARX1 I_4339 (I76768,I76751,I2966,I76539,);
nor I_4340 (I76785,I76768,I76607);
not I_4341 (I76802,I76768);
nand I_4342 (I76513,I76590,I76802);
DFFARX1 I_4343 (I76833,I70643,I2966,I76539,);
and I_4344 (I76850,I76833,I70619);
nor I_4345 (I76867,I76850,I76768);
nor I_4346 (I76884,I76850,I76802);
nand I_4347 (I76519,I76638,I76884);
not I_4348 (I76522,I76850);
DFFARX1 I_4349 (I76501,I76850,I2966,I76539,);
DFFARX1 I_4350 (I76943,I70646,I2966,I76539,);
nand I_4351 (I76960,I76943,I76655);
and I_4352 (I76977,I76638,I76960);
DFFARX1 I_4353 (I76531,I76977,I2966,I76539,);
nor I_4354 (I76528,I76943,I76850);
and I_4355 (I77022,I76943,I76785);
or I_4356 (I77039,I76638,I77022);
DFFARX1 I_4357 (I76516,I77039,I2966,I76539,);
nand I_4358 (I76525,I76943,I76867);
not I_4359 (I77117,I2973);
nand I_4360 (I77134,I69959,I69986);
and I_4361 (I77151,I77134,I69974);
DFFARX1 I_4362 (I77168,I77151,I2966,I77117,);
not I_4363 (I77185,I77168);
DFFARX1 I_4364 (I77085,I77168,I2966,I77117,);
nor I_4365 (I77216,I69962,I69986);
DFFARX1 I_4366 (I77233,I69977,I2966,I77117,);
DFFARX1 I_4367 (I77250,I77233,I2966,I77117,);
not I_4368 (I77088,I77250);
DFFARX1 I_4369 (I77281,I77233,I2966,I77117,);
and I_4370 (I77082,I77168,I77281);
nand I_4371 (I77312,I69971,I69968);
and I_4372 (I77329,I77312,I69965);
DFFARX1 I_4373 (I77346,I77329,I2966,I77117,);
nor I_4374 (I77363,I77346,I77185);
not I_4375 (I77380,I77346);
nand I_4376 (I77091,I77168,I77380);
DFFARX1 I_4377 (I77411,I69980,I2966,I77117,);
and I_4378 (I77428,I77411,I69956);
nor I_4379 (I77445,I77428,I77346);
nor I_4380 (I77462,I77428,I77380);
nand I_4381 (I77097,I77216,I77462);
not I_4382 (I77100,I77428);
DFFARX1 I_4383 (I77079,I77428,I2966,I77117,);
DFFARX1 I_4384 (I77521,I69983,I2966,I77117,);
nand I_4385 (I77538,I77521,I77233);
and I_4386 (I77555,I77216,I77538);
DFFARX1 I_4387 (I77109,I77555,I2966,I77117,);
nor I_4388 (I77106,I77521,I77428);
and I_4389 (I77600,I77521,I77363);
or I_4390 (I77617,I77216,I77600);
DFFARX1 I_4391 (I77094,I77617,I2966,I77117,);
nand I_4392 (I77103,I77521,I77445);
not I_4393 (I77695,I2973);
nand I_4394 (I77712,I67464,I67449);
and I_4395 (I77729,I77712,I67458);
DFFARX1 I_4396 (I77746,I77729,I2966,I77695,);
not I_4397 (I77763,I77746);
DFFARX1 I_4398 (I77663,I77746,I2966,I77695,);
nor I_4399 (I77794,I67467,I67449);
DFFARX1 I_4400 (I77811,I67446,I2966,I77695,);
DFFARX1 I_4401 (I77828,I77811,I2966,I77695,);
not I_4402 (I77666,I77828);
DFFARX1 I_4403 (I77859,I77811,I2966,I77695,);
and I_4404 (I77660,I77746,I77859);
nand I_4405 (I77890,I67470,I67443);
and I_4406 (I77907,I77890,I67461);
DFFARX1 I_4407 (I77924,I77907,I2966,I77695,);
nor I_4408 (I77941,I77924,I77763);
not I_4409 (I77958,I77924);
nand I_4410 (I77669,I77746,I77958);
DFFARX1 I_4411 (I77989,I67455,I2966,I77695,);
and I_4412 (I78006,I77989,I67440);
nor I_4413 (I78023,I78006,I77924);
nor I_4414 (I78040,I78006,I77958);
nand I_4415 (I77675,I77794,I78040);
not I_4416 (I77678,I78006);
DFFARX1 I_4417 (I77657,I78006,I2966,I77695,);
DFFARX1 I_4418 (I78099,I67452,I2966,I77695,);
nand I_4419 (I78116,I78099,I77811);
and I_4420 (I78133,I77794,I78116);
DFFARX1 I_4421 (I77687,I78133,I2966,I77695,);
nor I_4422 (I77684,I78099,I78006);
and I_4423 (I78178,I78099,I77941);
or I_4424 (I78195,I77794,I78178);
DFFARX1 I_4425 (I77672,I78195,I2966,I77695,);
nand I_4426 (I77681,I78099,I78023);
not I_4427 (I78273,I2973);
nand I_4428 (I78290,I57323,I57314);
and I_4429 (I78307,I78290,I57332);
DFFARX1 I_4430 (I78324,I78307,I2966,I78273,);
nor I_4431 (I78341,I57311,I57314);
nor I_4432 (I78358,I78341,I78324);
not I_4433 (I78256,I78341);
DFFARX1 I_4434 (I78389,I57320,I2966,I78273,);
not I_4435 (I78406,I78389);
nor I_4436 (I78423,I78341,I78406);
nand I_4437 (I78259,I78389,I78358);
DFFARX1 I_4438 (I78241,I78389,I2966,I78273,);
nand I_4439 (I78468,I57335,I57317);
and I_4440 (I78485,I78468,I57338);
DFFARX1 I_4441 (I78502,I78485,I2966,I78273,);
nor I_4442 (I78262,I78502,I78324);
nand I_4443 (I78253,I78502,I78423);
DFFARX1 I_4444 (I78547,I57326,I2966,I78273,);
and I_4445 (I78564,I78547,I57308);
DFFARX1 I_4446 (I78581,I78564,I2966,I78273,);
not I_4447 (I78244,I78581);
nand I_4448 (I78612,I78564,I78502);
and I_4449 (I78629,I78324,I78612);
DFFARX1 I_4450 (I78235,I78629,I2966,I78273,);
DFFARX1 I_4451 (I78660,I57329,I2966,I78273,);
nand I_4452 (I78677,I78660,I78324);
and I_4453 (I78694,I78502,I78677);
DFFARX1 I_4454 (I78265,I78694,I2966,I78273,);
not I_4455 (I78725,I78660);
nor I_4456 (I78742,I78341,I78725);
and I_4457 (I78759,I78660,I78742);
or I_4458 (I78776,I78564,I78759);
DFFARX1 I_4459 (I78250,I78776,I2966,I78273,);
nand I_4460 (I78247,I78660,I78406);
DFFARX1 I_4461 (I78238,I78660,I2966,I78273,);
not I_4462 (I78868,I2973);
nand I_4463 (I78885,I73289,I73301);
and I_4464 (I78902,I78885,I73283);
DFFARX1 I_4465 (I78919,I78902,I2966,I78868,);
nor I_4466 (I78936,I73295,I73301);
nor I_4467 (I78953,I78936,I78919);
not I_4468 (I78851,I78936);
DFFARX1 I_4469 (I78984,I73280,I2966,I78868,);
not I_4470 (I79001,I78984);
nor I_4471 (I79018,I78936,I79001);
nand I_4472 (I78854,I78984,I78953);
DFFARX1 I_4473 (I78836,I78984,I2966,I78868,);
nand I_4474 (I79063,I73271,I73286);
and I_4475 (I79080,I79063,I73277);
DFFARX1 I_4476 (I79097,I79080,I2966,I78868,);
nor I_4477 (I78857,I79097,I78919);
nand I_4478 (I78848,I79097,I79018);
DFFARX1 I_4479 (I79142,I73298,I2966,I78868,);
and I_4480 (I79159,I79142,I73292);
DFFARX1 I_4481 (I79176,I79159,I2966,I78868,);
not I_4482 (I78839,I79176);
nand I_4483 (I79207,I79159,I79097);
and I_4484 (I79224,I78919,I79207);
DFFARX1 I_4485 (I78830,I79224,I2966,I78868,);
DFFARX1 I_4486 (I79255,I73274,I2966,I78868,);
nand I_4487 (I79272,I79255,I78919);
and I_4488 (I79289,I79097,I79272);
DFFARX1 I_4489 (I78860,I79289,I2966,I78868,);
not I_4490 (I79320,I79255);
nor I_4491 (I79337,I78936,I79320);
and I_4492 (I79354,I79255,I79337);
or I_4493 (I79371,I79159,I79354);
DFFARX1 I_4494 (I78845,I79371,I2966,I78868,);
nand I_4495 (I78842,I79255,I79001);
DFFARX1 I_4496 (I78833,I79255,I2966,I78868,);
not I_4497 (I79463,I2973);
nand I_4498 (I79480,I64831,I64843);
and I_4499 (I79497,I79480,I64852);
DFFARX1 I_4500 (I79514,I79497,I2966,I79463,);
nor I_4501 (I79531,I64846,I64843);
nor I_4502 (I79548,I79531,I79514);
not I_4503 (I79446,I79531);
DFFARX1 I_4504 (I79579,I64840,I2966,I79463,);
not I_4505 (I79596,I79579);
nor I_4506 (I79613,I79531,I79596);
nand I_4507 (I79449,I79579,I79548);
DFFARX1 I_4508 (I79431,I79579,I2966,I79463,);
nand I_4509 (I79658,I64837,I64834);
and I_4510 (I79675,I79658,I64825);
DFFARX1 I_4511 (I79692,I79675,I2966,I79463,);
nor I_4512 (I79452,I79692,I79514);
nand I_4513 (I79443,I79692,I79613);
DFFARX1 I_4514 (I79737,I64849,I2966,I79463,);
and I_4515 (I79754,I79737,I64828);
DFFARX1 I_4516 (I79771,I79754,I2966,I79463,);
not I_4517 (I79434,I79771);
nand I_4518 (I79802,I79754,I79692);
and I_4519 (I79819,I79514,I79802);
DFFARX1 I_4520 (I79425,I79819,I2966,I79463,);
DFFARX1 I_4521 (I79850,I64822,I2966,I79463,);
nand I_4522 (I79867,I79850,I79514);
and I_4523 (I79884,I79692,I79867);
DFFARX1 I_4524 (I79455,I79884,I2966,I79463,);
not I_4525 (I79915,I79850);
nor I_4526 (I79932,I79531,I79915);
and I_4527 (I79949,I79850,I79932);
or I_4528 (I79966,I79754,I79949);
DFFARX1 I_4529 (I79440,I79966,I2966,I79463,);
nand I_4530 (I79437,I79850,I79596);
DFFARX1 I_4531 (I79428,I79850,I2966,I79463,);
not I_4532 (I80058,I2973);
nand I_4533 (I80075,I66132,I66144);
and I_4534 (I80092,I80075,I66123);
DFFARX1 I_4535 (I80109,I80092,I2966,I80058,);
nor I_4536 (I80126,I66114,I66144);
nor I_4537 (I80143,I80126,I80109);
not I_4538 (I80041,I80126);
DFFARX1 I_4539 (I80174,I66126,I2966,I80058,);
not I_4540 (I80191,I80174);
nor I_4541 (I80208,I80126,I80191);
nand I_4542 (I80044,I80174,I80143);
DFFARX1 I_4543 (I80026,I80174,I2966,I80058,);
nand I_4544 (I80253,I66141,I66129);
and I_4545 (I80270,I80253,I66117);
DFFARX1 I_4546 (I80287,I80270,I2966,I80058,);
nor I_4547 (I80047,I80287,I80109);
nand I_4548 (I80038,I80287,I80208);
DFFARX1 I_4549 (I80332,I66135,I2966,I80058,);
and I_4550 (I80349,I80332,I66120);
DFFARX1 I_4551 (I80366,I80349,I2966,I80058,);
not I_4552 (I80029,I80366);
nand I_4553 (I80397,I80349,I80287);
and I_4554 (I80414,I80109,I80397);
DFFARX1 I_4555 (I80020,I80414,I2966,I80058,);
DFFARX1 I_4556 (I80445,I66138,I2966,I80058,);
nand I_4557 (I80462,I80445,I80109);
and I_4558 (I80479,I80287,I80462);
DFFARX1 I_4559 (I80050,I80479,I2966,I80058,);
not I_4560 (I80510,I80445);
nor I_4561 (I80527,I80126,I80510);
and I_4562 (I80544,I80445,I80527);
or I_4563 (I80561,I80349,I80544);
DFFARX1 I_4564 (I80035,I80561,I2966,I80058,);
nand I_4565 (I80032,I80445,I80191);
DFFARX1 I_4566 (I80023,I80445,I2966,I80058,);
not I_4567 (I80653,I2973);
nand I_4568 (I80670,I75227,I75239);
and I_4569 (I80687,I80670,I75230);
DFFARX1 I_4570 (I80704,I80687,I2966,I80653,);
nor I_4571 (I80721,I75224,I75239);
DFFARX1 I_4572 (I80738,I75215,I2966,I80653,);
nand I_4573 (I80755,I80738,I80721);
DFFARX1 I_4574 (I80624,I80738,I2966,I80653,);
nand I_4575 (I80786,I75221,I75212);
and I_4576 (I80803,I80786,I75218);
DFFARX1 I_4577 (I80820,I80803,I2966,I80653,);
not I_4578 (I80837,I80820);
nor I_4579 (I80854,I80704,I80837);
and I_4580 (I80871,I80721,I80854);
and I_4581 (I80888,I80820,I80755);
DFFARX1 I_4582 (I80621,I80888,I2966,I80653,);
DFFARX1 I_4583 (I80615,I80820,I2966,I80653,);
DFFARX1 I_4584 (I80933,I75233,I2966,I80653,);
and I_4585 (I80950,I80933,I75209);
nand I_4586 (I80967,I80950,I80820);
nor I_4587 (I80642,I80950,I80721);
not I_4588 (I80998,I80950);
nor I_4589 (I81015,I80704,I80998);
nand I_4590 (I80633,I80738,I81015);
nand I_4591 (I80627,I80820,I80998);
or I_4592 (I81060,I80950,I80871);
DFFARX1 I_4593 (I80630,I81060,I2966,I80653,);
DFFARX1 I_4594 (I81091,I75236,I2966,I80653,);
and I_4595 (I81108,I81091,I80967);
DFFARX1 I_4596 (I80645,I81108,I2966,I80653,);
nor I_4597 (I81139,I81091,I80704);
nand I_4598 (I80639,I80950,I81139);
not I_4599 (I80636,I81091);
DFFARX1 I_4600 (I81184,I81091,I2966,I80653,);
and I_4601 (I80618,I81091,I81184);
not I_4602 (I81248,I2973);
nand I_4603 (I81265,I59157,I59145);
and I_4604 (I81282,I81265,I59130);
DFFARX1 I_4605 (I81299,I81282,I2966,I81248,);
nor I_4606 (I81316,I59142,I59145);
DFFARX1 I_4607 (I81333,I59154,I2966,I81248,);
nand I_4608 (I81350,I81333,I81316);
DFFARX1 I_4609 (I81219,I81333,I2966,I81248,);
nand I_4610 (I81381,I59127,I59151);
and I_4611 (I81398,I81381,I59136);
DFFARX1 I_4612 (I81415,I81398,I2966,I81248,);
not I_4613 (I81432,I81415);
nor I_4614 (I81449,I81299,I81432);
and I_4615 (I81466,I81316,I81449);
and I_4616 (I81483,I81415,I81350);
DFFARX1 I_4617 (I81216,I81483,I2966,I81248,);
DFFARX1 I_4618 (I81210,I81415,I2966,I81248,);
DFFARX1 I_4619 (I81528,I59139,I2966,I81248,);
and I_4620 (I81545,I81528,I59148);
nand I_4621 (I81562,I81545,I81415);
nor I_4622 (I81237,I81545,I81316);
not I_4623 (I81593,I81545);
nor I_4624 (I81610,I81299,I81593);
nand I_4625 (I81228,I81333,I81610);
nand I_4626 (I81222,I81415,I81593);
or I_4627 (I81655,I81545,I81466);
DFFARX1 I_4628 (I81225,I81655,I2966,I81248,);
DFFARX1 I_4629 (I81686,I59133,I2966,I81248,);
and I_4630 (I81703,I81686,I81562);
DFFARX1 I_4631 (I81240,I81703,I2966,I81248,);
nor I_4632 (I81734,I81686,I81299);
nand I_4633 (I81234,I81545,I81734);
not I_4634 (I81231,I81686);
DFFARX1 I_4635 (I81779,I81686,I2966,I81248,);
and I_4636 (I81213,I81686,I81779);
not I_4637 (I81843,I2973);
nand I_4638 (I81860,I79440,I79425);
and I_4639 (I81877,I81860,I79431);
DFFARX1 I_4640 (I81894,I81877,I2966,I81843,);
nor I_4641 (I81911,I79434,I79425);
DFFARX1 I_4642 (I81928,I79446,I2966,I81843,);
nand I_4643 (I81945,I81928,I81911);
DFFARX1 I_4644 (I81814,I81928,I2966,I81843,);
nand I_4645 (I81976,I79437,I79428);
and I_4646 (I81993,I81976,I79455);
DFFARX1 I_4647 (I82010,I81993,I2966,I81843,);
not I_4648 (I82027,I82010);
nor I_4649 (I82044,I81894,I82027);
and I_4650 (I82061,I81911,I82044);
and I_4651 (I82078,I82010,I81945);
DFFARX1 I_4652 (I81811,I82078,I2966,I81843,);
DFFARX1 I_4653 (I81805,I82010,I2966,I81843,);
DFFARX1 I_4654 (I82123,I79443,I2966,I81843,);
and I_4655 (I82140,I82123,I79449);
nand I_4656 (I82157,I82140,I82010);
nor I_4657 (I81832,I82140,I81911);
not I_4658 (I82188,I82140);
nor I_4659 (I82205,I81894,I82188);
nand I_4660 (I81823,I81928,I82205);
nand I_4661 (I81817,I82010,I82188);
or I_4662 (I82250,I82140,I82061);
DFFARX1 I_4663 (I81820,I82250,I2966,I81843,);
DFFARX1 I_4664 (I82281,I79452,I2966,I81843,);
and I_4665 (I82298,I82281,I82157);
DFFARX1 I_4666 (I81835,I82298,I2966,I81843,);
nor I_4667 (I82329,I82281,I81894);
nand I_4668 (I81829,I82140,I82329);
not I_4669 (I81826,I82281);
DFFARX1 I_4670 (I82374,I82281,I2966,I81843,);
and I_4671 (I81808,I82281,I82374);
not I_4672 (I82438,I2973);
nand I_4673 (I82455,I78250,I78235);
and I_4674 (I82472,I82455,I78241);
DFFARX1 I_4675 (I82489,I82472,I2966,I82438,);
nor I_4676 (I82506,I78244,I78235);
DFFARX1 I_4677 (I82523,I78256,I2966,I82438,);
nand I_4678 (I82540,I82523,I82506);
DFFARX1 I_4679 (I82409,I82523,I2966,I82438,);
nand I_4680 (I82571,I78247,I78238);
and I_4681 (I82588,I82571,I78265);
DFFARX1 I_4682 (I82605,I82588,I2966,I82438,);
not I_4683 (I82622,I82605);
nor I_4684 (I82639,I82489,I82622);
and I_4685 (I82656,I82506,I82639);
and I_4686 (I82673,I82605,I82540);
DFFARX1 I_4687 (I82406,I82673,I2966,I82438,);
DFFARX1 I_4688 (I82400,I82605,I2966,I82438,);
DFFARX1 I_4689 (I82718,I78253,I2966,I82438,);
and I_4690 (I82735,I82718,I78259);
nand I_4691 (I82752,I82735,I82605);
nor I_4692 (I82427,I82735,I82506);
not I_4693 (I82783,I82735);
nor I_4694 (I82800,I82489,I82783);
nand I_4695 (I82418,I82523,I82800);
nand I_4696 (I82412,I82605,I82783);
or I_4697 (I82845,I82735,I82656);
DFFARX1 I_4698 (I82415,I82845,I2966,I82438,);
DFFARX1 I_4699 (I82876,I78262,I2966,I82438,);
and I_4700 (I82893,I82876,I82752);
DFFARX1 I_4701 (I82430,I82893,I2966,I82438,);
nor I_4702 (I82924,I82876,I82489);
nand I_4703 (I82424,I82735,I82924);
not I_4704 (I82421,I82876);
DFFARX1 I_4705 (I82969,I82876,I2966,I82438,);
and I_4706 (I82403,I82876,I82969);
not I_4707 (I83033,I2973);
not I_4708 (I83050,I71963);
nor I_4709 (I83067,I71969,I71948);
nand I_4710 (I83084,I83067,I71954);
nor I_4711 (I83101,I83050,I71969);
nand I_4712 (I83118,I83101,I71960);
not I_4713 (I83135,I71969);
not I_4714 (I83152,I83135);
not I_4715 (I83169,I71957);
nor I_4716 (I83186,I83169,I71975);
and I_4717 (I83203,I83186,I71966);
or I_4718 (I83220,I83203,I71945);
DFFARX1 I_4719 (I83237,I83220,I2966,I83033,);
nand I_4720 (I83254,I83050,I71957);
or I_4721 (I83022,I83254,I83237);
not I_4722 (I83285,I83254);
nor I_4723 (I83302,I83237,I83285);
and I_4724 (I83319,I83135,I83302);
nand I_4725 (I82995,I83254,I83152);
DFFARX1 I_4726 (I83350,I71972,I2966,I83033,);
or I_4727 (I83016,I83350,I83237);
nor I_4728 (I83381,I83350,I83118);
nor I_4729 (I83398,I83350,I83152);
nand I_4730 (I83001,I83084,I83398);
or I_4731 (I83429,I83350,I83319);
DFFARX1 I_4732 (I82998,I83429,I2966,I83033,);
not I_4733 (I83004,I83350);
DFFARX1 I_4734 (I83474,I71951,I2966,I83033,);
not I_4735 (I83491,I83474);
nor I_4736 (I83508,I83491,I83084);
DFFARX1 I_4737 (I83010,I83508,I2966,I83033,);
nor I_4738 (I83025,I83350,I83491);
nor I_4739 (I83013,I83491,I83254);
not I_4740 (I83567,I83491);
and I_4741 (I83584,I83118,I83567);
nor I_4742 (I83019,I83254,I83584);
nand I_4743 (I83007,I83491,I83381);
not I_4744 (I83662,I2973);
not I_4745 (I83679,I73935);
nor I_4746 (I83696,I73944,I73947);
nand I_4747 (I83713,I83696,I73932);
nor I_4748 (I83730,I83679,I73944);
nand I_4749 (I83747,I83730,I73929);
not I_4750 (I83764,I73944);
not I_4751 (I83781,I83764);
not I_4752 (I83798,I73917);
nor I_4753 (I83815,I83798,I73923);
and I_4754 (I83832,I83815,I73920);
or I_4755 (I83849,I83832,I73941);
DFFARX1 I_4756 (I83866,I83849,I2966,I83662,);
nand I_4757 (I83883,I83679,I73917);
or I_4758 (I83651,I83883,I83866);
not I_4759 (I83914,I83883);
nor I_4760 (I83931,I83866,I83914);
and I_4761 (I83948,I83764,I83931);
nand I_4762 (I83624,I83883,I83781);
DFFARX1 I_4763 (I83979,I73926,I2966,I83662,);
or I_4764 (I83645,I83979,I83866);
nor I_4765 (I84010,I83979,I83747);
nor I_4766 (I84027,I83979,I83781);
nand I_4767 (I83630,I83713,I84027);
or I_4768 (I84058,I83979,I83948);
DFFARX1 I_4769 (I83627,I84058,I2966,I83662,);
not I_4770 (I83633,I83979);
DFFARX1 I_4771 (I84103,I73938,I2966,I83662,);
not I_4772 (I84120,I84103);
nor I_4773 (I84137,I84120,I83713);
DFFARX1 I_4774 (I83639,I84137,I2966,I83662,);
nor I_4775 (I83654,I83979,I84120);
nor I_4776 (I83642,I84120,I83883);
not I_4777 (I84196,I84120);
and I_4778 (I84213,I83747,I84196);
nor I_4779 (I83648,I83883,I84213);
nand I_4780 (I83636,I84120,I84010);
not I_4781 (I84291,I2973);
not I_4782 (I84308,I63536);
nor I_4783 (I84325,I63554,I63533);
nand I_4784 (I84342,I84325,I63551);
nor I_4785 (I84359,I84308,I63554);
nand I_4786 (I84376,I84359,I63545);
not I_4787 (I84393,I63554);
not I_4788 (I84410,I84393);
not I_4789 (I84427,I63548);
nor I_4790 (I84444,I84427,I63542);
and I_4791 (I84461,I84444,I63539);
or I_4792 (I84478,I84461,I63530);
DFFARX1 I_4793 (I84495,I84478,I2966,I84291,);
nand I_4794 (I84512,I84308,I63548);
or I_4795 (I84280,I84512,I84495);
not I_4796 (I84543,I84512);
nor I_4797 (I84560,I84495,I84543);
and I_4798 (I84577,I84393,I84560);
nand I_4799 (I84253,I84512,I84410);
DFFARX1 I_4800 (I84608,I63560,I2966,I84291,);
or I_4801 (I84274,I84608,I84495);
nor I_4802 (I84639,I84608,I84376);
nor I_4803 (I84656,I84608,I84410);
nand I_4804 (I84259,I84342,I84656);
or I_4805 (I84687,I84608,I84577);
DFFARX1 I_4806 (I84256,I84687,I2966,I84291,);
not I_4807 (I84262,I84608);
DFFARX1 I_4808 (I84732,I63557,I2966,I84291,);
not I_4809 (I84749,I84732);
nor I_4810 (I84766,I84749,I84342);
DFFARX1 I_4811 (I84268,I84766,I2966,I84291,);
nor I_4812 (I84283,I84608,I84749);
nor I_4813 (I84271,I84749,I84512);
not I_4814 (I84825,I84749);
and I_4815 (I84842,I84376,I84825);
nor I_4816 (I84277,I84512,I84842);
nand I_4817 (I84265,I84749,I84639);
not I_4818 (I84920,I2973);
not I_4819 (I84937,I74581);
nor I_4820 (I84954,I74590,I74593);
nand I_4821 (I84971,I84954,I74578);
nor I_4822 (I84988,I84937,I74590);
nand I_4823 (I85005,I84988,I74575);
not I_4824 (I85022,I74590);
not I_4825 (I85039,I85022);
not I_4826 (I85056,I74563);
nor I_4827 (I85073,I85056,I74569);
and I_4828 (I85090,I85073,I74566);
or I_4829 (I85107,I85090,I74587);
DFFARX1 I_4830 (I85124,I85107,I2966,I84920,);
nand I_4831 (I85141,I84937,I74563);
or I_4832 (I84909,I85141,I85124);
not I_4833 (I85172,I85141);
nor I_4834 (I85189,I85124,I85172);
and I_4835 (I85206,I85022,I85189);
nand I_4836 (I84882,I85141,I85039);
DFFARX1 I_4837 (I85237,I74572,I2966,I84920,);
or I_4838 (I84903,I85237,I85124);
nor I_4839 (I85268,I85237,I85005);
nor I_4840 (I85285,I85237,I85039);
nand I_4841 (I84888,I84971,I85285);
or I_4842 (I85316,I85237,I85206);
DFFARX1 I_4843 (I84885,I85316,I2966,I84920,);
not I_4844 (I84891,I85237);
DFFARX1 I_4845 (I85361,I74584,I2966,I84920,);
not I_4846 (I85378,I85361);
nor I_4847 (I85395,I85378,I84971);
DFFARX1 I_4848 (I84897,I85395,I2966,I84920,);
nor I_4849 (I84912,I85237,I85378);
nor I_4850 (I84900,I85378,I85141);
not I_4851 (I85454,I85378);
and I_4852 (I85471,I85005,I85454);
nor I_4853 (I84906,I85141,I85471);
nand I_4854 (I84894,I85378,I85268);
not I_4855 (I85549,I2973);
nand I_4856 (I85566,I61613,I61598);
and I_4857 (I85583,I85566,I61592);
DFFARX1 I_4858 (I85600,I85583,I2966,I85549,);
not I_4859 (I85538,I85600);
DFFARX1 I_4860 (I85631,I85600,I2966,I85549,);
not I_4861 (I85526,I85631);
nor I_4862 (I85662,I61619,I61598);
not I_4863 (I85679,I85662);
nor I_4864 (I85696,I85600,I85679);
DFFARX1 I_4865 (I85713,I61622,I2966,I85549,);
not I_4866 (I85730,I85713);
nand I_4867 (I85529,I85713,I85679);
DFFARX1 I_4868 (I85761,I85713,I2966,I85549,);
and I_4869 (I85514,I85600,I85761);
nand I_4870 (I85792,I61604,I61607);
and I_4871 (I85809,I85792,I61610);
DFFARX1 I_4872 (I85826,I85809,I2966,I85549,);
nor I_4873 (I85843,I85826,I85730);
and I_4874 (I85860,I85662,I85843);
nor I_4875 (I85877,I85826,I85600);
DFFARX1 I_4876 (I85520,I85826,I2966,I85549,);
DFFARX1 I_4877 (I85908,I61616,I2966,I85549,);
and I_4878 (I85925,I85908,I61601);
or I_4879 (I85942,I85925,I85860);
DFFARX1 I_4880 (I85532,I85942,I2966,I85549,);
nand I_4881 (I85541,I85925,I85877);
DFFARX1 I_4882 (I85511,I85925,I2966,I85549,);
DFFARX1 I_4883 (I86001,I61595,I2966,I85549,);
nand I_4884 (I85535,I86001,I85696);
DFFARX1 I_4885 (I85523,I86001,I2966,I85549,);
nand I_4886 (I86046,I86001,I85662);
and I_4887 (I86063,I85713,I86046);
DFFARX1 I_4888 (I85517,I86063,I2966,I85549,);
not I_4889 (I86127,I2973);
nand I_4890 (I86144,I76513,I76510);
and I_4891 (I86161,I86144,I76504);
DFFARX1 I_4892 (I86178,I86161,I2966,I86127,);
not I_4893 (I86195,I86178);
nor I_4894 (I86212,I76516,I76510);
or I_4895 (I86110,I86212,I86178);
not I_4896 (I86098,I86212);
DFFARX1 I_4897 (I86257,I76528,I2966,I86127,);
nor I_4898 (I86274,I86257,I86212);
nand I_4899 (I86291,I76519,I76501);
and I_4900 (I86308,I86291,I76531);
DFFARX1 I_4901 (I86325,I86308,I2966,I86127,);
nor I_4902 (I86107,I86325,I86178);
not I_4903 (I86356,I86325);
nor I_4904 (I86373,I86257,I86356);
DFFARX1 I_4905 (I86390,I76507,I2966,I86127,);
and I_4906 (I86407,I86390,I76525);
or I_4907 (I86116,I86407,I86212);
nand I_4908 (I86095,I86407,I86373);
DFFARX1 I_4909 (I86452,I76522,I2966,I86127,);
and I_4910 (I86469,I86452,I86195);
nor I_4911 (I86113,I86407,I86469);
nor I_4912 (I86500,I86452,I86257);
DFFARX1 I_4913 (I86104,I86500,I2966,I86127,);
nor I_4914 (I86119,I86452,I86178);
not I_4915 (I86545,I86452);
nor I_4916 (I86562,I86325,I86545);
and I_4917 (I86579,I86212,I86562);
or I_4918 (I86596,I86407,I86579);
DFFARX1 I_4919 (I86092,I86596,I2966,I86127,);
nand I_4920 (I86101,I86452,I86274);
nand I_4921 (I86089,I86452,I86356);
not I_4922 (I86688,I2973);
nand I_4923 (I86705,I62259,I62262);
and I_4924 (I86722,I86705,I62244);
DFFARX1 I_4925 (I86739,I86722,I2966,I86688,);
not I_4926 (I86756,I86739);
nor I_4927 (I86773,I62241,I62262);
or I_4928 (I86671,I86773,I86739);
not I_4929 (I86659,I86773);
DFFARX1 I_4930 (I86818,I62265,I2966,I86688,);
nor I_4931 (I86835,I86818,I86773);
nand I_4932 (I86852,I62250,I62256);
and I_4933 (I86869,I86852,I62268);
DFFARX1 I_4934 (I86886,I86869,I2966,I86688,);
nor I_4935 (I86668,I86886,I86739);
not I_4936 (I86917,I86886);
nor I_4937 (I86934,I86818,I86917);
DFFARX1 I_4938 (I86951,I62247,I2966,I86688,);
and I_4939 (I86968,I86951,I62238);
or I_4940 (I86677,I86968,I86773);
nand I_4941 (I86656,I86968,I86934);
DFFARX1 I_4942 (I87013,I62253,I2966,I86688,);
and I_4943 (I87030,I87013,I86756);
nor I_4944 (I86674,I86968,I87030);
nor I_4945 (I87061,I87013,I86818);
DFFARX1 I_4946 (I86665,I87061,I2966,I86688,);
nor I_4947 (I86680,I87013,I86739);
not I_4948 (I87106,I87013);
nor I_4949 (I87123,I86886,I87106);
and I_4950 (I87140,I86773,I87123);
or I_4951 (I87157,I86968,I87140);
DFFARX1 I_4952 (I86653,I87157,I2966,I86688,);
nand I_4953 (I86662,I87013,I86835);
nand I_4954 (I86650,I87013,I86917);
not I_4955 (I87249,I2973);
nand I_4956 (I87266,I71306,I71297);
and I_4957 (I87283,I87266,I71312);
DFFARX1 I_4958 (I87300,I87283,I2966,I87249,);
not I_4959 (I87317,I87300);
nor I_4960 (I87334,I71282,I71297);
or I_4961 (I87232,I87334,I87300);
not I_4962 (I87220,I87334);
DFFARX1 I_4963 (I87379,I71285,I2966,I87249,);
nor I_4964 (I87396,I87379,I87334);
nand I_4965 (I87413,I71303,I71300);
and I_4966 (I87430,I87413,I71288);
DFFARX1 I_4967 (I87447,I87430,I2966,I87249,);
nor I_4968 (I87229,I87447,I87300);
not I_4969 (I87478,I87447);
nor I_4970 (I87495,I87379,I87478);
DFFARX1 I_4971 (I87512,I71309,I2966,I87249,);
and I_4972 (I87529,I87512,I71294);
or I_4973 (I87238,I87529,I87334);
nand I_4974 (I87217,I87529,I87495);
DFFARX1 I_4975 (I87574,I71291,I2966,I87249,);
and I_4976 (I87591,I87574,I87317);
nor I_4977 (I87235,I87529,I87591);
nor I_4978 (I87622,I87574,I87379);
DFFARX1 I_4979 (I87226,I87622,I2966,I87249,);
nor I_4980 (I87241,I87574,I87300);
not I_4981 (I87667,I87574);
nor I_4982 (I87684,I87447,I87667);
and I_4983 (I87701,I87334,I87684);
or I_4984 (I87718,I87529,I87701);
DFFARX1 I_4985 (I87214,I87718,I2966,I87249,);
nand I_4986 (I87223,I87574,I87396);
nand I_4987 (I87211,I87574,I87478);
not I_4988 (I87810,I2973);
not I_4989 (I87827,I68648);
nor I_4990 (I87844,I68645,I68633);
nand I_4991 (I87861,I87844,I68636);
DFFARX1 I_4992 (I87784,I87861,I2966,I87810,);
nor I_4993 (I87892,I87827,I68645);
nand I_4994 (I87909,I87892,I68642);
not I_4995 (I87799,I87909);
DFFARX1 I_4996 (I87781,I87909,I2966,I87810,);
not I_4997 (I87954,I68645);
not I_4998 (I87971,I87954);
not I_4999 (I87988,I68654);
nor I_5000 (I88005,I87988,I68630);
and I_5001 (I88022,I88005,I68651);
or I_5002 (I88039,I88022,I68639);
DFFARX1 I_5003 (I88056,I88039,I2966,I87810,);
nor I_5004 (I88073,I88056,I87909);
nor I_5005 (I88090,I88056,I87971);
nand I_5006 (I87796,I87861,I88090);
nand I_5007 (I88121,I87827,I68654);
nand I_5008 (I88138,I88121,I88056);
and I_5009 (I88155,I88121,I88138);
DFFARX1 I_5010 (I87778,I88155,I2966,I87810,);
DFFARX1 I_5011 (I88186,I88121,I2966,I87810,);
and I_5012 (I87775,I87954,I88186);
DFFARX1 I_5013 (I88217,I68660,I2966,I87810,);
not I_5014 (I88234,I88217);
nor I_5015 (I88251,I87909,I88234);
and I_5016 (I88268,I88217,I88251);
nand I_5017 (I87790,I88217,I87971);
DFFARX1 I_5018 (I88299,I88217,I2966,I87810,);
not I_5019 (I87787,I88299);
DFFARX1 I_5020 (I88330,I68657,I2966,I87810,);
not I_5021 (I88347,I88330);
or I_5022 (I88364,I88347,I88268);
DFFARX1 I_5023 (I87793,I88364,I2966,I87810,);
nand I_5024 (I87802,I88347,I88073);
DFFARX1 I_5025 (I87772,I88347,I2966,I87810,);
not I_5026 (I88456,I2973);
not I_5027 (I88473,I82995);
nor I_5028 (I88490,I83010,I83025);
nand I_5029 (I88507,I88490,I83013);
DFFARX1 I_5030 (I88430,I88507,I2966,I88456,);
nor I_5031 (I88538,I88473,I83010);
nand I_5032 (I88555,I88538,I83016);
not I_5033 (I88445,I88555);
DFFARX1 I_5034 (I88427,I88555,I2966,I88456,);
not I_5035 (I88600,I83010);
not I_5036 (I88617,I88600);
not I_5037 (I88634,I83022);
nor I_5038 (I88651,I88634,I83019);
and I_5039 (I88668,I88651,I82998);
or I_5040 (I88685,I88668,I83007);
DFFARX1 I_5041 (I88702,I88685,I2966,I88456,);
nor I_5042 (I88719,I88702,I88555);
nor I_5043 (I88736,I88702,I88617);
nand I_5044 (I88442,I88507,I88736);
nand I_5045 (I88767,I88473,I83022);
nand I_5046 (I88784,I88767,I88702);
and I_5047 (I88801,I88767,I88784);
DFFARX1 I_5048 (I88424,I88801,I2966,I88456,);
DFFARX1 I_5049 (I88832,I88767,I2966,I88456,);
and I_5050 (I88421,I88600,I88832);
DFFARX1 I_5051 (I88863,I83004,I2966,I88456,);
not I_5052 (I88880,I88863);
nor I_5053 (I88897,I88555,I88880);
and I_5054 (I88914,I88863,I88897);
nand I_5055 (I88436,I88863,I88617);
DFFARX1 I_5056 (I88945,I88863,I2966,I88456,);
not I_5057 (I88433,I88945);
DFFARX1 I_5058 (I88976,I83001,I2966,I88456,);
not I_5059 (I88993,I88976);
or I_5060 (I89010,I88993,I88914);
DFFARX1 I_5061 (I88439,I89010,I2966,I88456,);
nand I_5062 (I88448,I88993,I88719);
DFFARX1 I_5063 (I88418,I88993,I2966,I88456,);
not I_5064 (I89102,I2973);
not I_5065 (I89119,I80047);
nor I_5066 (I89136,I80023,I80029);
nand I_5067 (I89153,I89136,I80032);
DFFARX1 I_5068 (I89076,I89153,I2966,I89102,);
nor I_5069 (I89184,I89119,I80023);
nand I_5070 (I89201,I89184,I80041);
not I_5071 (I89091,I89201);
DFFARX1 I_5072 (I89073,I89201,I2966,I89102,);
not I_5073 (I89246,I80023);
not I_5074 (I89263,I89246);
not I_5075 (I89280,I80020);
nor I_5076 (I89297,I89280,I80035);
and I_5077 (I89314,I89297,I80026);
or I_5078 (I89331,I89314,I80038);
DFFARX1 I_5079 (I89348,I89331,I2966,I89102,);
nor I_5080 (I89365,I89348,I89201);
nor I_5081 (I89382,I89348,I89263);
nand I_5082 (I89088,I89153,I89382);
nand I_5083 (I89413,I89119,I80020);
nand I_5084 (I89430,I89413,I89348);
and I_5085 (I89447,I89413,I89430);
DFFARX1 I_5086 (I89070,I89447,I2966,I89102,);
DFFARX1 I_5087 (I89478,I89413,I2966,I89102,);
and I_5088 (I89067,I89246,I89478);
DFFARX1 I_5089 (I89509,I80050,I2966,I89102,);
not I_5090 (I89526,I89509);
nor I_5091 (I89543,I89201,I89526);
and I_5092 (I89560,I89509,I89543);
nand I_5093 (I89082,I89509,I89263);
DFFARX1 I_5094 (I89591,I89509,I2966,I89102,);
not I_5095 (I89079,I89591);
DFFARX1 I_5096 (I89622,I80044,I2966,I89102,);
not I_5097 (I89639,I89622);
or I_5098 (I89656,I89639,I89560);
DFFARX1 I_5099 (I89085,I89656,I2966,I89102,);
nand I_5100 (I89094,I89639,I89365);
DFFARX1 I_5101 (I89064,I89639,I2966,I89102,);
not I_5102 (I89748,I2973);
not I_5103 (I89765,I83624);
nor I_5104 (I89782,I83639,I83654);
nand I_5105 (I89799,I89782,I83642);
DFFARX1 I_5106 (I89722,I89799,I2966,I89748,);
nor I_5107 (I89830,I89765,I83639);
nand I_5108 (I89847,I89830,I83645);
not I_5109 (I89737,I89847);
DFFARX1 I_5110 (I89719,I89847,I2966,I89748,);
not I_5111 (I89892,I83639);
not I_5112 (I89909,I89892);
not I_5113 (I89926,I83651);
nor I_5114 (I89943,I89926,I83648);
and I_5115 (I89960,I89943,I83627);
or I_5116 (I89977,I89960,I83636);
DFFARX1 I_5117 (I89994,I89977,I2966,I89748,);
nor I_5118 (I90011,I89994,I89847);
nor I_5119 (I90028,I89994,I89909);
nand I_5120 (I89734,I89799,I90028);
nand I_5121 (I90059,I89765,I83651);
nand I_5122 (I90076,I90059,I89994);
and I_5123 (I90093,I90059,I90076);
DFFARX1 I_5124 (I89716,I90093,I2966,I89748,);
DFFARX1 I_5125 (I90124,I90059,I2966,I89748,);
and I_5126 (I89713,I89892,I90124);
DFFARX1 I_5127 (I90155,I83633,I2966,I89748,);
not I_5128 (I90172,I90155);
nor I_5129 (I90189,I89847,I90172);
and I_5130 (I90206,I90155,I90189);
nand I_5131 (I89728,I90155,I89909);
DFFARX1 I_5132 (I90237,I90155,I2966,I89748,);
not I_5133 (I89725,I90237);
DFFARX1 I_5134 (I90268,I83630,I2966,I89748,);
not I_5135 (I90285,I90268);
or I_5136 (I90302,I90285,I90206);
DFFARX1 I_5137 (I89731,I90302,I2966,I89748,);
nand I_5138 (I89740,I90285,I90011);
DFFARX1 I_5139 (I89710,I90285,I2966,I89748,);
not I_5140 (I90394,I2973);
not I_5141 (I90411,I68059);
nor I_5142 (I90428,I68041,I68035);
nand I_5143 (I90445,I90428,I68038);
DFFARX1 I_5144 (I90365,I90445,I2966,I90394,);
nor I_5145 (I90476,I90411,I68041);
nand I_5146 (I90493,I90476,I68047);
nand I_5147 (I90510,I90493,I90445);
not I_5148 (I90527,I68041);
not I_5149 (I90544,I68056);
nor I_5150 (I90561,I90544,I68044);
and I_5151 (I90578,I90561,I68050);
or I_5152 (I90595,I90578,I68065);
DFFARX1 I_5153 (I90612,I90595,I2966,I90394,);
nor I_5154 (I90629,I90612,I90493);
nand I_5155 (I90380,I90527,I90629);
not I_5156 (I90377,I90612);
and I_5157 (I90674,I90612,I90510);
DFFARX1 I_5158 (I90362,I90674,I2966,I90394,);
DFFARX1 I_5159 (I90705,I90612,I2966,I90394,);
and I_5160 (I90359,I90527,I90705);
nand I_5161 (I90736,I90411,I68056);
not I_5162 (I90753,I90736);
nor I_5163 (I90770,I90612,I90753);
DFFARX1 I_5164 (I90787,I68053,I2966,I90394,);
nand I_5165 (I90804,I90787,I90736);
and I_5166 (I90821,I90527,I90804);
DFFARX1 I_5167 (I90386,I90821,I2966,I90394,);
not I_5168 (I90852,I90787);
nand I_5169 (I90374,I90787,I90770);
nand I_5170 (I90368,I90787,I90753);
DFFARX1 I_5171 (I90897,I68062,I2966,I90394,);
not I_5172 (I90914,I90897);
nor I_5173 (I90383,I90787,I90914);
nor I_5174 (I90945,I90914,I90852);
and I_5175 (I90962,I90493,I90945);
or I_5176 (I90979,I90736,I90962);
DFFARX1 I_5177 (I90371,I90979,I2966,I90394,);
DFFARX1 I_5178 (I90356,I90914,I2966,I90394,);
not I_5179 (I91057,I2973);
not I_5180 (I91074,I75873);
nor I_5181 (I91091,I75882,I75855);
nand I_5182 (I91108,I91091,I75867);
DFFARX1 I_5183 (I91028,I91108,I2966,I91057,);
nor I_5184 (I91139,I91074,I75882);
nand I_5185 (I91156,I91139,I75879);
nand I_5186 (I91173,I91156,I91108);
not I_5187 (I91190,I75882);
not I_5188 (I91207,I75858);
nor I_5189 (I91224,I91207,I75864);
and I_5190 (I91241,I91224,I75876);
or I_5191 (I91258,I91241,I75861);
DFFARX1 I_5192 (I91275,I91258,I2966,I91057,);
nor I_5193 (I91292,I91275,I91156);
nand I_5194 (I91043,I91190,I91292);
not I_5195 (I91040,I91275);
and I_5196 (I91337,I91275,I91173);
DFFARX1 I_5197 (I91025,I91337,I2966,I91057,);
DFFARX1 I_5198 (I91368,I91275,I2966,I91057,);
and I_5199 (I91022,I91190,I91368);
nand I_5200 (I91399,I91074,I75858);
not I_5201 (I91416,I91399);
nor I_5202 (I91433,I91275,I91416);
DFFARX1 I_5203 (I91450,I75885,I2966,I91057,);
nand I_5204 (I91467,I91450,I91399);
and I_5205 (I91484,I91190,I91467);
DFFARX1 I_5206 (I91049,I91484,I2966,I91057,);
not I_5207 (I91515,I91450);
nand I_5208 (I91037,I91450,I91433);
nand I_5209 (I91031,I91450,I91416);
DFFARX1 I_5210 (I91560,I75870,I2966,I91057,);
not I_5211 (I91577,I91560);
nor I_5212 (I91046,I91450,I91577);
nor I_5213 (I91608,I91577,I91515);
and I_5214 (I91625,I91156,I91608);
or I_5215 (I91642,I91399,I91625);
DFFARX1 I_5216 (I91034,I91642,I2966,I91057,);
DFFARX1 I_5217 (I91019,I91577,I2966,I91057,);
not I_5218 (I91720,I2973);
not I_5219 (I91737,I80621);
nor I_5220 (I91754,I80636,I80618);
nand I_5221 (I91771,I91754,I80630);
DFFARX1 I_5222 (I91691,I91771,I2966,I91720,);
nor I_5223 (I91802,I91737,I80636);
nand I_5224 (I91819,I91802,I80627);
nand I_5225 (I91836,I91819,I91771);
not I_5226 (I91853,I80636);
not I_5227 (I91870,I80645);
nor I_5228 (I91887,I91870,I80615);
and I_5229 (I91904,I91887,I80624);
or I_5230 (I91921,I91904,I80642);
DFFARX1 I_5231 (I91938,I91921,I2966,I91720,);
nor I_5232 (I91955,I91938,I91819);
nand I_5233 (I91706,I91853,I91955);
not I_5234 (I91703,I91938);
and I_5235 (I92000,I91938,I91836);
DFFARX1 I_5236 (I91688,I92000,I2966,I91720,);
DFFARX1 I_5237 (I92031,I91938,I2966,I91720,);
and I_5238 (I91685,I91853,I92031);
nand I_5239 (I92062,I91737,I80645);
not I_5240 (I92079,I92062);
nor I_5241 (I92096,I91938,I92079);
DFFARX1 I_5242 (I92113,I80633,I2966,I91720,);
nand I_5243 (I92130,I92113,I92062);
and I_5244 (I92147,I91853,I92130);
DFFARX1 I_5245 (I91712,I92147,I2966,I91720,);
not I_5246 (I92178,I92113);
nand I_5247 (I91700,I92113,I92096);
nand I_5248 (I91694,I92113,I92079);
DFFARX1 I_5249 (I92223,I80639,I2966,I91720,);
not I_5250 (I92240,I92223);
nor I_5251 (I91709,I92113,I92240);
nor I_5252 (I92271,I92240,I92178);
and I_5253 (I92288,I91819,I92271);
or I_5254 (I92305,I92062,I92288);
DFFARX1 I_5255 (I91697,I92305,I2966,I91720,);
DFFARX1 I_5256 (I91682,I92240,I2966,I91720,);
not I_5257 (I92383,I2973);
or I_5258 (I92400,I69293,I69308);
or I_5259 (I92417,I69296,I69293);
DFFARX1 I_5260 (I92357,I92417,I2966,I92383,);
nor I_5261 (I92448,I69299,I69314);
not I_5262 (I92465,I92448);
not I_5263 (I92482,I69299);
and I_5264 (I92499,I92482,I69302);
nor I_5265 (I92516,I92499,I69308);
nor I_5266 (I92533,I69305,I69323);
DFFARX1 I_5267 (I92550,I92533,I2966,I92383,);
nand I_5268 (I92567,I92550,I92400);
and I_5269 (I92584,I92516,I92567);
DFFARX1 I_5270 (I92351,I92584,I2966,I92383,);
nor I_5271 (I92615,I69305,I69296);
DFFARX1 I_5272 (I92632,I92615,I2966,I92383,);
and I_5273 (I92348,I92448,I92632);
DFFARX1 I_5274 (I92663,I69320,I2966,I92383,);
and I_5275 (I92680,I92663,I69311);
DFFARX1 I_5276 (I92697,I92680,I2966,I92383,);
not I_5277 (I92360,I92697);
DFFARX1 I_5278 (I92345,I92680,I2966,I92383,);
DFFARX1 I_5279 (I92742,I69317,I2966,I92383,);
not I_5280 (I92759,I92742);
nor I_5281 (I92776,I92417,I92759);
and I_5282 (I92793,I92680,I92776);
or I_5283 (I92810,I92400,I92793);
DFFARX1 I_5284 (I92366,I92810,I2966,I92383,);
nor I_5285 (I92841,I92742,I92550);
nand I_5286 (I92375,I92516,I92841);
nor I_5287 (I92872,I92742,I92465);
nand I_5288 (I92369,I92615,I92872);
not I_5289 (I92372,I92742);
nand I_5290 (I92363,I92742,I92465);
DFFARX1 I_5291 (I92354,I92742,I2966,I92383,);
not I_5292 (I92978,I2973);
not I_5293 (I92995,I77094);
nor I_5294 (I93012,I77106,I77088);
nand I_5295 (I93029,I93012,I77109);
nor I_5296 (I93046,I92995,I77106);
nand I_5297 (I93063,I93046,I77100);
not I_5298 (I93080,I93063);
not I_5299 (I93097,I77106);
nor I_5300 (I92967,I93063,I93097);
not I_5301 (I93128,I93097);
nand I_5302 (I92952,I93063,I93128);
not I_5303 (I93159,I77091);
nor I_5304 (I93176,I93159,I77085);
and I_5305 (I93193,I93176,I77097);
or I_5306 (I93210,I93193,I77082);
DFFARX1 I_5307 (I93227,I93210,I2966,I92978,);
nor I_5308 (I93244,I93227,I93080);
DFFARX1 I_5309 (I93261,I93227,I2966,I92978,);
not I_5310 (I92949,I93261);
nand I_5311 (I93292,I92995,I77091);
and I_5312 (I93309,I93292,I93244);
DFFARX1 I_5313 (I92946,I93292,I2966,I92978,);
DFFARX1 I_5314 (I93340,I77079,I2966,I92978,);
nor I_5315 (I93357,I93340,I93063);
nand I_5316 (I92964,I93227,I93357);
nor I_5317 (I93388,I93340,I93128);
not I_5318 (I92961,I93340);
nand I_5319 (I93419,I93340,I93029);
and I_5320 (I93436,I93097,I93419);
DFFARX1 I_5321 (I92940,I93436,I2966,I92978,);
DFFARX1 I_5322 (I92943,I93340,I2966,I92978,);
DFFARX1 I_5323 (I93481,I77103,I2966,I92978,);
not I_5324 (I93498,I93481);
nand I_5325 (I93515,I93498,I93063);
and I_5326 (I93532,I93292,I93515);
DFFARX1 I_5327 (I92970,I93532,I2966,I92978,);
or I_5328 (I93563,I93498,I93309);
DFFARX1 I_5329 (I92955,I93563,I2966,I92978,);
nand I_5330 (I92958,I93498,I93388);
not I_5331 (I93641,I2973);
not I_5332 (I93658,I91685);
nor I_5333 (I93675,I91691,I91697);
nand I_5334 (I93692,I93675,I91700);
nor I_5335 (I93709,I93658,I91691);
nand I_5336 (I93726,I93709,I91682);
not I_5337 (I93743,I93726);
not I_5338 (I93760,I91691);
nor I_5339 (I93630,I93726,I93760);
not I_5340 (I93791,I93760);
nand I_5341 (I93615,I93726,I93791);
not I_5342 (I93822,I91694);
nor I_5343 (I93839,I93822,I91688);
and I_5344 (I93856,I93839,I91703);
or I_5345 (I93873,I93856,I91709);
DFFARX1 I_5346 (I93890,I93873,I2966,I93641,);
nor I_5347 (I93907,I93890,I93743);
DFFARX1 I_5348 (I93924,I93890,I2966,I93641,);
not I_5349 (I93612,I93924);
nand I_5350 (I93955,I93658,I91694);
and I_5351 (I93972,I93955,I93907);
DFFARX1 I_5352 (I93609,I93955,I2966,I93641,);
DFFARX1 I_5353 (I94003,I91706,I2966,I93641,);
nor I_5354 (I94020,I94003,I93726);
nand I_5355 (I93627,I93890,I94020);
nor I_5356 (I94051,I94003,I93791);
not I_5357 (I93624,I94003);
nand I_5358 (I94082,I94003,I93692);
and I_5359 (I94099,I93760,I94082);
DFFARX1 I_5360 (I93603,I94099,I2966,I93641,);
DFFARX1 I_5361 (I93606,I94003,I2966,I93641,);
DFFARX1 I_5362 (I94144,I91712,I2966,I93641,);
not I_5363 (I94161,I94144);
nand I_5364 (I94178,I94161,I93726);
and I_5365 (I94195,I93955,I94178);
DFFARX1 I_5366 (I93633,I94195,I2966,I93641,);
or I_5367 (I94226,I94161,I93972);
DFFARX1 I_5368 (I93618,I94226,I2966,I93641,);
nand I_5369 (I93621,I94161,I94051);
not I_5370 (I94304,I2973);
not I_5371 (I94321,I81823);
nor I_5372 (I94338,I81811,I81820);
nand I_5373 (I94355,I94338,I81835);
nor I_5374 (I94372,I94321,I81811);
nand I_5375 (I94389,I94372,I81817);
DFFARX1 I_5376 (I94406,I94389,I2966,I94304,);
not I_5377 (I94275,I94406);
not I_5378 (I94437,I81811);
not I_5379 (I94454,I94437);
not I_5380 (I94471,I81805);
nor I_5381 (I94488,I94471,I81826);
and I_5382 (I94505,I94488,I81808);
or I_5383 (I94522,I94505,I81814);
DFFARX1 I_5384 (I94539,I94522,I2966,I94304,);
DFFARX1 I_5385 (I94272,I94539,I2966,I94304,);
DFFARX1 I_5386 (I94570,I94539,I2966,I94304,);
DFFARX1 I_5387 (I94266,I94539,I2966,I94304,);
nand I_5388 (I94601,I94321,I81805);
nand I_5389 (I94618,I94601,I94355);
and I_5390 (I94635,I94437,I94618);
DFFARX1 I_5391 (I94296,I94635,I2966,I94304,);
and I_5392 (I94269,I94601,I94570);
DFFARX1 I_5393 (I94680,I81832,I2966,I94304,);
nor I_5394 (I94293,I94680,I94601);
nor I_5395 (I94711,I94680,I94355);
nand I_5396 (I94290,I94389,I94711);
not I_5397 (I94287,I94680);
DFFARX1 I_5398 (I94756,I81829,I2966,I94304,);
not I_5399 (I94773,I94756);
nor I_5400 (I94790,I94773,I94454);
and I_5401 (I94807,I94680,I94790);
or I_5402 (I94824,I94601,I94807);
DFFARX1 I_5403 (I94281,I94824,I2966,I94304,);
not I_5404 (I94855,I94773);
nor I_5405 (I94872,I94680,I94855);
nand I_5406 (I94284,I94773,I94872);
nand I_5407 (I94278,I94437,I94855);
not I_5408 (I94950,I2973);
not I_5409 (I94967,I82418);
nor I_5410 (I94984,I82406,I82415);
nand I_5411 (I95001,I94984,I82430);
nor I_5412 (I95018,I94967,I82406);
nand I_5413 (I95035,I95018,I82412);
DFFARX1 I_5414 (I95052,I95035,I2966,I94950,);
not I_5415 (I94921,I95052);
not I_5416 (I95083,I82406);
not I_5417 (I95100,I95083);
not I_5418 (I95117,I82400);
nor I_5419 (I95134,I95117,I82421);
and I_5420 (I95151,I95134,I82403);
or I_5421 (I95168,I95151,I82409);
DFFARX1 I_5422 (I95185,I95168,I2966,I94950,);
DFFARX1 I_5423 (I94918,I95185,I2966,I94950,);
DFFARX1 I_5424 (I95216,I95185,I2966,I94950,);
DFFARX1 I_5425 (I94912,I95185,I2966,I94950,);
nand I_5426 (I95247,I94967,I82400);
nand I_5427 (I95264,I95247,I95001);
and I_5428 (I95281,I95083,I95264);
DFFARX1 I_5429 (I94942,I95281,I2966,I94950,);
and I_5430 (I94915,I95247,I95216);
DFFARX1 I_5431 (I95326,I82427,I2966,I94950,);
nor I_5432 (I94939,I95326,I95247);
nor I_5433 (I95357,I95326,I95001);
nand I_5434 (I94936,I95035,I95357);
not I_5435 (I94933,I95326);
DFFARX1 I_5436 (I95402,I82424,I2966,I94950,);
not I_5437 (I95419,I95402);
nor I_5438 (I95436,I95419,I95100);
and I_5439 (I95453,I95326,I95436);
or I_5440 (I95470,I95247,I95453);
DFFARX1 I_5441 (I94927,I95470,I2966,I94950,);
not I_5442 (I95501,I95419);
nor I_5443 (I95518,I95326,I95501);
nand I_5444 (I94930,I95419,I95518);
nand I_5445 (I94924,I95083,I95501);
not I_5446 (I95596,I2973);
not I_5447 (I95613,I77672);
nor I_5448 (I95630,I77675,I77657);
nand I_5449 (I95647,I95630,I77684);
nor I_5450 (I95664,I95613,I77675);
nand I_5451 (I95681,I95664,I77663);
DFFARX1 I_5452 (I95698,I95681,I2966,I95596,);
not I_5453 (I95567,I95698);
not I_5454 (I95729,I77675);
not I_5455 (I95746,I95729);
not I_5456 (I95763,I77669);
nor I_5457 (I95780,I95763,I77681);
and I_5458 (I95797,I95780,I77687);
or I_5459 (I95814,I95797,I77666);
DFFARX1 I_5460 (I95831,I95814,I2966,I95596,);
DFFARX1 I_5461 (I95564,I95831,I2966,I95596,);
DFFARX1 I_5462 (I95862,I95831,I2966,I95596,);
DFFARX1 I_5463 (I95558,I95831,I2966,I95596,);
nand I_5464 (I95893,I95613,I77669);
nand I_5465 (I95910,I95893,I95647);
and I_5466 (I95927,I95729,I95910);
DFFARX1 I_5467 (I95588,I95927,I2966,I95596,);
and I_5468 (I95561,I95893,I95862);
DFFARX1 I_5469 (I95972,I77678,I2966,I95596,);
nor I_5470 (I95585,I95972,I95893);
nor I_5471 (I96003,I95972,I95647);
nand I_5472 (I95582,I95681,I96003);
not I_5473 (I95579,I95972);
DFFARX1 I_5474 (I96048,I77660,I2966,I95596,);
not I_5475 (I96065,I96048);
nor I_5476 (I96082,I96065,I95746);
and I_5477 (I96099,I95972,I96082);
or I_5478 (I96116,I95893,I96099);
DFFARX1 I_5479 (I95573,I96116,I2966,I95596,);
not I_5480 (I96147,I96065);
nor I_5481 (I96164,I95972,I96147);
nand I_5482 (I95576,I96065,I96164);
nand I_5483 (I95570,I95729,I96147);
not I_5484 (I96242,I2973);
not I_5485 (I96259,I89085);
nor I_5486 (I96276,I89076,I89067);
nand I_5487 (I96293,I96276,I89082);
nor I_5488 (I96310,I96259,I89076);
nand I_5489 (I96327,I96310,I89079);
DFFARX1 I_5490 (I96344,I96327,I2966,I96242,);
not I_5491 (I96213,I96344);
not I_5492 (I96375,I89076);
not I_5493 (I96392,I96375);
not I_5494 (I96409,I89088);
nor I_5495 (I96426,I96409,I89073);
and I_5496 (I96443,I96426,I89091);
or I_5497 (I96460,I96443,I89064);
DFFARX1 I_5498 (I96477,I96460,I2966,I96242,);
DFFARX1 I_5499 (I96210,I96477,I2966,I96242,);
DFFARX1 I_5500 (I96508,I96477,I2966,I96242,);
DFFARX1 I_5501 (I96204,I96477,I2966,I96242,);
nand I_5502 (I96539,I96259,I89088);
nand I_5503 (I96556,I96539,I96293);
and I_5504 (I96573,I96375,I96556);
DFFARX1 I_5505 (I96234,I96573,I2966,I96242,);
and I_5506 (I96207,I96539,I96508);
DFFARX1 I_5507 (I96618,I89094,I2966,I96242,);
nor I_5508 (I96231,I96618,I96539);
nor I_5509 (I96649,I96618,I96293);
nand I_5510 (I96228,I96327,I96649);
not I_5511 (I96225,I96618);
DFFARX1 I_5512 (I96694,I89070,I2966,I96242,);
not I_5513 (I96711,I96694);
nor I_5514 (I96728,I96711,I96392);
and I_5515 (I96745,I96618,I96728);
or I_5516 (I96762,I96539,I96745);
DFFARX1 I_5517 (I96219,I96762,I2966,I96242,);
not I_5518 (I96793,I96711);
nor I_5519 (I96810,I96618,I96793);
nand I_5520 (I96222,I96711,I96810);
nand I_5521 (I96216,I96375,I96793);
not I_5522 (I96888,I2973);
not I_5523 (I96905,I78839);
nor I_5524 (I96922,I78851,I78845);
nand I_5525 (I96939,I96922,I78830);
nor I_5526 (I96956,I96905,I78851);
nand I_5527 (I96973,I96956,I78857);
DFFARX1 I_5528 (I96990,I96973,I2966,I96888,);
not I_5529 (I96859,I96990);
not I_5530 (I97021,I78851);
not I_5531 (I97038,I97021);
not I_5532 (I97055,I78854);
nor I_5533 (I97072,I97055,I78836);
and I_5534 (I97089,I97072,I78833);
or I_5535 (I97106,I97089,I78860);
DFFARX1 I_5536 (I97123,I97106,I2966,I96888,);
DFFARX1 I_5537 (I96856,I97123,I2966,I96888,);
DFFARX1 I_5538 (I97154,I97123,I2966,I96888,);
DFFARX1 I_5539 (I96850,I97123,I2966,I96888,);
nand I_5540 (I97185,I96905,I78854);
nand I_5541 (I97202,I97185,I96939);
and I_5542 (I97219,I97021,I97202);
DFFARX1 I_5543 (I96880,I97219,I2966,I96888,);
and I_5544 (I96853,I97185,I97154);
DFFARX1 I_5545 (I97264,I78848,I2966,I96888,);
nor I_5546 (I96877,I97264,I97185);
nor I_5547 (I97295,I97264,I96939);
nand I_5548 (I96874,I96973,I97295);
not I_5549 (I96871,I97264);
DFFARX1 I_5550 (I97340,I78842,I2966,I96888,);
not I_5551 (I97357,I97340);
nor I_5552 (I97374,I97357,I97038);
and I_5553 (I97391,I97264,I97374);
or I_5554 (I97408,I97185,I97391);
DFFARX1 I_5555 (I96865,I97408,I2966,I96888,);
not I_5556 (I97439,I97357);
nor I_5557 (I97456,I97264,I97439);
nand I_5558 (I96868,I97357,I97456);
nand I_5559 (I96862,I97021,I97439);
not I_5560 (I97534,I2973);
nand I_5561 (I97551,I84271,I84274);
and I_5562 (I97568,I97551,I84280);
DFFARX1 I_5563 (I97585,I97568,I2966,I97534,);
not I_5564 (I97602,I97585);
DFFARX1 I_5565 (I97502,I97585,I2966,I97534,);
nor I_5566 (I97633,I84277,I84274);
DFFARX1 I_5567 (I97650,I84256,I2966,I97534,);
DFFARX1 I_5568 (I97667,I97650,I2966,I97534,);
not I_5569 (I97505,I97667);
DFFARX1 I_5570 (I97698,I97650,I2966,I97534,);
and I_5571 (I97499,I97585,I97698);
nand I_5572 (I97729,I84253,I84268);
and I_5573 (I97746,I97729,I84265);
DFFARX1 I_5574 (I97763,I97746,I2966,I97534,);
nor I_5575 (I97780,I97763,I97602);
not I_5576 (I97797,I97763);
nand I_5577 (I97508,I97585,I97797);
DFFARX1 I_5578 (I97828,I84283,I2966,I97534,);
and I_5579 (I97845,I97828,I84262);
nor I_5580 (I97862,I97845,I97763);
nor I_5581 (I97879,I97845,I97797);
nand I_5582 (I97514,I97633,I97879);
not I_5583 (I97517,I97845);
DFFARX1 I_5584 (I97496,I97845,I2966,I97534,);
DFFARX1 I_5585 (I97938,I84259,I2966,I97534,);
nand I_5586 (I97955,I97938,I97650);
and I_5587 (I97972,I97633,I97955);
DFFARX1 I_5588 (I97526,I97972,I2966,I97534,);
nor I_5589 (I97523,I97938,I97845);
and I_5590 (I98017,I97938,I97780);
or I_5591 (I98034,I97633,I98017);
DFFARX1 I_5592 (I97511,I98034,I2966,I97534,);
nand I_5593 (I97520,I97938,I97862);
not I_5594 (I98112,I2973);
nand I_5595 (I98129,I84900,I84903);
and I_5596 (I98146,I98129,I84909);
DFFARX1 I_5597 (I98163,I98146,I2966,I98112,);
not I_5598 (I98180,I98163);
DFFARX1 I_5599 (I98080,I98163,I2966,I98112,);
nor I_5600 (I98211,I84906,I84903);
DFFARX1 I_5601 (I98228,I84885,I2966,I98112,);
DFFARX1 I_5602 (I98245,I98228,I2966,I98112,);
not I_5603 (I98083,I98245);
DFFARX1 I_5604 (I98276,I98228,I2966,I98112,);
and I_5605 (I98077,I98163,I98276);
nand I_5606 (I98307,I84882,I84897);
and I_5607 (I98324,I98307,I84894);
DFFARX1 I_5608 (I98341,I98324,I2966,I98112,);
nor I_5609 (I98358,I98341,I98180);
not I_5610 (I98375,I98341);
nand I_5611 (I98086,I98163,I98375);
DFFARX1 I_5612 (I98406,I84912,I2966,I98112,);
and I_5613 (I98423,I98406,I84891);
nor I_5614 (I98440,I98423,I98341);
nor I_5615 (I98457,I98423,I98375);
nand I_5616 (I98092,I98211,I98457);
not I_5617 (I98095,I98423);
DFFARX1 I_5618 (I98074,I98423,I2966,I98112,);
DFFARX1 I_5619 (I98516,I84888,I2966,I98112,);
nand I_5620 (I98533,I98516,I98228);
and I_5621 (I98550,I98211,I98533);
DFFARX1 I_5622 (I98104,I98550,I2966,I98112,);
nor I_5623 (I98101,I98516,I98423);
and I_5624 (I98595,I98516,I98358);
or I_5625 (I98612,I98211,I98595);
DFFARX1 I_5626 (I98089,I98612,I2966,I98112,);
nand I_5627 (I98098,I98516,I98440);
not I_5628 (I98690,I2973);
or I_5629 (I98707,I90365,I90356);
or I_5630 (I98724,I90368,I90365);
nor I_5631 (I98741,I90383,I90359);
not I_5632 (I98758,I98741);
DFFARX1 I_5633 (I98658,I98741,I2966,I98690,);
nand I_5634 (I98789,I98741,I98707);
not I_5635 (I98806,I90383);
and I_5636 (I98823,I98806,I90380);
nor I_5637 (I98840,I98823,I90356);
nor I_5638 (I98857,I90377,I90362);
DFFARX1 I_5639 (I98874,I98857,I2966,I98690,);
nor I_5640 (I98891,I98874,I98758);
not I_5641 (I98908,I98874);
nand I_5642 (I98664,I98741,I98908);
DFFARX1 I_5643 (I98655,I98874,I2966,I98690,);
nor I_5644 (I98953,I90377,I90368);
nand I_5645 (I98970,I98724,I98953);
nor I_5646 (I98679,I98707,I98953);
and I_5647 (I99001,I98953,I98891);
or I_5648 (I99018,I98840,I99001);
DFFARX1 I_5649 (I98667,I99018,I2966,I98690,);
DFFARX1 I_5650 (I99049,I90386,I2966,I98690,);
and I_5651 (I99066,I99049,I90371);
not I_5652 (I98673,I99066);
DFFARX1 I_5653 (I99097,I99066,I2966,I98690,);
not I_5654 (I98661,I99097);
and I_5655 (I99128,I99066,I98789);
DFFARX1 I_5656 (I98652,I99128,I2966,I98690,);
DFFARX1 I_5657 (I99159,I90374,I2966,I98690,);
and I_5658 (I99176,I99159,I98970);
DFFARX1 I_5659 (I98682,I99176,I2966,I98690,);
nor I_5660 (I99207,I99159,I99066);
nand I_5661 (I98676,I98840,I99207);
nor I_5662 (I99238,I99159,I98908);
nand I_5663 (I98670,I98724,I99238);
not I_5664 (I99302,I2973);
or I_5665 (I99319,I81231,I81228);
or I_5666 (I99336,I81216,I81231);
nor I_5667 (I99353,I81210,I81237);
or I_5668 (I99291,I99353,I99319);
not I_5669 (I99384,I81210);
and I_5670 (I99401,I99384,I81222);
nor I_5671 (I99418,I99401,I81228);
not I_5672 (I99435,I99418);
nor I_5673 (I99452,I81213,I81234);
DFFARX1 I_5674 (I99469,I99452,I2966,I99302,);
nor I_5675 (I99486,I99469,I99418);
nand I_5676 (I99276,I99319,I99486);
nor I_5677 (I99517,I99469,I99435);
not I_5678 (I99273,I99469);
nor I_5679 (I99548,I81213,I81216);
or I_5680 (I99285,I99319,I99548);
DFFARX1 I_5681 (I99579,I81225,I2966,I99302,);
and I_5682 (I99596,I99579,I81219);
nor I_5683 (I99613,I99596,I99469);
DFFARX1 I_5684 (I99279,I99613,I2966,I99302,);
nor I_5685 (I99294,I99596,I99548);
not I_5686 (I99658,I99596);
nor I_5687 (I99675,I99336,I99658);
nand I_5688 (I99264,I99596,I99435);
DFFARX1 I_5689 (I99706,I81240,I2966,I99302,);
nor I_5690 (I99282,I99706,I99336);
not I_5691 (I99737,I99706);
and I_5692 (I99754,I99548,I99737);
nor I_5693 (I99288,I99353,I99754);
and I_5694 (I99785,I99706,I99675);
or I_5695 (I99802,I99353,I99785);
DFFARX1 I_5696 (I99267,I99802,I2966,I99302,);
nand I_5697 (I99270,I99706,I99517);
not I_5698 (I99880,I2973);
nand I_5699 (I99897,I88427,I88439);
and I_5700 (I99914,I99897,I88448);
DFFARX1 I_5701 (I99931,I99914,I2966,I99880,);
nor I_5702 (I99948,I88442,I88439);
nor I_5703 (I99965,I99948,I99931);
not I_5704 (I99863,I99948);
DFFARX1 I_5705 (I99996,I88436,I2966,I99880,);
not I_5706 (I100013,I99996);
nor I_5707 (I100030,I99948,I100013);
nand I_5708 (I99866,I99996,I99965);
DFFARX1 I_5709 (I99848,I99996,I2966,I99880,);
nand I_5710 (I100075,I88433,I88430);
and I_5711 (I100092,I100075,I88421);
DFFARX1 I_5712 (I100109,I100092,I2966,I99880,);
nor I_5713 (I99869,I100109,I99931);
nand I_5714 (I99860,I100109,I100030);
DFFARX1 I_5715 (I100154,I88445,I2966,I99880,);
and I_5716 (I100171,I100154,I88424);
DFFARX1 I_5717 (I100188,I100171,I2966,I99880,);
not I_5718 (I99851,I100188);
nand I_5719 (I100219,I100171,I100109);
and I_5720 (I100236,I99931,I100219);
DFFARX1 I_5721 (I99842,I100236,I2966,I99880,);
DFFARX1 I_5722 (I100267,I88418,I2966,I99880,);
nand I_5723 (I100284,I100267,I99931);
and I_5724 (I100301,I100109,I100284);
DFFARX1 I_5725 (I99872,I100301,I2966,I99880,);
not I_5726 (I100332,I100267);
nor I_5727 (I100349,I99948,I100332);
and I_5728 (I100366,I100267,I100349);
or I_5729 (I100383,I100171,I100366);
DFFARX1 I_5730 (I99857,I100383,I2966,I99880,);
nand I_5731 (I99854,I100267,I100013);
DFFARX1 I_5732 (I99845,I100267,I2966,I99880,);
not I_5733 (I100475,I2973);
nand I_5734 (I100492,I89719,I89731);
and I_5735 (I100509,I100492,I89740);
DFFARX1 I_5736 (I100526,I100509,I2966,I100475,);
nor I_5737 (I100543,I89734,I89731);
nor I_5738 (I100560,I100543,I100526);
not I_5739 (I100458,I100543);
DFFARX1 I_5740 (I100591,I89728,I2966,I100475,);
not I_5741 (I100608,I100591);
nor I_5742 (I100625,I100543,I100608);
nand I_5743 (I100461,I100591,I100560);
DFFARX1 I_5744 (I100443,I100591,I2966,I100475,);
nand I_5745 (I100670,I89725,I89722);
and I_5746 (I100687,I100670,I89713);
DFFARX1 I_5747 (I100704,I100687,I2966,I100475,);
nor I_5748 (I100464,I100704,I100526);
nand I_5749 (I100455,I100704,I100625);
DFFARX1 I_5750 (I100749,I89737,I2966,I100475,);
and I_5751 (I100766,I100749,I89716);
DFFARX1 I_5752 (I100783,I100766,I2966,I100475,);
not I_5753 (I100446,I100783);
nand I_5754 (I100814,I100766,I100704);
and I_5755 (I100831,I100526,I100814);
DFFARX1 I_5756 (I100437,I100831,I2966,I100475,);
DFFARX1 I_5757 (I100862,I89710,I2966,I100475,);
nand I_5758 (I100879,I100862,I100526);
and I_5759 (I100896,I100704,I100879);
DFFARX1 I_5760 (I100467,I100896,I2966,I100475,);
not I_5761 (I100927,I100862);
nor I_5762 (I100944,I100543,I100927);
and I_5763 (I100961,I100862,I100944);
or I_5764 (I100978,I100766,I100961);
DFFARX1 I_5765 (I100452,I100978,I2966,I100475,);
nand I_5766 (I100449,I100862,I100608);
DFFARX1 I_5767 (I100440,I100862,I2966,I100475,);
not I_5768 (I101070,I2973);
nand I_5769 (I101087,I85523,I85529);
and I_5770 (I101104,I101087,I85520);
DFFARX1 I_5771 (I101121,I101104,I2966,I101070,);
nor I_5772 (I101138,I85532,I85529);
nor I_5773 (I101155,I101138,I101121);
not I_5774 (I101053,I101138);
DFFARX1 I_5775 (I101186,I85511,I2966,I101070,);
not I_5776 (I101203,I101186);
nor I_5777 (I101220,I101138,I101203);
nand I_5778 (I101056,I101186,I101155);
DFFARX1 I_5779 (I101038,I101186,I2966,I101070,);
nand I_5780 (I101265,I85535,I85517);
and I_5781 (I101282,I101265,I85526);
DFFARX1 I_5782 (I101299,I101282,I2966,I101070,);
nor I_5783 (I101059,I101299,I101121);
nand I_5784 (I101050,I101299,I101220);
DFFARX1 I_5785 (I101344,I85541,I2966,I101070,);
and I_5786 (I101361,I101344,I85514);
DFFARX1 I_5787 (I101378,I101361,I2966,I101070,);
not I_5788 (I101041,I101378);
nand I_5789 (I101409,I101361,I101299);
and I_5790 (I101426,I101121,I101409);
DFFARX1 I_5791 (I101032,I101426,I2966,I101070,);
DFFARX1 I_5792 (I101457,I85538,I2966,I101070,);
nand I_5793 (I101474,I101457,I101121);
and I_5794 (I101491,I101299,I101474);
DFFARX1 I_5795 (I101062,I101491,I2966,I101070,);
not I_5796 (I101522,I101457);
nor I_5797 (I101539,I101138,I101522);
and I_5798 (I101556,I101457,I101539);
or I_5799 (I101573,I101361,I101556);
DFFARX1 I_5800 (I101047,I101573,I2966,I101070,);
nand I_5801 (I101044,I101457,I101203);
DFFARX1 I_5802 (I101035,I101457,I2966,I101070,);
not I_5803 (I101665,I2973);
nand I_5804 (I101682,I93621,I93627);
and I_5805 (I101699,I101682,I93609);
DFFARX1 I_5806 (I101716,I101699,I2966,I101665,);
nor I_5807 (I101733,I93603,I93627);
nor I_5808 (I101750,I101733,I101716);
not I_5809 (I101648,I101733);
DFFARX1 I_5810 (I101781,I93633,I2966,I101665,);
not I_5811 (I101798,I101781);
nor I_5812 (I101815,I101733,I101798);
nand I_5813 (I101651,I101781,I101750);
DFFARX1 I_5814 (I101633,I101781,I2966,I101665,);
nand I_5815 (I101860,I93624,I93615);
and I_5816 (I101877,I101860,I93618);
DFFARX1 I_5817 (I101894,I101877,I2966,I101665,);
nor I_5818 (I101654,I101894,I101716);
nand I_5819 (I101645,I101894,I101815);
DFFARX1 I_5820 (I101939,I93630,I2966,I101665,);
and I_5821 (I101956,I101939,I93606);
DFFARX1 I_5822 (I101973,I101956,I2966,I101665,);
not I_5823 (I101636,I101973);
nand I_5824 (I102004,I101956,I101894);
and I_5825 (I102021,I101716,I102004);
DFFARX1 I_5826 (I101627,I102021,I2966,I101665,);
DFFARX1 I_5827 (I102052,I93612,I2966,I101665,);
nand I_5828 (I102069,I102052,I101716);
and I_5829 (I102086,I101894,I102069);
DFFARX1 I_5830 (I101657,I102086,I2966,I101665,);
not I_5831 (I102117,I102052);
nor I_5832 (I102134,I101733,I102117);
and I_5833 (I102151,I102052,I102134);
or I_5834 (I102168,I101956,I102151);
DFFARX1 I_5835 (I101642,I102168,I2966,I101665,);
nand I_5836 (I101639,I102052,I101798);
DFFARX1 I_5837 (I101630,I102052,I2966,I101665,);
not I_5838 (I102260,I2973);
nand I_5839 (I102277,I87781,I87793);
and I_5840 (I102294,I102277,I87802);
DFFARX1 I_5841 (I102311,I102294,I2966,I102260,);
nor I_5842 (I102328,I87796,I87793);
nor I_5843 (I102345,I102328,I102311);
not I_5844 (I102243,I102328);
DFFARX1 I_5845 (I102376,I87790,I2966,I102260,);
not I_5846 (I102393,I102376);
nor I_5847 (I102410,I102328,I102393);
nand I_5848 (I102246,I102376,I102345);
DFFARX1 I_5849 (I102228,I102376,I2966,I102260,);
nand I_5850 (I102455,I87787,I87784);
and I_5851 (I102472,I102455,I87775);
DFFARX1 I_5852 (I102489,I102472,I2966,I102260,);
nor I_5853 (I102249,I102489,I102311);
nand I_5854 (I102240,I102489,I102410);
DFFARX1 I_5855 (I102534,I87799,I2966,I102260,);
and I_5856 (I102551,I102534,I87778);
DFFARX1 I_5857 (I102568,I102551,I2966,I102260,);
not I_5858 (I102231,I102568);
nand I_5859 (I102599,I102551,I102489);
and I_5860 (I102616,I102311,I102599);
DFFARX1 I_5861 (I102222,I102616,I2966,I102260,);
DFFARX1 I_5862 (I102647,I87772,I2966,I102260,);
nand I_5863 (I102664,I102647,I102311);
and I_5864 (I102681,I102489,I102664);
DFFARX1 I_5865 (I102252,I102681,I2966,I102260,);
not I_5866 (I102712,I102647);
nor I_5867 (I102729,I102328,I102712);
and I_5868 (I102746,I102647,I102729);
or I_5869 (I102763,I102551,I102746);
DFFARX1 I_5870 (I102237,I102763,I2966,I102260,);
nand I_5871 (I102234,I102647,I102393);
DFFARX1 I_5872 (I102225,I102647,I2966,I102260,);
not I_5873 (I102855,I2973);
nand I_5874 (I102872,I87214,I87229);
and I_5875 (I102889,I102872,I87235);
DFFARX1 I_5876 (I102906,I102889,I2966,I102855,);
nor I_5877 (I102923,I87223,I87229);
DFFARX1 I_5878 (I102940,I87211,I2966,I102855,);
nand I_5879 (I102957,I102940,I102923);
DFFARX1 I_5880 (I102826,I102940,I2966,I102855,);
nand I_5881 (I102988,I87217,I87220);
and I_5882 (I103005,I102988,I87226);
DFFARX1 I_5883 (I103022,I103005,I2966,I102855,);
not I_5884 (I103039,I103022);
nor I_5885 (I103056,I102906,I103039);
and I_5886 (I103073,I102923,I103056);
and I_5887 (I103090,I103022,I102957);
DFFARX1 I_5888 (I102823,I103090,I2966,I102855,);
DFFARX1 I_5889 (I102817,I103022,I2966,I102855,);
DFFARX1 I_5890 (I103135,I87232,I2966,I102855,);
and I_5891 (I103152,I103135,I87241);
nand I_5892 (I103169,I103152,I103022);
nor I_5893 (I102844,I103152,I102923);
not I_5894 (I103200,I103152);
nor I_5895 (I103217,I102906,I103200);
nand I_5896 (I102835,I102940,I103217);
nand I_5897 (I102829,I103022,I103200);
or I_5898 (I103262,I103152,I103073);
DFFARX1 I_5899 (I102832,I103262,I2966,I102855,);
DFFARX1 I_5900 (I103293,I87238,I2966,I102855,);
and I_5901 (I103310,I103293,I103169);
DFFARX1 I_5902 (I102847,I103310,I2966,I102855,);
nor I_5903 (I103341,I103293,I102906);
nand I_5904 (I102841,I103152,I103341);
not I_5905 (I102838,I103293);
DFFARX1 I_5906 (I103386,I103293,I2966,I102855,);
and I_5907 (I102820,I103293,I103386);
not I_5908 (I103450,I2973);
nand I_5909 (I103467,I97508,I97523);
and I_5910 (I103484,I103467,I97520);
DFFARX1 I_5911 (I103501,I103484,I2966,I103450,);
nor I_5912 (I103518,I97496,I97523);
DFFARX1 I_5913 (I103535,I97514,I2966,I103450,);
nand I_5914 (I103552,I103535,I103518);
DFFARX1 I_5915 (I103421,I103535,I2966,I103450,);
nand I_5916 (I103583,I97517,I97505);
and I_5917 (I103600,I103583,I97511);
DFFARX1 I_5918 (I103617,I103600,I2966,I103450,);
not I_5919 (I103634,I103617);
nor I_5920 (I103651,I103501,I103634);
and I_5921 (I103668,I103518,I103651);
and I_5922 (I103685,I103617,I103552);
DFFARX1 I_5923 (I103418,I103685,I2966,I103450,);
DFFARX1 I_5924 (I103412,I103617,I2966,I103450,);
DFFARX1 I_5925 (I103730,I97502,I2966,I103450,);
and I_5926 (I103747,I103730,I97526);
nand I_5927 (I103764,I103747,I103617);
nor I_5928 (I103439,I103747,I103518);
not I_5929 (I103795,I103747);
nor I_5930 (I103812,I103501,I103795);
nand I_5931 (I103430,I103535,I103812);
nand I_5932 (I103424,I103617,I103795);
or I_5933 (I103857,I103747,I103668);
DFFARX1 I_5934 (I103427,I103857,I2966,I103450,);
DFFARX1 I_5935 (I103888,I97499,I2966,I103450,);
and I_5936 (I103905,I103888,I103764);
DFFARX1 I_5937 (I103442,I103905,I2966,I103450,);
nor I_5938 (I103936,I103888,I103501);
nand I_5939 (I103436,I103747,I103936);
not I_5940 (I103433,I103888);
DFFARX1 I_5941 (I103981,I103888,I2966,I103450,);
and I_5942 (I103415,I103888,I103981);
not I_5943 (I104045,I2973);
not I_5944 (I104062,I102228);
nor I_5945 (I104079,I102246,I102225);
nand I_5946 (I104096,I104079,I102249);
nor I_5947 (I104113,I104062,I102246);
nand I_5948 (I104130,I104113,I102243);
not I_5949 (I104147,I102246);
not I_5950 (I104164,I104147);
not I_5951 (I104181,I102234);
nor I_5952 (I104198,I104181,I102222);
and I_5953 (I104215,I104198,I102240);
or I_5954 (I104232,I104215,I102252);
DFFARX1 I_5955 (I104249,I104232,I2966,I104045,);
nand I_5956 (I104266,I104062,I102234);
or I_5957 (I104034,I104266,I104249);
not I_5958 (I104297,I104266);
nor I_5959 (I104314,I104249,I104297);
and I_5960 (I104331,I104147,I104314);
nand I_5961 (I104007,I104266,I104164);
DFFARX1 I_5962 (I104362,I102231,I2966,I104045,);
or I_5963 (I104028,I104362,I104249);
nor I_5964 (I104393,I104362,I104130);
nor I_5965 (I104410,I104362,I104164);
nand I_5966 (I104013,I104096,I104410);
or I_5967 (I104441,I104362,I104331);
DFFARX1 I_5968 (I104010,I104441,I2966,I104045,);
not I_5969 (I104016,I104362);
DFFARX1 I_5970 (I104486,I102237,I2966,I104045,);
not I_5971 (I104503,I104486);
nor I_5972 (I104520,I104503,I104096);
DFFARX1 I_5973 (I104022,I104520,I2966,I104045,);
nor I_5974 (I104037,I104362,I104503);
nor I_5975 (I104025,I104503,I104266);
not I_5976 (I104579,I104503);
and I_5977 (I104596,I104130,I104579);
nor I_5978 (I104031,I104266,I104596);
nand I_5979 (I104019,I104503,I104393);
not I_5980 (I104674,I2973);
not I_5981 (I104691,I92958);
nor I_5982 (I104708,I92964,I92943);
nand I_5983 (I104725,I104708,I92949);
nor I_5984 (I104742,I104691,I92964);
nand I_5985 (I104759,I104742,I92955);
not I_5986 (I104776,I92964);
not I_5987 (I104793,I104776);
not I_5988 (I104810,I92952);
nor I_5989 (I104827,I104810,I92970);
and I_5990 (I104844,I104827,I92961);
or I_5991 (I104861,I104844,I92940);
DFFARX1 I_5992 (I104878,I104861,I2966,I104674,);
nand I_5993 (I104895,I104691,I92952);
or I_5994 (I104663,I104895,I104878);
not I_5995 (I104926,I104895);
nor I_5996 (I104943,I104878,I104926);
and I_5997 (I104960,I104776,I104943);
nand I_5998 (I104636,I104895,I104793);
DFFARX1 I_5999 (I104991,I92967,I2966,I104674,);
or I_6000 (I104657,I104991,I104878);
nor I_6001 (I105022,I104991,I104759);
nor I_6002 (I105039,I104991,I104793);
nand I_6003 (I104642,I104725,I105039);
or I_6004 (I105070,I104991,I104960);
DFFARX1 I_6005 (I104639,I105070,I2966,I104674,);
not I_6006 (I104645,I104991);
DFFARX1 I_6007 (I105115,I92946,I2966,I104674,);
not I_6008 (I105132,I105115);
nor I_6009 (I105149,I105132,I104725);
DFFARX1 I_6010 (I104651,I105149,I2966,I104674,);
nor I_6011 (I104666,I104991,I105132);
nor I_6012 (I104654,I105132,I104895);
not I_6013 (I105208,I105132);
and I_6014 (I105225,I104759,I105208);
nor I_6015 (I104660,I104895,I105225);
nand I_6016 (I104648,I105132,I105022);
not I_6017 (I105303,I2973);
not I_6018 (I105320,I92375);
nor I_6019 (I105337,I92351,I92366);
nand I_6020 (I105354,I105337,I92348);
nor I_6021 (I105371,I105320,I92351);
nand I_6022 (I105388,I105371,I92363);
not I_6023 (I105405,I92351);
not I_6024 (I105422,I105405);
not I_6025 (I105439,I92354);
nor I_6026 (I105456,I105439,I92369);
and I_6027 (I105473,I105456,I92360);
or I_6028 (I105490,I105473,I92345);
DFFARX1 I_6029 (I105507,I105490,I2966,I105303,);
nand I_6030 (I105524,I105320,I92354);
or I_6031 (I105292,I105524,I105507);
not I_6032 (I105555,I105524);
nor I_6033 (I105572,I105507,I105555);
and I_6034 (I105589,I105405,I105572);
nand I_6035 (I105265,I105524,I105422);
DFFARX1 I_6036 (I105620,I92357,I2966,I105303,);
or I_6037 (I105286,I105620,I105507);
nor I_6038 (I105651,I105620,I105388);
nor I_6039 (I105668,I105620,I105422);
nand I_6040 (I105271,I105354,I105668);
or I_6041 (I105699,I105620,I105589);
DFFARX1 I_6042 (I105268,I105699,I2966,I105303,);
not I_6043 (I105274,I105620);
DFFARX1 I_6044 (I105744,I92372,I2966,I105303,);
not I_6045 (I105761,I105744);
nor I_6046 (I105778,I105761,I105354);
DFFARX1 I_6047 (I105280,I105778,I2966,I105303,);
nor I_6048 (I105295,I105620,I105761);
nor I_6049 (I105283,I105761,I105524);
not I_6050 (I105837,I105761);
and I_6051 (I105854,I105388,I105837);
nor I_6052 (I105289,I105524,I105854);
nand I_6053 (I105277,I105761,I105651);
not I_6054 (I105932,I2973);
not I_6055 (I105949,I102826);
nor I_6056 (I105966,I102829,I102838);
nand I_6057 (I105983,I105966,I102823);
nor I_6058 (I106000,I105949,I102829);
nand I_6059 (I106017,I106000,I102832);
not I_6060 (I106034,I102829);
not I_6061 (I106051,I106034);
not I_6062 (I106068,I102847);
nor I_6063 (I106085,I106068,I102835);
and I_6064 (I106102,I106085,I102820);
or I_6065 (I106119,I106102,I102817);
DFFARX1 I_6066 (I106136,I106119,I2966,I105932,);
nand I_6067 (I106153,I105949,I102847);
or I_6068 (I105921,I106153,I106136);
not I_6069 (I106184,I106153);
nor I_6070 (I106201,I106136,I106184);
and I_6071 (I106218,I106034,I106201);
nand I_6072 (I105894,I106153,I106051);
DFFARX1 I_6073 (I106249,I102841,I2966,I105932,);
or I_6074 (I105915,I106249,I106136);
nor I_6075 (I106280,I106249,I106017);
nor I_6076 (I106297,I106249,I106051);
nand I_6077 (I105900,I105983,I106297);
or I_6078 (I106328,I106249,I106218);
DFFARX1 I_6079 (I105897,I106328,I2966,I105932,);
not I_6080 (I105903,I106249);
DFFARX1 I_6081 (I106373,I102844,I2966,I105932,);
not I_6082 (I106390,I106373);
nor I_6083 (I106407,I106390,I105983);
DFFARX1 I_6084 (I105909,I106407,I2966,I105932,);
nor I_6085 (I105924,I106249,I106390);
nor I_6086 (I105912,I106390,I106153);
not I_6087 (I106466,I106390);
and I_6088 (I106483,I106017,I106466);
nor I_6089 (I105918,I106153,I106483);
nand I_6090 (I105906,I106390,I106280);
not I_6091 (I106561,I2973);
nand I_6092 (I106578,I86113,I86098);
and I_6093 (I106595,I106578,I86107);
DFFARX1 I_6094 (I106612,I106595,I2966,I106561,);
not I_6095 (I106550,I106612);
DFFARX1 I_6096 (I106643,I106612,I2966,I106561,);
not I_6097 (I106538,I106643);
nor I_6098 (I106674,I86119,I86098);
not I_6099 (I106691,I106674);
nor I_6100 (I106708,I106612,I106691);
DFFARX1 I_6101 (I106725,I86110,I2966,I106561,);
not I_6102 (I106742,I106725);
nand I_6103 (I106541,I106725,I106691);
DFFARX1 I_6104 (I106773,I106725,I2966,I106561,);
and I_6105 (I106526,I106612,I106773);
nand I_6106 (I106804,I86095,I86089);
and I_6107 (I106821,I106804,I86104);
DFFARX1 I_6108 (I106838,I106821,I2966,I106561,);
nor I_6109 (I106855,I106838,I106742);
and I_6110 (I106872,I106674,I106855);
nor I_6111 (I106889,I106838,I106612);
DFFARX1 I_6112 (I106532,I106838,I2966,I106561,);
DFFARX1 I_6113 (I106920,I86092,I2966,I106561,);
and I_6114 (I106937,I106920,I86116);
or I_6115 (I106954,I106937,I106872);
DFFARX1 I_6116 (I106544,I106954,I2966,I106561,);
nand I_6117 (I106553,I106937,I106889);
DFFARX1 I_6118 (I106523,I106937,I2966,I106561,);
DFFARX1 I_6119 (I107013,I86101,I2966,I106561,);
nand I_6120 (I106547,I107013,I106708);
DFFARX1 I_6121 (I106535,I107013,I2966,I106561,);
nand I_6122 (I107058,I107013,I106674);
and I_6123 (I107075,I106725,I107058);
DFFARX1 I_6124 (I106529,I107075,I2966,I106561,);
not I_6125 (I107139,I2973);
nand I_6126 (I107156,I86674,I86659);
and I_6127 (I107173,I107156,I86668);
DFFARX1 I_6128 (I107190,I107173,I2966,I107139,);
not I_6129 (I107128,I107190);
DFFARX1 I_6130 (I107221,I107190,I2966,I107139,);
not I_6131 (I107116,I107221);
nor I_6132 (I107252,I86680,I86659);
not I_6133 (I107269,I107252);
nor I_6134 (I107286,I107190,I107269);
DFFARX1 I_6135 (I107303,I86671,I2966,I107139,);
not I_6136 (I107320,I107303);
nand I_6137 (I107119,I107303,I107269);
DFFARX1 I_6138 (I107351,I107303,I2966,I107139,);
and I_6139 (I107104,I107190,I107351);
nand I_6140 (I107382,I86656,I86650);
and I_6141 (I107399,I107382,I86665);
DFFARX1 I_6142 (I107416,I107399,I2966,I107139,);
nor I_6143 (I107433,I107416,I107320);
and I_6144 (I107450,I107252,I107433);
nor I_6145 (I107467,I107416,I107190);
DFFARX1 I_6146 (I107110,I107416,I2966,I107139,);
DFFARX1 I_6147 (I107498,I86653,I2966,I107139,);
and I_6148 (I107515,I107498,I86677);
or I_6149 (I107532,I107515,I107450);
DFFARX1 I_6150 (I107122,I107532,I2966,I107139,);
nand I_6151 (I107131,I107515,I107467);
DFFARX1 I_6152 (I107101,I107515,I2966,I107139,);
DFFARX1 I_6153 (I107591,I86662,I2966,I107139,);
nand I_6154 (I107125,I107591,I107286);
DFFARX1 I_6155 (I107113,I107591,I2966,I107139,);
nand I_6156 (I107636,I107591,I107252);
and I_6157 (I107653,I107303,I107636);
DFFARX1 I_6158 (I107107,I107653,I2966,I107139,);
not I_6159 (I107717,I2973);
nand I_6160 (I107734,I104639,I104657);
and I_6161 (I107751,I107734,I104654);
DFFARX1 I_6162 (I107768,I107751,I2966,I107717,);
not I_6163 (I107706,I107768);
DFFARX1 I_6164 (I107799,I107768,I2966,I107717,);
not I_6165 (I107694,I107799);
nor I_6166 (I107830,I104660,I104657);
not I_6167 (I107847,I107830);
nor I_6168 (I107864,I107768,I107847);
DFFARX1 I_6169 (I107881,I104663,I2966,I107717,);
not I_6170 (I107898,I107881);
nand I_6171 (I107697,I107881,I107847);
DFFARX1 I_6172 (I107929,I107881,I2966,I107717,);
and I_6173 (I107682,I107768,I107929);
nand I_6174 (I107960,I104648,I104642);
and I_6175 (I107977,I107960,I104645);
DFFARX1 I_6176 (I107994,I107977,I2966,I107717,);
nor I_6177 (I108011,I107994,I107898);
and I_6178 (I108028,I107830,I108011);
nor I_6179 (I108045,I107994,I107768);
DFFARX1 I_6180 (I107688,I107994,I2966,I107717,);
DFFARX1 I_6181 (I108076,I104651,I2966,I107717,);
and I_6182 (I108093,I108076,I104636);
or I_6183 (I108110,I108093,I108028);
DFFARX1 I_6184 (I107700,I108110,I2966,I107717,);
nand I_6185 (I107709,I108093,I108045);
DFFARX1 I_6186 (I107679,I108093,I2966,I107717,);
DFFARX1 I_6187 (I108169,I104666,I2966,I107717,);
nand I_6188 (I107703,I108169,I107864);
DFFARX1 I_6189 (I107691,I108169,I2966,I107717,);
nand I_6190 (I108214,I108169,I107830);
and I_6191 (I108231,I107881,I108214);
DFFARX1 I_6192 (I107685,I108231,I2966,I107717,);
not I_6193 (I108295,I2973);
nand I_6194 (I108312,I91028,I91025);
and I_6195 (I108329,I108312,I91022);
DFFARX1 I_6196 (I108346,I108329,I2966,I108295,);
not I_6197 (I108363,I108346);
nor I_6198 (I108380,I91046,I91025);
or I_6199 (I108278,I108380,I108346);
not I_6200 (I108266,I108380);
DFFARX1 I_6201 (I108425,I91040,I2966,I108295,);
nor I_6202 (I108442,I108425,I108380);
nand I_6203 (I108459,I91019,I91031);
and I_6204 (I108476,I108459,I91034);
DFFARX1 I_6205 (I108493,I108476,I2966,I108295,);
nor I_6206 (I108275,I108493,I108346);
not I_6207 (I108524,I108493);
nor I_6208 (I108541,I108425,I108524);
DFFARX1 I_6209 (I108558,I91043,I2966,I108295,);
and I_6210 (I108575,I108558,I91049);
or I_6211 (I108284,I108575,I108380);
nand I_6212 (I108263,I108575,I108541);
DFFARX1 I_6213 (I108620,I91037,I2966,I108295,);
and I_6214 (I108637,I108620,I108363);
nor I_6215 (I108281,I108575,I108637);
nor I_6216 (I108668,I108620,I108425);
DFFARX1 I_6217 (I108272,I108668,I2966,I108295,);
nor I_6218 (I108287,I108620,I108346);
not I_6219 (I108713,I108620);
nor I_6220 (I108730,I108493,I108713);
and I_6221 (I108747,I108380,I108730);
or I_6222 (I108764,I108575,I108747);
DFFARX1 I_6223 (I108260,I108764,I2966,I108295,);
nand I_6224 (I108269,I108620,I108442);
nand I_6225 (I108257,I108620,I108524);
not I_6226 (I108856,I2973);
not I_6227 (I108873,I95576);
nor I_6228 (I108890,I95588,I95570);
nand I_6229 (I108907,I108890,I95585);
DFFARX1 I_6230 (I108830,I108907,I2966,I108856,);
nor I_6231 (I108938,I108873,I95588);
nand I_6232 (I108955,I108938,I95573);
not I_6233 (I108845,I108955);
DFFARX1 I_6234 (I108827,I108955,I2966,I108856,);
not I_6235 (I109000,I95588);
not I_6236 (I109017,I109000);
not I_6237 (I109034,I95582);
nor I_6238 (I109051,I109034,I95561);
and I_6239 (I109068,I109051,I95564);
or I_6240 (I109085,I109068,I95567);
DFFARX1 I_6241 (I109102,I109085,I2966,I108856,);
nor I_6242 (I109119,I109102,I108955);
nor I_6243 (I109136,I109102,I109017);
nand I_6244 (I108842,I108907,I109136);
nand I_6245 (I109167,I108873,I95582);
nand I_6246 (I109184,I109167,I109102);
and I_6247 (I109201,I109167,I109184);
DFFARX1 I_6248 (I108824,I109201,I2966,I108856,);
DFFARX1 I_6249 (I109232,I109167,I2966,I108856,);
and I_6250 (I108821,I109000,I109232);
DFFARX1 I_6251 (I109263,I95558,I2966,I108856,);
not I_6252 (I109280,I109263);
nor I_6253 (I109297,I108955,I109280);
and I_6254 (I109314,I109263,I109297);
nand I_6255 (I108836,I109263,I109017);
DFFARX1 I_6256 (I109345,I109263,I2966,I108856,);
not I_6257 (I108833,I109345);
DFFARX1 I_6258 (I109376,I95579,I2966,I108856,);
not I_6259 (I109393,I109376);
or I_6260 (I109410,I109393,I109314);
DFFARX1 I_6261 (I108839,I109410,I2966,I108856,);
nand I_6262 (I108848,I109393,I109119);
DFFARX1 I_6263 (I108818,I109393,I2966,I108856,);
not I_6264 (I109502,I2973);
not I_6265 (I109519,I98676);
nor I_6266 (I109536,I98658,I98667);
nand I_6267 (I109553,I109536,I98679);
DFFARX1 I_6268 (I109476,I109553,I2966,I109502,);
nor I_6269 (I109584,I109519,I98658);
nand I_6270 (I109601,I109584,I98664);
not I_6271 (I109491,I109601);
DFFARX1 I_6272 (I109473,I109601,I2966,I109502,);
not I_6273 (I109646,I98658);
not I_6274 (I109663,I109646);
not I_6275 (I109680,I98655);
nor I_6276 (I109697,I109680,I98673);
and I_6277 (I109714,I109697,I98661);
or I_6278 (I109731,I109714,I98682);
DFFARX1 I_6279 (I109748,I109731,I2966,I109502,);
nor I_6280 (I109765,I109748,I109601);
nor I_6281 (I109782,I109748,I109663);
nand I_6282 (I109488,I109553,I109782);
nand I_6283 (I109813,I109519,I98655);
nand I_6284 (I109830,I109813,I109748);
and I_6285 (I109847,I109813,I109830);
DFFARX1 I_6286 (I109470,I109847,I2966,I109502,);
DFFARX1 I_6287 (I109878,I109813,I2966,I109502,);
and I_6288 (I109467,I109646,I109878);
DFFARX1 I_6289 (I109909,I98670,I2966,I109502,);
not I_6290 (I109926,I109909);
nor I_6291 (I109943,I109601,I109926);
and I_6292 (I109960,I109909,I109943);
nand I_6293 (I109482,I109909,I109663);
DFFARX1 I_6294 (I109991,I109909,I2966,I109502,);
not I_6295 (I109479,I109991);
DFFARX1 I_6296 (I110022,I98652,I2966,I109502,);
not I_6297 (I110039,I110022);
or I_6298 (I110056,I110039,I109960);
DFFARX1 I_6299 (I109485,I110056,I2966,I109502,);
nand I_6300 (I109494,I110039,I109765);
DFFARX1 I_6301 (I109464,I110039,I2966,I109502,);
not I_6302 (I110148,I2973);
not I_6303 (I110165,I101059);
nor I_6304 (I110182,I101035,I101041);
nand I_6305 (I110199,I110182,I101044);
DFFARX1 I_6306 (I110122,I110199,I2966,I110148,);
nor I_6307 (I110230,I110165,I101035);
nand I_6308 (I110247,I110230,I101053);
not I_6309 (I110137,I110247);
DFFARX1 I_6310 (I110119,I110247,I2966,I110148,);
not I_6311 (I110292,I101035);
not I_6312 (I110309,I110292);
not I_6313 (I110326,I101032);
nor I_6314 (I110343,I110326,I101047);
and I_6315 (I110360,I110343,I101038);
or I_6316 (I110377,I110360,I101050);
DFFARX1 I_6317 (I110394,I110377,I2966,I110148,);
nor I_6318 (I110411,I110394,I110247);
nor I_6319 (I110428,I110394,I110309);
nand I_6320 (I110134,I110199,I110428);
nand I_6321 (I110459,I110165,I101032);
nand I_6322 (I110476,I110459,I110394);
and I_6323 (I110493,I110459,I110476);
DFFARX1 I_6324 (I110116,I110493,I2966,I110148,);
DFFARX1 I_6325 (I110524,I110459,I2966,I110148,);
and I_6326 (I110113,I110292,I110524);
DFFARX1 I_6327 (I110555,I101062,I2966,I110148,);
not I_6328 (I110572,I110555);
nor I_6329 (I110589,I110247,I110572);
and I_6330 (I110606,I110555,I110589);
nand I_6331 (I110128,I110555,I110309);
DFFARX1 I_6332 (I110637,I110555,I2966,I110148,);
not I_6333 (I110125,I110637);
DFFARX1 I_6334 (I110668,I101056,I2966,I110148,);
not I_6335 (I110685,I110668);
or I_6336 (I110702,I110685,I110606);
DFFARX1 I_6337 (I110131,I110702,I2966,I110148,);
nand I_6338 (I110140,I110685,I110411);
DFFARX1 I_6339 (I110110,I110685,I2966,I110148,);
not I_6340 (I110794,I2973);
not I_6341 (I110811,I99857);
nor I_6342 (I110828,I99869,I99872);
nand I_6343 (I110845,I110828,I99860);
DFFARX1 I_6344 (I110765,I110845,I2966,I110794,);
nor I_6345 (I110876,I110811,I99869);
nand I_6346 (I110893,I110876,I99845);
nand I_6347 (I110910,I110893,I110845);
not I_6348 (I110927,I99869);
not I_6349 (I110944,I99848);
nor I_6350 (I110961,I110944,I99851);
and I_6351 (I110978,I110961,I99854);
or I_6352 (I110995,I110978,I99863);
DFFARX1 I_6353 (I111012,I110995,I2966,I110794,);
nor I_6354 (I111029,I111012,I110893);
nand I_6355 (I110780,I110927,I111029);
not I_6356 (I110777,I111012);
and I_6357 (I111074,I111012,I110910);
DFFARX1 I_6358 (I110762,I111074,I2966,I110794,);
DFFARX1 I_6359 (I111105,I111012,I2966,I110794,);
and I_6360 (I110759,I110927,I111105);
nand I_6361 (I111136,I110811,I99848);
not I_6362 (I111153,I111136);
nor I_6363 (I111170,I111012,I111153);
DFFARX1 I_6364 (I111187,I99866,I2966,I110794,);
nand I_6365 (I111204,I111187,I111136);
and I_6366 (I111221,I110927,I111204);
DFFARX1 I_6367 (I110786,I111221,I2966,I110794,);
not I_6368 (I111252,I111187);
nand I_6369 (I110774,I111187,I111170);
nand I_6370 (I110768,I111187,I111153);
DFFARX1 I_6371 (I111297,I99842,I2966,I110794,);
not I_6372 (I111314,I111297);
nor I_6373 (I110783,I111187,I111314);
nor I_6374 (I111345,I111314,I111252);
and I_6375 (I111362,I110893,I111345);
or I_6376 (I111379,I111136,I111362);
DFFARX1 I_6377 (I110771,I111379,I2966,I110794,);
DFFARX1 I_6378 (I110756,I111314,I2966,I110794,);
not I_6379 (I111457,I2973);
not I_6380 (I111474,I107703);
nor I_6381 (I111491,I107682,I107694);
nand I_6382 (I111508,I111491,I107688);
DFFARX1 I_6383 (I111428,I111508,I2966,I111457,);
nor I_6384 (I111539,I111474,I107682);
nand I_6385 (I111556,I111539,I107709);
nand I_6386 (I111573,I111556,I111508);
not I_6387 (I111590,I107682);
not I_6388 (I111607,I107685);
nor I_6389 (I111624,I111607,I107697);
and I_6390 (I111641,I111624,I107700);
or I_6391 (I111658,I111641,I107706);
DFFARX1 I_6392 (I111675,I111658,I2966,I111457,);
nor I_6393 (I111692,I111675,I111556);
nand I_6394 (I111443,I111590,I111692);
not I_6395 (I111440,I111675);
and I_6396 (I111737,I111675,I111573);
DFFARX1 I_6397 (I111425,I111737,I2966,I111457,);
DFFARX1 I_6398 (I111768,I111675,I2966,I111457,);
and I_6399 (I111422,I111590,I111768);
nand I_6400 (I111799,I111474,I107685);
not I_6401 (I111816,I111799);
nor I_6402 (I111833,I111675,I111816);
DFFARX1 I_6403 (I111850,I107679,I2966,I111457,);
nand I_6404 (I111867,I111850,I111799);
and I_6405 (I111884,I111590,I111867);
DFFARX1 I_6406 (I111449,I111884,I2966,I111457,);
not I_6407 (I111915,I111850);
nand I_6408 (I111437,I111850,I111833);
nand I_6409 (I111431,I111850,I111816);
DFFARX1 I_6410 (I111960,I107691,I2966,I111457,);
not I_6411 (I111977,I111960);
nor I_6412 (I111446,I111850,I111977);
nor I_6413 (I112008,I111977,I111915);
and I_6414 (I112025,I111556,I112008);
or I_6415 (I112042,I111799,I112025);
DFFARX1 I_6416 (I111434,I112042,I2966,I111457,);
DFFARX1 I_6417 (I111419,I111977,I2966,I111457,);
not I_6418 (I112120,I2973);
not I_6419 (I112137,I96868);
nor I_6420 (I112154,I96877,I96850);
nand I_6421 (I112171,I112154,I96862);
DFFARX1 I_6422 (I112091,I112171,I2966,I112120,);
nor I_6423 (I112202,I112137,I96877);
nand I_6424 (I112219,I112202,I96874);
nand I_6425 (I112236,I112219,I112171);
not I_6426 (I112253,I96877);
not I_6427 (I112270,I96853);
nor I_6428 (I112287,I112270,I96859);
and I_6429 (I112304,I112287,I96871);
or I_6430 (I112321,I112304,I96856);
DFFARX1 I_6431 (I112338,I112321,I2966,I112120,);
nor I_6432 (I112355,I112338,I112219);
nand I_6433 (I112106,I112253,I112355);
not I_6434 (I112103,I112338);
and I_6435 (I112400,I112338,I112236);
DFFARX1 I_6436 (I112088,I112400,I2966,I112120,);
DFFARX1 I_6437 (I112431,I112338,I2966,I112120,);
and I_6438 (I112085,I112253,I112431);
nand I_6439 (I112462,I112137,I96853);
not I_6440 (I112479,I112462);
nor I_6441 (I112496,I112338,I112479);
DFFARX1 I_6442 (I112513,I96880,I2966,I112120,);
nand I_6443 (I112530,I112513,I112462);
and I_6444 (I112547,I112253,I112530);
DFFARX1 I_6445 (I112112,I112547,I2966,I112120,);
not I_6446 (I112578,I112513);
nand I_6447 (I112100,I112513,I112496);
nand I_6448 (I112094,I112513,I112479);
DFFARX1 I_6449 (I112623,I96865,I2966,I112120,);
not I_6450 (I112640,I112623);
nor I_6451 (I112109,I112513,I112640);
nor I_6452 (I112671,I112640,I112578);
and I_6453 (I112688,I112219,I112671);
or I_6454 (I112705,I112462,I112688);
DFFARX1 I_6455 (I112097,I112705,I2966,I112120,);
DFFARX1 I_6456 (I112082,I112640,I2966,I112120,);
not I_6457 (I112783,I2973);
not I_6458 (I112800,I94284);
nor I_6459 (I112817,I94293,I94266);
nand I_6460 (I112834,I112817,I94278);
DFFARX1 I_6461 (I112754,I112834,I2966,I112783,);
nor I_6462 (I112865,I112800,I94293);
nand I_6463 (I112882,I112865,I94290);
nand I_6464 (I112899,I112882,I112834);
not I_6465 (I112916,I94293);
not I_6466 (I112933,I94269);
nor I_6467 (I112950,I112933,I94275);
and I_6468 (I112967,I112950,I94287);
or I_6469 (I112984,I112967,I94272);
DFFARX1 I_6470 (I113001,I112984,I2966,I112783,);
nor I_6471 (I113018,I113001,I112882);
nand I_6472 (I112769,I112916,I113018);
not I_6473 (I112766,I113001);
and I_6474 (I113063,I113001,I112899);
DFFARX1 I_6475 (I112751,I113063,I2966,I112783,);
DFFARX1 I_6476 (I113094,I113001,I2966,I112783,);
and I_6477 (I112748,I112916,I113094);
nand I_6478 (I113125,I112800,I94269);
not I_6479 (I113142,I113125);
nor I_6480 (I113159,I113001,I113142);
DFFARX1 I_6481 (I113176,I94296,I2966,I112783,);
nand I_6482 (I113193,I113176,I113125);
and I_6483 (I113210,I112916,I113193);
DFFARX1 I_6484 (I112775,I113210,I2966,I112783,);
not I_6485 (I113241,I113176);
nand I_6486 (I112763,I113176,I113159);
nand I_6487 (I112757,I113176,I113142);
DFFARX1 I_6488 (I113286,I94281,I2966,I112783,);
not I_6489 (I113303,I113286);
nor I_6490 (I112772,I113176,I113303);
nor I_6491 (I113334,I113303,I113241);
and I_6492 (I113351,I112882,I113334);
or I_6493 (I113368,I113125,I113351);
DFFARX1 I_6494 (I112760,I113368,I2966,I112783,);
DFFARX1 I_6495 (I112745,I113303,I2966,I112783,);
not I_6496 (I113446,I2973);
not I_6497 (I113463,I96222);
nor I_6498 (I113480,I96231,I96204);
nand I_6499 (I113497,I113480,I96216);
DFFARX1 I_6500 (I113417,I113497,I2966,I113446,);
nor I_6501 (I113528,I113463,I96231);
nand I_6502 (I113545,I113528,I96228);
nand I_6503 (I113562,I113545,I113497);
not I_6504 (I113579,I96231);
not I_6505 (I113596,I96207);
nor I_6506 (I113613,I113596,I96213);
and I_6507 (I113630,I113613,I96225);
or I_6508 (I113647,I113630,I96210);
DFFARX1 I_6509 (I113664,I113647,I2966,I113446,);
nor I_6510 (I113681,I113664,I113545);
nand I_6511 (I113432,I113579,I113681);
not I_6512 (I113429,I113664);
and I_6513 (I113726,I113664,I113562);
DFFARX1 I_6514 (I113414,I113726,I2966,I113446,);
DFFARX1 I_6515 (I113757,I113664,I2966,I113446,);
and I_6516 (I113411,I113579,I113757);
nand I_6517 (I113788,I113463,I96207);
not I_6518 (I113805,I113788);
nor I_6519 (I113822,I113664,I113805);
DFFARX1 I_6520 (I113839,I96234,I2966,I113446,);
nand I_6521 (I113856,I113839,I113788);
and I_6522 (I113873,I113579,I113856);
DFFARX1 I_6523 (I113438,I113873,I2966,I113446,);
not I_6524 (I113904,I113839);
nand I_6525 (I113426,I113839,I113822);
nand I_6526 (I113420,I113839,I113805);
DFFARX1 I_6527 (I113949,I96219,I2966,I113446,);
not I_6528 (I113966,I113949);
nor I_6529 (I113435,I113839,I113966);
nor I_6530 (I113997,I113966,I113904);
and I_6531 (I114014,I113545,I113997);
or I_6532 (I114031,I113788,I114014);
DFFARX1 I_6533 (I113423,I114031,I2966,I113446,);
DFFARX1 I_6534 (I113408,I113966,I2966,I113446,);
not I_6535 (I114109,I2973);
or I_6536 (I114126,I103424,I103418);
or I_6537 (I114143,I103412,I103424);
DFFARX1 I_6538 (I114083,I114143,I2966,I114109,);
nor I_6539 (I114174,I103415,I103421);
not I_6540 (I114191,I114174);
not I_6541 (I114208,I103415);
and I_6542 (I114225,I114208,I103439);
nor I_6543 (I114242,I114225,I103418);
nor I_6544 (I114259,I103442,I103433);
DFFARX1 I_6545 (I114276,I114259,I2966,I114109,);
nand I_6546 (I114293,I114276,I114126);
and I_6547 (I114310,I114242,I114293);
DFFARX1 I_6548 (I114077,I114310,I2966,I114109,);
nor I_6549 (I114341,I103442,I103412);
DFFARX1 I_6550 (I114358,I114341,I2966,I114109,);
and I_6551 (I114074,I114174,I114358);
DFFARX1 I_6552 (I114389,I103430,I2966,I114109,);
and I_6553 (I114406,I114389,I103427);
DFFARX1 I_6554 (I114423,I114406,I2966,I114109,);
not I_6555 (I114086,I114423);
DFFARX1 I_6556 (I114071,I114406,I2966,I114109,);
DFFARX1 I_6557 (I114468,I103436,I2966,I114109,);
not I_6558 (I114485,I114468);
nor I_6559 (I114502,I114143,I114485);
and I_6560 (I114519,I114406,I114502);
or I_6561 (I114536,I114126,I114519);
DFFARX1 I_6562 (I114092,I114536,I2966,I114109,);
nor I_6563 (I114567,I114468,I114276);
nand I_6564 (I114101,I114242,I114567);
nor I_6565 (I114598,I114468,I114191);
nand I_6566 (I114095,I114341,I114598);
not I_6567 (I114098,I114468);
nand I_6568 (I114089,I114468,I114191);
DFFARX1 I_6569 (I114080,I114468,I2966,I114109,);
not I_6570 (I114704,I2973);
or I_6571 (I114721,I98074,I98104);
not I_6572 (I114687,I114721);
DFFARX1 I_6573 (I114666,I114721,I2966,I114704,);
or I_6574 (I114766,I98083,I98074);
nor I_6575 (I114783,I98089,I98086);
nor I_6576 (I114800,I114783,I114721);
not I_6577 (I114817,I98089);
and I_6578 (I114834,I114817,I98095);
nor I_6579 (I114851,I114834,I98104);
DFFARX1 I_6580 (I114868,I114851,I2966,I114704,);
nor I_6581 (I114885,I98080,I98098);
DFFARX1 I_6582 (I114902,I114885,I2966,I114704,);
nor I_6583 (I114693,I114902,I114851);
not I_6584 (I114933,I114902);
nor I_6585 (I114950,I98080,I98083);
nand I_6586 (I114967,I114851,I114950);
and I_6587 (I114984,I114766,I114967);
DFFARX1 I_6588 (I114696,I114984,I2966,I114704,);
DFFARX1 I_6589 (I115015,I98101,I2966,I114704,);
and I_6590 (I115032,I115015,I98092);
nor I_6591 (I115049,I115032,I114933);
and I_6592 (I115066,I114950,I115049);
or I_6593 (I115083,I114783,I115066);
DFFARX1 I_6594 (I114681,I115083,I2966,I114704,);
not I_6595 (I115114,I115032);
nor I_6596 (I115131,I114721,I115114);
nand I_6597 (I114684,I114766,I115131);
nand I_6598 (I114678,I114902,I115114);
DFFARX1 I_6599 (I114672,I115032,I2966,I114704,);
DFFARX1 I_6600 (I115190,I98077,I2966,I114704,);
nand I_6601 (I114690,I115190,I114800);
DFFARX1 I_6602 (I115221,I115190,I2966,I114704,);
not I_6603 (I114675,I115221);
and I_6604 (I114669,I115190,I114868);
not I_6605 (I115299,I2973);
or I_6606 (I115316,I99267,I99288);
not I_6607 (I115282,I115316);
DFFARX1 I_6608 (I115261,I115316,I2966,I115299,);
or I_6609 (I115361,I99264,I99267);
nor I_6610 (I115378,I99285,I99291);
nor I_6611 (I115395,I115378,I115316);
not I_6612 (I115412,I99285);
and I_6613 (I115429,I115412,I99279);
nor I_6614 (I115446,I115429,I99288);
DFFARX1 I_6615 (I115463,I115446,I2966,I115299,);
nor I_6616 (I115480,I99294,I99282);
DFFARX1 I_6617 (I115497,I115480,I2966,I115299,);
nor I_6618 (I115288,I115497,I115446);
not I_6619 (I115528,I115497);
nor I_6620 (I115545,I99294,I99264);
nand I_6621 (I115562,I115446,I115545);
and I_6622 (I115579,I115361,I115562);
DFFARX1 I_6623 (I115291,I115579,I2966,I115299,);
DFFARX1 I_6624 (I115610,I99276,I2966,I115299,);
and I_6625 (I115627,I115610,I99273);
nor I_6626 (I115644,I115627,I115528);
and I_6627 (I115661,I115545,I115644);
or I_6628 (I115678,I115378,I115661);
DFFARX1 I_6629 (I115276,I115678,I2966,I115299,);
not I_6630 (I115709,I115627);
nor I_6631 (I115726,I115316,I115709);
nand I_6632 (I115279,I115361,I115726);
nand I_6633 (I115273,I115497,I115709);
DFFARX1 I_6634 (I115267,I115627,I2966,I115299,);
DFFARX1 I_6635 (I115785,I99270,I2966,I115299,);
nand I_6636 (I115285,I115785,I115395);
DFFARX1 I_6637 (I115816,I115785,I2966,I115299,);
not I_6638 (I115270,I115816);
and I_6639 (I115264,I115785,I115463);
not I_6640 (I115894,I2973);
not I_6641 (I115911,I104013);
nor I_6642 (I115928,I104031,I104022);
nand I_6643 (I115945,I115928,I104028);
nor I_6644 (I115962,I115911,I104031);
nand I_6645 (I115979,I115962,I104034);
not I_6646 (I115996,I115979);
not I_6647 (I116013,I104031);
nor I_6648 (I115883,I115979,I116013);
not I_6649 (I116044,I116013);
nand I_6650 (I115868,I115979,I116044);
not I_6651 (I116075,I104010);
nor I_6652 (I116092,I116075,I104025);
and I_6653 (I116109,I116092,I104007);
or I_6654 (I116126,I116109,I104016);
DFFARX1 I_6655 (I116143,I116126,I2966,I115894,);
nor I_6656 (I116160,I116143,I115996);
DFFARX1 I_6657 (I116177,I116143,I2966,I115894,);
not I_6658 (I115865,I116177);
nand I_6659 (I116208,I115911,I104010);
and I_6660 (I116225,I116208,I116160);
DFFARX1 I_6661 (I115862,I116208,I2966,I115894,);
DFFARX1 I_6662 (I116256,I104019,I2966,I115894,);
nor I_6663 (I116273,I116256,I115979);
nand I_6664 (I115880,I116143,I116273);
nor I_6665 (I116304,I116256,I116044);
not I_6666 (I115877,I116256);
nand I_6667 (I116335,I116256,I115945);
and I_6668 (I116352,I116013,I116335);
DFFARX1 I_6669 (I115856,I116352,I2966,I115894,);
DFFARX1 I_6670 (I115859,I116256,I2966,I115894,);
DFFARX1 I_6671 (I116397,I104037,I2966,I115894,);
not I_6672 (I116414,I116397);
nand I_6673 (I116431,I116414,I115979);
and I_6674 (I116448,I116208,I116431);
DFFARX1 I_6675 (I115886,I116448,I2966,I115894,);
or I_6676 (I116479,I116414,I116225);
DFFARX1 I_6677 (I115871,I116479,I2966,I115894,);
nand I_6678 (I115874,I116414,I116304);
not I_6679 (I116557,I2973);
not I_6680 (I116574,I105271);
nor I_6681 (I116591,I105289,I105280);
nand I_6682 (I116608,I116591,I105286);
nor I_6683 (I116625,I116574,I105289);
nand I_6684 (I116642,I116625,I105292);
not I_6685 (I116659,I116642);
not I_6686 (I116676,I105289);
nor I_6687 (I116546,I116642,I116676);
not I_6688 (I116707,I116676);
nand I_6689 (I116531,I116642,I116707);
not I_6690 (I116738,I105268);
nor I_6691 (I116755,I116738,I105283);
and I_6692 (I116772,I116755,I105265);
or I_6693 (I116789,I116772,I105274);
DFFARX1 I_6694 (I116806,I116789,I2966,I116557,);
nor I_6695 (I116823,I116806,I116659);
DFFARX1 I_6696 (I116840,I116806,I2966,I116557,);
not I_6697 (I116528,I116840);
nand I_6698 (I116871,I116574,I105268);
and I_6699 (I116888,I116871,I116823);
DFFARX1 I_6700 (I116525,I116871,I2966,I116557,);
DFFARX1 I_6701 (I116919,I105277,I2966,I116557,);
nor I_6702 (I116936,I116919,I116642);
nand I_6703 (I116543,I116806,I116936);
nor I_6704 (I116967,I116919,I116707);
not I_6705 (I116540,I116919);
nand I_6706 (I116998,I116919,I116608);
and I_6707 (I117015,I116676,I116998);
DFFARX1 I_6708 (I116519,I117015,I2966,I116557,);
DFFARX1 I_6709 (I116522,I116919,I2966,I116557,);
DFFARX1 I_6710 (I117060,I105295,I2966,I116557,);
not I_6711 (I117077,I117060);
nand I_6712 (I117094,I117077,I116642);
and I_6713 (I117111,I116871,I117094);
DFFARX1 I_6714 (I116549,I117111,I2966,I116557,);
or I_6715 (I117142,I117077,I116888);
DFFARX1 I_6716 (I116534,I117142,I2966,I116557,);
nand I_6717 (I116537,I117077,I116967);
not I_6718 (I117220,I2973);
not I_6719 (I117237,I112748);
nor I_6720 (I117254,I112754,I112760);
nand I_6721 (I117271,I117254,I112763);
nor I_6722 (I117288,I117237,I112754);
nand I_6723 (I117305,I117288,I112745);
not I_6724 (I117322,I117305);
not I_6725 (I117339,I112754);
nor I_6726 (I117209,I117305,I117339);
not I_6727 (I117370,I117339);
nand I_6728 (I117194,I117305,I117370);
not I_6729 (I117401,I112757);
nor I_6730 (I117418,I117401,I112751);
and I_6731 (I117435,I117418,I112766);
or I_6732 (I117452,I117435,I112772);
DFFARX1 I_6733 (I117469,I117452,I2966,I117220,);
nor I_6734 (I117486,I117469,I117322);
DFFARX1 I_6735 (I117503,I117469,I2966,I117220,);
not I_6736 (I117191,I117503);
nand I_6737 (I117534,I117237,I112757);
and I_6738 (I117551,I117534,I117486);
DFFARX1 I_6739 (I117188,I117534,I2966,I117220,);
DFFARX1 I_6740 (I117582,I112769,I2966,I117220,);
nor I_6741 (I117599,I117582,I117305);
nand I_6742 (I117206,I117469,I117599);
nor I_6743 (I117630,I117582,I117370);
not I_6744 (I117203,I117582);
nand I_6745 (I117661,I117582,I117271);
and I_6746 (I117678,I117339,I117661);
DFFARX1 I_6747 (I117182,I117678,I2966,I117220,);
DFFARX1 I_6748 (I117185,I117582,I2966,I117220,);
DFFARX1 I_6749 (I117723,I112775,I2966,I117220,);
not I_6750 (I117740,I117723);
nand I_6751 (I117757,I117740,I117305);
and I_6752 (I117774,I117534,I117757);
DFFARX1 I_6753 (I117212,I117774,I2966,I117220,);
or I_6754 (I117805,I117740,I117551);
DFFARX1 I_6755 (I117197,I117805,I2966,I117220,);
nand I_6756 (I117200,I117740,I117630);
not I_6757 (I117883,I2973);
not I_6758 (I117900,I110759);
nor I_6759 (I117917,I110765,I110771);
nand I_6760 (I117934,I117917,I110774);
nor I_6761 (I117951,I117900,I110765);
nand I_6762 (I117968,I117951,I110756);
not I_6763 (I117985,I117968);
not I_6764 (I118002,I110765);
nor I_6765 (I117872,I117968,I118002);
not I_6766 (I118033,I118002);
nand I_6767 (I117857,I117968,I118033);
not I_6768 (I118064,I110768);
nor I_6769 (I118081,I118064,I110762);
and I_6770 (I118098,I118081,I110777);
or I_6771 (I118115,I118098,I110783);
DFFARX1 I_6772 (I118132,I118115,I2966,I117883,);
nor I_6773 (I118149,I118132,I117985);
DFFARX1 I_6774 (I118166,I118132,I2966,I117883,);
not I_6775 (I117854,I118166);
nand I_6776 (I118197,I117900,I110768);
and I_6777 (I118214,I118197,I118149);
DFFARX1 I_6778 (I117851,I118197,I2966,I117883,);
DFFARX1 I_6779 (I118245,I110780,I2966,I117883,);
nor I_6780 (I118262,I118245,I117968);
nand I_6781 (I117869,I118132,I118262);
nor I_6782 (I118293,I118245,I118033);
not I_6783 (I117866,I118245);
nand I_6784 (I118324,I118245,I117934);
and I_6785 (I118341,I118002,I118324);
DFFARX1 I_6786 (I117845,I118341,I2966,I117883,);
DFFARX1 I_6787 (I117848,I118245,I2966,I117883,);
DFFARX1 I_6788 (I118386,I110786,I2966,I117883,);
not I_6789 (I118403,I118386);
nand I_6790 (I118420,I118403,I117968);
and I_6791 (I118437,I118197,I118420);
DFFARX1 I_6792 (I117875,I118437,I2966,I117883,);
or I_6793 (I118468,I118403,I118214);
DFFARX1 I_6794 (I117860,I118468,I2966,I117883,);
nand I_6795 (I117863,I118403,I118293);
not I_6796 (I118546,I2973);
not I_6797 (I118563,I94924);
nor I_6798 (I118580,I94921,I94939);
nand I_6799 (I118597,I118580,I94942);
nor I_6800 (I118614,I118563,I94921);
nand I_6801 (I118631,I118614,I94927);
not I_6802 (I118648,I118631);
not I_6803 (I118665,I94921);
nor I_6804 (I118535,I118631,I118665);
not I_6805 (I118696,I118665);
nand I_6806 (I118520,I118631,I118696);
not I_6807 (I118727,I94936);
nor I_6808 (I118744,I118727,I94918);
and I_6809 (I118761,I118744,I94912);
or I_6810 (I118778,I118761,I94930);
DFFARX1 I_6811 (I118795,I118778,I2966,I118546,);
nor I_6812 (I118812,I118795,I118648);
DFFARX1 I_6813 (I118829,I118795,I2966,I118546,);
not I_6814 (I118517,I118829);
nand I_6815 (I118860,I118563,I94936);
and I_6816 (I118877,I118860,I118812);
DFFARX1 I_6817 (I118514,I118860,I2966,I118546,);
DFFARX1 I_6818 (I118908,I94915,I2966,I118546,);
nor I_6819 (I118925,I118908,I118631);
nand I_6820 (I118532,I118795,I118925);
nor I_6821 (I118956,I118908,I118696);
not I_6822 (I118529,I118908);
nand I_6823 (I118987,I118908,I118597);
and I_6824 (I119004,I118665,I118987);
DFFARX1 I_6825 (I118508,I119004,I2966,I118546,);
DFFARX1 I_6826 (I118511,I118908,I2966,I118546,);
DFFARX1 I_6827 (I119049,I94933,I2966,I118546,);
not I_6828 (I119066,I119049);
nand I_6829 (I119083,I119066,I118631);
and I_6830 (I119100,I118860,I119083);
DFFARX1 I_6831 (I118538,I119100,I2966,I118546,);
or I_6832 (I119131,I119066,I118877);
DFFARX1 I_6833 (I118523,I119131,I2966,I118546,);
nand I_6834 (I118526,I119066,I118956);
not I_6835 (I119209,I2973);
not I_6836 (I119226,I108266);
nor I_6837 (I119243,I108281,I108275);
nand I_6838 (I119260,I119243,I108284);
nor I_6839 (I119277,I119226,I108281);
nand I_6840 (I119294,I119277,I108260);
DFFARX1 I_6841 (I119311,I119294,I2966,I119209,);
not I_6842 (I119180,I119311);
not I_6843 (I119342,I108281);
not I_6844 (I119359,I119342);
not I_6845 (I119376,I108257);
nor I_6846 (I119393,I119376,I108272);
and I_6847 (I119410,I119393,I108278);
or I_6848 (I119427,I119410,I108287);
DFFARX1 I_6849 (I119444,I119427,I2966,I119209,);
DFFARX1 I_6850 (I119177,I119444,I2966,I119209,);
DFFARX1 I_6851 (I119475,I119444,I2966,I119209,);
DFFARX1 I_6852 (I119171,I119444,I2966,I119209,);
nand I_6853 (I119506,I119226,I108257);
nand I_6854 (I119523,I119506,I119260);
and I_6855 (I119540,I119342,I119523);
DFFARX1 I_6856 (I119201,I119540,I2966,I119209,);
and I_6857 (I119174,I119506,I119475);
DFFARX1 I_6858 (I119585,I108269,I2966,I119209,);
nor I_6859 (I119198,I119585,I119506);
nor I_6860 (I119616,I119585,I119260);
nand I_6861 (I119195,I119294,I119616);
not I_6862 (I119192,I119585);
DFFARX1 I_6863 (I119661,I108263,I2966,I119209,);
not I_6864 (I119678,I119661);
nor I_6865 (I119695,I119678,I119359);
and I_6866 (I119712,I119585,I119695);
or I_6867 (I119729,I119506,I119712);
DFFARX1 I_6868 (I119186,I119729,I2966,I119209,);
not I_6869 (I119760,I119678);
nor I_6870 (I119777,I119585,I119760);
nand I_6871 (I119189,I119678,I119777);
nand I_6872 (I119183,I119342,I119760);
not I_6873 (I119855,I2973);
or I_6874 (I119872,I108818,I108845);
or I_6875 (I119889,I108833,I108818);
nor I_6876 (I119906,I108842,I108821);
DFFARX1 I_6877 (I119923,I119906,I2966,I119855,);
DFFARX1 I_6878 (I119817,I119906,I2966,I119855,);
not I_6879 (I119954,I108842);
and I_6880 (I119971,I119954,I108839);
nor I_6881 (I119988,I119971,I108845);
nor I_6882 (I120005,I108836,I108824);
DFFARX1 I_6883 (I120022,I120005,I2966,I119855,);
not I_6884 (I120039,I120022);
DFFARX1 I_6885 (I119826,I120022,I2966,I119855,);
nor I_6886 (I120070,I108836,I108833);
and I_6887 (I119820,I120070,I119923);
DFFARX1 I_6888 (I120101,I108848,I2966,I119855,);
and I_6889 (I120118,I120101,I108830);
nand I_6890 (I120135,I120118,I119889);
and I_6891 (I120152,I120022,I120135);
DFFARX1 I_6892 (I119847,I120152,I2966,I119855,);
nor I_6893 (I119844,I120118,I119988);
not I_6894 (I120197,I120118);
nor I_6895 (I120214,I119872,I120197);
nor I_6896 (I120231,I120118,I120070);
nand I_6897 (I119841,I119889,I120231);
nor I_6898 (I120262,I120118,I120039);
not I_6899 (I119838,I120118);
nand I_6900 (I119829,I120118,I120039);
DFFARX1 I_6901 (I120307,I108827,I2966,I119855,);
and I_6902 (I120324,I120307,I120214);
or I_6903 (I120341,I119872,I120324);
DFFARX1 I_6904 (I119832,I120341,I2966,I119855,);
nand I_6905 (I119835,I120307,I120262);
nand I_6906 (I120386,I120307,I119988);
and I_6907 (I120403,I119906,I120386);
DFFARX1 I_6908 (I119823,I120403,I2966,I119855,);
not I_6909 (I120467,I2973);
nand I_6910 (I120484,I114666,I114669);
and I_6911 (I120501,I120484,I114675);
DFFARX1 I_6912 (I120518,I120501,I2966,I120467,);
not I_6913 (I120535,I120518);
DFFARX1 I_6914 (I120435,I120518,I2966,I120467,);
nor I_6915 (I120566,I114687,I114669);
DFFARX1 I_6916 (I120583,I114678,I2966,I120467,);
DFFARX1 I_6917 (I120600,I120583,I2966,I120467,);
not I_6918 (I120438,I120600);
DFFARX1 I_6919 (I120631,I120583,I2966,I120467,);
and I_6920 (I120432,I120518,I120631);
nand I_6921 (I120662,I114684,I114681);
and I_6922 (I120679,I120662,I114693);
DFFARX1 I_6923 (I120696,I120679,I2966,I120467,);
nor I_6924 (I120713,I120696,I120535);
not I_6925 (I120730,I120696);
nand I_6926 (I120441,I120518,I120730);
DFFARX1 I_6927 (I120761,I114690,I2966,I120467,);
and I_6928 (I120778,I120761,I114696);
nor I_6929 (I120795,I120778,I120696);
nor I_6930 (I120812,I120778,I120730);
nand I_6931 (I120447,I120566,I120812);
not I_6932 (I120450,I120778);
DFFARX1 I_6933 (I120429,I120778,I2966,I120467,);
DFFARX1 I_6934 (I120871,I114672,I2966,I120467,);
nand I_6935 (I120888,I120871,I120583);
and I_6936 (I120905,I120566,I120888);
DFFARX1 I_6937 (I120459,I120905,I2966,I120467,);
nor I_6938 (I120456,I120871,I120778);
and I_6939 (I120950,I120871,I120713);
or I_6940 (I120967,I120566,I120950);
DFFARX1 I_6941 (I120444,I120967,I2966,I120467,);
nand I_6942 (I120453,I120871,I120795);
not I_6943 (I121045,I2973);
nand I_6944 (I121062,I117848,I117875);
and I_6945 (I121079,I121062,I117863);
DFFARX1 I_6946 (I121096,I121079,I2966,I121045,);
not I_6947 (I121113,I121096);
DFFARX1 I_6948 (I121013,I121096,I2966,I121045,);
nor I_6949 (I121144,I117851,I117875);
DFFARX1 I_6950 (I121161,I117866,I2966,I121045,);
DFFARX1 I_6951 (I121178,I121161,I2966,I121045,);
not I_6952 (I121016,I121178);
DFFARX1 I_6953 (I121209,I121161,I2966,I121045,);
and I_6954 (I121010,I121096,I121209);
nand I_6955 (I121240,I117860,I117857);
and I_6956 (I121257,I121240,I117854);
DFFARX1 I_6957 (I121274,I121257,I2966,I121045,);
nor I_6958 (I121291,I121274,I121113);
not I_6959 (I121308,I121274);
nand I_6960 (I121019,I121096,I121308);
DFFARX1 I_6961 (I121339,I117869,I2966,I121045,);
and I_6962 (I121356,I121339,I117845);
nor I_6963 (I121373,I121356,I121274);
nor I_6964 (I121390,I121356,I121308);
nand I_6965 (I121025,I121144,I121390);
not I_6966 (I121028,I121356);
DFFARX1 I_6967 (I121007,I121356,I2966,I121045,);
DFFARX1 I_6968 (I121449,I117872,I2966,I121045,);
nand I_6969 (I121466,I121449,I121161);
and I_6970 (I121483,I121144,I121466);
DFFARX1 I_6971 (I121037,I121483,I2966,I121045,);
nor I_6972 (I121034,I121449,I121356);
and I_6973 (I121528,I121449,I121291);
or I_6974 (I121545,I121144,I121528);
DFFARX1 I_6975 (I121022,I121545,I2966,I121045,);
nand I_6976 (I121031,I121449,I121373);
not I_6977 (I121623,I2973);
nand I_6978 (I121640,I101654,I101642);
and I_6979 (I121657,I121640,I101636);
DFFARX1 I_6980 (I121674,I121657,I2966,I121623,);
not I_6981 (I121691,I121674);
DFFARX1 I_6982 (I121591,I121674,I2966,I121623,);
nor I_6983 (I121722,I101633,I101642);
DFFARX1 I_6984 (I121739,I101627,I2966,I121623,);
DFFARX1 I_6985 (I121756,I121739,I2966,I121623,);
not I_6986 (I121594,I121756);
DFFARX1 I_6987 (I121787,I121739,I2966,I121623,);
and I_6988 (I121588,I121674,I121787);
nand I_6989 (I121818,I101630,I101645);
and I_6990 (I121835,I121818,I101657);
DFFARX1 I_6991 (I121852,I121835,I2966,I121623,);
nor I_6992 (I121869,I121852,I121691);
not I_6993 (I121886,I121852);
nand I_6994 (I121597,I121674,I121886);
DFFARX1 I_6995 (I121917,I101648,I2966,I121623,);
and I_6996 (I121934,I121917,I101639);
nor I_6997 (I121951,I121934,I121852);
nor I_6998 (I121968,I121934,I121886);
nand I_6999 (I121603,I121722,I121968);
not I_7000 (I121606,I121934);
DFFARX1 I_7001 (I121585,I121934,I2966,I121623,);
DFFARX1 I_7002 (I122027,I101651,I2966,I121623,);
nand I_7003 (I122044,I122027,I121739);
and I_7004 (I122061,I121722,I122044);
DFFARX1 I_7005 (I121615,I122061,I2966,I121623,);
nor I_7006 (I121612,I122027,I121934);
and I_7007 (I122106,I122027,I121869);
or I_7008 (I122123,I121722,I122106);
DFFARX1 I_7009 (I121600,I122123,I2966,I121623,);
nand I_7010 (I121609,I122027,I121951);
not I_7011 (I122201,I2973);
nand I_7012 (I122218,I100464,I100452);
and I_7013 (I122235,I122218,I100446);
DFFARX1 I_7014 (I122252,I122235,I2966,I122201,);
not I_7015 (I122269,I122252);
DFFARX1 I_7016 (I122169,I122252,I2966,I122201,);
nor I_7017 (I122300,I100443,I100452);
DFFARX1 I_7018 (I122317,I100437,I2966,I122201,);
DFFARX1 I_7019 (I122334,I122317,I2966,I122201,);
not I_7020 (I122172,I122334);
DFFARX1 I_7021 (I122365,I122317,I2966,I122201,);
and I_7022 (I122166,I122252,I122365);
nand I_7023 (I122396,I100440,I100455);
and I_7024 (I122413,I122396,I100467);
DFFARX1 I_7025 (I122430,I122413,I2966,I122201,);
nor I_7026 (I122447,I122430,I122269);
not I_7027 (I122464,I122430);
nand I_7028 (I122175,I122252,I122464);
DFFARX1 I_7029 (I122495,I100458,I2966,I122201,);
and I_7030 (I122512,I122495,I100449);
nor I_7031 (I122529,I122512,I122430);
nor I_7032 (I122546,I122512,I122464);
nand I_7033 (I122181,I122300,I122546);
not I_7034 (I122184,I122512);
DFFARX1 I_7035 (I122163,I122512,I2966,I122201,);
DFFARX1 I_7036 (I122605,I100461,I2966,I122201,);
nand I_7037 (I122622,I122605,I122317);
and I_7038 (I122639,I122300,I122622);
DFFARX1 I_7039 (I122193,I122639,I2966,I122201,);
nor I_7040 (I122190,I122605,I122512);
and I_7041 (I122684,I122605,I122447);
or I_7042 (I122701,I122300,I122684);
DFFARX1 I_7043 (I122178,I122701,I2966,I122201,);
nand I_7044 (I122187,I122605,I122529);
not I_7045 (I122779,I2973);
or I_7046 (I122796,I109473,I109464);
or I_7047 (I122813,I109470,I109473);
nor I_7048 (I122830,I109479,I109488);
or I_7049 (I122768,I122830,I122796);
not I_7050 (I122861,I109479);
and I_7051 (I122878,I122861,I109491);
nor I_7052 (I122895,I122878,I109464);
not I_7053 (I122912,I122895);
nor I_7054 (I122929,I109482,I109485);
DFFARX1 I_7055 (I122946,I122929,I2966,I122779,);
nor I_7056 (I122963,I122946,I122895);
nand I_7057 (I122753,I122796,I122963);
nor I_7058 (I122994,I122946,I122912);
not I_7059 (I122750,I122946);
nor I_7060 (I123025,I109482,I109470);
or I_7061 (I122762,I122796,I123025);
DFFARX1 I_7062 (I123056,I109467,I2966,I122779,);
and I_7063 (I123073,I123056,I109476);
nor I_7064 (I123090,I123073,I122946);
DFFARX1 I_7065 (I122756,I123090,I2966,I122779,);
nor I_7066 (I122771,I123073,I123025);
not I_7067 (I123135,I123073);
nor I_7068 (I123152,I122813,I123135);
nand I_7069 (I122741,I123073,I122912);
DFFARX1 I_7070 (I123183,I109494,I2966,I122779,);
nor I_7071 (I122759,I123183,I122813);
not I_7072 (I123214,I123183);
and I_7073 (I123231,I123025,I123214);
nor I_7074 (I122765,I122830,I123231);
and I_7075 (I123262,I123183,I123152);
or I_7076 (I123279,I122830,I123262);
DFFARX1 I_7077 (I122744,I123279,I2966,I122779,);
nand I_7078 (I122747,I123183,I122994);
not I_7079 (I123357,I2973);
nand I_7080 (I123374,I110119,I110131);
and I_7081 (I123391,I123374,I110140);
DFFARX1 I_7082 (I123408,I123391,I2966,I123357,);
nor I_7083 (I123425,I110134,I110131);
nor I_7084 (I123442,I123425,I123408);
not I_7085 (I123340,I123425);
DFFARX1 I_7086 (I123473,I110128,I2966,I123357,);
not I_7087 (I123490,I123473);
nor I_7088 (I123507,I123425,I123490);
nand I_7089 (I123343,I123473,I123442);
DFFARX1 I_7090 (I123325,I123473,I2966,I123357,);
nand I_7091 (I123552,I110125,I110122);
and I_7092 (I123569,I123552,I110113);
DFFARX1 I_7093 (I123586,I123569,I2966,I123357,);
nor I_7094 (I123346,I123586,I123408);
nand I_7095 (I123337,I123586,I123507);
DFFARX1 I_7096 (I123631,I110137,I2966,I123357,);
and I_7097 (I123648,I123631,I110116);
DFFARX1 I_7098 (I123665,I123648,I2966,I123357,);
not I_7099 (I123328,I123665);
nand I_7100 (I123696,I123648,I123586);
and I_7101 (I123713,I123408,I123696);
DFFARX1 I_7102 (I123319,I123713,I2966,I123357,);
DFFARX1 I_7103 (I123744,I110110,I2966,I123357,);
nand I_7104 (I123761,I123744,I123408);
and I_7105 (I123778,I123586,I123761);
DFFARX1 I_7106 (I123349,I123778,I2966,I123357,);
not I_7107 (I123809,I123744);
nor I_7108 (I123826,I123425,I123809);
and I_7109 (I123843,I123744,I123826);
or I_7110 (I123860,I123648,I123843);
DFFARX1 I_7111 (I123334,I123860,I2966,I123357,);
nand I_7112 (I123331,I123744,I123490);
DFFARX1 I_7113 (I123322,I123744,I2966,I123357,);
not I_7114 (I123952,I2973);
nand I_7115 (I123969,I105912,I105903);
and I_7116 (I123986,I123969,I105921);
DFFARX1 I_7117 (I124003,I123986,I2966,I123952,);
nor I_7118 (I124020,I105918,I105903);
nor I_7119 (I124037,I124020,I124003);
not I_7120 (I123935,I124020);
DFFARX1 I_7121 (I124068,I105900,I2966,I123952,);
not I_7122 (I124085,I124068);
nor I_7123 (I124102,I124020,I124085);
nand I_7124 (I123938,I124068,I124037);
DFFARX1 I_7125 (I123920,I124068,I2966,I123952,);
nand I_7126 (I124147,I105909,I105924);
and I_7127 (I124164,I124147,I105915);
DFFARX1 I_7128 (I124181,I124164,I2966,I123952,);
nor I_7129 (I123941,I124181,I124003);
nand I_7130 (I123932,I124181,I124102);
DFFARX1 I_7131 (I124226,I105897,I2966,I123952,);
and I_7132 (I124243,I124226,I105906);
DFFARX1 I_7133 (I124260,I124243,I2966,I123952,);
not I_7134 (I123923,I124260);
nand I_7135 (I124291,I124243,I124181);
and I_7136 (I124308,I124003,I124291);
DFFARX1 I_7137 (I123914,I124308,I2966,I123952,);
DFFARX1 I_7138 (I124339,I105894,I2966,I123952,);
nand I_7139 (I124356,I124339,I124003);
and I_7140 (I124373,I124181,I124356);
DFFARX1 I_7141 (I123944,I124373,I2966,I123952,);
not I_7142 (I124404,I124339);
nor I_7143 (I124421,I124020,I124404);
and I_7144 (I124438,I124339,I124421);
or I_7145 (I124455,I124243,I124438);
DFFARX1 I_7146 (I123929,I124455,I2966,I123952,);
nand I_7147 (I123926,I124339,I124085);
DFFARX1 I_7148 (I123917,I124339,I2966,I123952,);
not I_7149 (I124547,I2973);
nand I_7150 (I124564,I119189,I119201);
and I_7151 (I124581,I124564,I119183);
DFFARX1 I_7152 (I124598,I124581,I2966,I124547,);
nor I_7153 (I124615,I119195,I119201);
nor I_7154 (I124632,I124615,I124598);
not I_7155 (I124530,I124615);
DFFARX1 I_7156 (I124663,I119180,I2966,I124547,);
not I_7157 (I124680,I124663);
nor I_7158 (I124697,I124615,I124680);
nand I_7159 (I124533,I124663,I124632);
DFFARX1 I_7160 (I124515,I124663,I2966,I124547,);
nand I_7161 (I124742,I119171,I119186);
and I_7162 (I124759,I124742,I119177);
DFFARX1 I_7163 (I124776,I124759,I2966,I124547,);
nor I_7164 (I124536,I124776,I124598);
nand I_7165 (I124527,I124776,I124697);
DFFARX1 I_7166 (I124821,I119198,I2966,I124547,);
and I_7167 (I124838,I124821,I119192);
DFFARX1 I_7168 (I124855,I124838,I2966,I124547,);
not I_7169 (I124518,I124855);
nand I_7170 (I124886,I124838,I124776);
and I_7171 (I124903,I124598,I124886);
DFFARX1 I_7172 (I124509,I124903,I2966,I124547,);
DFFARX1 I_7173 (I124934,I119174,I2966,I124547,);
nand I_7174 (I124951,I124934,I124598);
and I_7175 (I124968,I124776,I124951);
DFFARX1 I_7176 (I124539,I124968,I2966,I124547,);
not I_7177 (I124999,I124934);
nor I_7178 (I125016,I124615,I124999);
and I_7179 (I125033,I124934,I125016);
or I_7180 (I125050,I124838,I125033);
DFFARX1 I_7181 (I124524,I125050,I2966,I124547,);
nand I_7182 (I124521,I124934,I124680);
DFFARX1 I_7183 (I124512,I124934,I2966,I124547,);
not I_7184 (I125142,I2973);
nand I_7185 (I125159,I112085,I112106);
and I_7186 (I125176,I125159,I112091);
DFFARX1 I_7187 (I125193,I125176,I2966,I125142,);
nor I_7188 (I125210,I112109,I112106);
DFFARX1 I_7189 (I125227,I112112,I2966,I125142,);
nand I_7190 (I125244,I125227,I125210);
DFFARX1 I_7191 (I125113,I125227,I2966,I125142,);
nand I_7192 (I125275,I112082,I112094);
and I_7193 (I125292,I125275,I112103);
DFFARX1 I_7194 (I125309,I125292,I2966,I125142,);
not I_7195 (I125326,I125309);
nor I_7196 (I125343,I125193,I125326);
and I_7197 (I125360,I125210,I125343);
and I_7198 (I125377,I125309,I125244);
DFFARX1 I_7199 (I125110,I125377,I2966,I125142,);
DFFARX1 I_7200 (I125104,I125309,I2966,I125142,);
DFFARX1 I_7201 (I125422,I112097,I2966,I125142,);
and I_7202 (I125439,I125422,I112100);
nand I_7203 (I125456,I125439,I125309);
nor I_7204 (I125131,I125439,I125210);
not I_7205 (I125487,I125439);
nor I_7206 (I125504,I125193,I125487);
nand I_7207 (I125122,I125227,I125504);
nand I_7208 (I125116,I125309,I125487);
or I_7209 (I125549,I125439,I125360);
DFFARX1 I_7210 (I125119,I125549,I2966,I125142,);
DFFARX1 I_7211 (I125580,I112088,I2966,I125142,);
and I_7212 (I125597,I125580,I125456);
DFFARX1 I_7213 (I125134,I125597,I2966,I125142,);
nor I_7214 (I125628,I125580,I125193);
nand I_7215 (I125128,I125439,I125628);
not I_7216 (I125125,I125580);
DFFARX1 I_7217 (I125673,I125580,I2966,I125142,);
and I_7218 (I125107,I125580,I125673);
not I_7219 (I125737,I2973);
nand I_7220 (I125754,I106523,I106526);
and I_7221 (I125771,I125754,I106535);
DFFARX1 I_7222 (I125788,I125771,I2966,I125737,);
nor I_7223 (I125805,I106529,I106526);
DFFARX1 I_7224 (I125822,I106550,I2966,I125737,);
nand I_7225 (I125839,I125822,I125805);
DFFARX1 I_7226 (I125708,I125822,I2966,I125737,);
nand I_7227 (I125870,I106547,I106553);
and I_7228 (I125887,I125870,I106538);
DFFARX1 I_7229 (I125904,I125887,I2966,I125737,);
not I_7230 (I125921,I125904);
nor I_7231 (I125938,I125788,I125921);
and I_7232 (I125955,I125805,I125938);
and I_7233 (I125972,I125904,I125839);
DFFARX1 I_7234 (I125705,I125972,I2966,I125737,);
DFFARX1 I_7235 (I125699,I125904,I2966,I125737,);
DFFARX1 I_7236 (I126017,I106541,I2966,I125737,);
and I_7237 (I126034,I126017,I106544);
nand I_7238 (I126051,I126034,I125904);
nor I_7239 (I125726,I126034,I125805);
not I_7240 (I126082,I126034);
nor I_7241 (I126099,I125788,I126082);
nand I_7242 (I125717,I125822,I126099);
nand I_7243 (I125711,I125904,I126082);
or I_7244 (I126144,I126034,I125955);
DFFARX1 I_7245 (I125714,I126144,I2966,I125737,);
DFFARX1 I_7246 (I126175,I106532,I2966,I125737,);
and I_7247 (I126192,I126175,I126051);
DFFARX1 I_7248 (I125729,I126192,I2966,I125737,);
nor I_7249 (I126223,I126175,I125788);
nand I_7250 (I125723,I126034,I126223);
not I_7251 (I125720,I126175);
DFFARX1 I_7252 (I126268,I126175,I2966,I125737,);
and I_7253 (I125702,I126175,I126268);
not I_7254 (I126332,I2973);
nand I_7255 (I126349,I116549,I116519);
and I_7256 (I126366,I126349,I116537);
DFFARX1 I_7257 (I126383,I126366,I2966,I126332,);
nor I_7258 (I126400,I116531,I116519);
DFFARX1 I_7259 (I126417,I116528,I2966,I126332,);
nand I_7260 (I126434,I126417,I126400);
DFFARX1 I_7261 (I126303,I126417,I2966,I126332,);
nand I_7262 (I126465,I116522,I116525);
and I_7263 (I126482,I126465,I116543);
DFFARX1 I_7264 (I126499,I126482,I2966,I126332,);
not I_7265 (I126516,I126499);
nor I_7266 (I126533,I126383,I126516);
and I_7267 (I126550,I126400,I126533);
and I_7268 (I126567,I126499,I126434);
DFFARX1 I_7269 (I126300,I126567,I2966,I126332,);
DFFARX1 I_7270 (I126294,I126499,I2966,I126332,);
DFFARX1 I_7271 (I126612,I116546,I2966,I126332,);
and I_7272 (I126629,I126612,I116540);
nand I_7273 (I126646,I126629,I126499);
nor I_7274 (I126321,I126629,I126400);
not I_7275 (I126677,I126629);
nor I_7276 (I126694,I126383,I126677);
nand I_7277 (I126312,I126417,I126694);
nand I_7278 (I126306,I126499,I126677);
or I_7279 (I126739,I126629,I126550);
DFFARX1 I_7280 (I126309,I126739,I2966,I126332,);
DFFARX1 I_7281 (I126770,I116534,I2966,I126332,);
and I_7282 (I126787,I126770,I126646);
DFFARX1 I_7283 (I126324,I126787,I2966,I126332,);
nor I_7284 (I126818,I126770,I126383);
nand I_7285 (I126318,I126629,I126818);
not I_7286 (I126315,I126770);
DFFARX1 I_7287 (I126863,I126770,I2966,I126332,);
and I_7288 (I126297,I126770,I126863);
not I_7289 (I126927,I2973);
not I_7290 (I126944,I107107);
nor I_7291 (I126961,I107131,I107116);
nand I_7292 (I126978,I126961,I107101);
nor I_7293 (I126995,I126944,I107131);
nand I_7294 (I127012,I126995,I107128);
not I_7295 (I127029,I107131);
not I_7296 (I127046,I127029);
not I_7297 (I127063,I107110);
nor I_7298 (I127080,I127063,I107104);
and I_7299 (I127097,I127080,I107125);
or I_7300 (I127114,I127097,I107113);
DFFARX1 I_7301 (I127131,I127114,I2966,I126927,);
nand I_7302 (I127148,I126944,I107110);
or I_7303 (I126916,I127148,I127131);
not I_7304 (I127179,I127148);
nor I_7305 (I127196,I127131,I127179);
and I_7306 (I127213,I127029,I127196);
nand I_7307 (I126889,I127148,I127046);
DFFARX1 I_7308 (I127244,I107122,I2966,I126927,);
or I_7309 (I126910,I127244,I127131);
nor I_7310 (I127275,I127244,I127012);
nor I_7311 (I127292,I127244,I127046);
nand I_7312 (I126895,I126978,I127292);
or I_7313 (I127323,I127244,I127213);
DFFARX1 I_7314 (I126892,I127323,I2966,I126927,);
not I_7315 (I126898,I127244);
DFFARX1 I_7316 (I127368,I107119,I2966,I126927,);
not I_7317 (I127385,I127368);
nor I_7318 (I127402,I127385,I126978);
DFFARX1 I_7319 (I126904,I127402,I2966,I126927,);
nor I_7320 (I126919,I127244,I127385);
nor I_7321 (I126907,I127385,I127148);
not I_7322 (I127461,I127385);
and I_7323 (I127478,I127012,I127461);
nor I_7324 (I126913,I127148,I127478);
nand I_7325 (I126901,I127385,I127275);
not I_7326 (I127556,I2973);
nand I_7327 (I127573,I123340,I123322);
and I_7328 (I127590,I127573,I123337);
DFFARX1 I_7329 (I127607,I127590,I2966,I127556,);
not I_7330 (I127545,I127607);
DFFARX1 I_7331 (I127638,I127607,I2966,I127556,);
not I_7332 (I127533,I127638);
nor I_7333 (I127669,I123328,I123322);
not I_7334 (I127686,I127669);
nor I_7335 (I127703,I127607,I127686);
DFFARX1 I_7336 (I127720,I123343,I2966,I127556,);
not I_7337 (I127737,I127720);
nand I_7338 (I127536,I127720,I127686);
DFFARX1 I_7339 (I127768,I127720,I2966,I127556,);
and I_7340 (I127521,I127607,I127768);
nand I_7341 (I127799,I123319,I123325);
and I_7342 (I127816,I127799,I123331);
DFFARX1 I_7343 (I127833,I127816,I2966,I127556,);
nor I_7344 (I127850,I127833,I127737);
and I_7345 (I127867,I127669,I127850);
nor I_7346 (I127884,I127833,I127607);
DFFARX1 I_7347 (I127527,I127833,I2966,I127556,);
DFFARX1 I_7348 (I127915,I123346,I2966,I127556,);
and I_7349 (I127932,I127915,I123334);
or I_7350 (I127949,I127932,I127867);
DFFARX1 I_7351 (I127539,I127949,I2966,I127556,);
nand I_7352 (I127548,I127932,I127884);
DFFARX1 I_7353 (I127518,I127932,I2966,I127556,);
DFFARX1 I_7354 (I128008,I123349,I2966,I127556,);
nand I_7355 (I127542,I128008,I127703);
DFFARX1 I_7356 (I127530,I128008,I2966,I127556,);
nand I_7357 (I128053,I128008,I127669);
and I_7358 (I128070,I127720,I128053);
DFFARX1 I_7359 (I127524,I128070,I2966,I127556,);
not I_7360 (I128134,I2973);
nand I_7361 (I128151,I113408,I113438);
and I_7362 (I128168,I128151,I113420);
DFFARX1 I_7363 (I128185,I128168,I2966,I128134,);
not I_7364 (I128123,I128185);
DFFARX1 I_7365 (I128216,I128185,I2966,I128134,);
not I_7366 (I128111,I128216);
nor I_7367 (I128247,I113417,I113438);
not I_7368 (I128264,I128247);
nor I_7369 (I128281,I128185,I128264);
DFFARX1 I_7370 (I128298,I113411,I2966,I128134,);
not I_7371 (I128315,I128298);
nand I_7372 (I128114,I128298,I128264);
DFFARX1 I_7373 (I128346,I128298,I2966,I128134,);
and I_7374 (I128099,I128185,I128346);
nand I_7375 (I128377,I113414,I113429);
and I_7376 (I128394,I128377,I113426);
DFFARX1 I_7377 (I128411,I128394,I2966,I128134,);
nor I_7378 (I128428,I128411,I128315);
and I_7379 (I128445,I128247,I128428);
nor I_7380 (I128462,I128411,I128185);
DFFARX1 I_7381 (I128105,I128411,I2966,I128134,);
DFFARX1 I_7382 (I128493,I113423,I2966,I128134,);
and I_7383 (I128510,I128493,I113435);
or I_7384 (I128527,I128510,I128445);
DFFARX1 I_7385 (I128117,I128527,I2966,I128134,);
nand I_7386 (I128126,I128510,I128462);
DFFARX1 I_7387 (I128096,I128510,I2966,I128134,);
DFFARX1 I_7388 (I128586,I113432,I2966,I128134,);
nand I_7389 (I128120,I128586,I128281);
DFFARX1 I_7390 (I128108,I128586,I2966,I128134,);
nand I_7391 (I128631,I128586,I128247);
and I_7392 (I128648,I128298,I128631);
DFFARX1 I_7393 (I128102,I128648,I2966,I128134,);
not I_7394 (I128712,I2973);
nand I_7395 (I128729,I111419,I111449);
and I_7396 (I128746,I128729,I111431);
DFFARX1 I_7397 (I128763,I128746,I2966,I128712,);
not I_7398 (I128701,I128763);
DFFARX1 I_7399 (I128794,I128763,I2966,I128712,);
not I_7400 (I128689,I128794);
nor I_7401 (I128825,I111428,I111449);
not I_7402 (I128842,I128825);
nor I_7403 (I128859,I128763,I128842);
DFFARX1 I_7404 (I128876,I111422,I2966,I128712,);
not I_7405 (I128893,I128876);
nand I_7406 (I128692,I128876,I128842);
DFFARX1 I_7407 (I128924,I128876,I2966,I128712,);
and I_7408 (I128677,I128763,I128924);
nand I_7409 (I128955,I111425,I111440);
and I_7410 (I128972,I128955,I111437);
DFFARX1 I_7411 (I128989,I128972,I2966,I128712,);
nor I_7412 (I129006,I128989,I128893);
and I_7413 (I129023,I128825,I129006);
nor I_7414 (I129040,I128989,I128763);
DFFARX1 I_7415 (I128683,I128989,I2966,I128712,);
DFFARX1 I_7416 (I129071,I111434,I2966,I128712,);
and I_7417 (I129088,I129071,I111446);
or I_7418 (I129105,I129088,I129023);
DFFARX1 I_7419 (I128695,I129105,I2966,I128712,);
nand I_7420 (I128704,I129088,I129040);
DFFARX1 I_7421 (I128674,I129088,I2966,I128712,);
DFFARX1 I_7422 (I129164,I111443,I2966,I128712,);
nand I_7423 (I128698,I129164,I128859);
DFFARX1 I_7424 (I128686,I129164,I2966,I128712,);
nand I_7425 (I129209,I129164,I128825);
and I_7426 (I129226,I128876,I129209);
DFFARX1 I_7427 (I128680,I129226,I2966,I128712,);
not I_7428 (I129290,I2973);
nand I_7429 (I129307,I126315,I126303);
and I_7430 (I129324,I129307,I126300);
DFFARX1 I_7431 (I129341,I129324,I2966,I129290,);
not I_7432 (I129358,I129341);
nor I_7433 (I129375,I126321,I126303);
or I_7434 (I129273,I129375,I129341);
not I_7435 (I129261,I129375);
DFFARX1 I_7436 (I129420,I126324,I2966,I129290,);
nor I_7437 (I129437,I129420,I129375);
nand I_7438 (I129454,I126294,I126312);
and I_7439 (I129471,I129454,I126309);
DFFARX1 I_7440 (I129488,I129471,I2966,I129290,);
nor I_7441 (I129270,I129488,I129341);
not I_7442 (I129519,I129488);
nor I_7443 (I129536,I129420,I129519);
DFFARX1 I_7444 (I129553,I126318,I2966,I129290,);
and I_7445 (I129570,I129553,I126306);
or I_7446 (I129279,I129570,I129375);
nand I_7447 (I129258,I129570,I129536);
DFFARX1 I_7448 (I129615,I126297,I2966,I129290,);
and I_7449 (I129632,I129615,I129358);
nor I_7450 (I129276,I129570,I129632);
nor I_7451 (I129663,I129615,I129420);
DFFARX1 I_7452 (I129267,I129663,I2966,I129290,);
nor I_7453 (I129282,I129615,I129341);
not I_7454 (I129708,I129615);
nor I_7455 (I129725,I129488,I129708);
and I_7456 (I129742,I129375,I129725);
or I_7457 (I129759,I129570,I129742);
DFFARX1 I_7458 (I129255,I129759,I2966,I129290,);
nand I_7459 (I129264,I129615,I129437);
nand I_7460 (I129252,I129615,I129519);
not I_7461 (I129851,I2973);
nand I_7462 (I129868,I119838,I119832);
and I_7463 (I129885,I129868,I119844);
DFFARX1 I_7464 (I129902,I129885,I2966,I129851,);
not I_7465 (I129919,I129902);
nor I_7466 (I129936,I119841,I119832);
or I_7467 (I129834,I129936,I129902);
not I_7468 (I129822,I129936);
DFFARX1 I_7469 (I129981,I119820,I2966,I129851,);
nor I_7470 (I129998,I129981,I129936);
nand I_7471 (I130015,I119826,I119835);
and I_7472 (I130032,I130015,I119823);
DFFARX1 I_7473 (I130049,I130032,I2966,I129851,);
nor I_7474 (I129831,I130049,I129902);
not I_7475 (I130080,I130049);
nor I_7476 (I130097,I129981,I130080);
DFFARX1 I_7477 (I130114,I119847,I2966,I129851,);
and I_7478 (I130131,I130114,I119817);
or I_7479 (I129840,I130131,I129936);
nand I_7480 (I129819,I130131,I130097);
DFFARX1 I_7481 (I130176,I119829,I2966,I129851,);
and I_7482 (I130193,I130176,I129919);
nor I_7483 (I129837,I130131,I130193);
nor I_7484 (I130224,I130176,I129981);
DFFARX1 I_7485 (I129828,I130224,I2966,I129851,);
nor I_7486 (I129843,I130176,I129902);
not I_7487 (I130269,I130176);
nor I_7488 (I130286,I130049,I130269);
and I_7489 (I130303,I129936,I130286);
or I_7490 (I130320,I130131,I130303);
DFFARX1 I_7491 (I129816,I130320,I2966,I129851,);
nand I_7492 (I129825,I130176,I129998);
nand I_7493 (I129813,I130176,I130080);
not I_7494 (I130412,I2973);
nand I_7495 (I130429,I118532,I118523);
and I_7496 (I130446,I130429,I118538);
DFFARX1 I_7497 (I130463,I130446,I2966,I130412,);
not I_7498 (I130480,I130463);
nor I_7499 (I130497,I118508,I118523);
or I_7500 (I130395,I130497,I130463);
not I_7501 (I130383,I130497);
DFFARX1 I_7502 (I130542,I118511,I2966,I130412,);
nor I_7503 (I130559,I130542,I130497);
nand I_7504 (I130576,I118529,I118526);
and I_7505 (I130593,I130576,I118514);
DFFARX1 I_7506 (I130610,I130593,I2966,I130412,);
nor I_7507 (I130392,I130610,I130463);
not I_7508 (I130641,I130610);
nor I_7509 (I130658,I130542,I130641);
DFFARX1 I_7510 (I130675,I118535,I2966,I130412,);
and I_7511 (I130692,I130675,I118520);
or I_7512 (I130401,I130692,I130497);
nand I_7513 (I130380,I130692,I130658);
DFFARX1 I_7514 (I130737,I118517,I2966,I130412,);
and I_7515 (I130754,I130737,I130480);
nor I_7516 (I130398,I130692,I130754);
nor I_7517 (I130785,I130737,I130542);
DFFARX1 I_7518 (I130389,I130785,I2966,I130412,);
nor I_7519 (I130404,I130737,I130463);
not I_7520 (I130830,I130737);
nor I_7521 (I130847,I130610,I130830);
and I_7522 (I130864,I130497,I130847);
or I_7523 (I130881,I130692,I130864);
DFFARX1 I_7524 (I130377,I130881,I2966,I130412,);
nand I_7525 (I130386,I130737,I130559);
nand I_7526 (I130374,I130737,I130641);
not I_7527 (I130973,I2973);
not I_7528 (I130990,I125714);
nor I_7529 (I131007,I125699,I125726);
nand I_7530 (I131024,I131007,I125702);
DFFARX1 I_7531 (I130947,I131024,I2966,I130973,);
nor I_7532 (I131055,I130990,I125699);
nand I_7533 (I131072,I131055,I125717);
not I_7534 (I130962,I131072);
DFFARX1 I_7535 (I130944,I131072,I2966,I130973,);
not I_7536 (I131117,I125699);
not I_7537 (I131134,I131117);
not I_7538 (I131151,I125729);
nor I_7539 (I131168,I131151,I125711);
and I_7540 (I131185,I131168,I125720);
or I_7541 (I131202,I131185,I125705);
DFFARX1 I_7542 (I131219,I131202,I2966,I130973,);
nor I_7543 (I131236,I131219,I131072);
nor I_7544 (I131253,I131219,I131134);
nand I_7545 (I130959,I131024,I131253);
nand I_7546 (I131284,I130990,I125729);
nand I_7547 (I131301,I131284,I131219);
and I_7548 (I131318,I131284,I131301);
DFFARX1 I_7549 (I130941,I131318,I2966,I130973,);
DFFARX1 I_7550 (I131349,I131284,I2966,I130973,);
and I_7551 (I130938,I131117,I131349);
DFFARX1 I_7552 (I131380,I125708,I2966,I130973,);
not I_7553 (I131397,I131380);
nor I_7554 (I131414,I131072,I131397);
and I_7555 (I131431,I131380,I131414);
nand I_7556 (I130953,I131380,I131134);
DFFARX1 I_7557 (I131462,I131380,I2966,I130973,);
not I_7558 (I130950,I131462);
DFFARX1 I_7559 (I131493,I125723,I2966,I130973,);
not I_7560 (I131510,I131493);
or I_7561 (I131527,I131510,I131431);
DFFARX1 I_7562 (I130956,I131527,I2966,I130973,);
nand I_7563 (I130965,I131510,I131236);
DFFARX1 I_7564 (I130935,I131510,I2966,I130973,);
not I_7565 (I131619,I2973);
not I_7566 (I131636,I115273);
nor I_7567 (I131653,I115267,I115285);
nand I_7568 (I131670,I131653,I115261);
DFFARX1 I_7569 (I131590,I131670,I2966,I131619,);
nor I_7570 (I131701,I131636,I115267);
nand I_7571 (I131718,I131701,I115276);
nand I_7572 (I131735,I131718,I131670);
not I_7573 (I131752,I115267);
not I_7574 (I131769,I115291);
nor I_7575 (I131786,I131769,I115282);
and I_7576 (I131803,I131786,I115270);
or I_7577 (I131820,I131803,I115288);
DFFARX1 I_7578 (I131837,I131820,I2966,I131619,);
nor I_7579 (I131854,I131837,I131718);
nand I_7580 (I131605,I131752,I131854);
not I_7581 (I131602,I131837);
and I_7582 (I131899,I131837,I131735);
DFFARX1 I_7583 (I131587,I131899,I2966,I131619,);
DFFARX1 I_7584 (I131930,I131837,I2966,I131619,);
and I_7585 (I131584,I131752,I131930);
nand I_7586 (I131961,I131636,I115291);
not I_7587 (I131978,I131961);
nor I_7588 (I131995,I131837,I131978);
DFFARX1 I_7589 (I132012,I115279,I2966,I131619,);
nand I_7590 (I132029,I132012,I131961);
and I_7591 (I132046,I131752,I132029);
DFFARX1 I_7592 (I131611,I132046,I2966,I131619,);
not I_7593 (I132077,I132012);
nand I_7594 (I131599,I132012,I131995);
nand I_7595 (I131593,I132012,I131978);
DFFARX1 I_7596 (I132122,I115264,I2966,I131619,);
not I_7597 (I132139,I132122);
nor I_7598 (I131608,I132012,I132139);
nor I_7599 (I132170,I132139,I132077);
and I_7600 (I132187,I131718,I132170);
or I_7601 (I132204,I131961,I132187);
DFFARX1 I_7602 (I131596,I132204,I2966,I131619,);
DFFARX1 I_7603 (I131581,I132139,I2966,I131619,);
not I_7604 (I132282,I2973);
not I_7605 (I132299,I125110);
nor I_7606 (I132316,I125125,I125107);
nand I_7607 (I132333,I132316,I125119);
DFFARX1 I_7608 (I132253,I132333,I2966,I132282,);
nor I_7609 (I132364,I132299,I125125);
nand I_7610 (I132381,I132364,I125116);
nand I_7611 (I132398,I132381,I132333);
not I_7612 (I132415,I125125);
not I_7613 (I132432,I125134);
nor I_7614 (I132449,I132432,I125104);
and I_7615 (I132466,I132449,I125113);
or I_7616 (I132483,I132466,I125131);
DFFARX1 I_7617 (I132500,I132483,I2966,I132282,);
nor I_7618 (I132517,I132500,I132381);
nand I_7619 (I132268,I132415,I132517);
not I_7620 (I132265,I132500);
and I_7621 (I132562,I132500,I132398);
DFFARX1 I_7622 (I132250,I132562,I2966,I132282,);
DFFARX1 I_7623 (I132593,I132500,I2966,I132282,);
and I_7624 (I132247,I132415,I132593);
nand I_7625 (I132624,I132299,I125134);
not I_7626 (I132641,I132624);
nor I_7627 (I132658,I132500,I132641);
DFFARX1 I_7628 (I132675,I125122,I2966,I132282,);
nand I_7629 (I132692,I132675,I132624);
and I_7630 (I132709,I132415,I132692);
DFFARX1 I_7631 (I132274,I132709,I2966,I132282,);
not I_7632 (I132740,I132675);
nand I_7633 (I132262,I132675,I132658);
nand I_7634 (I132256,I132675,I132641);
DFFARX1 I_7635 (I132785,I125128,I2966,I132282,);
not I_7636 (I132802,I132785);
nor I_7637 (I132271,I132675,I132802);
nor I_7638 (I132833,I132802,I132740);
and I_7639 (I132850,I132381,I132833);
or I_7640 (I132867,I132624,I132850);
DFFARX1 I_7641 (I132259,I132867,I2966,I132282,);
DFFARX1 I_7642 (I132244,I132802,I2966,I132282,);
not I_7643 (I132945,I2973);
not I_7644 (I132962,I130389);
nor I_7645 (I132979,I130377,I130380);
nand I_7646 (I132996,I132979,I130395);
DFFARX1 I_7647 (I132916,I132996,I2966,I132945,);
nor I_7648 (I133027,I132962,I130377);
nand I_7649 (I133044,I133027,I130386);
nand I_7650 (I133061,I133044,I132996);
not I_7651 (I133078,I130377);
not I_7652 (I133095,I130398);
nor I_7653 (I133112,I133095,I130374);
and I_7654 (I133129,I133112,I130383);
or I_7655 (I133146,I133129,I130392);
DFFARX1 I_7656 (I133163,I133146,I2966,I132945,);
nor I_7657 (I133180,I133163,I133044);
nand I_7658 (I132931,I133078,I133180);
not I_7659 (I132928,I133163);
and I_7660 (I133225,I133163,I133061);
DFFARX1 I_7661 (I132913,I133225,I2966,I132945,);
DFFARX1 I_7662 (I133256,I133163,I2966,I132945,);
and I_7663 (I132910,I133078,I133256);
nand I_7664 (I133287,I132962,I130398);
not I_7665 (I133304,I133287);
nor I_7666 (I133321,I133163,I133304);
DFFARX1 I_7667 (I133338,I130404,I2966,I132945,);
nand I_7668 (I133355,I133338,I133287);
and I_7669 (I133372,I133078,I133355);
DFFARX1 I_7670 (I132937,I133372,I2966,I132945,);
not I_7671 (I133403,I133338);
nand I_7672 (I132925,I133338,I133321);
nand I_7673 (I132919,I133338,I133304);
DFFARX1 I_7674 (I133448,I130401,I2966,I132945,);
not I_7675 (I133465,I133448);
nor I_7676 (I132934,I133338,I133465);
nor I_7677 (I133496,I133465,I133403);
and I_7678 (I133513,I133044,I133496);
or I_7679 (I133530,I133287,I133513);
DFFARX1 I_7680 (I132922,I133530,I2966,I132945,);
DFFARX1 I_7681 (I132907,I133465,I2966,I132945,);
not I_7682 (I133608,I2973);
or I_7683 (I133625,I127518,I127536);
or I_7684 (I133642,I127521,I127518);
DFFARX1 I_7685 (I133582,I133642,I2966,I133608,);
nor I_7686 (I133673,I127530,I127533);
not I_7687 (I133690,I133673);
not I_7688 (I133707,I127530);
and I_7689 (I133724,I133707,I127539);
nor I_7690 (I133741,I133724,I127536);
nor I_7691 (I133758,I127545,I127524);
DFFARX1 I_7692 (I133775,I133758,I2966,I133608,);
nand I_7693 (I133792,I133775,I133625);
and I_7694 (I133809,I133741,I133792);
DFFARX1 I_7695 (I133576,I133809,I2966,I133608,);
nor I_7696 (I133840,I127545,I127521);
DFFARX1 I_7697 (I133857,I133840,I2966,I133608,);
and I_7698 (I133573,I133673,I133857);
DFFARX1 I_7699 (I133888,I127548,I2966,I133608,);
and I_7700 (I133905,I133888,I127542);
DFFARX1 I_7701 (I133922,I133905,I2966,I133608,);
not I_7702 (I133585,I133922);
DFFARX1 I_7703 (I133570,I133905,I2966,I133608,);
DFFARX1 I_7704 (I133967,I127527,I2966,I133608,);
not I_7705 (I133984,I133967);
nor I_7706 (I134001,I133642,I133984);
and I_7707 (I134018,I133905,I134001);
or I_7708 (I134035,I133625,I134018);
DFFARX1 I_7709 (I133591,I134035,I2966,I133608,);
nor I_7710 (I134066,I133967,I133775);
nand I_7711 (I133600,I133741,I134066);
nor I_7712 (I134097,I133967,I133690);
nand I_7713 (I133594,I133840,I134097);
not I_7714 (I133597,I133967);
nand I_7715 (I133588,I133967,I133690);
DFFARX1 I_7716 (I133579,I133967,I2966,I133608,);
not I_7717 (I134203,I2973);
or I_7718 (I134220,I129834,I129843);
or I_7719 (I134237,I129837,I129834);
DFFARX1 I_7720 (I134177,I134237,I2966,I134203,);
nor I_7721 (I134268,I129813,I129816);
not I_7722 (I134285,I134268);
not I_7723 (I134302,I129813);
and I_7724 (I134319,I134302,I129825);
nor I_7725 (I134336,I134319,I129843);
nor I_7726 (I134353,I129831,I129822);
DFFARX1 I_7727 (I134370,I134353,I2966,I134203,);
nand I_7728 (I134387,I134370,I134220);
and I_7729 (I134404,I134336,I134387);
DFFARX1 I_7730 (I134171,I134404,I2966,I134203,);
nor I_7731 (I134435,I129831,I129837);
DFFARX1 I_7732 (I134452,I134435,I2966,I134203,);
and I_7733 (I134168,I134268,I134452);
DFFARX1 I_7734 (I134483,I129828,I2966,I134203,);
and I_7735 (I134500,I134483,I129819);
DFFARX1 I_7736 (I134517,I134500,I2966,I134203,);
not I_7737 (I134180,I134517);
DFFARX1 I_7738 (I134165,I134500,I2966,I134203,);
DFFARX1 I_7739 (I134562,I129840,I2966,I134203,);
not I_7740 (I134579,I134562);
nor I_7741 (I134596,I134237,I134579);
and I_7742 (I134613,I134500,I134596);
or I_7743 (I134630,I134220,I134613);
DFFARX1 I_7744 (I134186,I134630,I2966,I134203,);
nor I_7745 (I134661,I134562,I134370);
nand I_7746 (I134195,I134336,I134661);
nor I_7747 (I134692,I134562,I134285);
nand I_7748 (I134189,I134435,I134692);
not I_7749 (I134192,I134562);
nand I_7750 (I134183,I134562,I134285);
DFFARX1 I_7751 (I134174,I134562,I2966,I134203,);
not I_7752 (I134798,I2973);
not I_7753 (I134815,I128686);
nor I_7754 (I134832,I128677,I128683);
nand I_7755 (I134849,I134832,I128695);
nor I_7756 (I134866,I134815,I128677);
nand I_7757 (I134883,I134866,I128680);
not I_7758 (I134900,I134883);
not I_7759 (I134917,I128677);
nor I_7760 (I134787,I134883,I134917);
not I_7761 (I134948,I134917);
nand I_7762 (I134772,I134883,I134948);
not I_7763 (I134979,I128704);
nor I_7764 (I134996,I134979,I128698);
and I_7765 (I135013,I134996,I128689);
or I_7766 (I135030,I135013,I128674);
DFFARX1 I_7767 (I135047,I135030,I2966,I134798,);
nor I_7768 (I135064,I135047,I134900);
DFFARX1 I_7769 (I135081,I135047,I2966,I134798,);
not I_7770 (I134769,I135081);
nand I_7771 (I135112,I134815,I128704);
and I_7772 (I135129,I135112,I135064);
DFFARX1 I_7773 (I134766,I135112,I2966,I134798,);
DFFARX1 I_7774 (I135160,I128692,I2966,I134798,);
nor I_7775 (I135177,I135160,I134883);
nand I_7776 (I134784,I135047,I135177);
nor I_7777 (I135208,I135160,I134948);
not I_7778 (I134781,I135160);
nand I_7779 (I135239,I135160,I134849);
and I_7780 (I135256,I134917,I135239);
DFFARX1 I_7781 (I134760,I135256,I2966,I134798,);
DFFARX1 I_7782 (I134763,I135160,I2966,I134798,);
DFFARX1 I_7783 (I135301,I128701,I2966,I134798,);
not I_7784 (I135318,I135301);
nand I_7785 (I135335,I135318,I134883);
and I_7786 (I135352,I135112,I135335);
DFFARX1 I_7787 (I134790,I135352,I2966,I134798,);
or I_7788 (I135383,I135318,I135129);
DFFARX1 I_7789 (I134775,I135383,I2966,I134798,);
nand I_7790 (I134778,I135318,I135208);
not I_7791 (I135461,I2973);
not I_7792 (I135478,I126895);
nor I_7793 (I135495,I126913,I126904);
nand I_7794 (I135512,I135495,I126910);
nor I_7795 (I135529,I135478,I126913);
nand I_7796 (I135546,I135529,I126916);
not I_7797 (I135563,I135546);
not I_7798 (I135580,I126913);
nor I_7799 (I135450,I135546,I135580);
not I_7800 (I135611,I135580);
nand I_7801 (I135435,I135546,I135611);
not I_7802 (I135642,I126892);
nor I_7803 (I135659,I135642,I126907);
and I_7804 (I135676,I135659,I126889);
or I_7805 (I135693,I135676,I126898);
DFFARX1 I_7806 (I135710,I135693,I2966,I135461,);
nor I_7807 (I135727,I135710,I135563);
DFFARX1 I_7808 (I135744,I135710,I2966,I135461,);
not I_7809 (I135432,I135744);
nand I_7810 (I135775,I135478,I126892);
and I_7811 (I135792,I135775,I135727);
DFFARX1 I_7812 (I135429,I135775,I2966,I135461,);
DFFARX1 I_7813 (I135823,I126901,I2966,I135461,);
nor I_7814 (I135840,I135823,I135546);
nand I_7815 (I135447,I135710,I135840);
nor I_7816 (I135871,I135823,I135611);
not I_7817 (I135444,I135823);
nand I_7818 (I135902,I135823,I135512);
and I_7819 (I135919,I135580,I135902);
DFFARX1 I_7820 (I135423,I135919,I2966,I135461,);
DFFARX1 I_7821 (I135426,I135823,I2966,I135461,);
DFFARX1 I_7822 (I135964,I126919,I2966,I135461,);
not I_7823 (I135981,I135964);
nand I_7824 (I135998,I135981,I135546);
and I_7825 (I136015,I135775,I135998);
DFFARX1 I_7826 (I135453,I136015,I2966,I135461,);
or I_7827 (I136046,I135981,I135792);
DFFARX1 I_7828 (I135438,I136046,I2966,I135461,);
nand I_7829 (I135441,I135981,I135871);
not I_7830 (I136124,I2973);
not I_7831 (I136141,I122178);
nor I_7832 (I136158,I122190,I122172);
nand I_7833 (I136175,I136158,I122193);
nor I_7834 (I136192,I136141,I122190);
nand I_7835 (I136209,I136192,I122184);
not I_7836 (I136226,I136209);
not I_7837 (I136243,I122190);
nor I_7838 (I136113,I136209,I136243);
not I_7839 (I136274,I136243);
nand I_7840 (I136098,I136209,I136274);
not I_7841 (I136305,I122175);
nor I_7842 (I136322,I136305,I122169);
and I_7843 (I136339,I136322,I122181);
or I_7844 (I136356,I136339,I122166);
DFFARX1 I_7845 (I136373,I136356,I2966,I136124,);
nor I_7846 (I136390,I136373,I136226);
DFFARX1 I_7847 (I136407,I136373,I2966,I136124,);
not I_7848 (I136095,I136407);
nand I_7849 (I136438,I136141,I122175);
and I_7850 (I136455,I136438,I136390);
DFFARX1 I_7851 (I136092,I136438,I2966,I136124,);
DFFARX1 I_7852 (I136486,I122163,I2966,I136124,);
nor I_7853 (I136503,I136486,I136209);
nand I_7854 (I136110,I136373,I136503);
nor I_7855 (I136534,I136486,I136274);
not I_7856 (I136107,I136486);
nand I_7857 (I136565,I136486,I136175);
and I_7858 (I136582,I136243,I136565);
DFFARX1 I_7859 (I136086,I136582,I2966,I136124,);
DFFARX1 I_7860 (I136089,I136486,I2966,I136124,);
DFFARX1 I_7861 (I136627,I122187,I2966,I136124,);
not I_7862 (I136644,I136627);
nand I_7863 (I136661,I136644,I136209);
and I_7864 (I136678,I136438,I136661);
DFFARX1 I_7865 (I136116,I136678,I2966,I136124,);
or I_7866 (I136709,I136644,I136455);
DFFARX1 I_7867 (I136101,I136709,I2966,I136124,);
nand I_7868 (I136104,I136644,I136534);
not I_7869 (I136787,I2973);
not I_7870 (I136804,I131584);
nor I_7871 (I136821,I131590,I131596);
nand I_7872 (I136838,I136821,I131599);
nor I_7873 (I136855,I136804,I131590);
nand I_7874 (I136872,I136855,I131581);
not I_7875 (I136889,I136872);
not I_7876 (I136906,I131590);
nor I_7877 (I136776,I136872,I136906);
not I_7878 (I136937,I136906);
nand I_7879 (I136761,I136872,I136937);
not I_7880 (I136968,I131593);
nor I_7881 (I136985,I136968,I131587);
and I_7882 (I137002,I136985,I131602);
or I_7883 (I137019,I137002,I131608);
DFFARX1 I_7884 (I137036,I137019,I2966,I136787,);
nor I_7885 (I137053,I137036,I136889);
DFFARX1 I_7886 (I137070,I137036,I2966,I136787,);
not I_7887 (I136758,I137070);
nand I_7888 (I137101,I136804,I131593);
and I_7889 (I137118,I137101,I137053);
DFFARX1 I_7890 (I136755,I137101,I2966,I136787,);
DFFARX1 I_7891 (I137149,I131605,I2966,I136787,);
nor I_7892 (I137166,I137149,I136872);
nand I_7893 (I136773,I137036,I137166);
nor I_7894 (I137197,I137149,I136937);
not I_7895 (I136770,I137149);
nand I_7896 (I137228,I137149,I136838);
and I_7897 (I137245,I136906,I137228);
DFFARX1 I_7898 (I136749,I137245,I2966,I136787,);
DFFARX1 I_7899 (I136752,I137149,I2966,I136787,);
DFFARX1 I_7900 (I137290,I131611,I2966,I136787,);
not I_7901 (I137307,I137290);
nand I_7902 (I137324,I137307,I136872);
and I_7903 (I137341,I137101,I137324);
DFFARX1 I_7904 (I136779,I137341,I2966,I136787,);
or I_7905 (I137372,I137307,I137118);
DFFARX1 I_7906 (I136764,I137372,I2966,I136787,);
nand I_7907 (I136767,I137307,I137197);
not I_7908 (I137450,I2973);
not I_7909 (I137467,I120444);
nor I_7910 (I137484,I120456,I120438);
nand I_7911 (I137501,I137484,I120459);
nor I_7912 (I137518,I137467,I120456);
nand I_7913 (I137535,I137518,I120450);
not I_7914 (I137552,I137535);
not I_7915 (I137569,I120456);
nor I_7916 (I137439,I137535,I137569);
not I_7917 (I137600,I137569);
nand I_7918 (I137424,I137535,I137600);
not I_7919 (I137631,I120441);
nor I_7920 (I137648,I137631,I120435);
and I_7921 (I137665,I137648,I120447);
or I_7922 (I137682,I137665,I120432);
DFFARX1 I_7923 (I137699,I137682,I2966,I137450,);
nor I_7924 (I137716,I137699,I137552);
DFFARX1 I_7925 (I137733,I137699,I2966,I137450,);
not I_7926 (I137421,I137733);
nand I_7927 (I137764,I137467,I120441);
and I_7928 (I137781,I137764,I137716);
DFFARX1 I_7929 (I137418,I137764,I2966,I137450,);
DFFARX1 I_7930 (I137812,I120429,I2966,I137450,);
nor I_7931 (I137829,I137812,I137535);
nand I_7932 (I137436,I137699,I137829);
nor I_7933 (I137860,I137812,I137600);
not I_7934 (I137433,I137812);
nand I_7935 (I137891,I137812,I137501);
and I_7936 (I137908,I137569,I137891);
DFFARX1 I_7937 (I137412,I137908,I2966,I137450,);
DFFARX1 I_7938 (I137415,I137812,I2966,I137450,);
DFFARX1 I_7939 (I137953,I120453,I2966,I137450,);
not I_7940 (I137970,I137953);
nand I_7941 (I137987,I137970,I137535);
and I_7942 (I138004,I137764,I137987);
DFFARX1 I_7943 (I137442,I138004,I2966,I137450,);
or I_7944 (I138035,I137970,I137781);
DFFARX1 I_7945 (I137427,I138035,I2966,I137450,);
nand I_7946 (I137430,I137970,I137860);
not I_7947 (I138113,I2973);
not I_7948 (I138130,I130941);
nor I_7949 (I138147,I130938,I130962);
nand I_7950 (I138164,I138147,I130959);
nor I_7951 (I138181,I138130,I130938);
nand I_7952 (I138198,I138181,I130965);
not I_7953 (I138215,I138198);
not I_7954 (I138232,I130938);
nor I_7955 (I138102,I138198,I138232);
not I_7956 (I138263,I138232);
nand I_7957 (I138087,I138198,I138263);
not I_7958 (I138294,I130956);
nor I_7959 (I138311,I138294,I130947);
and I_7960 (I138328,I138311,I130944);
or I_7961 (I138345,I138328,I130953);
DFFARX1 I_7962 (I138362,I138345,I2966,I138113,);
nor I_7963 (I138379,I138362,I138215);
DFFARX1 I_7964 (I138396,I138362,I2966,I138113,);
not I_7965 (I138084,I138396);
nand I_7966 (I138427,I138130,I130956);
and I_7967 (I138444,I138427,I138379);
DFFARX1 I_7968 (I138081,I138427,I2966,I138113,);
DFFARX1 I_7969 (I138475,I130935,I2966,I138113,);
nor I_7970 (I138492,I138475,I138198);
nand I_7971 (I138099,I138362,I138492);
nor I_7972 (I138523,I138475,I138263);
not I_7973 (I138096,I138475);
nand I_7974 (I138554,I138475,I138164);
and I_7975 (I138571,I138232,I138554);
DFFARX1 I_7976 (I138075,I138571,I2966,I138113,);
DFFARX1 I_7977 (I138078,I138475,I2966,I138113,);
DFFARX1 I_7978 (I138616,I130950,I2966,I138113,);
not I_7979 (I138633,I138616);
nand I_7980 (I138650,I138633,I138198);
and I_7981 (I138667,I138427,I138650);
DFFARX1 I_7982 (I138105,I138667,I2966,I138113,);
or I_7983 (I138698,I138633,I138444);
DFFARX1 I_7984 (I138090,I138698,I2966,I138113,);
nand I_7985 (I138093,I138633,I138523);
not I_7986 (I138776,I2973);
not I_7987 (I138793,I135447);
nor I_7988 (I138810,I135426,I135438);
nand I_7989 (I138827,I138810,I135441);
nor I_7990 (I138844,I138793,I135426);
nand I_7991 (I138861,I138844,I135423);
DFFARX1 I_7992 (I138878,I138861,I2966,I138776,);
not I_7993 (I138747,I138878);
not I_7994 (I138909,I135426);
not I_7995 (I138926,I138909);
not I_7996 (I138943,I135444);
nor I_7997 (I138960,I138943,I135435);
and I_7998 (I138977,I138960,I135429);
or I_7999 (I138994,I138977,I135453);
DFFARX1 I_8000 (I139011,I138994,I2966,I138776,);
DFFARX1 I_8001 (I138744,I139011,I2966,I138776,);
DFFARX1 I_8002 (I139042,I139011,I2966,I138776,);
DFFARX1 I_8003 (I138738,I139011,I2966,I138776,);
nand I_8004 (I139073,I138793,I135444);
nand I_8005 (I139090,I139073,I138827);
and I_8006 (I139107,I138909,I139090);
DFFARX1 I_8007 (I138768,I139107,I2966,I138776,);
and I_8008 (I138741,I139073,I139042);
DFFARX1 I_8009 (I139152,I135450,I2966,I138776,);
nor I_8010 (I138765,I139152,I139073);
nor I_8011 (I139183,I139152,I138827);
nand I_8012 (I138762,I138861,I139183);
not I_8013 (I138759,I139152);
DFFARX1 I_8014 (I139228,I135432,I2966,I138776,);
not I_8015 (I139245,I139228);
nor I_8016 (I139262,I139245,I138926);
and I_8017 (I139279,I139152,I139262);
or I_8018 (I139296,I139073,I139279);
DFFARX1 I_8019 (I138753,I139296,I2966,I138776,);
not I_8020 (I139327,I139245);
nor I_8021 (I139344,I139152,I139327);
nand I_8022 (I138756,I139245,I139344);
nand I_8023 (I138750,I138909,I139327);
not I_8024 (I139422,I2973);
not I_8025 (I139439,I124518);
nor I_8026 (I139456,I124530,I124524);
nand I_8027 (I139473,I139456,I124509);
nor I_8028 (I139490,I139439,I124530);
nand I_8029 (I139507,I139490,I124536);
DFFARX1 I_8030 (I139524,I139507,I2966,I139422,);
not I_8031 (I139393,I139524);
not I_8032 (I139555,I124530);
not I_8033 (I139572,I139555);
not I_8034 (I139589,I124533);
nor I_8035 (I139606,I139589,I124515);
and I_8036 (I139623,I139606,I124512);
or I_8037 (I139640,I139623,I124539);
DFFARX1 I_8038 (I139657,I139640,I2966,I139422,);
DFFARX1 I_8039 (I139390,I139657,I2966,I139422,);
DFFARX1 I_8040 (I139688,I139657,I2966,I139422,);
DFFARX1 I_8041 (I139384,I139657,I2966,I139422,);
nand I_8042 (I139719,I139439,I124533);
nand I_8043 (I139736,I139719,I139473);
and I_8044 (I139753,I139555,I139736);
DFFARX1 I_8045 (I139414,I139753,I2966,I139422,);
and I_8046 (I139387,I139719,I139688);
DFFARX1 I_8047 (I139798,I124527,I2966,I139422,);
nor I_8048 (I139411,I139798,I139719);
nor I_8049 (I139829,I139798,I139473);
nand I_8050 (I139408,I139507,I139829);
not I_8051 (I139405,I139798);
DFFARX1 I_8052 (I139874,I124521,I2966,I139422,);
not I_8053 (I139891,I139874);
nor I_8054 (I139908,I139891,I139572);
and I_8055 (I139925,I139798,I139908);
or I_8056 (I139942,I139719,I139925);
DFFARX1 I_8057 (I139399,I139942,I2966,I139422,);
not I_8058 (I139973,I139891);
nor I_8059 (I139990,I139798,I139973);
nand I_8060 (I139402,I139891,I139990);
nand I_8061 (I139396,I139555,I139973);
not I_8062 (I140068,I2973);
not I_8063 (I140085,I132247);
nor I_8064 (I140102,I132268,I132250);
nand I_8065 (I140119,I140102,I132274);
nor I_8066 (I140136,I140085,I132268);
nand I_8067 (I140153,I140136,I132271);
DFFARX1 I_8068 (I140170,I140153,I2966,I140068,);
not I_8069 (I140039,I140170);
not I_8070 (I140201,I132268);
not I_8071 (I140218,I140201);
not I_8072 (I140235,I132265);
nor I_8073 (I140252,I140235,I132244);
and I_8074 (I140269,I140252,I132256);
or I_8075 (I140286,I140269,I132253);
DFFARX1 I_8076 (I140303,I140286,I2966,I140068,);
DFFARX1 I_8077 (I140036,I140303,I2966,I140068,);
DFFARX1 I_8078 (I140334,I140303,I2966,I140068,);
DFFARX1 I_8079 (I140030,I140303,I2966,I140068,);
nand I_8080 (I140365,I140085,I132265);
nand I_8081 (I140382,I140365,I140119);
and I_8082 (I140399,I140201,I140382);
DFFARX1 I_8083 (I140060,I140399,I2966,I140068,);
and I_8084 (I140033,I140365,I140334);
DFFARX1 I_8085 (I140444,I132259,I2966,I140068,);
nor I_8086 (I140057,I140444,I140365);
nor I_8087 (I140475,I140444,I140119);
nand I_8088 (I140054,I140153,I140475);
not I_8089 (I140051,I140444);
DFFARX1 I_8090 (I140520,I132262,I2966,I140068,);
not I_8091 (I140537,I140520);
nor I_8092 (I140554,I140537,I140218);
and I_8093 (I140571,I140444,I140554);
or I_8094 (I140588,I140365,I140571);
DFFARX1 I_8095 (I140045,I140588,I2966,I140068,);
not I_8096 (I140619,I140537);
nor I_8097 (I140636,I140444,I140619);
nand I_8098 (I140048,I140537,I140636);
nand I_8099 (I140042,I140201,I140619);
not I_8100 (I140714,I2973);
nand I_8101 (I140731,I128111,I128123);
and I_8102 (I140748,I140731,I128096);
DFFARX1 I_8103 (I140765,I140748,I2966,I140714,);
not I_8104 (I140782,I140765);
DFFARX1 I_8105 (I140682,I140765,I2966,I140714,);
nor I_8106 (I140813,I128114,I128123);
DFFARX1 I_8107 (I140830,I128105,I2966,I140714,);
DFFARX1 I_8108 (I140847,I140830,I2966,I140714,);
not I_8109 (I140685,I140847);
DFFARX1 I_8110 (I140878,I140830,I2966,I140714,);
and I_8111 (I140679,I140765,I140878);
nand I_8112 (I140909,I128102,I128108);
and I_8113 (I140926,I140909,I128120);
DFFARX1 I_8114 (I140943,I140926,I2966,I140714,);
nor I_8115 (I140960,I140943,I140782);
not I_8116 (I140977,I140943);
nand I_8117 (I140688,I140765,I140977);
DFFARX1 I_8118 (I141008,I128126,I2966,I140714,);
and I_8119 (I141025,I141008,I128117);
nor I_8120 (I141042,I141025,I140943);
nor I_8121 (I141059,I141025,I140977);
nand I_8122 (I140694,I140813,I141059);
not I_8123 (I140697,I141025);
DFFARX1 I_8124 (I140676,I141025,I2966,I140714,);
DFFARX1 I_8125 (I141118,I128099,I2966,I140714,);
nand I_8126 (I141135,I141118,I140830);
and I_8127 (I141152,I140813,I141135);
DFFARX1 I_8128 (I140706,I141152,I2966,I140714,);
nor I_8129 (I140703,I141118,I141025);
and I_8130 (I141197,I141118,I140960);
or I_8131 (I141214,I140813,I141197);
DFFARX1 I_8132 (I140691,I141214,I2966,I140714,);
nand I_8133 (I140700,I141118,I141042);
not I_8134 (I141292,I2973);
nand I_8135 (I141309,I123941,I123929);
and I_8136 (I141326,I141309,I123923);
DFFARX1 I_8137 (I141343,I141326,I2966,I141292,);
not I_8138 (I141360,I141343);
DFFARX1 I_8139 (I141260,I141343,I2966,I141292,);
nor I_8140 (I141391,I123920,I123929);
DFFARX1 I_8141 (I141408,I123914,I2966,I141292,);
DFFARX1 I_8142 (I141425,I141408,I2966,I141292,);
not I_8143 (I141263,I141425);
DFFARX1 I_8144 (I141456,I141408,I2966,I141292,);
and I_8145 (I141257,I141343,I141456);
nand I_8146 (I141487,I123917,I123932);
and I_8147 (I141504,I141487,I123944);
DFFARX1 I_8148 (I141521,I141504,I2966,I141292,);
nor I_8149 (I141538,I141521,I141360);
not I_8150 (I141555,I141521);
nand I_8151 (I141266,I141343,I141555);
DFFARX1 I_8152 (I141586,I123935,I2966,I141292,);
and I_8153 (I141603,I141586,I123926);
nor I_8154 (I141620,I141603,I141521);
nor I_8155 (I141637,I141603,I141555);
nand I_8156 (I141272,I141391,I141637);
not I_8157 (I141275,I141603);
DFFARX1 I_8158 (I141254,I141603,I2966,I141292,);
DFFARX1 I_8159 (I141696,I123938,I2966,I141292,);
nand I_8160 (I141713,I141696,I141408);
and I_8161 (I141730,I141391,I141713);
DFFARX1 I_8162 (I141284,I141730,I2966,I141292,);
nor I_8163 (I141281,I141696,I141603);
and I_8164 (I141775,I141696,I141538);
or I_8165 (I141792,I141391,I141775);
DFFARX1 I_8166 (I141269,I141792,I2966,I141292,);
nand I_8167 (I141278,I141696,I141620);
not I_8168 (I141870,I2973);
nand I_8169 (I141887,I133585,I133582);
and I_8170 (I141904,I141887,I133579);
DFFARX1 I_8171 (I141921,I141904,I2966,I141870,);
nor I_8172 (I141938,I133570,I133582);
nor I_8173 (I141955,I141938,I141921);
not I_8174 (I141853,I141938);
DFFARX1 I_8175 (I141986,I133588,I2966,I141870,);
not I_8176 (I142003,I141986);
nor I_8177 (I142020,I141938,I142003);
nand I_8178 (I141856,I141986,I141955);
DFFARX1 I_8179 (I141838,I141986,I2966,I141870,);
nand I_8180 (I142065,I133573,I133597);
and I_8181 (I142082,I142065,I133576);
DFFARX1 I_8182 (I142099,I142082,I2966,I141870,);
nor I_8183 (I141859,I142099,I141921);
nand I_8184 (I141850,I142099,I142020);
DFFARX1 I_8185 (I142144,I133594,I2966,I141870,);
and I_8186 (I142161,I142144,I133591);
DFFARX1 I_8187 (I142178,I142161,I2966,I141870,);
not I_8188 (I141841,I142178);
nand I_8189 (I142209,I142161,I142099);
and I_8190 (I142226,I141921,I142209);
DFFARX1 I_8191 (I141832,I142226,I2966,I141870,);
DFFARX1 I_8192 (I142257,I133600,I2966,I141870,);
nand I_8193 (I142274,I142257,I141921);
and I_8194 (I142291,I142099,I142274);
DFFARX1 I_8195 (I141862,I142291,I2966,I141870,);
not I_8196 (I142322,I142257);
nor I_8197 (I142339,I141938,I142322);
and I_8198 (I142356,I142257,I142339);
or I_8199 (I142373,I142161,I142356);
DFFARX1 I_8200 (I141847,I142373,I2966,I141870,);
nand I_8201 (I141844,I142257,I142003);
DFFARX1 I_8202 (I141835,I142257,I2966,I141870,);
not I_8203 (I142465,I2973);
nand I_8204 (I142482,I140048,I140060);
and I_8205 (I142499,I142482,I140051);
DFFARX1 I_8206 (I142516,I142499,I2966,I142465,);
nor I_8207 (I142533,I140045,I140060);
DFFARX1 I_8208 (I142550,I140036,I2966,I142465,);
nand I_8209 (I142567,I142550,I142533);
DFFARX1 I_8210 (I142436,I142550,I2966,I142465,);
nand I_8211 (I142598,I140042,I140033);
and I_8212 (I142615,I142598,I140039);
DFFARX1 I_8213 (I142632,I142615,I2966,I142465,);
not I_8214 (I142649,I142632);
nor I_8215 (I142666,I142516,I142649);
and I_8216 (I142683,I142533,I142666);
and I_8217 (I142700,I142632,I142567);
DFFARX1 I_8218 (I142433,I142700,I2966,I142465,);
DFFARX1 I_8219 (I142427,I142632,I2966,I142465,);
DFFARX1 I_8220 (I142745,I140054,I2966,I142465,);
and I_8221 (I142762,I142745,I140030);
nand I_8222 (I142779,I142762,I142632);
nor I_8223 (I142454,I142762,I142533);
not I_8224 (I142810,I142762);
nor I_8225 (I142827,I142516,I142810);
nand I_8226 (I142445,I142550,I142827);
nand I_8227 (I142439,I142632,I142810);
or I_8228 (I142872,I142762,I142683);
DFFARX1 I_8229 (I142442,I142872,I2966,I142465,);
DFFARX1 I_8230 (I142903,I140057,I2966,I142465,);
and I_8231 (I142920,I142903,I142779);
DFFARX1 I_8232 (I142457,I142920,I2966,I142465,);
nor I_8233 (I142951,I142903,I142516);
nand I_8234 (I142451,I142762,I142951);
not I_8235 (I142448,I142903);
DFFARX1 I_8236 (I142996,I142903,I2966,I142465,);
and I_8237 (I142430,I142903,I142996);
not I_8238 (I143060,I2973);
nand I_8239 (I143077,I138756,I138759);
and I_8240 (I143094,I143077,I138738);
DFFARX1 I_8241 (I143111,I143094,I2966,I143060,);
not I_8242 (I143049,I143111);
DFFARX1 I_8243 (I143142,I143111,I2966,I143060,);
not I_8244 (I143037,I143142);
nor I_8245 (I143173,I138753,I138759);
not I_8246 (I143190,I143173);
nor I_8247 (I143207,I143111,I143190);
DFFARX1 I_8248 (I143224,I138762,I2966,I143060,);
not I_8249 (I143241,I143224);
nand I_8250 (I143040,I143224,I143190);
DFFARX1 I_8251 (I143272,I143224,I2966,I143060,);
and I_8252 (I143025,I143111,I143272);
nand I_8253 (I143303,I138750,I138768);
and I_8254 (I143320,I143303,I138744);
DFFARX1 I_8255 (I143337,I143320,I2966,I143060,);
nor I_8256 (I143354,I143337,I143241);
and I_8257 (I143371,I143173,I143354);
nor I_8258 (I143388,I143337,I143111);
DFFARX1 I_8259 (I143031,I143337,I2966,I143060,);
DFFARX1 I_8260 (I143419,I138741,I2966,I143060,);
and I_8261 (I143436,I143419,I138747);
or I_8262 (I143453,I143436,I143371);
DFFARX1 I_8263 (I143043,I143453,I2966,I143060,);
nand I_8264 (I143052,I143436,I143388);
DFFARX1 I_8265 (I143022,I143436,I2966,I143060,);
DFFARX1 I_8266 (I143512,I138765,I2966,I143060,);
nand I_8267 (I143046,I143512,I143207);
DFFARX1 I_8268 (I143034,I143512,I2966,I143060,);
nand I_8269 (I143557,I143512,I143173);
and I_8270 (I143574,I143224,I143557);
DFFARX1 I_8271 (I143028,I143574,I2966,I143060,);
not I_8272 (I143638,I2973);
nand I_8273 (I143655,I136773,I136764);
and I_8274 (I143672,I143655,I136779);
DFFARX1 I_8275 (I143689,I143672,I2966,I143638,);
not I_8276 (I143706,I143689);
nor I_8277 (I143723,I136749,I136764);
or I_8278 (I143621,I143723,I143689);
not I_8279 (I143609,I143723);
DFFARX1 I_8280 (I143768,I136752,I2966,I143638,);
nor I_8281 (I143785,I143768,I143723);
nand I_8282 (I143802,I136770,I136767);
and I_8283 (I143819,I143802,I136755);
DFFARX1 I_8284 (I143836,I143819,I2966,I143638,);
nor I_8285 (I143618,I143836,I143689);
not I_8286 (I143867,I143836);
nor I_8287 (I143884,I143768,I143867);
DFFARX1 I_8288 (I143901,I136776,I2966,I143638,);
and I_8289 (I143918,I143901,I136761);
or I_8290 (I143627,I143918,I143723);
nand I_8291 (I143606,I143918,I143884);
DFFARX1 I_8292 (I143963,I136758,I2966,I143638,);
and I_8293 (I143980,I143963,I143706);
nor I_8294 (I143624,I143918,I143980);
nor I_8295 (I144011,I143963,I143768);
DFFARX1 I_8296 (I143615,I144011,I2966,I143638,);
nor I_8297 (I143630,I143963,I143689);
not I_8298 (I144056,I143963);
nor I_8299 (I144073,I143836,I144056);
and I_8300 (I144090,I143723,I144073);
or I_8301 (I144107,I143918,I144090);
DFFARX1 I_8302 (I143603,I144107,I2966,I143638,);
nand I_8303 (I143612,I143963,I143785);
nand I_8304 (I143600,I143963,I143867);
not I_8305 (I144199,I2973);
nand I_8306 (I144216,I137436,I137427);
and I_8307 (I144233,I144216,I137442);
DFFARX1 I_8308 (I144250,I144233,I2966,I144199,);
not I_8309 (I144267,I144250);
nor I_8310 (I144284,I137412,I137427);
or I_8311 (I144182,I144284,I144250);
not I_8312 (I144170,I144284);
DFFARX1 I_8313 (I144329,I137415,I2966,I144199,);
nor I_8314 (I144346,I144329,I144284);
nand I_8315 (I144363,I137433,I137430);
and I_8316 (I144380,I144363,I137418);
DFFARX1 I_8317 (I144397,I144380,I2966,I144199,);
nor I_8318 (I144179,I144397,I144250);
not I_8319 (I144428,I144397);
nor I_8320 (I144445,I144329,I144428);
DFFARX1 I_8321 (I144462,I137439,I2966,I144199,);
and I_8322 (I144479,I144462,I137424);
or I_8323 (I144188,I144479,I144284);
nand I_8324 (I144167,I144479,I144445);
DFFARX1 I_8325 (I144524,I137421,I2966,I144199,);
and I_8326 (I144541,I144524,I144267);
nor I_8327 (I144185,I144479,I144541);
nor I_8328 (I144572,I144524,I144329);
DFFARX1 I_8329 (I144176,I144572,I2966,I144199,);
nor I_8330 (I144191,I144524,I144250);
not I_8331 (I144617,I144524);
nor I_8332 (I144634,I144397,I144617);
and I_8333 (I144651,I144284,I144634);
or I_8334 (I144668,I144479,I144651);
DFFARX1 I_8335 (I144164,I144668,I2966,I144199,);
nand I_8336 (I144173,I144524,I144346);
nand I_8337 (I144161,I144524,I144428);
not I_8338 (I144760,I2973);
nand I_8339 (I144777,I136110,I136101);
and I_8340 (I144794,I144777,I136116);
DFFARX1 I_8341 (I144811,I144794,I2966,I144760,);
not I_8342 (I144828,I144811);
nor I_8343 (I144845,I136086,I136101);
or I_8344 (I144743,I144845,I144811);
not I_8345 (I144731,I144845);
DFFARX1 I_8346 (I144890,I136089,I2966,I144760,);
nor I_8347 (I144907,I144890,I144845);
nand I_8348 (I144924,I136107,I136104);
and I_8349 (I144941,I144924,I136092);
DFFARX1 I_8350 (I144958,I144941,I2966,I144760,);
nor I_8351 (I144740,I144958,I144811);
not I_8352 (I144989,I144958);
nor I_8353 (I145006,I144890,I144989);
DFFARX1 I_8354 (I145023,I136113,I2966,I144760,);
and I_8355 (I145040,I145023,I136098);
or I_8356 (I144749,I145040,I144845);
nand I_8357 (I144728,I145040,I145006);
DFFARX1 I_8358 (I145085,I136095,I2966,I144760,);
and I_8359 (I145102,I145085,I144828);
nor I_8360 (I144746,I145040,I145102);
nor I_8361 (I145133,I145085,I144890);
DFFARX1 I_8362 (I144737,I145133,I2966,I144760,);
nor I_8363 (I144752,I145085,I144811);
not I_8364 (I145178,I145085);
nor I_8365 (I145195,I144958,I145178);
and I_8366 (I145212,I144845,I145195);
or I_8367 (I145229,I145040,I145212);
DFFARX1 I_8368 (I144725,I145229,I2966,I144760,);
nand I_8369 (I144734,I145085,I144907);
nand I_8370 (I144722,I145085,I144989);
not I_8371 (I145321,I2973);
not I_8372 (I145338,I138093);
nor I_8373 (I145355,I138090,I138078);
nand I_8374 (I145372,I145355,I138081);
DFFARX1 I_8375 (I145295,I145372,I2966,I145321,);
nor I_8376 (I145403,I145338,I138090);
nand I_8377 (I145420,I145403,I138087);
not I_8378 (I145310,I145420);
DFFARX1 I_8379 (I145292,I145420,I2966,I145321,);
not I_8380 (I145465,I138090);
not I_8381 (I145482,I145465);
not I_8382 (I145499,I138099);
nor I_8383 (I145516,I145499,I138075);
and I_8384 (I145533,I145516,I138096);
or I_8385 (I145550,I145533,I138084);
DFFARX1 I_8386 (I145567,I145550,I2966,I145321,);
nor I_8387 (I145584,I145567,I145420);
nor I_8388 (I145601,I145567,I145482);
nand I_8389 (I145307,I145372,I145601);
nand I_8390 (I145632,I145338,I138099);
nand I_8391 (I145649,I145632,I145567);
and I_8392 (I145666,I145632,I145649);
DFFARX1 I_8393 (I145289,I145666,I2966,I145321,);
DFFARX1 I_8394 (I145697,I145632,I2966,I145321,);
and I_8395 (I145286,I145465,I145697);
DFFARX1 I_8396 (I145728,I138105,I2966,I145321,);
not I_8397 (I145745,I145728);
nor I_8398 (I145762,I145420,I145745);
and I_8399 (I145779,I145728,I145762);
nand I_8400 (I145301,I145728,I145482);
DFFARX1 I_8401 (I145810,I145728,I2966,I145321,);
not I_8402 (I145298,I145810);
DFFARX1 I_8403 (I145841,I138102,I2966,I145321,);
not I_8404 (I145858,I145841);
or I_8405 (I145875,I145858,I145779);
DFFARX1 I_8406 (I145304,I145875,I2966,I145321,);
nand I_8407 (I145313,I145858,I145584);
DFFARX1 I_8408 (I145283,I145858,I2966,I145321,);
not I_8409 (I145967,I2973);
not I_8410 (I145984,I139402);
nor I_8411 (I146001,I139414,I139396);
nand I_8412 (I146018,I146001,I139411);
DFFARX1 I_8413 (I145941,I146018,I2966,I145967,);
nor I_8414 (I146049,I145984,I139414);
nand I_8415 (I146066,I146049,I139399);
not I_8416 (I145956,I146066);
DFFARX1 I_8417 (I145938,I146066,I2966,I145967,);
not I_8418 (I146111,I139414);
not I_8419 (I146128,I146111);
not I_8420 (I146145,I139408);
nor I_8421 (I146162,I146145,I139387);
and I_8422 (I146179,I146162,I139390);
or I_8423 (I146196,I146179,I139393);
DFFARX1 I_8424 (I146213,I146196,I2966,I145967,);
nor I_8425 (I146230,I146213,I146066);
nor I_8426 (I146247,I146213,I146128);
nand I_8427 (I145953,I146018,I146247);
nand I_8428 (I146278,I145984,I139408);
nand I_8429 (I146295,I146278,I146213);
and I_8430 (I146312,I146278,I146295);
DFFARX1 I_8431 (I145935,I146312,I2966,I145967,);
DFFARX1 I_8432 (I146343,I146278,I2966,I145967,);
and I_8433 (I145932,I146111,I146343);
DFFARX1 I_8434 (I146374,I139384,I2966,I145967,);
not I_8435 (I146391,I146374);
nor I_8436 (I146408,I146066,I146391);
and I_8437 (I146425,I146374,I146408);
nand I_8438 (I145947,I146374,I146128);
DFFARX1 I_8439 (I146456,I146374,I2966,I145967,);
not I_8440 (I145944,I146456);
DFFARX1 I_8441 (I146487,I139405,I2966,I145967,);
not I_8442 (I146504,I146487);
or I_8443 (I146521,I146504,I146425);
DFFARX1 I_8444 (I145950,I146521,I2966,I145967,);
nand I_8445 (I145959,I146504,I146230);
DFFARX1 I_8446 (I145929,I146504,I2966,I145967,);
not I_8447 (I146613,I2973);
or I_8448 (I146630,I143022,I143040);
or I_8449 (I146647,I143025,I143022);
DFFARX1 I_8450 (I146587,I146647,I2966,I146613,);
nor I_8451 (I146678,I143034,I143037);
not I_8452 (I146695,I146678);
not I_8453 (I146712,I143034);
and I_8454 (I146729,I146712,I143043);
nor I_8455 (I146746,I146729,I143040);
nor I_8456 (I146763,I143049,I143028);
DFFARX1 I_8457 (I146780,I146763,I2966,I146613,);
nand I_8458 (I146797,I146780,I146630);
and I_8459 (I146814,I146746,I146797);
DFFARX1 I_8460 (I146581,I146814,I2966,I146613,);
nor I_8461 (I146845,I143049,I143025);
DFFARX1 I_8462 (I146862,I146845,I2966,I146613,);
and I_8463 (I146578,I146678,I146862);
DFFARX1 I_8464 (I146893,I143052,I2966,I146613,);
and I_8465 (I146910,I146893,I143046);
DFFARX1 I_8466 (I146927,I146910,I2966,I146613,);
not I_8467 (I146590,I146927);
DFFARX1 I_8468 (I146575,I146910,I2966,I146613,);
DFFARX1 I_8469 (I146972,I143031,I2966,I146613,);
not I_8470 (I146989,I146972);
nor I_8471 (I147006,I146647,I146989);
and I_8472 (I147023,I146910,I147006);
or I_8473 (I147040,I146630,I147023);
DFFARX1 I_8474 (I146596,I147040,I2966,I146613,);
nor I_8475 (I147071,I146972,I146780);
nand I_8476 (I146605,I146746,I147071);
nor I_8477 (I147102,I146972,I146695);
nand I_8478 (I146599,I146845,I147102);
not I_8479 (I146602,I146972);
nand I_8480 (I146593,I146972,I146695);
DFFARX1 I_8481 (I146584,I146972,I2966,I146613,);
not I_8482 (I147208,I2973);
not I_8483 (I147225,I140691);
nor I_8484 (I147242,I140703,I140685);
nand I_8485 (I147259,I147242,I140706);
nor I_8486 (I147276,I147225,I140703);
nand I_8487 (I147293,I147276,I140697);
not I_8488 (I147310,I147293);
not I_8489 (I147327,I140703);
nor I_8490 (I147197,I147293,I147327);
not I_8491 (I147358,I147327);
nand I_8492 (I147182,I147293,I147358);
not I_8493 (I147389,I140688);
nor I_8494 (I147406,I147389,I140682);
and I_8495 (I147423,I147406,I140694);
or I_8496 (I147440,I147423,I140679);
DFFARX1 I_8497 (I147457,I147440,I2966,I147208,);
nor I_8498 (I147474,I147457,I147310);
DFFARX1 I_8499 (I147491,I147457,I2966,I147208,);
not I_8500 (I147179,I147491);
nand I_8501 (I147522,I147225,I140688);
and I_8502 (I147539,I147522,I147474);
DFFARX1 I_8503 (I147176,I147522,I2966,I147208,);
DFFARX1 I_8504 (I147570,I140676,I2966,I147208,);
nor I_8505 (I147587,I147570,I147293);
nand I_8506 (I147194,I147457,I147587);
nor I_8507 (I147618,I147570,I147358);
not I_8508 (I147191,I147570);
nand I_8509 (I147649,I147570,I147259);
and I_8510 (I147666,I147327,I147649);
DFFARX1 I_8511 (I147170,I147666,I2966,I147208,);
DFFARX1 I_8512 (I147173,I147570,I2966,I147208,);
DFFARX1 I_8513 (I147711,I140700,I2966,I147208,);
not I_8514 (I147728,I147711);
nand I_8515 (I147745,I147728,I147293);
and I_8516 (I147762,I147522,I147745);
DFFARX1 I_8517 (I147200,I147762,I2966,I147208,);
or I_8518 (I147793,I147728,I147539);
DFFARX1 I_8519 (I147185,I147793,I2966,I147208,);
nand I_8520 (I147188,I147728,I147618);
not I_8521 (I147871,I2973);
not I_8522 (I147888,I141269);
nor I_8523 (I147905,I141272,I141254);
nand I_8524 (I147922,I147905,I141281);
nor I_8525 (I147939,I147888,I141272);
nand I_8526 (I147956,I147939,I141260);
DFFARX1 I_8527 (I147973,I147956,I2966,I147871,);
not I_8528 (I147842,I147973);
not I_8529 (I148004,I141272);
not I_8530 (I148021,I148004);
not I_8531 (I148038,I141266);
nor I_8532 (I148055,I148038,I141278);
and I_8533 (I148072,I148055,I141284);
or I_8534 (I148089,I148072,I141263);
DFFARX1 I_8535 (I148106,I148089,I2966,I147871,);
DFFARX1 I_8536 (I147839,I148106,I2966,I147871,);
DFFARX1 I_8537 (I148137,I148106,I2966,I147871,);
DFFARX1 I_8538 (I147833,I148106,I2966,I147871,);
nand I_8539 (I148168,I147888,I141266);
nand I_8540 (I148185,I148168,I147922);
and I_8541 (I148202,I148004,I148185);
DFFARX1 I_8542 (I147863,I148202,I2966,I147871,);
and I_8543 (I147836,I148168,I148137);
DFFARX1 I_8544 (I148247,I141275,I2966,I147871,);
nor I_8545 (I147860,I148247,I148168);
nor I_8546 (I148278,I148247,I147922);
nand I_8547 (I147857,I147956,I148278);
not I_8548 (I147854,I148247);
DFFARX1 I_8549 (I148323,I141257,I2966,I147871,);
not I_8550 (I148340,I148323);
nor I_8551 (I148357,I148340,I148021);
and I_8552 (I148374,I148247,I148357);
or I_8553 (I148391,I148168,I148374);
DFFARX1 I_8554 (I147848,I148391,I2966,I147871,);
not I_8555 (I148422,I148340);
nor I_8556 (I148439,I148247,I148422);
nand I_8557 (I147851,I148340,I148439);
nand I_8558 (I147845,I148004,I148422);
not I_8559 (I148517,I2973);
nand I_8560 (I148534,I144176,I144191);
and I_8561 (I148551,I148534,I144179);
DFFARX1 I_8562 (I148568,I148551,I2966,I148517,);
not I_8563 (I148585,I148568);
DFFARX1 I_8564 (I148485,I148568,I2966,I148517,);
nor I_8565 (I148616,I144188,I144191);
DFFARX1 I_8566 (I148633,I144173,I2966,I148517,);
DFFARX1 I_8567 (I148650,I148633,I2966,I148517,);
not I_8568 (I148488,I148650);
DFFARX1 I_8569 (I148681,I148633,I2966,I148517,);
and I_8570 (I148482,I148568,I148681);
nand I_8571 (I148712,I144164,I144161);
and I_8572 (I148729,I148712,I144167);
DFFARX1 I_8573 (I148746,I148729,I2966,I148517,);
nor I_8574 (I148763,I148746,I148585);
not I_8575 (I148780,I148746);
nand I_8576 (I148491,I148568,I148780);
DFFARX1 I_8577 (I148811,I144170,I2966,I148517,);
and I_8578 (I148828,I148811,I144182);
nor I_8579 (I148845,I148828,I148746);
nor I_8580 (I148862,I148828,I148780);
nand I_8581 (I148497,I148616,I148862);
not I_8582 (I148500,I148828);
DFFARX1 I_8583 (I148479,I148828,I2966,I148517,);
DFFARX1 I_8584 (I148921,I144185,I2966,I148517,);
nand I_8585 (I148938,I148921,I148633);
and I_8586 (I148955,I148616,I148938);
DFFARX1 I_8587 (I148509,I148955,I2966,I148517,);
nor I_8588 (I148506,I148921,I148828);
and I_8589 (I149000,I148921,I148763);
or I_8590 (I149017,I148616,I149000);
DFFARX1 I_8591 (I148494,I149017,I2966,I148517,);
nand I_8592 (I148503,I148921,I148845);
not I_8593 (I149095,I2973);
not I_8594 (I149112,I147188);
nor I_8595 (I149129,I147194,I147173);
nand I_8596 (I149146,I149129,I147179);
nor I_8597 (I149163,I149112,I147194);
nand I_8598 (I149180,I149163,I147185);
not I_8599 (I149197,I147194);
not I_8600 (I149214,I149197);
not I_8601 (I149231,I147182);
nor I_8602 (I149248,I149231,I147200);
and I_8603 (I149265,I149248,I147191);
or I_8604 (I149282,I149265,I147170);
DFFARX1 I_8605 (I149299,I149282,I2966,I149095,);
nand I_8606 (I149316,I149112,I147182);
or I_8607 (I149084,I149316,I149299);
not I_8608 (I149347,I149316);
nor I_8609 (I149364,I149299,I149347);
and I_8610 (I149381,I149197,I149364);
nand I_8611 (I149057,I149316,I149214);
DFFARX1 I_8612 (I149412,I147197,I2966,I149095,);
or I_8613 (I149078,I149412,I149299);
nor I_8614 (I149443,I149412,I149180);
nor I_8615 (I149460,I149412,I149214);
nand I_8616 (I149063,I149146,I149460);
or I_8617 (I149491,I149412,I149381);
DFFARX1 I_8618 (I149060,I149491,I2966,I149095,);
not I_8619 (I149066,I149412);
DFFARX1 I_8620 (I149536,I147176,I2966,I149095,);
not I_8621 (I149553,I149536);
nor I_8622 (I149570,I149553,I149146);
DFFARX1 I_8623 (I149072,I149570,I2966,I149095,);
nor I_8624 (I149087,I149412,I149553);
nor I_8625 (I149075,I149553,I149316);
not I_8626 (I149629,I149553);
and I_8627 (I149646,I149180,I149629);
nor I_8628 (I149081,I149316,I149646);
nand I_8629 (I149069,I149553,I149443);
not I_8630 (I149724,I2973);
nand I_8631 (I149741,I144746,I144731);
and I_8632 (I149758,I149741,I144740);
DFFARX1 I_8633 (I149775,I149758,I2966,I149724,);
not I_8634 (I149713,I149775);
DFFARX1 I_8635 (I149806,I149775,I2966,I149724,);
not I_8636 (I149701,I149806);
nor I_8637 (I149837,I144752,I144731);
not I_8638 (I149854,I149837);
nor I_8639 (I149871,I149775,I149854);
DFFARX1 I_8640 (I149888,I144743,I2966,I149724,);
not I_8641 (I149905,I149888);
nand I_8642 (I149704,I149888,I149854);
DFFARX1 I_8643 (I149936,I149888,I2966,I149724,);
and I_8644 (I149689,I149775,I149936);
nand I_8645 (I149967,I144728,I144722);
and I_8646 (I149984,I149967,I144737);
DFFARX1 I_8647 (I150001,I149984,I2966,I149724,);
nor I_8648 (I150018,I150001,I149905);
and I_8649 (I150035,I149837,I150018);
nor I_8650 (I150052,I150001,I149775);
DFFARX1 I_8651 (I149695,I150001,I2966,I149724,);
DFFARX1 I_8652 (I150083,I144725,I2966,I149724,);
and I_8653 (I150100,I150083,I144749);
or I_8654 (I150117,I150100,I150035);
DFFARX1 I_8655 (I149707,I150117,I2966,I149724,);
nand I_8656 (I149716,I150100,I150052);
DFFARX1 I_8657 (I149686,I150100,I2966,I149724,);
DFFARX1 I_8658 (I150176,I144734,I2966,I149724,);
nand I_8659 (I149710,I150176,I149871);
DFFARX1 I_8660 (I149698,I150176,I2966,I149724,);
nand I_8661 (I150221,I150176,I149837);
and I_8662 (I150238,I149888,I150221);
DFFARX1 I_8663 (I149692,I150238,I2966,I149724,);
not I_8664 (I150302,I2973);
nand I_8665 (I150319,I147863,I147854);
and I_8666 (I150336,I150319,I147857);
DFFARX1 I_8667 (I150353,I150336,I2966,I150302,);
not I_8668 (I150370,I150353);
nor I_8669 (I150387,I147833,I147854);
or I_8670 (I150285,I150387,I150353);
not I_8671 (I150273,I150387);
DFFARX1 I_8672 (I150432,I147848,I2966,I150302,);
nor I_8673 (I150449,I150432,I150387);
nand I_8674 (I150466,I147836,I147851);
and I_8675 (I150483,I150466,I147845);
DFFARX1 I_8676 (I150500,I150483,I2966,I150302,);
nor I_8677 (I150282,I150500,I150353);
not I_8678 (I150531,I150500);
nor I_8679 (I150548,I150432,I150531);
DFFARX1 I_8680 (I150565,I147860,I2966,I150302,);
and I_8681 (I150582,I150565,I147839);
or I_8682 (I150291,I150582,I150387);
nand I_8683 (I150270,I150582,I150548);
DFFARX1 I_8684 (I150627,I147842,I2966,I150302,);
and I_8685 (I150644,I150627,I150370);
nor I_8686 (I150288,I150582,I150644);
nor I_8687 (I150675,I150627,I150432);
DFFARX1 I_8688 (I150279,I150675,I2966,I150302,);
nor I_8689 (I150294,I150627,I150353);
not I_8690 (I150720,I150627);
nor I_8691 (I150737,I150500,I150720);
and I_8692 (I150754,I150387,I150737);
or I_8693 (I150771,I150582,I150754);
DFFARX1 I_8694 (I150267,I150771,I2966,I150302,);
nand I_8695 (I150276,I150627,I150449);
nand I_8696 (I150264,I150627,I150531);
not I_8697 (I150863,I2973);
not I_8698 (I150880,I148494);
nor I_8699 (I150897,I148506,I148488);
nand I_8700 (I150914,I150897,I148509);
nor I_8701 (I150931,I150880,I148506);
nand I_8702 (I150948,I150931,I148500);
not I_8703 (I150965,I150948);
not I_8704 (I150982,I148506);
nor I_8705 (I150852,I150948,I150982);
not I_8706 (I151013,I150982);
nand I_8707 (I150837,I150948,I151013);
not I_8708 (I151044,I148491);
nor I_8709 (I151061,I151044,I148485);
and I_8710 (I151078,I151061,I148497);
or I_8711 (I151095,I151078,I148482);
DFFARX1 I_8712 (I151112,I151095,I2966,I150863,);
nor I_8713 (I151129,I151112,I150965);
DFFARX1 I_8714 (I151146,I151112,I2966,I150863,);
not I_8715 (I150834,I151146);
nand I_8716 (I151177,I150880,I148491);
and I_8717 (I151194,I151177,I151129);
DFFARX1 I_8718 (I150831,I151177,I2966,I150863,);
DFFARX1 I_8719 (I151225,I148479,I2966,I150863,);
nor I_8720 (I151242,I151225,I150948);
nand I_8721 (I150849,I151112,I151242);
nor I_8722 (I151273,I151225,I151013);
not I_8723 (I150846,I151225);
nand I_8724 (I151304,I151225,I150914);
and I_8725 (I151321,I150982,I151304);
DFFARX1 I_8726 (I150825,I151321,I2966,I150863,);
DFFARX1 I_8727 (I150828,I151225,I2966,I150863,);
DFFARX1 I_8728 (I151366,I148503,I2966,I150863,);
not I_8729 (I151383,I151366);
nand I_8730 (I151400,I151383,I150948);
and I_8731 (I151417,I151177,I151400);
DFFARX1 I_8732 (I150855,I151417,I2966,I150863,);
or I_8733 (I151448,I151383,I151194);
DFFARX1 I_8734 (I150840,I151448,I2966,I150863,);
nand I_8735 (I150843,I151383,I151273);
endmodule


