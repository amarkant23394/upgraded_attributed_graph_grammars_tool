module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_7_r_5,n7_5,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_5,n28_5,n46_5);
nand I_37(N1508_0_r_5,n26_5,n43_5);
not I_38(N1372_1_r_5,n43_5);
nor I_39(N1508_1_r_5,n30_5,n43_5);
nor I_40(N6147_2_r_5,n29_5,n32_5);
nor I_41(N1507_6_r_5,n26_5,n44_5);
nor I_42(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_43(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_44(n_572_7_r_5,n27_5,n28_5);
nand I_45(n_573_7_r_5,n26_5,n27_5);
nand I_46(n_549_7_r_5,N1372_1_r_3,N1508_1_r_3);
nand I_47(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_48(n_452_7_r_5,n29_5);
nor I_49(n4_7_r_5,n30_5,n31_5);
not I_50(n7_5,blif_reset_net_7_r_5);
not I_51(n26_5,n35_5);
nand I_52(n27_5,n40_5,n41_5);
nand I_53(n28_5,N1508_6_r_3,n_549_7_r_3);
nand I_54(n29_5,n27_5,n33_5);
nor I_55(n30_5,n45_5,N1372_1_r_3);
not I_56(n31_5,n_549_7_r_5);
nor I_57(n32_5,n34_5,n35_5);
not I_58(n33_5,n30_5);
nor I_59(n34_5,n31_5,n36_5);
nor I_60(n35_5,n28_5,n_569_7_r_3);
not I_61(n36_5,n28_5);
nand I_62(n37_5,n36_5,n38_5);
nand I_63(n38_5,n26_5,n39_5);
nand I_64(n39_5,n30_5,n31_5);
nor I_65(n40_5,N1507_6_r_3,G42_7_r_3);
or I_66(n41_5,n42_5,G42_7_r_3);
nor I_67(n42_5,n_573_7_r_3,N1508_6_r_3);
nand I_68(n43_5,n36_5,n46_5);
nor I_69(n44_5,n_549_7_r_5,n33_5);
or I_70(n45_5,N1508_1_r_3,n_452_7_r_3);
and I_71(n46_5,n31_5,n47_5);
or I_72(n47_5,N6134_9_r_3,N1507_6_r_3);
endmodule


