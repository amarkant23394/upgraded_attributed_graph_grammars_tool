module test_final(IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_102_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13,n4_7_l_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_13,n59_13,n61_13);
nor I_1(N1508_0_r_13,n59_13,n60_13);
not I_2(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_3(n_431_5_r_13,blif_clk_net_7_r_1,n9_1,G78_5_r_13,);
nand I_4(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_5(n_102_5_r_13,IN_9_7_l_13,IN_10_7_l_13);
nand I_6(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_7(n1_13,blif_clk_net_7_r_1,n9_1,G42_7_r_13,);
nor I_8(n_572_7_r_13,n40_13,n41_13);
nand I_9(n_573_7_r_13,n37_13,n38_13);
nor I_10(n_549_7_r_13,n46_13,n47_13);
nand I_11(n_569_7_r_13,n37_13,n43_13);
nand I_12(n_452_7_r_13,n52_13,n53_13);
nor I_13(n4_7_l_13,G18_7_l_13,IN_1_7_l_13);
DFFARX1 I_14(n4_7_l_13,blif_clk_net_7_r_1,n9_1,n62_13,);
not I_15(n33_13,n62_13);
nand I_16(n_431_5_r_13,n54_13,n55_13);
not I_17(n1_13,n52_13);
nor I_18(n34_13,n35_13,n36_13);
nor I_19(n35_13,G15_7_l_13,n42_13);
nand I_20(n36_13,n50_13,n58_13);
nand I_21(n37_13,n44_13,n45_13);
or I_22(n38_13,IN_3_1_l_13,n39_13);
nand I_23(n39_13,IN_1_1_l_13,IN_2_1_l_13);
not I_24(n40_13,n36_13);
nor I_25(n41_13,IN_10_7_l_13,n35_13);
not I_26(n42_13,IN_4_7_l_13);
or I_27(n43_13,G18_7_l_13,IN_5_7_l_13);
not I_28(n44_13,G15_7_l_13);
not I_29(n45_13,IN_7_7_l_13);
nor I_30(n46_13,n39_13,n40_13);
nor I_31(n47_13,G18_7_l_13,IN_5_7_l_13);
nor I_32(n48_13,n50_13,n51_13);
nor I_33(n49_13,G15_7_l_13,IN_7_7_l_13);
not I_34(n50_13,n59_13);
not I_35(n51_13,n_102_5_r_13);
nand I_36(n52_13,n33_13,n39_13);
nand I_37(n53_13,IN_3_1_l_13,n33_13);
nor I_38(n54_13,IN_5_7_l_13,IN_9_7_l_13);
nand I_39(n55_13,n62_13,n56_13);
nor I_40(n56_13,n39_13,n57_13);
not I_41(n57_13,G18_7_l_13);
or I_42(n58_13,IN_3_10_l_13,IN_4_10_l_13);
nand I_43(n59_13,IN_1_10_l_13,IN_2_10_l_13);
nor I_44(n60_13,IN_5_7_l_13,n51_13);
nor I_45(n61_13,IN_3_1_l_13,n39_13);
and I_46(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_47(N1508_0_r_1,n40_1,n44_1);
nor I_48(N1507_6_r_1,n43_1,n49_1);
nor I_49(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_50(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_51(n_572_7_r_1,n29_1,n30_1);
not I_52(n_573_7_r_1,n_452_7_r_1);
nor I_53(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_54(n_569_7_r_1,n30_1,n31_1);
nor I_55(n_452_7_r_1,n30_1,n32_1);
nor I_56(N6147_9_r_1,n35_1,n36_1);
nand I_57(N6134_9_r_1,n38_1,n39_1);
not I_58(I_BUFF_1_9_r_1,n40_1);
nor I_59(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_60(n9_1,blif_reset_net_7_r_1);
nor I_61(n29_1,n34_1,n_572_7_r_13);
nor I_62(n30_1,n33_1,n34_1);
nor I_63(n31_1,n54_1,N1508_0_r_13);
not I_64(n32_1,n48_1);
nor I_65(n33_1,n_429_or_0_5_r_13,G78_5_r_13);
not I_66(n34_1,N1371_0_r_13);
nor I_67(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_68(n36_1,n29_1);
not I_69(n37_1,n41_1);
nand I_70(n38_1,I_BUFF_1_9_r_1,N1508_0_r_13);
nand I_71(n39_1,n37_1,n40_1);
nand I_72(n40_1,n_547_5_r_13,n_569_7_r_13);
nand I_73(n41_1,n52_1,G42_7_r_13);
or I_74(n42_1,n36_1,n43_1);
nor I_75(n43_1,n32_1,n49_1);
nand I_76(n44_1,n45_1,n46_1);
nand I_77(n45_1,n47_1,n48_1);
not I_78(n46_1,N1508_0_r_13);
not I_79(n47_1,n31_1);
nand I_80(n48_1,n50_1,n_576_5_r_13);
nor I_81(n49_1,n41_1,n47_1);
and I_82(n50_1,n51_1,n_452_7_r_13);
nand I_83(n51_1,n52_1,n53_1);
nand I_84(n52_1,n_573_7_r_13,n_549_7_r_13);
not I_85(n53_1,G42_7_r_13);
or I_86(n54_1,N1371_0_r_13,n_429_or_0_5_r_13);
nor I_87(n55_1,n29_1,N1508_0_r_13);
endmodule


