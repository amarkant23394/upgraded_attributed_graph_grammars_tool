module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_5_r_11,n9_11,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
not I_41(N1372_1_r_11,n53_11);
nor I_42(N1508_1_r_11,n39_11,n53_11);
nor I_43(N6147_2_r_11,n48_11,n49_11);
nor I_44(N6147_3_r_11,n44_11,n45_11);
nand I_45(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_46(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_47(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_48(n_102_5_r_11,n39_11);
nand I_49(n_547_5_r_11,n36_11,n37_11);
nor I_50(N1507_6_r_11,n52_11,n57_11);
nor I_51(N1508_6_r_11,n46_11,n51_11);
nor I_52(N1372_10_r_11,n43_11,n47_11);
nor I_53(N1508_10_r_11,n55_11,n56_11);
nand I_54(n_431_5_r_11,n40_11,n41_11);
not I_55(n9_11,blif_reset_net_5_r_11);
nor I_56(n36_11,n38_11,n39_11);
not I_57(n37_11,n40_11);
nor I_58(n38_11,n60_11,N6134_9_r_1);
nor I_59(n39_11,n54_11,N1507_6_r_1);
nand I_60(n40_11,G42_7_r_1,n_572_7_r_1);
nand I_61(n41_11,n_102_5_r_11,n42_11);
and I_62(n42_11,n58_11,n_569_7_r_1);
not I_63(n43_11,n44_11);
nor I_64(n44_11,n40_11,N6147_9_r_1);
nand I_65(n45_11,n46_11,n47_11);
not I_66(n46_11,n38_11);
nand I_67(n47_11,n59_11,n62_11);
and I_68(n48_11,n37_11,n47_11);
or I_69(n49_11,n44_11,n50_11);
nor I_70(n50_11,n60_11,n61_11);
or I_71(n51_11,n_102_5_r_11,n52_11);
nor I_72(n52_11,n42_11,n57_11);
nand I_73(n53_11,n37_11,n50_11);
or I_74(n54_11,N1508_0_r_1,N1507_6_r_1);
nor I_75(n55_11,n38_11,n42_11);
not I_76(n56_11,N1372_10_r_11);
and I_77(n57_11,n38_11,n50_11);
and I_78(n58_11,n59_11,N1508_0_r_1);
or I_79(n59_11,n63_11,n_573_7_r_1);
not I_80(n60_11,n_549_7_r_1);
nor I_81(n61_11,n_572_7_r_1,n_573_7_r_1);
nand I_82(n62_11,N1508_6_r_1,G42_7_r_1);
and I_83(n63_11,N1508_6_r_1,G42_7_r_1);
endmodule


