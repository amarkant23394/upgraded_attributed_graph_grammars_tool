module test_I8267(I1477,I5785,I5864,I1470,I4691,I8267);
input I1477,I5785,I5864,I1470,I4691;
output I8267;
wire I5963,I4869,I5898,I5802,I5716,I4518,I5881,I5719,I8250,I5737,I6265,I6203,I5751,I5915,I6248;
DFFARX1 I_0(I5915,I1470,I5751,,,I5963,);
DFFARX1 I_1(I1470,,,I4869,);
nor I_2(I5898,I5802,I5881);
DFFARX1 I_3(I5785,I1470,I5751,,,I5802,);
and I_4(I5716,I5802,I5963);
nand I_5(I4518,I4869,I4691);
not I_6(I5881,I5864);
DFFARX1 I_7(I6265,I1470,I5751,,,I5719,);
nor I_8(I8250,I5719,I5716);
nand I_9(I5737,I6203,I5898);
and I_10(I6265,I5915,I6248);
DFFARX1 I_11(I4518,I1470,I5751,,,I6203,);
not I_12(I5751,I1477);
DFFARX1 I_13(I1470,I5751,,,I5915,);
nand I_14(I8267,I8250,I5737);
nand I_15(I6248,I6203,I5864);
endmodule


