module test_I8824(I7156,I6975,I7427,I7026,I5097,I8824);
input I7156,I6975,I7427,I7026,I5097;
output I8824;
wire I6893,I6992,I7317,I8981,I7057,I6881,I8879,I6887,I9083,I7286,I8964;
nand I_0(I8824,I9083,I8981);
nand I_1(I6893,I7156,I7286);
nand I_2(I6992,I6975,I5097);
nor I_3(I7317,I7057);
not I_4(I8981,I8964);
not I_5(I7057,I7026);
nand I_6(I6881,I6992,I7057);
not I_7(I8879,I6887);
nand I_8(I6887,I7427,I7317);
nand I_9(I9083,I8879,I6881);
nor I_10(I7286,I6992);
not I_11(I8964,I6893);
endmodule


