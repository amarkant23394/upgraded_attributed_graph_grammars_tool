module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_8_r_10,n11_10,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N1371_0_r_10,n37_10,n38_10);
nor I_42(N1508_0_r_10,n37_10,n58_10);
nand I_43(N6147_2_r_10,n39_10,n40_10);
not I_44(N6147_3_r_10,n39_10);
nor I_45(N1372_4_r_10,n46_10,n49_10);
nor I_46(N1508_4_r_10,n51_10,n52_10);
nor I_47(N1507_6_r_10,n49_10,n60_10);
nor I_48(N1508_6_r_10,n49_10,n50_10);
nor I_49(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_50(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_51(N6147_9_r_10,n36_10,n37_10);
nor I_52(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_53(I_BUFF_1_9_r_10,n48_10);
nor I_54(N3_8_r_10,n44_10,n47_10);
not I_55(n11_10,blif_reset_net_8_r_10);
not I_56(n35_10,n49_10);
nor I_57(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_58(n37_10,N6147_9_r_1);
not I_59(n38_10,n46_10);
nand I_60(n39_10,n43_10,n44_10);
nand I_61(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_62(n41_10,n42_10,N6147_9_r_1);
not I_63(n42_10,n44_10);
nor I_64(n43_10,n45_10,N6147_9_r_1);
nand I_65(n44_10,n54_10,N1507_6_r_1);
nor I_66(n45_10,n59_10,n_572_7_r_1);
nand I_67(n46_10,n61_10,N1508_0_r_1);
nor I_68(n47_10,n46_10,n48_10);
nand I_69(n48_10,n62_10,n63_10);
nand I_70(n49_10,n56_10,N1508_0_r_1);
not I_71(n50_10,n45_10);
nor I_72(n51_10,n42_10,n53_10);
not I_73(n52_10,N1372_4_r_10);
nor I_74(n53_10,n48_10,n50_10);
and I_75(n54_10,n55_10,n_572_7_r_1);
nand I_76(n55_10,n56_10,n57_10);
nand I_77(n56_10,n_573_7_r_1,N1508_6_r_1);
not I_78(n57_10,N1508_0_r_1);
nor I_79(n58_10,n35_10,n45_10);
nor I_80(n59_10,n_569_7_r_1,G42_7_r_1);
nor I_81(n60_10,n37_10,n46_10);
or I_82(n61_10,n_569_7_r_1,G42_7_r_1);
nor I_83(n62_10,N1508_6_r_1,G42_7_r_1);
or I_84(n63_10,n64_10,n_549_7_r_1);
nor I_85(n64_10,N1507_6_r_1,N6134_9_r_1);
endmodule


