module test_I8981(I7139,I6992,I1470,I6907,I8981);
input I7139,I6992,I1470,I6907;
output I8981;
wire I6893,I7156,I7269,I7286,I8964;
nand I_0(I6893,I7156,I7286);
DFFARX1 I_1(I7139,I1470,I6907,,,I7156,);
not I_2(I8981,I8964);
DFFARX1 I_3(I1470,I6907,,,I7269,);
nor I_4(I7286,I7269,I6992);
not I_5(I8964,I6893);
endmodule


