module test_I12024(I7556,I10349,I10270,I10154,I1477,I1470,I12024);
input I7556,I10349,I10270,I10154,I1477,I1470;
output I12024;
wire I10029,I10219,I12007,I10507,I10044,I10020,I10490,I10052,I10287,I10366,I10459;
DFFARX1 I_0(I10459,I1470,I10052,,,I10029,);
DFFARX1 I_1(I1470,I10052,,,I10219,);
nor I_2(I12007,I10020,I10029);
and I_3(I10507,I10490,I10366);
DFFARX1 I_4(I10507,I1470,I10052,,,I10044,);
DFFARX1 I_5(I10287,I1470,I10052,,,I10020,);
nand I_6(I12024,I12007,I10044);
DFFARX1 I_7(I7556,I1470,I10052,,,I10490,);
not I_8(I10052,I1477);
and I_9(I10287,I10219,I10154);
nand I_10(I10366,I10349,I10219);
or I_11(I10459,I10349,I10270);
endmodule


