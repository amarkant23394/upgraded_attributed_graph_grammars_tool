module test_I8377(I6248,I1477,I1470,I8377);
input I6248,I1477,I1470;
output I8377;
wire I6265,I8360,I5751,I5915,I5719;
and I_0(I6265,I5915,I6248);
not I_1(I8360,I5719);
not I_2(I5751,I1477);
DFFARX1 I_3(I1470,I5751,,,I5915,);
DFFARX1 I_4(I6265,I1470,I5751,,,I5719,);
not I_5(I8377,I8360);
endmodule


