module test_I3297(I1902,I2702,I1294,I1920,I2914,I1301,I3297);
input I1902,I2702,I1294,I1920,I2914,I1301;
output I3297;
wire I2563,I2733,I3103,I3168,I2548,I2560,I2583,I3280,I2993,I2945,I3086;
nand I_0(I2563,I3103,I2993);
not I_1(I2733,I2702);
not I_2(I3103,I3086);
or I_3(I3168,I3103,I2914);
DFFARX1 I_4(I2945,I1294,I2583,,,I2548,);
DFFARX1 I_5(I3168,I1294,I2583,,,I2560,);
not I_6(I2583,I1301);
nor I_7(I3280,I2548,I2560);
nor I_8(I2993,I2945,I2733);
DFFARX1 I_9(I1902,I1294,I2583,,,I2945,);
DFFARX1 I_10(I1920,I1294,I2583,,,I3086,);
nand I_11(I3297,I3280,I2563);
endmodule


