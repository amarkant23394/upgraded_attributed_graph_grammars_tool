module test_I2251(I1749,I1294,I1492,I1301,I1704,I2251);
input I1749,I1294,I1492,I1301,I1704;
output I2251;
wire I1797,I1322,I1656,I1971,I2234,I1334,I1310,I1577,I1319,I1427,I1954,I1780,I1342,I1988,I1509,I1304;
and I_0(I1797,I1780,I1656);
nand I_1(I1322,I1427,I1704);
nand I_2(I1656,I1509);
nor I_3(I1971,I1310,I1319);
nand I_4(I2234,I1954,I1304);
DFFARX1 I_5(I1797,I1294,I1342,,,I1334,);
DFFARX1 I_6(I1577,I1294,I1342,,,I1310,);
and I_7(I1577,I1509);
DFFARX1 I_8(I1749,I1294,I1342,,,I1319,);
DFFARX1 I_9(I1294,I1342,,,I1427,);
not I_10(I1954,I1322);
DFFARX1 I_11(I1294,I1342,,,I1780,);
nand I_12(I2251,I2234,I1988);
not I_13(I1342,I1301);
nand I_14(I1988,I1971,I1334);
DFFARX1 I_15(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_16(I1509,I1294,I1342,,,I1304,);
endmodule


