module test_I14338(I13177,I1477,I14503,I1470,I13186,I14338);
input I13177,I1477,I14503,I1470,I13186;
output I14338;
wire I14438,I14472,I14520,I14455,I13174,I14537,I13159,I14605,I14370;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
nor I_1(I14438,I13159,I13186);
nand I_2(I14472,I14455,I14438);
and I_3(I14520,I14503,I13174);
DFFARX1 I_4(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_5(I1470,,,I13174,);
DFFARX1 I_6(I14520,I1470,I14370,,,I14537,);
DFFARX1 I_7(I1470,,,I13159,);
and I_8(I14605,I14537,I14472);
not I_9(I14370,I1477);
endmodule


