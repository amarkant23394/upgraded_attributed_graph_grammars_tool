module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_7_r_1,n9_1,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
and I_39(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_40(N1508_0_r_1,n40_1,n44_1);
nor I_41(N1507_6_r_1,n43_1,n49_1);
nor I_42(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_43(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_44(n_572_7_r_1,n29_1,n30_1);
not I_45(n_573_7_r_1,n_452_7_r_1);
nor I_46(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_47(n_569_7_r_1,n30_1,n31_1);
nor I_48(n_452_7_r_1,n30_1,n32_1);
nor I_49(N6147_9_r_1,n35_1,n36_1);
nand I_50(N6134_9_r_1,n38_1,n39_1);
not I_51(I_BUFF_1_9_r_1,n40_1);
nor I_52(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_53(n9_1,blif_reset_net_7_r_1);
nor I_54(n29_1,n34_1,N1508_6_r_6);
nor I_55(n30_1,n33_1,n34_1);
nor I_56(n31_1,n54_1,n_42_8_r_6);
not I_57(n32_1,n48_1);
nor I_58(n33_1,N1371_0_r_6,N1372_1_r_6);
not I_59(n34_1,N1508_10_r_6);
nor I_60(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_61(n36_1,n29_1);
not I_62(n37_1,n41_1);
nand I_63(n38_1,I_BUFF_1_9_r_1,G199_8_r_6);
nand I_64(n39_1,n37_1,n40_1);
nand I_65(n40_1,N1372_1_r_6,N1508_0_r_6);
nand I_66(n41_1,n52_1,N1507_6_r_6);
or I_67(n42_1,n36_1,n43_1);
nor I_68(n43_1,n32_1,n49_1);
nand I_69(n44_1,n45_1,n46_1);
nand I_70(n45_1,n47_1,n48_1);
not I_71(n46_1,G199_8_r_6);
not I_72(n47_1,n31_1);
nand I_73(n48_1,n50_1,N6134_9_r_6);
nor I_74(n49_1,n41_1,n47_1);
and I_75(n50_1,n51_1,N1508_0_r_6);
nand I_76(n51_1,n52_1,n53_1);
nand I_77(n52_1,N6147_9_r_6,N1372_10_r_6);
not I_78(n53_1,N1507_6_r_6);
or I_79(n54_1,N1508_1_r_6,N1371_0_r_6);
nor I_80(n55_1,n29_1,G199_8_r_6);
endmodule


