module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n_102_5_r_0,n_452_7_r_0,n_431_5_r_0,n6_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_5_r_0,n6_0,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_5_r_0,n6_0,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_41(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_42(n_429_or_0_5_r_0,n38_0,N1372_1_r_16);
DFFARX1 I_43(n_431_5_r_0,blif_clk_net_5_r_0,n6_0,G78_5_r_0,);
nand I_44(n_576_5_r_0,n26_0,N1372_1_r_16);
not I_45(n_102_5_r_0,n27_0);
nand I_46(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_47(n4_7_r_0,blif_clk_net_5_r_0,n6_0,G42_7_r_0,);
nor I_48(n_572_7_r_0,n31_0,N1372_1_r_16);
or I_49(n_573_7_r_0,n29_0,n30_0);
nor I_50(n_549_7_r_0,n29_0,n33_0);
nand I_51(n_569_7_r_0,n28_0,n32_0);
nor I_52(n_452_7_r_0,n30_0,n31_0);
nand I_53(n_431_5_r_0,n_102_5_r_0,n35_0);
not I_54(n6_0,blif_reset_net_5_r_0);
nor I_55(n4_7_r_0,n31_0,n37_0);
nor I_56(n26_0,n27_0,n28_0);
nor I_57(n27_0,n28_0,n44_0);
nand I_58(n28_0,G42_7_r_16,n_573_7_r_16);
not I_59(n29_0,n32_0);
nor I_60(n30_0,n39_0,N1508_6_r_16);
not I_61(n31_0,n38_0);
nand I_62(n32_0,n41_0,n42_0);
nor I_63(n33_0,n_102_5_r_0,N1372_1_r_16);
nor I_64(n34_0,n27_0,N1372_1_r_16);
nand I_65(n35_0,n29_0,n36_0);
nor I_66(n36_0,n37_0,n38_0);
not I_67(n37_0,n28_0);
nand I_68(n38_0,n40_0,N1508_1_r_16);
nor I_69(n39_0,N1507_6_r_16,n_452_7_r_16);
or I_70(n40_0,N1507_6_r_16,n_452_7_r_16);
nor I_71(n41_0,n_572_7_r_16,n_569_7_r_16);
or I_72(n42_0,n43_0,N1371_0_r_16);
nor I_73(n43_0,N1508_0_r_16,N1372_1_r_16);
nor I_74(n44_0,n45_0,N1508_0_r_16);
and I_75(n45_0,N6147_2_r_16,N1371_0_r_16);
endmodule


