module test_I5334(I1477,I3685,I3877,I1976,I1470,I5334);
input I1477,I3685,I3877,I1976,I1470;
output I5334;
wire I3422,I3356,I1483,I5300,I3388,I3365,I5317,I5283,I1518,I3620,I3362,I1480,I1880,I3374,I3702;
or I_0(I3422,I1483,I1480);
DFFARX1 I_1(I1470,I3388,,,I3356,);
DFFARX1 I_2(I1880,I1470,I1518,,,I1483,);
nor I_3(I5300,I5283,I3374);
not I_4(I3388,I1477);
not I_5(I3365,I3702);
and I_6(I5317,I5300,I3365);
not I_7(I5283,I3356);
not I_8(I1518,I1477);
nor I_9(I3620,I1483);
DFFARX1 I_10(I3422,I1470,I3388,,,I3362,);
DFFARX1 I_11(I1976,I1470,I1518,,,I1480,);
or I_12(I5334,I5317,I3362);
DFFARX1 I_13(I1470,I1518,,,I1880,);
nand I_14(I3374,I3620,I3877);
DFFARX1 I_15(I3685,I1470,I3388,,,I3702,);
endmodule


