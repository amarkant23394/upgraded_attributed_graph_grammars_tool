module test_I3107(I1351,I1447,I1477,I1470,I1359,I1407,I3107);
input I1351,I1447,I1477,I1470,I1359,I1407;
output I3107;
wire I2759,I3076,I2844,I2827,I2776;
not I_0(I2759,I1477);
nor I_1(I3107,I3076,I2844);
DFFARX1 I_2(I1447,I1470,I2759,,,I3076,);
nand I_3(I2844,I2827,I1359);
nor I_4(I2827,I2776,I1351);
not I_5(I2776,I1407);
endmodule


