module test_I9689(I8267,I1477,I1470,I8377,I8315,I9689);
input I8267,I1477,I1470,I8377,I8315;
output I9689;
wire I8479,I8462,I8216,I9672,I8753,I8623,I8196,I9655,I8736,I8190,I9491,I8208;
nor I_0(I8479,I8462,I8315);
DFFARX1 I_1(I1470,I8216,,,I8462,);
not I_2(I8216,I1477);
and I_3(I9672,I9655,I8208);
not I_4(I8753,I8736);
DFFARX1 I_5(I1470,I8216,,,I8623,);
nand I_6(I8196,I8623,I8377);
nand I_7(I9655,I8190,I8196);
DFFARX1 I_8(I1470,I8216,,,I8736,);
DFFARX1 I_9(I9672,I1470,I9491,,,I9689,);
DFFARX1 I_10(I8267,I1470,I8216,,,I8190,);
not I_11(I9491,I1477);
nand I_12(I8208,I8753,I8479);
endmodule


