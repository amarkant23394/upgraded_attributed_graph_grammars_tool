module test_I8879(I7026,I1470,I6907,I5082,I8879);
input I7026,I1470,I6907,I5082;
output I8879;
wire I7427,I7317,I7057,I5067,I7410,I7269,I6887;
not I_0(I7427,I7410);
nor I_1(I7317,I7269,I7057);
not I_2(I7057,I7026);
DFFARX1 I_3(I1470,,,I5067,);
DFFARX1 I_4(I5082,I1470,I6907,,,I7410,);
not I_5(I8879,I6887);
DFFARX1 I_6(I5067,I1470,I6907,,,I7269,);
nand I_7(I6887,I7427,I7317);
endmodule


