module test_I3235(I1902,I1908,I1294,I1301,I3235);
input I1902,I1908,I1294,I1301;
output I3235;
wire I3263,I3622,I2668,I2962,I1914,I2583,I2651,I2569,I3246,I2566,I2945,I2702,I3543,I2832,I2572;
not I_0(I3263,I2569);
DFFARX1 I_1(I2572,I1294,I3246,,,I3622,);
nand I_2(I2668,I2651,I1914);
nor I_3(I2962,I2945,I2668);
DFFARX1 I_4(I1294,,,I1914,);
not I_5(I2583,I1301);
nor I_6(I2651,I1908);
nor I_7(I3235,I3622,I3543);
nand I_8(I2569,I2832,I2962);
not I_9(I3246,I1301);
not I_10(I2566,I2945);
DFFARX1 I_11(I1902,I1294,I2583,,,I2945,);
not I_12(I2702,I1908);
nand I_13(I3543,I3263,I2566);
DFFARX1 I_14(I1294,I2583,,,I2832,);
nor I_15(I2572,I2668,I2702);
endmodule


