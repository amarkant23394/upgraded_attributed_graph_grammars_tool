module test_I15160(I12930,I1477,I1470,I12882,I15160);
input I12930,I1477,I1470,I12882;
output I15160;
wire I12619,I13040,I13023,I12718,I10615,I10639,I15143,I12599,I13057,I12735,I12964,I12611;
not I_0(I12619,I1477);
nand I_1(I13040,I13023,I12735);
DFFARX1 I_2(I1470,I12619,,,I13023,);
nor I_3(I12718,I10615,I10639);
DFFARX1 I_4(I1470,,,I10615,);
DFFARX1 I_5(I1470,,,I10639,);
nor I_6(I15160,I15143,I12611);
not I_7(I15143,I12599);
nand I_8(I12599,I12718,I12964);
and I_9(I13057,I12718,I13040);
DFFARX1 I_10(I1470,I12619,,,I12735,);
nor I_11(I12964,I12930,I12882);
DFFARX1 I_12(I13057,I1470,I12619,,,I12611,);
endmodule


