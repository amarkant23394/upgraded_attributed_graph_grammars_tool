module test_I15976(I1477,I13860,I14066,I1470,I15976);
input I1477,I13860,I14066,I1470;
output I15976;
wire I14083,I15713,I13761,I15730,I13746,I13891,I13775,I15611,I15928;
DFFARX1 I_0(I14066,I1470,I13775,,,I14083,);
not I_1(I15713,I13761);
nand I_2(I13761,I13891,I13860);
not I_3(I15730,I15713);
not I_4(I13746,I14083);
DFFARX1 I_5(I1470,I13775,,,I13891,);
not I_6(I13775,I1477);
not I_7(I15611,I1477);
nor I_8(I15976,I15928,I15730);
DFFARX1 I_9(I13746,I1470,I15611,,,I15928,);
endmodule


