module test_I5994(I1477,I2695,I2170,I2557,I1470,I4725,I5994);
input I1477,I2695,I2170,I2557,I1470,I4725;
output I5994;
wire I4544,I4869,I2149,I4790,I2143,I4674,I2155,I4807,I2181,I4506,I4512,I4742,I4824,I4773;
not I_0(I4544,I1477);
DFFARX1 I_1(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_2(I2695,I1470,I2181,,,I2149,);
nor I_3(I4790,I4674,I4773);
nand I_4(I5994,I4512,I4506);
DFFARX1 I_5(I2557,I1470,I2181,,,I2143,);
DFFARX1 I_6(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_7(I1470,I2181,,,I2155,);
DFFARX1 I_8(I2170,I1470,I4544,,,I4807,);
not I_9(I2181,I1477);
nand I_10(I4506,I4869,I4773);
nand I_11(I4512,I4824,I4790);
DFFARX1 I_12(I4725,I1470,I4544,,,I4742,);
and I_13(I4824,I4807,I2143);
not I_14(I4773,I4742);
endmodule


