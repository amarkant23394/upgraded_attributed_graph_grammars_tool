module test_I7238(I7122,I5085,I1477,I5563,I5642,I5450,I1470,I7238);
input I7122,I5085,I1477,I5563,I5642,I5450,I1470;
output I7238;
wire I7173,I5659,I5088,I6907,I7221,I5097,I7139,I6975,I7009,I5073,I6992,I5105,I6924,I7156;
nor I_0(I7173,I7156,I7009);
or I_1(I5659,I5642,I5563);
DFFARX1 I_2(I5659,I1470,I5105,,,I5088,);
not I_3(I6907,I1477);
nand I_4(I7221,I6924,I5088);
nand I_5(I5097,I5642);
or I_6(I7139,I7122,I5085);
and I_7(I7238,I7221,I7173);
nor I_8(I6975,I6924);
not I_9(I7009,I6992);
DFFARX1 I_10(I5450,I1470,I5105,,,I5073,);
nand I_11(I6992,I6975,I5097);
not I_12(I5105,I1477);
not I_13(I6924,I5073);
DFFARX1 I_14(I7139,I1470,I6907,,,I7156,);
endmodule


