module test_I13186(I8851,I1477,I1470,I8848,I11751,I13186);
input I8851,I1477,I1470,I8848,I11751;
output I13186;
wire I11378,I13601,I11429,I11296,I13197,I11299,I11559,I11768,I11272,I11395,I13508,I11689,I13491,I11310;
nor I_0(I11378,I8848);
DFFARX1 I_1(I11299,I1470,I13197,,,I13601,);
not I_2(I11429,I8848);
nand I_3(I11296,I11559,I11689);
not I_4(I13197,I1477);
nor I_5(I11299,I11395,I11429);
DFFARX1 I_6(I1470,I11310,,,I11559,);
and I_7(I11768,I11429,I11751);
DFFARX1 I_8(I11768,I1470,I11310,,,I11272,);
nor I_9(I13186,I13601,I13508);
nand I_10(I11395,I11378,I8851);
and I_11(I13508,I13491,I11272);
nor I_12(I11689,I11395);
DFFARX1 I_13(I11296,I1470,I13197,,,I13491,);
not I_14(I11310,I1477);
endmodule


