module test_I7748(I1477,I1470,I4263,I4068,I7748);
input I1477,I1470,I4263,I4068;
output I7748;
wire I3948,I6329,I6688,I6705,I6291,I3972;
DFFARX1 I_0(I1470,,,I3948,);
not I_1(I6329,I1477);
DFFARX1 I_2(I3948,I1470,I6329,,,I6688,);
and I_3(I6705,I6688,I3972);
DFFARX1 I_4(I6705,I1470,I6329,,,I6291,);
or I_5(I3972,I4263,I4068);
not I_6(I7748,I6291);
endmodule


