module test_I6476(I1477,I1470,I4068,I3969,I6476);
input I1477,I1470,I4068,I3969;
output I6476;
wire I3963,I3975,I3954,I6346,I6442,I6363,I6380,I6329,I4308,I4181,I4034,I6459;
nor I_0(I3963,I4181,I4034);
nor I_1(I3975,I4308,I4034);
nor I_2(I6476,I6380,I6459);
not I_3(I3954,I4068);
nand I_4(I6346,I3969,I3954);
nor I_5(I6442,I3975,I3954);
and I_6(I6363,I6346,I3963);
DFFARX1 I_7(I6363,I1470,I6329,,,I6380,);
not I_8(I6329,I1477);
DFFARX1 I_9(I1470,,,I4308,);
DFFARX1 I_10(I1470,,,I4181,);
DFFARX1 I_11(I1470,,,I4034,);
not I_12(I6459,I6442);
endmodule


