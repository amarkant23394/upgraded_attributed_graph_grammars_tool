module test_final(IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_2,blif_reset_net_1_r_2,G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2);
input IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_2,blif_reset_net_1_r_2;
output G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2;
wire G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5,N3_2_l_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5,n_573_1_r_2,N3_2_l_2,n5_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2;
DFFARX1 I_0(n4_1_r_5,blif_clk_net_1_r_2,n5_2,G42_1_r_5,);
nor I_1(n_572_1_r_5,n21_5,n22_5);
nand I_2(n_573_1_r_5,n13_5,n16_5);
nor I_3(n_549_1_r_5,n21_5,n17_5);
nand I_4(n_569_1_r_5,n13_5,n15_5);
nor I_5(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_6(G199_2_l_5,blif_clk_net_1_r_2,n5_2,ACVQN2_3_r_5,);
nor I_7(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_8(n_42_2_l_5,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_5,);
not I_9(P6_5_r_5,P6_5_r_internal_5);
and I_10(N3_2_l_5,IN_6_2_l_5,n19_5);
DFFARX1 I_11(N3_2_l_5,blif_clk_net_1_r_2,n5_2,G199_2_l_5,);
DFFARX1 I_12(IN_1_3_l_5,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_5,);
not I_13(n13_5,ACVQN2_3_l_5);
DFFARX1 I_14(IN_2_3_l_5,blif_clk_net_1_r_2,n5_2,ACVQN1_3_l_5,);
and I_15(N1_4_l_5,IN_6_4_l_5,n20_5);
DFFARX1 I_16(N1_4_l_5,blif_clk_net_1_r_2,n5_2,n21_5,);
not I_17(n15_5,n21_5);
DFFARX1 I_18(IN_3_4_l_5,blif_clk_net_1_r_2,n5_2,n22_5,);
nor I_19(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_20(ACVQN2_3_l_5,blif_clk_net_1_r_2,n5_2,n11_internal_5,);
not I_21(n11_5,n11_internal_5);
nor I_22(n_42_2_l_5,IN_1_2_l_5,IN_3_2_l_5);
not I_23(n1_5,n18_5);
DFFARX1 I_24(n1_5,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_5,);
not I_25(n16_5,n_42_2_l_5);
nor I_26(n17_5,n22_5,n18_5);
nand I_27(n18_5,IN_4_3_l_5,ACVQN1_3_l_5);
nand I_28(n19_5,IN_2_2_l_5,IN_3_2_l_5);
nand I_29(n20_5,IN_1_4_l_5,IN_2_4_l_5);
DFFARX1 I_30(n4_1_r_2,blif_clk_net_1_r_2,n5_2,G42_1_r_2,);
nor I_31(n_572_1_r_2,n26_2,n18_2);
nand I_32(n_573_1_r_2,n17_2,n19_2);
nor I_33(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_34(n_569_1_r_2,n13_2,n19_2);
not I_35(n_452_1_r_2,n_573_1_r_2);
nor I_36(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_37(N3_2_r_2,blif_clk_net_1_r_2,n5_2,G199_2_r_2,);
DFFARX1 I_38(ACVQN2_3_l_2,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_2,);
not I_39(P6_5_r_2,P6_5_r_internal_2);
and I_40(N3_2_l_2,n24_2,n_572_1_r_5);
not I_41(n5_2,blif_reset_net_1_r_2);
DFFARX1 I_42(N3_2_l_2,blif_clk_net_1_r_2,n5_2,G199_2_l_2,);
not I_43(n13_2,G199_2_l_2);
DFFARX1 I_44(P6_5_r_5,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_2,);
DFFARX1 I_45(n_266_and_0_3_r_5,blif_clk_net_1_r_2,n5_2,n16_2,);
and I_46(N1_4_l_2,n25_2,n_549_1_r_5);
DFFARX1 I_47(N1_4_l_2,blif_clk_net_1_r_2,n5_2,n26_2,);
DFFARX1 I_48(n_573_1_r_5,blif_clk_net_1_r_2,n5_2,n17_internal_2,);
not I_49(n17_2,n17_internal_2);
nor I_50(n4_1_r_2,n26_2,n22_2);
nor I_51(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_52(G199_2_l_2,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_2,);
nor I_53(n18_2,G42_1_r_5,n_569_1_r_5);
nand I_54(n19_2,n16_2,ACVQN1_5_r_5);
nor I_55(n20_2,n26_2,n21_2);
not I_56(n21_2,n18_2);
and I_57(n22_2,n16_2,ACVQN1_5_r_5);
nor I_58(n23_2,n13_2,n21_2);
nand I_59(n24_2,n_569_1_r_5,G42_1_r_5);
nand I_60(n25_2,n_452_1_r_5,ACVQN2_3_r_5);
endmodule


