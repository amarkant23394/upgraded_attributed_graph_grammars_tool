module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_8_r_10,n11_10,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_10,n37_10,n38_10);
nor I_43(N1508_0_r_10,n37_10,n58_10);
nand I_44(N6147_2_r_10,n39_10,n40_10);
not I_45(N6147_3_r_10,n39_10);
nor I_46(N1372_4_r_10,n46_10,n49_10);
nor I_47(N1508_4_r_10,n51_10,n52_10);
nor I_48(N1507_6_r_10,n49_10,n60_10);
nor I_49(N1508_6_r_10,n49_10,n50_10);
nor I_50(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_51(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_52(N6147_9_r_10,n36_10,n37_10);
nor I_53(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_54(I_BUFF_1_9_r_10,n48_10);
nor I_55(N3_8_r_10,n44_10,n47_10);
not I_56(n11_10,blif_reset_net_8_r_10);
not I_57(n35_10,n49_10);
nor I_58(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_59(n37_10,N1507_6_r_11);
not I_60(n38_10,n46_10);
nand I_61(n39_10,n43_10,n44_10);
nand I_62(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_63(n41_10,n42_10,N1507_6_r_11);
not I_64(n42_10,n44_10);
nor I_65(n43_10,n45_10,N1507_6_r_11);
nand I_66(n44_10,n54_10,N6147_3_r_11);
nor I_67(n45_10,n59_10,N1508_1_r_11);
nand I_68(n46_10,n61_10,n_429_or_0_5_r_11);
nor I_69(n47_10,n46_10,n48_10);
nand I_70(n48_10,n62_10,n63_10);
nand I_71(n49_10,n56_10,n_547_5_r_11);
not I_72(n50_10,n45_10);
nor I_73(n51_10,n42_10,n53_10);
not I_74(n52_10,N1372_4_r_10);
nor I_75(n53_10,n48_10,n50_10);
and I_76(n54_10,n55_10,N6147_2_r_11);
nand I_77(n55_10,n56_10,n57_10);
nand I_78(n56_10,N1372_1_r_11,N1508_6_r_11);
not I_79(n57_10,n_547_5_r_11);
nor I_80(n58_10,n35_10,n45_10);
nor I_81(n59_10,n_576_5_r_11,N1372_1_r_11);
nor I_82(n60_10,n37_10,n46_10);
or I_83(n61_10,n_576_5_r_11,N1372_1_r_11);
nor I_84(n62_10,N1508_1_r_11,G78_5_r_11);
or I_85(n63_10,n64_10,N6147_2_r_11);
nor I_86(n64_10,N1508_10_r_11,N6147_3_r_11);
endmodule


