module Benchmark_testing100(I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I163,I170,I2006,I2087,I2123,I2294,I2312,I2339,I2429,I2519,I2537);
input I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I163,I170;
output I2006,I2087,I2123,I2294,I2312,I2339,I2429,I2519,I2537;
wire I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I163,I170,I179,I206,I224,I233,I251,I269,I287,I314,I323,I350,I359,I377,I395,I422,I431,I458,I467,I485,I503,I530,I539,I557,I575,I593,I620,I629,I647,I665,I683,I701,I728,I746,I755,I782,I800,I809,I836,I845,I863,I881,I899,I917,I935,I953,I980,I989,I1007,I1025,I1043,I1070,I1079,I1097,I1115,I1133,I1151,I1178,I1187,I1205,I1223,I1250,I1259,I1277,I1295,I1313,I1340,I1349,I1367,I1385,I1412,I1421,I1439,I1457,I1484,I1502,I1511,I1529,I1556,I1565,I1583,I1601,I1628,I1646,I1655,I1673,I1700,I1718,I1727,I1745,I1763,I1781,I1799,I1817,I1835,I1862,I1871,I1889,I1907,I1925,I1943,I1970,I1979,I2024,I2033,I2051,I2069,I2114,I2141,I2159,I2186,I2195,I2213,I2231,I2249,I2267,I2321,I2357,I2375,I2402,I2411,I2447,I2465,I2483,I2501;
not I_0 (I179,I170);
DFFARX1 I_1 (I108,I163,I179,I206,);
DFFARX1 I_2 (I206,I163,I179,I224,);
not I_3 (I233,I224);
not I_4 (I251,I206);
nand I_5 (I269,I148,I156);
and I_6 (I287,I269,I92);
DFFARX1 I_7 (I287,I163,I179,I314,);
not I_8 (I323,I314);
DFFARX1 I_9 (I124,I163,I179,I350,);
and I_10 (I359,I350,I100);
nand I_11 (I377,I350,I100);
nand I_12 (I395,I323,I377);
DFFARX1 I_13 (I84,I163,I179,I422,);
nor I_14 (I431,I422,I359);
DFFARX1 I_15 (I431,I163,I179,I458,);
nor I_16 (I467,I422,I314);
nand I_17 (I485,I76,I116);
and I_18 (I503,I485,I140);
DFFARX1 I_19 (I503,I163,I179,I530,);
nor I_20 (I539,I530,I422);
not I_21 (I557,I530);
nor I_22 (I575,I557,I323);
nor I_23 (I593,I251,I575);
DFFARX1 I_24 (I593,I163,I179,I620,);
nor I_25 (I629,I557,I422);
nor I_26 (I647,I132,I116);
nor I_27 (I665,I647,I629);
not I_28 (I683,I647);
nand I_29 (I701,I377,I683);
DFFARX1 I_30 (I647,I163,I179,I728,);
DFFARX1 I_31 (I647,I163,I179,I746,);
not I_32 (I755,I170);
DFFARX1 I_33 (I458,I163,I755,I782,);
DFFARX1 I_34 (I782,I163,I755,I800,);
not I_35 (I809,I800);
DFFARX1 I_36 (I728,I163,I755,I836,);
not I_37 (I845,I539);
nor I_38 (I863,I782,I845);
not I_39 (I881,I665);
not I_40 (I899,I467);
nand I_41 (I917,I899,I665);
nor I_42 (I935,I845,I917);
nor I_43 (I953,I836,I935);
DFFARX1 I_44 (I899,I163,I755,I980,);
nor I_45 (I989,I467,I233);
nand I_46 (I1007,I989,I746);
nor I_47 (I1025,I1007,I881);
nand I_48 (I1043,I1025,I539);
DFFARX1 I_49 (I1007,I163,I755,I1070,);
nand I_50 (I1079,I881,I467);
nor I_51 (I1097,I881,I467);
nand I_52 (I1115,I863,I1097);
not I_53 (I1133,I395);
nor I_54 (I1151,I1133,I1079);
DFFARX1 I_55 (I1151,I163,I755,I1178,);
nor I_56 (I1187,I1133,I458);
and I_57 (I1205,I1187,I620);
or I_58 (I1223,I1205,I701);
DFFARX1 I_59 (I1223,I163,I755,I1250,);
nor I_60 (I1259,I1250,I836);
nor I_61 (I1277,I782,I1259);
not I_62 (I1295,I1250);
nor I_63 (I1313,I1295,I953);
DFFARX1 I_64 (I1313,I163,I755,I1340,);
nand I_65 (I1349,I1295,I881);
nor I_66 (I1367,I1133,I1349);
not I_67 (I1385,I170);
DFFARX1 I_68 (I1367,I163,I1385,I1412,);
not I_69 (I1421,I1412);
nand I_70 (I1439,I809,I1070);
and I_71 (I1457,I1439,I1178);
DFFARX1 I_72 (I1457,I163,I1385,I1484,);
DFFARX1 I_73 (I1367,I163,I1385,I1502,);
and I_74 (I1511,I1502,I1115);
nor I_75 (I1529,I1484,I1511);
DFFARX1 I_76 (I1529,I163,I1385,I1556,);
nand I_77 (I1565,I1502,I1115);
nand I_78 (I1583,I1421,I1565);
not I_79 (I1601,I1583);
DFFARX1 I_80 (I1277,I163,I1385,I1628,);
DFFARX1 I_81 (I1628,I163,I1385,I1646,);
nand I_82 (I1655,I1340,I1043);
and I_83 (I1673,I1655,I1178);
DFFARX1 I_84 (I1673,I163,I1385,I1700,);
DFFARX1 I_85 (I1700,I163,I1385,I1718,);
not I_86 (I1727,I1718);
not I_87 (I1745,I1700);
nand I_88 (I1763,I1745,I1565);
nor I_89 (I1781,I980,I1043);
not I_90 (I1799,I1781);
nor I_91 (I1817,I1745,I1799);
nor I_92 (I1835,I1421,I1817);
DFFARX1 I_93 (I1835,I163,I1385,I1862,);
nor I_94 (I1871,I1484,I1799);
nor I_95 (I1889,I1700,I1871);
nor I_96 (I1907,I1628,I1781);
nor I_97 (I1925,I1484,I1781);
not I_98 (I1943,I170);
DFFARX1 I_99 (I1727,I163,I1943,I1970,);
and I_100 (I1979,I1970,I1556);
DFFARX1 I_101 (I1979,I163,I1943,I2006,);
DFFARX1 I_102 (I1862,I163,I1943,I2024,);
not I_103 (I2033,I1889);
not I_104 (I2051,I1925);
nand I_105 (I2069,I2051,I2033);
nor I_106 (I2087,I2024,I2069);
DFFARX1 I_107 (I2069,I163,I1943,I2114,);
not I_108 (I2123,I2114);
not I_109 (I2141,I1601);
nand I_110 (I2159,I2051,I2141);
DFFARX1 I_111 (I2159,I163,I1943,I2186,);
not I_112 (I2195,I2186);
not I_113 (I2213,I1925);
nand I_114 (I2231,I2213,I1646);
and I_115 (I2249,I2033,I2231);
nor I_116 (I2267,I2159,I2249);
DFFARX1 I_117 (I2267,I163,I1943,I2294,);
DFFARX1 I_118 (I2249,I163,I1943,I2312,);
nor I_119 (I2321,I1925,I1907);
nor I_120 (I2339,I2159,I2321);
or I_121 (I2357,I1925,I1907);
nor I_122 (I2375,I1763,I1556);
DFFARX1 I_123 (I2375,I163,I1943,I2402,);
not I_124 (I2411,I2402);
nor I_125 (I2429,I2411,I2195);
nand I_126 (I2447,I2411,I2024);
not I_127 (I2465,I1763);
nand I_128 (I2483,I2465,I2141);
nand I_129 (I2501,I2411,I2483);
nand I_130 (I2519,I2501,I2447);
nand I_131 (I2537,I2483,I2357);
endmodule


