module test_I10618(I9462,I10862,I1477,I1470,I10618);
input I9462,I10862,I1477,I1470;
output I10618;
wire I10879,I10647,I10896,I10930;
or I_0(I10879,I10862,I9462);
not I_1(I10647,I1477);
not I_2(I10618,I10930);
DFFARX1 I_3(I10879,I1470,I10647,,,I10896,);
DFFARX1 I_4(I10896,I1470,I10647,,,I10930,);
endmodule


