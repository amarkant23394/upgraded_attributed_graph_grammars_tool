module test_I2038(I1477,I1295,I1470,I2038);
input I1477,I1295,I1470;
output I2038;
wire I1518,I2021;
not I_0(I1518,I1477);
not I_1(I2038,I2021);
DFFARX1 I_2(I1295,I1470,I1518,,,I2021,);
endmodule


