module test_I5546(I1477,I3521,I3620,I1470,I1501,I5546);
input I1477,I3521,I3620,I1470,I1501;
output I5546;
wire I1486,I3470,I3637,I5512,I3747,I3388,I3846,I5122,I5204,I5187,I3380,I3453,I5105,I3368,I3350,I3353,I5529;
DFFARX1 I_0(I1470,,,I1486,);
not I_1(I3470,I3453);
DFFARX1 I_2(I3620,I1470,I3388,,,I3637,);
DFFARX1 I_3(I3368,I1470,I5105,,,I5512,);
DFFARX1 I_4(I1470,I3388,,,I3747,);
not I_5(I3388,I1477);
nor I_6(I5546,I5204,I5529);
nor I_7(I3846,I3747);
not I_8(I5122,I3350);
nand I_9(I5204,I5187,I3353);
nor I_10(I5187,I5122,I3380);
nand I_11(I3380,I3521,I3846);
nor I_12(I3453,I1486,I1501);
not I_13(I5105,I1477);
nand I_14(I3368,I3747,I3470);
DFFARX1 I_15(I1470,I3388,,,I3350,);
and I_16(I3353,I3453,I3637);
not I_17(I5529,I5512);
endmodule


