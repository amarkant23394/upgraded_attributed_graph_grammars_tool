module test_I6722(I2733,I1477,I2742,I6589,I1470,I6722);
input I2733,I1477,I2742,I6589,I1470;
output I6722;
wire I6640,I6442,I6705,I3972,I3983,I6510,I3954,I6329,I4068,I4263,I2724,I3975,I6688,I6493,I4308,I4452,I4034,I6606,I3948,I6623,I4246;
or I_0(I6722,I6705,I6640);
and I_1(I6640,I6442,I6623);
nor I_2(I6442,I3975,I3954);
and I_3(I6705,I6688,I3972);
or I_4(I3972,I4263,I4068);
not I_5(I3983,I1477);
not I_6(I6510,I6493);
not I_7(I3954,I4068);
not I_8(I6329,I1477);
nor I_9(I4068,I2742,I2724);
and I_10(I4263,I4246,I2733);
DFFARX1 I_11(I1470,,,I2724,);
nor I_12(I3975,I4308,I4034);
DFFARX1 I_13(I3948,I1470,I6329,,,I6688,);
DFFARX1 I_14(I1470,I6329,,,I6493,);
DFFARX1 I_15(I1470,I3983,,,I4308,);
or I_16(I4452,I4263);
DFFARX1 I_17(I1470,I3983,,,I4034,);
DFFARX1 I_18(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_19(I4452,I1470,I3983,,,I3948,);
nor I_20(I6623,I6606,I6510);
DFFARX1 I_21(I1470,I3983,,,I4246,);
endmodule


