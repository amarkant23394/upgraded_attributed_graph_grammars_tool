module test_I1926(I1239,I1207,I1294,I1492,I1301,I1704,I1223,I1926);
input I1239,I1207,I1294,I1492,I1301,I1704,I1223;
output I1926;
wire I2313,I1322,I2234,I1639,I1410,I1427,I1331,I1954,I1622,I1937,I1342,I1509,I1304;
DFFARX1 I_0(I1331,I1294,I1937,,,I2313,);
nand I_1(I1322,I1427,I1704);
nand I_2(I2234,I1954,I1304);
and I_3(I1639,I1622,I1207);
nor I_4(I1410,I1223,I1239);
DFFARX1 I_5(I1294,I1342,,,I1427,);
nor I_6(I1331,I1639,I1410);
not I_7(I1954,I1322);
nor I_8(I1926,I2313,I2234);
DFFARX1 I_9(I1294,I1342,,,I1622,);
not I_10(I1937,I1301);
not I_11(I1342,I1301);
DFFARX1 I_12(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_13(I1509,I1294,I1342,,,I1304,);
endmodule


