module test_I2678(I1231,I1477,I1470,I1239,I1287,I2678);
input I1231,I1477,I1470,I1239,I1287;
output I2678;
wire I2181,I2294,I2633;
not I_0(I2181,I1477);
nor I_1(I2294,I1287,I1231);
nand I_2(I2678,I2633,I2294);
DFFARX1 I_3(I1239,I1470,I2181,,,I2633,);
endmodule


