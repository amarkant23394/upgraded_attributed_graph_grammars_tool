module test_I16052(I11956,I1477,I14244,I1470,I16052);
input I11956,I1477,I14244,I1470;
output I16052;
wire I13752,I14162,I13775,I15611,I14049,I14261,I14278,I14066;
DFFARX1 I_0(I14278,I1470,I13775,,,I13752,);
DFFARX1 I_1(I1470,I13775,,,I14162,);
DFFARX1 I_2(I13752,I1470,I15611,,,I16052,);
not I_3(I13775,I1477);
not I_4(I15611,I1477);
DFFARX1 I_5(I1470,I13775,,,I14049,);
and I_6(I14261,I14162,I14244);
or I_7(I14278,I14066,I14261);
and I_8(I14066,I14049,I11956);
endmodule


