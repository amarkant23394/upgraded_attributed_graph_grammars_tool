module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_5_r_7,n6_7,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_7,n53_7,n52_7);
nor I_40(N1508_0_r_7,n51_7,n52_7);
nand I_41(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_42(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_43(n_576_5_r_7,n31_7,n32_7);
nor I_44(n_102_5_r_7,N1372_4_r_15,N1507_6_r_15);
nand I_45(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_46(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_47(n_572_7_r_7,n54_7,n33_7);
nand I_48(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_49(n_549_7_r_7,n53_7,n36_7);
nand I_50(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_51(n_452_7_r_7,N1508_1_r_15,n_547_5_r_15);
nor I_52(n4_7_l_7,N1508_4_r_15,n_576_5_r_15);
not I_53(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_54(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_55(n30_7,n53_7);
and I_56(N3_8_l_7,n50_7,N1508_1_r_15);
DFFARX1 I_57(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_58(n_431_5_r_7,n40_7,n41_7);
nor I_59(n4_7_r_7,n54_7,n49_7);
and I_60(n31_7,n_102_5_r_7,n39_7);
not I_61(n32_7,N1508_4_r_15);
nor I_62(n33_7,n34_7,N1372_4_r_15);
and I_63(n34_7,n35_7,G78_5_r_15);
not I_64(n35_7,n_429_or_0_5_r_15);
nor I_65(n36_7,n37_7,N1508_4_r_15);
or I_66(n37_7,n54_7,N1507_6_r_15);
or I_67(n38_7,n_547_5_r_15,N1508_6_r_15);
nor I_68(n39_7,n_452_7_r_7,n_429_or_0_5_r_15);
nand I_69(n40_7,n46_7,n47_7);
nand I_70(n41_7,n42_7,n43_7);
nor I_71(n42_7,n44_7,n45_7);
nor I_72(n43_7,n_547_5_r_15,N1508_6_r_15);
nor I_73(n44_7,n_429_or_0_5_r_15,n_576_5_r_15);
nor I_74(n45_7,N1372_4_r_15,N1508_4_r_15);
nand I_75(n46_7,n35_7,G78_5_r_15);
not I_76(n47_7,N1372_4_r_15);
or I_77(n48_7,n_452_7_r_7,n_429_or_0_5_r_15);
not I_78(n49_7,n_452_7_r_7);
nand I_79(n50_7,N1508_6_r_15,G78_5_r_15);
and I_80(n51_7,n_452_7_r_7,n45_7);
not I_81(n52_7,n44_7);
endmodule


