module test_I4017(I1415,I1447,I1477,I1470,I2861,I2776,I4017);
input I1415,I1447,I1477,I1470,I2861,I2776;
output I4017;
wire I2730,I2721,I2878,I2759,I3045,I3155,I4000,I3076,I2980,I2724;
not I_0(I2730,I3076);
nand I_1(I2721,I2980,I2878);
not I_2(I2878,I2861);
not I_3(I2759,I1477);
and I_4(I3045,I2861);
and I_5(I4017,I4000,I2730);
or I_6(I3155,I3076,I3045);
nand I_7(I4000,I2721,I2724);
DFFARX1 I_8(I1447,I1470,I2759,,,I3076,);
nand I_9(I2980,I2776,I1415);
DFFARX1 I_10(I3155,I1470,I2759,,,I2724,);
endmodule


