module test_I11935(I1477,I1470,I12157,I10017,I11935);
input I1477,I1470,I12157,I10017;
output I11935;
wire I12208,I10023,I10052,I10137,I11973,I12174,I12191;
DFFARX1 I_0(I12208,I1470,I11973,,,I11935,);
DFFARX1 I_1(I12191,I1470,I11973,,,I12208,);
DFFARX1 I_2(I10137,I1470,I10052,,,I10023,);
not I_3(I10052,I1477);
DFFARX1 I_4(I1470,I10052,,,I10137,);
not I_5(I11973,I1477);
and I_6(I12174,I12157,I10017);
or I_7(I12191,I12174,I10023);
endmodule


