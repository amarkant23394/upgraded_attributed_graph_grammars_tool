module test_I5283(I1477,I3504,I1470,I5283);
input I1477,I3504,I1470;
output I5283;
wire I3388,I3521,I3405,I3555,I3589,I1495,I3356,I3572;
not I_0(I3388,I1477);
nor I_1(I3521,I3504,I1495);
or I_2(I3405,I1495);
DFFARX1 I_3(I1470,I3388,,,I3555,);
and I_4(I3589,I3521,I3572);
DFFARX1 I_5(I1470,,,I1495,);
not I_6(I5283,I3356);
DFFARX1 I_7(I3589,I1470,I3388,,,I3356,);
nand I_8(I3572,I3555,I3405);
endmodule


