module test_I8411(I1477,I4533,I1470,I4691,I8411);
input I1477,I4533,I1470,I4691;
output I8411;
wire I8394,I6203,I5713,I5751,I4518,I5725,I6127,I6110,I4869;
not I_0(I8394,I5713);
DFFARX1 I_1(I4518,I1470,I5751,,,I6203,);
DFFARX1 I_2(I6127,I1470,I5751,,,I5713,);
not I_3(I5751,I1477);
nor I_4(I8411,I8394,I5725);
nand I_5(I4518,I4869,I4691);
DFFARX1 I_6(I6203,I1470,I5751,,,I5725,);
and I_7(I6127,I6110,I4533);
DFFARX1 I_8(I1470,I5751,,,I6110,);
DFFARX1 I_9(I1470,,,I4869,);
endmodule


