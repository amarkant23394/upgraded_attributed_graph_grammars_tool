module test_I12493(I1477,I10202,I10120,I10349,I10414,I12106,I1470,I12493);
input I1477,I10202,I10120,I10349,I10414,I12106,I1470;
output I12493;
wire I12123,I10032,I10219,I12476,I10014,I10041,I12425,I10052,I12270,I12349,I11990,I10137,I11973,I12442,I12459;
not I_0(I12123,I12106);
nand I_1(I10032,I10137,I10414);
DFFARX1 I_2(I10202,I1470,I10052,,,I10219,);
and I_3(I12476,I12349,I12459);
DFFARX1 I_4(I10219,I1470,I10052,,,I10014,);
nor I_5(I10041,I10349,I10120);
DFFARX1 I_6(I1470,I11973,,,I12425,);
not I_7(I10052,I1477);
nand I_8(I12270,I11990,I10014);
DFFARX1 I_9(I10041,I1470,I11973,,,I12349,);
or I_10(I12493,I12270,I12476);
not I_11(I11990,I10032);
DFFARX1 I_12(I1470,I10052,,,I10137,);
not I_13(I11973,I1477);
not I_14(I12442,I12425);
nor I_15(I12459,I12442,I12123);
endmodule


