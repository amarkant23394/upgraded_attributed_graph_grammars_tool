module test_I9926(I8479,I8753,I1477,I8196,I1470,I9926);
input I8479,I8753,I1477,I8196,I1470;
output I9926;
wire I9491,I9816,I8705,I9909,I9655,I9689,I8193,I8190,I9672,I8208;
nor I_0(I9926,I9689,I9909);
not I_1(I9491,I1477);
DFFARX1 I_2(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_3(I1470,,,I8705,);
not I_4(I9909,I9816);
nand I_5(I9655,I8190,I8196);
DFFARX1 I_6(I9672,I1470,I9491,,,I9689,);
not I_7(I8193,I8705);
DFFARX1 I_8(I1470,,,I8190,);
and I_9(I9672,I9655,I8208);
nand I_10(I8208,I8753,I8479);
endmodule


