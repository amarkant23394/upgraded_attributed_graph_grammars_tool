module test_final(IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_6,blif_reset_net_1_r_6,G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6);
input IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_6_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_4_3_l_5,IN_1_4_l_5,IN_2_4_l_5,IN_3_4_l_5,IN_6_4_l_5,blif_clk_net_1_r_6,blif_reset_net_1_r_6;
output G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6;
wire G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5,N3_2_l_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5,N3_2_l_6,n4_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6;
DFFARX1 I_0(n4_1_r_5,blif_clk_net_1_r_6,n4_6,G42_1_r_5,);
nor I_1(n_572_1_r_5,n21_5,n22_5);
nand I_2(n_573_1_r_5,n13_5,n16_5);
nor I_3(n_549_1_r_5,n21_5,n17_5);
nand I_4(n_569_1_r_5,n13_5,n15_5);
nor I_5(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_6(G199_2_l_5,blif_clk_net_1_r_6,n4_6,ACVQN2_3_r_5,);
nor I_7(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_8(n_42_2_l_5,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_5,);
not I_9(P6_5_r_5,P6_5_r_internal_5);
and I_10(N3_2_l_5,IN_6_2_l_5,n19_5);
DFFARX1 I_11(N3_2_l_5,blif_clk_net_1_r_6,n4_6,G199_2_l_5,);
DFFARX1 I_12(IN_1_3_l_5,blif_clk_net_1_r_6,n4_6,ACVQN2_3_l_5,);
not I_13(n13_5,ACVQN2_3_l_5);
DFFARX1 I_14(IN_2_3_l_5,blif_clk_net_1_r_6,n4_6,ACVQN1_3_l_5,);
and I_15(N1_4_l_5,IN_6_4_l_5,n20_5);
DFFARX1 I_16(N1_4_l_5,blif_clk_net_1_r_6,n4_6,n21_5,);
not I_17(n15_5,n21_5);
DFFARX1 I_18(IN_3_4_l_5,blif_clk_net_1_r_6,n4_6,n22_5,);
nor I_19(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_20(ACVQN2_3_l_5,blif_clk_net_1_r_6,n4_6,n11_internal_5,);
not I_21(n11_5,n11_internal_5);
nor I_22(n_42_2_l_5,IN_1_2_l_5,IN_3_2_l_5);
not I_23(n1_5,n18_5);
DFFARX1 I_24(n1_5,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_5,);
not I_25(n16_5,n_42_2_l_5);
nor I_26(n17_5,n22_5,n18_5);
nand I_27(n18_5,IN_4_3_l_5,ACVQN1_3_l_5);
nand I_28(n19_5,IN_2_2_l_5,IN_3_2_l_5);
nand I_29(n20_5,IN_1_4_l_5,IN_2_4_l_5);
DFFARX1 I_30(n4_1_r_6,blif_clk_net_1_r_6,n4_6,G42_1_r_6,);
nor I_31(n_572_1_r_6,n27_6,n28_6);
nand I_32(n_573_1_r_6,n18_6,n19_6);
nor I_33(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_34(n_569_1_r_6,n19_6,n20_6);
nor I_35(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_36(N1_4_r_6,blif_clk_net_1_r_6,n4_6,G199_4_r_6,);
DFFARX1 I_37(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,G214_4_r_6,);
DFFARX1 I_38(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_6,);
not I_39(P6_5_r_6,P6_5_r_internal_6);
and I_40(N3_2_l_6,n23_6,ACVQN1_5_r_5);
not I_41(n4_6,blif_reset_net_1_r_6);
DFFARX1 I_42(N3_2_l_6,blif_clk_net_1_r_6,n4_6,n27_6,);
not I_43(n17_6,n27_6);
DFFARX1 I_44(n_569_1_r_5,blif_clk_net_1_r_6,n4_6,n28_6,);
DFFARX1 I_45(n_572_1_r_5,blif_clk_net_1_r_6,n4_6,n26_6,);
and I_46(N1_4_l_6,n25_6,G42_1_r_5);
DFFARX1 I_47(N1_4_l_6,blif_clk_net_1_r_6,n4_6,n29_6,);
not I_48(n18_6,n29_6);
DFFARX1 I_49(P6_5_r_5,blif_clk_net_1_r_6,n4_6,G214_4_l_6,);
not I_50(n12_6,G214_4_l_6);
nor I_51(n4_1_r_6,n28_6,n22_6);
nor I_52(N1_4_r_6,n12_6,n24_6);
nor I_53(n_42_2_l_6,n_573_1_r_5,n_266_and_0_3_r_5);
DFFARX1 I_54(G214_4_l_6,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_6,);
nand I_55(n19_6,n26_6,ACVQN2_3_r_5);
not I_56(n20_6,n_42_2_l_6);
nor I_57(n21_6,n17_6,n28_6);
and I_58(n22_6,n26_6,ACVQN2_3_r_5);
nand I_59(n23_6,G42_1_r_5,n_266_and_0_3_r_5);
nor I_60(n24_6,n17_6,n18_6);
nand I_61(n25_6,n_549_1_r_5,n_452_1_r_5);
endmodule


