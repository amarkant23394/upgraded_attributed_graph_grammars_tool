module test_I2389(I1255,I1376,I1215,I1207,I1294,I1301,I2389);
input I1255,I1376,I1215,I1207,I1294,I1301;
output I2389;
wire I1328,I1622,I1937,I1342,I1393,I1828,I1639,I1780;
nand I_0(I1328,I1639,I1828);
DFFARX1 I_1(I1255,I1294,I1342,,,I1622,);
not I_2(I1937,I1301);
not I_3(I1342,I1301);
DFFARX1 I_4(I1376,I1294,I1342,,,I1393,);
nor I_5(I1828,I1780,I1393);
DFFARX1 I_6(I1328,I1294,I1937,,,I2389,);
and I_7(I1639,I1622,I1207);
DFFARX1 I_8(I1215,I1294,I1342,,,I1780,);
endmodule


