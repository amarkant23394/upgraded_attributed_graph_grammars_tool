module test_I16240_rst(I1477_rst,I16240_rst);
,I16240_rst);
input I1477_rst;
output I16240_rst;
wire ;
not I_0(I16240_rst,I1477_rst);
endmodule


