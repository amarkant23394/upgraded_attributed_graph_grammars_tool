module test_I16869(I15064,I1477,I1470,I16869);
input I15064,I1477,I1470;
output I16869;
wire I14948,I15502,I15211,I14936,I16835,I16818,I16852,I15519,I14965,I15228,I15485,I14957;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
not I_1(I15502,I15485);
DFFARX1 I_2(I1470,I14965,,,I15211,);
DFFARX1 I_3(I15064,I1470,I14965,,,I14936,);
nand I_4(I16835,I14936,I14948);
DFFARX1 I_5(I16852,I1470,I16818,,,I16869,);
not I_6(I16818,I1477);
and I_7(I16852,I16835,I14957);
or I_8(I15519,I15502);
not I_9(I14965,I1477);
nor I_10(I15228,I15211,I15064);
DFFARX1 I_11(I1470,I14965,,,I15485,);
nand I_12(I14957,I15502,I15228);
endmodule


