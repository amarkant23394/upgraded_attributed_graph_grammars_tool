module test_final(G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G18_1_l_15,G15_1_l_15,IN_1_1_l_15,IN_4_1_l_15,IN_5_1_l_15,IN_7_1_l_15,IN_9_1_l_15,IN_10_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_4_3_l_15,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,n_452_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15,n4_1_l_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n_452_1_r_15,blif_clk_net_1_r_7,n8_7,G42_1_r_15,);
and I_1(n_572_1_r_15,n17_15,n19_15);
nand I_2(n_573_1_r_15,n15_15,n18_15);
nor I_3(n_549_1_r_15,n21_15,n22_15);
nand I_4(n_569_1_r_15,n15_15,n20_15);
nor I_5(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_6(G42_1_l_15,blif_clk_net_1_r_7,n8_7,ACVQN2_3_r_15,);
nor I_7(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_8(N1_4_r_15,blif_clk_net_1_r_7,n8_7,G199_4_r_15,);
DFFARX1 I_9(n_573_1_l_15,blif_clk_net_1_r_7,n8_7,G214_4_r_15,);
nor I_10(n4_1_l_15,G18_1_l_15,IN_1_1_l_15);
DFFARX1 I_11(n4_1_l_15,blif_clk_net_1_r_7,n8_7,G42_1_l_15,);
not I_12(n15_15,G42_1_l_15);
DFFARX1 I_13(IN_1_3_l_15,blif_clk_net_1_r_7,n8_7,n17_internal_15,);
not I_14(n17_15,n17_internal_15);
DFFARX1 I_15(IN_2_3_l_15,blif_clk_net_1_r_7,n8_7,n30_15,);
nor I_16(n_572_1_l_15,G15_1_l_15,IN_7_1_l_15);
DFFARX1 I_17(n_572_1_l_15,blif_clk_net_1_r_7,n8_7,n14_internal_15,);
not I_18(n14_15,n14_internal_15);
nand I_19(N1_4_r_15,n25_15,n26_15);
or I_20(n_573_1_l_15,IN_5_1_l_15,IN_9_1_l_15);
nor I_21(n18_15,IN_9_1_l_15,IN_10_1_l_15);
nand I_22(n19_15,n27_15,n28_15);
nand I_23(n20_15,IN_4_3_l_15,n30_15);
not I_24(n21_15,n20_15);
and I_25(n22_15,n17_15,n_572_1_l_15);
nor I_26(n23_15,G18_1_l_15,IN_5_1_l_15);
or I_27(n24_15,IN_9_1_l_15,IN_10_1_l_15);
or I_28(n25_15,G18_1_l_15,n_573_1_l_15);
nand I_29(n26_15,n19_15,n23_15);
not I_30(n27_15,IN_10_1_l_15);
nand I_31(n28_15,IN_4_1_l_15,n29_15);
not I_32(n29_15,G15_1_l_15);
DFFARX1 I_33(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_34(n_572_1_r_7,n30_7,n31_7);
nand I_35(n_573_1_r_7,n28_7,n_572_1_r_15);
nor I_36(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_37(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_38(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_39(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_40(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_41(P6_5_r_7,P6_5_r_internal_7);
or I_42(n_431_0_l_7,n36_7,n_266_and_0_3_r_15);
not I_43(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_44(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_45(n27_7,n43_7);
DFFARX1 I_46(n_549_1_r_15,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_47(ACVQN2_3_r_15,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_48(n4_1_r_7,n30_7,n38_7);
nor I_49(N1_4_r_7,n27_7,n40_7);
nand I_50(n26_7,n39_7,G199_4_r_15);
not I_51(n5_7,n_569_1_r_15);
DFFARX1 I_52(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_53(n28_7,n26_7,n29_7);
not I_54(n29_7,n_573_1_r_15);
not I_55(n30_7,G42_1_r_15);
nand I_56(n31_7,n27_7,n29_7);
nor I_57(n32_7,ACVQN1_5_l_7,n34_7);
nor I_58(n33_7,n29_7,n_569_1_r_15);
not I_59(n34_7,n_572_1_r_15);
nor I_60(n35_7,n43_7,n44_7);
and I_61(n36_7,n37_7,G42_1_r_15);
nor I_62(n37_7,n30_7,G214_4_r_15);
nand I_63(n38_7,n29_7,n_569_1_r_15);
nor I_64(n39_7,n_569_1_r_15,n_572_1_r_15);
nor I_65(n40_7,n44_7,n41_7);
nor I_66(n41_7,n34_7,n42_7);
nand I_67(n42_7,n5_7,n_573_1_r_15);
endmodule


