module test_I10766(I8216,I8753,I1470,I8193,I9491,I10766);
input I8216,I8753,I1470,I8193,I9491;
output I10766;
wire I9477,I8187,I9542,I9754,I9816,I9559,I9771,I8178,I9833;
nor I_0(I9477,I9771,I9833);
DFFARX1 I_1(I1470,I8216,,,I8187,);
DFFARX1 I_2(I1470,I9491,,,I9542,);
DFFARX1 I_3(I8187,I1470,I9491,,,I9754,);
DFFARX1 I_4(I8193,I1470,I9491,,,I9816,);
not I_5(I9559,I9542);
not I_6(I10766,I9477);
and I_7(I9771,I9754,I8178);
DFFARX1 I_8(I8753,I1470,I8216,,,I8178,);
and I_9(I9833,I9816,I9559);
endmodule


