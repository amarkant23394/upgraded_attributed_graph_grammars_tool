module test_I3453(I1477,I1470,I1207,I1455,I1383,I3453);
input I1477,I1470,I1207,I1455,I1383;
output I3453;
wire I1518,I1486,I1880,I1501,I1832,I1535;
not I_0(I1518,I1477);
DFFARX1 I_1(I1832,I1470,I1518,,,I1486,);
DFFARX1 I_2(I1383,I1470,I1518,,,I1880,);
not I_3(I1501,I1880);
nor I_4(I3453,I1486,I1501);
nand I_5(I1832,I1535,I1207);
not I_6(I1535,I1455);
endmodule


