module test_I1480(I1463,I1477,I1215,I1470,I1383,I1480);
input I1463,I1477,I1215,I1470,I1383;
output I1480;
wire I1518,I1637,I1552,I1976,I1880,I1569,I1959;
not I_0(I1518,I1477);
not I_1(I1637,I1215);
nor I_2(I1552,I1215);
DFFARX1 I_3(I1976,I1470,I1518,,,I1480,);
and I_4(I1976,I1637,I1959);
DFFARX1 I_5(I1383,I1470,I1518,,,I1880,);
nand I_6(I1569,I1552,I1463);
nand I_7(I1959,I1880,I1569);
endmodule


