module test_I5139(I3487,I1477,I1470,I1489,I2103,I3538,I1897,I5139);
input I3487,I1477,I1470,I1489,I2103,I3538,I1897;
output I5139;
wire I1518,I3388,I1504,I3846,I3521,I3380,I3504,I1495,I3555,I3747,I3359,I1767;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
nand I_2(I1504,I1767,I1897);
nor I_3(I3846,I3747,I3555);
nor I_4(I3521,I3504,I1495);
nand I_5(I3380,I3521,I3846);
and I_6(I3504,I3487,I1489);
DFFARX1 I_7(I2103,I1470,I1518,,,I1495,);
DFFARX1 I_8(I3538,I1470,I3388,,,I3555,);
nor I_9(I5139,I3380,I3359);
DFFARX1 I_10(I1504,I1470,I3388,,,I3747,);
DFFARX1 I_11(I3747,I1470,I3388,,,I3359,);
DFFARX1 I_12(I1470,I1518,,,I1767,);
endmodule


