module test_I5088(I3368,I1477,I5204,I1470,I3377,I5088);
input I3368,I1477,I5204,I1470,I3377;
output I5088;
wire I5659,I5625,I5546,I5563,I5529,I5512,I5105,I5642;
or I_0(I5659,I5642,I5563);
DFFARX1 I_1(I3377,I1470,I5105,,,I5625,);
nor I_2(I5546,I5204,I5529);
DFFARX1 I_3(I5659,I1470,I5105,,,I5088,);
and I_4(I5563,I5512,I5546);
not I_5(I5529,I5512);
DFFARX1 I_6(I3368,I1470,I5105,,,I5512,);
not I_7(I5105,I1477);
not I_8(I5642,I5625);
endmodule


