module test_I10639(I9465,I1477,I9771,I1470,I9737,I9471,I10639);
input I9465,I1477,I9771,I1470,I9737,I9471;
output I10639;
wire I10647,I10715,I10961,I11184,I10664,I11167,I9459,I11201,I11150,I10732;
not I_0(I10647,I1477);
nor I_1(I10715,I10664);
nand I_2(I10961,I10664,I9459);
nand I_3(I11184,I11167,I10732);
not I_4(I10664,I9471);
not I_5(I11167,I11150);
DFFARX1 I_6(I11201,I1470,I10647,,,I10639,);
nand I_7(I9459,I9771,I9737);
and I_8(I11201,I10961,I11184);
DFFARX1 I_9(I1470,I10647,,,I11150,);
nand I_10(I10732,I10715,I9465);
endmodule


