module test_I1716(I1207,I1367,I1716);
input I1207,I1367;
output I1716;
wire I1699;
nor I_0(I1716,I1699,I1367);
not I_1(I1699,I1207);
endmodule


