module test_I6589(I2733,I2727,I1477,I1470,I2751,I6589);
input I2733,I2727,I1477,I1470,I2751;
output I6589;
wire I3945,I3960,I3951,I4246,I4113,I6572,I4263,I4308,I4181,I4229,I4212,I4356,I3983;
nand I_0(I3945,I4308,I4212);
DFFARX1 I_1(I4356,I1470,I3983,,,I3960,);
nand I_2(I3951,I4263,I4229);
DFFARX1 I_3(I1470,I3983,,,I4246,);
and I_4(I6589,I6572,I3960);
DFFARX1 I_5(I2751,I1470,I3983,,,I4113,);
nand I_6(I6572,I3951,I3945);
and I_7(I4263,I4246,I2733);
DFFARX1 I_8(I2727,I1470,I3983,,,I4308,);
DFFARX1 I_9(I1470,I3983,,,I4181,);
nor I_10(I4229,I4113,I4212);
not I_11(I4212,I4181);
nor I_12(I4356,I4308,I4113);
not I_13(I3983,I1477);
endmodule


