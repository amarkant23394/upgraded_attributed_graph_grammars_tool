module test_final(IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_1_l_13,IN_2_1_l_13,IN_3_1_l_13,G18_7_l_13,G15_7_l_13,IN_1_7_l_13,IN_4_7_l_13,IN_5_7_l_13,IN_7_7_l_13,IN_9_7_l_13,IN_10_7_l_13,IN_1_10_l_13,IN_2_10_l_13,IN_3_10_l_13,IN_4_10_l_13,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_102_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13,n4_7_l_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
nor I_0(N1371_0_r_13,n59_13,n61_13);
nor I_1(N1508_0_r_13,n59_13,n60_13);
not I_2(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_3(n_431_5_r_13,blif_clk_net_7_r_16,n8_16,G78_5_r_13,);
nand I_4(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_5(n_102_5_r_13,IN_9_7_l_13,IN_10_7_l_13);
nand I_6(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_7(n1_13,blif_clk_net_7_r_16,n8_16,G42_7_r_13,);
nor I_8(n_572_7_r_13,n40_13,n41_13);
nand I_9(n_573_7_r_13,n37_13,n38_13);
nor I_10(n_549_7_r_13,n46_13,n47_13);
nand I_11(n_569_7_r_13,n37_13,n43_13);
nand I_12(n_452_7_r_13,n52_13,n53_13);
nor I_13(n4_7_l_13,G18_7_l_13,IN_1_7_l_13);
DFFARX1 I_14(n4_7_l_13,blif_clk_net_7_r_16,n8_16,n62_13,);
not I_15(n33_13,n62_13);
nand I_16(n_431_5_r_13,n54_13,n55_13);
not I_17(n1_13,n52_13);
nor I_18(n34_13,n35_13,n36_13);
nor I_19(n35_13,G15_7_l_13,n42_13);
nand I_20(n36_13,n50_13,n58_13);
nand I_21(n37_13,n44_13,n45_13);
or I_22(n38_13,IN_3_1_l_13,n39_13);
nand I_23(n39_13,IN_1_1_l_13,IN_2_1_l_13);
not I_24(n40_13,n36_13);
nor I_25(n41_13,IN_10_7_l_13,n35_13);
not I_26(n42_13,IN_4_7_l_13);
or I_27(n43_13,G18_7_l_13,IN_5_7_l_13);
not I_28(n44_13,G15_7_l_13);
not I_29(n45_13,IN_7_7_l_13);
nor I_30(n46_13,n39_13,n40_13);
nor I_31(n47_13,G18_7_l_13,IN_5_7_l_13);
nor I_32(n48_13,n50_13,n51_13);
nor I_33(n49_13,G15_7_l_13,IN_7_7_l_13);
not I_34(n50_13,n59_13);
not I_35(n51_13,n_102_5_r_13);
nand I_36(n52_13,n33_13,n39_13);
nand I_37(n53_13,IN_3_1_l_13,n33_13);
nor I_38(n54_13,IN_5_7_l_13,IN_9_7_l_13);
nand I_39(n55_13,n62_13,n56_13);
nor I_40(n56_13,n39_13,n57_13);
not I_41(n57_13,G18_7_l_13);
or I_42(n58_13,IN_3_10_l_13,IN_4_10_l_13);
nand I_43(n59_13,IN_1_10_l_13,IN_2_10_l_13);
nor I_44(n60_13,IN_5_7_l_13,n51_13);
nor I_45(n61_13,IN_3_1_l_13,n39_13);
nor I_46(N1371_0_r_16,n35_16,n39_16);
nor I_47(N1508_0_r_16,n39_16,n46_16);
not I_48(N1372_1_r_16,n45_16);
nor I_49(N1508_1_r_16,n53_16,n45_16);
nor I_50(N6147_2_r_16,n37_16,n38_16);
nor I_51(N1507_6_r_16,n44_16,n49_16);
nor I_52(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_53(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_54(n_572_7_r_16,n32_16,n33_16);
nand I_55(n_573_7_r_16,n30_16,n31_16);
nand I_56(n_549_7_r_16,n47_16,G42_7_r_13);
nand I_57(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_58(n_452_7_r_16,n34_16,n35_16);
and I_59(N3_8_l_16,n41_16,n_452_7_r_13);
not I_60(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_61(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_62(n29_16,n53_16);
nor I_63(n4_7_r_16,n35_16,n36_16);
nand I_64(n30_16,n_429_or_0_5_r_13,N1371_0_r_13);
not I_65(n31_16,n34_16);
nor I_66(n32_16,n30_16,n_576_5_r_13);
not I_67(n33_16,n_549_7_r_16);
nor I_68(n34_16,n48_16,n_429_or_0_5_r_13);
and I_69(n35_16,n50_16,N1508_0_r_13);
not I_70(n36_16,n30_16);
nor I_71(n37_16,n31_16,n40_16);
nand I_72(n38_16,n29_16,n39_16);
not I_73(n39_16,n32_16);
nor I_74(n40_16,G78_5_r_13,n_549_7_r_13);
nand I_75(n41_16,n_547_5_r_13,n_549_7_r_13);
nand I_76(n42_16,n35_16,n43_16);
not I_77(n43_16,n44_16);
nor I_78(n44_16,n32_16,n49_16);
nand I_79(n45_16,n36_16,n40_16);
nor I_80(n46_16,n33_16,n34_16);
nand I_81(n47_16,N1371_0_r_13,n_573_7_r_13);
or I_82(n48_16,n_569_7_r_13,N1508_0_r_13);
and I_83(n49_16,n35_16,n36_16);
and I_84(n50_16,n51_16,n_572_7_r_13);
nand I_85(n51_16,n47_16,n52_16);
not I_86(n52_16,G42_7_r_13);
endmodule


