module test_I2963(I1391,I1263,I1477,I1470,I2895,I1311,I2963);
input I1391,I1263,I1477,I1470,I2895,I1311;
output I2963;
wire I2759,I2946,I2929,I2912;
not I_0(I2759,I1477);
or I_1(I2946,I2929,I1263);
and I_2(I2929,I2912,I1391);
DFFARX1 I_3(I2946,I1470,I2759,,,I2963,);
nor I_4(I2912,I2895,I1311);
endmodule


