module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7,n_452_7_r_7,n4_7_l_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_7,n53_7,n52_7);
nor I_1(N1508_0_r_7,n51_7,n52_7);
nand I_2(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_3(n_431_5_r_7,blif_clk_net_8_r_10,n11_10,G78_5_r_7,);
nand I_4(n_576_5_r_7,n31_7,n32_7);
nor I_5(n_102_5_r_7,IN_5_7_l_7,IN_9_7_l_7);
nand I_6(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_7(n4_7_r_7,blif_clk_net_8_r_10,n11_10,G42_7_r_7,);
nor I_8(n_572_7_r_7,n54_7,n33_7);
nand I_9(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_10(n_549_7_r_7,n53_7,n36_7);
nand I_11(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_12(n_452_7_r_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_13(n4_7_l_7,G18_7_l_7,IN_1_7_l_7);
DFFARX1 I_14(n4_7_l_7,blif_clk_net_8_r_10,n11_10,n53_7,);
not I_15(n30_7,n53_7);
and I_16(N3_8_l_7,IN_6_8_l_7,n50_7);
DFFARX1 I_17(N3_8_l_7,blif_clk_net_8_r_10,n11_10,n54_7,);
nand I_18(n_431_5_r_7,n40_7,n41_7);
nor I_19(n4_7_r_7,n54_7,n49_7);
and I_20(n31_7,n_102_5_r_7,n39_7);
not I_21(n32_7,G18_7_l_7);
nor I_22(n33_7,IN_10_7_l_7,n34_7);
and I_23(n34_7,IN_4_7_l_7,n35_7);
not I_24(n35_7,G15_7_l_7);
nor I_25(n36_7,G18_7_l_7,n37_7);
or I_26(n37_7,IN_5_7_l_7,n54_7);
or I_27(n38_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_28(n39_7,IN_3_1_l_7,n_452_7_r_7);
nand I_29(n40_7,n46_7,n47_7);
nand I_30(n41_7,n42_7,n43_7);
nor I_31(n42_7,n44_7,n45_7);
nor I_32(n43_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_33(n44_7,G15_7_l_7,IN_7_7_l_7);
nor I_34(n45_7,IN_9_7_l_7,IN_10_7_l_7);
nand I_35(n46_7,IN_4_7_l_7,n35_7);
not I_36(n47_7,IN_10_7_l_7);
or I_37(n48_7,IN_3_1_l_7,n_452_7_r_7);
not I_38(n49_7,n_452_7_r_7);
nand I_39(n50_7,IN_2_8_l_7,IN_3_8_l_7);
and I_40(n51_7,n_452_7_r_7,n45_7);
not I_41(n52_7,n44_7);
nor I_42(N1371_0_r_10,n37_10,n38_10);
nor I_43(N1508_0_r_10,n37_10,n58_10);
nand I_44(N6147_2_r_10,n39_10,n40_10);
not I_45(N6147_3_r_10,n39_10);
nor I_46(N1372_4_r_10,n46_10,n49_10);
nor I_47(N1508_4_r_10,n51_10,n52_10);
nor I_48(N1507_6_r_10,n49_10,n60_10);
nor I_49(N1508_6_r_10,n49_10,n50_10);
nor I_50(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_51(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_52(N6147_9_r_10,n36_10,n37_10);
nor I_53(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_54(I_BUFF_1_9_r_10,n48_10);
nor I_55(N3_8_r_10,n44_10,n47_10);
not I_56(n11_10,blif_reset_net_8_r_10);
not I_57(n35_10,n49_10);
nor I_58(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_59(n37_10,N1371_0_r_7);
not I_60(n38_10,n46_10);
nand I_61(n39_10,n43_10,n44_10);
nand I_62(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_63(n41_10,n42_10,N1371_0_r_7);
not I_64(n42_10,n44_10);
nor I_65(n43_10,n45_10,N1371_0_r_7);
nand I_66(n44_10,n54_10,G78_5_r_7);
nor I_67(n45_10,n59_10,G78_5_r_7);
nand I_68(n46_10,n61_10,N1371_0_r_7);
nor I_69(n47_10,n46_10,n48_10);
nand I_70(n48_10,n62_10,n63_10);
nand I_71(n49_10,n56_10,n_429_or_0_5_r_7);
not I_72(n50_10,n45_10);
nor I_73(n51_10,n42_10,n53_10);
not I_74(n52_10,N1372_4_r_10);
nor I_75(n53_10,n48_10,n50_10);
and I_76(n54_10,n55_10,N1508_0_r_7);
nand I_77(n55_10,n56_10,n57_10);
nand I_78(n56_10,n_547_5_r_7,n_549_7_r_7);
not I_79(n57_10,n_429_or_0_5_r_7);
nor I_80(n58_10,n35_10,n45_10);
nor I_81(n59_10,n_576_5_r_7,G42_7_r_7);
nor I_82(n60_10,n37_10,n46_10);
or I_83(n61_10,n_576_5_r_7,G42_7_r_7);
nor I_84(n62_10,n_569_7_r_7,N1508_0_r_7);
or I_85(n63_10,n64_10,n_572_7_r_7);
nor I_86(n64_10,n_573_7_r_7,n_429_or_0_5_r_7);
endmodule


