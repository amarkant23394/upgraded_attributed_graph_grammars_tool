module test_final(G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_13,blif_reset_net_1_r_13,G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13);
input G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_13,blif_reset_net_1_r_13;
output G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13;
wire G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_569_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0,n4_1_l_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n_569_1_r_13,n4_1_l_13,n7_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13;
DFFARX1 I_0(n4_1_r_0,blif_clk_net_1_r_13,n7_13,G42_1_r_0,);
nor I_1(n_572_1_r_0,IN_5_1_l_0,n23_0);
nand I_2(n_573_1_r_0,n21_0,n22_0);
nand I_3(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_4(n_569_1_r_0,n21_0,n26_0);
nor I_5(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_6(N3_2_r_0,blif_clk_net_1_r_13,n7_13,G199_2_r_0,);
DFFARX1 I_7(N1_4_r_0,blif_clk_net_1_r_13,n7_13,G199_4_r_0,);
DFFARX1 I_8(n2_0,blif_clk_net_1_r_13,n7_13,G214_4_r_0,);
nor I_9(n4_1_l_0,G18_1_l_0,IN_1_1_l_0);
DFFARX1 I_10(n4_1_l_0,blif_clk_net_1_r_13,n7_13,n37_0,);
DFFARX1 I_11(IN_1_3_l_0,blif_clk_net_1_r_13,n7_13,n38_0,);
not I_12(n20_0,n38_0);
DFFARX1 I_13(IN_2_3_l_0,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_0,);
nor I_14(n4_1_r_0,IN_10_1_l_0,n23_0);
nor I_15(N3_2_r_0,n31_0,n32_0);
nor I_16(N1_4_r_0,n29_0,n32_0);
not I_17(n2_0,n31_0);
nor I_18(n21_0,IN_9_1_l_0,n37_0);
not I_19(n22_0,IN_5_1_l_0);
nand I_20(n23_0,n20_0,n30_0);
nand I_21(n24_0,n38_0,n25_0);
nor I_22(n25_0,IN_9_1_l_0,IN_10_1_l_0);
not I_23(n26_0,IN_10_1_l_0);
not I_24(n27_0,n29_0);
nor I_25(n28_0,G15_1_l_0,IN_7_1_l_0);
nand I_26(n29_0,n26_0,n33_0);
not I_27(n30_0,IN_9_1_l_0);
nand I_28(n31_0,IN_4_3_l_0,ACVQN1_3_l_0);
and I_29(n32_0,n35_0,n36_0);
nand I_30(n33_0,IN_4_1_l_0,n34_0);
not I_31(n34_0,G15_1_l_0);
nor I_32(n35_0,G18_1_l_0,G15_1_l_0);
nor I_33(n36_0,IN_5_1_l_0,IN_7_1_l_0);
DFFARX1 I_34(n4_1_r_13,blif_clk_net_1_r_13,n7_13,G42_1_r_13,);
nor I_35(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_36(n_573_1_r_13,n18_13,n19_13);
nand I_37(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_38(n_569_1_r_13,n17_13,n18_13);
nor I_39(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_40(n_266_and_0_3_l_13,blif_clk_net_1_r_13,n7_13,ACVQN2_3_r_13,);
nor I_41(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_42(n_549_1_l_13,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_13,);
not I_43(P6_5_r_13,P6_5_r_internal_13);
nor I_44(n4_1_l_13,G42_1_r_0,n_573_1_r_0);
not I_45(n7_13,blif_reset_net_1_r_13);
DFFARX1 I_46(n4_1_l_13,blif_clk_net_1_r_13,n7_13,n17_internal_13,);
not I_47(n17_13,n17_internal_13);
DFFARX1 I_48(n_573_1_r_0,blif_clk_net_1_r_13,n7_13,n28_13,);
DFFARX1 I_49(G199_2_r_0,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_13,);
nor I_50(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_51(n_266_and_0_3_l_13,ACVQN1_3_l_13,G42_1_r_0);
nand I_52(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_53(n_573_1_l_13,blif_clk_net_1_r_13,n7_13,n14_internal_13,);
not I_54(n14_13,n14_internal_13);
and I_55(n_549_1_l_13,n21_13,n26_13);
nand I_56(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_57(n_569_1_l_13,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_13,);
nand I_58(n18_13,n23_13,n24_13);
or I_59(n19_13,n_42_2_r_0,G199_4_r_0);
not I_60(n20_13,n_572_1_r_0);
not I_61(n21_13,n_572_1_r_0);
nand I_62(n22_13,n17_13,n28_13);
not I_63(n23_13,G42_1_r_0);
not I_64(n24_13,G214_4_r_0);
nor I_65(n25_13,n_42_2_r_0,G199_4_r_0);
nand I_66(n26_13,n27_13,n_549_1_r_0);
not I_67(n27_13,G199_4_r_0);
endmodule


