module test_I12208(I12140,I1477,I1470,I12208);
input I12140,I1477,I1470;
output I12208;
wire I10583,I10023,I10052,I10137,I10490,I11973,I12157,I10017,I12174,I7553,I12191,I10035;
DFFARX1 I_0(I10490,I1470,I10052,,,I10583,);
DFFARX1 I_1(I12191,I1470,I11973,,,I12208,);
DFFARX1 I_2(I10137,I1470,I10052,,,I10023,);
not I_3(I10052,I1477);
DFFARX1 I_4(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_5(I1470,I10052,,,I10490,);
not I_6(I11973,I1477);
nor I_7(I12157,I12140,I10035);
and I_8(I10017,I10490,I10583);
and I_9(I12174,I12157,I10017);
DFFARX1 I_10(I1470,,,I7553,);
or I_11(I12191,I12174,I10023);
not I_12(I10035,I10490);
endmodule


