module test_I7057(I5416,I3380,I1470,I5105,I7057);
input I5416,I3380,I1470,I5105;
output I7057;
wire I5070,I7026,I5249,I5481;
and I_0(I5070,I5249,I5481);
not I_1(I7026,I5070);
not I_2(I7057,I7026);
not I_3(I5249,I3380);
DFFARX1 I_4(I5416,I1470,I5105,,,I5481,);
endmodule


