module test_I3749(I2554,I1908,I1294,I1301,I3749);
input I2554,I1908,I1294,I1301;
output I3749;
wire I3622,I3396,I2668,I3379,I1914,I2651,I2548,I2702,I3246,I3715,I3732,I3698,I2572;
and I_0(I3749,I3622,I3732);
DFFARX1 I_1(I2572,I1294,I3246,,,I3622,);
not I_2(I3396,I3379);
nand I_3(I2668,I2651,I1914);
not I_4(I3379,I2548);
DFFARX1 I_5(I1294,,,I1914,);
nor I_6(I2651,I1908);
DFFARX1 I_7(I1294,,,I2548,);
not I_8(I2702,I1908);
not I_9(I3246,I1301);
not I_10(I3715,I3698);
nor I_11(I3732,I3715,I3396);
DFFARX1 I_12(I2554,I1294,I3246,,,I3698,);
nor I_13(I2572,I2668,I2702);
endmodule


