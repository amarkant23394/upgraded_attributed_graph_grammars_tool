module test_I14196(I1477,I13792,I12270,I11947,I1470,I14196);
input I1477,I13792,I12270,I11947,I1470;
output I14196;
wire I11935,I14004,I11941,I12208,I13987,I13775,I14179,I11950,I12239,I11938,I13809,I13826,I14162,I11973,I13970;
DFFARX1 I_0(I12208,I1470,I11973,,,I11935,);
DFFARX1 I_1(I13987,I1470,I13775,,,I14004,);
DFFARX1 I_2(I12208,I1470,I11973,,,I11941,);
DFFARX1 I_3(I1470,I11973,,,I12208,);
and I_4(I13987,I13970,I11941);
not I_5(I13775,I1477);
and I_6(I14196,I14004,I14179);
nand I_7(I14179,I14162,I13826);
DFFARX1 I_8(I1470,I11973,,,I11950,);
DFFARX1 I_9(I12208,I1470,I11973,,,I12239,);
and I_10(I11938,I12270,I12239);
and I_11(I13809,I13792,I11947);
DFFARX1 I_12(I13809,I1470,I13775,,,I13826,);
DFFARX1 I_13(I11938,I1470,I13775,,,I14162,);
not I_14(I11973,I1477);
nand I_15(I13970,I11935,I11950);
endmodule


