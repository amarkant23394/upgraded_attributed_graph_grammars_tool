module test_I2021(I1477,I1295,I1470,I2021);
input I1477,I1295,I1470;
output I2021;
wire I1518;
not I_0(I1518,I1477);
DFFARX1 I_1(I1295,I1470,I1518,,,I2021,);
endmodule


