module test_I6045(I4917,I4629,I1477,I4512,I4506,I1470,I6045);
input I4917,I4629,I1477,I4512,I4506,I1470;
output I6045;
wire I5994,I6028,I6011,I5751,I4521,I4527,I4544,I5932,I5915,I4595;
nand I_0(I5994,I4512,I4506);
nor I_1(I6045,I6028,I5932);
DFFARX1 I_2(I6011,I1470,I5751,,,I6028,);
and I_3(I6011,I5994,I4521);
not I_4(I5751,I1477);
DFFARX1 I_5(I4917,I1470,I4544,,,I4521,);
or I_6(I4527,I4629,I4595);
not I_7(I4544,I1477);
not I_8(I5932,I5915);
DFFARX1 I_9(I4527,I1470,I5751,,,I5915,);
DFFARX1 I_10(I1470,I4544,,,I4595,);
endmodule


