module Benchmark_testing85000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2507,I2514,I30115,I30106,I30103,I30109,I30097,I30091,I30112,I30100,I30094,I184764,I184740,I184752,I184746,I184761,I184755,I184749,I184743,I184758,I236529,I236505,I236517,I236511,I236526,I236520,I236514,I236508,I236523,I443626,I443605,I443599,I443614,I443602,I443617,I443608,I443611,I443623,I443620,I470282,I470261,I470255,I470270,I470258,I470273,I470264,I470267,I470279,I470276,I553284,I553281,I553272,I553275,I553269,I553278,I553266,I553290,I553287,I674083,I674086,I674068,I674077,I674089,I674080,I674071,I674074,I674092,I759049,I759052,I759034,I759043,I759055,I759046,I759037,I759040,I759058,I892114,I892117,I892093,I892105,I892120,I892108,I892102,I892096,I892099,I892111,I1110405,I1110393,I1110414,I1110390,I1110411,I1110402,I1110408,I1110399,I1110396,I1263448,I1263427,I1263433,I1263442,I1263445,I1263424,I1263439,I1263436,I1263430,I1281944,I1281923,I1281929,I1281938,I1281941,I1281920,I1281935,I1281932,I1281926,I1303684,I1303687,I1303672,I1303675,I1303669,I1303666,I1303690,I1303681,I1303663,I1303678);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2507,I2514;
output I30115,I30106,I30103,I30109,I30097,I30091,I30112,I30100,I30094,I184764,I184740,I184752,I184746,I184761,I184755,I184749,I184743,I184758,I236529,I236505,I236517,I236511,I236526,I236520,I236514,I236508,I236523,I443626,I443605,I443599,I443614,I443602,I443617,I443608,I443611,I443623,I443620,I470282,I470261,I470255,I470270,I470258,I470273,I470264,I470267,I470279,I470276,I553284,I553281,I553272,I553275,I553269,I553278,I553266,I553290,I553287,I674083,I674086,I674068,I674077,I674089,I674080,I674071,I674074,I674092,I759049,I759052,I759034,I759043,I759055,I759046,I759037,I759040,I759058,I892114,I892117,I892093,I892105,I892120,I892108,I892102,I892096,I892099,I892111,I1110405,I1110393,I1110414,I1110390,I1110411,I1110402,I1110408,I1110399,I1110396,I1263448,I1263427,I1263433,I1263442,I1263445,I1263424,I1263439,I1263436,I1263430,I1281944,I1281923,I1281929,I1281938,I1281941,I1281920,I1281935,I1281932,I1281926,I1303684,I1303687,I1303672,I1303675,I1303669,I1303666,I1303690,I1303681,I1303663,I1303678;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2507,I2514,I2546,I208543,I2572,I2580,I2597,I2538,I208549,I2637,I2645,I2662,I208558,I2679,I208552,I2696,I2713,I2517,I2744,I2761,I2778,I208555,I208561,I2520,I2809,I2826,I208564,I2843,I208540,I2860,I2877,I2894,I2529,I2925,I208546,I2942,I2959,I2535,I2990,I2532,I3021,I3047,I3055,I3072,I2526,I2523,I3141,I775242,I3167,I3175,I775221,I3192,I3133,I775230,I3232,I3240,I3257,I775236,I3274,I775233,I3291,I3308,I3112,I3339,I3356,I3373,I775224,I775218,I3115,I3404,I3421,I775239,I3438,I3455,I3472,I3489,I3124,I3520,I775227,I3537,I3554,I3130,I3585,I3127,I3616,I3642,I3650,I3667,I3121,I3118,I3736,I740562,I3762,I3770,I740541,I3787,I3728,I740550,I3827,I3835,I3852,I740556,I3869,I740553,I3886,I3903,I3707,I3934,I3951,I3968,I740544,I740538,I3710,I3999,I4016,I740559,I4033,I4050,I4067,I4084,I3719,I4115,I740547,I4132,I4149,I3725,I4180,I3722,I4211,I4237,I4245,I4262,I3716,I3713,I4331,I696634,I4357,I4365,I696613,I4382,I4323,I696622,I4422,I4430,I4447,I696628,I4464,I696625,I4481,I4498,I4302,I4529,I4546,I4563,I696616,I696610,I4305,I4594,I4611,I696631,I4628,I4645,I4662,I4679,I4314,I4710,I696619,I4727,I4744,I4320,I4775,I4317,I4806,I4832,I4840,I4857,I4311,I4308,I4926,I765416,I4952,I4960,I765395,I4977,I4918,I765404,I5017,I5025,I5042,I765410,I5059,I765407,I5076,I5093,I4897,I5124,I5141,I5158,I765398,I765392,I4900,I5189,I5206,I765413,I5223,I5240,I5257,I5274,I4909,I5305,I765401,I5322,I5339,I4915,I5370,I4912,I5401,I5427,I5435,I5452,I4906,I4903,I5521,I1043246,I5547,I5555,I1043258,I5572,I5513,I1043243,I5612,I5620,I5637,I5654,I1043240,I5671,I5688,I5492,I5719,I5736,I5753,I1043249,I5495,I5784,I5801,I1043255,I5818,I5835,I5852,I5869,I5504,I5900,I1043252,I5917,I5934,I5510,I5965,I5507,I5996,I1043261,I6022,I6030,I6047,I5501,I5498,I6116,I48548,I6142,I6150,I48539,I6167,I6108,I48560,I6207,I6215,I6232,I48536,I6249,I6266,I6283,I6087,I6314,I6331,I6348,I48545,I6090,I6379,I6396,I48557,I6413,I48554,I6430,I6447,I6464,I6099,I6495,I48551,I6512,I6529,I6105,I6560,I6102,I6591,I48542,I6617,I6625,I6642,I6096,I6093,I6711,I359294,I6737,I6745,I359285,I6762,I6703,I359288,I6802,I6810,I6827,I359282,I6844,I359291,I6861,I6878,I6682,I6909,I6926,I6943,I359279,I359297,I6685,I6974,I6991,I7008,I359303,I7025,I7042,I7059,I6694,I7090,I359300,I7107,I7124,I6700,I7155,I6697,I7186,I359306,I7212,I7220,I7237,I6691,I6688,I7306,I273393,I7332,I7340,I273384,I7357,I7298,I273387,I7397,I7405,I7422,I273381,I7439,I273390,I7456,I7473,I7277,I7504,I7521,I7538,I273378,I273396,I7280,I7569,I7586,I7603,I273402,I7620,I7637,I7654,I7289,I7685,I273399,I7702,I7719,I7295,I7750,I7292,I7781,I273405,I7807,I7815,I7832,I7286,I7283,I7901,I854430,I7927,I7935,I854421,I7952,I7893,I854427,I7992,I8000,I8017,I8034,I854433,I8051,I8068,I7872,I8099,I8116,I8133,I854442,I854439,I7875,I8164,I8181,I8198,I854424,I8215,I8232,I8249,I7884,I8280,I8297,I8314,I7890,I8345,I7887,I8376,I854436,I8402,I8410,I8427,I7881,I7878,I8496,I604133,I8522,I8530,I604151,I8547,I8488,I604145,I8587,I8595,I8612,I604136,I8629,I8646,I8663,I8467,I8694,I8711,I8728,I604142,I604130,I8470,I8759,I8776,I604148,I8793,I604154,I8810,I8827,I8844,I8479,I8875,I8892,I8909,I8485,I8940,I8482,I8971,I604139,I8997,I9005,I9022,I8476,I8473,I9091,I600665,I9117,I9125,I600683,I9142,I9083,I600677,I9182,I9190,I9207,I600668,I9224,I9241,I9258,I9062,I9289,I9306,I9323,I600674,I600662,I9065,I9354,I9371,I600680,I9388,I600686,I9405,I9422,I9439,I9074,I9470,I9487,I9504,I9080,I9535,I9077,I9566,I600671,I9592,I9600,I9617,I9071,I9068,I9686,I624363,I9712,I9720,I624381,I9737,I9678,I624375,I9777,I9785,I9802,I624366,I9819,I9836,I9853,I9657,I9884,I9901,I9918,I624372,I624360,I9660,I9949,I9966,I624378,I9983,I624384,I10000,I10017,I10034,I9669,I10065,I10082,I10099,I9675,I10130,I9672,I10161,I624369,I10187,I10195,I10212,I9666,I9663,I10281,I60669,I10307,I10315,I60660,I10332,I10273,I60681,I10372,I10380,I10397,I60657,I10414,I10431,I10448,I10252,I10479,I10496,I10513,I60666,I10255,I10544,I10561,I60678,I10578,I60675,I10595,I10612,I10629,I10264,I10660,I60672,I10677,I10694,I10270,I10725,I10267,I10756,I60663,I10782,I10790,I10807,I10261,I10258,I10876,I904388,I10902,I10910,I904379,I10927,I10868,I904382,I10967,I10975,I10992,I904394,I11009,I904373,I11026,I11043,I10847,I11074,I11091,I11108,I904385,I904391,I10850,I11139,I11156,I904376,I11173,I904367,I11190,I11207,I11224,I10859,I11255,I11272,I11289,I10865,I11320,I10862,I11351,I904370,I11377,I11385,I11402,I10856,I10853,I11471,I383780,I11497,I11505,I383762,I11522,I11463,I383774,I11562,I11570,I11587,I383759,I11604,I383768,I11621,I11638,I11442,I11669,I11686,I11703,I383765,I383786,I11445,I11734,I11751,I383777,I11768,I383783,I11785,I11802,I11819,I11454,I11850,I11867,I11884,I11460,I11915,I11457,I11946,I383771,I11972,I11980,I11997,I11451,I11448,I12066,I12092,I12100,I12117,I12058,I12157,I12165,I12182,I12199,I12216,I12233,I12037,I12264,I12281,I12298,I12040,I12329,I12346,I12363,I12380,I12397,I12414,I12049,I12445,I12462,I12479,I12055,I12510,I12052,I12541,I12567,I12575,I12592,I12046,I12043,I12661,I903096,I12687,I12695,I903087,I12712,I12653,I903090,I12752,I12760,I12777,I903102,I12794,I903081,I12811,I12828,I12632,I12859,I12876,I12893,I903093,I903099,I12635,I12924,I12941,I903084,I12958,I903075,I12975,I12992,I13009,I12644,I13040,I13057,I13074,I12650,I13105,I12647,I13136,I903078,I13162,I13170,I13187,I12641,I12638,I13259,I224016,I13285,I13302,I13310,I13327,I224034,I224019,I13344,I224022,I13370,I13251,I13242,I224010,I13415,I13423,I224013,I13440,I13239,I224025,I13480,I13488,I13245,I13233,I13533,I224031,I224028,I13550,I13576,I13584,I13227,I13615,I13632,I13649,I13666,I13683,I13248,I13714,I13236,I13230,I13786,I1039880,I13812,I13829,I13837,I13854,I1039874,I1039895,I13871,I13897,I13778,I13769,I1039877,I13942,I13950,I1039886,I13967,I13766,I14007,I14015,I13772,I13760,I14060,I1039892,I14077,I1039883,I14103,I14111,I13754,I14142,I14159,I1039889,I14176,I14193,I14210,I13775,I14241,I13763,I13757,I14313,I859700,I14339,I14356,I14364,I14381,I859691,I859712,I14398,I859694,I14424,I14305,I14296,I14469,I14477,I859709,I14494,I14293,I859703,I14534,I14542,I14299,I14287,I14587,I859697,I859706,I14604,I14630,I14638,I14281,I14669,I14686,I14703,I14720,I14737,I14302,I14768,I14290,I14284,I14840,I53282,I14866,I14883,I14891,I14908,I53297,I14925,I53300,I14951,I14832,I14823,I53294,I14996,I15004,I53303,I15021,I14820,I53279,I15061,I15069,I14826,I14814,I15114,I53285,I15131,I53288,I15157,I15165,I14808,I15196,I15213,I53291,I15230,I15247,I15264,I14829,I15295,I14817,I14811,I15367,I1136424,I15393,I15410,I15418,I15435,I1136412,I1136403,I15452,I1136400,I15478,I15359,I15350,I1136406,I15523,I15531,I1136418,I15548,I15347,I1136415,I15588,I15596,I15353,I15341,I15641,I1136409,I15658,I1136421,I15684,I15692,I15335,I15723,I15740,I15757,I15774,I15791,I15356,I15822,I15344,I15338,I15894,I205571,I15920,I15937,I15945,I15962,I205589,I205574,I15979,I205577,I16005,I15886,I15877,I205565,I16050,I16058,I205568,I16075,I15874,I205580,I16115,I16123,I15880,I15868,I16168,I205586,I205583,I16185,I16211,I16219,I15862,I16250,I16267,I16284,I16301,I16318,I15883,I16349,I15871,I15865,I16421,I649220,I16447,I16464,I16472,I16489,I649235,I649238,I16506,I649217,I16532,I16413,I16404,I649223,I16577,I16585,I649229,I16602,I16401,I16642,I16650,I16407,I16395,I16695,I649232,I649214,I16712,I649226,I16738,I16746,I16389,I16777,I16794,I16811,I16828,I16845,I16410,I16876,I16398,I16392,I16948,I818594,I16974,I16991,I16999,I17016,I818585,I818606,I17033,I818588,I17059,I16940,I16931,I17104,I17112,I818603,I17129,I16928,I818597,I17169,I17177,I16934,I16922,I17222,I818591,I818600,I17239,I17265,I17273,I16916,I17304,I17321,I17338,I17355,I17372,I16937,I17403,I16925,I16919,I17475,I853903,I17501,I17518,I17526,I17543,I853894,I853915,I17560,I853897,I17586,I17467,I17458,I17631,I17639,I853912,I17656,I17455,I853906,I17696,I17704,I17461,I17449,I17749,I853900,I853909,I17766,I17792,I17800,I17443,I17831,I17848,I17865,I17882,I17899,I17464,I17930,I17452,I17446,I18002,I375643,I18028,I18045,I18053,I18070,I375640,I375634,I18087,I375628,I18113,I17994,I17985,I375616,I18158,I18166,I375625,I18183,I17982,I375622,I18223,I18231,I17988,I17976,I18276,I375619,I375637,I18293,I18319,I18327,I17970,I18358,I18375,I375631,I18392,I18409,I18426,I17991,I18457,I17979,I17973,I18529,I493103,I18555,I18572,I18580,I18597,I493106,I18614,I493127,I18640,I18521,I18512,I493115,I18685,I18693,I493118,I18710,I18509,I493124,I18750,I18758,I18515,I18503,I18803,I493121,I493109,I18820,I493112,I18846,I18854,I18497,I18885,I18902,I493130,I18919,I18936,I18953,I18518,I18984,I18506,I18500,I19056,I252325,I19082,I19099,I19107,I19124,I252322,I252316,I19141,I252310,I19167,I19048,I19039,I252298,I19212,I19220,I252307,I19237,I19036,I252304,I19277,I19285,I19042,I19030,I19330,I252301,I252319,I19347,I19373,I19381,I19024,I19412,I19429,I252313,I19446,I19463,I19480,I19045,I19511,I19033,I19027,I19583,I351928,I19609,I19626,I19634,I19651,I351925,I351919,I19668,I351913,I19694,I19575,I19566,I351901,I19739,I19747,I351910,I19764,I19563,I351907,I19804,I19812,I19569,I19557,I19857,I351904,I351922,I19874,I19900,I19908,I19551,I19939,I19956,I351916,I19973,I19990,I20007,I19572,I20038,I19560,I19554,I20110,I354563,I20136,I20153,I20161,I20178,I354560,I354554,I20195,I354548,I20221,I20102,I20093,I354536,I20266,I20274,I354545,I20291,I20090,I354542,I20331,I20339,I20096,I20084,I20384,I354539,I354557,I20401,I20427,I20435,I20078,I20466,I20483,I354551,I20500,I20517,I20534,I20099,I20565,I20087,I20081,I20637,I90172,I20663,I20680,I20688,I20705,I90187,I20722,I90190,I20748,I20629,I20620,I90184,I20793,I20801,I90193,I20818,I20617,I90169,I20858,I20866,I20623,I20611,I20911,I90175,I20928,I90178,I20954,I20962,I20605,I20993,I21010,I90181,I21027,I21044,I21061,I20626,I21092,I20614,I20608,I21164,I1300882,I21190,I21207,I21215,I21232,I1300873,I1300879,I21249,I1300858,I21275,I21156,I21147,I1300876,I21320,I21328,I21345,I21144,I1300870,I21385,I21393,I21150,I21138,I21438,I1300864,I1300885,I21455,I1300867,I21481,I21489,I21132,I21520,I21537,I1300861,I21554,I21571,I21588,I21153,I21619,I21141,I21135,I21691,I671184,I21717,I21734,I21742,I21759,I671199,I671202,I21776,I671181,I21802,I21683,I21674,I671187,I21847,I21855,I671193,I21872,I21671,I21912,I21920,I21677,I21665,I21965,I671196,I671178,I21982,I671190,I22008,I22016,I21659,I22047,I22064,I22081,I22098,I22115,I21680,I22146,I21668,I21662,I22218,I749214,I22244,I22261,I22269,I22286,I749229,I749232,I22303,I749211,I22329,I22210,I22201,I749217,I22374,I22382,I749223,I22399,I22198,I22439,I22447,I22204,I22192,I22492,I749226,I749208,I22509,I749220,I22535,I22543,I22186,I22574,I22591,I22608,I22625,I22642,I22207,I22673,I22195,I22189,I22745,I1157810,I22771,I22788,I22796,I22813,I1157798,I1157789,I22830,I1157786,I22856,I22737,I22728,I1157792,I22901,I22909,I1157804,I22926,I22725,I1157801,I22966,I22974,I22731,I22719,I23019,I1157795,I23036,I1157807,I23062,I23070,I22713,I23101,I23118,I23135,I23152,I23169,I22734,I23200,I22722,I22716,I23272,I771178,I23298,I23315,I23323,I23340,I771193,I771196,I23357,I771175,I23383,I23264,I23255,I771181,I23428,I23436,I771187,I23453,I23252,I23493,I23501,I23258,I23246,I23546,I771190,I771172,I23563,I771184,I23589,I23597,I23240,I23628,I23645,I23662,I23679,I23696,I23261,I23727,I23249,I23243,I23799,I444143,I23825,I23842,I23850,I23867,I444146,I23884,I444167,I23910,I23791,I23782,I444155,I23955,I23963,I444158,I23980,I23779,I444164,I24020,I24028,I23785,I23773,I24073,I444161,I444149,I24090,I444152,I24116,I24124,I23767,I24155,I24172,I444170,I24189,I24206,I24223,I23788,I24254,I23776,I23770,I24326,I610503,I24352,I24369,I24377,I24394,I610488,I610506,I24411,I610500,I24437,I24318,I24309,I610497,I24482,I24490,I24507,I24306,I610491,I24547,I24555,I24312,I24300,I24600,I610512,I610494,I24617,I610509,I24643,I24651,I24294,I24682,I24699,I24716,I24733,I24750,I24315,I24781,I24303,I24297,I24853,I1109836,I24879,I24896,I24904,I24921,I1109824,I1109815,I24938,I1109812,I24964,I24845,I24836,I1109818,I25009,I25017,I1109830,I25034,I24833,I1109827,I25074,I25082,I24839,I24827,I25127,I1109821,I25144,I1109833,I25170,I25178,I24821,I25209,I25226,I25243,I25260,I25277,I24842,I25308,I24830,I24824,I25380,I113360,I25406,I25423,I25431,I25448,I113375,I25465,I113378,I25491,I25372,I25363,I113372,I25536,I25544,I113381,I25561,I25360,I113357,I25601,I25609,I25366,I25354,I25654,I113363,I25671,I113366,I25697,I25705,I25348,I25736,I25753,I113369,I25770,I25787,I25804,I25369,I25835,I25357,I25351,I25907,I972867,I25933,I25950,I25958,I25975,I972843,I972870,I25992,I972855,I26018,I25899,I25890,I972861,I26063,I26071,I972846,I26088,I25887,I972864,I26128,I26136,I25893,I25881,I26181,I972849,I972852,I26198,I26224,I26232,I25875,I26263,I26280,I972858,I26297,I26314,I26331,I25896,I26362,I25884,I25878,I26434,I143105,I26460,I26477,I26485,I26502,I143108,I143090,I26519,I143096,I26545,I26426,I26417,I143099,I26590,I26598,I26615,I26414,I143111,I26655,I26663,I26420,I26408,I26708,I143114,I143102,I26725,I143093,I26751,I26759,I26402,I26790,I26807,I143117,I26824,I26841,I26858,I26423,I26889,I26411,I26405,I26961,I728984,I26987,I27004,I27012,I27029,I728999,I729002,I27046,I728981,I27072,I26953,I26944,I728987,I27117,I27125,I728993,I27142,I26941,I27182,I27190,I26947,I26935,I27235,I728996,I728978,I27252,I728990,I27278,I27286,I26929,I27317,I27334,I27351,I27368,I27385,I26950,I27416,I26938,I26932,I27488,I336645,I27514,I27531,I27539,I27556,I336642,I336636,I27573,I336630,I27599,I27480,I27471,I336618,I27644,I27652,I336627,I27669,I27468,I336624,I27709,I27717,I27474,I27462,I27762,I336621,I336639,I27779,I27805,I27813,I27456,I27844,I27861,I336633,I27878,I27895,I27912,I27477,I27943,I27465,I27459,I28015,I557327,I28041,I28058,I28066,I28083,I557312,I557330,I28100,I557324,I28126,I28007,I27998,I557321,I28171,I28179,I28196,I27995,I557315,I28236,I28244,I28001,I27989,I28289,I557336,I557318,I28306,I557333,I28332,I28340,I27983,I28371,I28388,I28405,I28422,I28439,I28004,I28470,I27992,I27986,I28542,I1024172,I28568,I28585,I28593,I28610,I1024166,I1024187,I28627,I28653,I28534,I28525,I1024169,I28698,I28706,I1024178,I28723,I28522,I28763,I28771,I28528,I28516,I28816,I1024184,I28833,I1024175,I28859,I28867,I28510,I28898,I28915,I1024181,I28932,I28949,I28966,I28531,I28997,I28519,I28513,I29069,I804892,I29095,I29112,I29120,I29137,I804883,I804904,I29154,I804886,I29180,I29061,I29052,I29225,I29233,I804901,I29250,I29049,I804895,I29290,I29298,I29055,I29043,I29343,I804889,I804898,I29360,I29386,I29394,I29037,I29425,I29442,I29459,I29476,I29493,I29058,I29524,I29046,I29040,I29596,I1119662,I29622,I29639,I29647,I29664,I1119650,I1119641,I29681,I1119638,I29707,I29588,I29579,I1119644,I29752,I29760,I1119656,I29777,I29576,I1119653,I29817,I29825,I29582,I29570,I29870,I1119647,I29887,I1119659,I29913,I29921,I29564,I29952,I29969,I29986,I30003,I30020,I29585,I30051,I29573,I29567,I30123,I724938,I30149,I30166,I30174,I30191,I724953,I724956,I30208,I724935,I30234,I724941,I30279,I30287,I724947,I30304,I30344,I30352,I30397,I724950,I724932,I30414,I724944,I30440,I30448,I30479,I30496,I30513,I30530,I30547,I30578,I30650,I395183,I30676,I30693,I30701,I30718,I395186,I30735,I395207,I30761,I30642,I30633,I395195,I30806,I30814,I395198,I30831,I30630,I395204,I30871,I30879,I30636,I30624,I30924,I395201,I395189,I30941,I395192,I30967,I30975,I30618,I31006,I31023,I395210,I31040,I31057,I31074,I30639,I31105,I30627,I30621,I31177,I561951,I31203,I31220,I31228,I31245,I561936,I561954,I31262,I561948,I31288,I31169,I31160,I561945,I31333,I31341,I31358,I31157,I561939,I31398,I31406,I31163,I31151,I31451,I561960,I561942,I31468,I561957,I31494,I31502,I31145,I31533,I31550,I31567,I31584,I31601,I31166,I31632,I31154,I31148,I31704,I1132378,I31730,I31747,I31755,I31772,I1132366,I1132357,I31789,I1132354,I31815,I31696,I31687,I1132360,I31860,I31868,I1132372,I31885,I31684,I1132369,I31925,I31933,I31690,I31678,I31978,I1132363,I31995,I1132375,I32021,I32029,I31672,I32060,I32077,I32094,I32111,I32128,I31693,I32159,I31681,I31675,I32231,I725516,I32257,I32274,I32282,I32299,I725531,I725534,I32316,I725513,I32342,I32223,I32214,I725519,I32387,I32395,I725525,I32412,I32211,I32452,I32460,I32217,I32205,I32505,I725528,I725510,I32522,I725522,I32548,I32556,I32199,I32587,I32604,I32621,I32638,I32655,I32220,I32686,I32208,I32202,I32758,I302390,I32784,I32801,I32809,I32826,I302387,I302381,I32843,I302375,I32869,I32750,I32741,I302363,I32914,I32922,I302372,I32939,I32738,I302369,I32979,I32987,I32744,I32732,I33032,I302366,I302384,I33049,I33075,I33083,I32726,I33114,I33131,I302378,I33148,I33165,I33182,I32747,I33213,I32735,I32729,I33285,I315565,I33311,I33328,I33336,I33353,I315562,I315556,I33370,I315550,I33396,I33277,I33268,I315538,I33441,I33449,I315547,I33466,I33265,I315544,I33506,I33514,I33271,I33259,I33559,I315541,I315559,I33576,I33602,I33610,I33253,I33641,I33658,I315553,I33675,I33692,I33709,I33274,I33740,I33262,I33256,I33812,I1280779,I33838,I33855,I33863,I33880,I1280782,I1280776,I33897,I1280785,I33923,I33804,I33795,I1280773,I33968,I33976,I1280788,I33993,I33792,I1280764,I34033,I34041,I33798,I33786,I34086,I1280767,I34103,I34129,I34137,I33780,I34168,I34185,I1280770,I34202,I34219,I34236,I33801,I34267,I33789,I33783,I34339,I1264595,I34365,I34382,I34390,I34407,I1264598,I1264592,I34424,I1264601,I34450,I34331,I34322,I1264589,I34495,I34503,I1264604,I34520,I34319,I1264580,I34560,I34568,I34325,I34313,I34613,I1264583,I34630,I34656,I34664,I34307,I34695,I34712,I1264586,I34729,I34746,I34763,I34328,I34794,I34316,I34310,I34866,I1026977,I34892,I34909,I34917,I34934,I1026971,I1026992,I34951,I34977,I34858,I34849,I1026974,I35022,I35030,I1026983,I35047,I34846,I35087,I35095,I34852,I34840,I35140,I1026989,I35157,I1026980,I35183,I35191,I34834,I35222,I35239,I1026986,I35256,I35273,I35290,I34855,I35321,I34843,I34837,I35393,I897285,I35419,I35436,I35444,I35461,I897261,I897288,I35478,I897273,I35504,I35385,I35376,I897279,I35549,I35557,I897264,I35574,I35373,I897282,I35614,I35622,I35379,I35367,I35667,I897267,I897270,I35684,I35710,I35718,I35361,I35749,I35766,I897276,I35783,I35800,I35817,I35382,I35848,I35370,I35364,I35920,I901807,I35946,I35963,I35971,I35988,I901783,I901810,I36005,I901795,I36031,I35912,I35903,I901801,I36076,I36084,I901786,I36101,I35900,I901804,I36141,I36149,I35906,I35894,I36194,I901789,I901792,I36211,I36237,I36245,I35888,I36276,I36293,I901798,I36310,I36327,I36344,I35909,I36375,I35897,I35891,I36447,I866024,I36473,I36490,I36498,I36515,I866015,I866036,I36532,I866018,I36558,I36439,I36430,I36603,I36611,I866033,I36628,I36427,I866027,I36668,I36676,I36433,I36421,I36721,I866021,I866030,I36738,I36764,I36772,I36415,I36803,I36820,I36837,I36854,I36871,I36436,I36902,I36424,I36418,I36974,I1299199,I37000,I37017,I37025,I37042,I1299190,I1299196,I37059,I1299175,I37085,I36966,I36957,I1299193,I37130,I37138,I37155,I36954,I1299187,I37195,I37203,I36960,I36948,I37248,I1299181,I1299202,I37265,I1299184,I37291,I37299,I36942,I37330,I37347,I1299178,I37364,I37381,I37398,I36963,I37429,I36951,I36945,I37501,I689680,I37527,I37544,I37552,I37569,I689695,I689698,I37586,I689677,I37612,I37493,I37484,I689683,I37657,I37665,I689689,I37682,I37481,I37722,I37730,I37487,I37475,I37775,I689692,I689674,I37792,I689686,I37818,I37826,I37469,I37857,I37874,I37891,I37908,I37925,I37490,I37956,I37478,I37472,I38028,I503023,I38054,I38071,I38079,I38096,I503029,I503017,I38113,I503014,I38139,I38020,I38011,I503026,I38184,I38192,I503020,I38209,I38008,I503038,I38249,I38257,I38014,I38002,I38302,I503032,I503035,I38319,I38345,I38353,I37996,I38384,I38401,I38418,I38435,I38452,I38017,I38483,I38005,I37999,I38555,I273932,I38581,I38598,I38606,I38623,I273929,I273923,I38640,I273917,I38666,I38547,I38538,I273905,I38711,I38719,I273914,I38736,I38535,I273911,I38776,I38784,I38541,I38529,I38829,I273908,I273926,I38846,I38872,I38880,I38523,I38911,I38928,I273920,I38945,I38962,I38979,I38544,I39010,I38532,I38526,I39082,I148451,I39108,I39125,I39133,I39150,I148469,I148454,I39167,I148457,I39193,I39074,I39065,I148445,I39238,I39246,I148448,I39263,I39062,I148460,I39303,I39311,I39068,I39056,I39356,I148466,I148463,I39373,I39399,I39407,I39050,I39438,I39455,I39472,I39489,I39506,I39071,I39537,I39059,I39053,I39609,I1130644,I39635,I39652,I39660,I39677,I1130632,I1130623,I39694,I1130620,I39720,I39601,I39592,I1130626,I39765,I39773,I1130638,I39790,I39589,I1130635,I39830,I39838,I39595,I39583,I39883,I1130629,I39900,I1130641,I39926,I39934,I39577,I39965,I39982,I39999,I40016,I40033,I39598,I40064,I39586,I39580,I40136,I514328,I40162,I40179,I40187,I40204,I514334,I514322,I40221,I514319,I40247,I40128,I40119,I514331,I40292,I40300,I514325,I40317,I40116,I514343,I40357,I40365,I40122,I40110,I40410,I514337,I514340,I40427,I40453,I40461,I40104,I40492,I40509,I40526,I40543,I40560,I40125,I40591,I40113,I40107,I40663,I49593,I40689,I40706,I40714,I40731,I49608,I40748,I49611,I40774,I40655,I40646,I49605,I40819,I40827,I49614,I40844,I40643,I49590,I40884,I40892,I40649,I40637,I40937,I49596,I40954,I49599,I40980,I40988,I40631,I41019,I41036,I49602,I41053,I41070,I41087,I40652,I41118,I40640,I40634,I41190,I1132956,I41216,I41233,I41241,I41258,I1132944,I1132935,I41275,I1132932,I41301,I41182,I41173,I1132938,I41346,I41354,I1132950,I41371,I41170,I1132947,I41411,I41419,I41176,I41164,I41464,I1132941,I41481,I1132953,I41507,I41515,I41158,I41546,I41563,I41580,I41597,I41614,I41179,I41645,I41167,I41161,I41717,I757306,I41743,I41760,I41768,I41785,I757321,I757324,I41802,I757303,I41828,I41709,I41700,I757309,I41873,I41881,I757315,I41898,I41697,I41938,I41946,I41703,I41691,I41991,I757318,I757300,I42008,I757312,I42034,I42042,I41685,I42073,I42090,I42107,I42124,I42141,I41706,I42172,I41694,I41688,I42244,I168086,I42270,I42287,I42295,I42312,I168104,I168089,I42329,I168092,I42355,I42236,I42227,I168080,I42400,I42408,I168083,I42425,I42224,I168095,I42465,I42473,I42230,I42218,I42518,I168101,I168098,I42535,I42561,I42569,I42212,I42600,I42617,I42634,I42651,I42668,I42233,I42699,I42221,I42215,I42771,I295012,I42797,I42814,I42822,I42839,I295009,I295003,I42856,I294997,I42882,I42763,I42754,I294985,I42927,I42935,I294994,I42952,I42751,I294991,I42992,I43000,I42757,I42745,I43045,I294988,I295006,I43062,I43088,I43096,I42739,I43127,I43144,I295000,I43161,I43178,I43195,I42760,I43226,I42748,I42742,I43298,I564841,I43324,I43341,I43349,I43366,I564826,I564844,I43383,I564838,I43409,I43290,I43281,I564835,I43454,I43462,I43479,I43278,I564829,I43519,I43527,I43284,I43272,I43572,I564850,I564832,I43589,I564847,I43615,I43623,I43266,I43654,I43671,I43688,I43705,I43722,I43287,I43753,I43275,I43269,I43825,I1131800,I43851,I43868,I43876,I43893,I1131788,I1131779,I43910,I1131776,I43936,I43817,I43808,I1131782,I43981,I43989,I1131794,I44006,I43805,I1131791,I44046,I44054,I43811,I43799,I44099,I1131785,I44116,I1131797,I44142,I44150,I43793,I44181,I44198,I44215,I44232,I44249,I43814,I44280,I43802,I43796,I44352,I679854,I44378,I44395,I44403,I44420,I679869,I679872,I44437,I679851,I44463,I44344,I44335,I679857,I44508,I44516,I679863,I44533,I44332,I44573,I44581,I44338,I44326,I44626,I679866,I679848,I44643,I679860,I44669,I44677,I44320,I44708,I44725,I44742,I44759,I44776,I44341,I44807,I44329,I44323,I44879,I1013513,I44905,I44922,I44930,I44947,I1013507,I1013528,I44964,I44990,I44871,I44862,I1013510,I45035,I45043,I1013519,I45060,I44859,I45100,I45108,I44865,I44853,I45153,I1013525,I45170,I1013516,I45196,I45204,I44847,I45235,I45252,I1013522,I45269,I45286,I45303,I44868,I45334,I44856,I44850,I45406,I655000,I45432,I45449,I45457,I45474,I655015,I655018,I45491,I654997,I45517,I45398,I45389,I655003,I45562,I45570,I655009,I45587,I45386,I45627,I45635,I45392,I45380,I45680,I655012,I654994,I45697,I655006,I45723,I45731,I45374,I45762,I45779,I45796,I45813,I45830,I45395,I45861,I45383,I45377,I45933,I565997,I45959,I45976,I45984,I46001,I565982,I566000,I46018,I565994,I46044,I45925,I45916,I565991,I46089,I46097,I46114,I45913,I565985,I46154,I46162,I45919,I45907,I46207,I566006,I565988,I46224,I566003,I46250,I46258,I45901,I46289,I46306,I46323,I46340,I46357,I45922,I46388,I45910,I45904,I46460,I415855,I46486,I46503,I46511,I46528,I415858,I46545,I415879,I46571,I46452,I46443,I415867,I46616,I46624,I415870,I46641,I46440,I415876,I46681,I46689,I46446,I46434,I46734,I415873,I415861,I46751,I415864,I46777,I46785,I46428,I46816,I46833,I415882,I46850,I46867,I46884,I46449,I46915,I46437,I46431,I46987,I1076890,I47013,I47030,I47038,I47055,I1076878,I1076869,I47072,I1076866,I47098,I46979,I46970,I1076872,I47143,I47151,I1076884,I47168,I46967,I1076881,I47208,I47216,I46973,I46961,I47261,I1076875,I47278,I1076887,I47304,I47312,I46955,I47343,I47360,I47377,I47394,I47411,I46976,I47442,I46964,I46958,I47514,I140130,I47540,I47557,I47565,I47582,I140133,I140115,I47599,I140121,I47625,I47506,I47497,I140124,I47670,I47678,I47695,I47494,I140136,I47735,I47743,I47500,I47488,I47788,I140139,I140127,I47805,I140118,I47831,I47839,I47482,I47870,I47887,I140142,I47904,I47921,I47938,I47503,I47969,I47491,I47485,I48041,I943151,I48067,I48084,I48092,I48109,I943127,I943154,I48126,I943139,I48152,I48033,I48024,I943145,I48197,I48205,I943130,I48222,I48021,I943148,I48262,I48270,I48027,I48015,I48315,I943133,I943136,I48332,I48358,I48366,I48009,I48397,I48414,I943142,I48431,I48448,I48465,I48030,I48496,I48018,I48012,I48568,I611653,I48594,I48602,I48619,I611665,I611650,I48636,I611644,I48662,I611659,I48679,I48687,I611647,I48704,I48735,I48752,I611656,I48792,I48814,I611662,I611668,I48831,I48857,I48874,I48896,I48927,I48944,I48961,I48978,I49009,I49095,I757890,I49121,I49129,I49146,I757881,I757899,I49163,I757878,I49189,I49206,I49214,I757884,I49231,I49063,I49262,I49279,I49075,I49319,I49084,I49341,I757896,I757887,I49358,I757902,I49384,I49401,I49087,I49423,I49072,I49454,I757893,I49471,I49488,I49505,I49081,I49536,I49069,I49078,I49066,I49622,I1138718,I49648,I49656,I49673,I1138733,I1138712,I49690,I1138715,I49716,I1138736,I49733,I49741,I49758,I49789,I49806,I49846,I49868,I1138724,I1138721,I49885,I1138727,I49911,I49928,I49950,I49981,I1138730,I49998,I50015,I50032,I50063,I50149,I306079,I50175,I50183,I50200,I306061,I306076,I50217,I306052,I50243,I306055,I50260,I50268,I306070,I50285,I50117,I50316,I50333,I50129,I306073,I50373,I50138,I50395,I306064,I50412,I306058,I50438,I50455,I50141,I50477,I50126,I50508,I306067,I50525,I50542,I50559,I50135,I50590,I50123,I50132,I50120,I50676,I1286565,I50702,I50710,I50727,I1286568,I1286562,I50744,I1286559,I50770,I1286544,I50787,I50795,I1286553,I50812,I50644,I50843,I50860,I50656,I50900,I50665,I50922,I1286547,I1286550,I50939,I1286556,I50965,I50982,I50668,I51004,I50653,I51035,I51052,I51069,I51086,I50662,I51117,I50650,I50659,I50647,I51203,I1141030,I51229,I51237,I51254,I1141045,I1141024,I51271,I1141027,I51297,I1141048,I51314,I51322,I51339,I51171,I51370,I51387,I51183,I51427,I51192,I51449,I1141036,I1141033,I51466,I1141039,I51492,I51509,I51195,I51531,I51180,I51562,I1141042,I51579,I51596,I51613,I51189,I51644,I51177,I51186,I51174,I51730,I1118488,I51756,I51764,I51781,I1118503,I1118482,I51798,I1118485,I51824,I1118506,I51841,I51849,I51866,I51698,I51897,I51914,I51710,I51954,I51719,I51976,I1118494,I1118491,I51993,I1118497,I52019,I52036,I51722,I52058,I51707,I52089,I1118500,I52106,I52123,I52140,I51716,I52171,I51704,I51713,I51701,I52257,I991586,I52283,I52291,I52308,I991604,I991598,I52325,I991577,I52351,I991595,I52368,I52376,I991580,I52393,I52225,I52424,I52441,I52237,I991592,I52481,I52246,I52503,I991601,I991589,I52520,I991583,I52546,I52563,I52249,I52585,I52234,I52616,I52633,I52650,I52667,I52243,I52698,I52231,I52240,I52228,I52784,I1327934,I52810,I52818,I52835,I1327928,I1327949,I52852,I1327925,I52878,I1327946,I52895,I52903,I1327943,I52920,I52752,I52951,I52968,I52764,I1327931,I53008,I52773,I53030,I1327940,I1327937,I53047,I1327922,I53073,I53090,I52776,I53112,I52761,I53143,I53160,I53177,I53194,I52770,I53225,I52758,I52767,I52755,I53311,I53337,I53345,I53362,I53379,I53405,I53422,I53430,I53447,I53478,I53495,I53535,I53557,I53574,I53600,I53617,I53639,I53670,I53687,I53704,I53721,I53752,I53838,I1030901,I53864,I53872,I53889,I1030898,I1030904,I53906,I53932,I53949,I53957,I53974,I53806,I54005,I54022,I53818,I1030907,I54062,I53827,I54084,I1030910,I1030919,I54101,I1030913,I54127,I54144,I53830,I54166,I53815,I54197,I1030916,I54214,I54231,I54248,I53824,I54279,I53812,I53821,I53809,I54365,I669456,I54391,I54399,I54416,I669447,I669465,I54433,I669444,I54459,I54476,I54484,I669450,I54501,I54333,I54532,I54549,I54345,I54589,I54354,I54611,I669462,I669453,I54628,I669468,I54654,I54671,I54357,I54693,I54342,I54724,I669459,I54741,I54758,I54775,I54351,I54806,I54339,I54348,I54336,I54892,I883942,I54918,I54926,I54943,I883939,I883954,I54960,I883936,I54986,I883933,I55003,I55011,I55028,I54860,I55059,I55076,I54872,I55116,I54881,I55138,I883948,I55155,I883951,I55181,I55198,I54884,I55220,I54869,I55251,I883945,I55268,I55285,I55302,I54878,I55333,I54866,I54875,I54863,I55419,I536337,I55445,I55453,I55470,I536358,I536352,I55487,I536334,I55513,I55530,I55538,I536346,I55555,I55387,I55586,I55603,I55399,I536343,I55643,I55408,I55665,I536349,I536340,I55682,I55708,I55725,I55411,I55747,I55396,I55778,I536355,I55795,I55812,I55829,I55405,I55860,I55393,I55402,I55390,I55946,I219262,I55972,I55980,I55997,I219256,I219250,I56014,I219271,I56040,I219268,I56057,I56065,I219265,I56082,I55914,I56113,I56130,I55926,I56170,I55935,I56192,I219253,I56209,I219274,I56235,I56252,I55938,I56274,I55923,I56305,I219259,I56322,I56339,I56356,I55932,I56387,I55920,I55929,I55917,I56473,I819121,I56499,I56507,I56524,I819118,I819133,I56541,I819115,I56567,I819112,I56584,I56592,I56609,I56441,I56640,I56657,I56453,I56697,I56462,I56719,I819127,I56736,I819130,I56762,I56779,I56465,I56801,I56450,I56832,I819124,I56849,I56866,I56883,I56459,I56914,I56447,I56456,I56444,I57000,I713384,I57026,I57034,I57051,I713375,I713393,I57068,I713372,I57094,I57111,I57119,I713378,I57136,I56968,I57167,I57184,I56980,I57224,I56989,I57246,I713390,I713381,I57263,I713396,I57289,I57306,I56992,I57328,I56977,I57359,I713387,I57376,I57393,I57410,I56986,I57441,I56974,I56983,I56971,I57527,I832296,I57553,I57561,I57578,I832293,I832308,I57595,I832290,I57621,I832287,I57638,I57646,I57663,I57495,I57694,I57711,I57507,I57751,I57516,I57773,I832302,I57790,I832305,I57816,I57833,I57519,I57855,I57504,I57886,I832299,I57903,I57920,I57937,I57513,I57968,I57501,I57510,I57498,I58054,I457761,I58080,I58088,I58105,I457755,I457746,I58122,I457767,I58148,I457749,I58165,I58173,I457743,I58190,I58022,I58221,I58238,I58034,I58278,I58043,I58300,I457770,I457752,I58317,I457758,I58343,I58360,I58046,I58382,I58031,I58413,I457764,I58430,I58447,I58464,I58040,I58495,I58028,I58037,I58025,I58581,I846525,I58607,I58615,I58632,I846522,I846537,I58649,I846519,I58675,I846516,I58692,I58700,I58717,I58549,I58748,I58765,I58561,I58805,I58570,I58827,I846531,I58844,I846534,I58870,I58887,I58573,I58909,I58558,I58940,I846528,I58957,I58974,I58991,I58567,I59022,I58555,I58564,I58552,I59108,I877091,I59134,I59142,I59159,I877088,I877103,I59176,I877085,I59202,I877082,I59219,I59227,I59244,I59076,I59275,I59292,I59088,I59332,I59097,I59354,I877097,I59371,I877100,I59397,I59414,I59100,I59436,I59085,I59467,I877094,I59484,I59501,I59518,I59094,I59549,I59082,I59091,I59079,I59635,I360887,I59661,I59669,I59686,I360869,I360884,I59703,I360860,I59729,I360863,I59746,I59754,I360878,I59771,I59603,I59802,I59819,I59615,I360881,I59859,I59624,I59881,I360872,I59898,I360866,I59924,I59941,I59627,I59963,I59612,I59994,I360875,I60011,I60028,I60045,I59621,I60076,I59609,I59618,I59606,I60162,I592001,I60188,I60196,I60213,I592013,I591998,I60230,I591992,I60256,I592007,I60273,I60281,I591995,I60298,I60130,I60329,I60346,I60142,I592004,I60386,I60151,I60408,I592010,I592016,I60425,I60451,I60468,I60154,I60490,I60139,I60521,I60538,I60555,I60572,I60148,I60603,I60136,I60145,I60133,I60689,I339807,I60715,I60723,I60740,I339789,I339804,I60757,I339780,I60783,I339783,I60800,I60808,I339798,I60825,I60856,I60873,I339801,I60913,I60935,I339792,I60952,I339786,I60978,I60995,I61017,I61048,I339795,I61065,I61082,I61099,I61130,I61216,I61242,I61250,I61267,I61284,I61310,I61327,I61335,I61352,I61184,I61383,I61400,I61196,I61440,I61205,I61462,I61479,I61505,I61522,I61208,I61544,I61193,I61575,I61592,I61609,I61626,I61202,I61657,I61190,I61199,I61187,I61743,I715118,I61769,I61777,I61794,I715109,I715127,I61811,I715106,I61837,I61854,I61862,I715112,I61879,I61711,I61910,I61927,I61723,I61967,I61732,I61989,I715124,I715115,I62006,I715130,I62032,I62049,I61735,I62071,I61720,I62102,I715121,I62119,I62136,I62153,I61729,I62184,I61717,I61726,I61714,I62270,I196652,I62296,I62304,I62321,I196646,I196640,I62338,I196661,I62364,I196658,I62381,I62389,I196655,I62406,I62238,I62437,I62454,I62250,I62494,I62259,I62516,I196643,I62533,I196664,I62559,I62576,I62262,I62598,I62247,I62629,I196649,I62646,I62663,I62680,I62256,I62711,I62244,I62253,I62241,I62797,I1253672,I62823,I62831,I62848,I1253666,I1253687,I62865,I1253678,I62891,I1253669,I62908,I62916,I1253681,I62933,I62765,I62964,I62981,I62777,I63021,I62786,I63043,I1253690,I1253675,I63060,I63086,I63103,I62789,I63125,I62774,I63156,I1253684,I63173,I63190,I63207,I62783,I63238,I62771,I62780,I62768,I63324,I209742,I63350,I63358,I63375,I209736,I209730,I63392,I209751,I63418,I209748,I63435,I63443,I209745,I63460,I63292,I63491,I63508,I63304,I63548,I63313,I63570,I209733,I63587,I209754,I63613,I63630,I63316,I63652,I63301,I63683,I209739,I63700,I63717,I63734,I63310,I63765,I63298,I63307,I63295,I63851,I479521,I63877,I63885,I63902,I479515,I479506,I63919,I479527,I63945,I479509,I63962,I63970,I479503,I63987,I63819,I64018,I64035,I63831,I64075,I63840,I64097,I479530,I479512,I64114,I479518,I64140,I64157,I63843,I64179,I63828,I64210,I479524,I64227,I64244,I64261,I63837,I64292,I63825,I63834,I63822,I64378,I268135,I64404,I64412,I64429,I268117,I268132,I64446,I268108,I64472,I268111,I64489,I64497,I268126,I64514,I64346,I64545,I64562,I64358,I268129,I64602,I64367,I64624,I268120,I64641,I268114,I64667,I64684,I64370,I64706,I64355,I64737,I268123,I64754,I64771,I64788,I64364,I64819,I64352,I64361,I64349,I64905,I143706,I64931,I64939,I64956,I143703,I143685,I64973,I143691,I64999,I143700,I65016,I65024,I143694,I65041,I64873,I65072,I65089,I64885,I143709,I65129,I64894,I65151,I143697,I143688,I65168,I65194,I65211,I64897,I65233,I64882,I65264,I143712,I65281,I65298,I65315,I64891,I65346,I64879,I64888,I64876,I65432,I1290033,I65458,I65466,I65483,I1290036,I1290030,I65500,I1290027,I65526,I1290012,I65543,I65551,I1290021,I65568,I65400,I65599,I65616,I65412,I65656,I65421,I65678,I1290015,I1290018,I65695,I1290024,I65721,I65738,I65424,I65760,I65409,I65791,I65808,I65825,I65842,I65418,I65873,I65406,I65415,I65403,I65959,I181777,I65985,I65993,I66010,I181771,I181765,I66027,I181786,I66053,I181783,I66070,I66078,I181780,I66095,I65927,I66126,I66143,I65939,I66183,I65948,I66205,I181768,I66222,I181789,I66248,I66265,I65951,I66287,I65936,I66318,I181774,I66335,I66352,I66369,I65945,I66400,I65933,I65942,I65930,I66486,I399009,I66512,I66520,I66537,I399003,I398994,I66554,I399015,I66580,I398997,I66597,I66605,I398991,I66622,I66454,I66653,I66670,I66466,I66710,I66475,I66732,I399018,I399000,I66749,I399006,I66775,I66792,I66478,I66814,I66463,I66845,I399012,I66862,I66879,I66896,I66472,I66927,I66460,I66469,I66457,I67013,I907606,I67039,I67047,I67064,I907624,I907618,I67081,I907597,I67107,I907615,I67124,I67132,I907600,I67149,I66981,I67180,I67197,I66993,I907612,I67237,I67002,I67259,I907621,I907609,I67276,I907603,I67302,I67319,I67005,I67341,I66990,I67372,I67389,I67406,I67423,I66999,I67454,I66987,I66996,I66984,I67540,I685062,I67566,I67574,I67591,I685053,I685071,I67608,I685050,I67634,I67651,I67659,I685056,I67676,I67508,I67707,I67724,I67520,I67764,I67529,I67786,I685068,I685059,I67803,I685074,I67829,I67846,I67532,I67868,I67517,I67899,I685065,I67916,I67933,I67950,I67526,I67981,I67514,I67523,I67511,I68067,I144301,I68093,I68101,I68118,I144298,I144280,I68135,I144286,I68161,I144295,I68178,I68186,I144289,I68203,I68035,I68234,I68251,I68047,I144304,I68291,I68056,I68313,I144292,I144283,I68330,I68356,I68373,I68059,I68395,I68044,I68426,I144307,I68443,I68460,I68477,I68053,I68508,I68041,I68050,I68038,I68594,I476257,I68620,I68628,I68645,I476251,I476242,I68662,I476263,I68688,I476245,I68705,I68713,I476239,I68730,I68562,I68761,I68778,I68574,I68818,I68583,I68840,I476266,I476248,I68857,I476254,I68883,I68900,I68586,I68922,I68571,I68953,I476260,I68970,I68987,I69004,I68580,I69035,I68568,I68577,I68565,I69121,I1033145,I69147,I69155,I69172,I1033142,I1033148,I69189,I69215,I69232,I69240,I69257,I69089,I69288,I69305,I69101,I1033151,I69345,I69110,I69367,I1033154,I1033163,I69384,I1033157,I69410,I69427,I69113,I69449,I69098,I69480,I1033160,I69497,I69514,I69531,I69107,I69562,I69095,I69104,I69092,I69648,I797514,I69674,I69682,I69699,I797511,I797526,I69716,I797508,I69742,I797505,I69759,I69767,I69784,I69616,I69815,I69832,I69628,I69872,I69637,I69894,I797520,I69911,I797523,I69937,I69954,I69640,I69976,I69625,I70007,I797517,I70024,I70041,I70058,I69634,I70089,I69622,I69631,I69619,I70175,I872875,I70201,I70209,I70226,I872872,I872887,I70243,I872869,I70269,I872866,I70286,I70294,I70311,I70143,I70342,I70359,I70155,I70399,I70164,I70421,I872881,I70438,I872884,I70464,I70481,I70167,I70503,I70152,I70534,I872878,I70551,I70568,I70585,I70161,I70616,I70149,I70158,I70146,I70702,I1287143,I70728,I70736,I70753,I1287146,I1287140,I70770,I1287137,I70796,I1287122,I70813,I70821,I1287131,I70838,I70670,I70869,I70886,I70682,I70926,I70691,I70948,I1287125,I1287128,I70965,I1287134,I70991,I71008,I70694,I71030,I70679,I71061,I71078,I71095,I71112,I70688,I71143,I70676,I70685,I70673,I71229,I71255,I71263,I71280,I71297,I71323,I71340,I71348,I71365,I71197,I71396,I71413,I71209,I71453,I71218,I71475,I71492,I71518,I71535,I71221,I71557,I71206,I71588,I71605,I71622,I71639,I71215,I71670,I71203,I71212,I71200,I71756,I1345189,I71782,I71790,I71807,I1345183,I1345204,I71824,I1345180,I71850,I1345201,I71867,I71875,I1345198,I71892,I71724,I71923,I71940,I71736,I1345186,I71980,I71745,I72002,I1345195,I1345192,I72019,I1345177,I72045,I72062,I71748,I72084,I71733,I72115,I72132,I72149,I72166,I71742,I72197,I71730,I71739,I71727,I72283,I484961,I72309,I72317,I72334,I484955,I484946,I72351,I484967,I72377,I484949,I72394,I72402,I484943,I72419,I72251,I72450,I72467,I72263,I72507,I72272,I72529,I484970,I484952,I72546,I484958,I72572,I72589,I72275,I72611,I72260,I72642,I484964,I72659,I72676,I72693,I72269,I72724,I72257,I72266,I72254,I72810,I473537,I72836,I72844,I72861,I473531,I473522,I72878,I473543,I72904,I473525,I72921,I72929,I473519,I72946,I72778,I72977,I72994,I72790,I73034,I72799,I73056,I473546,I473528,I73073,I473534,I73099,I73116,I72802,I73138,I72787,I73169,I473540,I73186,I73203,I73220,I72796,I73251,I72784,I72793,I72781,I73337,I1243880,I73363,I73371,I73388,I1243874,I1243895,I73405,I1243886,I73431,I1243877,I73448,I73456,I1243889,I73473,I73305,I73504,I73521,I73317,I73561,I73326,I73583,I1243898,I1243883,I73600,I73626,I73643,I73329,I73665,I73314,I73696,I1243892,I73713,I73730,I73747,I73323,I73778,I73311,I73320,I73308,I73864,I280783,I73890,I73898,I73915,I280765,I280780,I73932,I280756,I73958,I280759,I73975,I73983,I280774,I74000,I73832,I74031,I74048,I73844,I280777,I74088,I73853,I74110,I280768,I74127,I280762,I74153,I74170,I73856,I74192,I73841,I74223,I280771,I74240,I74257,I74274,I73850,I74305,I73838,I73847,I73835,I74391,I254960,I74417,I74425,I74442,I254942,I254957,I74459,I254933,I74485,I254936,I74502,I74510,I254951,I74527,I74359,I74558,I74575,I74371,I254954,I74615,I74380,I74637,I254945,I74654,I254939,I74680,I74697,I74383,I74719,I74368,I74750,I254948,I74767,I74784,I74801,I74377,I74832,I74365,I74374,I74362,I74918,I835985,I74944,I74952,I74969,I835982,I835997,I74986,I835979,I75012,I835976,I75029,I75037,I75054,I74886,I75085,I75102,I74898,I75142,I74907,I75164,I835991,I75181,I835994,I75207,I75224,I74910,I75246,I74895,I75277,I835988,I75294,I75311,I75328,I74904,I75359,I74892,I74901,I74889,I75445,I223427,I75471,I75479,I75496,I223421,I223415,I75513,I223436,I75539,I223433,I75556,I75564,I223430,I75581,I75413,I75612,I75629,I75425,I75669,I75434,I75691,I223418,I75708,I223439,I75734,I75751,I75437,I75773,I75422,I75804,I223424,I75821,I75838,I75855,I75431,I75886,I75419,I75428,I75416,I75972,I1157214,I75998,I76006,I76023,I1157229,I1157208,I76040,I1157211,I76066,I1157232,I76083,I76091,I76108,I75940,I76139,I76156,I75952,I76196,I75961,I76218,I1157220,I1157217,I76235,I1157223,I76261,I76278,I75964,I76300,I75949,I76331,I1157226,I76348,I76365,I76382,I75958,I76413,I75946,I75955,I75943,I76499,I306606,I76525,I76533,I76550,I306588,I306603,I76567,I306579,I76593,I306582,I76610,I76618,I306597,I76635,I76467,I76666,I76683,I76479,I306600,I76723,I76488,I76745,I306591,I76762,I306585,I76788,I76805,I76491,I76827,I76476,I76858,I306594,I76875,I76892,I76909,I76485,I76940,I76473,I76482,I76470,I77026,I908898,I77052,I77060,I77077,I908916,I908910,I77094,I908889,I77120,I908907,I77137,I77145,I908892,I77162,I76994,I77193,I77210,I77006,I908904,I77250,I77015,I77272,I908913,I908901,I77289,I908895,I77315,I77332,I77018,I77354,I77003,I77385,I77402,I77419,I77436,I77012,I77467,I77000,I77009,I76997,I77553,I77579,I77587,I77604,I77621,I77647,I77664,I77672,I77689,I77521,I77720,I77737,I77533,I77777,I77542,I77799,I77816,I77842,I77859,I77545,I77881,I77530,I77912,I77929,I77946,I77963,I77539,I77994,I77527,I77536,I77524,I78080,I1095946,I78106,I78114,I78131,I1095961,I1095940,I78148,I1095943,I78174,I1095964,I78191,I78199,I78216,I78048,I78247,I78264,I78060,I78304,I78069,I78326,I1095952,I1095949,I78343,I1095955,I78369,I78386,I78072,I78408,I78057,I78439,I1095958,I78456,I78473,I78490,I78066,I78521,I78054,I78063,I78051,I78607,I78633,I78641,I78658,I78675,I78701,I78718,I78726,I78743,I78575,I78774,I78791,I78587,I78831,I78596,I78853,I78870,I78896,I78913,I78599,I78935,I78584,I78966,I78983,I79000,I79017,I78593,I79048,I78581,I78590,I78578,I79134,I529792,I79160,I79168,I79185,I529813,I529807,I79202,I529789,I79228,I79245,I79253,I529801,I79270,I79102,I79301,I79318,I79114,I529798,I79358,I79123,I79380,I529804,I529795,I79397,I79423,I79440,I79126,I79462,I79111,I79493,I529810,I79510,I79527,I79544,I79120,I79575,I79108,I79117,I79105,I79661,I1086120,I79687,I79695,I79712,I1086135,I1086114,I79729,I1086117,I79755,I1086138,I79772,I79780,I79797,I79629,I79828,I79845,I79641,I79885,I79650,I79907,I1086126,I1086123,I79924,I1086129,I79950,I79967,I79653,I79989,I79638,I80020,I1086132,I80037,I80054,I80071,I79647,I80102,I79635,I79644,I79632,I80188,I867078,I80214,I80222,I80239,I867075,I867090,I80256,I867072,I80282,I867069,I80299,I80307,I80324,I80156,I80355,I80372,I80168,I80412,I80177,I80434,I867084,I80451,I867087,I80477,I80494,I80180,I80516,I80165,I80547,I867081,I80564,I80581,I80598,I80174,I80629,I80162,I80171,I80159,I80715,I293958,I80741,I80749,I80766,I293940,I293955,I80783,I293931,I80809,I293934,I80826,I80834,I293949,I80851,I80683,I80882,I80899,I80695,I293952,I80939,I80704,I80961,I293943,I80978,I293937,I81004,I81021,I80707,I81043,I80692,I81074,I293946,I81091,I81108,I81125,I80701,I81156,I80689,I80698,I80686,I81242,I508967,I81268,I81276,I81293,I508988,I508982,I81310,I508964,I81336,I81353,I81361,I508976,I81378,I81210,I81409,I81426,I81222,I508973,I81466,I81231,I81488,I508979,I508970,I81505,I81531,I81548,I81234,I81570,I81219,I81601,I508985,I81618,I81635,I81652,I81228,I81683,I81216,I81225,I81213,I81769,I468097,I81795,I81803,I81820,I468091,I468082,I81837,I468103,I81863,I468085,I81880,I81888,I468079,I81905,I81737,I81936,I81953,I81749,I81993,I81758,I82015,I468106,I468088,I82032,I468094,I82058,I82075,I81761,I82097,I81746,I82128,I468100,I82145,I82162,I82179,I81755,I82210,I81743,I81752,I81740,I82296,I329794,I82322,I82330,I82347,I329776,I329791,I82364,I329767,I82390,I329770,I82407,I82415,I329785,I82432,I82264,I82463,I82480,I82276,I329788,I82520,I82285,I82542,I329779,I82559,I329773,I82585,I82602,I82288,I82624,I82273,I82655,I329782,I82672,I82689,I82706,I82282,I82737,I82270,I82279,I82267,I82823,I1164728,I82849,I82857,I82874,I1164743,I1164722,I82891,I1164725,I82917,I1164746,I82934,I82942,I82959,I82791,I82990,I83007,I82803,I83047,I82812,I83069,I1164734,I1164731,I83086,I1164737,I83112,I83129,I82815,I83151,I82800,I83182,I1164740,I83199,I83216,I83233,I82809,I83264,I82797,I82806,I82794,I83350,I760202,I83376,I83384,I83401,I760193,I760211,I83418,I760190,I83444,I83461,I83469,I760196,I83486,I83318,I83517,I83534,I83330,I83574,I83339,I83596,I760208,I760199,I83613,I760214,I83639,I83656,I83342,I83678,I83327,I83709,I760205,I83726,I83743,I83760,I83336,I83791,I83324,I83333,I83321,I83877,I191297,I83903,I83911,I83928,I191291,I191285,I83945,I191306,I83971,I191303,I83988,I83996,I191300,I84013,I83845,I84044,I84061,I83857,I84101,I83866,I84123,I191288,I84140,I191309,I84166,I84183,I83869,I84205,I83854,I84236,I191294,I84253,I84270,I84287,I83863,I84318,I83851,I83860,I83848,I84404,I1091900,I84430,I84438,I84455,I1091915,I1091894,I84472,I1091897,I84498,I1091918,I84515,I84523,I84540,I84372,I84571,I84588,I84384,I84628,I84393,I84650,I1091906,I1091903,I84667,I1091909,I84693,I84710,I84396,I84732,I84381,I84763,I1091912,I84780,I84797,I84814,I84390,I84845,I84378,I84387,I84375,I84931,I1278473,I84957,I84965,I84982,I1278476,I1278470,I84999,I1278467,I85025,I1278452,I85042,I85050,I1278461,I85067,I84899,I85098,I85115,I84911,I85155,I84920,I85177,I1278455,I1278458,I85194,I1278464,I85220,I85237,I84923,I85259,I84908,I85290,I85307,I85324,I85341,I84917,I85372,I84905,I84914,I84902,I85458,I390305,I85484,I85492,I85509,I390299,I390290,I85526,I390311,I85552,I390293,I85569,I85577,I390287,I85594,I85426,I85625,I85642,I85438,I85682,I85447,I85704,I390314,I390296,I85721,I390302,I85747,I85764,I85450,I85786,I85435,I85817,I390308,I85834,I85851,I85868,I85444,I85899,I85432,I85441,I85429,I85985,I607607,I86011,I86019,I86036,I607619,I607604,I86053,I607598,I86079,I607613,I86096,I86104,I607601,I86121,I85953,I86152,I86169,I85965,I607610,I86209,I85974,I86231,I607616,I607622,I86248,I86274,I86291,I85977,I86313,I85962,I86344,I86361,I86378,I86395,I85971,I86426,I85959,I85968,I85956,I86512,I1147388,I86538,I86546,I86563,I1147403,I1147382,I86580,I1147385,I86606,I1147406,I86623,I86631,I86648,I86480,I86679,I86696,I86492,I86736,I86501,I86758,I1147394,I1147391,I86775,I1147397,I86801,I86818,I86504,I86840,I86489,I86871,I1147400,I86888,I86905,I86922,I86498,I86953,I86486,I86495,I86483,I87039,I1151434,I87065,I87073,I87090,I1151449,I1151428,I87107,I1151431,I87133,I1151452,I87150,I87158,I87175,I87007,I87206,I87223,I87019,I87263,I87028,I87285,I1151440,I1151437,I87302,I1151443,I87328,I87345,I87031,I87367,I87016,I87398,I1151446,I87415,I87432,I87449,I87025,I87480,I87013,I87022,I87010,I87566,I1252584,I87592,I87600,I87617,I1252578,I1252599,I87634,I1252590,I87660,I1252581,I87677,I87685,I1252593,I87702,I87534,I87733,I87750,I87546,I87790,I87555,I87812,I1252602,I1252587,I87829,I87855,I87872,I87558,I87894,I87543,I87925,I1252596,I87942,I87959,I87976,I87552,I88007,I87540,I87549,I87537,I88093,I1336264,I88119,I88127,I88144,I1336258,I1336279,I88161,I1336255,I88187,I1336276,I88204,I88212,I1336273,I88229,I88061,I88260,I88277,I88073,I1336261,I88317,I88082,I88339,I1336270,I1336267,I88356,I1336252,I88382,I88399,I88085,I88421,I88070,I88452,I88469,I88486,I88503,I88079,I88534,I88067,I88076,I88064,I88620,I533957,I88646,I88654,I88671,I533978,I533972,I88688,I533954,I88714,I88731,I88739,I533966,I88756,I88588,I88787,I88804,I88600,I533963,I88844,I88609,I88866,I533969,I533960,I88883,I88909,I88926,I88612,I88948,I88597,I88979,I533975,I88996,I89013,I89030,I88606,I89061,I88594,I88603,I88591,I89147,I663098,I89173,I89181,I89198,I663089,I663107,I89215,I663086,I89241,I89258,I89266,I663092,I89283,I89115,I89314,I89331,I89127,I89371,I89136,I89393,I663104,I663095,I89410,I663110,I89436,I89453,I89139,I89475,I89124,I89506,I663101,I89523,I89540,I89557,I89133,I89588,I89121,I89130,I89118,I89674,I467009,I89700,I89708,I89725,I467003,I466994,I89742,I467015,I89768,I466997,I89785,I89793,I466991,I89810,I89642,I89841,I89858,I89654,I89898,I89663,I89920,I467018,I467000,I89937,I467006,I89963,I89980,I89666,I90002,I89651,I90033,I467012,I90050,I90067,I90084,I89660,I90115,I89648,I89657,I89645,I90201,I90227,I90235,I90252,I90269,I90295,I90312,I90320,I90337,I90368,I90385,I90425,I90447,I90464,I90490,I90507,I90529,I90560,I90577,I90594,I90611,I90642,I90728,I905668,I90754,I90762,I90779,I905686,I905680,I90796,I905659,I90822,I905677,I90839,I90847,I905662,I90864,I90696,I90895,I90912,I90708,I905674,I90952,I90717,I90974,I905683,I905671,I90991,I905665,I91017,I91034,I90720,I91056,I90705,I91087,I91104,I91121,I91138,I90714,I91169,I90702,I90711,I90699,I91255,I1247688,I91281,I91289,I91306,I1247682,I1247703,I91323,I1247694,I91349,I1247685,I91366,I91374,I1247697,I91391,I91223,I91422,I91439,I91235,I91479,I91244,I91501,I1247706,I1247691,I91518,I91544,I91561,I91247,I91583,I91232,I91614,I1247700,I91631,I91648,I91665,I91241,I91696,I91229,I91238,I91226,I91782,I152622,I91808,I91816,I91833,I152616,I152610,I91850,I152631,I91876,I152628,I91893,I91901,I152625,I91918,I91750,I91949,I91966,I91762,I92006,I91771,I92028,I152613,I92045,I152634,I92071,I92088,I91774,I92110,I91759,I92141,I152619,I92158,I92175,I92192,I91768,I92223,I91756,I91765,I91753,I92309,I747486,I92335,I92343,I92360,I747477,I747495,I92377,I747474,I92403,I92420,I92428,I747480,I92445,I92277,I92476,I92493,I92289,I92533,I92298,I92555,I747492,I747483,I92572,I747498,I92598,I92615,I92301,I92637,I92286,I92668,I747489,I92685,I92702,I92719,I92295,I92750,I92283,I92292,I92280,I92836,I1234088,I92862,I92870,I92887,I1234082,I1234103,I92904,I1234094,I92930,I1234085,I92947,I92955,I1234097,I92972,I92804,I93003,I93020,I92816,I93060,I92825,I93082,I1234106,I1234091,I93099,I93125,I93142,I92828,I93164,I92813,I93195,I1234100,I93212,I93229,I93246,I92822,I93277,I92810,I92819,I92807,I93363,I246037,I93389,I93397,I93414,I246031,I246025,I93431,I246046,I93457,I246043,I93474,I93482,I246040,I93499,I93331,I93530,I93547,I93343,I93587,I93352,I93609,I246028,I93626,I246049,I93652,I93669,I93355,I93691,I93340,I93722,I246034,I93739,I93756,I93773,I93349,I93804,I93337,I93346,I93334,I93890,I895978,I93916,I93924,I93941,I895996,I895990,I93958,I895969,I93984,I895987,I94001,I94009,I895972,I94026,I93858,I94057,I94074,I93870,I895984,I94114,I93879,I94136,I895993,I895981,I94153,I895975,I94179,I94196,I93882,I94218,I93867,I94249,I94266,I94283,I94300,I93876,I94331,I93864,I93873,I93861,I94417,I955410,I94443,I94451,I94468,I955428,I955422,I94485,I955401,I94511,I955419,I94528,I94536,I955404,I94553,I94385,I94584,I94601,I94397,I955416,I94641,I94406,I94663,I955425,I955413,I94680,I955407,I94706,I94723,I94409,I94745,I94394,I94776,I94793,I94810,I94827,I94403,I94858,I94391,I94400,I94388,I94944,I553853,I94970,I94978,I94995,I553865,I553850,I95012,I553844,I95038,I553859,I95055,I95063,I553847,I95080,I94912,I95111,I95128,I94924,I553856,I95168,I94933,I95190,I553862,I553868,I95207,I95233,I95250,I94936,I95272,I94921,I95303,I95320,I95337,I95354,I94930,I95385,I94918,I94927,I94915,I95471,I272878,I95497,I95505,I95522,I272860,I272875,I95539,I272851,I95565,I272854,I95582,I95590,I272869,I95607,I95439,I95638,I95655,I95451,I272872,I95695,I95460,I95717,I272863,I95734,I272857,I95760,I95777,I95463,I95799,I95448,I95830,I272866,I95847,I95864,I95881,I95457,I95912,I95445,I95454,I95442,I95998,I370373,I96024,I96032,I96049,I370355,I370370,I96066,I370346,I96092,I370349,I96109,I96117,I370364,I96134,I95966,I96165,I96182,I95978,I370367,I96222,I95987,I96244,I370358,I96261,I370352,I96287,I96304,I95990,I96326,I95975,I96357,I370361,I96374,I96391,I96408,I95984,I96439,I95972,I95981,I95969,I96525,I1261133,I96551,I96559,I96576,I1261136,I1261130,I96593,I1261127,I96619,I1261112,I96636,I96644,I1261121,I96661,I96493,I96692,I96709,I96505,I96749,I96514,I96771,I1261115,I1261118,I96788,I1261124,I96814,I96831,I96517,I96853,I96502,I96884,I96901,I96918,I96935,I96511,I96966,I96499,I96508,I96496,I97052,I750376,I97078,I97086,I97103,I750367,I750385,I97120,I750364,I97146,I97163,I97171,I750370,I97188,I97020,I97219,I97236,I97032,I97276,I97041,I97298,I750382,I750373,I97315,I750388,I97341,I97358,I97044,I97380,I97029,I97411,I750379,I97428,I97445,I97462,I97038,I97493,I97026,I97035,I97023,I97579,I672346,I97605,I97613,I97630,I672337,I672355,I97647,I672334,I97673,I97690,I97698,I672340,I97715,I97547,I97746,I97763,I97559,I97803,I97568,I97825,I672352,I672343,I97842,I672358,I97868,I97885,I97571,I97907,I97556,I97938,I672349,I97955,I97972,I97989,I97565,I98020,I97553,I97562,I97550,I98106,I847052,I98132,I98140,I98157,I847049,I847064,I98174,I847046,I98200,I847043,I98217,I98225,I98242,I98074,I98273,I98290,I98086,I98330,I98095,I98352,I847058,I98369,I847061,I98395,I98412,I98098,I98434,I98083,I98465,I847055,I98482,I98499,I98516,I98092,I98547,I98080,I98089,I98077,I98633,I509562,I98659,I98667,I98684,I509583,I509577,I98701,I509559,I98727,I98744,I98752,I509571,I98769,I98601,I98800,I98817,I98613,I509568,I98857,I98622,I98879,I509574,I509565,I98896,I98922,I98939,I98625,I98961,I98610,I98992,I509580,I99009,I99026,I99043,I98619,I99074,I98607,I98616,I98604,I99160,I565413,I99186,I99194,I99211,I565425,I565410,I99228,I565404,I99254,I565419,I99271,I99279,I565407,I99296,I99128,I99327,I99344,I99140,I565416,I99384,I99149,I99406,I565422,I565428,I99423,I99449,I99466,I99152,I99488,I99137,I99519,I99536,I99553,I99570,I99146,I99601,I99134,I99143,I99131,I99687,I99713,I99721,I99738,I99755,I99781,I99798,I99806,I99823,I99655,I99854,I99871,I99667,I99911,I99676,I99933,I99950,I99976,I99993,I99679,I100015,I99664,I100046,I100063,I100080,I100097,I99673,I100128,I99661,I99670,I99658,I100214,I938614,I100240,I100248,I100265,I938632,I938626,I100282,I938605,I100308,I938623,I100325,I100333,I938608,I100350,I100182,I100381,I100398,I100194,I938620,I100438,I100203,I100460,I938629,I938617,I100477,I938611,I100503,I100520,I100206,I100542,I100191,I100573,I100590,I100607,I100624,I100200,I100655,I100188,I100197,I100185,I100741,I1167040,I100767,I100775,I100792,I1167055,I1167034,I100809,I1167037,I100835,I1167058,I100852,I100860,I100877,I100709,I100908,I100925,I100721,I100965,I100730,I100987,I1167046,I1167043,I101004,I1167049,I101030,I101047,I100733,I101069,I100718,I101100,I1167052,I101117,I101134,I101151,I100727,I101182,I100715,I100724,I100712,I101268,I1340429,I101294,I101302,I101319,I1340423,I1340444,I101336,I1340420,I101362,I1340441,I101379,I101387,I1340438,I101404,I101236,I101435,I101452,I101248,I1340426,I101492,I101257,I101514,I1340435,I1340432,I101531,I1340417,I101557,I101574,I101260,I101596,I101245,I101627,I101644,I101661,I101678,I101254,I101709,I101242,I101251,I101239,I101795,I188322,I101821,I101829,I101846,I188316,I188310,I101863,I188331,I101889,I188328,I101906,I101914,I188325,I101931,I101763,I101962,I101979,I101775,I102019,I101784,I102041,I188313,I102058,I188334,I102084,I102101,I101787,I102123,I101772,I102154,I188319,I102171,I102188,I102205,I101781,I102236,I101769,I101778,I101766,I102322,I1336859,I102348,I102356,I102373,I1336853,I1336874,I102390,I1336850,I102416,I1336871,I102433,I102441,I1336868,I102458,I102290,I102489,I102506,I102302,I1336856,I102546,I102311,I102568,I1336865,I1336862,I102585,I1336847,I102611,I102628,I102314,I102650,I102299,I102681,I102698,I102715,I102732,I102308,I102763,I102296,I102305,I102293,I102849,I235922,I102875,I102883,I102900,I235916,I235910,I102917,I235931,I102943,I235928,I102960,I102968,I235925,I102985,I102817,I103016,I103033,I102829,I103073,I102838,I103095,I235913,I103112,I235934,I103138,I103155,I102841,I103177,I102826,I103208,I235919,I103225,I103242,I103259,I102835,I103290,I102823,I102832,I102820,I103376,I923756,I103402,I103410,I103427,I923774,I923768,I103444,I923747,I103470,I923765,I103487,I103495,I923750,I103512,I103344,I103543,I103560,I103356,I923762,I103600,I103365,I103622,I923771,I923759,I103639,I923753,I103665,I103682,I103368,I103704,I103353,I103735,I103752,I103769,I103786,I103362,I103817,I103350,I103359,I103347,I103903,I1028096,I103929,I103937,I103954,I1028093,I1028099,I103971,I103997,I104014,I104022,I104039,I103871,I104070,I104087,I103883,I1028102,I104127,I103892,I104149,I1028105,I1028114,I104166,I1028108,I104192,I104209,I103895,I104231,I103880,I104262,I1028111,I104279,I104296,I104313,I103889,I104344,I103877,I103886,I103874,I104430,I1356494,I104456,I104464,I104481,I1356488,I1356509,I104498,I1356485,I104524,I1356506,I104541,I104549,I1356503,I104566,I104398,I104597,I104614,I104410,I1356491,I104654,I104419,I104676,I1356500,I1356497,I104693,I1356482,I104719,I104736,I104422,I104758,I104407,I104789,I104806,I104823,I104840,I104416,I104871,I104404,I104413,I104401,I104957,I911482,I104983,I104991,I105008,I911500,I911494,I105025,I911473,I105051,I911491,I105068,I105076,I911476,I105093,I104925,I105124,I105141,I104937,I911488,I105181,I104946,I105203,I911497,I911485,I105220,I911479,I105246,I105263,I104949,I105285,I104934,I105316,I105333,I105350,I105367,I104943,I105398,I104931,I104940,I104928,I105484,I1360659,I105510,I105518,I105535,I1360653,I1360674,I105552,I1360650,I105578,I1360671,I105595,I105603,I1360668,I105620,I105452,I105651,I105668,I105464,I1360656,I105708,I105473,I105730,I1360665,I1360662,I105747,I1360647,I105773,I105790,I105476,I105812,I105461,I105843,I105860,I105877,I105894,I105470,I105925,I105458,I105467,I105455,I106011,I377249,I106037,I106045,I106062,I377243,I377234,I106079,I377255,I106105,I377237,I106122,I106130,I377231,I106147,I105979,I106178,I106195,I105991,I106235,I106000,I106257,I377258,I377240,I106274,I377246,I106300,I106317,I106003,I106339,I105988,I106370,I377252,I106387,I106404,I106421,I105997,I106452,I105985,I105994,I105982,I106538,I312930,I106564,I106572,I106589,I312912,I312927,I106606,I312903,I106632,I312906,I106649,I106657,I312921,I106674,I106506,I106705,I106722,I106518,I312924,I106762,I106527,I106784,I312915,I106801,I312909,I106827,I106844,I106530,I106866,I106515,I106897,I312918,I106914,I106931,I106948,I106524,I106979,I106512,I106521,I106509,I107065,I523247,I107091,I107099,I107116,I523268,I523262,I107133,I523244,I107159,I107176,I107184,I523256,I107201,I107033,I107232,I107249,I107045,I523253,I107289,I107054,I107311,I523259,I523250,I107328,I107354,I107371,I107057,I107393,I107042,I107424,I523265,I107441,I107458,I107475,I107051,I107506,I107039,I107048,I107036,I107592,I888872,I107618,I107626,I107643,I888890,I888884,I107660,I888863,I107686,I888881,I107703,I107711,I888866,I107728,I107560,I107759,I107776,I107572,I888878,I107816,I107581,I107838,I888887,I888875,I107855,I888869,I107881,I107898,I107584,I107920,I107569,I107951,I107968,I107985,I108002,I107578,I108033,I107566,I107575,I107563,I108119,I778542,I108145,I108153,I108170,I778539,I778554,I108187,I778536,I108213,I778533,I108230,I108238,I108255,I108087,I108286,I108303,I108099,I108343,I108108,I108365,I778548,I108382,I778551,I108408,I108425,I108111,I108447,I108096,I108478,I778545,I108495,I108512,I108529,I108105,I108560,I108093,I108102,I108090,I108646,I513132,I108672,I108680,I108697,I513153,I513147,I108714,I513129,I108740,I108757,I108765,I513141,I108782,I108614,I108813,I108830,I108626,I513138,I108870,I108635,I108892,I513144,I513135,I108909,I108935,I108952,I108638,I108974,I108623,I109005,I513150,I109022,I109039,I109056,I108632,I109087,I108620,I108629,I108617,I109173,I839674,I109199,I109207,I109224,I839671,I839686,I109241,I839668,I109267,I839665,I109284,I109292,I109309,I109141,I109340,I109357,I109153,I109397,I109162,I109419,I839680,I109436,I839683,I109462,I109479,I109165,I109501,I109150,I109532,I839677,I109549,I109566,I109583,I109159,I109614,I109147,I109156,I109144,I109700,I822283,I109726,I109734,I109751,I822280,I822295,I109768,I822277,I109794,I822274,I109811,I109819,I109836,I109668,I109867,I109884,I109680,I109924,I109689,I109946,I822289,I109963,I822292,I109989,I110006,I109692,I110028,I109677,I110059,I822286,I110076,I110093,I110110,I109686,I110141,I109674,I109683,I109671,I110227,I391393,I110253,I110261,I110278,I391387,I391378,I110295,I391399,I110321,I391381,I110338,I110346,I391375,I110363,I110195,I110394,I110411,I110207,I110451,I110216,I110473,I391402,I391384,I110490,I391390,I110516,I110533,I110219,I110555,I110204,I110586,I391396,I110603,I110620,I110637,I110213,I110668,I110201,I110210,I110198,I110754,I809108,I110780,I110788,I110805,I809105,I809120,I110822,I809102,I110848,I809099,I110865,I110873,I110890,I110722,I110921,I110938,I110734,I110978,I110743,I111000,I809114,I111017,I809117,I111043,I111060,I110746,I111082,I110731,I111113,I809111,I111130,I111147,I111164,I110740,I111195,I110728,I110737,I110725,I111281,I814905,I111307,I111315,I111332,I814902,I814917,I111349,I814899,I111375,I814896,I111392,I111400,I111417,I111249,I111448,I111465,I111261,I111505,I111270,I111527,I814911,I111544,I814914,I111570,I111587,I111273,I111609,I111258,I111640,I814908,I111657,I111674,I111691,I111267,I111722,I111255,I111264,I111252,I111808,I1386244,I111834,I111842,I111859,I1386238,I1386259,I111876,I1386235,I111902,I1386256,I111919,I111927,I1386253,I111944,I111776,I111975,I111992,I111788,I1386241,I112032,I111797,I112054,I1386250,I1386247,I112071,I1386232,I112097,I112114,I111800,I112136,I111785,I112167,I112184,I112201,I112218,I111794,I112249,I111782,I111791,I111779,I112335,I410977,I112361,I112369,I112386,I410971,I410962,I112403,I410983,I112429,I410965,I112446,I112454,I410959,I112471,I112303,I112502,I112519,I112315,I112559,I112324,I112581,I410986,I410968,I112598,I410974,I112624,I112641,I112327,I112663,I112312,I112694,I410980,I112711,I112728,I112745,I112321,I112776,I112309,I112318,I112306,I112862,I1329719,I112888,I112896,I112913,I1329713,I1329734,I112930,I1329710,I112956,I1329731,I112973,I112981,I1329728,I112998,I112830,I113029,I113046,I112842,I1329716,I113086,I112851,I113108,I1329725,I1329722,I113125,I1329707,I113151,I113168,I112854,I113190,I112839,I113221,I113238,I113255,I113272,I112848,I113303,I112836,I112845,I112833,I113389,I113415,I113423,I113440,I113457,I113483,I113500,I113508,I113525,I113556,I113573,I113613,I113635,I113652,I113678,I113695,I113717,I113748,I113765,I113782,I113799,I113830,I113916,I705292,I113942,I113950,I113967,I705283,I705301,I113984,I705280,I114010,I114027,I114035,I705286,I114052,I113884,I114083,I114100,I113896,I114140,I113905,I114162,I705298,I705289,I114179,I705304,I114205,I114222,I113908,I114244,I113893,I114275,I705295,I114292,I114309,I114326,I113902,I114357,I113890,I113899,I113887,I114443,I1241704,I114469,I114477,I114494,I1241698,I1241719,I114511,I1241710,I114537,I1241701,I114554,I114562,I1241713,I114579,I114411,I114610,I114627,I114423,I114667,I114432,I114689,I1241722,I1241707,I114706,I114732,I114749,I114435,I114771,I114420,I114802,I1241716,I114819,I114836,I114853,I114429,I114884,I114417,I114426,I114414,I114970,I326105,I114996,I115004,I115021,I326087,I326102,I115038,I326078,I115064,I326081,I115081,I115089,I326096,I115106,I114938,I115137,I115154,I114950,I326099,I115194,I114959,I115216,I326090,I115233,I326084,I115259,I115276,I114962,I115298,I114947,I115329,I326093,I115346,I115363,I115380,I114956,I115411,I114944,I114953,I114941,I115497,I376705,I115523,I115531,I115548,I376699,I376690,I115565,I376711,I115591,I376693,I115608,I115616,I376687,I115633,I115465,I115664,I115681,I115477,I115721,I115486,I115743,I376714,I376696,I115760,I376702,I115786,I115803,I115489,I115825,I115474,I115856,I376708,I115873,I115890,I115907,I115483,I115938,I115471,I115480,I115468,I116024,I157977,I116050,I116058,I116075,I157971,I157965,I116092,I157986,I116118,I157983,I116135,I116143,I157980,I116160,I115992,I116191,I116208,I116004,I116248,I116013,I116270,I157968,I116287,I157989,I116313,I116330,I116016,I116352,I116001,I116383,I157974,I116400,I116417,I116434,I116010,I116465,I115998,I116007,I115995,I116551,I798568,I116577,I116585,I116602,I798565,I798580,I116619,I798562,I116645,I798559,I116662,I116670,I116687,I116519,I116718,I116735,I116531,I116775,I116540,I116797,I798574,I116814,I798577,I116840,I116857,I116543,I116879,I116528,I116910,I798571,I116927,I116944,I116961,I116537,I116992,I116525,I116534,I116522,I117078,I494209,I117104,I117112,I117129,I494203,I494194,I117146,I494215,I117172,I494197,I117189,I117197,I494191,I117214,I117046,I117245,I117262,I117058,I117302,I117067,I117324,I494218,I494200,I117341,I494206,I117367,I117384,I117070,I117406,I117055,I117437,I494212,I117454,I117471,I117488,I117064,I117519,I117052,I117061,I117049,I117605,I894040,I117631,I117639,I117656,I894058,I894052,I117673,I894031,I117699,I894049,I117716,I117724,I894034,I117741,I117573,I117772,I117789,I117585,I894046,I117829,I117594,I117851,I894055,I894043,I117868,I894037,I117894,I117911,I117597,I117933,I117582,I117964,I117981,I117998,I118015,I117591,I118046,I117579,I117588,I117576,I118132,I843890,I118158,I118166,I118183,I843887,I843902,I118200,I843884,I118226,I843881,I118243,I118251,I118268,I118100,I118299,I118316,I118112,I118356,I118121,I118378,I843896,I118395,I843899,I118421,I118438,I118124,I118460,I118109,I118491,I843893,I118508,I118525,I118542,I118118,I118573,I118106,I118115,I118103,I118659,I380513,I118685,I118693,I118710,I380507,I380498,I118727,I380519,I118753,I380501,I118770,I118778,I380495,I118795,I118627,I118826,I118843,I118639,I118883,I118648,I118905,I380522,I380504,I118922,I380510,I118948,I118965,I118651,I118987,I118636,I119018,I380516,I119035,I119052,I119069,I118645,I119100,I118633,I118642,I118630,I119186,I1192472,I119212,I119220,I119237,I1192487,I1192466,I119254,I1192469,I119280,I1192490,I119297,I119305,I119322,I119154,I119353,I119370,I119166,I119410,I119175,I119432,I1192478,I1192475,I119449,I1192481,I119475,I119492,I119178,I119514,I119163,I119545,I1192484,I119562,I119579,I119596,I119172,I119627,I119160,I119169,I119157,I119713,I300809,I119739,I119747,I119764,I300791,I300806,I119781,I300782,I119807,I300785,I119824,I119832,I300800,I119849,I119681,I119880,I119897,I119693,I300803,I119937,I119702,I119959,I300794,I119976,I300788,I120002,I120019,I119705,I120041,I119690,I120072,I300797,I120089,I120106,I120123,I119699,I120154,I119687,I119696,I119684,I120240,I503612,I120266,I120274,I120291,I503633,I503627,I120308,I503609,I120334,I120351,I120359,I503621,I120376,I120208,I120407,I120424,I120220,I503618,I120464,I120229,I120486,I503624,I503615,I120503,I120529,I120546,I120232,I120568,I120217,I120599,I503630,I120616,I120633,I120650,I120226,I120681,I120214,I120223,I120211,I120767,I375116,I120793,I120801,I120818,I375098,I375113,I120835,I375089,I120861,I375092,I120878,I120886,I375107,I120903,I120735,I120934,I120951,I120747,I375110,I120991,I120756,I121013,I375101,I121030,I375095,I121056,I121073,I120759,I121095,I120744,I121126,I375104,I121143,I121160,I121177,I120753,I121208,I120741,I120750,I120738,I121294,I812270,I121320,I121328,I121345,I812267,I812282,I121362,I812264,I121388,I812261,I121405,I121413,I121430,I121262,I121461,I121478,I121274,I121518,I121283,I121540,I812276,I121557,I812279,I121583,I121600,I121286,I121622,I121271,I121653,I812273,I121670,I121687,I121704,I121280,I121735,I121268,I121277,I121265,I121821,I800676,I121847,I121855,I121872,I800673,I800688,I121889,I800670,I121915,I800667,I121932,I121940,I121957,I121789,I121988,I122005,I121801,I122045,I121810,I122067,I800682,I122084,I800685,I122110,I122127,I121813,I122149,I121798,I122180,I800679,I122197,I122214,I122231,I121807,I122262,I121795,I121804,I121792,I122348,I1223752,I122374,I122382,I122399,I1223746,I1223767,I122416,I1223758,I122442,I1223749,I122459,I122467,I1223761,I122484,I122316,I122515,I122532,I122328,I122572,I122337,I122594,I1223770,I1223755,I122611,I122637,I122654,I122340,I122676,I122325,I122707,I1223764,I122724,I122741,I122758,I122334,I122789,I122322,I122331,I122319,I122875,I948950,I122901,I122909,I122926,I948968,I948962,I122943,I948941,I122969,I948959,I122986,I122994,I948944,I123011,I122843,I123042,I123059,I122855,I948956,I123099,I122864,I123121,I948965,I948953,I123138,I948947,I123164,I123181,I122867,I123203,I122852,I123234,I123251,I123268,I123285,I122861,I123316,I122849,I122858,I122846,I123402,I580441,I123428,I123436,I123453,I580453,I580438,I123470,I580432,I123496,I580447,I123513,I123521,I580435,I123538,I123370,I123569,I123586,I123382,I580444,I123626,I123391,I123648,I580450,I580456,I123665,I123691,I123708,I123394,I123730,I123379,I123761,I123778,I123795,I123812,I123388,I123843,I123376,I123385,I123373,I123929,I217477,I123955,I123963,I123980,I217471,I217465,I123997,I217486,I124023,I217483,I124040,I124048,I217480,I124065,I123897,I124096,I124113,I123909,I124153,I123918,I124175,I217468,I124192,I217489,I124218,I124235,I123921,I124257,I123906,I124288,I217474,I124305,I124322,I124339,I123915,I124370,I123903,I123912,I123900,I124456,I1031462,I124482,I124490,I124507,I1031459,I1031465,I124524,I124550,I124567,I124575,I124592,I124424,I124623,I124640,I124436,I1031468,I124680,I124445,I124702,I1031471,I1031480,I124719,I1031474,I124745,I124762,I124448,I124784,I124433,I124815,I1031477,I124832,I124849,I124866,I124442,I124897,I124430,I124439,I124427,I124983,I878145,I125009,I125017,I125034,I878142,I878157,I125051,I878139,I125077,I878136,I125094,I125102,I125119,I124951,I125150,I125167,I124963,I125207,I124972,I125229,I878151,I125246,I878154,I125272,I125289,I124975,I125311,I124960,I125342,I878148,I125359,I125376,I125393,I124969,I125424,I124957,I124966,I124954,I125510,I671768,I125536,I125544,I125561,I671759,I671777,I125578,I671756,I125604,I125621,I125629,I671762,I125646,I125478,I125677,I125694,I125490,I125734,I125499,I125756,I671774,I671765,I125773,I671780,I125799,I125816,I125502,I125838,I125487,I125869,I671771,I125886,I125903,I125920,I125496,I125951,I125484,I125493,I125481,I126037,I418049,I126063,I126071,I126088,I418043,I418034,I126105,I418055,I126131,I418037,I126148,I126156,I418031,I126173,I126005,I126204,I126221,I126017,I126261,I126026,I126283,I418058,I418040,I126300,I418046,I126326,I126343,I126029,I126365,I126014,I126396,I418052,I126413,I126430,I126447,I126023,I126478,I126011,I126020,I126008,I126564,I1079762,I126590,I126598,I126615,I1079777,I1079756,I126632,I1079759,I126658,I1079780,I126675,I126683,I126700,I126532,I126731,I126748,I126544,I126788,I126553,I126810,I1079768,I1079765,I126827,I1079771,I126853,I126870,I126556,I126892,I126541,I126923,I1079774,I126940,I126957,I126974,I126550,I127005,I126538,I126547,I126535,I127091,I1291767,I127117,I127125,I127142,I1291770,I1291764,I127159,I1291761,I127185,I1291746,I127202,I127210,I1291755,I127227,I127059,I127258,I127275,I127071,I127315,I127080,I127337,I1291749,I1291752,I127354,I1291758,I127380,I127397,I127083,I127419,I127068,I127450,I127467,I127484,I127501,I127077,I127532,I127065,I127074,I127062,I127618,I494753,I127644,I127652,I127669,I494747,I494738,I127686,I494759,I127712,I494741,I127729,I127737,I494735,I127754,I127586,I127785,I127802,I127598,I127842,I127607,I127864,I494762,I494744,I127881,I494750,I127907,I127924,I127610,I127946,I127595,I127977,I494756,I127994,I128011,I128028,I127604,I128059,I127592,I127601,I127589,I128145,I235327,I128171,I128179,I128196,I235321,I235315,I128213,I235336,I128239,I235333,I128256,I128264,I235330,I128281,I128113,I128312,I128329,I128125,I128369,I128134,I128391,I235318,I128408,I235339,I128434,I128451,I128137,I128473,I128122,I128504,I235324,I128521,I128538,I128555,I128131,I128586,I128119,I128128,I128116,I128672,I128698,I128706,I128723,I128740,I128766,I128783,I128791,I128808,I128640,I128839,I128856,I128652,I128896,I128661,I128918,I128935,I128961,I128978,I128664,I129000,I128649,I129031,I129048,I129065,I129082,I128658,I129113,I128646,I128655,I128643,I129199,I798041,I129225,I129233,I129250,I798038,I798053,I129267,I798035,I129293,I798032,I129310,I129318,I129335,I129167,I129366,I129383,I129179,I129423,I129188,I129445,I798047,I129462,I798050,I129488,I129505,I129191,I129527,I129176,I129558,I798044,I129575,I129592,I129609,I129185,I129640,I129173,I129182,I129170,I129726,I753266,I129752,I129760,I129777,I753257,I753275,I129794,I753254,I129820,I129837,I129845,I753260,I129862,I129694,I129893,I129910,I129706,I129950,I129715,I129972,I753272,I753263,I129989,I753278,I130015,I130032,I129718,I130054,I129703,I130085,I753269,I130102,I130119,I130136,I129712,I130167,I129700,I129709,I129697,I130253,I1064156,I130279,I130287,I130304,I1064171,I1064150,I130321,I1064153,I130347,I1064174,I130364,I130372,I130389,I130221,I130420,I130437,I130233,I130477,I130242,I130499,I1064162,I1064159,I130516,I1064165,I130542,I130559,I130245,I130581,I130230,I130612,I1064168,I130629,I130646,I130663,I130239,I130694,I130227,I130236,I130224,I130780,I1209064,I130806,I130814,I130831,I1209058,I1209079,I130848,I1209070,I130874,I1209061,I130891,I130899,I1209073,I130916,I130748,I130947,I130964,I130760,I131004,I130769,I131026,I1209082,I1209067,I131043,I131069,I131086,I130772,I131108,I130757,I131139,I1209076,I131156,I131173,I131190,I130766,I131221,I130754,I130763,I130751,I131307,I131333,I131341,I131358,I131375,I131401,I131418,I131426,I131443,I131275,I131474,I131491,I131287,I131531,I131296,I131553,I131570,I131596,I131613,I131299,I131635,I131284,I131666,I131683,I131700,I131717,I131293,I131748,I131281,I131290,I131278,I131834,I1353519,I131860,I131868,I131885,I1353513,I1353534,I131902,I1353510,I131928,I1353531,I131945,I131953,I1353528,I131970,I131802,I132001,I132018,I131814,I1353516,I132058,I131823,I132080,I1353525,I1353522,I132097,I1353507,I132123,I132140,I131826,I132162,I131811,I132193,I132210,I132227,I132244,I131820,I132275,I131808,I131817,I131805,I132361,I596047,I132387,I132395,I132412,I596059,I596044,I132429,I596038,I132455,I596053,I132472,I132480,I596041,I132497,I132329,I132528,I132545,I132341,I596050,I132585,I132350,I132607,I596056,I596062,I132624,I132650,I132667,I132353,I132689,I132338,I132720,I132737,I132754,I132771,I132347,I132802,I132335,I132344,I132332,I132888,I1098836,I132914,I132922,I132939,I1098851,I1098830,I132956,I1098833,I132982,I1098854,I132999,I133007,I133024,I132856,I133055,I133072,I132868,I133112,I132877,I133134,I1098842,I1098839,I133151,I1098845,I133177,I133194,I132880,I133216,I132865,I133247,I1098848,I133264,I133281,I133298,I132874,I133329,I132862,I132871,I132859,I133415,I864443,I133441,I133449,I133466,I864440,I864455,I133483,I864437,I133509,I864434,I133526,I133534,I133551,I133383,I133582,I133599,I133395,I133639,I133404,I133661,I864449,I133678,I864452,I133704,I133721,I133407,I133743,I133392,I133774,I864446,I133791,I133808,I133825,I133401,I133856,I133389,I133398,I133386,I133942,I956056,I133968,I133976,I133993,I956074,I956068,I134010,I956047,I134036,I956065,I134053,I134061,I956050,I134078,I133910,I134109,I134126,I133922,I956062,I134166,I133931,I134188,I956071,I956059,I134205,I956053,I134231,I134248,I133934,I134270,I133919,I134301,I134318,I134335,I134352,I133928,I134383,I133916,I133925,I133913,I134469,I1112708,I134495,I134503,I134520,I1112723,I1112702,I134537,I1112705,I134563,I1112726,I134580,I134588,I134605,I134437,I134636,I134653,I134449,I134693,I134458,I134715,I1112714,I1112711,I134732,I1112717,I134758,I134775,I134461,I134797,I134446,I134828,I1112720,I134845,I134862,I134879,I134455,I134910,I134443,I134452,I134440,I134996,I549229,I135022,I135030,I135047,I549241,I549226,I135064,I549220,I135090,I549235,I135107,I135115,I549223,I135132,I134964,I135163,I135180,I134976,I549232,I135220,I134985,I135242,I549238,I549244,I135259,I135285,I135302,I134988,I135324,I134973,I135355,I135372,I135389,I135406,I134982,I135437,I134970,I134979,I134967,I135523,I365630,I135549,I135557,I135574,I365612,I365627,I135591,I365603,I135617,I365606,I135634,I135642,I365621,I135659,I135491,I135690,I135707,I135503,I365624,I135747,I135512,I135769,I365615,I135786,I365609,I135812,I135829,I135515,I135851,I135500,I135882,I365618,I135899,I135916,I135933,I135509,I135964,I135497,I135506,I135494,I136050,I605873,I136076,I136084,I136101,I605885,I605870,I136118,I605864,I136144,I605879,I136161,I136169,I605867,I136186,I136018,I136217,I136234,I136030,I605876,I136274,I136039,I136296,I605882,I605888,I136313,I136339,I136356,I136042,I136378,I136027,I136409,I136426,I136443,I136460,I136036,I136491,I136024,I136033,I136021,I136580,I460487,I136606,I136614,I460481,I136640,I136648,I460478,I136665,I460469,I136682,I136557,I136713,I460472,I136551,I136744,I460475,I136761,I136778,I460463,I460490,I136795,I136812,I136829,I136566,I136563,I136569,I136888,I136905,I136922,I460466,I136948,I136548,I136979,I136987,I460484,I136572,I137018,I137035,I137052,I136554,I137083,I137100,I136545,I136560,I137175,I197259,I137201,I137209,I197253,I137235,I137243,I197238,I137260,I197247,I137277,I137152,I137308,I197235,I137146,I137339,I197241,I137356,I137373,I197244,I197256,I137390,I137407,I137424,I137161,I137158,I137164,I137483,I137500,I137517,I197250,I137543,I137143,I137574,I137582,I137167,I137613,I137630,I137647,I137149,I137678,I137695,I137140,I137155,I137770,I526231,I137796,I137804,I526237,I137830,I137838,I526219,I137855,I526243,I137872,I137747,I137903,I526234,I137741,I137934,I526225,I137951,I137968,I526228,I526222,I137985,I138002,I138019,I137756,I137753,I137759,I138078,I138095,I138112,I526240,I138138,I137738,I138169,I138177,I137762,I138208,I138225,I138242,I137744,I138273,I138290,I137735,I137750,I138365,I601255,I138391,I138399,I601240,I138425,I138433,I601264,I138450,I601243,I138467,I138342,I138498,I601246,I138336,I138529,I601249,I138546,I138563,I601252,I601258,I138580,I138597,I138614,I138351,I138348,I138354,I138673,I138690,I138707,I601261,I138733,I138333,I138764,I138772,I138357,I138803,I138820,I138837,I138339,I138868,I138885,I138330,I138345,I138960,I279711,I138986,I138994,I279708,I139020,I139028,I279705,I139045,I279717,I139062,I138937,I139093,I279726,I138931,I139124,I279723,I139141,I139158,I279702,I139175,I139192,I139209,I138946,I138943,I138949,I139268,I139285,I139302,I279714,I279729,I139328,I138928,I139359,I139367,I279720,I138952,I139398,I139415,I139432,I138934,I139463,I139480,I138925,I138940,I139555,I489863,I139581,I139589,I489857,I139615,I139623,I489854,I139640,I489845,I139657,I139532,I139688,I489848,I139526,I139719,I489851,I139736,I139753,I489839,I489866,I139770,I139787,I139804,I139541,I139538,I139544,I139863,I139880,I139897,I489842,I139923,I139523,I139954,I139962,I489860,I139547,I139993,I140010,I140027,I139529,I140058,I140075,I139520,I139535,I140150,I140176,I140184,I140210,I140218,I140235,I140252,I140283,I140314,I140331,I140348,I140365,I140382,I140399,I140458,I140475,I140492,I140518,I140549,I140557,I140588,I140605,I140622,I140653,I140670,I140745,I140771,I140779,I140805,I140813,I140830,I140847,I140722,I140878,I140716,I140909,I140926,I140943,I140960,I140977,I140994,I140731,I140728,I140734,I141053,I141070,I141087,I141113,I140713,I141144,I141152,I140737,I141183,I141200,I141217,I140719,I141248,I141265,I140710,I140725,I141340,I449063,I141366,I141374,I449057,I141400,I141408,I449054,I141425,I449045,I141442,I141317,I141473,I449048,I141311,I141504,I449051,I141521,I141538,I449039,I449066,I141555,I141572,I141589,I141326,I141323,I141329,I141648,I141665,I141682,I449042,I141708,I141308,I141739,I141747,I449060,I141332,I141778,I141795,I141812,I141314,I141843,I141860,I141305,I141320,I141935,I1084383,I141961,I141969,I1084380,I141995,I142003,I1084389,I142020,I142037,I141912,I142068,I1084392,I141906,I142099,I1084386,I142116,I142133,I1084401,I142150,I142167,I142184,I141921,I141918,I141924,I142243,I142260,I142277,I1084404,I1084398,I142303,I141903,I142334,I142342,I1084395,I141927,I142373,I142390,I142407,I141909,I142438,I142455,I141900,I141915,I142530,I712216,I142556,I142564,I712237,I142590,I142598,I142615,I712228,I142632,I142507,I142663,I712225,I142501,I142694,I712234,I142711,I142728,I712219,I142745,I142762,I142779,I142516,I142513,I142519,I142838,I142855,I142872,I712240,I712222,I142898,I142498,I142929,I142937,I712231,I142522,I142968,I142985,I143002,I142504,I143033,I143050,I142495,I142510,I143125,I697188,I143151,I143159,I697209,I143185,I143193,I143210,I697200,I143227,I143258,I697197,I143289,I697206,I143306,I143323,I697191,I143340,I143357,I143374,I143433,I143450,I143467,I697212,I697194,I143493,I143524,I143532,I697203,I143563,I143580,I143597,I143628,I143645,I143720,I652104,I143746,I143754,I652125,I143780,I143788,I143805,I652116,I143822,I143853,I652113,I143884,I652122,I143901,I143918,I652107,I143935,I143952,I143969,I144028,I144045,I144062,I652128,I652110,I144088,I144119,I144127,I652119,I144158,I144175,I144192,I144223,I144240,I144315,I604723,I144341,I144349,I604708,I144375,I144383,I604732,I144400,I604711,I144417,I144448,I604714,I144479,I604717,I144496,I144513,I604720,I604726,I144530,I144547,I144564,I144623,I144640,I144657,I604729,I144683,I144714,I144722,I144753,I144770,I144787,I144818,I144835,I144910,I567731,I144936,I144944,I567716,I144970,I144978,I567740,I144995,I567719,I145012,I144887,I145043,I567722,I144881,I145074,I567725,I145091,I145108,I567728,I567734,I145125,I145142,I145159,I144896,I144893,I144899,I145218,I145235,I145252,I567737,I145278,I144878,I145309,I145317,I144902,I145348,I145365,I145382,I144884,I145413,I145430,I144875,I144890,I145505,I231769,I145531,I145539,I231763,I145565,I145573,I231748,I145590,I231757,I145607,I145482,I145638,I231745,I145476,I145669,I231751,I145686,I145703,I231754,I231766,I145720,I145737,I145754,I145491,I145488,I145494,I145813,I145830,I145847,I231760,I145873,I145473,I145904,I145912,I145497,I145943,I145960,I145977,I145479,I146008,I146025,I145470,I145485,I146100,I498266,I146126,I146134,I498272,I146160,I146168,I498254,I146185,I498278,I146202,I146077,I146233,I498269,I146071,I146264,I498260,I146281,I146298,I498263,I498257,I146315,I146332,I146349,I146086,I146083,I146089,I146408,I146425,I146442,I498275,I146468,I146068,I146499,I146507,I146092,I146538,I146555,I146572,I146074,I146603,I146620,I146065,I146080,I146695,I850738,I146721,I146729,I146755,I146763,I850735,I146780,I850747,I146797,I146672,I146828,I850741,I146666,I146859,I850753,I146876,I146893,I850744,I850732,I146910,I146927,I146944,I146681,I146678,I146684,I147003,I147020,I147037,I147063,I146663,I147094,I147102,I850750,I146687,I147133,I147150,I147167,I146669,I147198,I147215,I146660,I146675,I147290,I225224,I147316,I147324,I225218,I147350,I147358,I225203,I147375,I225212,I147392,I147267,I147423,I225200,I147261,I147454,I225206,I147471,I147488,I225209,I225221,I147505,I147522,I147539,I147276,I147273,I147279,I147598,I147615,I147632,I225215,I147658,I147258,I147689,I147697,I147282,I147728,I147745,I147762,I147264,I147793,I147810,I147255,I147270,I147885,I147911,I147919,I147945,I147953,I147970,I147987,I147862,I148018,I147856,I148049,I148066,I148083,I148100,I148117,I148134,I147871,I147868,I147874,I148193,I148210,I148227,I148253,I147853,I148284,I148292,I147877,I148323,I148340,I148357,I147859,I148388,I148405,I147850,I147865,I148477,I621485,I148503,I148520,I148542,I621476,I148568,I148576,I148593,I621494,I148610,I621491,I148627,I148644,I621470,I148661,I621473,I148678,I621482,I148695,I148726,I148743,I148760,I148777,I148822,I621488,I148867,I148884,I148901,I621479,I148918,I148944,I148952,I149006,I149014,I149072,I490951,I149098,I149115,I149064,I149137,I490939,I149163,I149171,I149188,I490948,I149205,I490945,I149222,I149239,I490936,I149256,I490942,I149273,I490927,I149290,I149040,I149321,I149338,I149355,I149372,I149052,I149046,I149417,I149061,I149055,I149462,I149479,I490933,I149496,I490930,I149513,I490954,I149539,I149547,I149049,I149043,I149601,I149609,I149058,I149667,I1134666,I149693,I149710,I149659,I149732,I149758,I149766,I149783,I1134669,I149800,I1134681,I149817,I149834,I1134687,I149851,I1134678,I149868,I1134684,I149885,I149635,I149916,I149933,I149950,I149967,I149647,I149641,I150012,I1134675,I149656,I149650,I150057,I150074,I1134672,I150091,I1134690,I150108,I150134,I150142,I149644,I149638,I150196,I150204,I149653,I150262,I510166,I150288,I150305,I150254,I150327,I510160,I150353,I150361,I150378,I510175,I150395,I510172,I150412,I150429,I510163,I150446,I510154,I150463,I510157,I150480,I150230,I150511,I150528,I150545,I150562,I150242,I150236,I150607,I510178,I150251,I150245,I150652,I150669,I510169,I150686,I150703,I150729,I150737,I150239,I150233,I150791,I150799,I150248,I150857,I335564,I150883,I150900,I150849,I150922,I335579,I150948,I150956,I150973,I335576,I150990,I151007,I151024,I335573,I151041,I335588,I151058,I335585,I151075,I150825,I151106,I151123,I151140,I151157,I150837,I150831,I151202,I335582,I150846,I150840,I151247,I151264,I335570,I151281,I335591,I151298,I335567,I151324,I151332,I150834,I150828,I151386,I151394,I150843,I151452,I786444,I151478,I151495,I151444,I151517,I786438,I151543,I151551,I151568,I786456,I151585,I151602,I151619,I151636,I786450,I151653,I786441,I151670,I151420,I151701,I151718,I151735,I151752,I151432,I151426,I151797,I786453,I151441,I151435,I151842,I151859,I786459,I151876,I151893,I786447,I151919,I151927,I151429,I151423,I151981,I151989,I151438,I152047,I890170,I152073,I152090,I152039,I152112,I890179,I152138,I152146,I152163,I890167,I152180,I890158,I152197,I152214,I890164,I152231,I890182,I152248,I890155,I152265,I152015,I152296,I152313,I152330,I152347,I152027,I152021,I152392,I890161,I152036,I152030,I152437,I152454,I890173,I152471,I152488,I890176,I152514,I152522,I152024,I152018,I152576,I152584,I152033,I152642,I1376733,I152668,I152685,I152707,I1376724,I152733,I152741,I152758,I1376718,I152775,I1376712,I152792,I152809,I1376739,I152826,I152843,I1376736,I152860,I152891,I152908,I152925,I152942,I152987,I1376721,I153032,I153049,I1376727,I153066,I1376730,I153083,I1376715,I153109,I153117,I153171,I153179,I153237,I323443,I153263,I153280,I153229,I153302,I323458,I153328,I153336,I153353,I323455,I153370,I153387,I153404,I323452,I153421,I323467,I153438,I323464,I153455,I153205,I153486,I153503,I153520,I153537,I153217,I153211,I153582,I323461,I153226,I153220,I153627,I153644,I323449,I153661,I323470,I153678,I323446,I153704,I153712,I153214,I153208,I153766,I153774,I153223,I153832,I935390,I153858,I153875,I153824,I153897,I935399,I153923,I153931,I153948,I935387,I153965,I935378,I153982,I153999,I935384,I154016,I935402,I154033,I935375,I154050,I153800,I154081,I154098,I154115,I154132,I153812,I153806,I154177,I935381,I153821,I153815,I154222,I154239,I935393,I154256,I154273,I935396,I154299,I154307,I153809,I153803,I154361,I154369,I153818,I154427,I1080334,I154453,I154470,I154419,I154492,I154518,I154526,I154543,I1080337,I154560,I1080349,I154577,I154594,I1080355,I154611,I1080346,I154628,I1080352,I154645,I154395,I154676,I154693,I154710,I154727,I154407,I154401,I154772,I1080343,I154416,I154410,I154817,I154834,I1080340,I154851,I1080358,I154868,I154894,I154902,I154404,I154398,I154956,I154964,I154413,I155022,I155048,I155065,I155014,I155087,I155113,I155121,I155138,I155155,I155172,I155189,I155206,I155223,I155240,I154990,I155271,I155288,I155305,I155322,I155002,I154996,I155367,I155011,I155005,I155412,I155429,I155446,I155463,I155489,I155497,I154999,I154993,I155551,I155559,I155008,I155617,I1071086,I155643,I155660,I155609,I155682,I155708,I155716,I155733,I1071089,I155750,I1071101,I155767,I155784,I1071107,I155801,I1071098,I155818,I1071104,I155835,I155585,I155866,I155883,I155900,I155917,I155597,I155591,I155962,I1071095,I155606,I155600,I156007,I156024,I1071092,I156041,I1071110,I156058,I156084,I156092,I155594,I155588,I156146,I156154,I155603,I156212,I1382088,I156238,I156255,I156204,I156277,I1382079,I156303,I156311,I156328,I1382073,I156345,I1382067,I156362,I156379,I1382094,I156396,I156413,I1382091,I156430,I156180,I156461,I156478,I156495,I156512,I156192,I156186,I156557,I1382076,I156201,I156195,I156602,I156619,I1382082,I156636,I1382085,I156653,I1382070,I156679,I156687,I156189,I156183,I156741,I156749,I156198,I156807,I392487,I156833,I156850,I156799,I156872,I392475,I156898,I156906,I156923,I392484,I156940,I392481,I156957,I156974,I392472,I156991,I392478,I157008,I392463,I157025,I156775,I157056,I157073,I157090,I157107,I156787,I156781,I157152,I156796,I156790,I157197,I157214,I392469,I157231,I392466,I157248,I392490,I157274,I157282,I156784,I156778,I157336,I157344,I156793,I157402,I1246612,I157428,I157445,I157394,I157467,I1246597,I157493,I157501,I157518,I1246615,I157535,I157552,I157569,I1246618,I157586,I1246609,I157603,I1246606,I157620,I157370,I157651,I157668,I157685,I157702,I157382,I157376,I157747,I1246603,I157391,I157385,I157792,I157809,I1246594,I157826,I1246600,I157843,I157869,I157877,I157379,I157373,I157931,I157939,I157388,I157997,I638822,I158023,I158040,I158062,I638819,I158088,I158096,I158113,I638825,I158130,I638810,I158147,I158164,I638813,I158181,I638834,I158198,I638831,I158215,I158246,I158263,I158280,I158297,I158342,I158387,I158404,I638816,I158421,I638828,I158438,I158464,I158472,I158526,I158534,I158592,I1149116,I158618,I158635,I158584,I158657,I158683,I158691,I158708,I1149119,I158725,I1149131,I158742,I158759,I1149137,I158776,I1149128,I158793,I1149134,I158810,I158560,I158841,I158858,I158875,I158892,I158572,I158566,I158937,I1149125,I158581,I158575,I158982,I158999,I1149122,I159016,I1149140,I159033,I159059,I159067,I158569,I158563,I159121,I159129,I158578,I159187,I1359478,I159213,I159230,I159179,I159252,I1359469,I159278,I159286,I159303,I1359463,I159320,I1359457,I159337,I159354,I1359484,I159371,I159388,I1359481,I159405,I159155,I159436,I159453,I159470,I159487,I159167,I159161,I159532,I1359466,I159176,I159170,I159577,I159594,I1359472,I159611,I1359475,I159628,I1359460,I159654,I159662,I159164,I159158,I159716,I159724,I159173,I159782,I1129464,I159808,I159825,I159774,I159847,I159873,I159881,I159898,I1129467,I159915,I1129479,I159932,I159949,I1129485,I159966,I1129476,I159983,I1129482,I160000,I159750,I160031,I160048,I160065,I160082,I159762,I159756,I160127,I1129473,I159771,I159765,I160172,I160189,I1129470,I160206,I1129488,I160223,I160249,I160257,I159759,I159753,I160311,I160319,I159768,I160377,I1360073,I160403,I160420,I160369,I160442,I1360064,I160468,I160476,I160493,I1360058,I160510,I1360052,I160527,I160544,I1360079,I160561,I160578,I1360076,I160595,I160345,I160626,I160643,I160660,I160677,I160357,I160351,I160722,I1360061,I160366,I160360,I160767,I160784,I1360067,I160801,I1360070,I160818,I1360055,I160844,I160852,I160354,I160348,I160906,I160914,I160363,I160972,I160998,I161015,I160964,I161037,I161063,I161071,I161088,I161105,I161122,I161139,I161156,I161173,I161190,I160940,I161221,I161238,I161255,I161272,I160952,I160946,I161317,I160961,I160955,I161362,I161379,I161396,I161413,I161439,I161447,I160949,I160943,I161501,I161509,I160958,I161567,I161593,I161610,I161559,I161632,I161658,I161666,I161683,I161700,I161717,I161734,I161751,I161768,I161785,I161535,I161816,I161833,I161850,I161867,I161547,I161541,I161912,I161556,I161550,I161957,I161974,I161991,I162008,I162034,I162042,I161544,I161538,I162096,I162104,I161553,I162162,I642290,I162188,I162205,I162154,I162227,I642287,I162253,I162261,I162278,I642293,I162295,I642278,I162312,I162329,I642281,I162346,I642302,I162363,I642299,I162380,I162130,I162411,I162428,I162445,I162462,I162142,I162136,I162507,I162151,I162145,I162552,I162569,I642284,I162586,I642296,I162603,I162629,I162637,I162139,I162133,I162691,I162699,I162148,I162757,I1313663,I162783,I162800,I162749,I162822,I1313654,I162848,I162856,I162873,I1313648,I162890,I1313642,I162907,I162924,I1313669,I162941,I162958,I1313666,I162975,I162725,I163006,I163023,I163040,I163057,I162737,I162731,I163102,I1313651,I162746,I162740,I163147,I163164,I1313657,I163181,I1313660,I163198,I1313645,I163224,I163232,I162734,I162728,I163286,I163294,I162743,I163352,I686218,I163378,I163395,I163344,I163417,I686215,I163443,I163451,I163468,I686221,I163485,I686206,I163502,I163519,I686209,I163536,I686230,I163553,I686227,I163570,I163320,I163601,I163618,I163635,I163652,I163332,I163326,I163697,I163341,I163335,I163742,I163759,I686212,I163776,I686224,I163793,I163819,I163827,I163329,I163323,I163881,I163889,I163338,I163947,I1395178,I163973,I163990,I163939,I164012,I1395169,I164038,I164046,I164063,I1395163,I164080,I1395157,I164097,I164114,I1395184,I164131,I164148,I1395181,I164165,I163915,I164196,I164213,I164230,I164247,I163927,I163921,I164292,I1395166,I163936,I163930,I164337,I164354,I1395172,I164371,I1395175,I164388,I1395160,I164414,I164422,I163924,I163918,I164476,I164484,I163933,I164542,I620329,I164568,I164585,I164534,I164607,I620320,I164633,I164641,I164658,I620338,I164675,I620335,I164692,I164709,I620314,I164726,I620317,I164743,I620326,I164760,I164510,I164791,I164808,I164825,I164842,I164522,I164516,I164887,I620332,I164531,I164525,I164932,I164949,I164966,I620323,I164983,I165009,I165017,I164519,I164513,I165071,I165079,I164528,I165137,I346104,I165163,I165180,I165129,I165202,I346119,I165228,I165236,I165253,I346116,I165270,I165287,I165304,I346113,I165321,I346128,I165338,I346125,I165355,I165105,I165386,I165403,I165420,I165437,I165117,I165111,I165482,I346122,I165126,I165120,I165527,I165544,I346110,I165561,I346131,I165578,I346107,I165604,I165612,I165114,I165108,I165666,I165674,I165123,I165732,I1395773,I165758,I165775,I165724,I165797,I1395764,I165823,I165831,I165848,I1395758,I165865,I1395752,I165882,I165899,I1395779,I165916,I165933,I1395776,I165950,I165700,I165981,I165998,I166015,I166032,I165712,I165706,I166077,I1395761,I165721,I165715,I166122,I166139,I1395767,I166156,I1395770,I166173,I1395755,I166199,I166207,I165709,I165703,I166261,I166269,I165718,I166327,I166353,I166370,I166319,I166392,I166418,I166426,I166443,I166460,I166477,I166494,I166511,I166528,I166545,I166295,I166576,I166593,I166610,I166627,I166307,I166301,I166672,I166316,I166310,I166717,I166734,I166751,I166768,I166794,I166802,I166304,I166298,I166856,I166864,I166313,I166922,I643446,I166948,I166965,I166914,I166987,I643443,I167013,I167021,I167038,I643449,I167055,I643434,I167072,I167089,I643437,I167106,I643458,I167123,I643455,I167140,I166890,I167171,I167188,I167205,I167222,I166902,I166896,I167267,I166911,I166905,I167312,I167329,I643440,I167346,I643452,I167363,I167389,I167397,I166899,I166893,I167451,I167459,I166908,I167517,I388135,I167543,I167560,I167509,I167582,I388123,I167608,I167616,I167633,I388132,I167650,I388129,I167667,I167684,I388120,I167701,I388126,I167718,I388111,I167735,I167485,I167766,I167783,I167800,I167817,I167497,I167491,I167862,I167506,I167500,I167907,I167924,I388117,I167941,I388114,I167958,I388138,I167984,I167992,I167494,I167488,I168046,I168054,I167503,I168112,I1190732,I168138,I168155,I168177,I168203,I168211,I168228,I1190735,I168245,I1190747,I168262,I168279,I1190753,I168296,I1190744,I168313,I1190750,I168330,I168361,I168378,I168395,I168412,I168457,I1190741,I168502,I168519,I1190738,I168536,I1190756,I168553,I168579,I168587,I168641,I168649,I168707,I257041,I168733,I168750,I168699,I168772,I257056,I168798,I168806,I168823,I257053,I168840,I168857,I168874,I257050,I168891,I257065,I168908,I257062,I168925,I168675,I168956,I168973,I168990,I169007,I168687,I168681,I169052,I257059,I168696,I168690,I169097,I169114,I257047,I169131,I257068,I169148,I257044,I169174,I169182,I168684,I168678,I169236,I169244,I168693,I169302,I430023,I169328,I169345,I169294,I169367,I430011,I169393,I169401,I169418,I430020,I169435,I430017,I169452,I169469,I430008,I169486,I430014,I169503,I429999,I169520,I169270,I169551,I169568,I169585,I169602,I169282,I169276,I169647,I169291,I169285,I169692,I169709,I430005,I169726,I430002,I169743,I430026,I169769,I169777,I169279,I169273,I169831,I169839,I169288,I169897,I847576,I169923,I169940,I169889,I169962,I847570,I169988,I169996,I170013,I847588,I170030,I170047,I170064,I170081,I847582,I170098,I847573,I170115,I169865,I170146,I170163,I170180,I170197,I169877,I169871,I170242,I847585,I169886,I169880,I170287,I170304,I847591,I170321,I170338,I847579,I170364,I170372,I169874,I169868,I170426,I170434,I169883,I170492,I170518,I170535,I170484,I170557,I170583,I170591,I170608,I170625,I170642,I170659,I170676,I170693,I170710,I170460,I170741,I170758,I170775,I170792,I170472,I170466,I170837,I170481,I170475,I170882,I170899,I170916,I170933,I170959,I170967,I170469,I170463,I171021,I171029,I170478,I171087,I171113,I171130,I171079,I171152,I171178,I171186,I171203,I171220,I171237,I171254,I171271,I171288,I171305,I171055,I171336,I171353,I171370,I171387,I171067,I171061,I171432,I171076,I171070,I171477,I171494,I171511,I171528,I171554,I171562,I171064,I171058,I171616,I171624,I171073,I171682,I660786,I171708,I171725,I171674,I171747,I660783,I171773,I171781,I171798,I660789,I171815,I660774,I171832,I171849,I660777,I171866,I660798,I171883,I660795,I171900,I171650,I171931,I171948,I171965,I171982,I171662,I171656,I172027,I171671,I171665,I172072,I172089,I660780,I172106,I660792,I172123,I172149,I172157,I171659,I171653,I172211,I172219,I171668,I172277,I1272097,I172303,I172320,I172269,I172342,I1272109,I172368,I172376,I172393,I1272103,I172410,I1272115,I172427,I172444,I1272100,I172461,I1272112,I172478,I1272094,I172495,I172245,I172526,I172543,I172560,I172577,I172257,I172251,I172622,I1272106,I172266,I172260,I172667,I172684,I172701,I172718,I1272118,I172744,I172752,I172254,I172248,I172806,I172814,I172263,I172872,I1073398,I172898,I172915,I172864,I172937,I172963,I172971,I172988,I1073401,I173005,I1073413,I173022,I173039,I1073419,I173056,I1073410,I173073,I1073416,I173090,I172840,I173121,I173138,I173155,I173172,I172852,I172846,I173217,I1073407,I172861,I172855,I173262,I173279,I1073404,I173296,I1073422,I173313,I173339,I173347,I172849,I172843,I173401,I173409,I172858,I173467,I444711,I173493,I173510,I173459,I173532,I444699,I173558,I173566,I173583,I444708,I173600,I444705,I173617,I173634,I444696,I173651,I444702,I173668,I444687,I173685,I173435,I173716,I173733,I173750,I173767,I173447,I173441,I173812,I173456,I173450,I173857,I173874,I444693,I173891,I444690,I173908,I444714,I173934,I173942,I173444,I173438,I173996,I174004,I173453,I174062,I1012949,I174088,I174105,I174054,I174127,I1012958,I174153,I174161,I174178,I1012952,I174195,I1012946,I174212,I174229,I1012961,I174246,I174263,I1012955,I174280,I174030,I174311,I174328,I174345,I174362,I174042,I174036,I174407,I174051,I174045,I174452,I174469,I1012967,I174486,I1012964,I174503,I174529,I174537,I174039,I174033,I174591,I174599,I174048,I174657,I575245,I174683,I174700,I174649,I174722,I575236,I174748,I174756,I174773,I575254,I174790,I575251,I174807,I174824,I575230,I174841,I575233,I174858,I575242,I174875,I174625,I174906,I174923,I174940,I174957,I174637,I174631,I175002,I575248,I174646,I174640,I175047,I175064,I175081,I575239,I175098,I175124,I175132,I174634,I174628,I175186,I175194,I174643,I175252,I521471,I175278,I175295,I175244,I175317,I521465,I175343,I175351,I175368,I521480,I175385,I521477,I175402,I175419,I521468,I175436,I521459,I175453,I521462,I175470,I175220,I175501,I175518,I175535,I175552,I175232,I175226,I175597,I521483,I175241,I175235,I175642,I175659,I521474,I175676,I175693,I175719,I175727,I175229,I175223,I175781,I175789,I175238,I175847,I607035,I175873,I175890,I175839,I175912,I607026,I175938,I175946,I175963,I607044,I175980,I607041,I175997,I176014,I607020,I176031,I607023,I176048,I607032,I176065,I175815,I176096,I176113,I176130,I176147,I175827,I175821,I176192,I607038,I175836,I175830,I176237,I176254,I176271,I607029,I176288,I176314,I176322,I175824,I175818,I176376,I176384,I175833,I176442,I1314853,I176468,I176485,I176434,I176507,I1314844,I176533,I176541,I176558,I1314838,I176575,I1314832,I176592,I176609,I1314859,I176626,I176643,I1314856,I176660,I176410,I176691,I176708,I176725,I176742,I176422,I176416,I176787,I1314841,I176431,I176425,I176832,I176849,I1314847,I176866,I1314850,I176883,I1314835,I176909,I176917,I176419,I176413,I176971,I176979,I176428,I177037,I519686,I177063,I177080,I177029,I177102,I519680,I177128,I177136,I177153,I519695,I177170,I519692,I177187,I177204,I519683,I177221,I519674,I177238,I519677,I177255,I177005,I177286,I177303,I177320,I177337,I177017,I177011,I177382,I519698,I177026,I177020,I177427,I177444,I519689,I177461,I177478,I177504,I177512,I177014,I177008,I177566,I177574,I177023,I177632,I687952,I177658,I177675,I177624,I177697,I687949,I177723,I177731,I177748,I687955,I177765,I687940,I177782,I177799,I687943,I177816,I687964,I177833,I687961,I177850,I177600,I177881,I177898,I177915,I177932,I177612,I177606,I177977,I177621,I177615,I178022,I178039,I687946,I178056,I687958,I178073,I178099,I178107,I177609,I177603,I178161,I178169,I177618,I178227,I1051658,I178253,I178270,I178219,I178292,I1051667,I178318,I178326,I178343,I1051661,I178360,I1051655,I178377,I178394,I1051670,I178411,I178428,I1051664,I178445,I178195,I178476,I178493,I178510,I178527,I178207,I178201,I178572,I178216,I178210,I178617,I178634,I1051676,I178651,I1051673,I178668,I178694,I178702,I178204,I178198,I178756,I178764,I178213,I178822,I976734,I178848,I178865,I178814,I178887,I976743,I178913,I178921,I178938,I976731,I178955,I976722,I178972,I178989,I976728,I179006,I976746,I179023,I976719,I179040,I178790,I179071,I179088,I179105,I179122,I178802,I178796,I179167,I976725,I178811,I178805,I179212,I179229,I976737,I179246,I179263,I976740,I179289,I179297,I178799,I178793,I179351,I179359,I178808,I179417,I842833,I179443,I179460,I179409,I179482,I842827,I179508,I179516,I179533,I842845,I179550,I179567,I179584,I179601,I842839,I179618,I842830,I179635,I179385,I179666,I179683,I179700,I179717,I179397,I179391,I179762,I842842,I179406,I179400,I179807,I179824,I842848,I179841,I179858,I842836,I179884,I179892,I179394,I179388,I179946,I179954,I179403,I180012,I180038,I180055,I180004,I180077,I180103,I180111,I180128,I180145,I180162,I180179,I180196,I180213,I180230,I179980,I180261,I180278,I180295,I180312,I179992,I179986,I180357,I180001,I179995,I180402,I180419,I180436,I180453,I180479,I180487,I179989,I179983,I180541,I180549,I179998,I180607,I686796,I180633,I180650,I180599,I180672,I686793,I180698,I180706,I180723,I686799,I180740,I686784,I180757,I180774,I686787,I180791,I686808,I180808,I686805,I180825,I180575,I180856,I180873,I180890,I180907,I180587,I180581,I180952,I180596,I180590,I180997,I181014,I686790,I181031,I686802,I181048,I181074,I181082,I180584,I180578,I181136,I181144,I180593,I181202,I414791,I181228,I181245,I181194,I181267,I414779,I181293,I181301,I181318,I414788,I181335,I414785,I181352,I181369,I414776,I181386,I414782,I181403,I414767,I181420,I181170,I181451,I181468,I181485,I181502,I181182,I181176,I181547,I181191,I181185,I181592,I181609,I414773,I181626,I414770,I181643,I414794,I181669,I181677,I181179,I181173,I181731,I181739,I181188,I181797,I310268,I181823,I181840,I181862,I310283,I181888,I181896,I181913,I310280,I181930,I181947,I181964,I310277,I181981,I310292,I181998,I310289,I182015,I182046,I182063,I182080,I182097,I182142,I310286,I182187,I182204,I310274,I182221,I310295,I182238,I310271,I182264,I182272,I182326,I182334,I182392,I1121950,I182418,I182435,I182384,I182457,I182483,I182491,I182508,I1121953,I182525,I1121965,I182542,I182559,I1121971,I182576,I1121962,I182593,I1121968,I182610,I182360,I182641,I182658,I182675,I182692,I182372,I182366,I182737,I1121959,I182381,I182375,I182782,I182799,I1121956,I182816,I1121974,I182833,I182859,I182867,I182369,I182363,I182921,I182929,I182378,I182987,I668878,I183013,I183030,I182979,I183052,I668875,I183078,I183086,I183103,I668881,I183120,I668866,I183137,I183154,I668869,I183171,I668890,I183188,I668887,I183205,I182955,I183236,I183253,I183270,I183287,I182967,I182961,I183332,I182976,I182970,I183377,I183394,I668872,I183411,I668884,I183428,I183454,I183462,I182964,I182958,I183516,I183524,I182973,I183582,I1168768,I183608,I183625,I183574,I183647,I183673,I183681,I183698,I1168771,I183715,I1168783,I183732,I183749,I1168789,I183766,I1168780,I183783,I1168786,I183800,I183550,I183831,I183848,I183865,I183882,I183562,I183556,I183927,I1168777,I183571,I183565,I183972,I183989,I1168774,I184006,I1168792,I184023,I184049,I184057,I183559,I183553,I184111,I184119,I183568,I184177,I184203,I184220,I184169,I184242,I184268,I184276,I184293,I184310,I184327,I184344,I184361,I184378,I184395,I184145,I184426,I184443,I184460,I184477,I184157,I184151,I184522,I184166,I184160,I184567,I184584,I184601,I184618,I184644,I184652,I184154,I184148,I184706,I184714,I184163,I184772,I280229,I184798,I184815,I184837,I280244,I184863,I184871,I184888,I280241,I184905,I184922,I184939,I280238,I184956,I280253,I184973,I280250,I184990,I185021,I185038,I185055,I185072,I185117,I280247,I185162,I185179,I280235,I185196,I280256,I185213,I280232,I185239,I185247,I185301,I185309,I185367,I185393,I185410,I185359,I185432,I185458,I185466,I185483,I185500,I185517,I185534,I185551,I185568,I185585,I185335,I185616,I185633,I185650,I185667,I185347,I185341,I185712,I185356,I185350,I185757,I185774,I185791,I185808,I185834,I185842,I185344,I185338,I185896,I185904,I185353,I185962,I316065,I185988,I186005,I185954,I186027,I316080,I186053,I186061,I186078,I316077,I186095,I186112,I186129,I316074,I186146,I316089,I186163,I316086,I186180,I185930,I186211,I186228,I186245,I186262,I185942,I185936,I186307,I316083,I185951,I185945,I186352,I186369,I316071,I186386,I316092,I186403,I316068,I186429,I186437,I185939,I185933,I186491,I186499,I185948,I186557,I1301446,I186583,I186600,I186549,I186622,I1301419,I186648,I186656,I186673,I1301443,I186690,I1301440,I186707,I186724,I186741,I1301437,I186758,I1301425,I186775,I186525,I186806,I186823,I186840,I186857,I186537,I186531,I186902,I1301431,I186546,I186540,I186947,I186964,I1301434,I186981,I1301422,I186998,I1301428,I187024,I187032,I186534,I186528,I187086,I187094,I186543,I187152,I1321398,I187178,I187195,I187144,I187217,I1321389,I187243,I187251,I187268,I1321383,I187285,I1321377,I187302,I187319,I1321404,I187336,I187353,I1321401,I187370,I187120,I187401,I187418,I187435,I187452,I187132,I187126,I187497,I1321386,I187141,I187135,I187542,I187559,I1321392,I187576,I1321395,I187593,I1321380,I187619,I187627,I187129,I187123,I187681,I187689,I187138,I187747,I1065306,I187773,I187790,I187739,I187812,I187838,I187846,I187863,I1065309,I187880,I1065321,I187897,I187914,I1065327,I187931,I1065318,I187948,I1065324,I187965,I187715,I187996,I188013,I188030,I188047,I187727,I187721,I188092,I1065315,I187736,I187730,I188137,I188154,I1065312,I188171,I1065330,I188188,I188214,I188222,I187724,I187718,I188276,I188284,I187733,I188342,I188368,I188385,I188407,I188433,I188441,I188458,I188475,I188492,I188509,I188526,I188543,I188560,I188591,I188608,I188625,I188642,I188687,I188732,I188749,I188766,I188783,I188809,I188817,I188871,I188879,I188937,I1043804,I188963,I188980,I188929,I189002,I1043813,I189028,I189036,I189053,I1043807,I189070,I1043801,I189087,I189104,I1043816,I189121,I189138,I1043810,I189155,I188905,I189186,I189203,I189220,I189237,I188917,I188911,I189282,I188926,I188920,I189327,I189344,I1043822,I189361,I1043819,I189378,I189404,I189412,I188914,I188908,I189466,I189474,I188923,I189532,I590273,I189558,I189575,I189524,I189597,I590264,I189623,I189631,I189648,I590282,I189665,I590279,I189682,I189699,I590258,I189716,I590261,I189733,I590270,I189750,I189500,I189781,I189798,I189815,I189832,I189512,I189506,I189877,I590276,I189521,I189515,I189922,I189939,I189956,I590267,I189973,I189999,I190007,I189509,I189503,I190061,I190069,I189518,I190127,I796457,I190153,I190170,I190119,I190192,I796451,I190218,I190226,I190243,I796469,I190260,I190277,I190294,I190311,I796463,I190328,I796454,I190345,I190095,I190376,I190393,I190410,I190427,I190107,I190101,I190472,I796466,I190116,I190110,I190517,I190534,I796472,I190551,I190568,I796460,I190594,I190602,I190104,I190098,I190656,I190664,I190113,I190722,I1155474,I190748,I190765,I190714,I190787,I190813,I190821,I190838,I1155477,I190855,I1155489,I190872,I190889,I1155495,I190906,I1155486,I190923,I1155492,I190940,I190690,I190971,I190988,I191005,I191022,I190702,I190696,I191067,I1155483,I190711,I190705,I191112,I191129,I1155480,I191146,I1155498,I191163,I191189,I191197,I190699,I190693,I191251,I191259,I190708,I191317,I366130,I191343,I191360,I191382,I366145,I191408,I191416,I191433,I366142,I191450,I191467,I191484,I366139,I191501,I366154,I191518,I366151,I191535,I191566,I191583,I191600,I191617,I191662,I366148,I191707,I191724,I366136,I191741,I366157,I191758,I366133,I191784,I191792,I191846,I191854,I191912,I258095,I191938,I191955,I191904,I191977,I258110,I192003,I192011,I192028,I258107,I192045,I192062,I192079,I258104,I192096,I258119,I192113,I258116,I192130,I191880,I192161,I192178,I192195,I192212,I191892,I191886,I192257,I258113,I191901,I191895,I192302,I192319,I258101,I192336,I258122,I192353,I258098,I192379,I192387,I191889,I191883,I192441,I192449,I191898,I192507,I524446,I192533,I192550,I192499,I192572,I524440,I192598,I192606,I192623,I524455,I192640,I524452,I192657,I192674,I524443,I192691,I524434,I192708,I524437,I192725,I192475,I192756,I192773,I192790,I192807,I192487,I192481,I192852,I524458,I192496,I192490,I192897,I192914,I524449,I192931,I192948,I192974,I192982,I192484,I192478,I193036,I193044,I192493,I193102,I844941,I193128,I193145,I193094,I193167,I844935,I193193,I193201,I193218,I844953,I193235,I193252,I193269,I193286,I844947,I193303,I844938,I193320,I193070,I193351,I193368,I193385,I193402,I193082,I193076,I193447,I844950,I193091,I193085,I193492,I193509,I844956,I193526,I193543,I844944,I193569,I193577,I193079,I193073,I193631,I193639,I193088,I193697,I670612,I193723,I193740,I193689,I193762,I670609,I193788,I193796,I193813,I670615,I193830,I670600,I193847,I193864,I670603,I193881,I670624,I193898,I670621,I193915,I193665,I193946,I193963,I193980,I193997,I193677,I193671,I194042,I193686,I193680,I194087,I194104,I670606,I194121,I670618,I194138,I194164,I194172,I193674,I193668,I194226,I194234,I193683,I194292,I1342818,I194318,I194335,I194284,I194357,I1342809,I194383,I194391,I194408,I1342803,I194425,I1342797,I194442,I194459,I1342824,I194476,I194493,I1342821,I194510,I194260,I194541,I194558,I194575,I194592,I194272,I194266,I194637,I1342806,I194281,I194275,I194682,I194699,I1342812,I194716,I1342815,I194733,I1342800,I194759,I194767,I194269,I194263,I194821,I194829,I194278,I194887,I1184374,I194913,I194930,I194879,I194952,I194978,I194986,I195003,I1184377,I195020,I1184389,I195037,I195054,I1184395,I195071,I1184386,I195088,I1184392,I195105,I194855,I195136,I195153,I195170,I195187,I194867,I194861,I195232,I1184383,I194876,I194870,I195277,I195294,I1184380,I195311,I1184398,I195328,I195354,I195362,I194864,I194858,I195416,I195424,I194873,I195482,I574667,I195508,I195525,I195474,I195547,I574658,I195573,I195581,I195598,I574676,I195615,I574673,I195632,I195649,I574652,I195666,I574655,I195683,I574664,I195700,I195450,I195731,I195748,I195765,I195782,I195462,I195456,I195827,I574670,I195471,I195465,I195872,I195889,I195906,I574661,I195923,I195949,I195957,I195459,I195453,I196011,I196019,I195468,I196077,I874980,I196103,I196120,I196069,I196142,I874974,I196168,I196176,I196193,I874992,I196210,I196227,I196244,I196261,I874986,I196278,I874977,I196295,I196045,I196326,I196343,I196360,I196377,I196057,I196051,I196422,I874989,I196066,I196060,I196467,I196484,I874995,I196501,I196518,I874983,I196544,I196552,I196054,I196048,I196606,I196614,I196063,I196672,I545189,I196698,I196715,I196737,I545180,I196763,I196771,I196788,I545198,I196805,I545195,I196822,I196839,I545174,I196856,I545177,I196873,I545186,I196890,I196921,I196938,I196955,I196972,I197017,I545192,I197062,I197079,I197096,I545183,I197113,I197139,I197147,I197201,I197209,I197267,I308160,I197293,I197310,I197332,I308175,I197358,I197366,I197383,I308172,I197400,I197417,I197434,I308169,I197451,I308184,I197468,I308181,I197485,I197516,I197533,I197550,I197567,I197612,I308178,I197657,I197674,I308166,I197691,I308187,I197708,I308163,I197734,I197742,I197796,I197804,I197862,I992238,I197888,I197905,I197854,I197927,I992247,I197953,I197961,I197978,I992235,I197995,I992226,I198012,I198029,I992232,I198046,I992250,I198063,I992223,I198080,I197830,I198111,I198128,I198145,I198162,I197842,I197836,I198207,I992229,I197851,I197845,I198252,I198269,I992241,I198286,I198303,I992244,I198329,I198337,I197839,I197833,I198391,I198399,I197848,I198457,I634776,I198483,I198500,I198449,I198522,I634773,I198548,I198556,I198573,I634779,I198590,I634764,I198607,I198624,I634767,I198641,I634788,I198658,I634785,I198675,I198425,I198706,I198723,I198740,I198757,I198437,I198431,I198802,I198446,I198440,I198847,I198864,I634770,I198881,I634782,I198898,I198924,I198932,I198434,I198428,I198986,I198994,I198443,I199052,I1273831,I199078,I199095,I199044,I199117,I1273843,I199143,I199151,I199168,I1273837,I199185,I1273849,I199202,I199219,I1273834,I199236,I1273846,I199253,I1273828,I199270,I199020,I199301,I199318,I199335,I199352,I199032,I199026,I199397,I1273840,I199041,I199035,I199442,I199459,I199476,I199493,I1273852,I199519,I199527,I199029,I199023,I199581,I199589,I199038,I199647,I1258803,I199673,I199690,I199639,I199712,I1258815,I199738,I199746,I199763,I1258809,I199780,I1258821,I199797,I199814,I1258806,I199831,I1258818,I199848,I1258800,I199865,I199615,I199896,I199913,I199930,I199947,I199627,I199621,I199992,I1258812,I199636,I199630,I200037,I200054,I200071,I200088,I1258824,I200114,I200122,I199624,I199618,I200176,I200184,I199633,I200242,I1312473,I200268,I200285,I200234,I200307,I1312464,I200333,I200341,I200358,I1312458,I200375,I1312452,I200392,I200409,I1312479,I200426,I200443,I1312476,I200460,I200210,I200491,I200508,I200525,I200542,I200222,I200216,I200587,I1312461,I200231,I200225,I200632,I200649,I1312467,I200666,I1312470,I200683,I1312455,I200709,I200717,I200219,I200213,I200771,I200779,I200228,I200837,I372981,I200863,I200880,I200829,I200902,I372996,I200928,I200936,I200953,I372993,I200970,I200987,I201004,I372990,I201021,I373005,I201038,I373002,I201055,I200805,I201086,I201103,I201120,I201137,I200817,I200811,I201182,I372999,I200826,I200820,I201227,I201244,I372987,I201261,I373008,I201278,I372984,I201304,I201312,I200814,I200808,I201366,I201374,I200823,I201432,I525041,I201458,I201475,I201424,I201497,I525035,I201523,I201531,I201548,I525050,I201565,I525047,I201582,I201599,I525038,I201616,I525029,I201633,I525032,I201650,I201400,I201681,I201698,I201715,I201732,I201412,I201406,I201777,I525053,I201421,I201415,I201822,I201839,I525044,I201856,I201873,I201899,I201907,I201409,I201403,I201961,I201969,I201418,I202027,I1161832,I202053,I202070,I202019,I202092,I202118,I202126,I202143,I1161835,I202160,I1161847,I202177,I202194,I1161853,I202211,I1161844,I202228,I1161850,I202245,I201995,I202276,I202293,I202310,I202327,I202007,I202001,I202372,I1161841,I202016,I202010,I202417,I202434,I1161838,I202451,I1161856,I202468,I202494,I202502,I202004,I201998,I202556,I202564,I202013,I202622,I829131,I202648,I202665,I202614,I202687,I829125,I202713,I202721,I202738,I829143,I202755,I202772,I202789,I202806,I829137,I202823,I829128,I202840,I202590,I202871,I202888,I202905,I202922,I202602,I202596,I202967,I829140,I202611,I202605,I203012,I203029,I829146,I203046,I203063,I829134,I203089,I203097,I202599,I202593,I203151,I203159,I202608,I203217,I1375543,I203243,I203260,I203209,I203282,I1375534,I203308,I203316,I203333,I1375528,I203350,I1375522,I203367,I203384,I1375549,I203401,I203418,I1375546,I203435,I203185,I203466,I203483,I203500,I203517,I203197,I203191,I203562,I1375531,I203206,I203200,I203607,I203624,I1375537,I203641,I1375540,I203658,I1375525,I203684,I203692,I203194,I203188,I203746,I203754,I203203,I203812,I483335,I203838,I203855,I203804,I203877,I483323,I203903,I203911,I203928,I483332,I203945,I483329,I203962,I203979,I483320,I203996,I483326,I204013,I483311,I204030,I203780,I204061,I204078,I204095,I204112,I203792,I203786,I204157,I203801,I203795,I204202,I204219,I483317,I204236,I483314,I204253,I483338,I204279,I204287,I203789,I203783,I204341,I204349,I203798,I204407,I838090,I204433,I204450,I204399,I204472,I838084,I204498,I204506,I204523,I838102,I204540,I204557,I204574,I204591,I838096,I204608,I838087,I204625,I204375,I204656,I204673,I204690,I204707,I204387,I204381,I204752,I838099,I204396,I204390,I204797,I204814,I838105,I204831,I204848,I838093,I204874,I204882,I204384,I204378,I204936,I204944,I204393,I205002,I608769,I205028,I205045,I204994,I205067,I608760,I205093,I205101,I205118,I608778,I205135,I608775,I205152,I205169,I608754,I205186,I608757,I205203,I608766,I205220,I204970,I205251,I205268,I205285,I205302,I204982,I204976,I205347,I608772,I204991,I204985,I205392,I205409,I205426,I608763,I205443,I205469,I205477,I204979,I204973,I205531,I205539,I204988,I205597,I1300324,I205623,I205640,I205662,I1300297,I205688,I205696,I205713,I1300321,I205730,I1300318,I205747,I205764,I205781,I1300315,I205798,I1300303,I205815,I205846,I205863,I205880,I205897,I205942,I1300309,I205987,I206004,I1300312,I206021,I1300300,I206038,I1300306,I206064,I206072,I206126,I206134,I206192,I866548,I206218,I206235,I206184,I206257,I866542,I206283,I206291,I206308,I866560,I206325,I206342,I206359,I206376,I866554,I206393,I866545,I206410,I206160,I206441,I206458,I206475,I206492,I206172,I206166,I206537,I866557,I206181,I206175,I206582,I206599,I866563,I206616,I206633,I866551,I206659,I206667,I206169,I206163,I206721,I206729,I206178,I206787,I562529,I206813,I206830,I206779,I206852,I562520,I206878,I206886,I206903,I562538,I206920,I562535,I206937,I206954,I562514,I206971,I562517,I206988,I562526,I207005,I206755,I207036,I207053,I207070,I207087,I206767,I206761,I207132,I562532,I206776,I206770,I207177,I207194,I207211,I562523,I207228,I207254,I207262,I206764,I206758,I207316,I207324,I206773,I207382,I1352933,I207408,I207425,I207374,I207447,I1352924,I207473,I207481,I207498,I1352918,I207515,I1352912,I207532,I207549,I1352939,I207566,I207583,I1352936,I207600,I207350,I207631,I207648,I207665,I207682,I207362,I207356,I207727,I1352921,I207371,I207365,I207772,I207789,I1352927,I207806,I1352930,I207823,I1352915,I207849,I207857,I207359,I207353,I207911,I207919,I207368,I207977,I1267473,I208003,I208020,I207969,I208042,I1267485,I208068,I208076,I208093,I1267479,I208110,I1267491,I208127,I208144,I1267476,I208161,I1267488,I208178,I1267470,I208195,I207945,I208226,I208243,I208260,I208277,I207957,I207951,I208322,I1267482,I207966,I207960,I208367,I208384,I208401,I208418,I1267494,I208444,I208452,I207954,I207948,I208506,I208514,I207963,I208572,I1269785,I208598,I208615,I208637,I1269797,I208663,I208671,I208688,I1269791,I208705,I1269803,I208722,I208739,I1269788,I208756,I1269800,I208773,I1269782,I208790,I208821,I208838,I208855,I208872,I208917,I1269794,I208962,I208979,I208996,I209013,I1269806,I209039,I209047,I209101,I209109,I209167,I874453,I209193,I209210,I209159,I209232,I874447,I209258,I209266,I209283,I874465,I209300,I209317,I209334,I209351,I874459,I209368,I874450,I209385,I209135,I209416,I209433,I209450,I209467,I209147,I209141,I209512,I874462,I209156,I209150,I209557,I209574,I874468,I209591,I209608,I874456,I209634,I209642,I209144,I209138,I209696,I209704,I209153,I209762,I548657,I209788,I209805,I209827,I548648,I209853,I209861,I209878,I548666,I209895,I548663,I209912,I209929,I548642,I209946,I548645,I209963,I548654,I209980,I210011,I210028,I210045,I210062,I210107,I548660,I210152,I210169,I210186,I548651,I210203,I210229,I210237,I210291,I210299,I210357,I1114436,I210383,I210400,I210349,I210422,I210448,I210456,I210473,I1114439,I210490,I1114451,I210507,I210524,I1114457,I210541,I1114448,I210558,I1114454,I210575,I210325,I210606,I210623,I210640,I210657,I210337,I210331,I210702,I1114445,I210346,I210340,I210747,I210764,I1114442,I210781,I1114460,I210798,I210824,I210832,I210334,I210328,I210886,I210894,I210343,I210952,I1086692,I210978,I210995,I210944,I211017,I211043,I211051,I211068,I1086695,I211085,I1086707,I211102,I211119,I1086713,I211136,I1086704,I211153,I1086710,I211170,I210920,I211201,I211218,I211235,I211252,I210932,I210926,I211297,I1086701,I210941,I210935,I211342,I211359,I1086698,I211376,I1086716,I211393,I211419,I211427,I210929,I210923,I211481,I211489,I210938,I211547,I648648,I211573,I211590,I211539,I211612,I648645,I211638,I211646,I211663,I648651,I211680,I648636,I211697,I211714,I648639,I211731,I648660,I211748,I648657,I211765,I211515,I211796,I211813,I211830,I211847,I211527,I211521,I211892,I211536,I211530,I211937,I211954,I648642,I211971,I648654,I211988,I212014,I212022,I211524,I211518,I212076,I212084,I211533,I212142,I447431,I212168,I212185,I212134,I212207,I447419,I212233,I212241,I212258,I447428,I212275,I447425,I212292,I212309,I447416,I212326,I447422,I212343,I447407,I212360,I212110,I212391,I212408,I212425,I212442,I212122,I212116,I212487,I212131,I212125,I212532,I212549,I447413,I212566,I447410,I212583,I447434,I212609,I212617,I212119,I212113,I212671,I212679,I212128,I212737,I886294,I212763,I212780,I212729,I212802,I886303,I212828,I212836,I212853,I886291,I212870,I886282,I212887,I212904,I886288,I212921,I886306,I212938,I886279,I212955,I212705,I212986,I213003,I213020,I213037,I212717,I212711,I213082,I886285,I212726,I212720,I213127,I213144,I886297,I213161,I213178,I886300,I213204,I213212,I212714,I212708,I213266,I213274,I212723,I213332,I213358,I213375,I213324,I213397,I213423,I213431,I213448,I213465,I213482,I213499,I213516,I213533,I213550,I213300,I213581,I213598,I213615,I213632,I213312,I213306,I213677,I213321,I213315,I213722,I213739,I213756,I213773,I213799,I213807,I213309,I213303,I213861,I213869,I213318,I213927,I1334488,I213953,I213970,I213919,I213992,I1334479,I214018,I214026,I214043,I1334473,I214060,I1334467,I214077,I214094,I1334494,I214111,I214128,I1334491,I214145,I213895,I214176,I214193,I214210,I214227,I213907,I213901,I214272,I1334476,I213916,I213910,I214317,I214334,I1334482,I214351,I1334485,I214368,I1334470,I214394,I214402,I213904,I213898,I214456,I214464,I213913,I214522,I522066,I214548,I214565,I214514,I214587,I522060,I214613,I214621,I214638,I522075,I214655,I522072,I214672,I214689,I522063,I214706,I522054,I214723,I522057,I214740,I214490,I214771,I214788,I214805,I214822,I214502,I214496,I214867,I522078,I214511,I214505,I214912,I214929,I522069,I214946,I214963,I214989,I214997,I214499,I214493,I215051,I215059,I214508,I215117,I215143,I215160,I215109,I215182,I215208,I215216,I215233,I215250,I215267,I215284,I215301,I215318,I215335,I215085,I215366,I215383,I215400,I215417,I215097,I215091,I215462,I215106,I215100,I215507,I215524,I215541,I215558,I215584,I215592,I215094,I215088,I215646,I215654,I215103,I215712,I1044926,I215738,I215755,I215704,I215777,I1044935,I215803,I215811,I215828,I1044929,I215845,I1044923,I215862,I215879,I1044938,I215896,I215913,I1044932,I215930,I215680,I215961,I215978,I215995,I216012,I215692,I215686,I216057,I215701,I215695,I216102,I216119,I1044944,I216136,I1044941,I216153,I216179,I216187,I215689,I215683,I216241,I216249,I215698,I216307,I696044,I216333,I216350,I216299,I216372,I696041,I216398,I216406,I216423,I696047,I216440,I696032,I216457,I216474,I696035,I216491,I696056,I216508,I696053,I216525,I216275,I216556,I216573,I216590,I216607,I216287,I216281,I216652,I216296,I216290,I216697,I216714,I696038,I216731,I696050,I216748,I216774,I216782,I216284,I216278,I216836,I216844,I216293,I216902,I1198824,I216928,I216945,I216894,I216967,I216993,I217001,I217018,I1198827,I217035,I1198839,I217052,I217069,I1198845,I217086,I1198836,I217103,I1198842,I217120,I216870,I217151,I217168,I217185,I217202,I216882,I216876,I217247,I1198833,I216891,I216885,I217292,I217309,I1198830,I217326,I1198848,I217343,I217369,I217377,I216879,I216873,I217431,I217439,I216888,I217497,I217523,I217540,I217562,I217588,I217596,I217613,I217630,I217647,I217664,I217681,I217698,I217715,I217746,I217763,I217780,I217797,I217842,I217887,I217904,I217921,I217938,I217964,I217972,I218026,I218034,I218092,I852319,I218118,I218135,I218084,I218157,I852313,I218183,I218191,I218208,I852331,I218225,I218242,I218259,I218276,I852325,I218293,I852316,I218310,I218060,I218341,I218358,I218375,I218392,I218072,I218066,I218437,I852328,I218081,I218075,I218482,I218499,I852334,I218516,I218533,I852322,I218559,I218567,I218069,I218063,I218621,I218629,I218078,I218687,I1209620,I218713,I218730,I218679,I218752,I1209605,I218778,I218786,I218803,I1209623,I218820,I218837,I218854,I1209626,I218871,I1209617,I218888,I1209614,I218905,I218655,I218936,I218953,I218970,I218987,I218667,I218661,I219032,I1209611,I218676,I218670,I219077,I219094,I1209602,I219111,I1209608,I219128,I219154,I219162,I218664,I218658,I219216,I219224,I218673,I219282,I760780,I219308,I219325,I219347,I760777,I219373,I219381,I219398,I760783,I219415,I760768,I219432,I219449,I760771,I219466,I760792,I219483,I760789,I219500,I219531,I219548,I219565,I219582,I219627,I219672,I219689,I760774,I219706,I760786,I219723,I219749,I219757,I219811,I219819,I219877,I488231,I219903,I219920,I219869,I219942,I488219,I219968,I219976,I219993,I488228,I220010,I488225,I220027,I220044,I488216,I220061,I488222,I220078,I488207,I220095,I219845,I220126,I220143,I220160,I220177,I219857,I219851,I220222,I219866,I219860,I220267,I220284,I488213,I220301,I488210,I220318,I488234,I220344,I220352,I219854,I219848,I220406,I220414,I219863,I220472,I1262849,I220498,I220515,I220464,I220537,I1262861,I220563,I220571,I220588,I1262855,I220605,I1262867,I220622,I220639,I1262852,I220656,I1262864,I220673,I1262846,I220690,I220440,I220721,I220738,I220755,I220772,I220452,I220446,I220817,I1262858,I220461,I220455,I220862,I220879,I220896,I220913,I1262870,I220939,I220947,I220449,I220443,I221001,I221009,I220458,I221067,I1160676,I221093,I221110,I221059,I221132,I221158,I221166,I221183,I1160679,I221200,I1160691,I221217,I221234,I1160697,I221251,I1160688,I221268,I1160694,I221285,I221035,I221316,I221333,I221350,I221367,I221047,I221041,I221412,I1160685,I221056,I221050,I221457,I221474,I1160682,I221491,I1160700,I221508,I221534,I221542,I221044,I221038,I221596,I221604,I221053,I221662,I723788,I221688,I221705,I221654,I221727,I723785,I221753,I221761,I221778,I723791,I221795,I723776,I221812,I221829,I723779,I221846,I723800,I221863,I723797,I221880,I221630,I221911,I221928,I221945,I221962,I221642,I221636,I222007,I221651,I221645,I222052,I222069,I723782,I222086,I723794,I222103,I222129,I222137,I221639,I221633,I222191,I222199,I221648,I222257,I871818,I222283,I222300,I222249,I222322,I871812,I222348,I222356,I222373,I871830,I222390,I222407,I222424,I222441,I871824,I222458,I871815,I222475,I222225,I222506,I222523,I222540,I222557,I222237,I222231,I222602,I871827,I222246,I222240,I222647,I222664,I871833,I222681,I222698,I871821,I222724,I222732,I222234,I222228,I222786,I222794,I222243,I222852,I470823,I222878,I222895,I222844,I222917,I470811,I222943,I222951,I222968,I470820,I222985,I470817,I223002,I223019,I470808,I223036,I470814,I223053,I470799,I223070,I222820,I223101,I223118,I223135,I223152,I222832,I222826,I223197,I222841,I222835,I223242,I223259,I470805,I223276,I470802,I223293,I470826,I223319,I223327,I222829,I222823,I223381,I223389,I222838,I223447,I1088426,I223473,I223490,I223512,I223538,I223546,I223563,I1088429,I223580,I1088441,I223597,I223614,I1088447,I223631,I1088438,I223648,I1088444,I223665,I223696,I223713,I223730,I223747,I223792,I1088435,I223837,I223854,I1088432,I223871,I1088450,I223888,I223914,I223922,I223976,I223984,I224042,I850211,I224068,I224085,I224107,I850205,I224133,I224141,I224158,I850223,I224175,I224192,I224209,I224226,I850217,I224243,I850208,I224260,I224291,I224308,I224325,I224342,I224387,I850220,I224432,I224449,I850226,I224466,I224483,I850214,I224509,I224517,I224571,I224579,I224637,I785390,I224663,I224680,I224629,I224702,I785384,I224728,I224736,I224753,I785402,I224770,I224787,I224804,I224821,I785396,I224838,I785387,I224855,I224605,I224886,I224903,I224920,I224937,I224617,I224611,I224982,I785399,I224626,I224620,I225027,I225044,I785405,I225061,I225078,I785393,I225104,I225112,I224614,I224608,I225166,I225174,I224623,I225232,I361914,I225258,I225275,I225297,I361929,I225323,I225331,I225348,I361926,I225365,I225382,I225399,I361923,I225416,I361938,I225433,I361935,I225450,I225481,I225498,I225515,I225532,I225577,I361932,I225622,I225639,I361920,I225656,I361941,I225673,I361917,I225699,I225707,I225761,I225769,I225827,I1058948,I225853,I225870,I225819,I225892,I225918,I225926,I225943,I1058951,I225960,I1058963,I225977,I225994,I1058969,I226011,I1058960,I226028,I1058966,I226045,I225795,I226076,I226093,I226110,I226127,I225807,I225801,I226172,I1058957,I225816,I225810,I226217,I226234,I1058954,I226251,I1058972,I226268,I226294,I226302,I225804,I225798,I226356,I226364,I225813,I226422,I381607,I226448,I226465,I226414,I226487,I381595,I226513,I226521,I226538,I381604,I226555,I381601,I226572,I226589,I381592,I226606,I381598,I226623,I381583,I226640,I226390,I226671,I226688,I226705,I226722,I226402,I226396,I226767,I226411,I226405,I226812,I226829,I381589,I226846,I381586,I226863,I381610,I226889,I226897,I226399,I226393,I226951,I226959,I226408,I227017,I628418,I227043,I227060,I227009,I227082,I628415,I227108,I227116,I227133,I628421,I227150,I628406,I227167,I227184,I628409,I227201,I628430,I227218,I628427,I227235,I226985,I227266,I227283,I227300,I227317,I226997,I226991,I227362,I227006,I227000,I227407,I227424,I628412,I227441,I628424,I227458,I227484,I227492,I226994,I226988,I227546,I227554,I227003,I227612,I1319613,I227638,I227655,I227604,I227677,I1319604,I227703,I227711,I227728,I1319598,I227745,I1319592,I227762,I227779,I1319619,I227796,I227813,I1319616,I227830,I227580,I227861,I227878,I227895,I227912,I227592,I227586,I227957,I1319601,I227601,I227595,I228002,I228019,I1319607,I228036,I1319610,I228053,I1319595,I228079,I228087,I227589,I227583,I228141,I228149,I227598,I228207,I541106,I228233,I228250,I228199,I228272,I541100,I228298,I228306,I228323,I541115,I228340,I541112,I228357,I228374,I541103,I228391,I541094,I228408,I541097,I228425,I228175,I228456,I228473,I228490,I228507,I228187,I228181,I228552,I541118,I228196,I228190,I228597,I228614,I541109,I228631,I228648,I228674,I228682,I228184,I228178,I228736,I228744,I228193,I228802,I715696,I228828,I228845,I228794,I228867,I715693,I228893,I228901,I228918,I715699,I228935,I715684,I228952,I228969,I715687,I228986,I715708,I229003,I715705,I229020,I228770,I229051,I229068,I229085,I229102,I228782,I228776,I229147,I228791,I228785,I229192,I229209,I715690,I229226,I715702,I229243,I229269,I229277,I228779,I228773,I229331,I229339,I228788,I229397,I917302,I229423,I229440,I229389,I229462,I917311,I229488,I229496,I229513,I917299,I229530,I917290,I229547,I229564,I917296,I229581,I917314,I229598,I917287,I229615,I229365,I229646,I229663,I229680,I229697,I229377,I229371,I229742,I917293,I229386,I229380,I229787,I229804,I917305,I229821,I229838,I917308,I229864,I229872,I229374,I229368,I229926,I229934,I229383,I229992,I919240,I230018,I230035,I229984,I230057,I919249,I230083,I230091,I230108,I919237,I230125,I919228,I230142,I230159,I919234,I230176,I919252,I230193,I919225,I230210,I229960,I230241,I230258,I230275,I230292,I229972,I229966,I230337,I919231,I229981,I229975,I230382,I230399,I919243,I230416,I230433,I919246,I230459,I230467,I229969,I229963,I230521,I230529,I229978,I230587,I1222676,I230613,I230630,I230579,I230652,I1222661,I230678,I230686,I230703,I1222679,I230720,I230737,I230754,I1222682,I230771,I1222673,I230788,I1222670,I230805,I230555,I230836,I230853,I230870,I230887,I230567,I230561,I230932,I1222667,I230576,I230570,I230977,I230994,I1222658,I231011,I1222664,I231028,I231054,I231062,I230564,I230558,I231116,I231124,I230573,I231182,I903736,I231208,I231225,I231174,I231247,I903745,I231273,I231281,I231298,I903733,I231315,I903724,I231332,I231349,I903730,I231366,I903748,I231383,I903721,I231400,I231150,I231431,I231448,I231465,I231482,I231162,I231156,I231527,I903727,I231171,I231165,I231572,I231589,I903739,I231606,I231623,I903742,I231649,I231657,I231159,I231153,I231711,I231719,I231168,I231777,I596631,I231803,I231820,I231842,I596622,I231868,I231876,I231893,I596640,I231910,I596637,I231927,I231944,I596616,I231961,I596619,I231978,I596628,I231995,I232026,I232043,I232060,I232077,I232122,I596634,I232167,I232184,I232201,I596625,I232218,I232244,I232252,I232306,I232314,I232372,I1266895,I232398,I232415,I232364,I232437,I1266907,I232463,I232471,I232488,I1266901,I232505,I1266913,I232522,I232539,I1266898,I232556,I1266910,I232573,I1266892,I232590,I232340,I232621,I232638,I232655,I232672,I232352,I232346,I232717,I1266904,I232361,I232355,I232762,I232779,I232796,I232813,I1266916,I232839,I232847,I232349,I232343,I232901,I232909,I232358,I232967,I1383278,I232993,I233010,I232959,I233032,I1383269,I233058,I233066,I233083,I1383263,I233100,I1383257,I233117,I233134,I1383284,I233151,I233168,I1383281,I233185,I232935,I233216,I233233,I233250,I233267,I232947,I232941,I233312,I1383266,I232956,I232950,I233357,I233374,I1383272,I233391,I1383275,I233408,I1383260,I233434,I233442,I232944,I232938,I233496,I233504,I232953,I233562,I358752,I233588,I233605,I233554,I233627,I358767,I233653,I233661,I233678,I358764,I233695,I233712,I233729,I358761,I233746,I358776,I233763,I358773,I233780,I233530,I233811,I233828,I233845,I233862,I233542,I233536,I233907,I358770,I233551,I233545,I233952,I233969,I358758,I233986,I358779,I234003,I358755,I234029,I234037,I233539,I233533,I234091,I234099,I233548,I234157,I624953,I234183,I234200,I234149,I234222,I624944,I234248,I234256,I234273,I624962,I234290,I624959,I234307,I234324,I624938,I234341,I624941,I234358,I624950,I234375,I234125,I234406,I234423,I234440,I234457,I234137,I234131,I234502,I624956,I234146,I234140,I234547,I234564,I234581,I624947,I234598,I234624,I234632,I234134,I234128,I234686,I234694,I234143,I234752,I461575,I234778,I234795,I234744,I234817,I461563,I234843,I234851,I234868,I461572,I234885,I461569,I234902,I234919,I461560,I234936,I461566,I234953,I461551,I234970,I234720,I235001,I235018,I235035,I235052,I234732,I234726,I235097,I234741,I234735,I235142,I235159,I461557,I235176,I461554,I235193,I461578,I235219,I235227,I234729,I234723,I235281,I235289,I234738,I235347,I487687,I235373,I235390,I235412,I487675,I235438,I235446,I235463,I487684,I235480,I487681,I235497,I235514,I487672,I235531,I487678,I235548,I487663,I235565,I235596,I235613,I235630,I235647,I235692,I235737,I235754,I487669,I235771,I487666,I235788,I487690,I235814,I235822,I235876,I235884,I235942,I378343,I235968,I235985,I236007,I378331,I236033,I236041,I236058,I378340,I236075,I378337,I236092,I236109,I378328,I236126,I378334,I236143,I378319,I236160,I236191,I236208,I236225,I236242,I236287,I236332,I236349,I378325,I236366,I378322,I236383,I378346,I236409,I236417,I236471,I236479,I236537,I974150,I236563,I236580,I236602,I974159,I236628,I236636,I236653,I974147,I236670,I974138,I236687,I236704,I974144,I236721,I974162,I236738,I974135,I236755,I236786,I236803,I236820,I236837,I236882,I974141,I236927,I236944,I974153,I236961,I236978,I974156,I237004,I237012,I237066,I237074,I237132,I1074554,I237158,I237175,I237124,I237197,I237223,I237231,I237248,I1074557,I237265,I1074569,I237282,I237299,I1074575,I237316,I1074566,I237333,I1074572,I237350,I237100,I237381,I237398,I237415,I237432,I237112,I237106,I237477,I1074563,I237121,I237115,I237522,I237539,I1074560,I237556,I1074578,I237573,I237599,I237607,I237109,I237103,I237661,I237669,I237118,I237727,I937974,I237753,I237770,I237719,I237792,I937983,I237818,I237826,I237843,I937971,I237860,I937962,I237877,I237894,I937968,I237911,I937986,I237928,I937959,I237945,I237695,I237976,I237993,I238010,I238027,I237707,I237701,I238072,I937965,I237716,I237710,I238117,I238134,I937977,I238151,I238168,I937980,I238194,I238202,I237704,I237698,I238256,I238264,I237713,I238322,I266527,I238348,I238365,I238314,I238387,I266542,I238413,I238421,I238438,I266539,I238455,I238472,I238489,I266536,I238506,I266551,I238523,I266548,I238540,I238290,I238571,I238588,I238605,I238622,I238302,I238296,I238667,I266545,I238311,I238305,I238712,I238729,I266533,I238746,I266554,I238763,I266530,I238789,I238797,I238299,I238293,I238851,I238859,I238308,I238917,I493671,I238943,I238960,I238909,I238982,I493659,I239008,I239016,I239033,I493668,I239050,I493665,I239067,I239084,I493656,I239101,I493662,I239118,I493647,I239135,I238885,I239166,I239183,I239200,I239217,I238897,I238891,I239262,I238906,I238900,I239307,I239324,I493653,I239341,I493650,I239358,I493674,I239384,I239392,I238894,I238888,I239446,I239454,I238903,I239512,I239538,I239555,I239504,I239577,I239603,I239611,I239628,I239645,I239662,I239679,I239696,I239713,I239730,I239480,I239761,I239778,I239795,I239812,I239492,I239486,I239857,I239501,I239495,I239902,I239919,I239936,I239953,I239979,I239987,I239489,I239483,I240041,I240049,I239498,I240107,I1290593,I240133,I240150,I240099,I240172,I1290605,I240198,I240206,I240223,I1290599,I240240,I1290611,I240257,I240274,I1290596,I240291,I1290608,I240308,I1290590,I240325,I240075,I240356,I240373,I240390,I240407,I240087,I240081,I240452,I1290602,I240096,I240090,I240497,I240514,I240531,I240548,I1290614,I240574,I240582,I240084,I240078,I240636,I240644,I240093,I240702,I894692,I240728,I240745,I240694,I240767,I894701,I240793,I240801,I240818,I894689,I240835,I894680,I240852,I240869,I894686,I240886,I894704,I240903,I894677,I240920,I240670,I240951,I240968,I240985,I241002,I240682,I240676,I241047,I894683,I240691,I240685,I241092,I241109,I894695,I241126,I241143,I894698,I241169,I241177,I240679,I240673,I241231,I241239,I240688,I241297,I241323,I241340,I241289,I241362,I241388,I241396,I241413,I241430,I241447,I241464,I241481,I241498,I241515,I241265,I241546,I241563,I241580,I241597,I241277,I241271,I241642,I241286,I241280,I241687,I241704,I241721,I241738,I241764,I241772,I241274,I241268,I241826,I241834,I241283,I241892,I241918,I241935,I241884,I241957,I241983,I241991,I242008,I242025,I242042,I242059,I242076,I242093,I242110,I241860,I242141,I242158,I242175,I242192,I241872,I241866,I242237,I241881,I241875,I242282,I242299,I242316,I242333,I242359,I242367,I241869,I241863,I242421,I242429,I241878,I242487,I331875,I242513,I242530,I242479,I242552,I331890,I242578,I242586,I242603,I331887,I242620,I242637,I242654,I331884,I242671,I331899,I242688,I331896,I242705,I242455,I242736,I242753,I242770,I242787,I242467,I242461,I242832,I331893,I242476,I242470,I242877,I242894,I331881,I242911,I331902,I242928,I331878,I242954,I242962,I242464,I242458,I243016,I243024,I242473,I243082,I243108,I243125,I243074,I243147,I243173,I243181,I243198,I243215,I243232,I243249,I243266,I243283,I243300,I243050,I243331,I243348,I243365,I243382,I243062,I243056,I243427,I243071,I243065,I243472,I243489,I243506,I243523,I243549,I243557,I243059,I243053,I243611,I243619,I243068,I243677,I901152,I243703,I243720,I243669,I243742,I901161,I243768,I243776,I243793,I901149,I243810,I901140,I243827,I243844,I901146,I243861,I901164,I243878,I901137,I243895,I243645,I243926,I243943,I243960,I243977,I243657,I243651,I244022,I901143,I243666,I243660,I244067,I244084,I901155,I244101,I244118,I901158,I244144,I244152,I243654,I243648,I244206,I244214,I243663,I244272,I1351148,I244298,I244315,I244264,I244337,I1351139,I244363,I244371,I244388,I1351133,I244405,I1351127,I244422,I244439,I1351154,I244456,I244473,I1351151,I244490,I244240,I244521,I244538,I244555,I244572,I244252,I244246,I244617,I1351136,I244261,I244255,I244662,I244679,I1351142,I244696,I1351145,I244713,I1351130,I244739,I244747,I244249,I244243,I244801,I244809,I244258,I244867,I482247,I244893,I244910,I244859,I244932,I482235,I244958,I244966,I244983,I482244,I245000,I482241,I245017,I245034,I482232,I245051,I482238,I245068,I482223,I245085,I244835,I245116,I245133,I245150,I245167,I244847,I244841,I245212,I244856,I244850,I245257,I245274,I482229,I245291,I482226,I245308,I482250,I245334,I245342,I244844,I244838,I245396,I245404,I244853,I245462,I419143,I245488,I245505,I245454,I245527,I419131,I245553,I245561,I245578,I419140,I245595,I419137,I245612,I245629,I419128,I245646,I419134,I245663,I419119,I245680,I245430,I245711,I245728,I245745,I245762,I245442,I245436,I245807,I245451,I245445,I245852,I245869,I419125,I245886,I419122,I245903,I419146,I245929,I245937,I245439,I245433,I245991,I245999,I245448,I246057,I246083,I246100,I246122,I246148,I246156,I246173,I246190,I246207,I246224,I246241,I246258,I246275,I246306,I246323,I246340,I246357,I246402,I246447,I246464,I246481,I246498,I246524,I246532,I246586,I246594,I246652,I303944,I246678,I246695,I246644,I246717,I303959,I246743,I246751,I246768,I303956,I246785,I246802,I246819,I303953,I246836,I303968,I246853,I303965,I246870,I246620,I246901,I246918,I246935,I246952,I246632,I246626,I246997,I303962,I246641,I246635,I247042,I247059,I303950,I247076,I303971,I247093,I303947,I247119,I247127,I246629,I246623,I247181,I247189,I246638,I247247,I247273,I247290,I247239,I247312,I247338,I247346,I247363,I247380,I247397,I247414,I247431,I247448,I247465,I247215,I247496,I247513,I247530,I247547,I247227,I247221,I247592,I247236,I247230,I247637,I247654,I247671,I247688,I247714,I247722,I247224,I247218,I247776,I247784,I247233,I247842,I264946,I247868,I247885,I247834,I247907,I264961,I247933,I247941,I247958,I264958,I247975,I247992,I248009,I264955,I248026,I264970,I248043,I264967,I248060,I247810,I248091,I248108,I248125,I248142,I247822,I247816,I248187,I264964,I247831,I247825,I248232,I248249,I264952,I248266,I264973,I248283,I264949,I248309,I248317,I247819,I247813,I248371,I248379,I247828,I248437,I1349958,I248463,I248480,I248429,I248502,I1349949,I248528,I248536,I248553,I1349943,I248570,I1349937,I248587,I248604,I1349964,I248621,I248638,I1349961,I248655,I248405,I248686,I248703,I248720,I248737,I248417,I248411,I248782,I1349946,I248426,I248420,I248827,I248844,I1349952,I248861,I1349955,I248878,I1349940,I248904,I248912,I248414,I248408,I248966,I248974,I248423,I249032,I464295,I249058,I249075,I249024,I249097,I464283,I249123,I249131,I249148,I464292,I249165,I464289,I249182,I249199,I464280,I249216,I464286,I249233,I464271,I249250,I249000,I249281,I249298,I249315,I249332,I249012,I249006,I249377,I249021,I249015,I249422,I249439,I464277,I249456,I464274,I249473,I464298,I249499,I249507,I249009,I249003,I249561,I249569,I249018,I249627,I1186686,I249653,I249670,I249619,I249692,I249718,I249726,I249743,I1186689,I249760,I1186701,I249777,I249794,I1186707,I249811,I1186698,I249828,I1186704,I249845,I249595,I249876,I249893,I249910,I249927,I249607,I249601,I249972,I1186695,I249616,I249610,I250017,I250034,I1186692,I250051,I1186710,I250068,I250094,I250102,I249604,I249598,I250156,I250164,I249613,I250225,I1320208,I250251,I250259,I1320187,I250276,I1320214,I250302,I250193,I250324,I1320202,I250350,I250358,I1320205,I250375,I250401,I250217,I250423,I250199,I1320196,I250463,I250480,I250488,I250505,I250202,I250536,I1320193,I1320190,I250553,I1320211,I250579,I250587,I250190,I250208,I250632,I1320199,I250649,I250211,I250196,I250205,I250214,I250752,I1244980,I250778,I250786,I1244962,I1244986,I250803,I1244977,I250829,I250720,I250851,I1244983,I250877,I250885,I1244971,I250902,I250928,I250744,I250950,I250726,I250990,I251007,I251015,I251032,I250729,I251063,I1244968,I1244965,I251080,I1244974,I251106,I251114,I250717,I250735,I251159,I251176,I250738,I250723,I250732,I250741,I251279,I805413,I251305,I251313,I805416,I805410,I251330,I805422,I251356,I251247,I251378,I805425,I251404,I251412,I251429,I251455,I251271,I251477,I251253,I805428,I251517,I251534,I251542,I251559,I251256,I251590,I805419,I251607,I251633,I251641,I251244,I251262,I251686,I805431,I251703,I251265,I251250,I251259,I251268,I251806,I251832,I251840,I251857,I251883,I251774,I251905,I251931,I251939,I251956,I251982,I251798,I252004,I251780,I252044,I252061,I252069,I252086,I251783,I252117,I252134,I252160,I252168,I251771,I251789,I252213,I252230,I251792,I251777,I251786,I251795,I252333,I851789,I252359,I252367,I851792,I851786,I252384,I851798,I252410,I252432,I851801,I252458,I252466,I252483,I252509,I252531,I851804,I252571,I252588,I252596,I252613,I252644,I851795,I252661,I252687,I252695,I252740,I851807,I252757,I252860,I252886,I252894,I252911,I252937,I252828,I252959,I252985,I252993,I253010,I253036,I252852,I253058,I252834,I253098,I253115,I253123,I253140,I252837,I253171,I253188,I253214,I253222,I252825,I252843,I253267,I253284,I252846,I252831,I252840,I252849,I253387,I584493,I253413,I253421,I584478,I584481,I253438,I584496,I253464,I253355,I253486,I584490,I253512,I253520,I253537,I253563,I253379,I253585,I253361,I584487,I253625,I253642,I253650,I253667,I253364,I253698,I584502,I253715,I584499,I253741,I253749,I253352,I253370,I253794,I584484,I253811,I253373,I253358,I253367,I253376,I253914,I1060682,I253940,I253948,I1060697,I253965,I1060700,I253991,I253882,I254013,I1060706,I254039,I254047,I1060688,I254064,I254090,I253906,I254112,I253888,I1060685,I254152,I254169,I254177,I254194,I253891,I254225,I1060691,I254242,I1060703,I254268,I254276,I253879,I253897,I254321,I1060694,I254338,I253900,I253885,I253894,I253903,I254441,I1341033,I254467,I254475,I1341012,I254492,I1341039,I254518,I254409,I254540,I1341027,I254566,I254574,I1341030,I254591,I254617,I254433,I254639,I254415,I1341021,I254679,I254696,I254704,I254721,I254418,I254752,I1341018,I1341015,I254769,I1341036,I254795,I254803,I254406,I254424,I254848,I1341024,I254865,I254427,I254412,I254421,I254430,I254968,I925042,I254994,I255002,I925039,I925057,I255019,I925048,I255045,I255067,I925063,I255093,I255101,I925045,I255118,I255144,I255166,I925051,I255206,I255223,I255231,I255248,I255279,I925066,I255296,I925054,I255322,I255330,I255375,I925060,I255392,I255495,I1082646,I255521,I255529,I1082661,I255546,I1082664,I255572,I255463,I255594,I1082670,I255620,I255628,I1082652,I255645,I255671,I255487,I255693,I255469,I1082649,I255733,I255750,I255758,I255775,I255472,I255806,I1082655,I255823,I1082667,I255849,I255857,I255460,I255478,I255902,I1082658,I255919,I255481,I255466,I255475,I255484,I256022,I1231380,I256048,I256056,I1231362,I1231386,I256073,I1231377,I256099,I255990,I256121,I1231383,I256147,I256155,I1231371,I256172,I256198,I256014,I256220,I255996,I256260,I256277,I256285,I256302,I255999,I256333,I1231368,I1231365,I256350,I1231374,I256376,I256384,I255987,I256005,I256429,I256446,I256008,I255993,I256002,I256011,I256549,I256575,I256583,I256600,I256626,I256517,I256648,I256674,I256682,I256699,I256725,I256541,I256747,I256523,I256787,I256804,I256812,I256829,I256526,I256860,I256877,I256903,I256911,I256514,I256532,I256956,I256973,I256535,I256520,I256529,I256538,I257076,I549813,I257102,I257110,I549798,I549801,I257127,I549816,I257153,I257175,I549810,I257201,I257209,I257226,I257252,I257274,I549807,I257314,I257331,I257339,I257356,I257387,I549822,I257404,I549819,I257430,I257438,I257483,I549804,I257500,I257603,I1321993,I257629,I257637,I1321972,I257654,I1321999,I257680,I257571,I257702,I1321987,I257728,I257736,I1321990,I257753,I257779,I257595,I257801,I257577,I1321981,I257841,I257858,I257866,I257883,I257580,I257914,I1321978,I1321975,I257931,I1321996,I257957,I257965,I257568,I257586,I258010,I1321984,I258027,I257589,I257574,I257583,I257592,I258130,I633042,I258156,I258164,I633033,I633048,I258181,I633054,I258207,I258229,I633039,I258255,I258263,I258280,I258306,I258328,I633036,I258368,I258385,I258393,I258410,I258441,I633030,I633045,I258458,I258484,I258492,I258537,I633051,I258554,I258657,I258683,I258691,I258708,I258734,I258625,I258756,I258782,I258790,I258807,I258833,I258649,I258855,I258631,I258895,I258912,I258920,I258937,I258634,I258968,I258985,I259011,I259019,I258622,I258640,I259064,I259081,I258643,I258628,I258637,I258646,I259184,I259210,I259218,I259235,I259261,I259152,I259283,I259309,I259317,I259334,I259360,I259176,I259382,I259158,I259422,I259439,I259447,I259464,I259161,I259495,I259512,I259538,I259546,I259149,I259167,I259591,I259608,I259170,I259155,I259164,I259173,I259711,I259737,I259745,I259762,I259788,I259679,I259810,I259836,I259844,I259861,I259887,I259703,I259909,I259685,I259949,I259966,I259974,I259991,I259688,I260022,I260039,I260065,I260073,I259676,I259694,I260118,I260135,I259697,I259682,I259691,I259700,I260238,I1295229,I260264,I260272,I1295226,I1295217,I260289,I1295214,I260315,I260206,I260337,I1295223,I260363,I260371,I1295232,I260388,I260414,I260230,I260436,I260212,I1295235,I260476,I260493,I260501,I260518,I260215,I260549,I1295220,I260566,I1295238,I260592,I260600,I260203,I260221,I260645,I260662,I260224,I260209,I260218,I260227,I260765,I260791,I260799,I260816,I260842,I260733,I260864,I260890,I260898,I260915,I260941,I260757,I260963,I260739,I261003,I261020,I261028,I261045,I260742,I261076,I261093,I261119,I261127,I260730,I260748,I261172,I261189,I260751,I260736,I260745,I260754,I261292,I705870,I261318,I261326,I705861,I705876,I261343,I705882,I261369,I261260,I261391,I705867,I261417,I261425,I261442,I261468,I261284,I261490,I261266,I705864,I261530,I261547,I261555,I261572,I261269,I261603,I705858,I705873,I261620,I261646,I261654,I261257,I261275,I261699,I705879,I261716,I261278,I261263,I261272,I261281,I261819,I972200,I261845,I261853,I972197,I972215,I261870,I972206,I261896,I261787,I261918,I972221,I261944,I261952,I972203,I261969,I261995,I261811,I262017,I261793,I972209,I262057,I262074,I262082,I262099,I261796,I262130,I972224,I262147,I972212,I262173,I262181,I261784,I261802,I262226,I972218,I262243,I261805,I261790,I261799,I261808,I262346,I512537,I262372,I262380,I512549,I262397,I512534,I262423,I262314,I262445,I512558,I262471,I262479,I512555,I262496,I262522,I262338,I262544,I262320,I512546,I262584,I262601,I262609,I262626,I262323,I262657,I512543,I262674,I512552,I262700,I262708,I262311,I262329,I262753,I512540,I262770,I262332,I262317,I262326,I262335,I262873,I674658,I262899,I262907,I674649,I674664,I262924,I674670,I262950,I262841,I262972,I674655,I262998,I263006,I263023,I263049,I262865,I263071,I262847,I674652,I263111,I263128,I263136,I263153,I262850,I263184,I674646,I674661,I263201,I263227,I263235,I262838,I262856,I263280,I674667,I263297,I262859,I262844,I262853,I262862,I263400,I965740,I263426,I263434,I965737,I965755,I263451,I965746,I263477,I263368,I263499,I965761,I263525,I263533,I965743,I263550,I263576,I263392,I263598,I263374,I965749,I263638,I263655,I263663,I263680,I263377,I263711,I965764,I263728,I965752,I263754,I263762,I263365,I263383,I263807,I965758,I263824,I263386,I263371,I263380,I263389,I263927,I704714,I263953,I263961,I704705,I704720,I263978,I704726,I264004,I263895,I264026,I704711,I264052,I264060,I264077,I264103,I263919,I264125,I263901,I704708,I264165,I264182,I264190,I264207,I263904,I264238,I704702,I704717,I264255,I264281,I264289,I263892,I263910,I264334,I704723,I264351,I263913,I263898,I263907,I263916,I264454,I912122,I264480,I264488,I912119,I912137,I264505,I912128,I264531,I264422,I264553,I912143,I264579,I264587,I912125,I264604,I264630,I264446,I264652,I264428,I912131,I264692,I264709,I264717,I264734,I264431,I264765,I912146,I264782,I912134,I264808,I264816,I264419,I264437,I264861,I912140,I264878,I264440,I264425,I264434,I264443,I264981,I597787,I265007,I265015,I597772,I597775,I265032,I597790,I265058,I265080,I597784,I265106,I265114,I265131,I265157,I265179,I597781,I265219,I265236,I265244,I265261,I265292,I597796,I265309,I597793,I265335,I265343,I265388,I597778,I265405,I265508,I925688,I265534,I265542,I925685,I925703,I265559,I925694,I265585,I265476,I265607,I925709,I265633,I265641,I925691,I265658,I265684,I265500,I265706,I265482,I925697,I265746,I265763,I265771,I265788,I265485,I265819,I925712,I265836,I925700,I265862,I265870,I265473,I265491,I265915,I925706,I265932,I265494,I265479,I265488,I265497,I266035,I1063572,I266061,I266069,I1063587,I266086,I1063590,I266112,I266003,I266134,I1063596,I266160,I266168,I1063578,I266185,I266211,I266027,I266233,I266009,I1063575,I266273,I266290,I266298,I266315,I266012,I266346,I1063581,I266363,I1063593,I266389,I266397,I266000,I266018,I266442,I1063584,I266459,I266021,I266006,I266015,I266024,I266562,I441435,I266588,I266596,I441447,I441426,I266613,I441450,I266639,I266661,I441441,I266687,I266695,I441423,I266712,I266738,I266760,I441438,I266800,I266817,I266825,I266842,I266873,I441429,I266890,I441432,I266916,I266924,I266969,I441444,I266986,I267089,I267115,I267123,I267140,I267166,I267057,I267188,I267214,I267222,I267239,I267265,I267081,I267287,I267063,I267327,I267344,I267352,I267369,I267066,I267400,I267417,I267443,I267451,I267054,I267072,I267496,I267513,I267075,I267060,I267069,I267078,I267616,I1011827,I267642,I267650,I1011824,I267667,I1011836,I267693,I267584,I267715,I267741,I267749,I1011842,I267766,I267792,I267608,I267814,I267590,I1011830,I267854,I267871,I267879,I267896,I267593,I267927,I1011839,I1011845,I267944,I267970,I267978,I267581,I267599,I268023,I1011833,I268040,I267602,I267587,I267596,I267605,I268143,I1119060,I268169,I268177,I1119075,I268194,I1119078,I268220,I268242,I1119084,I268268,I268276,I1119066,I268293,I268319,I268341,I1119063,I268381,I268398,I268406,I268423,I268454,I1119069,I268471,I1119081,I268497,I268505,I268550,I1119072,I268567,I268670,I378875,I268696,I268704,I378887,I378866,I268721,I378890,I268747,I268638,I268769,I378881,I268795,I268803,I378863,I268820,I268846,I268662,I268868,I268644,I378878,I268908,I268925,I268933,I268950,I268647,I268981,I378869,I268998,I378872,I269024,I269032,I268635,I268653,I269077,I378884,I269094,I268656,I268641,I268650,I268659,I269197,I499447,I269223,I269231,I499459,I269248,I499444,I269274,I269165,I269296,I499468,I269322,I269330,I499465,I269347,I269373,I269189,I269395,I269171,I499456,I269435,I269452,I269460,I269477,I269174,I269508,I499453,I269525,I499462,I269551,I269559,I269162,I269180,I269604,I499450,I269621,I269183,I269168,I269177,I269186,I269724,I603567,I269750,I269758,I603552,I603555,I269775,I603570,I269801,I269692,I269823,I603564,I269849,I269857,I269874,I269900,I269716,I269922,I269698,I603561,I269962,I269979,I269987,I270004,I269701,I270035,I603576,I270052,I603573,I270078,I270086,I269689,I269707,I270131,I603558,I270148,I269710,I269695,I269704,I269713,I270251,I761358,I270277,I270285,I761349,I761364,I270302,I761370,I270328,I270219,I270350,I761355,I270376,I270384,I270401,I270427,I270243,I270449,I270225,I761352,I270489,I270506,I270514,I270531,I270228,I270562,I761346,I761361,I270579,I270605,I270613,I270216,I270234,I270658,I761367,I270675,I270237,I270222,I270231,I270240,I270778,I270804,I270812,I270829,I270855,I270746,I270877,I270903,I270911,I270928,I270954,I270770,I270976,I270752,I271016,I271033,I271041,I271058,I270755,I271089,I271106,I271132,I271140,I270743,I270761,I271185,I271202,I270764,I270749,I270758,I270767,I271305,I915998,I271331,I271339,I915995,I916013,I271356,I916004,I271382,I271273,I271404,I916019,I271430,I271438,I916001,I271455,I271481,I271297,I271503,I271279,I916007,I271543,I271560,I271568,I271585,I271282,I271616,I916022,I271633,I916010,I271659,I271667,I271270,I271288,I271712,I916016,I271729,I271291,I271276,I271285,I271294,I271832,I568887,I271858,I271866,I568872,I568875,I271883,I568890,I271909,I271800,I271931,I568884,I271957,I271965,I271982,I272008,I271824,I272030,I271806,I568881,I272070,I272087,I272095,I272112,I271809,I272143,I568896,I272160,I568893,I272186,I272194,I271797,I271815,I272239,I568878,I272256,I271818,I271803,I271812,I271821,I272359,I906954,I272385,I272393,I906951,I906969,I272410,I906960,I272436,I272327,I272458,I906975,I272484,I272492,I906957,I272509,I272535,I272351,I272557,I272333,I906963,I272597,I272614,I272622,I272639,I272336,I272670,I906978,I272687,I906966,I272713,I272721,I272324,I272342,I272766,I906972,I272783,I272345,I272330,I272339,I272348,I272886,I1093050,I272912,I272920,I1093065,I272937,I1093068,I272963,I272985,I1093074,I273011,I273019,I1093056,I273036,I273062,I273084,I1093053,I273124,I273141,I273149,I273166,I273197,I1093059,I273214,I1093071,I273240,I273248,I273293,I1093062,I273310,I273413,I273439,I273447,I273464,I273490,I273512,I273538,I273546,I273563,I273589,I273611,I273651,I273668,I273676,I273693,I273724,I273741,I273767,I273775,I273820,I273837,I273940,I273966,I273974,I273991,I274017,I274039,I274065,I274073,I274090,I274116,I274138,I274178,I274195,I274203,I274220,I274251,I274268,I274294,I274302,I274347,I274364,I274467,I542877,I274493,I274501,I542862,I542865,I274518,I542880,I274544,I274435,I274566,I542874,I274592,I274600,I274617,I274643,I274459,I274665,I274441,I542871,I274705,I274722,I274730,I274747,I274444,I274778,I542886,I274795,I542883,I274821,I274829,I274432,I274450,I274874,I542868,I274891,I274453,I274438,I274447,I274456,I274994,I823858,I275020,I275028,I823861,I823855,I275045,I823867,I275071,I274962,I275093,I823870,I275119,I275127,I275144,I275170,I274986,I275192,I274968,I823873,I275232,I275249,I275257,I275274,I274971,I275305,I823864,I275322,I275348,I275356,I274959,I274977,I275401,I823876,I275418,I274980,I274965,I274974,I274983,I275521,I594319,I275547,I275555,I594304,I594307,I275572,I594322,I275598,I275489,I275620,I594316,I275646,I275654,I275671,I275697,I275513,I275719,I275495,I594313,I275759,I275776,I275784,I275801,I275498,I275832,I594328,I275849,I594325,I275875,I275883,I275486,I275504,I275928,I594310,I275945,I275507,I275492,I275501,I275510,I276048,I1130042,I276074,I276082,I1130057,I276099,I1130060,I276125,I276016,I276147,I1130066,I276173,I276181,I1130048,I276198,I276224,I276040,I276246,I276022,I1130045,I276286,I276303,I276311,I276328,I276025,I276359,I1130051,I276376,I1130063,I276402,I276410,I276013,I276031,I276455,I1130054,I276472,I276034,I276019,I276028,I276037,I276575,I1036511,I276601,I276609,I1036508,I276626,I1036520,I276652,I276543,I276674,I276700,I276708,I1036526,I276725,I276751,I276567,I276773,I276549,I1036514,I276813,I276830,I276838,I276855,I276552,I276886,I1036523,I1036529,I276903,I276929,I276937,I276540,I276558,I276982,I1036517,I276999,I276561,I276546,I276555,I276564,I277102,I277128,I277136,I277153,I277179,I277070,I277201,I277227,I277235,I277252,I277278,I277094,I277300,I277076,I277340,I277357,I277365,I277382,I277079,I277413,I277430,I277456,I277464,I277067,I277085,I277509,I277526,I277088,I277073,I277082,I277091,I277629,I277655,I277663,I277680,I277706,I277597,I277728,I277754,I277762,I277779,I277805,I277621,I277827,I277603,I277867,I277884,I277892,I277909,I277606,I277940,I277957,I277983,I277991,I277594,I277612,I278036,I278053,I277615,I277600,I277609,I277618,I278156,I453403,I278182,I278190,I453415,I453394,I278207,I453418,I278233,I278124,I278255,I453409,I278281,I278289,I453391,I278306,I278332,I278148,I278354,I278130,I453406,I278394,I278411,I278419,I278436,I278133,I278467,I453397,I278484,I453400,I278510,I278518,I278121,I278139,I278563,I453412,I278580,I278142,I278127,I278136,I278145,I278683,I1188998,I278709,I278717,I1189013,I278734,I1189016,I278760,I278651,I278782,I1189022,I278808,I278816,I1189004,I278833,I278859,I278675,I278881,I278657,I1189001,I278921,I278938,I278946,I278963,I278660,I278994,I1189007,I279011,I1189019,I279037,I279045,I278648,I278666,I279090,I1189010,I279107,I278669,I278654,I278663,I278672,I279210,I1148538,I279236,I279244,I1148553,I279261,I1148556,I279287,I279178,I279309,I1148562,I279335,I279343,I1148544,I279360,I279386,I279202,I279408,I279184,I1148541,I279448,I279465,I279473,I279490,I279187,I279521,I1148547,I279538,I1148559,I279564,I279572,I279175,I279193,I279617,I1148550,I279634,I279196,I279181,I279190,I279199,I279737,I1364238,I279763,I279771,I1364217,I279788,I1364244,I279814,I279836,I1364232,I279862,I279870,I1364235,I279887,I279913,I279935,I1364226,I279975,I279992,I280000,I280017,I280048,I1364223,I1364220,I280065,I1364241,I280091,I280099,I280144,I1364229,I280161,I280264,I832817,I280290,I280298,I832820,I832814,I280315,I832826,I280341,I280363,I832829,I280389,I280397,I280414,I280440,I280462,I832832,I280502,I280519,I280527,I280544,I280575,I832823,I280592,I280618,I280626,I280671,I832835,I280688,I280791,I280817,I280825,I280842,I280868,I280890,I280916,I280924,I280941,I280967,I280989,I281029,I281046,I281054,I281071,I281102,I281119,I281145,I281153,I281198,I281215,I281318,I683328,I281344,I281352,I683319,I683334,I281369,I683340,I281395,I281286,I281417,I683325,I281443,I281451,I281468,I281494,I281310,I281516,I281292,I683322,I281556,I281573,I281581,I281598,I281295,I281629,I683316,I683331,I281646,I281672,I281680,I281283,I281301,I281725,I683337,I281742,I281304,I281289,I281298,I281307,I281845,I791184,I281871,I281879,I791187,I791181,I281896,I791193,I281922,I281813,I281944,I791196,I281970,I281978,I281995,I282021,I281837,I282043,I281819,I791199,I282083,I282100,I282108,I282125,I281822,I282156,I791190,I282173,I282199,I282207,I281810,I281828,I282252,I791202,I282269,I281831,I281816,I281825,I281834,I282372,I637088,I282398,I282406,I637079,I637094,I282423,I637100,I282449,I282340,I282471,I637085,I282497,I282505,I282522,I282548,I282364,I282570,I282346,I637082,I282610,I282627,I282635,I282652,I282349,I282683,I637076,I637091,I282700,I282726,I282734,I282337,I282355,I282779,I637097,I282796,I282358,I282343,I282352,I282361,I282899,I738816,I282925,I282933,I738807,I738822,I282950,I738828,I282976,I282867,I282998,I738813,I283024,I283032,I283049,I283075,I282891,I283097,I282873,I738810,I283137,I283154,I283162,I283179,I282876,I283210,I738804,I738819,I283227,I283253,I283261,I282864,I282882,I283306,I738825,I283323,I282885,I282870,I282879,I282888,I283426,I283452,I283460,I283477,I283503,I283394,I283525,I283551,I283559,I283576,I283602,I283418,I283624,I283400,I283664,I283681,I283689,I283706,I283403,I283737,I283754,I283780,I283788,I283391,I283409,I283833,I283850,I283412,I283397,I283406,I283415,I283953,I1179172,I283979,I283987,I1179187,I284004,I1179190,I284030,I283921,I284052,I1179196,I284078,I284086,I1179178,I284103,I284129,I283945,I284151,I283927,I1179175,I284191,I284208,I284216,I284233,I283930,I284264,I1179181,I284281,I1179193,I284307,I284315,I283918,I283936,I284360,I1179184,I284377,I283939,I283924,I283933,I283942,I284480,I1097096,I284506,I284514,I1097111,I284531,I1097114,I284557,I284448,I284579,I1097120,I284605,I284613,I1097102,I284630,I284656,I284472,I284678,I284454,I1097099,I284718,I284735,I284743,I284760,I284457,I284791,I1097105,I284808,I1097117,I284834,I284842,I284445,I284463,I284887,I1097108,I284904,I284466,I284451,I284460,I284469,I285007,I285033,I285041,I285058,I285084,I284975,I285106,I285132,I285140,I285157,I285183,I284999,I285205,I284981,I285245,I285262,I285270,I285287,I284984,I285318,I285335,I285361,I285369,I284972,I284990,I285414,I285431,I284993,I284978,I284987,I284996,I285534,I1199980,I285560,I285568,I1199995,I285585,I1199998,I285611,I285502,I285633,I1200004,I285659,I285667,I1199986,I285684,I285710,I285526,I285732,I285508,I1199983,I285772,I285789,I285797,I285814,I285511,I285845,I1199989,I285862,I1200001,I285888,I285896,I285499,I285517,I285941,I1199992,I285958,I285520,I285505,I285514,I285523,I286061,I480603,I286087,I286095,I480615,I480594,I286112,I480618,I286138,I286029,I286160,I480609,I286186,I286194,I480591,I286211,I286237,I286053,I286259,I286035,I480606,I286299,I286316,I286324,I286341,I286038,I286372,I480597,I286389,I480600,I286415,I286423,I286026,I286044,I286468,I480612,I286485,I286047,I286032,I286041,I286050,I286588,I1288293,I286614,I286622,I1288290,I1288281,I286639,I1288278,I286665,I286556,I286687,I1288287,I286713,I286721,I1288296,I286738,I286764,I286580,I286786,I286562,I1288299,I286826,I286843,I286851,I286868,I286565,I286899,I1288284,I286916,I1288302,I286942,I286950,I286553,I286571,I286995,I287012,I286574,I286559,I286568,I286577,I287115,I1030340,I287141,I287149,I1030337,I287166,I1030349,I287192,I287083,I287214,I287240,I287248,I1030355,I287265,I287291,I287107,I287313,I287089,I1030343,I287353,I287370,I287378,I287395,I287092,I287426,I1030352,I1030358,I287443,I287469,I287477,I287080,I287098,I287522,I1030346,I287539,I287101,I287086,I287095,I287104,I287642,I456123,I287668,I287676,I456135,I456114,I287693,I456138,I287719,I287610,I287741,I456129,I287767,I287775,I456111,I287792,I287818,I287634,I287840,I287616,I456126,I287880,I287897,I287905,I287922,I287619,I287953,I456117,I287970,I456120,I287996,I288004,I287607,I287625,I288049,I456132,I288066,I287628,I287613,I287622,I287631,I288169,I1123684,I288195,I288203,I1123699,I288220,I1123702,I288246,I288137,I288268,I1123708,I288294,I288302,I1123690,I288319,I288345,I288161,I288367,I288143,I1123687,I288407,I288424,I288432,I288449,I288146,I288480,I1123693,I288497,I1123705,I288523,I288531,I288134,I288152,I288576,I1123696,I288593,I288155,I288140,I288149,I288158,I288696,I792238,I288722,I288730,I792241,I792235,I288747,I792247,I288773,I288664,I288795,I792250,I288821,I288829,I288846,I288872,I288688,I288894,I288670,I792253,I288934,I288951,I288959,I288976,I288673,I289007,I792244,I289024,I289050,I289058,I288661,I288679,I289103,I792256,I289120,I288682,I288667,I288676,I288685,I289223,I289249,I289257,I289274,I289300,I289191,I289322,I289348,I289356,I289373,I289399,I289215,I289421,I289197,I289461,I289478,I289486,I289503,I289200,I289534,I289551,I289577,I289585,I289188,I289206,I289630,I289647,I289209,I289194,I289203,I289212,I289750,I400635,I289776,I289784,I400647,I400626,I289801,I400650,I289827,I289718,I289849,I400641,I289875,I289883,I400623,I289900,I289926,I289742,I289948,I289724,I400638,I289988,I290005,I290013,I290030,I289727,I290061,I400629,I290078,I400632,I290104,I290112,I289715,I289733,I290157,I400644,I290174,I289736,I289721,I289730,I289739,I290277,I891450,I290303,I290311,I891447,I891465,I290328,I891456,I290354,I290245,I290376,I891471,I290402,I290410,I891453,I290427,I290453,I290269,I290475,I290251,I891459,I290515,I290532,I290540,I290557,I290254,I290588,I891474,I290605,I891462,I290631,I290639,I290242,I290260,I290684,I891468,I290701,I290263,I290248,I290257,I290266,I290804,I462107,I290830,I290838,I462119,I462098,I290855,I462122,I290881,I290772,I290903,I462113,I290929,I290937,I462095,I290954,I290980,I290796,I291002,I290778,I462110,I291042,I291059,I291067,I291084,I290781,I291115,I462101,I291132,I462104,I291158,I291166,I290769,I290787,I291211,I462116,I291228,I290790,I290775,I290784,I290793,I291331,I843357,I291357,I291365,I843360,I843354,I291382,I843366,I291408,I291299,I291430,I843369,I291456,I291464,I291481,I291507,I291323,I291529,I291305,I843372,I291569,I291586,I291594,I291611,I291308,I291642,I843363,I291659,I291685,I291693,I291296,I291314,I291738,I843375,I291755,I291317,I291302,I291311,I291320,I291858,I291884,I291892,I291909,I291935,I291826,I291957,I291983,I291991,I292008,I292034,I291850,I292056,I291832,I292096,I292113,I292121,I292138,I291835,I292169,I292186,I292212,I292220,I291823,I291841,I292265,I292282,I291844,I291829,I291838,I291847,I292385,I1116170,I292411,I292419,I1116185,I292436,I1116188,I292462,I292353,I292484,I1116194,I292510,I292518,I1116176,I292535,I292561,I292377,I292583,I292359,I1116173,I292623,I292640,I292648,I292665,I292362,I292696,I1116179,I292713,I1116191,I292739,I292747,I292350,I292368,I292792,I1116182,I292809,I292371,I292356,I292365,I292374,I292912,I480059,I292938,I292946,I480071,I480050,I292963,I480074,I292989,I292880,I293011,I480065,I293037,I293045,I480047,I293062,I293088,I292904,I293110,I292886,I480062,I293150,I293167,I293175,I293192,I292889,I293223,I480053,I293240,I480056,I293266,I293274,I292877,I292895,I293319,I480068,I293336,I292898,I292883,I292892,I292901,I293439,I589117,I293465,I293473,I589102,I589105,I293490,I589120,I293516,I293407,I293538,I589114,I293564,I293572,I293589,I293615,I293431,I293637,I293413,I589111,I293677,I293694,I293702,I293719,I293416,I293750,I589126,I293767,I589123,I293793,I293801,I293404,I293422,I293846,I589108,I293863,I293425,I293410,I293419,I293428,I293966,I910184,I293992,I294000,I910181,I910199,I294017,I910190,I294043,I294065,I910205,I294091,I294099,I910187,I294116,I294142,I294164,I910193,I294204,I294221,I294229,I294246,I294277,I910208,I294294,I910196,I294320,I294328,I294373,I910202,I294390,I294493,I1217236,I294519,I294527,I1217218,I1217242,I294544,I1217233,I294570,I294461,I294592,I1217239,I294618,I294626,I1217227,I294643,I294669,I294485,I294691,I294467,I294731,I294748,I294756,I294773,I294470,I294804,I1217224,I1217221,I294821,I1217230,I294847,I294855,I294458,I294476,I294900,I294917,I294479,I294464,I294473,I294482,I295020,I295046,I295054,I295071,I295097,I295119,I295145,I295153,I295170,I295196,I295218,I295258,I295275,I295283,I295300,I295331,I295348,I295374,I295382,I295427,I295444,I295547,I295573,I295581,I295598,I295624,I295515,I295646,I295672,I295680,I295697,I295723,I295539,I295745,I295521,I295785,I295802,I295810,I295827,I295524,I295858,I295875,I295901,I295909,I295512,I295530,I295954,I295971,I295533,I295518,I295527,I295536,I296074,I713962,I296100,I296108,I713953,I713968,I296125,I713974,I296151,I296042,I296173,I713959,I296199,I296207,I296224,I296250,I296066,I296272,I296048,I713956,I296312,I296329,I296337,I296354,I296051,I296385,I713950,I713965,I296402,I296428,I296436,I296039,I296057,I296481,I713971,I296498,I296060,I296045,I296054,I296063,I296601,I1392798,I296627,I296635,I1392777,I296652,I1392804,I296678,I296569,I296700,I1392792,I296726,I296734,I1392795,I296751,I296777,I296593,I296799,I296575,I1392786,I296839,I296856,I296864,I296881,I296578,I296912,I1392783,I1392780,I296929,I1392801,I296955,I296963,I296566,I296584,I297008,I1392789,I297025,I296587,I296572,I296581,I296590,I297128,I905016,I297154,I297162,I905013,I905031,I297179,I905022,I297205,I297096,I297227,I905037,I297253,I297261,I905019,I297278,I297304,I297120,I297326,I297102,I905025,I297366,I297383,I297391,I297408,I297105,I297439,I905040,I297456,I905028,I297482,I297490,I297093,I297111,I297535,I905034,I297552,I297114,I297099,I297108,I297117,I297655,I388667,I297681,I297689,I388679,I388658,I297706,I388682,I297732,I297623,I297754,I388673,I297780,I297788,I388655,I297805,I297831,I297647,I297853,I297629,I388670,I297893,I297910,I297918,I297935,I297632,I297966,I388661,I297983,I388664,I298009,I298017,I297620,I297638,I298062,I388676,I298079,I297641,I297626,I297635,I297644,I298182,I611081,I298208,I298216,I611066,I611069,I298233,I611084,I298259,I298150,I298281,I611078,I298307,I298315,I298332,I298358,I298174,I298380,I298156,I611075,I298420,I298437,I298445,I298462,I298159,I298493,I611090,I298510,I611087,I298536,I298544,I298147,I298165,I298589,I611072,I298606,I298168,I298153,I298162,I298171,I298709,I576401,I298735,I298743,I576386,I576389,I298760,I576404,I298786,I298677,I298808,I576398,I298834,I298842,I298859,I298885,I298701,I298907,I298683,I576395,I298947,I298964,I298972,I298989,I298686,I299020,I576410,I299037,I576407,I299063,I299071,I298674,I298692,I299116,I576392,I299133,I298695,I298680,I298689,I298698,I299236,I474619,I299262,I299270,I474631,I474610,I299287,I474634,I299313,I299204,I299335,I474625,I299361,I299369,I474607,I299386,I299412,I299228,I299434,I299210,I474622,I299474,I299491,I299499,I299516,I299213,I299547,I474613,I299564,I474616,I299590,I299598,I299201,I299219,I299643,I474628,I299660,I299222,I299207,I299216,I299225,I299763,I731880,I299789,I299797,I731871,I731886,I299814,I731892,I299840,I299731,I299862,I731877,I299888,I299896,I299913,I299939,I299755,I299961,I299737,I731874,I300001,I300018,I300026,I300043,I299740,I300074,I731868,I731883,I300091,I300117,I300125,I299728,I299746,I300170,I731889,I300187,I299749,I299734,I299743,I299752,I300290,I990934,I300316,I300324,I990931,I990949,I300341,I990940,I300367,I300258,I300389,I990955,I300415,I300423,I990937,I300440,I300466,I300282,I300488,I300264,I990943,I300528,I300545,I300553,I300570,I300267,I300601,I990958,I300618,I990946,I300644,I300652,I300255,I300273,I300697,I990952,I300714,I300276,I300261,I300270,I300279,I300817,I394651,I300843,I300851,I394663,I394642,I300868,I394666,I300894,I300916,I394657,I300942,I300950,I394639,I300967,I300993,I301015,I394654,I301055,I301072,I301080,I301097,I301128,I394645,I301145,I394648,I301171,I301179,I301224,I394660,I301241,I301344,I638244,I301370,I301378,I638235,I638250,I301395,I638256,I301421,I301312,I301443,I638241,I301469,I301477,I301494,I301520,I301336,I301542,I301318,I638238,I301582,I301599,I301607,I301624,I301321,I301655,I638232,I638247,I301672,I301698,I301706,I301309,I301327,I301751,I638253,I301768,I301330,I301315,I301324,I301333,I301871,I814372,I301897,I301905,I814375,I814369,I301922,I814381,I301948,I301839,I301970,I814384,I301996,I302004,I302021,I302047,I301863,I302069,I301845,I814387,I302109,I302126,I302134,I302151,I301848,I302182,I814378,I302199,I302225,I302233,I301836,I301854,I302278,I814390,I302295,I301857,I301842,I301851,I301860,I302398,I978660,I302424,I302432,I978657,I978675,I302449,I978666,I302475,I302497,I978681,I302523,I302531,I978663,I302548,I302574,I302596,I978669,I302636,I302653,I302661,I302678,I302709,I978684,I302726,I978672,I302752,I302760,I302805,I978678,I302822,I302925,I302951,I302959,I302976,I303002,I302893,I303024,I303050,I303058,I303075,I303101,I302917,I303123,I302899,I303163,I303180,I303188,I303205,I302902,I303236,I303253,I303279,I303287,I302890,I302908,I303332,I303349,I302911,I302896,I302905,I302914,I303452,I411515,I303478,I303486,I411527,I411506,I303503,I411530,I303529,I303420,I303551,I411521,I303577,I303585,I411503,I303602,I303628,I303444,I303650,I303426,I411518,I303690,I303707,I303715,I303732,I303429,I303763,I411509,I303780,I411512,I303806,I303814,I303417,I303435,I303859,I411524,I303876,I303438,I303423,I303432,I303441,I303979,I863910,I304005,I304013,I863913,I863907,I304030,I863919,I304056,I304078,I863922,I304104,I304112,I304129,I304155,I304177,I863925,I304217,I304234,I304242,I304259,I304290,I863916,I304307,I304333,I304341,I304386,I863928,I304403,I304506,I304532,I304540,I304557,I304583,I304474,I304605,I304631,I304639,I304656,I304682,I304498,I304704,I304480,I304744,I304761,I304769,I304786,I304483,I304817,I304834,I304860,I304868,I304471,I304489,I304913,I304930,I304492,I304477,I304486,I304495,I305033,I495877,I305059,I305067,I495889,I305084,I495874,I305110,I305001,I305132,I495898,I305158,I305166,I495895,I305183,I305209,I305025,I305231,I305007,I495886,I305271,I305288,I305296,I305313,I305010,I305344,I495883,I305361,I495892,I305387,I305395,I304998,I305016,I305440,I495880,I305457,I305019,I305004,I305013,I305022,I305560,I305586,I305594,I305611,I305637,I305528,I305659,I305685,I305693,I305710,I305736,I305552,I305758,I305534,I305798,I305815,I305823,I305840,I305537,I305871,I305888,I305914,I305922,I305525,I305543,I305967,I305984,I305546,I305531,I305540,I305549,I306087,I664254,I306113,I306121,I664245,I664260,I306138,I664266,I306164,I306186,I664251,I306212,I306220,I306237,I306263,I306285,I664248,I306325,I306342,I306350,I306367,I306398,I664242,I664257,I306415,I306441,I306449,I306494,I664263,I306511,I306614,I873923,I306640,I306648,I873926,I873920,I306665,I873932,I306691,I306713,I873935,I306739,I306747,I306764,I306790,I306812,I873938,I306852,I306869,I306877,I306894,I306925,I873929,I306942,I306968,I306976,I307021,I873941,I307038,I307141,I778009,I307167,I307175,I778012,I778006,I307192,I778018,I307218,I307109,I307240,I778021,I307266,I307274,I307291,I307317,I307133,I307339,I307115,I778024,I307379,I307396,I307404,I307421,I307118,I307452,I778015,I307469,I307495,I307503,I307106,I307124,I307548,I778027,I307565,I307127,I307112,I307121,I307130,I307668,I876031,I307694,I307702,I876034,I876028,I307719,I876040,I307745,I307636,I307767,I876043,I307793,I307801,I307818,I307844,I307660,I307866,I307642,I876046,I307906,I307923,I307931,I307948,I307645,I307979,I876037,I307996,I308022,I308030,I307633,I307651,I308075,I876049,I308092,I307654,I307639,I307648,I307657,I308195,I551547,I308221,I308229,I551532,I551535,I308246,I551550,I308272,I308294,I551544,I308320,I308328,I308345,I308371,I308393,I551541,I308433,I308450,I308458,I308475,I308506,I551556,I308523,I551553,I308549,I308557,I308602,I551538,I308619,I308722,I968324,I308748,I308756,I968321,I968339,I308773,I968330,I308799,I308690,I308821,I968345,I308847,I308855,I968327,I308872,I308898,I308714,I308920,I308696,I968333,I308960,I308977,I308985,I309002,I308699,I309033,I968348,I309050,I968336,I309076,I309084,I308687,I308705,I309129,I968342,I309146,I308708,I308693,I308702,I308711,I309249,I711072,I309275,I309283,I711063,I711078,I309300,I711084,I309326,I309217,I309348,I711069,I309374,I309382,I309399,I309425,I309241,I309447,I309223,I711066,I309487,I309504,I309512,I309529,I309226,I309560,I711060,I711075,I309577,I309603,I309611,I309214,I309232,I309656,I711081,I309673,I309235,I309220,I309229,I309238,I309776,I966386,I309802,I309810,I966383,I966401,I309827,I966392,I309853,I309744,I309875,I966407,I309901,I309909,I966389,I309926,I309952,I309768,I309974,I309750,I966395,I310014,I310031,I310039,I310056,I309753,I310087,I966410,I310104,I966398,I310130,I310138,I309741,I309759,I310183,I966404,I310200,I309762,I309747,I309756,I309765,I310303,I436539,I310329,I310337,I436551,I436530,I310354,I436554,I310380,I310402,I436545,I310428,I310436,I436527,I310453,I310479,I310501,I436542,I310541,I310558,I310566,I310583,I310614,I436533,I310631,I436536,I310657,I310665,I310710,I436548,I310727,I310830,I1099408,I310856,I310864,I1099423,I310881,I1099426,I310907,I310798,I310929,I1099432,I310955,I310963,I1099414,I310980,I311006,I310822,I311028,I310804,I1099411,I311068,I311085,I311093,I311110,I310807,I311141,I1099417,I311158,I1099429,I311184,I311192,I310795,I310813,I311237,I1099420,I311254,I310816,I310801,I310810,I310819,I311357,I311383,I311391,I311408,I311434,I311325,I311456,I311482,I311490,I311507,I311533,I311349,I311555,I311331,I311595,I311612,I311620,I311637,I311334,I311668,I311685,I311711,I311719,I311322,I311340,I311764,I311781,I311343,I311328,I311337,I311346,I311884,I1250964,I311910,I311918,I1250946,I1250970,I311935,I1250961,I311961,I311852,I311983,I1250967,I312009,I312017,I1250955,I312034,I312060,I311876,I312082,I311858,I312122,I312139,I312147,I312164,I311861,I312195,I1250952,I1250949,I312212,I1250958,I312238,I312246,I311849,I311867,I312291,I312308,I311870,I311855,I311864,I311873,I312411,I1061838,I312437,I312445,I1061853,I312462,I1061856,I312488,I312379,I312510,I1061862,I312536,I312544,I1061844,I312561,I312587,I312403,I312609,I312385,I1061841,I312649,I312666,I312674,I312691,I312388,I312722,I1061847,I312739,I1061859,I312765,I312773,I312376,I312394,I312818,I1061850,I312835,I312397,I312382,I312391,I312400,I312938,I952174,I312964,I312972,I952171,I952189,I312989,I952180,I313015,I313037,I952195,I313063,I313071,I952177,I313088,I313114,I313136,I952183,I313176,I313193,I313201,I313218,I313249,I952198,I313266,I952186,I313292,I313300,I313345,I952192,I313362,I313465,I572933,I313491,I313499,I572918,I572921,I313516,I572936,I313542,I313433,I313564,I572930,I313590,I313598,I313615,I313641,I313457,I313663,I313439,I572927,I313703,I313720,I313728,I313745,I313442,I313776,I572942,I313793,I572939,I313819,I313827,I313430,I313448,I313872,I572924,I313889,I313451,I313436,I313445,I313454,I313992,I314018,I314026,I314043,I314069,I313960,I314091,I314117,I314125,I314142,I314168,I313984,I314190,I313966,I314230,I314247,I314255,I314272,I313969,I314303,I314320,I314346,I314354,I313957,I313975,I314399,I314416,I313978,I313963,I313972,I313981,I314519,I953466,I314545,I314553,I953463,I953481,I314570,I953472,I314596,I314487,I314618,I953487,I314644,I314652,I953469,I314669,I314695,I314511,I314717,I314493,I953475,I314757,I314774,I314782,I314799,I314496,I314830,I953490,I314847,I953478,I314873,I314881,I314484,I314502,I314926,I953484,I314943,I314505,I314490,I314499,I314508,I315046,I315072,I315080,I315097,I315123,I315014,I315145,I315171,I315179,I315196,I315222,I315038,I315244,I315020,I315284,I315301,I315309,I315326,I315023,I315357,I315374,I315400,I315408,I315011,I315029,I315453,I315470,I315032,I315017,I315026,I315035,I315573,I804359,I315599,I315607,I804362,I804356,I315624,I804368,I315650,I315672,I804371,I315698,I315706,I315723,I315749,I315771,I804374,I315811,I315828,I315836,I315853,I315884,I804365,I315901,I315927,I315935,I315980,I804377,I315997,I316100,I1311878,I316126,I316134,I1311857,I316151,I1311884,I316177,I316199,I1311872,I316225,I316233,I1311875,I316250,I316276,I316298,I1311866,I316338,I316355,I316363,I316380,I316411,I1311863,I1311860,I316428,I1311881,I316454,I316462,I316507,I1311869,I316524,I316627,I1384468,I316653,I316661,I1384447,I316678,I1384474,I316704,I316595,I316726,I1384462,I316752,I316760,I1384465,I316777,I316803,I316619,I316825,I316601,I1384456,I316865,I316882,I316890,I316907,I316604,I316938,I1384453,I1384450,I316955,I1384471,I316981,I316989,I316592,I316610,I317034,I1384459,I317051,I316613,I316598,I316607,I316616,I317154,I1052219,I317180,I317188,I1052216,I317205,I1052228,I317231,I317122,I317253,I317279,I317287,I1052234,I317304,I317330,I317146,I317352,I317128,I1052222,I317392,I317409,I317417,I317434,I317131,I317465,I1052231,I1052237,I317482,I317508,I317516,I317119,I317137,I317561,I1052225,I317578,I317140,I317125,I317134,I317143,I317681,I317707,I317715,I317732,I317758,I317649,I317780,I317806,I317814,I317831,I317857,I317673,I317879,I317655,I317919,I317936,I317944,I317961,I317658,I317992,I318009,I318035,I318043,I317646,I317664,I318088,I318105,I317667,I317652,I317661,I317670,I318208,I1179750,I318234,I318242,I1179765,I318259,I1179768,I318285,I318176,I318307,I1179774,I318333,I318341,I1179756,I318358,I318384,I318200,I318406,I318182,I1179753,I318446,I318463,I318471,I318488,I318185,I318519,I1179759,I318536,I1179771,I318562,I318570,I318173,I318191,I318615,I1179762,I318632,I318194,I318179,I318188,I318197,I318735,I1003854,I318761,I318769,I1003851,I1003869,I318786,I1003860,I318812,I318703,I318834,I1003875,I318860,I318868,I1003857,I318885,I318911,I318727,I318933,I318709,I1003863,I318973,I318990,I318998,I319015,I318712,I319046,I1003878,I319063,I1003866,I319089,I319097,I318700,I318718,I319142,I1003872,I319159,I318721,I318706,I318715,I318724,I319262,I1152006,I319288,I319296,I1152021,I319313,I1152024,I319339,I319230,I319361,I1152030,I319387,I319395,I1152012,I319412,I319438,I319254,I319460,I319236,I1152009,I319500,I319517,I319525,I319542,I319239,I319573,I1152015,I319590,I1152027,I319616,I319624,I319227,I319245,I319669,I1152018,I319686,I319248,I319233,I319242,I319251,I319789,I412059,I319815,I319823,I412071,I412050,I319840,I412074,I319866,I319757,I319888,I412065,I319914,I319922,I412047,I319939,I319965,I319781,I319987,I319763,I412062,I320027,I320044,I320052,I320069,I319766,I320100,I412053,I320117,I412056,I320143,I320151,I319754,I319772,I320196,I412068,I320213,I319775,I319760,I319769,I319778,I320316,I535742,I320342,I320350,I535754,I320367,I535739,I320393,I320284,I320415,I535763,I320441,I320449,I535760,I320466,I320492,I320308,I320514,I320290,I535751,I320554,I320571,I320579,I320596,I320293,I320627,I535748,I320644,I535757,I320670,I320678,I320281,I320299,I320723,I535745,I320740,I320302,I320287,I320296,I320305,I320843,I1145648,I320869,I320877,I1145663,I320894,I1145666,I320920,I320811,I320942,I1145672,I320968,I320976,I1145654,I320993,I321019,I320835,I321041,I320817,I1145651,I321081,I321098,I321106,I321123,I320820,I321154,I1145657,I321171,I1145669,I321197,I321205,I320808,I320826,I321250,I1145660,I321267,I320829,I320814,I320823,I320832,I321370,I849154,I321396,I321404,I849157,I849151,I321421,I849163,I321447,I321338,I321469,I849166,I321495,I321503,I321520,I321546,I321362,I321568,I321344,I849169,I321608,I321625,I321633,I321650,I321347,I321681,I849160,I321698,I321724,I321732,I321335,I321353,I321777,I849172,I321794,I321356,I321341,I321350,I321359,I321897,I382139,I321923,I321931,I382151,I382130,I321948,I382154,I321974,I321865,I321996,I382145,I322022,I322030,I382127,I322047,I322073,I321889,I322095,I321871,I382142,I322135,I322152,I322160,I322177,I321874,I322208,I382133,I322225,I382136,I322251,I322259,I321862,I321880,I322304,I382148,I322321,I321883,I321868,I321877,I321886,I322424,I322450,I322458,I322475,I322501,I322392,I322523,I322549,I322557,I322574,I322600,I322416,I322622,I322398,I322662,I322679,I322687,I322704,I322401,I322735,I322752,I322778,I322786,I322389,I322407,I322831,I322848,I322410,I322395,I322404,I322413,I322951,I322977,I322985,I323002,I323028,I322919,I323050,I323076,I323084,I323101,I323127,I322943,I323149,I322925,I323189,I323206,I323214,I323231,I322928,I323262,I323279,I323305,I323313,I322916,I322934,I323358,I323375,I322937,I322922,I322931,I322940,I323478,I1367213,I323504,I323512,I1367192,I323529,I1367219,I323555,I323577,I1367207,I323603,I323611,I1367210,I323628,I323654,I323676,I1367201,I323716,I323733,I323741,I323758,I323789,I1367198,I1367195,I323806,I1367216,I323832,I323840,I323885,I1367204,I323902,I324005,I451227,I324031,I324039,I451239,I451218,I324056,I451242,I324082,I323973,I324104,I451233,I324130,I324138,I451215,I324155,I324181,I323997,I324203,I323979,I451230,I324243,I324260,I324268,I324285,I323982,I324316,I451221,I324333,I451224,I324359,I324367,I323970,I323988,I324412,I451236,I324429,I323991,I323976,I323985,I323994,I324532,I774652,I324558,I324566,I774643,I774658,I324583,I774664,I324609,I324500,I324631,I774649,I324657,I324665,I324682,I324708,I324524,I324730,I324506,I774646,I324770,I324787,I324795,I324812,I324509,I324843,I774640,I774655,I324860,I324886,I324894,I324497,I324515,I324939,I774661,I324956,I324518,I324503,I324512,I324521,I325059,I325085,I325093,I325110,I325136,I325027,I325158,I325184,I325192,I325209,I325235,I325051,I325257,I325033,I325297,I325314,I325322,I325339,I325036,I325370,I325387,I325413,I325421,I325024,I325042,I325466,I325483,I325045,I325030,I325039,I325048,I325586,I387035,I325612,I325620,I387047,I387026,I325637,I387050,I325663,I325554,I325685,I387041,I325711,I325719,I387023,I325736,I325762,I325578,I325784,I325560,I387038,I325824,I325841,I325849,I325866,I325563,I325897,I387029,I325914,I387032,I325940,I325948,I325551,I325569,I325993,I387044,I326010,I325572,I325557,I325566,I325575,I326113,I1165300,I326139,I326147,I1165315,I326164,I1165318,I326190,I326212,I1165324,I326238,I326246,I1165306,I326263,I326289,I326311,I1165303,I326351,I326368,I326376,I326393,I326424,I1165309,I326441,I1165321,I326467,I326475,I326520,I1165312,I326537,I326640,I627262,I326666,I326674,I627253,I627268,I326691,I627274,I326717,I326608,I326739,I627259,I326765,I326773,I326790,I326816,I326632,I326838,I326614,I627256,I326878,I326895,I326903,I326920,I326617,I326951,I627250,I627265,I326968,I326994,I327002,I326605,I326623,I327047,I627271,I327064,I326626,I326611,I326620,I326629,I327167,I327193,I327201,I327218,I327244,I327135,I327266,I327292,I327300,I327317,I327343,I327159,I327365,I327141,I327405,I327422,I327430,I327447,I327144,I327478,I327495,I327521,I327529,I327132,I327150,I327574,I327591,I327153,I327138,I327147,I327156,I327694,I1313068,I327720,I327728,I1313047,I327745,I1313074,I327771,I327662,I327793,I1313062,I327819,I327827,I1313065,I327844,I327870,I327686,I327892,I327668,I1313056,I327932,I327949,I327957,I327974,I327671,I328005,I1313053,I1313050,I328022,I1313071,I328048,I328056,I327659,I327677,I328101,I1313059,I328118,I327680,I327665,I327674,I327683,I328221,I657318,I328247,I328255,I657309,I657324,I328272,I657330,I328298,I328189,I328320,I657315,I328346,I328354,I328371,I328397,I328213,I328419,I328195,I657312,I328459,I328476,I328484,I328501,I328198,I328532,I657306,I657321,I328549,I328575,I328583,I328186,I328204,I328628,I657327,I328645,I328207,I328192,I328201,I328210,I328748,I328774,I328782,I328799,I328825,I328716,I328847,I328873,I328881,I328898,I328924,I328740,I328946,I328722,I328986,I329003,I329011,I329028,I328725,I329059,I329076,I329102,I329110,I328713,I328731,I329155,I329172,I328734,I328719,I328728,I328737,I329275,I329301,I329309,I329326,I329352,I329243,I329374,I329400,I329408,I329425,I329451,I329267,I329473,I329249,I329513,I329530,I329538,I329555,I329252,I329586,I329603,I329629,I329637,I329240,I329258,I329682,I329699,I329261,I329246,I329255,I329264,I329802,I1007730,I329828,I329836,I1007727,I1007745,I329853,I1007736,I329879,I329901,I1007751,I329927,I329935,I1007733,I329952,I329978,I330000,I1007739,I330040,I330057,I330065,I330082,I330113,I1007754,I330130,I1007742,I330156,I330164,I330209,I1007748,I330226,I330329,I1206356,I330355,I330363,I1206338,I1206362,I330380,I1206353,I330406,I330297,I330428,I1206359,I330454,I330462,I1206347,I330479,I330505,I330321,I330527,I330303,I330567,I330584,I330592,I330609,I330306,I330640,I1206344,I1206341,I330657,I1206350,I330683,I330691,I330294,I330312,I330736,I330753,I330315,I330300,I330309,I330318,I330856,I394107,I330882,I330890,I394119,I394098,I330907,I394122,I330933,I330824,I330955,I394113,I330981,I330989,I394095,I331006,I331032,I330848,I331054,I330830,I394110,I331094,I331111,I331119,I331136,I330833,I331167,I394101,I331184,I394104,I331210,I331218,I330821,I330839,I331263,I394116,I331280,I330842,I330827,I330836,I330845,I331383,I1072820,I331409,I331417,I1072835,I331434,I1072838,I331460,I331351,I331482,I1072844,I331508,I331516,I1072826,I331533,I331559,I331375,I331581,I331357,I1072823,I331621,I331638,I331646,I331663,I331360,I331694,I1072829,I331711,I1072841,I331737,I331745,I331348,I331366,I331790,I1072832,I331807,I331369,I331354,I331363,I331372,I331910,I735926,I331936,I331944,I735917,I735932,I331961,I735938,I331987,I332009,I735923,I332035,I332043,I332060,I332086,I332108,I735920,I332148,I332165,I332173,I332190,I332221,I735914,I735929,I332238,I332264,I332272,I332317,I735935,I332334,I332437,I332463,I332471,I332488,I332514,I332405,I332536,I332562,I332570,I332587,I332613,I332429,I332635,I332411,I332675,I332692,I332700,I332717,I332414,I332748,I332765,I332791,I332799,I332402,I332420,I332844,I332861,I332423,I332408,I332417,I332426,I332964,I332990,I332998,I333015,I333041,I332932,I333063,I333089,I333097,I333114,I333140,I332956,I333162,I332938,I333202,I333219,I333227,I333244,I332941,I333275,I333292,I333318,I333326,I332929,I332947,I333371,I333388,I332950,I332935,I332944,I332953,I333491,I333517,I333525,I333542,I333568,I333459,I333590,I333616,I333624,I333641,I333667,I333483,I333689,I333465,I333729,I333746,I333754,I333771,I333468,I333802,I333819,I333845,I333853,I333456,I333474,I333898,I333915,I333477,I333462,I333471,I333480,I334018,I861802,I334044,I334052,I861805,I861799,I334069,I861811,I334095,I333986,I334117,I861814,I334143,I334151,I334168,I334194,I334010,I334216,I333992,I861817,I334256,I334273,I334281,I334298,I333995,I334329,I861808,I334346,I334372,I334380,I333983,I334001,I334425,I861820,I334442,I334004,I333989,I333998,I334007,I334545,I452315,I334571,I334579,I452327,I452306,I334596,I452330,I334622,I334513,I334644,I452321,I334670,I334678,I452303,I334695,I334721,I334537,I334743,I334519,I452318,I334783,I334800,I334808,I334825,I334522,I334856,I452309,I334873,I452312,I334899,I334907,I334510,I334528,I334952,I452324,I334969,I334531,I334516,I334525,I334534,I335072,I915352,I335098,I335106,I915349,I915367,I335123,I915358,I335149,I335040,I335171,I915373,I335197,I335205,I915355,I335222,I335248,I335064,I335270,I335046,I915361,I335310,I335327,I335335,I335352,I335049,I335383,I915376,I335400,I915364,I335426,I335434,I335037,I335055,I335479,I915370,I335496,I335058,I335043,I335052,I335061,I335599,I1056146,I335625,I335633,I1056143,I335650,I1056155,I335676,I335698,I335724,I335732,I1056161,I335749,I335775,I335797,I1056149,I335837,I335854,I335862,I335879,I335910,I1056158,I1056164,I335927,I335953,I335961,I336006,I1056152,I336023,I336126,I909538,I336152,I336160,I909535,I909553,I336177,I909544,I336203,I336094,I336225,I909559,I336251,I336259,I909541,I336276,I336302,I336118,I336324,I336100,I909547,I336364,I336381,I336389,I336406,I336103,I336437,I909562,I336454,I909550,I336480,I336488,I336091,I336109,I336533,I909556,I336550,I336112,I336097,I336106,I336115,I336653,I1149694,I336679,I336687,I1149709,I336704,I1149712,I336730,I336752,I1149718,I336778,I336786,I1149700,I336803,I336829,I336851,I1149697,I336891,I336908,I336916,I336933,I336964,I1149703,I336981,I1149715,I337007,I337015,I337060,I1149706,I337077,I337180,I1190154,I337206,I337214,I1190169,I337231,I1190172,I337257,I337148,I337279,I1190178,I337305,I337313,I1190160,I337330,I337356,I337172,I337378,I337154,I1190157,I337418,I337435,I337443,I337460,I337157,I337491,I1190163,I337508,I1190175,I337534,I337542,I337145,I337163,I337587,I1190166,I337604,I337166,I337151,I337160,I337169,I337707,I508372,I337733,I337741,I508384,I337758,I508369,I337784,I337675,I337806,I508393,I337832,I337840,I508390,I337857,I337883,I337699,I337905,I337681,I508381,I337945,I337962,I337970,I337987,I337684,I338018,I508378,I338035,I508387,I338061,I338069,I337672,I337690,I338114,I508375,I338131,I337693,I337678,I337687,I337696,I338234,I1175126,I338260,I338268,I1175141,I338285,I1175144,I338311,I338202,I338333,I1175150,I338359,I338367,I1175132,I338384,I338410,I338226,I338432,I338208,I1175129,I338472,I338489,I338497,I338514,I338211,I338545,I1175135,I338562,I1175147,I338588,I338596,I338199,I338217,I338641,I1175138,I338658,I338220,I338205,I338214,I338223,I338761,I573511,I338787,I338795,I573496,I573499,I338812,I573514,I338838,I338729,I338860,I573508,I338886,I338894,I338911,I338937,I338753,I338959,I338735,I573505,I338999,I339016,I339024,I339041,I338738,I339072,I573520,I339089,I573517,I339115,I339123,I338726,I338744,I339168,I573502,I339185,I338747,I338732,I338741,I338750,I339288,I1164144,I339314,I339322,I1164159,I339339,I1164162,I339365,I339256,I339387,I1164168,I339413,I339421,I1164150,I339438,I339464,I339280,I339486,I339262,I1164147,I339526,I339543,I339551,I339568,I339265,I339599,I1164153,I339616,I1164165,I339642,I339650,I339253,I339271,I339695,I1164156,I339712,I339274,I339259,I339268,I339277,I339815,I1165878,I339841,I339849,I1165893,I339866,I1165896,I339892,I339914,I1165902,I339940,I339948,I1165884,I339965,I339991,I340013,I1165881,I340053,I340070,I340078,I340095,I340126,I1165887,I340143,I1165899,I340169,I340177,I340222,I1165890,I340239,I340342,I739394,I340368,I340376,I739385,I739400,I340393,I739406,I340419,I340310,I340441,I739391,I340467,I340475,I340492,I340518,I340334,I340540,I340316,I739388,I340580,I340597,I340605,I340622,I340319,I340653,I739382,I739397,I340670,I340696,I340704,I340307,I340325,I340749,I739403,I340766,I340328,I340313,I340322,I340331,I340869,I1296370,I340895,I340903,I1296397,I1296373,I340920,I1296382,I340946,I340837,I340968,I340994,I341002,I1296394,I341019,I341045,I340861,I341067,I340843,I1296376,I341107,I341124,I341132,I341149,I340846,I341180,I1296391,I1296379,I341197,I1296385,I341223,I341231,I340834,I340852,I341276,I1296388,I341293,I340855,I340840,I340849,I340858,I341396,I1322588,I341422,I341430,I1322567,I341447,I1322594,I341473,I341364,I341495,I1322582,I341521,I341529,I1322585,I341546,I341572,I341388,I341594,I341370,I1322576,I341634,I341651,I341659,I341676,I341373,I341707,I1322573,I1322570,I341724,I1322591,I341750,I341758,I341361,I341379,I341803,I1322579,I341820,I341382,I341367,I341376,I341385,I341923,I341949,I341957,I341974,I342000,I341891,I342022,I342048,I342056,I342073,I342099,I341915,I342121,I341897,I342161,I342178,I342186,I342203,I341900,I342234,I342251,I342277,I342285,I341888,I341906,I342330,I342347,I341909,I341894,I341903,I341912,I342450,I920520,I342476,I342484,I920517,I920535,I342501,I920526,I342527,I342418,I342549,I920541,I342575,I342583,I920523,I342600,I342626,I342442,I342648,I342424,I920529,I342688,I342705,I342713,I342730,I342427,I342761,I920544,I342778,I920532,I342804,I342812,I342415,I342433,I342857,I920538,I342874,I342436,I342421,I342430,I342439,I342977,I397915,I343003,I343011,I397927,I397906,I343028,I397930,I343054,I342945,I343076,I397921,I343102,I343110,I397903,I343127,I343153,I342969,I343175,I342951,I397918,I343215,I343232,I343240,I343257,I342954,I343288,I397909,I343305,I397912,I343331,I343339,I342942,I342960,I343384,I397924,I343401,I342963,I342948,I342957,I342966,I343504,I413691,I343530,I343538,I413703,I413682,I343555,I413706,I343581,I343472,I343603,I413697,I343629,I343637,I413679,I343654,I343680,I343496,I343702,I343478,I413694,I343742,I343759,I343767,I343784,I343481,I343815,I413685,I343832,I413688,I343858,I343866,I343469,I343487,I343911,I413700,I343928,I343490,I343475,I343484,I343493,I344031,I384315,I344057,I344065,I384327,I384306,I344082,I384330,I344108,I343999,I344130,I384321,I344156,I344164,I384303,I344181,I344207,I344023,I344229,I344005,I384318,I344269,I344286,I344294,I344311,I344008,I344342,I384309,I344359,I384312,I344385,I344393,I343996,I344014,I344438,I384324,I344455,I344017,I344002,I344011,I344020,I344558,I1101720,I344584,I344592,I1101735,I344609,I1101738,I344635,I344526,I344657,I1101744,I344683,I344691,I1101726,I344708,I344734,I344550,I344756,I344532,I1101723,I344796,I344813,I344821,I344838,I344535,I344869,I1101729,I344886,I1101741,I344912,I344920,I344523,I344541,I344965,I1101732,I344982,I344544,I344529,I344538,I344547,I345085,I914706,I345111,I345119,I914703,I914721,I345136,I914712,I345162,I345053,I345184,I914727,I345210,I345218,I914709,I345235,I345261,I345077,I345283,I345059,I914715,I345323,I345340,I345348,I345365,I345062,I345396,I914730,I345413,I914718,I345439,I345447,I345050,I345068,I345492,I914724,I345509,I345071,I345056,I345065,I345074,I345612,I1303102,I345638,I345646,I1303129,I1303105,I345663,I1303114,I345689,I345580,I345711,I345737,I345745,I1303126,I345762,I345788,I345604,I345810,I345586,I1303108,I345850,I345867,I345875,I345892,I345589,I345923,I1303123,I1303111,I345940,I1303117,I345966,I345974,I345577,I345595,I346019,I1303120,I346036,I345598,I345583,I345592,I345601,I346139,I346165,I346173,I346190,I346216,I346238,I346264,I346272,I346289,I346315,I346337,I346377,I346394,I346402,I346419,I346450,I346467,I346493,I346501,I346546,I346563,I346666,I346692,I346700,I346717,I346743,I346634,I346765,I346791,I346799,I346816,I346842,I346658,I346864,I346640,I346904,I346921,I346929,I346946,I346643,I346977,I346994,I347020,I347028,I346631,I346649,I347073,I347090,I346652,I346637,I346646,I346655,I347193,I347219,I347227,I347244,I347270,I347161,I347292,I347318,I347326,I347343,I347369,I347185,I347391,I347167,I347431,I347448,I347456,I347473,I347170,I347504,I347521,I347547,I347555,I347158,I347176,I347600,I347617,I347179,I347164,I347173,I347182,I347720,I347746,I347754,I347771,I347797,I347688,I347819,I347845,I347853,I347870,I347896,I347712,I347918,I347694,I347958,I347975,I347983,I348000,I347697,I348031,I348048,I348074,I348082,I347685,I347703,I348127,I348144,I347706,I347691,I347700,I347709,I348247,I635354,I348273,I348281,I635345,I635360,I348298,I635366,I348324,I348215,I348346,I635351,I348372,I348380,I348397,I348423,I348239,I348445,I348221,I635348,I348485,I348502,I348510,I348527,I348224,I348558,I635342,I635357,I348575,I348601,I348609,I348212,I348230,I348654,I635363,I348671,I348233,I348218,I348227,I348236,I348774,I1002562,I348800,I348808,I1002559,I1002577,I348825,I1002568,I348851,I348742,I348873,I1002583,I348899,I348907,I1002565,I348924,I348950,I348766,I348972,I348748,I1002571,I349012,I349029,I349037,I349054,I348751,I349085,I1002586,I349102,I1002574,I349128,I349136,I348739,I348757,I349181,I1002580,I349198,I348760,I348745,I348754,I348763,I349301,I828074,I349327,I349335,I828077,I828071,I349352,I828083,I349378,I349269,I349400,I828086,I349426,I349434,I349451,I349477,I349293,I349499,I349275,I828089,I349539,I349556,I349564,I349581,I349278,I349612,I828080,I349629,I349655,I349663,I349266,I349284,I349708,I828092,I349725,I349287,I349272,I349281,I349290,I349828,I1078600,I349854,I349862,I1078615,I349879,I1078618,I349905,I349796,I349927,I1078624,I349953,I349961,I1078606,I349978,I350004,I349820,I350026,I349802,I1078603,I350066,I350083,I350091,I350108,I349805,I350139,I1078609,I350156,I1078621,I350182,I350190,I349793,I349811,I350235,I1078612,I350252,I349814,I349799,I349808,I349817,I350355,I983182,I350381,I350389,I983179,I983197,I350406,I983188,I350432,I350323,I350454,I983203,I350480,I350488,I983185,I350505,I350531,I350347,I350553,I350329,I983191,I350593,I350610,I350618,I350635,I350332,I350666,I983206,I350683,I983194,I350709,I350717,I350320,I350338,I350762,I983200,I350779,I350341,I350326,I350335,I350344,I350882,I833344,I350908,I350916,I833347,I833341,I350933,I833353,I350959,I350850,I350981,I833356,I351007,I351015,I351032,I351058,I350874,I351080,I350856,I833359,I351120,I351137,I351145,I351162,I350859,I351193,I833350,I351210,I351236,I351244,I350847,I350865,I351289,I833362,I351306,I350868,I350853,I350862,I350871,I351409,I385947,I351435,I351443,I385959,I385938,I351460,I385962,I351486,I351377,I351508,I385953,I351534,I351542,I385935,I351559,I351585,I351401,I351607,I351383,I385950,I351647,I351664,I351672,I351689,I351386,I351720,I385941,I351737,I385944,I351763,I351771,I351374,I351392,I351816,I385956,I351833,I351395,I351380,I351389,I351398,I351936,I351962,I351970,I351987,I352013,I352035,I352061,I352069,I352086,I352112,I352134,I352174,I352191,I352199,I352216,I352247,I352264,I352290,I352298,I352343,I352360,I352463,I352489,I352497,I352514,I352540,I352431,I352562,I352588,I352596,I352613,I352639,I352455,I352661,I352437,I352701,I352718,I352726,I352743,I352440,I352774,I352791,I352817,I352825,I352428,I352446,I352870,I352887,I352449,I352434,I352443,I352452,I352990,I353016,I353024,I353041,I353067,I352958,I353089,I353115,I353123,I353140,I353166,I352982,I353188,I352964,I353228,I353245,I353253,I353270,I352967,I353301,I353318,I353344,I353352,I352955,I352973,I353397,I353414,I352976,I352961,I352970,I352979,I353517,I353543,I353551,I353568,I353594,I353485,I353616,I353642,I353650,I353667,I353693,I353509,I353715,I353491,I353755,I353772,I353780,I353797,I353494,I353828,I353845,I353871,I353879,I353482,I353500,I353924,I353941,I353503,I353488,I353497,I353506,I354044,I354070,I354078,I354095,I354121,I354012,I354143,I354169,I354177,I354194,I354220,I354036,I354242,I354018,I354282,I354299,I354307,I354324,I354021,I354355,I354372,I354398,I354406,I354009,I354027,I354451,I354468,I354030,I354015,I354024,I354033,I354571,I451771,I354597,I354605,I451783,I451762,I354622,I451786,I354648,I354670,I451777,I354696,I354704,I451759,I354721,I354747,I354769,I451774,I354809,I354826,I354834,I354851,I354882,I451765,I354899,I451768,I354925,I354933,I354978,I451780,I354995,I355098,I526817,I355124,I355132,I526829,I355149,I526814,I355175,I355066,I355197,I526838,I355223,I355231,I526835,I355248,I355274,I355090,I355296,I355072,I526826,I355336,I355353,I355361,I355378,I355075,I355409,I526823,I355426,I526832,I355452,I355460,I355063,I355081,I355505,I526820,I355522,I355084,I355069,I355078,I355087,I355625,I768872,I355651,I355659,I768863,I768878,I355676,I768884,I355702,I355593,I355724,I768869,I355750,I355758,I355775,I355801,I355617,I355823,I355599,I768866,I355863,I355880,I355888,I355905,I355602,I355936,I768860,I768875,I355953,I355979,I355987,I355590,I355608,I356032,I768881,I356049,I355611,I355596,I355605,I355614,I356152,I1126574,I356178,I356186,I1126589,I356203,I1126592,I356229,I356120,I356251,I1126598,I356277,I356285,I1126580,I356302,I356328,I356144,I356350,I356126,I1126577,I356390,I356407,I356415,I356432,I356129,I356463,I1126583,I356480,I1126595,I356506,I356514,I356117,I356135,I356559,I1126586,I356576,I356138,I356123,I356132,I356141,I356679,I1244436,I356705,I356713,I1244418,I1244442,I356730,I1244433,I356756,I356647,I356778,I1244439,I356804,I356812,I1244427,I356829,I356855,I356671,I356877,I356653,I356917,I356934,I356942,I356959,I356656,I356990,I1244424,I1244421,I357007,I1244430,I357033,I357041,I356644,I356662,I357086,I357103,I356665,I356650,I356659,I356668,I357206,I357232,I357240,I357257,I357283,I357174,I357305,I357331,I357339,I357356,I357382,I357198,I357404,I357180,I357444,I357461,I357469,I357486,I357183,I357517,I357534,I357560,I357568,I357171,I357189,I357613,I357630,I357192,I357177,I357186,I357195,I357733,I458299,I357759,I357767,I458311,I458290,I357784,I458314,I357810,I357701,I357832,I458305,I357858,I357866,I458287,I357883,I357909,I357725,I357931,I357707,I458302,I357971,I357988,I357996,I358013,I357710,I358044,I458293,I358061,I458296,I358087,I358095,I357698,I357716,I358140,I458308,I358157,I357719,I357704,I357713,I357722,I358260,I358286,I358294,I358311,I358337,I358228,I358359,I358385,I358393,I358410,I358436,I358252,I358458,I358234,I358498,I358515,I358523,I358540,I358237,I358571,I358588,I358614,I358622,I358225,I358243,I358667,I358684,I358246,I358231,I358240,I358249,I358787,I358813,I358821,I358838,I358864,I358886,I358912,I358920,I358937,I358963,I358985,I359025,I359042,I359050,I359067,I359098,I359115,I359141,I359149,I359194,I359211,I359314,I1347578,I359340,I359348,I1347557,I359365,I1347584,I359391,I359413,I1347572,I359439,I359447,I1347575,I359464,I359490,I359512,I1347566,I359552,I359569,I359577,I359594,I359625,I1347563,I1347560,I359642,I1347581,I359668,I359676,I359721,I1347569,I359738,I359841,I431643,I359867,I359875,I431655,I431634,I359892,I431658,I359918,I359809,I359940,I431649,I359966,I359974,I431631,I359991,I360017,I359833,I360039,I359815,I431646,I360079,I360096,I360104,I360121,I359818,I360152,I431637,I360169,I431640,I360195,I360203,I359806,I359824,I360248,I431652,I360265,I359827,I359812,I359821,I359830,I360368,I360394,I360402,I360419,I360445,I360336,I360467,I360493,I360501,I360518,I360544,I360360,I360566,I360342,I360606,I360623,I360631,I360648,I360345,I360679,I360696,I360722,I360730,I360333,I360351,I360775,I360792,I360354,I360339,I360348,I360357,I360895,I360921,I360929,I360946,I360972,I360994,I361020,I361028,I361045,I361071,I361093,I361133,I361150,I361158,I361175,I361206,I361223,I361249,I361257,I361302,I361319,I361422,I745174,I361448,I361456,I745165,I745180,I361473,I745186,I361499,I361390,I361521,I745171,I361547,I361555,I361572,I361598,I361414,I361620,I361396,I745168,I361660,I361677,I361685,I361702,I361399,I361733,I745162,I745177,I361750,I361776,I361784,I361387,I361405,I361829,I745183,I361846,I361408,I361393,I361402,I361411,I361949,I941192,I361975,I361983,I941189,I941207,I362000,I941198,I362026,I362048,I941213,I362074,I362082,I941195,I362099,I362125,I362147,I941201,I362187,I362204,I362212,I362229,I362260,I941216,I362277,I941204,I362303,I362311,I362356,I941210,I362373,I362476,I749798,I362502,I362510,I749789,I749804,I362527,I749810,I362553,I362444,I362575,I749795,I362601,I362609,I362626,I362652,I362468,I362674,I362450,I749792,I362714,I362731,I362739,I362756,I362453,I362787,I749786,I749801,I362804,I362830,I362838,I362441,I362459,I362883,I749807,I362900,I362462,I362447,I362456,I362465,I363003,I548079,I363029,I363037,I548064,I548067,I363054,I548082,I363080,I362971,I363102,I548076,I363128,I363136,I363153,I363179,I362995,I363201,I362977,I548073,I363241,I363258,I363266,I363283,I362980,I363314,I548088,I363331,I548085,I363357,I363365,I362968,I362986,I363410,I548070,I363427,I362989,I362974,I362983,I362992,I363530,I1108656,I363556,I363564,I1108671,I363581,I1108674,I363607,I363498,I363629,I1108680,I363655,I363663,I1108662,I363680,I363706,I363522,I363728,I363504,I1108659,I363768,I363785,I363793,I363810,I363507,I363841,I1108665,I363858,I1108677,I363884,I363892,I363495,I363513,I363937,I1108668,I363954,I363516,I363501,I363510,I363519,I364057,I1062416,I364083,I364091,I1062431,I364108,I1062434,I364134,I364025,I364156,I1062440,I364182,I364190,I1062422,I364207,I364233,I364049,I364255,I364031,I1062419,I364295,I364312,I364320,I364337,I364034,I364368,I1062425,I364385,I1062437,I364411,I364419,I364022,I364040,I364464,I1062428,I364481,I364043,I364028,I364037,I364046,I364584,I364610,I364618,I364635,I364661,I364552,I364683,I364709,I364717,I364734,I364760,I364576,I364782,I364558,I364822,I364839,I364847,I364864,I364561,I364895,I364912,I364938,I364946,I364549,I364567,I364991,I365008,I364570,I364555,I364564,I364573,I365111,I1386848,I365137,I365145,I1386827,I365162,I1386854,I365188,I365079,I365210,I1386842,I365236,I365244,I1386845,I365261,I365287,I365103,I365309,I365085,I1386836,I365349,I365366,I365374,I365391,I365088,I365422,I1386833,I1386830,I365439,I1386851,I365465,I365473,I365076,I365094,I365518,I1386839,I365535,I365097,I365082,I365091,I365100,I365638,I644602,I365664,I365672,I644593,I644608,I365689,I644614,I365715,I365737,I644599,I365763,I365771,I365788,I365814,I365836,I644596,I365876,I365893,I365901,I365918,I365949,I644590,I644605,I365966,I365992,I366000,I366045,I644611,I366062,I366165,I1184952,I366191,I366199,I1184967,I366216,I1184970,I366242,I366264,I1184976,I366290,I366298,I1184958,I366315,I366341,I366363,I1184955,I366403,I366420,I366428,I366445,I366476,I1184961,I366493,I1184973,I366519,I366527,I366572,I1184964,I366589,I366692,I1208532,I366718,I366726,I1208514,I1208538,I366743,I1208529,I366769,I366660,I366791,I1208535,I366817,I366825,I1208523,I366842,I366868,I366684,I366890,I366666,I366930,I366947,I366955,I366972,I366669,I367003,I1208520,I1208517,I367020,I1208526,I367046,I367054,I366657,I366675,I367099,I367116,I366678,I366663,I366672,I366681,I367219,I1195356,I367245,I367253,I1195371,I367270,I1195374,I367296,I367187,I367318,I1195380,I367344,I367352,I1195362,I367369,I367395,I367211,I367417,I367193,I1195359,I367457,I367474,I367482,I367499,I367196,I367530,I1195365,I367547,I1195377,I367573,I367581,I367184,I367202,I367626,I1195368,I367643,I367205,I367190,I367199,I367208,I367746,I770606,I367772,I367780,I770597,I770612,I367797,I770618,I367823,I367714,I367845,I770603,I367871,I367879,I367896,I367922,I367738,I367944,I367720,I770600,I367984,I368001,I368009,I368026,I367723,I368057,I770594,I770609,I368074,I368100,I368108,I367711,I367729,I368153,I770615,I368170,I367732,I367717,I367726,I367735,I368273,I1123106,I368299,I368307,I1123121,I368324,I1123124,I368350,I368241,I368372,I1123130,I368398,I368406,I1123112,I368423,I368449,I368265,I368471,I368247,I1123109,I368511,I368528,I368536,I368553,I368250,I368584,I1123115,I368601,I1123127,I368627,I368635,I368238,I368256,I368680,I1123118,I368697,I368259,I368244,I368253,I368262,I368800,I875504,I368826,I368834,I875507,I875501,I368851,I875513,I368877,I368768,I368899,I875516,I368925,I368933,I368950,I368976,I368792,I368998,I368774,I875519,I369038,I369055,I369063,I369080,I368777,I369111,I875510,I369128,I369154,I369162,I368765,I368783,I369207,I875522,I369224,I368786,I368771,I368780,I368789,I369327,I369353,I369361,I369378,I369404,I369295,I369426,I369452,I369460,I369477,I369503,I369319,I369525,I369301,I369565,I369582,I369590,I369607,I369304,I369638,I369655,I369681,I369689,I369292,I369310,I369734,I369751,I369313,I369298,I369307,I369316,I369854,I1069930,I369880,I369888,I1069945,I369905,I1069948,I369931,I369822,I369953,I1069954,I369979,I369987,I1069936,I370004,I370030,I369846,I370052,I369828,I1069933,I370092,I370109,I370117,I370134,I369831,I370165,I1069939,I370182,I1069951,I370208,I370216,I369819,I369837,I370261,I1069942,I370278,I369840,I369825,I369834,I369843,I370381,I1055024,I370407,I370415,I1055021,I370432,I1055033,I370458,I370480,I370506,I370514,I1055039,I370531,I370557,I370579,I1055027,I370619,I370636,I370644,I370661,I370692,I1055036,I1055042,I370709,I370735,I370743,I370788,I1055030,I370805,I370908,I627840,I370934,I370942,I627831,I627846,I370959,I627852,I370985,I370876,I371007,I627837,I371033,I371041,I371058,I371084,I370900,I371106,I370882,I627834,I371146,I371163,I371171,I371188,I370885,I371219,I627828,I627843,I371236,I371262,I371270,I370873,I370891,I371315,I627849,I371332,I370894,I370879,I370888,I370897,I371435,I1198246,I371461,I371469,I1198261,I371486,I1198264,I371512,I371403,I371534,I1198270,I371560,I371568,I1198252,I371585,I371611,I371427,I371633,I371409,I1198249,I371673,I371690,I371698,I371715,I371412,I371746,I1198255,I371763,I1198267,I371789,I371797,I371400,I371418,I371842,I1198258,I371859,I371421,I371406,I371415,I371424,I371962,I1298614,I371988,I371996,I1298641,I1298617,I372013,I1298626,I372039,I371930,I372061,I372087,I372095,I1298638,I372112,I372138,I371954,I372160,I371936,I1298620,I372200,I372217,I372225,I372242,I371939,I372273,I1298635,I1298623,I372290,I1298629,I372316,I372324,I371927,I371945,I372369,I1298632,I372386,I371948,I371933,I371942,I371951,I372489,I870234,I372515,I372523,I870237,I870231,I372540,I870243,I372566,I372457,I372588,I870246,I372614,I372622,I372639,I372665,I372481,I372687,I372463,I870249,I372727,I372744,I372752,I372769,I372466,I372800,I870240,I372817,I372843,I372851,I372454,I372472,I372896,I870252,I372913,I372475,I372460,I372469,I372478,I373016,I728412,I373042,I373050,I728403,I728418,I373067,I728424,I373093,I373115,I728409,I373141,I373149,I373166,I373192,I373214,I728406,I373254,I373271,I373279,I373296,I373327,I728400,I728415,I373344,I373370,I373378,I373423,I728421,I373440,I373543,I1037072,I373569,I373577,I1037069,I373594,I1037081,I373620,I373511,I373642,I373668,I373676,I1037087,I373693,I373719,I373535,I373741,I373517,I1037075,I373781,I373798,I373806,I373823,I373520,I373854,I1037084,I1037090,I373871,I373897,I373905,I373508,I373526,I373950,I1037078,I373967,I373529,I373514,I373523,I373532,I374070,I983828,I374096,I374104,I983825,I983843,I374121,I983834,I374147,I374038,I374169,I983849,I374195,I374203,I983831,I374220,I374246,I374062,I374268,I374044,I983837,I374308,I374325,I374333,I374350,I374047,I374381,I983852,I374398,I983840,I374424,I374432,I374035,I374053,I374477,I983846,I374494,I374056,I374041,I374050,I374059,I374597,I374623,I374631,I374648,I374674,I374565,I374696,I374722,I374730,I374747,I374773,I374589,I374795,I374571,I374835,I374852,I374860,I374877,I374574,I374908,I374925,I374951,I374959,I374562,I374580,I375004,I375021,I374583,I374568,I374577,I374586,I375124,I1308308,I375150,I375158,I1308287,I375175,I1308314,I375201,I375223,I1308302,I375249,I375257,I1308305,I375274,I375300,I375322,I1308296,I375362,I375379,I375387,I375404,I375435,I1308293,I1308290,I375452,I1308311,I375478,I375486,I375531,I1308299,I375548,I375651,I1124262,I375677,I375685,I1124277,I375702,I1124280,I375728,I375750,I1124286,I375776,I375784,I1124268,I375801,I375827,I375849,I1124265,I375889,I375906,I375914,I375931,I375962,I1124271,I375979,I1124283,I376005,I376013,I376058,I1124274,I376075,I376178,I376204,I376221,I376170,I376243,I376260,I376277,I376303,I376311,I376337,I376345,I376362,I376149,I376402,I376410,I376143,I376158,I376455,I376472,I376498,I376146,I376520,I376537,I376554,I376161,I376585,I376602,I376152,I376633,I376155,I376167,I376164,I376722,I961221,I376748,I376765,I376787,I376804,I961236,I961224,I376821,I961215,I376847,I376855,I961227,I376881,I376889,I961218,I376906,I961233,I376946,I376954,I376999,I961242,I961230,I377016,I961239,I377042,I377064,I377081,I377098,I377129,I377146,I377177,I377266,I1238437,I377292,I377309,I377331,I377348,I1238449,I1238452,I377365,I1238455,I377391,I377399,I1238440,I377425,I377433,I1238446,I377450,I1238434,I377490,I377498,I377543,I1238458,I377560,I1238443,I377586,I377608,I377625,I377642,I377673,I377690,I377721,I377810,I578123,I377836,I377853,I377802,I377875,I377892,I578120,I578141,I377909,I578144,I377935,I377943,I578129,I377969,I377977,I578132,I377994,I377781,I578135,I378034,I378042,I377775,I377790,I378087,I578126,I378104,I578138,I378130,I377778,I378152,I378169,I378186,I377793,I378217,I378234,I377784,I378265,I377787,I377799,I377796,I378354,I1213957,I378380,I378397,I378419,I378436,I1213969,I1213972,I378453,I1213975,I378479,I378487,I1213960,I378513,I378521,I1213966,I378538,I1213954,I378578,I378586,I378631,I1213978,I378648,I1213963,I378674,I378696,I378713,I378730,I378761,I378778,I378809,I378898,I863392,I378924,I378941,I378963,I378980,I863386,I863383,I378997,I863398,I379023,I379031,I379057,I379065,I863380,I379082,I379122,I379130,I379175,I863395,I863389,I379192,I379218,I379240,I379257,I379274,I379305,I379322,I863401,I379353,I379442,I1207973,I379468,I379485,I379434,I379507,I379524,I1207985,I1207988,I379541,I1207991,I379567,I379575,I1207976,I379601,I379609,I1207982,I379626,I379413,I1207970,I379666,I379674,I379407,I379422,I379719,I1207994,I379736,I1207979,I379762,I379410,I379784,I379801,I379818,I379425,I379849,I379866,I379416,I379897,I379419,I379431,I379428,I379986,I380012,I380029,I379978,I380051,I380068,I380085,I380111,I380119,I380145,I380153,I380170,I379957,I380210,I380218,I379951,I379966,I380263,I380280,I380306,I379954,I380328,I380345,I380362,I379969,I380393,I380410,I379960,I380441,I379963,I379975,I379972,I380530,I1249861,I380556,I380573,I380595,I380612,I1249873,I1249876,I380629,I1249879,I380655,I380663,I1249864,I380689,I380697,I1249870,I380714,I1249858,I380754,I380762,I380807,I1249882,I380824,I1249867,I380850,I380872,I380889,I380906,I380937,I380954,I380985,I381074,I1258240,I381100,I381117,I381066,I381139,I381156,I1258237,I1258234,I381173,I1258222,I381199,I381207,I1258246,I381233,I381241,I1258231,I381258,I381045,I1258225,I381298,I381306,I381039,I381054,I381351,I1258228,I381368,I1258243,I381394,I381042,I381416,I381433,I381450,I381057,I381481,I381498,I381048,I381529,I381051,I381063,I381060,I381618,I381644,I381661,I381683,I381700,I381717,I381743,I381751,I381777,I381785,I381802,I381842,I381850,I381895,I381912,I381938,I381960,I381977,I381994,I382025,I382042,I382073,I382162,I545755,I382188,I382205,I382227,I382244,I545752,I545773,I382261,I545776,I382287,I382295,I545761,I382321,I382329,I545764,I382346,I545767,I382386,I382394,I382439,I545758,I382456,I545770,I382482,I382504,I382521,I382538,I382569,I382586,I382617,I382706,I382732,I382749,I382698,I382771,I382788,I382805,I382831,I382839,I382865,I382873,I382890,I382677,I382930,I382938,I382671,I382686,I382983,I383000,I383026,I382674,I383048,I383065,I383082,I382689,I383113,I383130,I382680,I383161,I382683,I382695,I382692,I383250,I383276,I383293,I383242,I383315,I383332,I383349,I383375,I383383,I383409,I383417,I383434,I383221,I383474,I383482,I383215,I383230,I383527,I383544,I383570,I383218,I383592,I383609,I383626,I383233,I383657,I383674,I383224,I383705,I383227,I383239,I383236,I383794,I1259974,I383820,I383837,I383859,I383876,I1259971,I1259968,I383893,I1259956,I383919,I383927,I1259980,I383953,I383961,I1259965,I383978,I1259959,I384018,I384026,I384071,I1259962,I384088,I1259977,I384114,I384136,I384153,I384170,I384201,I384218,I384249,I384338,I1108081,I384364,I384381,I384403,I384420,I1108093,I384437,I1108084,I384463,I384471,I1108102,I384497,I384505,I1108078,I384522,I1108096,I384562,I384570,I384615,I1108090,I1108087,I384632,I1108099,I384658,I384680,I384697,I384714,I384745,I384762,I384793,I384882,I384908,I384925,I384874,I384947,I384964,I384981,I385007,I385015,I385041,I385049,I385066,I384853,I385106,I385114,I384847,I384862,I385159,I385176,I385202,I384850,I385224,I385241,I385258,I384865,I385289,I385306,I384856,I385337,I384859,I384871,I384868,I385426,I1363649,I385452,I385469,I385418,I385491,I385508,I1363625,I1363646,I385525,I1363643,I385551,I385559,I1363622,I385585,I385593,I1363634,I385610,I385397,I1363637,I385650,I385658,I385391,I385406,I385703,I1363640,I1363628,I385720,I1363631,I385746,I385394,I385768,I385785,I385802,I385409,I385833,I385850,I385400,I385881,I385403,I385415,I385412,I385970,I819651,I385996,I386013,I386035,I386052,I819645,I819642,I386069,I819657,I386095,I386103,I386129,I386137,I819639,I386154,I386194,I386202,I386247,I819654,I819648,I386264,I386290,I386312,I386329,I386346,I386377,I386394,I819660,I386425,I386514,I386540,I386557,I386506,I386579,I386596,I386613,I386639,I386647,I386673,I386681,I386698,I386485,I386738,I386746,I386479,I386494,I386791,I386808,I386834,I386482,I386856,I386873,I386890,I386497,I386921,I386938,I386488,I386969,I386491,I386503,I386500,I387058,I1060107,I387084,I387101,I387123,I387140,I1060119,I387157,I1060110,I387183,I387191,I1060128,I387217,I387225,I1060104,I387242,I1060122,I387282,I387290,I387335,I1060116,I1060113,I387352,I1060125,I387378,I387400,I387417,I387434,I387465,I387482,I387513,I387602,I387628,I387645,I387594,I387667,I387684,I387701,I387727,I387735,I387761,I387769,I387786,I387573,I387826,I387834,I387567,I387582,I387879,I387896,I387922,I387570,I387944,I387961,I387978,I387585,I388009,I388026,I387576,I388057,I387579,I387591,I387588,I388146,I1275580,I388172,I388189,I388211,I388228,I1275577,I1275574,I388245,I1275562,I388271,I388279,I1275586,I388305,I388313,I1275571,I388330,I1275565,I388370,I388378,I388423,I1275568,I388440,I1275583,I388466,I388488,I388505,I388522,I388553,I388570,I388601,I388690,I939257,I388716,I388733,I388755,I388772,I939272,I939260,I388789,I939251,I388815,I388823,I939263,I388849,I388857,I939254,I388874,I939269,I388914,I388922,I388967,I939278,I939266,I388984,I939275,I389010,I389032,I389049,I389066,I389097,I389114,I389145,I389234,I389260,I389277,I389226,I389299,I389316,I389333,I389359,I389367,I389393,I389401,I389418,I389205,I389458,I389466,I389199,I389214,I389511,I389528,I389554,I389202,I389576,I389593,I389610,I389217,I389641,I389658,I389208,I389689,I389211,I389223,I389220,I389778,I389804,I389821,I389770,I389843,I389860,I389877,I389903,I389911,I389937,I389945,I389962,I389749,I390002,I390010,I389743,I389758,I390055,I390072,I390098,I389746,I390120,I390137,I390154,I389761,I390185,I390202,I389752,I390233,I389755,I389767,I389764,I390322,I390348,I390365,I390387,I390404,I390421,I390447,I390455,I390481,I390489,I390506,I390546,I390554,I390599,I390616,I390642,I390664,I390681,I390698,I390729,I390746,I390777,I390866,I912771,I390892,I390909,I390858,I390931,I390948,I912786,I912774,I390965,I912765,I390991,I390999,I912777,I391025,I391033,I912768,I391050,I390837,I912783,I391090,I391098,I390831,I390846,I391143,I912792,I912780,I391160,I912789,I391186,I390834,I391208,I391225,I391242,I390849,I391273,I391290,I390840,I391321,I390843,I390855,I390852,I391410,I1302556,I391436,I391453,I391475,I391492,I1302562,I1302565,I391509,I1302541,I391535,I391543,I1302568,I391569,I391577,I1302550,I391594,I1302547,I391634,I391642,I391687,I1302544,I1302553,I391704,I1302559,I391730,I391752,I391769,I391786,I391817,I391834,I391865,I391954,I745743,I391980,I391997,I391946,I392019,I392036,I745764,I745755,I392053,I392079,I392087,I745749,I392113,I392121,I745746,I392138,I391925,I745740,I392178,I392186,I391919,I391934,I392231,I745752,I392248,I745761,I392274,I391922,I392296,I392313,I392330,I391937,I392361,I392378,I745758,I391928,I392409,I391931,I391943,I391940,I392498,I582747,I392524,I392541,I392563,I392580,I582744,I582765,I392597,I582768,I392623,I392631,I582753,I392657,I392665,I582756,I392682,I582759,I392722,I392730,I392775,I582750,I392792,I582762,I392818,I392840,I392857,I392874,I392905,I392922,I392953,I393042,I667135,I393068,I393085,I393034,I393107,I393124,I667156,I667147,I393141,I393167,I393175,I667141,I393201,I393209,I667138,I393226,I393013,I667132,I393266,I393274,I393007,I393022,I393319,I667144,I393336,I667153,I393362,I393010,I393384,I393401,I393418,I393025,I393449,I393466,I667150,I393016,I393497,I393019,I393031,I393028,I393586,I1120797,I393612,I393629,I393578,I393651,I393668,I1120809,I393685,I1120800,I393711,I393719,I1120818,I393745,I393753,I1120794,I393770,I393557,I1120812,I393810,I393818,I393551,I393566,I393863,I1120806,I1120803,I393880,I1120815,I393906,I393554,I393928,I393945,I393962,I393569,I393993,I394010,I393560,I394041,I393563,I393575,I393572,I394130,I970265,I394156,I394173,I394195,I394212,I970280,I970268,I394229,I970259,I394255,I394263,I970271,I394289,I394297,I970262,I394314,I970277,I394354,I394362,I394407,I970286,I970274,I394424,I970283,I394450,I394472,I394489,I394506,I394537,I394554,I394585,I394674,I1357104,I394700,I394717,I394739,I394756,I1357080,I1357101,I394773,I1357098,I394799,I394807,I1357077,I394833,I394841,I1357089,I394858,I1357092,I394898,I394906,I394951,I1357095,I1357083,I394968,I1357086,I394994,I395016,I395033,I395050,I395081,I395098,I395129,I395218,I735339,I395244,I395261,I395283,I395300,I735360,I735351,I395317,I395343,I395351,I735345,I395377,I395385,I735342,I395402,I735336,I395442,I395450,I395495,I735348,I395512,I735357,I395538,I395560,I395577,I395594,I395625,I395642,I735354,I395673,I395762,I939903,I395788,I395805,I395754,I395827,I395844,I939918,I939906,I395861,I939897,I395887,I395895,I939909,I395921,I395929,I939900,I395946,I395733,I939915,I395986,I395994,I395727,I395742,I396039,I939924,I939912,I396056,I939921,I396082,I395730,I396104,I396121,I396138,I395745,I396169,I396186,I395736,I396217,I395739,I395751,I395748,I396306,I1139871,I396332,I396349,I396298,I396371,I396388,I1139883,I396405,I1139874,I396431,I396439,I1139892,I396465,I396473,I1139868,I396490,I396277,I1139886,I396530,I396538,I396271,I396286,I396583,I1139880,I1139877,I396600,I1139889,I396626,I396274,I396648,I396665,I396682,I396289,I396713,I396730,I396280,I396761,I396283,I396295,I396292,I396850,I985123,I396876,I396893,I396842,I396915,I396932,I985138,I985126,I396949,I985117,I396975,I396983,I985129,I397009,I397017,I985120,I397034,I396821,I985135,I397074,I397082,I396815,I396830,I397127,I985144,I985132,I397144,I985141,I397170,I396818,I397192,I397209,I397226,I396833,I397257,I397274,I396824,I397305,I396827,I396839,I396836,I397394,I397420,I397437,I397386,I397459,I397476,I397493,I397519,I397527,I397553,I397561,I397578,I397365,I397618,I397626,I397359,I397374,I397671,I397688,I397714,I397362,I397736,I397753,I397770,I397377,I397801,I397818,I397368,I397849,I397371,I397383,I397380,I397938,I706439,I397964,I397981,I398003,I398020,I706460,I706451,I398037,I398063,I398071,I706445,I398097,I398105,I706442,I398122,I706436,I398162,I398170,I398215,I706448,I398232,I706457,I398258,I398280,I398297,I398314,I398345,I398362,I706454,I398393,I398482,I1390424,I398508,I398525,I398474,I398547,I398564,I1390400,I1390421,I398581,I1390418,I398607,I398615,I1390397,I398641,I398649,I1390409,I398666,I398453,I1390412,I398706,I398714,I398447,I398462,I398759,I1390415,I1390403,I398776,I1390406,I398802,I398450,I398824,I398841,I398858,I398465,I398889,I398906,I398456,I398937,I398459,I398471,I398468,I399026,I752679,I399052,I399069,I399091,I399108,I752700,I752691,I399125,I399151,I399159,I752685,I399185,I399193,I752682,I399210,I752676,I399250,I399258,I399303,I752688,I399320,I752697,I399346,I399368,I399385,I399402,I399433,I399450,I752694,I399481,I399570,I881310,I399596,I399613,I399562,I399635,I399652,I881304,I881301,I399669,I881316,I399695,I399703,I399729,I399737,I881298,I399754,I399541,I399794,I399802,I399535,I399550,I399847,I881313,I881307,I399864,I399890,I399538,I399912,I399929,I399946,I399553,I399977,I399994,I881319,I399544,I400025,I399547,I399559,I399556,I400114,I937319,I400140,I400157,I400106,I400179,I400196,I937334,I937322,I400213,I937313,I400239,I400247,I937325,I400273,I400281,I937316,I400298,I400085,I937331,I400338,I400346,I400079,I400094,I400391,I937340,I937328,I400408,I937337,I400434,I400082,I400456,I400473,I400490,I400097,I400521,I400538,I400088,I400569,I400091,I400103,I400100,I400658,I1029215,I400684,I400701,I400723,I400740,I1029233,I400757,I1029227,I400783,I400791,I1029221,I400817,I400825,I1029230,I400842,I1029218,I400882,I400890,I400935,I1029236,I400952,I400978,I401000,I401017,I401034,I401065,I401082,I1029224,I401113,I401202,I401228,I401245,I401194,I401267,I401284,I401301,I401327,I401335,I401361,I401369,I401386,I401173,I401426,I401434,I401167,I401182,I401479,I401496,I401522,I401170,I401544,I401561,I401578,I401185,I401609,I401626,I401176,I401657,I401179,I401191,I401188,I401746,I1201139,I401772,I401789,I401738,I401811,I401828,I1201151,I401845,I1201142,I401871,I401879,I1201160,I401905,I401913,I1201136,I401930,I401717,I1201154,I401970,I401978,I401711,I401726,I402023,I1201148,I1201145,I402040,I1201157,I402066,I401714,I402088,I402105,I402122,I401729,I402153,I402170,I401720,I402201,I401723,I401735,I401732,I402290,I402316,I402333,I402282,I402355,I402372,I402389,I402415,I402423,I402449,I402457,I402474,I402261,I402514,I402522,I402255,I402270,I402567,I402584,I402610,I402258,I402632,I402649,I402666,I402273,I402697,I402714,I402264,I402745,I402267,I402279,I402276,I402834,I1217765,I402860,I402877,I402826,I402899,I402916,I1217777,I1217780,I402933,I1217783,I402959,I402967,I1217768,I402993,I403001,I1217774,I403018,I402805,I1217762,I403058,I403066,I402799,I402814,I403111,I1217786,I403128,I1217771,I403154,I402802,I403176,I403193,I403210,I402817,I403241,I403258,I402808,I403289,I402811,I402823,I402820,I403378,I879202,I403404,I403421,I403370,I403443,I403460,I879196,I879193,I403477,I879208,I403503,I403511,I403537,I403545,I879190,I403562,I403349,I403602,I403610,I403343,I403358,I403655,I879205,I879199,I403672,I403698,I403346,I403720,I403737,I403754,I403361,I403785,I403802,I879211,I403352,I403833,I403355,I403367,I403364,I403922,I554425,I403948,I403965,I403914,I403987,I404004,I554422,I554443,I404021,I554446,I404047,I404055,I554431,I404081,I404089,I554434,I404106,I403893,I554437,I404146,I404154,I403887,I403902,I404199,I554428,I404216,I554440,I404242,I403890,I404264,I404281,I404298,I403905,I404329,I404346,I403896,I404377,I403899,I403911,I403908,I404466,I947655,I404492,I404509,I404458,I404531,I404548,I947670,I947658,I404565,I947649,I404591,I404599,I947661,I404625,I404633,I947652,I404650,I404437,I947667,I404690,I404698,I404431,I404446,I404743,I947676,I947664,I404760,I947673,I404786,I404434,I404808,I404825,I404842,I404449,I404873,I404890,I404440,I404921,I404443,I404455,I404452,I405010,I405036,I405053,I405002,I405075,I405092,I405109,I405135,I405143,I405169,I405177,I405194,I404981,I405234,I405242,I404975,I404990,I405287,I405304,I405330,I404978,I405352,I405369,I405386,I404993,I405417,I405434,I404984,I405465,I404987,I404999,I404996,I405554,I405580,I405597,I405546,I405619,I405636,I405653,I405679,I405687,I405713,I405721,I405738,I405525,I405778,I405786,I405519,I405534,I405831,I405848,I405874,I405522,I405896,I405913,I405930,I405537,I405961,I405978,I405528,I406009,I405531,I405543,I405540,I406098,I683897,I406124,I406141,I406090,I406163,I406180,I683918,I683909,I406197,I406223,I406231,I683903,I406257,I406265,I683900,I406282,I406069,I683894,I406322,I406330,I406063,I406078,I406375,I683906,I406392,I683915,I406418,I406066,I406440,I406457,I406474,I406081,I406505,I406522,I683912,I406072,I406553,I406075,I406087,I406084,I406642,I406668,I406685,I406634,I406707,I406724,I406741,I406767,I406775,I406801,I406809,I406826,I406613,I406866,I406874,I406607,I406622,I406919,I406936,I406962,I406610,I406984,I407001,I407018,I406625,I407049,I407066,I406616,I407097,I406619,I406631,I406628,I407186,I1080915,I407212,I407229,I407178,I407251,I407268,I1080927,I407285,I1080918,I407311,I407319,I1080936,I407345,I407353,I1080912,I407370,I407157,I1080930,I407410,I407418,I407151,I407166,I407463,I1080924,I1080921,I407480,I1080933,I407506,I407154,I407528,I407545,I407562,I407169,I407593,I407610,I407160,I407641,I407163,I407175,I407172,I407730,I517892,I407756,I407773,I407722,I407795,I407812,I517895,I517913,I407829,I517901,I407855,I407863,I407889,I407897,I517910,I407914,I407701,I517904,I407954,I407962,I407695,I407710,I408007,I517907,I517889,I408024,I517898,I408050,I407698,I408072,I408089,I408106,I407713,I408137,I408154,I407704,I408185,I407707,I407719,I407716,I408274,I1380309,I408300,I408317,I408266,I408339,I408356,I1380285,I1380306,I408373,I1380303,I408399,I408407,I1380282,I408433,I408441,I1380294,I408458,I408245,I1380297,I408498,I408506,I408239,I408254,I408551,I1380300,I1380288,I408568,I1380291,I408594,I408242,I408616,I408633,I408650,I408257,I408681,I408698,I408248,I408729,I408251,I408263,I408260,I408818,I408844,I408861,I408810,I408883,I408900,I408917,I408943,I408951,I408977,I408985,I409002,I408789,I409042,I409050,I408783,I408798,I409095,I409112,I409138,I408786,I409160,I409177,I409194,I408801,I409225,I409242,I408792,I409273,I408795,I408807,I408804,I409362,I801206,I409388,I409405,I409354,I409427,I409444,I801200,I801197,I409461,I801212,I409487,I409495,I409521,I409529,I801194,I409546,I409333,I409586,I409594,I409327,I409342,I409639,I801209,I801203,I409656,I409682,I409330,I409704,I409721,I409738,I409345,I409769,I409786,I801215,I409336,I409817,I409339,I409351,I409348,I409906,I409932,I409949,I409898,I409971,I409988,I410005,I410031,I410039,I410065,I410073,I410090,I409877,I410130,I410138,I409871,I409886,I410183,I410200,I410226,I409874,I410248,I410265,I410282,I409889,I410313,I410330,I409880,I410361,I409883,I409895,I409892,I410450,I1234629,I410476,I410493,I410442,I410515,I410532,I1234641,I1234644,I410549,I1234647,I410575,I410583,I1234632,I410609,I410617,I1234638,I410634,I410421,I1234626,I410674,I410682,I410415,I410430,I410727,I1234650,I410744,I1234635,I410770,I410418,I410792,I410809,I410826,I410433,I410857,I410874,I410424,I410905,I410427,I410439,I410436,I410994,I1143917,I411020,I411037,I411059,I411076,I1143929,I411093,I1143920,I411119,I411127,I1143938,I411153,I411161,I1143914,I411178,I1143932,I411218,I411226,I411271,I1143926,I1143923,I411288,I1143935,I411314,I411336,I411353,I411370,I411401,I411418,I411449,I411538,I1101145,I411564,I411581,I411603,I411620,I1101157,I411637,I1101148,I411663,I411671,I1101166,I411697,I411705,I1101142,I411722,I1101160,I411762,I411770,I411815,I1101154,I1101151,I411832,I1101163,I411858,I411880,I411897,I411914,I411945,I411962,I411993,I412082,I412108,I412125,I412147,I412164,I412181,I412207,I412215,I412241,I412249,I412266,I412306,I412314,I412359,I412376,I412402,I412424,I412441,I412458,I412489,I412506,I412537,I412626,I412652,I412669,I412618,I412691,I412708,I412725,I412751,I412759,I412785,I412793,I412810,I412597,I412850,I412858,I412591,I412606,I412903,I412920,I412946,I412594,I412968,I412985,I413002,I412609,I413033,I413050,I412600,I413081,I412603,I412615,I412612,I413170,I1255350,I413196,I413213,I413162,I413235,I413252,I1255347,I1255344,I413269,I1255332,I413295,I413303,I1255356,I413329,I413337,I1255341,I413354,I413141,I1255335,I413394,I413402,I413135,I413150,I413447,I1255338,I413464,I1255353,I413490,I413138,I413512,I413529,I413546,I413153,I413577,I413594,I413144,I413625,I413147,I413159,I413156,I413714,I1373764,I413740,I413757,I413779,I413796,I1373740,I1373761,I413813,I1373758,I413839,I413847,I1373737,I413873,I413881,I1373749,I413898,I1373752,I413938,I413946,I413991,I1373755,I1373743,I414008,I1373746,I414034,I414056,I414073,I414090,I414121,I414138,I414169,I414258,I414284,I414301,I414250,I414323,I414340,I414357,I414383,I414391,I414417,I414425,I414442,I414229,I414482,I414490,I414223,I414238,I414535,I414552,I414578,I414226,I414600,I414617,I414634,I414241,I414665,I414682,I414232,I414713,I414235,I414247,I414244,I414802,I1106347,I414828,I414845,I414867,I414884,I1106359,I414901,I1106350,I414927,I414935,I1106368,I414961,I414969,I1106344,I414986,I1106362,I415026,I415034,I415079,I1106356,I1106353,I415096,I1106365,I415122,I415144,I415161,I415178,I415209,I415226,I415257,I415346,I1237893,I415372,I415389,I415338,I415411,I415428,I1237905,I1237908,I415445,I1237911,I415471,I415479,I1237896,I415505,I415513,I1237902,I415530,I415317,I1237890,I415570,I415578,I415311,I415326,I415623,I1237914,I415640,I1237899,I415666,I415314,I415688,I415705,I415722,I415329,I415753,I415770,I415320,I415801,I415323,I415335,I415332,I415890,I860757,I415916,I415933,I415955,I415972,I860751,I860748,I415989,I860763,I416015,I416023,I416049,I416057,I860745,I416074,I416114,I416122,I416167,I860760,I860754,I416184,I416210,I416232,I416249,I416266,I416297,I416314,I860766,I416345,I416434,I685631,I416460,I416477,I416426,I416499,I416516,I685652,I685643,I416533,I416559,I416567,I685637,I416593,I416601,I685634,I416618,I416405,I685628,I416658,I416666,I416399,I416414,I416711,I685640,I416728,I685649,I416754,I416402,I416776,I416793,I416810,I416417,I416841,I416858,I685646,I416408,I416889,I416411,I416423,I416420,I416978,I1374954,I417004,I417021,I416970,I417043,I417060,I1374930,I1374951,I417077,I1374948,I417103,I417111,I1374927,I417137,I417145,I1374939,I417162,I416949,I1374942,I417202,I417210,I416943,I416958,I417255,I1374945,I1374933,I417272,I1374936,I417298,I416946,I417320,I417337,I417354,I416961,I417385,I417402,I416952,I417433,I416955,I416967,I416964,I417522,I736495,I417548,I417565,I417514,I417587,I417604,I736516,I736507,I417621,I417647,I417655,I736501,I417681,I417689,I736498,I417706,I417493,I736492,I417746,I417754,I417487,I417502,I417799,I736504,I417816,I736513,I417842,I417490,I417864,I417881,I417898,I417505,I417929,I417946,I736510,I417496,I417977,I417499,I417511,I417508,I418066,I815962,I418092,I418109,I418131,I418148,I815956,I815953,I418165,I815968,I418191,I418199,I418225,I418233,I815950,I418250,I418290,I418298,I418343,I815965,I815959,I418360,I418386,I418408,I418425,I418442,I418473,I418490,I815971,I418521,I418610,I418636,I418653,I418602,I418675,I418692,I418709,I418735,I418743,I418769,I418777,I418794,I418581,I418834,I418842,I418575,I418590,I418887,I418904,I418930,I418578,I418952,I418969,I418986,I418593,I419017,I419034,I418584,I419065,I418587,I418599,I418596,I419154,I1023605,I419180,I419197,I419219,I419236,I1023623,I419253,I1023617,I419279,I419287,I1023611,I419313,I419321,I1023620,I419338,I1023608,I419378,I419386,I419431,I1023626,I419448,I419474,I419496,I419513,I419530,I419561,I419578,I1023614,I419609,I419698,I597197,I419724,I419741,I419690,I419763,I419780,I597194,I597215,I419797,I597218,I419823,I419831,I597203,I419857,I419865,I597206,I419882,I419669,I597209,I419922,I419930,I419663,I419678,I419975,I597200,I419992,I597212,I420018,I419666,I420040,I420057,I420074,I419681,I420105,I420122,I419672,I420153,I419675,I419687,I419684,I420242,I1154321,I420268,I420285,I420234,I420307,I420324,I1154333,I420341,I1154324,I420367,I420375,I1154342,I420401,I420409,I1154318,I420426,I420213,I1154336,I420466,I420474,I420207,I420222,I420519,I1154330,I1154327,I420536,I1154339,I420562,I420210,I420584,I420601,I420618,I420225,I420649,I420666,I420216,I420697,I420219,I420231,I420228,I420786,I420812,I420829,I420778,I420851,I420868,I420885,I420911,I420919,I420945,I420953,I420970,I420757,I421010,I421018,I420751,I420766,I421063,I421080,I421106,I420754,I421128,I421145,I421162,I420769,I421193,I421210,I420760,I421241,I420763,I420775,I420772,I421330,I855487,I421356,I421373,I421322,I421395,I421412,I855481,I855478,I421429,I855493,I421455,I421463,I421489,I421497,I855475,I421514,I421301,I421554,I421562,I421295,I421310,I421607,I855490,I855484,I421624,I421650,I421298,I421672,I421689,I421706,I421313,I421737,I421754,I855496,I421304,I421785,I421307,I421319,I421316,I421874,I421900,I421917,I421866,I421939,I421956,I421973,I421999,I422007,I422033,I422041,I422058,I421845,I422098,I422106,I421839,I421854,I422151,I422168,I422194,I421842,I422216,I422233,I422250,I421857,I422281,I422298,I421848,I422329,I421851,I421863,I421860,I422418,I602399,I422444,I422461,I422410,I422483,I422500,I602396,I602417,I422517,I602420,I422543,I422551,I602405,I422577,I422585,I602408,I422602,I422389,I602411,I422642,I422650,I422383,I422398,I422695,I602402,I422712,I602414,I422738,I422386,I422760,I422777,I422794,I422401,I422825,I422842,I422392,I422873,I422395,I422407,I422404,I422962,I1076291,I422988,I423005,I422954,I423027,I423044,I1076303,I423061,I1076294,I423087,I423095,I1076312,I423121,I423129,I1076288,I423146,I422933,I1076306,I423186,I423194,I422927,I422942,I423239,I1076300,I1076297,I423256,I1076309,I423282,I422930,I423304,I423321,I423338,I422945,I423369,I423386,I422936,I423417,I422939,I422951,I422948,I423506,I581591,I423532,I423549,I423498,I423571,I423588,I581588,I581609,I423605,I581612,I423631,I423639,I581597,I423665,I423673,I581600,I423690,I423477,I581603,I423730,I423738,I423471,I423486,I423783,I581594,I423800,I581606,I423826,I423474,I423848,I423865,I423882,I423489,I423913,I423930,I423480,I423961,I423483,I423495,I423492,I424050,I1355319,I424076,I424093,I424042,I424115,I424132,I1355295,I1355316,I424149,I1355313,I424175,I424183,I1355292,I424209,I424217,I1355304,I424234,I424021,I1355307,I424274,I424282,I424015,I424030,I424327,I1355310,I1355298,I424344,I1355301,I424370,I424018,I424392,I424409,I424426,I424033,I424457,I424474,I424024,I424505,I424027,I424039,I424036,I424594,I1221573,I424620,I424637,I424586,I424659,I424676,I1221585,I1221588,I424693,I1221591,I424719,I424727,I1221576,I424753,I424761,I1221582,I424778,I424565,I1221570,I424818,I424826,I424559,I424574,I424871,I1221594,I424888,I1221579,I424914,I424562,I424936,I424953,I424970,I424577,I425001,I425018,I424568,I425049,I424571,I424583,I424580,I425138,I856014,I425164,I425181,I425130,I425203,I425220,I856008,I856005,I425237,I856020,I425263,I425271,I425297,I425305,I856002,I425322,I425109,I425362,I425370,I425103,I425118,I425415,I856017,I856011,I425432,I425458,I425106,I425480,I425497,I425514,I425121,I425545,I425562,I856023,I425112,I425593,I425115,I425127,I425124,I425682,I716265,I425708,I425725,I425674,I425747,I425764,I716286,I716277,I425781,I425807,I425815,I716271,I425841,I425849,I716268,I425866,I425653,I716262,I425906,I425914,I425647,I425662,I425959,I716274,I425976,I716283,I426002,I425650,I426024,I426041,I426058,I425665,I426089,I426106,I716280,I425656,I426137,I425659,I425671,I425668,I426226,I759615,I426252,I426269,I426218,I426291,I426308,I759636,I759627,I426325,I426351,I426359,I759621,I426385,I426393,I759618,I426410,I426197,I759612,I426450,I426458,I426191,I426206,I426503,I759624,I426520,I759633,I426546,I426194,I426568,I426585,I426602,I426209,I426633,I426650,I759630,I426200,I426681,I426203,I426215,I426212,I426770,I426796,I426813,I426762,I426835,I426852,I426869,I426895,I426903,I426929,I426937,I426954,I426741,I426994,I427002,I426735,I426750,I427047,I427064,I427090,I426738,I427112,I427129,I427146,I426753,I427177,I427194,I426744,I427225,I426747,I426759,I426756,I427314,I1366029,I427340,I427357,I427306,I427379,I427396,I1366005,I1366026,I427413,I1366023,I427439,I427447,I1366002,I427473,I427481,I1366014,I427498,I427285,I1366017,I427538,I427546,I427279,I427294,I427591,I1366020,I1366008,I427608,I1366011,I427634,I427282,I427656,I427673,I427690,I427297,I427721,I427738,I427288,I427769,I427291,I427303,I427300,I427858,I427884,I427901,I427850,I427923,I427940,I427957,I427983,I427991,I428017,I428025,I428042,I427829,I428082,I428090,I427823,I427838,I428135,I428152,I428178,I427826,I428200,I428217,I428234,I427841,I428265,I428282,I427832,I428313,I427835,I427847,I427844,I428402,I428428,I428445,I428394,I428467,I428484,I428501,I428527,I428535,I428561,I428569,I428586,I428373,I428626,I428634,I428367,I428382,I428679,I428696,I428722,I428370,I428744,I428761,I428778,I428385,I428809,I428826,I428376,I428857,I428379,I428391,I428388,I428946,I746899,I428972,I428989,I428938,I429011,I429028,I746920,I746911,I429045,I429071,I429079,I746905,I429105,I429113,I746902,I429130,I428917,I746896,I429170,I429178,I428911,I428926,I429223,I746908,I429240,I746917,I429266,I428914,I429288,I429305,I429322,I428929,I429353,I429370,I746914,I428920,I429401,I428923,I428935,I428932,I429490,I1354724,I429516,I429533,I429482,I429555,I429572,I1354700,I1354721,I429589,I1354718,I429615,I429623,I1354697,I429649,I429657,I1354709,I429674,I429461,I1354712,I429714,I429722,I429455,I429470,I429767,I1354715,I1354703,I429784,I1354706,I429810,I429458,I429832,I429849,I429866,I429473,I429897,I429914,I429464,I429945,I429467,I429479,I429476,I430034,I560783,I430060,I430077,I430099,I430116,I560780,I560801,I430133,I560804,I430159,I430167,I560789,I430193,I430201,I560792,I430218,I560795,I430258,I430266,I430311,I560786,I430328,I560798,I430354,I430376,I430393,I430410,I430441,I430458,I430489,I430578,I717999,I430604,I430621,I430570,I430643,I430660,I718020,I718011,I430677,I430703,I430711,I718005,I430737,I430745,I718002,I430762,I430549,I717996,I430802,I430810,I430543,I430558,I430855,I718008,I430872,I718017,I430898,I430546,I430920,I430937,I430954,I430561,I430985,I431002,I718014,I430552,I431033,I430555,I430567,I430564,I431122,I1158367,I431148,I431165,I431114,I431187,I431204,I1158379,I431221,I1158370,I431247,I431255,I1158388,I431281,I431289,I1158364,I431306,I431093,I1158382,I431346,I431354,I431087,I431102,I431399,I1158376,I1158373,I431416,I1158385,I431442,I431090,I431464,I431481,I431498,I431105,I431529,I431546,I431096,I431577,I431099,I431111,I431108,I431666,I431692,I431709,I431731,I431748,I431765,I431791,I431799,I431825,I431833,I431850,I431890,I431898,I431943,I431960,I431986,I432008,I432025,I432042,I432073,I432090,I432121,I432210,I432236,I432253,I432202,I432275,I432292,I432309,I432335,I432343,I432369,I432377,I432394,I432181,I432434,I432442,I432175,I432190,I432487,I432504,I432530,I432178,I432552,I432569,I432586,I432193,I432617,I432634,I432184,I432665,I432187,I432199,I432196,I432754,I1125999,I432780,I432797,I432746,I432819,I432836,I1126011,I432853,I1126002,I432879,I432887,I1126020,I432913,I432921,I1125996,I432938,I432725,I1126014,I432978,I432986,I432719,I432734,I433031,I1126008,I1126005,I433048,I1126017,I433074,I432722,I433096,I433113,I433130,I432737,I433161,I433178,I432728,I433209,I432731,I432743,I432740,I433298,I782761,I433324,I433341,I433290,I433363,I433380,I782755,I782752,I433397,I782767,I433423,I433431,I433457,I433465,I782749,I433482,I433269,I433522,I433530,I433263,I433278,I433575,I782764,I782758,I433592,I433618,I433266,I433640,I433657,I433674,I433281,I433705,I433722,I782770,I433272,I433753,I433275,I433287,I433284,I433842,I1307124,I433868,I433885,I433834,I433907,I433924,I1307100,I1307121,I433941,I1307118,I433967,I433975,I1307097,I434001,I434009,I1307109,I434026,I433813,I1307112,I434066,I434074,I433807,I433822,I434119,I1307115,I1307103,I434136,I1307106,I434162,I433810,I434184,I434201,I434218,I433825,I434249,I434266,I433816,I434297,I433819,I433831,I433828,I434386,I434412,I434429,I434378,I434451,I434468,I434485,I434511,I434519,I434545,I434553,I434570,I434357,I434610,I434618,I434351,I434366,I434663,I434680,I434706,I434354,I434728,I434745,I434762,I434369,I434793,I434810,I434360,I434841,I434363,I434375,I434372,I434930,I967035,I434956,I434973,I434922,I434995,I435012,I967050,I967038,I435029,I967029,I435055,I435063,I967041,I435089,I435097,I967032,I435114,I434901,I967047,I435154,I435162,I434895,I434910,I435207,I967056,I967044,I435224,I967053,I435250,I434898,I435272,I435289,I435306,I434913,I435337,I435354,I434904,I435385,I434907,I434919,I434916,I435474,I1223205,I435500,I435517,I435466,I435539,I435556,I1223217,I1223220,I435573,I1223223,I435599,I435607,I1223208,I435633,I435641,I1223214,I435658,I435445,I1223202,I435698,I435706,I435439,I435454,I435751,I1223226,I435768,I1223211,I435794,I435442,I435816,I435833,I435850,I435457,I435881,I435898,I435448,I435929,I435451,I435463,I435460,I436018,I1389829,I436044,I436061,I436010,I436083,I436100,I1389805,I1389826,I436117,I1389823,I436143,I436151,I1389802,I436177,I436185,I1389814,I436202,I435989,I1389817,I436242,I436250,I435983,I435998,I436295,I1389820,I1389808,I436312,I1389811,I436338,I435986,I436360,I436377,I436394,I436001,I436425,I436442,I435992,I436473,I435995,I436007,I436004,I436562,I1194781,I436588,I436605,I436627,I436644,I1194793,I436661,I1194784,I436687,I436695,I1194802,I436721,I436729,I1194778,I436746,I1194796,I436786,I436794,I436839,I1194790,I1194787,I436856,I1194799,I436882,I436904,I436921,I436938,I436969,I436986,I437017,I437106,I437132,I437149,I437098,I437171,I437188,I437205,I437231,I437239,I437265,I437273,I437290,I437077,I437330,I437338,I437071,I437086,I437383,I437400,I437426,I437074,I437448,I437465,I437482,I437089,I437513,I437530,I437080,I437561,I437083,I437095,I437092,I437650,I781707,I437676,I437693,I437642,I437715,I437732,I781701,I781698,I437749,I781713,I437775,I437783,I437809,I437817,I781695,I437834,I437621,I437874,I437882,I437615,I437630,I437927,I781710,I781704,I437944,I437970,I437618,I437992,I438009,I438026,I437633,I438057,I438074,I781716,I437624,I438105,I437627,I437639,I437636,I438194,I976079,I438220,I438237,I438186,I438259,I438276,I976094,I976082,I438293,I976073,I438319,I438327,I976085,I438353,I438361,I976076,I438378,I438165,I976091,I438418,I438426,I438159,I438174,I438471,I976100,I976088,I438488,I976097,I438514,I438162,I438536,I438553,I438570,I438177,I438601,I438618,I438168,I438649,I438171,I438183,I438180,I438738,I438764,I438781,I438730,I438803,I438820,I438837,I438863,I438871,I438897,I438905,I438922,I438709,I438962,I438970,I438703,I438718,I439015,I439032,I439058,I438706,I439080,I439097,I439114,I438721,I439145,I439162,I438712,I439193,I438715,I438727,I438724,I439282,I782234,I439308,I439325,I439274,I439347,I439364,I782228,I782225,I439381,I782240,I439407,I439415,I439441,I439449,I782222,I439466,I439253,I439506,I439514,I439247,I439262,I439559,I782237,I782231,I439576,I439602,I439250,I439624,I439641,I439658,I439265,I439689,I439706,I782243,I439256,I439737,I439259,I439271,I439268,I439826,I884993,I439852,I439869,I439818,I439891,I439908,I885008,I884996,I439925,I884987,I439951,I439959,I884999,I439985,I439993,I884990,I440010,I439797,I885005,I440050,I440058,I439791,I439806,I440103,I885014,I885002,I440120,I885011,I440146,I439794,I440168,I440185,I440202,I439809,I440233,I440250,I439800,I440281,I439803,I439815,I439812,I440370,I440396,I440413,I440362,I440435,I440452,I440469,I440495,I440503,I440529,I440537,I440554,I440341,I440594,I440602,I440335,I440350,I440647,I440664,I440690,I440338,I440712,I440729,I440746,I440353,I440777,I440794,I440344,I440825,I440347,I440359,I440356,I440914,I1177441,I440940,I440957,I440906,I440979,I440996,I1177453,I441013,I1177444,I441039,I441047,I1177462,I441073,I441081,I1177438,I441098,I440885,I1177456,I441138,I441146,I440879,I440894,I441191,I1177450,I1177447,I441208,I1177459,I441234,I440882,I441256,I441273,I441290,I440897,I441321,I441338,I440888,I441369,I440891,I440903,I440900,I441458,I755569,I441484,I441501,I441523,I441540,I755590,I755581,I441557,I441583,I441591,I755575,I441617,I441625,I755572,I441642,I755566,I441682,I441690,I441735,I755578,I441752,I755587,I441778,I441800,I441817,I441834,I441865,I441882,I755584,I441913,I442002,I1166459,I442028,I442045,I441994,I442067,I442084,I1166471,I442101,I1166462,I442127,I442135,I1166480,I442161,I442169,I1166456,I442186,I441973,I1166474,I442226,I442234,I441967,I441982,I442279,I1166468,I1166465,I442296,I1166477,I442322,I441970,I442344,I442361,I442378,I441985,I442409,I442426,I441976,I442457,I441979,I441991,I441988,I442546,I650951,I442572,I442589,I442538,I442611,I442628,I650972,I650963,I442645,I442671,I442679,I650957,I442705,I442713,I650954,I442730,I442517,I650948,I442770,I442778,I442511,I442526,I442823,I650960,I442840,I650969,I442866,I442514,I442888,I442905,I442922,I442529,I442953,I442970,I650966,I442520,I443001,I442523,I442535,I442532,I443090,I899851,I443116,I443133,I443082,I443155,I443172,I899866,I899854,I443189,I899845,I443215,I443223,I899857,I443249,I443257,I899848,I443274,I443061,I899863,I443314,I443322,I443055,I443070,I443367,I899872,I899860,I443384,I899869,I443410,I443058,I443432,I443449,I443466,I443073,I443497,I443514,I443064,I443545,I443067,I443079,I443076,I443634,I707017,I443660,I443677,I443699,I443716,I707038,I707029,I443733,I443759,I443767,I707023,I443793,I443801,I707020,I443818,I707014,I443858,I443866,I443911,I707026,I443928,I707035,I443954,I443976,I443993,I444010,I444041,I444058,I707032,I444089,I444178,I444204,I444221,I444243,I444260,I444277,I444303,I444311,I444337,I444345,I444362,I444402,I444410,I444455,I444472,I444498,I444520,I444537,I444554,I444585,I444602,I444633,I444722,I1242789,I444748,I444765,I444787,I444804,I1242801,I1242804,I444821,I1242807,I444847,I444855,I1242792,I444881,I444889,I1242798,I444906,I1242786,I444946,I444954,I444999,I1242810,I445016,I1242795,I445042,I445064,I445081,I445098,I445129,I445146,I445177,I445266,I851271,I445292,I445309,I445258,I445331,I445348,I851265,I851262,I445365,I851277,I445391,I445399,I445425,I445433,I851259,I445450,I445237,I445490,I445498,I445231,I445246,I445543,I851274,I851268,I445560,I445586,I445234,I445608,I445625,I445642,I445249,I445673,I445690,I851280,I445240,I445721,I445243,I445255,I445252,I445810,I734183,I445836,I445853,I445802,I445875,I445892,I734204,I734195,I445909,I445935,I445943,I734189,I445969,I445977,I734186,I445994,I445781,I734180,I446034,I446042,I445775,I445790,I446087,I734192,I446104,I734201,I446130,I445778,I446152,I446169,I446186,I445793,I446217,I446234,I734198,I445784,I446265,I445787,I445799,I445796,I446354,I446380,I446397,I446346,I446419,I446436,I446453,I446479,I446487,I446513,I446521,I446538,I446325,I446578,I446586,I446319,I446334,I446631,I446648,I446674,I446322,I446696,I446713,I446730,I446337,I446761,I446778,I446328,I446809,I446331,I446343,I446340,I446898,I564251,I446924,I446941,I446890,I446963,I446980,I564248,I564269,I446997,I564272,I447023,I447031,I564257,I447057,I447065,I564260,I447082,I446869,I564263,I447122,I447130,I446863,I446878,I447175,I564254,I447192,I564266,I447218,I446866,I447240,I447257,I447274,I446881,I447305,I447322,I446872,I447353,I446875,I446887,I446884,I447442,I810165,I447468,I447485,I447507,I447524,I810159,I810156,I447541,I810171,I447567,I447575,I447601,I447609,I810153,I447626,I447666,I447674,I447719,I810168,I810162,I447736,I447762,I447784,I447801,I447818,I447849,I447866,I810174,I447897,I447986,I921815,I448012,I448029,I447978,I448051,I448068,I921830,I921818,I448085,I921809,I448111,I448119,I921821,I448145,I448153,I921812,I448170,I447957,I921827,I448210,I448218,I447951,I447966,I448263,I921836,I921824,I448280,I921833,I448306,I447954,I448328,I448345,I448362,I447969,I448393,I448410,I447960,I448441,I447963,I447975,I447972,I448530,I525627,I448556,I448573,I448522,I448595,I448612,I525630,I525648,I448629,I525636,I448655,I448663,I448689,I448697,I525645,I448714,I448501,I525639,I448754,I448762,I448495,I448510,I448807,I525642,I525624,I448824,I525633,I448850,I448498,I448872,I448889,I448906,I448513,I448937,I448954,I448504,I448985,I448507,I448519,I448516,I449074,I449100,I449117,I449139,I449156,I449173,I449199,I449207,I449233,I449241,I449258,I449298,I449306,I449351,I449368,I449394,I449416,I449433,I449450,I449481,I449498,I449529,I449618,I946363,I449644,I449661,I449610,I449683,I449700,I946378,I946366,I449717,I946357,I449743,I449751,I946369,I449777,I449785,I946360,I449802,I449589,I946375,I449842,I449850,I449583,I449598,I449895,I946384,I946372,I449912,I946381,I449938,I449586,I449960,I449977,I449994,I449601,I450025,I450042,I449592,I450073,I449595,I449607,I449604,I450162,I720311,I450188,I450205,I450154,I450227,I450244,I720332,I720323,I450261,I450287,I450295,I720317,I450321,I450329,I720314,I450346,I450133,I720308,I450386,I450394,I450127,I450142,I450439,I720320,I450456,I720329,I450482,I450130,I450504,I450521,I450538,I450145,I450569,I450586,I720326,I450136,I450617,I450139,I450151,I450148,I450706,I744009,I450732,I450749,I450698,I450771,I450788,I744030,I744021,I450805,I450831,I450839,I744015,I450865,I450873,I744012,I450890,I450677,I744006,I450930,I450938,I450671,I450686,I450983,I744018,I451000,I744027,I451026,I450674,I451048,I451065,I451082,I450689,I451113,I451130,I744024,I450680,I451161,I450683,I450695,I450692,I451250,I922461,I451276,I451293,I451315,I451332,I922476,I922464,I451349,I922455,I451375,I451383,I922467,I451409,I451417,I922458,I451434,I922473,I451474,I451482,I451527,I922482,I922470,I451544,I922479,I451570,I451592,I451609,I451626,I451657,I451674,I451705,I451794,I1241157,I451820,I451837,I451859,I451876,I1241169,I1241172,I451893,I1241175,I451919,I451927,I1241160,I451953,I451961,I1241166,I451978,I1241154,I452018,I452026,I452071,I1241178,I452088,I1241163,I452114,I452136,I452153,I452170,I452201,I452218,I452249,I452338,I1116751,I452364,I452381,I452403,I452420,I1116763,I452437,I1116754,I452463,I452471,I1116772,I452497,I452505,I1116748,I452522,I1116766,I452562,I452570,I452615,I1116760,I1116757,I452632,I1116769,I452658,I452680,I452697,I452714,I452745,I452762,I452793,I452882,I452908,I452925,I452874,I452947,I452964,I452981,I453007,I453015,I453041,I453049,I453066,I452853,I453106,I453114,I452847,I452862,I453159,I453176,I453202,I452850,I453224,I453241,I453258,I452865,I453289,I453306,I452856,I453337,I452859,I452871,I452868,I453426,I1228645,I453452,I453469,I453491,I453508,I1228657,I1228660,I453525,I1228663,I453551,I453559,I1228648,I453585,I453593,I1228654,I453610,I1228642,I453650,I453658,I453703,I1228666,I453720,I1228651,I453746,I453768,I453785,I453802,I453833,I453850,I453881,I453970,I722045,I453996,I454013,I453962,I454035,I454052,I722066,I722057,I454069,I454095,I454103,I722051,I454129,I454137,I722048,I454154,I453941,I722042,I454194,I454202,I453935,I453950,I454247,I722054,I454264,I722063,I454290,I453938,I454312,I454329,I454346,I453953,I454377,I454394,I722060,I453944,I454425,I453947,I453959,I453956,I454514,I454540,I454557,I454506,I454579,I454596,I454613,I454639,I454647,I454673,I454681,I454698,I454485,I454738,I454746,I454479,I454494,I454791,I454808,I454834,I454482,I454856,I454873,I454890,I454497,I454921,I454938,I454488,I454969,I454491,I454503,I454500,I455058,I1274424,I455084,I455101,I455050,I455123,I455140,I1274421,I1274418,I455157,I1274406,I455183,I455191,I1274430,I455217,I455225,I1274415,I455242,I455029,I1274409,I455282,I455290,I455023,I455038,I455335,I1274412,I455352,I1274427,I455378,I455026,I455400,I455417,I455434,I455041,I455465,I455482,I455032,I455513,I455035,I455047,I455044,I455602,I570031,I455628,I455645,I455594,I455667,I455684,I570028,I570049,I455701,I570052,I455727,I455735,I570037,I455761,I455769,I570040,I455786,I455573,I570043,I455826,I455834,I455567,I455582,I455879,I570034,I455896,I570046,I455922,I455570,I455944,I455961,I455978,I455585,I456009,I456026,I455576,I456057,I455579,I455591,I455588,I456146,I764817,I456172,I456189,I456211,I456228,I764838,I764829,I456245,I456271,I456279,I764823,I456305,I456313,I764820,I456330,I764814,I456370,I456378,I456423,I764826,I456440,I764835,I456466,I456488,I456505,I456522,I456553,I456570,I764832,I456601,I456690,I752101,I456716,I456733,I456682,I456755,I456772,I752122,I752113,I456789,I456815,I456823,I752107,I456849,I456857,I752104,I456874,I456661,I752098,I456914,I456922,I456655,I456670,I456967,I752110,I456984,I752119,I457010,I456658,I457032,I457049,I457066,I456673,I457097,I457114,I752116,I456664,I457145,I456667,I456679,I456676,I457234,I691411,I457260,I457277,I457226,I457299,I457316,I691432,I691423,I457333,I457359,I457367,I691417,I457393,I457401,I691414,I457418,I457205,I691408,I457458,I457466,I457199,I457214,I457511,I691420,I457528,I691429,I457554,I457202,I457576,I457593,I457610,I457217,I457641,I457658,I691426,I457208,I457689,I457211,I457223,I457220,I457778,I1089585,I457804,I457821,I457843,I457860,I1089597,I457877,I1089588,I457903,I457911,I1089606,I457937,I457945,I1089582,I457962,I1089600,I458002,I458010,I458055,I1089594,I1089591,I458072,I1089603,I458098,I458120,I458137,I458154,I458185,I458202,I458233,I458322,I590839,I458348,I458365,I458387,I458404,I590836,I590857,I458421,I590860,I458447,I458455,I590845,I458481,I458489,I590848,I458506,I590851,I458546,I458554,I458599,I590842,I458616,I590854,I458642,I458664,I458681,I458698,I458729,I458746,I458777,I458866,I1171083,I458892,I458909,I458858,I458931,I458948,I1171095,I458965,I1171086,I458991,I458999,I1171104,I459025,I459033,I1171080,I459050,I458837,I1171098,I459090,I459098,I458831,I458846,I459143,I1171092,I1171089,I459160,I1171101,I459186,I458834,I459208,I459225,I459242,I458849,I459273,I459290,I458840,I459321,I458843,I458855,I458852,I459410,I1061263,I459436,I459453,I459402,I459475,I459492,I1061275,I459509,I1061266,I459535,I459543,I1061284,I459569,I459577,I1061260,I459594,I459381,I1061278,I459634,I459642,I459375,I459390,I459687,I1061272,I1061269,I459704,I1061281,I459730,I459378,I459752,I459769,I459786,I459393,I459817,I459834,I459384,I459865,I459387,I459399,I459396,I459954,I504207,I459980,I459997,I459946,I460019,I460036,I504210,I504228,I460053,I504216,I460079,I460087,I460113,I460121,I504225,I460138,I459925,I504219,I460178,I460186,I459919,I459934,I460231,I504222,I504204,I460248,I504213,I460274,I459922,I460296,I460313,I460330,I459937,I460361,I460378,I459928,I460409,I459931,I459943,I459940,I460498,I1003211,I460524,I460541,I460563,I460580,I1003226,I1003214,I460597,I1003205,I460623,I460631,I1003217,I460657,I460665,I1003208,I460682,I1003223,I460722,I460730,I460775,I1003232,I1003220,I460792,I1003229,I460818,I460840,I460857,I460874,I460905,I460922,I460953,I461042,I461068,I461085,I461034,I461107,I461124,I461141,I461167,I461175,I461201,I461209,I461226,I461013,I461266,I461274,I461007,I461022,I461319,I461336,I461362,I461010,I461384,I461401,I461418,I461025,I461449,I461466,I461016,I461497,I461019,I461031,I461028,I461586,I1168193,I461612,I461629,I461651,I461668,I1168205,I461685,I1168196,I461711,I461719,I1168214,I461745,I461753,I1168190,I461770,I1168208,I461810,I461818,I461863,I1168202,I1168199,I461880,I1168211,I461906,I461928,I461945,I461962,I461993,I462010,I462041,I462130,I816489,I462156,I462173,I462195,I462212,I816483,I816480,I462229,I816495,I462255,I462263,I462289,I462297,I816477,I462314,I462354,I462362,I462407,I816492,I816486,I462424,I462450,I462472,I462489,I462506,I462537,I462554,I816498,I462585,I462674,I523842,I462700,I462717,I462666,I462739,I462756,I523845,I523863,I462773,I523851,I462799,I462807,I462833,I462841,I523860,I462858,I462645,I523854,I462898,I462906,I462639,I462654,I462951,I523857,I523839,I462968,I523848,I462994,I462642,I463016,I463033,I463050,I462657,I463081,I463098,I462648,I463129,I462651,I462663,I462660,I463218,I963805,I463244,I463261,I463210,I463283,I463300,I963820,I963808,I463317,I963799,I463343,I463351,I963811,I463377,I463385,I963802,I463402,I463189,I963817,I463442,I463450,I463183,I463198,I463495,I963826,I963814,I463512,I963823,I463538,I463186,I463560,I463577,I463594,I463201,I463625,I463642,I463192,I463673,I463195,I463207,I463204,I463762,I463788,I463805,I463754,I463827,I463844,I463861,I463887,I463895,I463921,I463929,I463946,I463733,I463986,I463994,I463727,I463742,I464039,I464056,I464082,I463730,I464104,I464121,I464138,I463745,I464169,I464186,I463736,I464217,I463739,I463751,I463748,I464306,I464332,I464349,I464371,I464388,I464405,I464431,I464439,I464465,I464473,I464490,I464530,I464538,I464583,I464600,I464626,I464648,I464665,I464682,I464713,I464730,I464761,I464850,I769441,I464876,I464893,I464842,I464915,I464932,I769462,I769453,I464949,I464975,I464983,I769447,I465009,I465017,I769444,I465034,I464821,I769438,I465074,I465082,I464815,I464830,I465127,I769450,I465144,I769459,I465170,I464818,I465192,I465209,I465226,I464833,I465257,I465274,I769456,I464824,I465305,I464827,I464839,I464836,I465394,I959283,I465420,I465437,I465386,I465459,I465476,I959298,I959286,I465493,I959277,I465519,I465527,I959289,I465553,I465561,I959280,I465578,I465365,I959295,I465618,I465626,I465359,I465374,I465671,I959304,I959292,I465688,I959301,I465714,I465362,I465736,I465753,I465770,I465377,I465801,I465818,I465368,I465849,I465371,I465383,I465380,I465938,I877621,I465964,I465981,I465930,I466003,I466020,I877615,I877612,I466037,I877627,I466063,I466071,I466097,I466105,I877609,I466122,I465909,I466162,I466170,I465903,I465918,I466215,I877624,I877618,I466232,I466258,I465906,I466280,I466297,I466314,I465921,I466345,I466362,I877630,I465912,I466393,I465915,I465927,I465924,I466482,I466508,I466525,I466474,I466547,I466564,I466581,I466607,I466615,I466641,I466649,I466666,I466453,I466706,I466714,I466447,I466462,I466759,I466776,I466802,I466450,I466824,I466841,I466858,I466465,I466889,I466906,I466456,I466937,I466459,I466471,I466468,I467026,I934089,I467052,I467069,I467091,I467108,I934104,I934092,I467125,I934083,I467151,I467159,I934095,I467185,I467193,I934086,I467210,I934101,I467250,I467258,I467303,I934110,I934098,I467320,I934107,I467346,I467368,I467385,I467402,I467433,I467450,I467481,I467570,I602977,I467596,I467613,I467562,I467635,I467652,I602974,I602995,I467669,I602998,I467695,I467703,I602983,I467729,I467737,I602986,I467754,I467541,I602989,I467794,I467802,I467535,I467550,I467847,I602980,I467864,I602992,I467890,I467538,I467912,I467929,I467946,I467553,I467977,I467994,I467544,I468025,I467547,I467559,I467556,I468114,I1008379,I468140,I468157,I468179,I468196,I1008394,I1008382,I468213,I1008373,I468239,I468247,I1008385,I468273,I468281,I1008376,I468298,I1008391,I468338,I468346,I468391,I1008400,I1008388,I468408,I1008397,I468434,I468456,I468473,I468490,I468521,I468538,I468569,I468658,I967681,I468684,I468701,I468650,I468723,I468740,I967696,I967684,I468757,I967675,I468783,I468791,I967687,I468817,I468825,I967678,I468842,I468629,I967693,I468882,I468890,I468623,I468638,I468935,I967702,I967690,I468952,I967699,I468978,I468626,I469000,I469017,I469034,I468641,I469065,I469082,I468632,I469113,I468635,I468647,I468644,I469202,I469228,I469245,I469194,I469267,I469284,I469301,I469327,I469335,I469361,I469369,I469386,I469173,I469426,I469434,I469167,I469182,I469479,I469496,I469522,I469170,I469544,I469561,I469578,I469185,I469609,I469626,I469176,I469657,I469179,I469191,I469188,I469746,I469772,I469789,I469738,I469811,I469828,I469845,I469871,I469879,I469905,I469913,I469930,I469717,I469970,I469978,I469711,I469726,I470023,I470040,I470066,I469714,I470088,I470105,I470122,I469729,I470153,I470170,I469720,I470201,I469723,I469735,I469732,I470290,I470316,I470333,I470355,I470372,I470389,I470415,I470423,I470449,I470457,I470474,I470514,I470522,I470567,I470584,I470610,I470632,I470649,I470666,I470697,I470714,I470745,I470834,I470860,I470877,I470899,I470916,I470933,I470959,I470967,I470993,I471001,I471018,I471058,I471066,I471111,I471128,I471154,I471176,I471193,I471210,I471241,I471258,I471289,I471378,I687365,I471404,I471421,I471370,I471443,I471460,I687386,I687377,I471477,I471503,I471511,I687371,I471537,I471545,I687368,I471562,I471349,I687362,I471602,I471610,I471343,I471358,I471655,I687374,I471672,I687383,I471698,I471346,I471720,I471737,I471754,I471361,I471785,I471802,I687380,I471352,I471833,I471355,I471367,I471364,I471922,I471948,I471965,I471914,I471987,I472004,I472021,I472047,I472055,I472081,I472089,I472106,I471893,I472146,I472154,I471887,I471902,I472199,I472216,I472242,I471890,I472264,I472281,I472298,I471905,I472329,I472346,I471896,I472377,I471899,I471911,I471908,I472466,I1283094,I472492,I472509,I472458,I472531,I472548,I1283091,I1283088,I472565,I1283076,I472591,I472599,I1283100,I472625,I472633,I1283085,I472650,I472437,I1283079,I472690,I472698,I472431,I472446,I472743,I1283082,I472760,I1283097,I472786,I472434,I472808,I472825,I472842,I472449,I472873,I472890,I472440,I472921,I472443,I472455,I472452,I473010,I996105,I473036,I473053,I473002,I473075,I473092,I996120,I996108,I473109,I996099,I473135,I473143,I996111,I473169,I473177,I996102,I473194,I472981,I996117,I473234,I473242,I472975,I472990,I473287,I996126,I996114,I473304,I996123,I473330,I472978,I473352,I473369,I473386,I472993,I473417,I473434,I472984,I473465,I472987,I472999,I472996,I473554,I934735,I473580,I473597,I473619,I473636,I934750,I934738,I473653,I934729,I473679,I473687,I934741,I473713,I473721,I934732,I473738,I934747,I473778,I473786,I473831,I934756,I934744,I473848,I934753,I473874,I473896,I473913,I473930,I473961,I473978,I474009,I474098,I474124,I474141,I474090,I474163,I474180,I474197,I474223,I474231,I474257,I474265,I474282,I474069,I474322,I474330,I474063,I474078,I474375,I474392,I474418,I474066,I474440,I474457,I474474,I474081,I474505,I474522,I474072,I474553,I474075,I474087,I474084,I474642,I1096521,I474668,I474685,I474707,I474724,I1096533,I474741,I1096524,I474767,I474775,I1096542,I474801,I474809,I1096518,I474826,I1096536,I474866,I474874,I474919,I1096530,I1096527,I474936,I1096539,I474962,I474984,I475001,I475018,I475049,I475066,I475097,I475186,I1230821,I475212,I475229,I475178,I475251,I475268,I1230833,I1230836,I475285,I1230839,I475311,I475319,I1230824,I475345,I475353,I1230830,I475370,I475157,I1230818,I475410,I475418,I475151,I475166,I475463,I1230842,I475480,I1230827,I475506,I475154,I475528,I475545,I475562,I475169,I475593,I475610,I475160,I475641,I475163,I475175,I475172,I475730,I475756,I475773,I475722,I475795,I475812,I475829,I475855,I475863,I475889,I475897,I475914,I475701,I475954,I475962,I475695,I475710,I476007,I476024,I476050,I475698,I476072,I476089,I476106,I475713,I476137,I476154,I475704,I476185,I475707,I475719,I475716,I476274,I1287718,I476300,I476317,I476339,I476356,I1287715,I1287712,I476373,I1287700,I476399,I476407,I1287724,I476433,I476441,I1287709,I476458,I1287703,I476498,I476506,I476551,I1287706,I476568,I1287721,I476594,I476616,I476633,I476650,I476681,I476698,I476729,I476818,I476844,I476861,I476810,I476883,I476900,I476917,I476943,I476951,I476977,I476985,I477002,I476789,I477042,I477050,I476783,I476798,I477095,I477112,I477138,I476786,I477160,I477177,I477194,I476801,I477225,I477242,I476792,I477273,I476795,I476807,I476804,I477362,I477388,I477405,I477354,I477427,I477444,I477461,I477487,I477495,I477521,I477529,I477546,I477333,I477586,I477594,I477327,I477342,I477639,I477656,I477682,I477330,I477704,I477721,I477738,I477345,I477769,I477786,I477336,I477817,I477339,I477351,I477348,I477906,I829664,I477932,I477949,I477898,I477971,I477988,I829658,I829655,I478005,I829670,I478031,I478039,I478065,I478073,I829652,I478090,I477877,I478130,I478138,I477871,I477886,I478183,I829667,I829661,I478200,I478226,I477874,I478248,I478265,I478282,I477889,I478313,I478330,I829673,I477880,I478361,I477883,I477895,I477892,I478450,I1106925,I478476,I478493,I478442,I478515,I478532,I1106937,I478549,I1106928,I478575,I478583,I1106946,I478609,I478617,I1106922,I478634,I478421,I1106940,I478674,I478682,I478415,I478430,I478727,I1106934,I1106931,I478744,I1106943,I478770,I478418,I478792,I478809,I478826,I478433,I478857,I478874,I478424,I478905,I478427,I478439,I478436,I478994,I1120219,I479020,I479037,I478986,I479059,I479076,I1120231,I479093,I1120222,I479119,I479127,I1120240,I479153,I479161,I1120216,I479178,I478965,I1120234,I479218,I479226,I478959,I478974,I479271,I1120228,I1120225,I479288,I1120237,I479314,I478962,I479336,I479353,I479370,I478977,I479401,I479418,I478968,I479449,I478971,I478983,I478980,I479538,I479564,I479581,I479603,I479620,I479637,I479663,I479671,I479697,I479705,I479722,I479762,I479770,I479815,I479832,I479858,I479880,I479897,I479914,I479945,I479962,I479993,I480082,I542287,I480108,I480125,I480147,I480164,I542284,I542305,I480181,I542308,I480207,I480215,I542293,I480241,I480249,I542296,I480266,I542299,I480306,I480314,I480359,I542290,I480376,I542302,I480402,I480424,I480441,I480458,I480489,I480506,I480537,I480626,I916647,I480652,I480669,I480691,I480708,I916662,I916650,I480725,I916641,I480751,I480759,I916653,I480785,I480793,I916644,I480810,I916659,I480850,I480858,I480903,I916668,I916656,I480920,I916665,I480946,I480968,I480985,I481002,I481033,I481050,I481081,I481170,I963159,I481196,I481213,I481162,I481235,I481252,I963174,I963162,I481269,I963153,I481295,I481303,I963165,I481329,I481337,I963156,I481354,I481141,I963171,I481394,I481402,I481135,I481150,I481447,I963180,I963168,I481464,I963177,I481490,I481138,I481512,I481529,I481546,I481153,I481577,I481594,I481144,I481625,I481147,I481159,I481156,I481714,I1260552,I481740,I481757,I481706,I481779,I481796,I1260549,I1260546,I481813,I1260534,I481839,I481847,I1260558,I481873,I481881,I1260543,I481898,I481685,I1260537,I481938,I481946,I481679,I481694,I481991,I1260540,I482008,I1260555,I482034,I481682,I482056,I482073,I482090,I481697,I482121,I482138,I481688,I482169,I481691,I481703,I481700,I482258,I482284,I482301,I482323,I482340,I482357,I482383,I482391,I482417,I482425,I482442,I482482,I482490,I482535,I482552,I482578,I482600,I482617,I482634,I482665,I482682,I482713,I482802,I945717,I482828,I482845,I482794,I482867,I482884,I945732,I945720,I482901,I945711,I482927,I482935,I945723,I482961,I482969,I945714,I482986,I482773,I945729,I483026,I483034,I482767,I482782,I483079,I945738,I945726,I483096,I945735,I483122,I482770,I483144,I483161,I483178,I482785,I483209,I483226,I482776,I483257,I482779,I482791,I482788,I483346,I1005795,I483372,I483389,I483411,I483428,I1005810,I1005798,I483445,I1005789,I483471,I483479,I1005801,I483505,I483513,I1005792,I483530,I1005807,I483570,I483578,I483623,I1005816,I1005804,I483640,I1005813,I483666,I483688,I483705,I483722,I483753,I483770,I483801,I483890,I1343419,I483916,I483933,I483882,I483955,I483972,I1343395,I1343416,I483989,I1343413,I484015,I484023,I1343392,I484049,I484057,I1343404,I484074,I483861,I1343407,I484114,I484122,I483855,I483870,I484167,I1343410,I1343398,I484184,I1343401,I484210,I483858,I484232,I484249,I484266,I483873,I484297,I484314,I483864,I484345,I483867,I483879,I483876,I484434,I1083227,I484460,I484477,I484426,I484499,I484516,I1083239,I484533,I1083230,I484559,I484567,I1083248,I484593,I484601,I1083224,I484618,I484405,I1083242,I484658,I484666,I484399,I484414,I484711,I1083236,I1083233,I484728,I1083245,I484754,I484402,I484776,I484793,I484810,I484417,I484841,I484858,I484408,I484889,I484411,I484423,I484420,I484978,I870770,I485004,I485021,I485043,I485060,I870764,I870761,I485077,I870776,I485103,I485111,I485137,I485145,I870758,I485162,I485202,I485210,I485255,I870773,I870767,I485272,I485298,I485320,I485337,I485354,I485385,I485402,I870779,I485433,I485522,I1021922,I485548,I485565,I485514,I485587,I485604,I1021940,I485621,I1021934,I485647,I485655,I1021928,I485681,I485689,I1021937,I485706,I485493,I1021925,I485746,I485754,I485487,I485502,I485799,I1021943,I485816,I485842,I485490,I485864,I485881,I485898,I485505,I485929,I485946,I1021931,I485496,I485977,I485499,I485511,I485508,I486066,I676961,I486092,I486109,I486058,I486131,I486148,I676982,I676973,I486165,I486191,I486199,I676967,I486225,I486233,I676964,I486250,I486037,I676958,I486290,I486298,I486031,I486046,I486343,I676970,I486360,I676979,I486386,I486034,I486408,I486425,I486442,I486049,I486473,I486490,I676976,I486040,I486521,I486043,I486055,I486052,I486610,I943779,I486636,I486653,I486602,I486675,I486692,I943794,I943782,I486709,I943773,I486735,I486743,I943785,I486769,I486777,I943776,I486794,I486581,I943791,I486834,I486842,I486575,I486590,I486887,I943800,I943788,I486904,I943797,I486930,I486578,I486952,I486969,I486986,I486593,I487017,I487034,I486584,I487065,I486587,I486599,I486596,I487154,I487180,I487197,I487146,I487219,I487236,I487253,I487279,I487287,I487313,I487321,I487338,I487125,I487378,I487386,I487119,I487134,I487431,I487448,I487474,I487122,I487496,I487513,I487530,I487137,I487561,I487578,I487128,I487609,I487131,I487143,I487140,I487698,I965097,I487724,I487741,I487763,I487780,I965112,I965100,I487797,I965091,I487823,I487831,I965103,I487857,I487865,I965094,I487882,I965109,I487922,I487930,I487975,I965118,I965106,I487992,I965115,I488018,I488040,I488057,I488074,I488105,I488122,I488153,I488242,I1001919,I488268,I488285,I488307,I488324,I1001934,I1001922,I488341,I1001913,I488367,I488375,I1001925,I488401,I488409,I1001916,I488426,I1001931,I488466,I488474,I488519,I1001940,I1001928,I488536,I1001937,I488562,I488584,I488601,I488618,I488649,I488666,I488697,I488786,I536932,I488812,I488829,I488778,I488851,I488868,I536935,I536953,I488885,I536941,I488911,I488919,I488945,I488953,I536950,I488970,I488757,I536944,I489010,I489018,I488751,I488766,I489063,I536947,I536929,I489080,I536938,I489106,I488754,I489128,I489145,I489162,I488769,I489193,I489210,I488760,I489241,I488763,I488775,I488772,I489330,I652685,I489356,I489373,I489322,I489395,I489412,I652706,I652697,I489429,I489455,I489463,I652691,I489489,I489497,I652688,I489514,I489301,I652682,I489554,I489562,I489295,I489310,I489607,I652694,I489624,I652703,I489650,I489298,I489672,I489689,I489706,I489313,I489737,I489754,I652700,I489304,I489785,I489307,I489319,I489316,I489874,I489900,I489917,I489939,I489956,I489973,I489999,I490007,I490033,I490041,I490058,I490098,I490106,I490151,I490168,I490194,I490216,I490233,I490250,I490281,I490298,I490329,I490418,I490444,I490461,I490410,I490483,I490500,I490517,I490543,I490551,I490577,I490585,I490602,I490389,I490642,I490650,I490383,I490398,I490695,I490712,I490738,I490386,I490760,I490777,I490794,I490401,I490825,I490842,I490392,I490873,I490395,I490407,I490404,I490962,I1138137,I490988,I491005,I491027,I491044,I1138149,I491061,I1138140,I491087,I491095,I1138158,I491121,I491129,I1138134,I491146,I1138152,I491186,I491194,I491239,I1138146,I1138143,I491256,I1138155,I491282,I491304,I491321,I491338,I491369,I491386,I491417,I491506,I783288,I491532,I491549,I491498,I491571,I491588,I783282,I783279,I491605,I783294,I491631,I491639,I491665,I491673,I783276,I491690,I491477,I491730,I491738,I491471,I491486,I491783,I783291,I783285,I491800,I491826,I491474,I491848,I491865,I491882,I491489,I491913,I491930,I783297,I491480,I491961,I491483,I491495,I491492,I492050,I648061,I492076,I492093,I492042,I492115,I492132,I648082,I648073,I492149,I492175,I492183,I648067,I492209,I492217,I648064,I492234,I492021,I648058,I492274,I492282,I492015,I492030,I492327,I648070,I492344,I648079,I492370,I492018,I492392,I492409,I492426,I492033,I492457,I492474,I648076,I492024,I492505,I492027,I492039,I492036,I492594,I1348179,I492620,I492637,I492586,I492659,I492676,I1348155,I1348176,I492693,I1348173,I492719,I492727,I1348152,I492753,I492761,I1348164,I492778,I492565,I1348167,I492818,I492826,I492559,I492574,I492871,I1348170,I1348158,I492888,I1348161,I492914,I492562,I492936,I492953,I492970,I492577,I493001,I493018,I492568,I493049,I492571,I492583,I492580,I493138,I1229733,I493164,I493181,I493203,I493220,I1229745,I1229748,I493237,I1229751,I493263,I493271,I1229736,I493297,I493305,I1229742,I493322,I1229730,I493362,I493370,I493415,I1229754,I493432,I1229739,I493458,I493480,I493497,I493514,I493545,I493562,I493593,I493682,I1373169,I493708,I493725,I493747,I493764,I1373145,I1373166,I493781,I1373163,I493807,I493815,I1373142,I493841,I493849,I1373154,I493866,I1373157,I493906,I493914,I493959,I1373160,I1373148,I493976,I1373151,I494002,I494024,I494041,I494058,I494089,I494106,I494137,I494226,I1344609,I494252,I494269,I494291,I494308,I1344585,I1344606,I494325,I1344603,I494351,I494359,I1344582,I494385,I494393,I1344594,I494410,I1344597,I494450,I494458,I494503,I1344600,I1344588,I494520,I1344591,I494546,I494568,I494585,I494602,I494633,I494650,I494681,I494770,I494796,I494813,I494835,I494852,I494869,I494895,I494903,I494929,I494937,I494954,I494994,I495002,I495047,I495064,I495090,I495112,I495129,I495146,I495177,I495194,I495225,I495311,I932160,I495337,I495354,I495303,I932148,I495385,I495393,I932145,I495410,I495427,I932157,I495444,I932154,I495461,I495478,I495495,I495300,I495526,I932163,I495543,I932166,I495560,I495285,I495297,I495605,I495622,I495291,I495653,I932169,I495670,I495279,I495701,I932172,I495718,I932151,I495735,I495761,I495769,I495288,I495800,I495817,I495294,I495848,I495282,I495906,I1097692,I495932,I495949,I1097674,I495980,I495988,I1097680,I496005,I496022,I1097695,I496039,I1097686,I496056,I496073,I496090,I496121,I1097698,I496138,I1097677,I496155,I496200,I496217,I496248,I1097683,I496265,I496296,I1097689,I496313,I496330,I496356,I496364,I496395,I496412,I496443,I496501,I864970,I496527,I496544,I496493,I864967,I496575,I496583,I496600,I496617,I864964,I496634,I864979,I496651,I496668,I496685,I496490,I496716,I864973,I496733,I864961,I496750,I496475,I496487,I496795,I496812,I496481,I496843,I864982,I496860,I496469,I496891,I496908,I864976,I496925,I496951,I496959,I496478,I496990,I497007,I496484,I497038,I496472,I497096,I1067636,I497122,I497139,I497088,I1067618,I497170,I497178,I1067624,I497195,I497212,I1067639,I497229,I1067630,I497246,I497263,I497280,I497085,I497311,I1067642,I497328,I1067621,I497345,I497070,I497082,I497390,I497407,I497076,I497438,I1067627,I497455,I497064,I497486,I1067633,I497503,I497520,I497546,I497554,I497073,I497585,I497602,I497079,I497633,I497067,I497691,I792771,I497717,I497734,I497683,I792768,I497765,I497773,I497790,I497807,I792765,I497824,I792780,I497841,I497858,I497875,I497680,I497906,I792774,I497923,I792762,I497940,I497665,I497677,I497985,I498002,I497671,I498033,I792783,I498050,I497659,I498081,I498098,I792777,I498115,I498141,I498149,I497668,I498180,I498197,I497674,I498228,I497662,I498286,I956708,I498312,I498329,I956696,I498360,I498368,I956693,I498385,I498402,I956705,I498419,I956702,I498436,I498453,I498470,I498501,I956711,I498518,I956714,I498535,I498580,I498597,I498628,I956717,I498645,I498676,I956720,I498693,I956699,I498710,I498736,I498744,I498775,I498792,I498823,I498881,I1113298,I498907,I498924,I498873,I1113280,I498955,I498963,I1113286,I498980,I498997,I1113301,I499014,I1113292,I499031,I499048,I499065,I498870,I499096,I1113304,I499113,I1113283,I499130,I498855,I498867,I499175,I499192,I498861,I499223,I1113289,I499240,I498849,I499271,I1113295,I499288,I499305,I499331,I499339,I498858,I499370,I499387,I498864,I499418,I498852,I499476,I998052,I499502,I499519,I998040,I499550,I499558,I998037,I499575,I499592,I998049,I499609,I998046,I499626,I499643,I499660,I499691,I998055,I499708,I998058,I499725,I499770,I499787,I499818,I998061,I499835,I499866,I998064,I499883,I998043,I499900,I499926,I499934,I499965,I499982,I500013,I500071,I500097,I500114,I500063,I500145,I500153,I500170,I500187,I500204,I500221,I500238,I500255,I500060,I500286,I500303,I500320,I500045,I500057,I500365,I500382,I500051,I500413,I500430,I500039,I500461,I500478,I500495,I500521,I500529,I500048,I500560,I500577,I500054,I500608,I500042,I500666,I500692,I500709,I500658,I500740,I500748,I500765,I500782,I500799,I500816,I500833,I500850,I500655,I500881,I500898,I500915,I500640,I500652,I500960,I500977,I500646,I501008,I501025,I500634,I501056,I501073,I501090,I501116,I501124,I500643,I501155,I501172,I500649,I501203,I500637,I501261,I563673,I501287,I501304,I501253,I563685,I501335,I501343,I563670,I501360,I501377,I563688,I501394,I563679,I501411,I501428,I501445,I501250,I501476,I563691,I501493,I563694,I501510,I501235,I501247,I501555,I501572,I501241,I501603,I501620,I501229,I501651,I563682,I501668,I563676,I501685,I501711,I501719,I501238,I501750,I501767,I501244,I501798,I501232,I501856,I1225922,I501882,I501899,I501848,I1225937,I501930,I501938,I1225946,I501955,I501972,I1225925,I501989,I1225931,I502006,I502023,I502040,I501845,I502071,I1225943,I502088,I1225940,I502105,I501830,I501842,I502150,I502167,I501836,I502198,I502215,I501824,I502246,I1225934,I502263,I1225928,I502280,I502306,I502314,I501833,I502345,I502362,I501839,I502393,I501827,I502451,I656737,I502477,I502494,I502443,I656731,I502525,I502533,I656728,I502550,I502567,I656740,I502584,I656743,I502601,I502618,I502635,I502440,I502666,I656752,I502683,I656746,I502700,I502425,I502437,I502745,I502762,I502431,I502793,I656734,I502810,I502419,I502841,I656749,I502858,I502875,I502901,I502909,I502428,I502940,I502957,I502434,I502988,I502422,I503046,I503072,I503089,I503120,I503128,I503145,I503162,I503179,I503196,I503213,I503230,I503261,I503278,I503295,I503340,I503357,I503388,I503405,I503436,I503453,I503470,I503496,I503504,I503535,I503552,I503583,I503641,I503667,I503684,I503715,I503723,I503740,I503757,I503774,I503791,I503808,I503825,I503856,I503873,I503890,I503935,I503952,I503983,I504000,I504031,I504048,I504065,I504091,I504099,I504130,I504147,I504178,I504236,I820175,I504262,I504279,I820172,I504310,I504318,I504335,I504352,I820169,I504369,I820184,I504386,I504403,I504420,I504451,I820178,I504468,I820166,I504485,I504530,I504547,I504578,I820187,I504595,I504626,I504643,I820181,I504660,I504686,I504694,I504725,I504742,I504773,I504831,I1310072,I504857,I504874,I504823,I1310078,I504905,I504913,I1310093,I504930,I504947,I1310084,I504964,I1310081,I504981,I504998,I505015,I504820,I505046,I505063,I1310096,I505080,I504805,I504817,I505125,I505142,I504811,I505173,I1310090,I505190,I504799,I505221,I1310075,I505238,I1310087,I505255,I1310099,I505281,I505289,I504808,I505320,I505337,I504814,I505368,I504802,I505426,I505452,I505469,I505418,I505500,I505508,I505525,I505542,I505559,I505576,I505593,I505610,I505415,I505641,I505658,I505675,I505400,I505412,I505720,I505737,I505406,I505768,I505785,I505394,I505816,I505833,I505850,I505876,I505884,I505403,I505915,I505932,I505409,I505963,I505397,I506021,I899214,I506047,I506064,I506013,I899202,I506095,I506103,I899199,I506120,I506137,I899211,I506154,I899208,I506171,I506188,I506205,I506010,I506236,I899217,I506253,I899220,I506270,I505995,I506007,I506315,I506332,I506001,I506363,I899223,I506380,I505989,I506411,I899226,I506428,I899205,I506445,I506471,I506479,I505998,I506510,I506527,I506004,I506558,I505992,I506616,I506642,I506659,I506608,I506690,I506698,I506715,I506732,I506749,I506766,I506783,I506800,I506605,I506831,I506848,I506865,I506590,I506602,I506910,I506927,I506596,I506958,I506975,I506584,I507006,I507023,I507040,I507066,I507074,I506593,I507105,I507122,I506599,I507153,I506587,I507211,I1025288,I507237,I507254,I507203,I1025291,I507285,I507293,I1025294,I507310,I507327,I1025306,I507344,I1025297,I507361,I507378,I507395,I507200,I507426,I1025303,I507443,I507460,I507185,I507197,I507505,I507522,I507191,I507553,I507570,I507179,I507601,I1025300,I507618,I507635,I1025309,I507661,I507669,I507188,I507700,I507717,I507194,I507748,I507182,I507806,I1257075,I507832,I507849,I507798,I1257081,I507880,I507888,I1257069,I507905,I507922,I1257072,I507939,I1257078,I507956,I507973,I507990,I507795,I508021,I508038,I1257087,I508055,I507780,I507792,I508100,I508117,I507786,I508148,I1257066,I508165,I507774,I508196,I1257090,I508213,I508230,I1257084,I508256,I508264,I507783,I508295,I508312,I507789,I508343,I507777,I508401,I586793,I508427,I508444,I586805,I508475,I508483,I586790,I508500,I508517,I586808,I508534,I586799,I508551,I508568,I508585,I508616,I586811,I508633,I586814,I508650,I508695,I508712,I508743,I508760,I508791,I586802,I508808,I586796,I508825,I508851,I508859,I508890,I508907,I508938,I508996,I1178034,I509022,I509039,I1178016,I509070,I509078,I1178022,I509095,I509112,I1178037,I509129,I1178028,I509146,I509163,I509180,I509211,I1178040,I509228,I1178019,I509245,I509290,I509307,I509338,I1178025,I509355,I509386,I1178031,I509403,I509420,I509446,I509454,I509485,I509502,I509533,I509591,I509617,I509634,I509665,I509673,I509690,I509707,I509724,I509741,I509758,I509775,I509806,I509823,I509840,I509885,I509902,I509933,I509950,I509981,I509998,I510015,I510041,I510049,I510080,I510097,I510128,I510186,I510212,I510229,I510260,I510268,I510285,I510302,I510319,I510336,I510353,I510370,I510401,I510418,I510435,I510480,I510497,I510528,I510545,I510576,I510593,I510610,I510636,I510644,I510675,I510692,I510723,I510781,I510807,I510824,I510773,I510855,I510863,I510880,I510897,I510914,I510931,I510948,I510965,I510770,I510996,I511013,I511030,I510755,I510767,I511075,I511092,I510761,I511123,I511140,I510749,I511171,I511188,I511205,I511231,I511239,I510758,I511270,I511287,I510764,I511318,I510752,I511376,I511402,I511419,I511368,I511450,I511458,I511475,I511492,I511509,I511526,I511543,I511560,I511365,I511591,I511608,I511625,I511350,I511362,I511670,I511687,I511356,I511718,I511735,I511344,I511766,I511783,I511800,I511826,I511834,I511353,I511865,I511882,I511359,I511913,I511347,I511971,I511997,I512014,I511963,I512045,I512053,I512070,I512087,I512104,I512121,I512138,I512155,I511960,I512186,I512203,I512220,I511945,I511957,I512265,I512282,I511951,I512313,I512330,I511939,I512361,I512378,I512395,I512421,I512429,I511948,I512460,I512477,I511954,I512508,I511942,I512566,I1213410,I512592,I512609,I1213425,I512640,I512648,I1213434,I512665,I512682,I1213413,I512699,I1213419,I512716,I512733,I512750,I512781,I1213431,I512798,I1213428,I512815,I512860,I512877,I512908,I512925,I512956,I1213422,I512973,I1213416,I512990,I513016,I513024,I513055,I513072,I513103,I513161,I513187,I513204,I513235,I513243,I513260,I513277,I513294,I513311,I513328,I513345,I513376,I513393,I513410,I513455,I513472,I513503,I513520,I513551,I513568,I513585,I513611,I513619,I513650,I513667,I513698,I513756,I1377902,I513782,I513799,I513748,I1377908,I513830,I513838,I1377923,I513855,I513872,I1377914,I513889,I1377911,I513906,I513923,I513940,I513745,I513971,I513988,I1377926,I514005,I513730,I513742,I514050,I514067,I513736,I514098,I1377920,I514115,I513724,I514146,I1377905,I514163,I1377917,I514180,I1377929,I514206,I514214,I513733,I514245,I514262,I513739,I514293,I513727,I514351,I514377,I514394,I514425,I514433,I514450,I514467,I514484,I514501,I514518,I514535,I514566,I514583,I514600,I514645,I514662,I514693,I514710,I514741,I514758,I514775,I514801,I514809,I514840,I514857,I514888,I514946,I514972,I514989,I514938,I515020,I515028,I515045,I515062,I515079,I515096,I515113,I515130,I514935,I515161,I515178,I515195,I514920,I514932,I515240,I515257,I514926,I515288,I515305,I514914,I515336,I515353,I515370,I515396,I515404,I514923,I515435,I515452,I514929,I515483,I514917,I515541,I682169,I515567,I515584,I515533,I682163,I515615,I515623,I682160,I515640,I515657,I682172,I515674,I682175,I515691,I515708,I515725,I515530,I515756,I682184,I515773,I682178,I515790,I515515,I515527,I515835,I515852,I515521,I515883,I682166,I515900,I515509,I515931,I682181,I515948,I515965,I515991,I515999,I515518,I516030,I516047,I515524,I516078,I515512,I516136,I910842,I516162,I516179,I516128,I910830,I516210,I516218,I910827,I516235,I516252,I910839,I516269,I910836,I516286,I516303,I516320,I516125,I516351,I910845,I516368,I910848,I516385,I516110,I516122,I516430,I516447,I516116,I516478,I910851,I516495,I516104,I516526,I910854,I516543,I910833,I516560,I516586,I516594,I516113,I516625,I516642,I516119,I516673,I516107,I516731,I1327327,I516757,I516774,I516723,I1327333,I516805,I516813,I1327348,I516830,I516847,I1327339,I516864,I1327336,I516881,I516898,I516915,I516720,I516946,I516963,I1327351,I516980,I516705,I516717,I517025,I517042,I516711,I517073,I1327345,I517090,I516699,I517121,I1327330,I517138,I1327342,I517155,I1327354,I517181,I517189,I516708,I517220,I517237,I516714,I517268,I516702,I517326,I1318402,I517352,I517369,I517318,I1318408,I517400,I517408,I1318423,I517425,I517442,I1318414,I517459,I1318411,I517476,I517493,I517510,I517315,I517541,I517558,I1318426,I517575,I517300,I517312,I517620,I517637,I517306,I517668,I1318420,I517685,I517294,I517716,I1318405,I517733,I1318417,I517750,I1318429,I517776,I517784,I517303,I517815,I517832,I517309,I517863,I517297,I517921,I1183814,I517947,I517964,I1183796,I517995,I518003,I1183802,I518020,I518037,I1183817,I518054,I1183808,I518071,I518088,I518105,I518136,I1183820,I518153,I1183799,I518170,I518215,I518232,I518263,I1183805,I518280,I518311,I1183811,I518328,I518345,I518371,I518379,I518410,I518427,I518458,I518516,I1237346,I518542,I518559,I518508,I1237361,I518590,I518598,I1237370,I518615,I518632,I1237349,I518649,I1237355,I518666,I518683,I518700,I518505,I518731,I1237367,I518748,I1237364,I518765,I518490,I518502,I518810,I518827,I518496,I518858,I518875,I518484,I518906,I1237358,I518923,I1237352,I518940,I518966,I518974,I518493,I519005,I519022,I518499,I519053,I518487,I519111,I519137,I519154,I519103,I519185,I519193,I519210,I519227,I519244,I519261,I519278,I519295,I519100,I519326,I519343,I519360,I519085,I519097,I519405,I519422,I519091,I519453,I519470,I519079,I519501,I519518,I519535,I519561,I519569,I519088,I519600,I519617,I519094,I519648,I519082,I519706,I665407,I519732,I519749,I665401,I519780,I519788,I665398,I519805,I519822,I665410,I519839,I665413,I519856,I519873,I519890,I519921,I665422,I519938,I665416,I519955,I520000,I520017,I520048,I665404,I520065,I520096,I665419,I520113,I520130,I520156,I520164,I520195,I520212,I520243,I520301,I520327,I520344,I520293,I520375,I520383,I520400,I520417,I520434,I520451,I520468,I520485,I520290,I520516,I520533,I520550,I520275,I520287,I520595,I520612,I520281,I520643,I520660,I520269,I520691,I520708,I520725,I520751,I520759,I520278,I520790,I520807,I520284,I520838,I520272,I520896,I520922,I520939,I520888,I520970,I520978,I520995,I521012,I521029,I521046,I521063,I521080,I520885,I521111,I521128,I521145,I520870,I520882,I521190,I521207,I520876,I521238,I521255,I520864,I521286,I521303,I521320,I521346,I521354,I520873,I521385,I521402,I520879,I521433,I520867,I521491,I521517,I521534,I521565,I521573,I521590,I521607,I521624,I521641,I521658,I521675,I521706,I521723,I521740,I521785,I521802,I521833,I521850,I521881,I521898,I521915,I521941,I521949,I521980,I521997,I522028,I522086,I522112,I522129,I522160,I522168,I522185,I522202,I522219,I522236,I522253,I522270,I522301,I522318,I522335,I522380,I522397,I522428,I522445,I522476,I522493,I522510,I522536,I522544,I522575,I522592,I522623,I522681,I522707,I522724,I522673,I522755,I522763,I522780,I522797,I522814,I522831,I522848,I522865,I522670,I522896,I522913,I522930,I522655,I522667,I522975,I522992,I522661,I523023,I523040,I522649,I523071,I523088,I523105,I523131,I523139,I522658,I523170,I523187,I522664,I523218,I522652,I523276,I714537,I523302,I523319,I714531,I523350,I523358,I714528,I523375,I523392,I714540,I523409,I714543,I523426,I523443,I523460,I523491,I714552,I523508,I714546,I523525,I523570,I523587,I523618,I714534,I523635,I523666,I714549,I523683,I523700,I523726,I523734,I523765,I523782,I523813,I523871,I547489,I523897,I523914,I547501,I523945,I523953,I547486,I523970,I523987,I547504,I524004,I547495,I524021,I524038,I524055,I524086,I547507,I524103,I547510,I524120,I524165,I524182,I524213,I524230,I524261,I547498,I524278,I547492,I524295,I524321,I524329,I524360,I524377,I524408,I524466,I524492,I524509,I524540,I524548,I524565,I524582,I524599,I524616,I524633,I524650,I524681,I524698,I524715,I524760,I524777,I524808,I524825,I524856,I524873,I524890,I524916,I524924,I524955,I524972,I525003,I525061,I678701,I525087,I525104,I678695,I525135,I525143,I678692,I525160,I525177,I678704,I525194,I678707,I525211,I525228,I525245,I525276,I678716,I525293,I678710,I525310,I525355,I525372,I525403,I678698,I525420,I525451,I678713,I525468,I525485,I525511,I525519,I525550,I525567,I525598,I525656,I1048850,I525682,I525699,I1048853,I525730,I525738,I1048856,I525755,I525772,I1048868,I525789,I1048859,I525806,I525823,I525840,I525871,I1048865,I525888,I525905,I525950,I525967,I525998,I526015,I526046,I1048862,I526063,I526080,I1048871,I526106,I526114,I526145,I526162,I526193,I526251,I526277,I526294,I526325,I526333,I526350,I526367,I526384,I526401,I526418,I526435,I526466,I526483,I526500,I526545,I526562,I526593,I526610,I526641,I526658,I526675,I526701,I526709,I526740,I526757,I526788,I526846,I526872,I526889,I526920,I526928,I526945,I526962,I526979,I526996,I527013,I527030,I527061,I527078,I527095,I527140,I527157,I527188,I527205,I527236,I527253,I527270,I527296,I527304,I527335,I527352,I527383,I527441,I527467,I527484,I527433,I527515,I527523,I527540,I527557,I527574,I527591,I527608,I527625,I527430,I527656,I527673,I527690,I527415,I527427,I527735,I527752,I527421,I527783,I527800,I527409,I527831,I527848,I527865,I527891,I527899,I527418,I527930,I527947,I527424,I527978,I527412,I528036,I1019117,I528062,I528079,I528028,I1019120,I528110,I528118,I1019123,I528135,I528152,I1019135,I528169,I1019126,I528186,I528203,I528220,I528025,I528251,I1019132,I528268,I528285,I528010,I528022,I528330,I528347,I528016,I528378,I528395,I528004,I528426,I1019129,I528443,I528460,I1019138,I528486,I528494,I528013,I528525,I528542,I528019,I528573,I528007,I528631,I528657,I528674,I528623,I528705,I528713,I528730,I528747,I528764,I528781,I528798,I528815,I528620,I528846,I528863,I528880,I528605,I528617,I528925,I528942,I528611,I528973,I528990,I528599,I529021,I529038,I529055,I529081,I529089,I528608,I529120,I529137,I528614,I529168,I528602,I529226,I1235714,I529252,I529269,I529218,I1235729,I529300,I529308,I1235738,I529325,I529342,I1235717,I529359,I1235723,I529376,I529393,I529410,I529215,I529441,I1235735,I529458,I1235732,I529475,I529200,I529212,I529520,I529537,I529206,I529568,I529585,I529194,I529616,I1235726,I529633,I1235720,I529650,I529676,I529684,I529203,I529715,I529732,I529209,I529763,I529197,I529821,I529847,I529864,I529895,I529903,I529920,I529937,I529954,I529971,I529988,I530005,I530036,I530053,I530070,I530115,I530132,I530163,I530180,I530211,I530228,I530245,I530271,I530279,I530310,I530327,I530358,I530416,I1176878,I530442,I530459,I530408,I1176860,I530490,I530498,I1176866,I530515,I530532,I1176881,I530549,I1176872,I530566,I530583,I530600,I530405,I530631,I1176884,I530648,I1176863,I530665,I530390,I530402,I530710,I530727,I530396,I530758,I1176869,I530775,I530384,I530806,I1176875,I530823,I530840,I530866,I530874,I530393,I530905,I530922,I530399,I530953,I530387,I531011,I1057265,I531037,I531054,I531003,I1057268,I531085,I531093,I1057271,I531110,I531127,I1057283,I531144,I1057274,I531161,I531178,I531195,I531000,I531226,I1057280,I531243,I531260,I530985,I530997,I531305,I531322,I530991,I531353,I531370,I530979,I531401,I1057277,I531418,I531435,I1057286,I531461,I531469,I530988,I531500,I531517,I530994,I531548,I530982,I531606,I1047167,I531632,I531649,I531598,I1047170,I531680,I531688,I1047173,I531705,I531722,I1047185,I531739,I1047176,I531756,I531773,I531790,I531595,I531821,I1047182,I531838,I531855,I531580,I531592,I531900,I531917,I531586,I531948,I531965,I531574,I531996,I1047179,I532013,I532030,I1047188,I532056,I532064,I531583,I532095,I532112,I531589,I532143,I531577,I532201,I1391587,I532227,I532244,I532193,I1391593,I532275,I532283,I1391608,I532300,I532317,I1391599,I532334,I1391596,I532351,I532368,I532385,I532190,I532416,I532433,I1391611,I532450,I532175,I532187,I532495,I532512,I532181,I532543,I1391605,I532560,I532169,I532591,I1391590,I532608,I1391602,I532625,I1391614,I532651,I532659,I532178,I532690,I532707,I532184,I532738,I532172,I532796,I532822,I532839,I532788,I532870,I532878,I532895,I532912,I532929,I532946,I532963,I532980,I532785,I533011,I533028,I533045,I532770,I532782,I533090,I533107,I532776,I533138,I533155,I532764,I533186,I533203,I533220,I533246,I533254,I532773,I533285,I533302,I532779,I533333,I532767,I533391,I533417,I533434,I533383,I533465,I533473,I533490,I533507,I533524,I533541,I533558,I533575,I533380,I533606,I533623,I533640,I533365,I533377,I533685,I533702,I533371,I533733,I533750,I533359,I533781,I533798,I533815,I533841,I533849,I533368,I533880,I533897,I533374,I533928,I533362,I533986,I534012,I534029,I534060,I534068,I534085,I534102,I534119,I534136,I534153,I534170,I534201,I534218,I534235,I534280,I534297,I534328,I534345,I534376,I534393,I534410,I534436,I534444,I534475,I534492,I534523,I534581,I620895,I534607,I534624,I534573,I620907,I534655,I534663,I620892,I534680,I534697,I620910,I534714,I620901,I534731,I534748,I534765,I534570,I534796,I620913,I534813,I620916,I534830,I534555,I534567,I534875,I534892,I534561,I534923,I534940,I534549,I534971,I620904,I534988,I620898,I535005,I535031,I535039,I534558,I535070,I535087,I534564,I535118,I534552,I535176,I633617,I535202,I535219,I535168,I633611,I535250,I535258,I633608,I535275,I535292,I633620,I535309,I633623,I535326,I535343,I535360,I535165,I535391,I633632,I535408,I633626,I535425,I535150,I535162,I535470,I535487,I535156,I535518,I633614,I535535,I535144,I535566,I633629,I535583,I535600,I535626,I535634,I535153,I535665,I535682,I535159,I535713,I535147,I535771,I1016312,I535797,I535814,I1016315,I535845,I535853,I1016318,I535870,I535887,I1016330,I535904,I1016321,I535921,I535938,I535955,I535986,I1016327,I536003,I536020,I536065,I536082,I536113,I536130,I536161,I1016324,I536178,I536195,I1016333,I536221,I536229,I536260,I536277,I536308,I536366,I536392,I536409,I536440,I536448,I536465,I536482,I536499,I536516,I536533,I536550,I536581,I536598,I536615,I536660,I536677,I536708,I536725,I536756,I536773,I536790,I536816,I536824,I536855,I536872,I536903,I536961,I1019678,I536987,I537004,I1019681,I537035,I537043,I1019684,I537060,I537077,I1019696,I537094,I1019687,I537111,I537128,I537145,I537176,I1019693,I537193,I537210,I537255,I537272,I537303,I537320,I537351,I1019690,I537368,I537385,I1019699,I537411,I537419,I537450,I537467,I537498,I537556,I537582,I537599,I537548,I537630,I537638,I537655,I537672,I537689,I537706,I537723,I537740,I537545,I537771,I537788,I537805,I537530,I537542,I537850,I537867,I537536,I537898,I537915,I537524,I537946,I537963,I537980,I538006,I538014,I537533,I538045,I538062,I537539,I538093,I537527,I538151,I1115032,I538177,I538194,I538143,I1115014,I538225,I538233,I1115020,I538250,I538267,I1115035,I538284,I1115026,I538301,I538318,I538335,I538140,I538366,I1115038,I538383,I1115017,I538400,I538125,I538137,I538445,I538462,I538131,I538493,I1115023,I538510,I538119,I538541,I1115029,I538558,I538575,I538601,I538609,I538128,I538640,I538657,I538134,I538688,I538122,I538746,I538772,I538789,I538738,I538820,I538828,I538845,I538862,I538879,I538896,I538913,I538930,I538735,I538961,I538978,I538995,I538720,I538732,I539040,I539057,I538726,I539088,I539105,I538714,I539136,I539153,I539170,I539196,I539204,I538723,I539235,I539252,I538729,I539283,I538717,I539341,I1254210,I539367,I539384,I539333,I1254225,I539415,I539423,I1254234,I539440,I539457,I1254213,I539474,I1254219,I539491,I539508,I539525,I539330,I539556,I1254231,I539573,I1254228,I539590,I539315,I539327,I539635,I539652,I539321,I539683,I539700,I539309,I539731,I1254222,I539748,I1254216,I539765,I539791,I539799,I539318,I539830,I539847,I539324,I539878,I539312,I539936,I539962,I539979,I539928,I540010,I540018,I540035,I540052,I540069,I540086,I540103,I540120,I539925,I540151,I540168,I540185,I539910,I539922,I540230,I540247,I539916,I540278,I540295,I539904,I540326,I540343,I540360,I540386,I540394,I539913,I540425,I540442,I539919,I540473,I539907,I540531,I1020239,I540557,I540574,I540523,I1020242,I540605,I540613,I1020245,I540630,I540647,I1020257,I540664,I1020248,I540681,I540698,I540715,I540520,I540746,I1020254,I540763,I540780,I540505,I540517,I540825,I540842,I540511,I540873,I540890,I540499,I540921,I1020251,I540938,I540955,I1020260,I540981,I540989,I540508,I541020,I541037,I540514,I541068,I540502,I541126,I841255,I541152,I541169,I841252,I541200,I541208,I541225,I541242,I841249,I541259,I841264,I541276,I541293,I541310,I541341,I841258,I541358,I841246,I541375,I541420,I541437,I541468,I841267,I541485,I541516,I541533,I841261,I541550,I541576,I541584,I541615,I541632,I541663,I541721,I609913,I541747,I541764,I541713,I609925,I541795,I541803,I609910,I541820,I541837,I609928,I541854,I609919,I541871,I541888,I541905,I541710,I541936,I609931,I541953,I609934,I541970,I541695,I541707,I542015,I542032,I541701,I542063,I542080,I541689,I542111,I609922,I542128,I609916,I542145,I542171,I542179,I541698,I542210,I542227,I541704,I542258,I541692,I542316,I936027,I542342,I542350,I936024,I542376,I542384,I936021,I542401,I936048,I542418,I542435,I936036,I542452,I542483,I542500,I542517,I936042,I542534,I936033,I542579,I542624,I936030,I542641,I542658,I542689,I936045,I542706,I936039,I542723,I542749,I542757,I542802,I542819,I542836,I542894,I542920,I542928,I542954,I542962,I542979,I542996,I543013,I543030,I543061,I543078,I543095,I543112,I543157,I543202,I543219,I543236,I543267,I543284,I543301,I543327,I543335,I543380,I543397,I543414,I543472,I1117904,I543498,I543506,I1117910,I543532,I543540,I543557,I1117907,I543574,I543591,I1117925,I543608,I543458,I543639,I543656,I543673,I1117928,I543690,I543455,I543446,I543735,I543449,I543443,I543780,I1117913,I543797,I543814,I543452,I543845,I1117919,I543862,I1117916,I543879,I1117922,I543905,I543913,I543440,I543464,I543958,I543975,I543992,I543461,I544050,I1169346,I544076,I544084,I1169352,I544110,I544118,I544135,I1169349,I544152,I544169,I1169367,I544186,I544036,I544217,I544234,I544251,I1169370,I544268,I544033,I544024,I544313,I544027,I544021,I544358,I1169355,I544375,I544392,I544030,I544423,I1169361,I544440,I1169358,I544457,I1169364,I544483,I544491,I544018,I544042,I544536,I544553,I544570,I544039,I544628,I1082068,I544654,I544662,I1082074,I544688,I544696,I544713,I1082071,I544730,I544747,I1082089,I544764,I544614,I544795,I544812,I544829,I1082092,I544846,I544611,I544602,I544891,I544605,I544599,I544936,I1082077,I544953,I544970,I544608,I545001,I1082083,I545018,I1082080,I545035,I1082086,I545061,I545069,I544596,I544620,I545114,I545131,I545148,I544617,I545206,I639388,I545232,I545240,I639400,I545266,I545274,I639391,I545291,I639394,I545308,I545325,I639397,I545342,I545373,I545390,I545407,I545424,I639403,I545469,I545514,I639409,I545531,I545548,I545579,I545596,I639406,I545613,I639412,I545639,I545647,I545692,I545709,I545726,I545784,I545810,I545818,I545844,I545852,I545869,I545886,I545903,I545920,I545951,I545968,I545985,I546002,I546047,I546092,I546109,I546126,I546157,I546174,I546191,I546217,I546225,I546270,I546287,I546304,I546362,I710482,I546388,I546396,I710494,I546422,I546430,I710485,I546447,I710488,I546464,I546481,I710491,I546498,I546348,I546529,I546546,I546563,I546580,I710497,I546345,I546336,I546625,I546339,I546333,I546670,I710503,I546687,I546704,I546342,I546735,I546752,I710500,I546769,I710506,I546795,I546803,I546330,I546354,I546848,I546865,I546882,I546351,I546940,I1292336,I546966,I546974,I1292348,I547000,I547008,I1292339,I547025,I1292327,I547042,I547059,I1292324,I547076,I546926,I547107,I547124,I547141,I1292330,I547158,I546923,I546914,I547203,I546917,I546911,I547248,I1292345,I547265,I547282,I546920,I547313,I1292333,I547330,I547347,I1292342,I547373,I547381,I546908,I546932,I547426,I547443,I547460,I546929,I547518,I1262280,I547544,I547552,I1262292,I547578,I547586,I1262283,I547603,I1262271,I547620,I547637,I1262268,I547654,I547685,I547702,I547719,I1262274,I547736,I547781,I547826,I1262289,I547843,I547860,I547891,I1262277,I547908,I547925,I1262286,I547951,I547959,I548004,I548021,I548038,I548096,I776374,I548122,I548130,I776386,I548156,I548164,I776377,I548181,I776380,I548198,I548215,I776383,I548232,I548263,I548280,I548297,I548314,I776389,I548359,I548404,I776395,I548421,I548438,I548469,I548486,I776392,I548503,I776398,I548529,I548537,I548582,I548599,I548616,I548674,I548700,I548708,I548734,I548742,I548759,I548776,I548793,I548810,I548841,I548858,I548875,I548892,I548937,I548982,I548999,I549016,I549047,I549064,I549081,I549107,I549115,I549160,I549177,I549194,I549252,I834401,I549278,I549286,I549312,I549320,I834398,I549337,I834413,I549354,I549371,I834407,I549388,I549419,I549436,I549453,I834404,I549470,I834395,I549515,I549560,I834416,I549577,I549594,I549625,I549642,I549659,I834410,I549685,I549693,I549738,I549755,I549772,I549830,I641122,I549856,I549864,I641134,I549890,I549898,I641125,I549915,I641128,I549932,I549949,I641131,I549966,I549997,I550014,I550031,I550048,I641137,I550093,I550138,I641143,I550155,I550172,I550203,I550220,I641140,I550237,I641146,I550263,I550271,I550316,I550333,I550350,I550408,I1039334,I550434,I550442,I1039325,I550468,I550476,I1039319,I550493,I1039331,I550510,I550527,I1039322,I550544,I550394,I550575,I550592,I550609,I1039328,I550626,I1039313,I550391,I550382,I550671,I550385,I550379,I550716,I550733,I550750,I550388,I550781,I1039316,I550798,I550815,I550841,I550849,I550376,I550400,I550894,I550911,I550928,I550397,I550986,I1004503,I551012,I551020,I1004500,I551046,I551054,I1004497,I551071,I1004524,I551088,I551105,I1004512,I551122,I550972,I551153,I551170,I551187,I1004518,I551204,I1004509,I550969,I550960,I551249,I550963,I550957,I551294,I1004506,I551311,I551328,I550966,I551359,I1004521,I551376,I1004515,I551393,I551419,I551427,I550954,I550978,I551472,I551489,I551506,I550975,I551564,I551590,I551598,I551624,I551632,I551649,I551666,I551683,I551700,I551731,I551748,I551765,I551782,I551827,I551872,I551889,I551906,I551937,I551954,I551971,I551997,I552005,I552050,I552067,I552084,I552142,I737070,I552168,I552176,I737082,I552202,I552210,I737073,I552227,I737076,I552244,I552261,I737079,I552278,I552128,I552309,I552326,I552343,I552360,I737085,I552125,I552116,I552405,I552119,I552113,I552450,I737091,I552467,I552484,I552122,I552515,I552532,I737088,I552549,I737094,I552575,I552583,I552110,I552134,I552628,I552645,I552662,I552131,I552720,I552746,I552754,I552780,I552788,I552805,I552822,I552839,I552856,I552706,I552887,I552904,I552921,I552938,I552703,I552694,I552983,I552697,I552691,I553028,I553045,I553062,I552700,I553093,I553110,I553127,I553153,I553161,I552688,I552712,I553206,I553223,I553240,I552709,I553298,I553324,I553332,I553358,I553366,I553383,I553400,I553417,I553434,I553465,I553482,I553499,I553516,I553561,I553606,I553623,I553640,I553671,I553688,I553705,I553731,I553739,I553784,I553801,I553818,I553876,I1170502,I553902,I553910,I1170508,I553936,I553944,I553961,I1170505,I553978,I553995,I1170523,I554012,I554043,I554060,I554077,I1170526,I554094,I554139,I554184,I1170511,I554201,I554218,I554249,I1170517,I554266,I1170514,I554283,I1170520,I554309,I554317,I554362,I554379,I554396,I554454,I1125418,I554480,I554488,I1125424,I554514,I554522,I554539,I1125421,I554556,I554573,I1125439,I554590,I554621,I554638,I554655,I1125442,I554672,I554717,I554762,I1125427,I554779,I554796,I554827,I1125433,I554844,I1125430,I554861,I1125436,I554887,I554895,I554940,I554957,I554974,I555032,I1045505,I555058,I555066,I1045496,I555092,I555100,I1045490,I555117,I1045502,I555134,I555151,I1045493,I555168,I555018,I555199,I555216,I555233,I1045499,I555250,I1045484,I555015,I555006,I555295,I555009,I555003,I555340,I555357,I555374,I555012,I555405,I1045487,I555422,I555439,I555465,I555473,I555000,I555024,I555518,I555535,I555552,I555021,I555610,I1122528,I555636,I555644,I1122534,I555670,I555678,I555695,I1122531,I555712,I555729,I1122549,I555746,I555596,I555777,I555794,I555811,I1122552,I555828,I555593,I555584,I555873,I555587,I555581,I555918,I1122537,I555935,I555952,I555590,I555983,I1122543,I556000,I1122540,I556017,I1122546,I556043,I556051,I555578,I555602,I556096,I556113,I556130,I555599,I556188,I1211796,I556214,I556222,I1211790,I556248,I556256,I1211799,I556273,I1211778,I556290,I556307,I1211787,I556324,I556174,I556355,I556372,I556389,I1211802,I556406,I1211781,I556171,I556162,I556451,I556165,I556159,I556496,I1211784,I556513,I556530,I556168,I556561,I1211793,I556578,I556595,I556621,I556629,I556156,I556180,I556674,I556691,I556708,I556177,I556766,I556792,I556800,I556826,I556834,I556851,I556868,I556885,I556902,I556752,I556933,I556950,I556967,I556984,I556749,I556740,I557029,I556743,I556737,I557074,I557091,I557108,I556746,I557139,I557156,I557173,I557199,I557207,I556734,I556758,I557252,I557269,I557286,I556755,I557344,I557370,I557378,I557404,I557412,I557429,I557446,I557463,I557480,I557511,I557528,I557545,I557562,I557607,I557652,I557669,I557686,I557717,I557734,I557751,I557777,I557785,I557830,I557847,I557864,I557922,I557948,I557956,I557982,I557990,I558007,I558024,I558041,I558058,I557908,I558089,I558106,I558123,I558140,I557905,I557896,I558185,I557899,I557893,I558230,I558247,I558264,I557902,I558295,I558312,I558329,I558355,I558363,I557890,I557914,I558408,I558425,I558442,I557911,I558500,I762502,I558526,I558534,I762514,I558560,I558568,I762505,I558585,I762508,I558602,I558619,I762511,I558636,I558486,I558667,I558684,I558701,I558718,I762517,I558483,I558474,I558763,I558477,I558471,I558808,I762523,I558825,I558842,I558480,I558873,I558890,I762520,I558907,I762526,I558933,I558941,I558468,I558492,I558986,I559003,I559020,I558489,I559078,I559104,I559112,I559138,I559146,I559163,I559180,I559197,I559214,I559064,I559245,I559262,I559279,I559296,I559061,I559052,I559341,I559055,I559049,I559386,I559403,I559420,I559058,I559451,I559468,I559485,I559511,I559519,I559046,I559070,I559564,I559581,I559598,I559067,I559656,I559682,I559690,I559716,I559724,I559741,I559758,I559775,I559792,I559642,I559823,I559840,I559857,I559874,I559639,I559630,I559919,I559633,I559627,I559964,I559981,I559998,I559636,I560029,I560046,I560063,I560089,I560097,I559624,I559648,I560142,I560159,I560176,I559645,I560234,I793295,I560260,I560268,I560294,I560302,I793292,I560319,I793307,I560336,I560353,I793301,I560370,I560220,I560401,I560418,I560435,I793298,I560452,I793289,I560217,I560208,I560497,I560211,I560205,I560542,I793310,I560559,I560576,I560214,I560607,I560624,I560641,I793304,I560667,I560675,I560202,I560226,I560720,I560737,I560754,I560223,I560812,I560838,I560846,I560872,I560880,I560897,I560914,I560931,I560948,I560979,I560996,I561013,I561030,I561075,I561120,I561137,I561154,I561185,I561202,I561219,I561245,I561253,I561298,I561315,I561332,I561390,I561416,I561424,I561450,I561458,I561475,I561492,I561509,I561526,I561376,I561557,I561574,I561591,I561608,I561373,I561364,I561653,I561367,I561361,I561698,I561715,I561732,I561370,I561763,I561780,I561797,I561823,I561831,I561358,I561382,I561876,I561893,I561910,I561379,I561968,I561994,I562002,I562028,I562036,I562053,I562070,I562087,I562104,I562135,I562152,I562169,I562186,I562231,I562276,I562293,I562310,I562341,I562358,I562375,I562401,I562409,I562454,I562471,I562488,I562546,I881831,I562572,I562580,I562606,I562614,I881828,I562631,I881843,I562648,I562665,I881837,I562682,I562713,I562730,I562747,I881834,I562764,I881825,I562809,I562854,I881846,I562871,I562888,I562919,I562936,I562953,I881840,I562979,I562987,I563032,I563049,I563066,I563124,I563150,I563158,I563184,I563192,I563209,I563226,I563243,I563260,I563110,I563291,I563308,I563325,I563342,I563107,I563098,I563387,I563101,I563095,I563432,I563449,I563466,I563104,I563497,I563514,I563531,I563557,I563565,I563092,I563116,I563610,I563627,I563644,I563113,I563702,I734758,I563728,I563736,I734770,I563762,I563770,I734761,I563787,I734764,I563804,I563821,I734767,I563838,I563869,I563886,I563903,I563920,I734773,I563965,I564010,I734779,I564027,I564044,I564075,I564092,I734776,I564109,I734782,I564135,I564143,I564188,I564205,I564222,I564280,I1098252,I564306,I564314,I1098258,I564340,I564348,I564365,I1098255,I564382,I564399,I1098273,I564416,I564447,I564464,I564481,I1098276,I564498,I564543,I564588,I1098261,I564605,I564622,I564653,I1098267,I564670,I1098264,I564687,I1098270,I564713,I564721,I564766,I564783,I564800,I564858,I564884,I564892,I564918,I564926,I564943,I564960,I564977,I564994,I565025,I565042,I565059,I565076,I565121,I565166,I565183,I565200,I565231,I565248,I565265,I565291,I565299,I565344,I565361,I565378,I565436,I698344,I565462,I565470,I698356,I565496,I565504,I698347,I565521,I698350,I565538,I565555,I698353,I565572,I565603,I565620,I565637,I565654,I698359,I565699,I565744,I698365,I565761,I565778,I565809,I565826,I698362,I565843,I698368,I565869,I565877,I565922,I565939,I565956,I566014,I914063,I566040,I566048,I914060,I566074,I566082,I914057,I566099,I914084,I566116,I566133,I914072,I566150,I566181,I566198,I566215,I914078,I566232,I914069,I566277,I566322,I914066,I566339,I566356,I566387,I914081,I566404,I914075,I566421,I566447,I566455,I566500,I566517,I566534,I566592,I886931,I566618,I566626,I886928,I566652,I566660,I886925,I566677,I886952,I566694,I566711,I886940,I566728,I566578,I566759,I566776,I566793,I886946,I566810,I886937,I566575,I566566,I566855,I566569,I566563,I566900,I886934,I566917,I566934,I566572,I566965,I886949,I566982,I886943,I566999,I567025,I567033,I566560,I566584,I567078,I567095,I567112,I566581,I567170,I1295804,I567196,I567204,I1295816,I567230,I567238,I1295807,I567255,I1295795,I567272,I567289,I1295792,I567306,I567156,I567337,I567354,I567371,I1295798,I567388,I567153,I567144,I567433,I567147,I567141,I567478,I1295813,I567495,I567512,I567150,I567543,I1295801,I567560,I567577,I1295810,I567603,I567611,I567138,I567162,I567656,I567673,I567690,I567159,I567748,I1050554,I567774,I567782,I1050545,I567808,I567816,I1050539,I567833,I1050551,I567850,I567867,I1050542,I567884,I567915,I567932,I567949,I1050548,I567966,I1050533,I568011,I568056,I568073,I568090,I568121,I1050536,I568138,I568155,I568181,I568189,I568234,I568251,I568268,I568326,I913417,I568352,I568360,I913414,I568386,I568394,I913411,I568411,I913438,I568428,I568445,I913426,I568462,I568312,I568493,I568510,I568527,I913432,I568544,I913423,I568309,I568300,I568589,I568303,I568297,I568634,I913420,I568651,I568668,I568306,I568699,I913435,I568716,I913429,I568733,I568759,I568767,I568294,I568318,I568812,I568829,I568846,I568315,I568904,I568930,I568938,I568964,I568972,I568989,I569006,I569023,I569040,I569071,I569088,I569105,I569122,I569167,I569212,I569229,I569246,I569277,I569294,I569311,I569337,I569345,I569390,I569407,I569424,I569482,I569508,I569516,I569542,I569550,I569567,I569584,I569601,I569618,I569468,I569649,I569666,I569683,I569700,I569465,I569456,I569745,I569459,I569453,I569790,I569807,I569824,I569462,I569855,I569872,I569889,I569915,I569923,I569450,I569474,I569968,I569985,I570002,I569471,I570060,I570086,I570094,I570120,I570128,I570145,I570162,I570179,I570196,I570227,I570244,I570261,I570278,I570323,I570368,I570385,I570402,I570433,I570450,I570467,I570493,I570501,I570546,I570563,I570580,I570638,I570664,I570672,I570698,I570706,I570723,I570740,I570757,I570774,I570624,I570805,I570822,I570839,I570856,I570621,I570612,I570901,I570615,I570609,I570946,I570963,I570980,I570618,I571011,I571028,I571045,I571071,I571079,I570606,I570630,I571124,I571141,I571158,I570627,I571216,I571242,I571250,I571276,I571284,I571301,I571318,I571335,I571352,I571202,I571383,I571400,I571417,I571434,I571199,I571190,I571479,I571193,I571187,I571524,I571541,I571558,I571196,I571589,I571606,I571623,I571649,I571657,I571184,I571208,I571702,I571719,I571736,I571205,I571794,I811740,I571820,I571828,I571854,I571862,I811737,I571879,I811752,I571896,I571913,I811746,I571930,I571780,I571961,I571978,I571995,I811743,I572012,I811734,I571777,I571768,I572057,I571771,I571765,I572102,I811755,I572119,I572136,I571774,I572167,I572184,I572201,I811749,I572227,I572235,I571762,I571786,I572280,I572297,I572314,I571783,I572372,I1363027,I572398,I572406,I572432,I572440,I1363051,I572457,I1363033,I572474,I572491,I1363048,I572508,I572358,I572539,I572556,I572573,I1363030,I572590,I1363039,I572355,I572346,I572635,I572349,I572343,I572680,I1363036,I572697,I572714,I572352,I572745,I1363045,I572762,I1363054,I572779,I1363042,I572805,I572813,I572340,I572364,I572858,I572875,I572892,I572361,I572950,I572976,I572984,I573010,I573018,I573035,I573052,I573069,I573086,I573117,I573134,I573151,I573168,I573213,I573258,I573275,I573292,I573323,I573340,I573357,I573383,I573391,I573436,I573453,I573470,I573528,I573554,I573562,I573588,I573596,I573613,I573630,I573647,I573664,I573695,I573712,I573729,I573746,I573791,I573836,I573853,I573870,I573901,I573918,I573935,I573961,I573969,I574014,I574031,I574048,I574106,I1387422,I574132,I574140,I574166,I574174,I1387446,I574191,I1387428,I574208,I574225,I1387443,I574242,I574092,I574273,I574290,I574307,I1387425,I574324,I1387434,I574089,I574080,I574369,I574083,I574077,I574414,I1387431,I574431,I574448,I574086,I574479,I1387440,I574496,I1387449,I574513,I1387437,I574539,I574547,I574074,I574098,I574592,I574609,I574626,I574095,I574684,I1091316,I574710,I574718,I1091322,I574744,I574752,I574769,I1091319,I574786,I574803,I1091337,I574820,I574851,I574868,I574885,I1091340,I574902,I574947,I574992,I1091325,I575009,I575026,I575057,I1091331,I575074,I1091328,I575091,I1091334,I575117,I575125,I575170,I575187,I575204,I575262,I575288,I575296,I575322,I575330,I575347,I575364,I575381,I575398,I575429,I575446,I575463,I575480,I575525,I575570,I575587,I575604,I575635,I575652,I575669,I575695,I575703,I575748,I575765,I575782,I575840,I1205760,I575866,I575874,I1205766,I575900,I575908,I575925,I1205763,I575942,I575959,I1205781,I575976,I575826,I576007,I576024,I576041,I1205784,I576058,I575823,I575814,I576103,I575817,I575811,I576148,I1205769,I576165,I576182,I575820,I576213,I1205775,I576230,I1205772,I576247,I1205778,I576273,I576281,I575808,I575832,I576326,I576343,I576360,I575829,I576418,I576444,I576452,I576478,I576486,I576503,I576520,I576537,I576554,I576585,I576602,I576619,I576636,I576681,I576726,I576743,I576760,I576791,I576808,I576825,I576851,I576859,I576904,I576921,I576938,I576996,I577022,I577030,I577056,I577064,I577081,I577098,I577115,I577132,I576982,I577163,I577180,I577197,I577214,I576979,I576970,I577259,I576973,I576967,I577304,I577321,I577338,I576976,I577369,I577386,I577403,I577429,I577437,I576964,I576988,I577482,I577499,I577516,I576985,I577574,I577600,I577608,I577634,I577642,I577659,I577676,I577693,I577710,I577560,I577741,I577758,I577775,I577792,I577557,I577548,I577837,I577551,I577545,I577882,I577899,I577916,I577554,I577947,I577964,I577981,I578007,I578015,I577542,I577566,I578060,I578077,I578094,I577563,I578152,I1200558,I578178,I578186,I1200564,I578212,I578220,I578237,I1200561,I578254,I578271,I1200579,I578288,I578319,I578336,I578353,I1200582,I578370,I578415,I578460,I1200567,I578477,I578494,I578525,I1200573,I578542,I1200570,I578559,I1200576,I578585,I578593,I578638,I578655,I578672,I578730,I653260,I578756,I578764,I653272,I578790,I578798,I653263,I578815,I653266,I578832,I578849,I653269,I578866,I578716,I578897,I578914,I578931,I578948,I653275,I578713,I578704,I578993,I578707,I578701,I579038,I653281,I579055,I579072,I578710,I579103,I579120,I653278,I579137,I653284,I579163,I579171,I578698,I578722,I579216,I579233,I579250,I578719,I579308,I579334,I579342,I579368,I579376,I579393,I579410,I579427,I579444,I579294,I579475,I579492,I579509,I579526,I579291,I579282,I579571,I579285,I579279,I579616,I579633,I579650,I579288,I579681,I579698,I579715,I579741,I579749,I579276,I579300,I579794,I579811,I579828,I579297,I579886,I579912,I579920,I579946,I579954,I579971,I579988,I580005,I580022,I579872,I580053,I580070,I580087,I580104,I579869,I579860,I580149,I579863,I579857,I580194,I580211,I580228,I579866,I580259,I580276,I580293,I580319,I580327,I579854,I579878,I580372,I580389,I580406,I579875,I580464,I580490,I580498,I580524,I580532,I580549,I580566,I580583,I580600,I580631,I580648,I580665,I580682,I580727,I580772,I580789,I580806,I580837,I580854,I580871,I580897,I580905,I580950,I580967,I580984,I581042,I581068,I581076,I581102,I581110,I581127,I581144,I581161,I581178,I581028,I581209,I581226,I581243,I581260,I581025,I581016,I581305,I581019,I581013,I581350,I581367,I581384,I581022,I581415,I581432,I581449,I581475,I581483,I581010,I581034,I581528,I581545,I581562,I581031,I581620,I1371952,I581646,I581654,I581680,I581688,I1371976,I581705,I1371958,I581722,I581739,I1371973,I581756,I581787,I581804,I581821,I1371955,I581838,I1371964,I581883,I581928,I1371961,I581945,I581962,I581993,I1371970,I582010,I1371979,I582027,I1371967,I582053,I582061,I582106,I582123,I582140,I582198,I582224,I582232,I582258,I582266,I582283,I582300,I582317,I582334,I582184,I582365,I582382,I582399,I582416,I582181,I582172,I582461,I582175,I582169,I582506,I582523,I582540,I582178,I582571,I582588,I582605,I582631,I582639,I582166,I582190,I582684,I582701,I582718,I582187,I582776,I694876,I582802,I582810,I694888,I582836,I582844,I694879,I582861,I694882,I582878,I582895,I694885,I582912,I582943,I582960,I582977,I582994,I694891,I583039,I583084,I694897,I583101,I583118,I583149,I583166,I694894,I583183,I694900,I583209,I583217,I583262,I583279,I583296,I583354,I583380,I583388,I583414,I583422,I583439,I583456,I583473,I583490,I583340,I583521,I583538,I583555,I583572,I583337,I583328,I583617,I583331,I583325,I583662,I583679,I583696,I583334,I583727,I583744,I583761,I583787,I583795,I583322,I583346,I583840,I583857,I583874,I583343,I583932,I984477,I583958,I583966,I984474,I583992,I584000,I984471,I584017,I984498,I584034,I584051,I984486,I584068,I583918,I584099,I584116,I584133,I984492,I584150,I984483,I583915,I583906,I584195,I583909,I583903,I584240,I984480,I584257,I584274,I583912,I584305,I984495,I584322,I984489,I584339,I584365,I584373,I583900,I583924,I584418,I584435,I584452,I583921,I584510,I584536,I584544,I584570,I584578,I584595,I584612,I584629,I584646,I584677,I584694,I584711,I584728,I584773,I584818,I584835,I584852,I584883,I584900,I584917,I584943,I584951,I584996,I585013,I585030,I585088,I585114,I585122,I585148,I585156,I585173,I585190,I585207,I585224,I585074,I585255,I585272,I585289,I585306,I585071,I585062,I585351,I585065,I585059,I585396,I585413,I585430,I585068,I585461,I585478,I585495,I585521,I585529,I585056,I585080,I585574,I585591,I585608,I585077,I585666,I811213,I585692,I585700,I585726,I585734,I811210,I585751,I811225,I585768,I585785,I811219,I585802,I585652,I585833,I585850,I585867,I811216,I585884,I811207,I585649,I585640,I585929,I585643,I585637,I585974,I811228,I585991,I586008,I585646,I586039,I586056,I586073,I811222,I586099,I586107,I585634,I585658,I586152,I586169,I586186,I585655,I586244,I783809,I586270,I586278,I586304,I586312,I783806,I586329,I783821,I586346,I586363,I783815,I586380,I586230,I586411,I586428,I586445,I783812,I586462,I783803,I586227,I586218,I586507,I586221,I586215,I586552,I783824,I586569,I586586,I586224,I586617,I586634,I586651,I783818,I586677,I586685,I586212,I586236,I586730,I586747,I586764,I586233,I586822,I1255922,I586848,I586856,I1255934,I586882,I586890,I1255925,I586907,I1255913,I586924,I586941,I1255910,I586958,I586989,I587006,I587023,I1255916,I587040,I587085,I587130,I1255931,I587147,I587164,I587195,I1255919,I587212,I587229,I1255928,I587255,I587263,I587308,I587325,I587342,I587400,I743428,I587426,I587434,I743440,I587460,I587468,I743431,I587485,I743434,I587502,I587519,I743437,I587536,I587386,I587567,I587584,I587601,I587618,I743443,I587383,I587374,I587663,I587377,I587371,I587708,I743449,I587725,I587742,I587380,I587773,I587790,I743446,I587807,I743452,I587833,I587841,I587368,I587392,I587886,I587903,I587920,I587389,I587978,I588004,I588012,I588038,I588046,I588063,I588080,I588097,I588114,I587964,I588145,I588162,I588179,I588196,I587961,I587952,I588241,I587955,I587949,I588286,I588303,I588320,I587958,I588351,I588368,I588385,I588411,I588419,I587946,I587970,I588464,I588481,I588498,I587967,I588556,I1128886,I588582,I588590,I1128892,I588616,I588624,I588641,I1128889,I588658,I588675,I1128907,I588692,I588542,I588723,I588740,I588757,I1128910,I588774,I588539,I588530,I588819,I588533,I588527,I588864,I1128895,I588881,I588898,I588536,I588929,I1128901,I588946,I1128898,I588963,I1128904,I588989,I588997,I588524,I588548,I589042,I589059,I589076,I588545,I589134,I589160,I589168,I589194,I589202,I589219,I589236,I589253,I589270,I589301,I589318,I589335,I589352,I589397,I589442,I589459,I589476,I589507,I589524,I589541,I589567,I589575,I589620,I589637,I589654,I589712,I1378497,I589738,I589746,I589772,I589780,I1378521,I589797,I1378503,I589814,I589831,I1378518,I589848,I589698,I589879,I589896,I589913,I1378500,I589930,I1378509,I589695,I589686,I589975,I589689,I589683,I590020,I1378506,I590037,I590054,I589692,I590085,I1378515,I590102,I1378524,I590119,I1378512,I590145,I590153,I589680,I589704,I590198,I590215,I590232,I589701,I590290,I1330897,I590316,I590324,I590350,I590358,I1330921,I590375,I1330903,I590392,I590409,I1330918,I590426,I590457,I590474,I590491,I1330900,I590508,I1330909,I590553,I590598,I1330906,I590615,I590632,I590663,I1330915,I590680,I1330924,I590697,I1330912,I590723,I590731,I590776,I590793,I590810,I590868,I590894,I590902,I590928,I590936,I590953,I590970,I590987,I591004,I591035,I591052,I591069,I591086,I591131,I591176,I591193,I591210,I591241,I591258,I591275,I591301,I591309,I591354,I591371,I591388,I591446,I591472,I591480,I591506,I591514,I591531,I591548,I591565,I591582,I591432,I591613,I591630,I591647,I591664,I591429,I591420,I591709,I591423,I591417,I591754,I591771,I591788,I591426,I591819,I591836,I591853,I591879,I591887,I591414,I591438,I591932,I591949,I591966,I591435,I592024,I592050,I592058,I592084,I592092,I592109,I592126,I592143,I592160,I592191,I592208,I592225,I592242,I592287,I592332,I592349,I592366,I592397,I592414,I592431,I592457,I592465,I592510,I592527,I592544,I592602,I628984,I592628,I592636,I628996,I592662,I592670,I628987,I592687,I628990,I592704,I592721,I628993,I592738,I592588,I592769,I592786,I592803,I592820,I628999,I592585,I592576,I592865,I592579,I592573,I592910,I629005,I592927,I592944,I592582,I592975,I592992,I629002,I593009,I629008,I593035,I593043,I592570,I592594,I593088,I593105,I593122,I592591,I593180,I1281354,I593206,I593214,I1281366,I593240,I593248,I1281357,I593265,I1281345,I593282,I593299,I1281342,I593316,I593166,I593347,I593364,I593381,I1281348,I593398,I593163,I593154,I593443,I593157,I593151,I593488,I1281363,I593505,I593522,I593160,I593553,I1281351,I593570,I593587,I1281360,I593613,I593621,I593148,I593172,I593666,I593683,I593700,I593169,I593758,I884466,I593784,I593792,I593818,I593826,I884463,I593843,I884478,I593860,I593877,I884472,I593894,I593744,I593925,I593942,I593959,I884469,I593976,I884460,I593741,I593732,I594021,I593735,I593729,I594066,I884481,I594083,I594100,I593738,I594131,I594148,I594165,I884475,I594191,I594199,I593726,I593750,I594244,I594261,I594278,I593747,I594336,I663664,I594362,I594370,I663676,I594396,I594404,I663667,I594421,I663670,I594438,I594455,I663673,I594472,I594503,I594520,I594537,I594554,I663679,I594599,I594644,I663685,I594661,I594678,I594709,I594726,I663682,I594743,I663688,I594769,I594777,I594822,I594839,I594856,I594914,I1379092,I594940,I594948,I594974,I594982,I1379116,I594999,I1379098,I595016,I595033,I1379113,I595050,I594900,I595081,I595098,I595115,I1379095,I595132,I1379104,I594897,I594888,I595177,I594891,I594885,I595222,I1379101,I595239,I595256,I594894,I595287,I1379110,I595304,I1379119,I595321,I1379107,I595347,I595355,I594882,I594906,I595400,I595417,I595434,I594903,I595492,I595518,I595526,I595552,I595560,I595577,I595594,I595611,I595628,I595478,I595659,I595676,I595693,I595710,I595475,I595466,I595755,I595469,I595463,I595800,I595817,I595834,I595472,I595865,I595882,I595899,I595925,I595933,I595460,I595484,I595978,I595995,I596012,I595481,I596070,I596096,I596104,I596130,I596138,I596155,I596172,I596189,I596206,I596237,I596254,I596271,I596288,I596333,I596378,I596395,I596412,I596443,I596460,I596477,I596503,I596511,I596556,I596573,I596590,I596648,I1014089,I596674,I596682,I1014080,I596708,I596716,I1014074,I596733,I1014086,I596750,I596767,I1014077,I596784,I596815,I596832,I596849,I1014083,I596866,I1014068,I596911,I596956,I596973,I596990,I597021,I1014071,I597038,I597055,I597081,I597089,I597134,I597151,I597168,I597226,I806997,I597252,I597260,I597286,I597294,I806994,I597311,I807009,I597328,I597345,I807003,I597362,I597393,I597410,I597427,I807000,I597444,I806991,I597489,I597534,I807012,I597551,I597568,I597599,I597616,I597633,I807006,I597659,I597667,I597712,I597729,I597746,I597804,I1206900,I597830,I597838,I1206894,I597864,I597872,I1206903,I597889,I1206882,I597906,I597923,I1206891,I597940,I597971,I597988,I598005,I1206906,I598022,I1206885,I598067,I598112,I1206888,I598129,I598146,I598177,I1206897,I598194,I598211,I598237,I598245,I598290,I598307,I598324,I598382,I852846,I598408,I598416,I598442,I598450,I852843,I598467,I852858,I598484,I598501,I852852,I598518,I598368,I598549,I598566,I598583,I852849,I598600,I852840,I598365,I598356,I598645,I598359,I598353,I598690,I852861,I598707,I598724,I598362,I598755,I598772,I598789,I852855,I598815,I598823,I598350,I598374,I598868,I598885,I598902,I598371,I598960,I1385637,I598986,I598994,I599020,I599028,I1385661,I599045,I1385643,I599062,I599079,I1385658,I599096,I598946,I599127,I599144,I599161,I1385640,I599178,I1385649,I598943,I598934,I599223,I598937,I598931,I599268,I1385646,I599285,I599302,I598940,I599333,I1385655,I599350,I1385664,I599367,I1385652,I599393,I599401,I598928,I598952,I599446,I599463,I599480,I598949,I599538,I1296931,I599564,I599572,I1296949,I599598,I599606,I1296946,I599623,I1296937,I599640,I599657,I1296934,I599674,I599524,I599705,I599722,I599739,I1296940,I599756,I1296955,I599521,I599512,I599801,I599515,I599509,I599846,I599863,I599880,I599518,I599911,I1296952,I599928,I1296943,I599945,I1296958,I599971,I599979,I599506,I599530,I600024,I600041,I600058,I599527,I600116,I973495,I600142,I600150,I973492,I600176,I600184,I973489,I600201,I973516,I600218,I600235,I973504,I600252,I600102,I600283,I600300,I600317,I973510,I600334,I973501,I600099,I600090,I600379,I600093,I600087,I600424,I973498,I600441,I600458,I600096,I600489,I973513,I600506,I973507,I600523,I600549,I600557,I600084,I600108,I600602,I600619,I600636,I600105,I600694,I794349,I600720,I600728,I600754,I600762,I794346,I600779,I794361,I600796,I600813,I794355,I600830,I600861,I600878,I600895,I794352,I600912,I794343,I600957,I601002,I794364,I601019,I601036,I601067,I601084,I601101,I794358,I601127,I601135,I601180,I601197,I601214,I601272,I858643,I601298,I601306,I601332,I601340,I858640,I601357,I858655,I601374,I601391,I858649,I601408,I601439,I601456,I601473,I858646,I601490,I858637,I601535,I601580,I858658,I601597,I601614,I601645,I601662,I601679,I858652,I601705,I601713,I601758,I601775,I601792,I601850,I601876,I601884,I601910,I601918,I601935,I601952,I601969,I601986,I601836,I602017,I602034,I602051,I602068,I601833,I601824,I602113,I601827,I601821,I602158,I602175,I602192,I601830,I602223,I602240,I602257,I602283,I602291,I601818,I601842,I602336,I602353,I602370,I601839,I602428,I1227572,I602454,I602462,I1227566,I602488,I602496,I1227575,I602513,I1227554,I602530,I602547,I1227563,I602564,I602595,I602612,I602629,I1227578,I602646,I1227557,I602691,I602736,I1227560,I602753,I602770,I602801,I1227569,I602818,I602835,I602861,I602869,I602914,I602931,I602948,I603006,I926337,I603032,I603040,I926334,I603066,I603074,I926331,I603091,I926358,I603108,I603125,I926346,I603142,I603173,I603190,I603207,I926352,I603224,I926343,I603269,I603314,I926340,I603331,I603348,I603379,I926355,I603396,I926349,I603413,I603439,I603447,I603492,I603509,I603526,I603584,I603610,I603618,I603644,I603652,I603669,I603686,I603703,I603720,I603751,I603768,I603785,I603802,I603847,I603892,I603909,I603926,I603957,I603974,I603991,I604017,I604025,I604070,I604087,I604104,I604162,I1280198,I604188,I604196,I1280210,I604222,I604230,I1280201,I604247,I1280189,I604264,I604281,I1280186,I604298,I604329,I604346,I604363,I1280192,I604380,I604425,I604470,I1280207,I604487,I604504,I604535,I1280195,I604552,I604569,I1280204,I604595,I604603,I604648,I604665,I604682,I604740,I1383852,I604766,I604774,I604800,I604808,I1383876,I604825,I1383858,I604842,I604859,I1383873,I604876,I604907,I604924,I604941,I1383855,I604958,I1383864,I605003,I605048,I1383861,I605065,I605082,I605113,I1383870,I605130,I1383879,I605147,I1383867,I605173,I605181,I605226,I605243,I605260,I605318,I689096,I605344,I605352,I689108,I605378,I605386,I689099,I605403,I689102,I605420,I605437,I689105,I605454,I605304,I605485,I605502,I605519,I605536,I689111,I605301,I605292,I605581,I605295,I605289,I605626,I689117,I605643,I605660,I605298,I605691,I605708,I689114,I605725,I689120,I605751,I605759,I605286,I605310,I605804,I605821,I605838,I605307,I605896,I605922,I605930,I605956,I605964,I605981,I605998,I606015,I606032,I606063,I606080,I606097,I606114,I606159,I606204,I606221,I606238,I606269,I606286,I606303,I606329,I606337,I606382,I606399,I606416,I606474,I606500,I606508,I606534,I606542,I606559,I606576,I606593,I606610,I606460,I606641,I606658,I606675,I606692,I606457,I606448,I606737,I606451,I606445,I606782,I606799,I606816,I606454,I606847,I606864,I606881,I606907,I606915,I606442,I606466,I606960,I606977,I606994,I606463,I607052,I607078,I607086,I607112,I607120,I607137,I607154,I607171,I607188,I607219,I607236,I607253,I607270,I607315,I607360,I607377,I607394,I607425,I607442,I607459,I607485,I607493,I607538,I607555,I607572,I607630,I1204026,I607656,I607664,I1204032,I607690,I607698,I607715,I1204029,I607732,I607749,I1204047,I607766,I607797,I607814,I607831,I1204050,I607848,I607893,I607938,I1204035,I607955,I607972,I608003,I1204041,I608020,I1204038,I608037,I1204044,I608063,I608071,I608116,I608133,I608150,I608208,I842306,I608234,I608242,I608268,I608276,I842303,I608293,I842318,I608310,I608327,I842312,I608344,I608194,I608375,I608392,I608409,I842309,I608426,I842300,I608191,I608182,I608471,I608185,I608179,I608516,I842321,I608533,I608550,I608188,I608581,I608598,I608615,I842315,I608641,I608649,I608176,I608200,I608694,I608711,I608728,I608197,I608786,I1078022,I608812,I608820,I1078028,I608846,I608854,I608871,I1078025,I608888,I608905,I1078043,I608922,I608953,I608970,I608987,I1078046,I609004,I609049,I609094,I1078031,I609111,I609128,I609159,I1078037,I609176,I1078034,I609193,I1078040,I609219,I609227,I609272,I609289,I609306,I609364,I609390,I609398,I609424,I609432,I609449,I609466,I609483,I609500,I609350,I609531,I609548,I609565,I609582,I609347,I609338,I609627,I609341,I609335,I609672,I609689,I609706,I609344,I609737,I609754,I609771,I609797,I609805,I609332,I609356,I609850,I609867,I609884,I609353,I609942,I609968,I609976,I610002,I610010,I610027,I610044,I610061,I610078,I610109,I610126,I610143,I610160,I610205,I610250,I610267,I610284,I610315,I610332,I610349,I610375,I610383,I610428,I610445,I610462,I610520,I610546,I610554,I610580,I610588,I610605,I610622,I610639,I610656,I610687,I610704,I610721,I610738,I610783,I610828,I610845,I610862,I610893,I610910,I610927,I610953,I610961,I611006,I611023,I611040,I611098,I630718,I611124,I611132,I630730,I611158,I611166,I630721,I611183,I630724,I611200,I611217,I630727,I611234,I611265,I611282,I611299,I611316,I630733,I611361,I611406,I630739,I611423,I611440,I611471,I611488,I630736,I611505,I630742,I611531,I611539,I611584,I611601,I611618,I611676,I1283666,I611702,I611710,I1283678,I611736,I611744,I1283669,I611761,I1283657,I611778,I611795,I1283654,I611812,I611843,I611860,I611877,I1283660,I611894,I611939,I611984,I1283675,I612001,I612018,I612049,I1283663,I612066,I612083,I1283672,I612109,I612117,I612162,I612179,I612196,I612254,I1370167,I612280,I612288,I612314,I612322,I1370191,I612339,I1370173,I612356,I612373,I1370188,I612390,I612240,I612421,I612438,I612455,I1370170,I612472,I1370179,I612237,I612228,I612517,I612231,I612225,I612562,I1370176,I612579,I612596,I612234,I612627,I1370185,I612644,I1370194,I612661,I1370182,I612687,I612695,I612222,I612246,I612740,I612757,I612774,I612243,I612832,I1048310,I612858,I612866,I1048301,I612892,I612900,I1048295,I612917,I1048307,I612934,I612951,I1048298,I612968,I612818,I612999,I613016,I613033,I1048304,I613050,I1048289,I612815,I612806,I613095,I612809,I612803,I613140,I613157,I613174,I612812,I613205,I1048292,I613222,I613239,I613265,I613273,I612800,I612824,I613318,I613335,I613352,I612821,I613410,I1169924,I613436,I613444,I1169930,I613470,I613478,I613495,I1169927,I613512,I613529,I1169945,I613546,I613396,I613577,I613594,I613611,I1169948,I613628,I613393,I613384,I613673,I613387,I613381,I613718,I1169933,I613735,I613752,I613390,I613783,I1169939,I613800,I1169936,I613817,I1169942,I613843,I613851,I613378,I613402,I613896,I613913,I613930,I613399,I613988,I614014,I614022,I614048,I614056,I614073,I614090,I614107,I614124,I613974,I614155,I614172,I614189,I614206,I613971,I613962,I614251,I613965,I613959,I614296,I614313,I614330,I613968,I614361,I614378,I614395,I614421,I614429,I613956,I613980,I614474,I614491,I614508,I613977,I614566,I614592,I614600,I614626,I614634,I614651,I614668,I614685,I614702,I614552,I614733,I614750,I614767,I614784,I614549,I614540,I614829,I614543,I614537,I614874,I614891,I614908,I614546,I614939,I614956,I614973,I614999,I615007,I614534,I614558,I615052,I615069,I615086,I614555,I615144,I954761,I615170,I615178,I954758,I615204,I615212,I954755,I615229,I954782,I615246,I615263,I954770,I615280,I615130,I615311,I615328,I615345,I954776,I615362,I954767,I615127,I615118,I615407,I615121,I615115,I615452,I954764,I615469,I615486,I615124,I615517,I954779,I615534,I954773,I615551,I615577,I615585,I615112,I615136,I615630,I615647,I615664,I615133,I615722,I1389207,I615748,I615756,I615782,I615790,I1389231,I615807,I1389213,I615824,I615841,I1389228,I615858,I615708,I615889,I615906,I615923,I1389210,I615940,I1389219,I615705,I615696,I615985,I615699,I615693,I616030,I1389216,I616047,I616064,I615702,I616095,I1389225,I616112,I1389234,I616129,I1389222,I616155,I616163,I615690,I615714,I616208,I616225,I616242,I615711,I616300,I616326,I616334,I616360,I616368,I616385,I616402,I616419,I616436,I616286,I616467,I616484,I616501,I616518,I616283,I616274,I616563,I616277,I616271,I616608,I616625,I616642,I616280,I616673,I616690,I616707,I616733,I616741,I616268,I616292,I616786,I616803,I616820,I616289,I616878,I1041578,I616904,I616912,I1041569,I616938,I616946,I1041563,I616963,I1041575,I616980,I616997,I1041566,I617014,I616864,I617045,I617062,I617079,I1041572,I617096,I1041557,I616861,I616852,I617141,I616855,I616849,I617186,I617203,I617220,I616858,I617251,I1041560,I617268,I617285,I617311,I617319,I616846,I616870,I617364,I617381,I617398,I616867,I617456,I647480,I617482,I617490,I647492,I617516,I617524,I647483,I617541,I647486,I617558,I617575,I647489,I617592,I617442,I617623,I617640,I617657,I617674,I647495,I617439,I617430,I617719,I617433,I617427,I617764,I647501,I617781,I617798,I617436,I617829,I617846,I647498,I617863,I647504,I617889,I617897,I617424,I617448,I617942,I617959,I617976,I617445,I618034,I732446,I618060,I618068,I732458,I618094,I618102,I732449,I618119,I732452,I618136,I618153,I732455,I618170,I618020,I618201,I618218,I618235,I618252,I732461,I618017,I618008,I618297,I618011,I618005,I618342,I732467,I618359,I618376,I618014,I618407,I618424,I732464,I618441,I732470,I618467,I618475,I618002,I618026,I618520,I618537,I618554,I618023,I618612,I618638,I618646,I618672,I618680,I618697,I618714,I618731,I618748,I618598,I618779,I618796,I618813,I618830,I618595,I618586,I618875,I618589,I618583,I618920,I618937,I618954,I618592,I618985,I619002,I619019,I619045,I619053,I618580,I618604,I619098,I619115,I619132,I618601,I619190,I619216,I619224,I619250,I619258,I619275,I619292,I619309,I619326,I619176,I619357,I619374,I619391,I619408,I619173,I619164,I619453,I619167,I619161,I619498,I619515,I619532,I619170,I619563,I619580,I619597,I619623,I619631,I619158,I619182,I619676,I619693,I619710,I619179,I619768,I753832,I619794,I619802,I753844,I619828,I619836,I753835,I619853,I753838,I619870,I619887,I753841,I619904,I619754,I619935,I619952,I619969,I619986,I753847,I619751,I619742,I620031,I619745,I619739,I620076,I753853,I620093,I620110,I619748,I620141,I620158,I753850,I620175,I753856,I620201,I620209,I619736,I619760,I620254,I620271,I620288,I619757,I620346,I1150272,I620372,I620380,I1150278,I620406,I620414,I620431,I1150275,I620448,I620465,I1150293,I620482,I620513,I620530,I620547,I1150296,I620564,I620609,I620654,I1150281,I620671,I620688,I620719,I1150287,I620736,I1150284,I620753,I1150290,I620779,I620787,I620832,I620849,I620866,I620924,I1362432,I620950,I620958,I620984,I620992,I1362456,I621009,I1362438,I621026,I621043,I1362453,I621060,I621091,I621108,I621125,I1362435,I621142,I1362444,I621187,I621232,I1362441,I621249,I621266,I621297,I1362450,I621314,I1362459,I621331,I1362447,I621357,I621365,I621410,I621427,I621444,I621502,I1231924,I621528,I621536,I1231918,I621562,I621570,I1231927,I621587,I1231906,I621604,I621621,I1231915,I621638,I621669,I621686,I621703,I1231930,I621720,I1231909,I621765,I621810,I1231912,I621827,I621844,I621875,I1231921,I621892,I621909,I621935,I621943,I621988,I622005,I622022,I622080,I622106,I622114,I622140,I622148,I622165,I622182,I622199,I622216,I622066,I622247,I622264,I622281,I622298,I622063,I622054,I622343,I622057,I622051,I622388,I622405,I622422,I622060,I622453,I622470,I622487,I622513,I622521,I622048,I622072,I622566,I622583,I622600,I622069,I622658,I1167612,I622684,I622692,I1167618,I622718,I622726,I622743,I1167615,I622760,I622777,I1167633,I622794,I622644,I622825,I622842,I622859,I1167636,I622876,I622641,I622632,I622921,I622635,I622629,I622966,I1167621,I622983,I623000,I622638,I623031,I1167627,I623048,I1167624,I623065,I1167630,I623091,I623099,I622626,I622650,I623144,I623161,I623178,I622647,I623236,I1370762,I623262,I623270,I623296,I623304,I1370786,I623321,I1370768,I623338,I623355,I1370783,I623372,I623222,I623403,I623420,I623437,I1370765,I623454,I1370774,I623219,I623210,I623499,I623213,I623207,I623544,I1370771,I623561,I623578,I623216,I623609,I1370780,I623626,I1370789,I623643,I1370777,I623669,I623677,I623204,I623228,I623722,I623739,I623756,I623225,I623814,I682738,I623840,I623848,I682750,I623874,I623882,I682741,I623899,I682744,I623916,I623933,I682747,I623950,I623800,I623981,I623998,I624015,I624032,I682753,I623797,I623788,I624077,I623791,I623785,I624122,I682759,I624139,I624156,I623794,I624187,I624204,I682756,I624221,I682762,I624247,I624255,I623782,I623806,I624300,I624317,I624334,I623803,I624392,I838617,I624418,I624426,I624452,I624460,I838614,I624477,I838629,I624494,I624511,I838623,I624528,I624559,I624576,I624593,I838620,I624610,I838611,I624655,I624700,I838632,I624717,I624734,I624765,I624782,I624799,I838626,I624825,I624833,I624878,I624895,I624912,I624970,I1365407,I624996,I625004,I625030,I625038,I1365431,I625055,I1365413,I625072,I625089,I1365428,I625106,I625137,I625154,I625171,I1365410,I625188,I1365419,I625233,I625278,I1365416,I625295,I625312,I625343,I1365425,I625360,I1365434,I625377,I1365422,I625403,I625411,I625456,I625473,I625490,I625548,I977371,I625574,I625582,I977368,I625608,I625616,I977365,I625633,I977392,I625650,I625667,I977380,I625684,I625534,I625715,I625732,I625749,I977386,I625766,I977377,I625531,I625522,I625811,I625525,I625519,I625856,I977374,I625873,I625890,I625528,I625921,I977389,I625938,I977383,I625955,I625981,I625989,I625516,I625540,I626034,I626051,I626068,I625537,I626126,I1201714,I626152,I626160,I1201720,I626186,I626194,I626211,I1201717,I626228,I626245,I1201735,I626262,I626112,I626293,I626310,I626327,I1201738,I626344,I626109,I626100,I626389,I626103,I626097,I626434,I1201723,I626451,I626468,I626106,I626499,I1201729,I626516,I1201726,I626533,I1201732,I626559,I626567,I626094,I626118,I626612,I626629,I626646,I626115,I626704,I626730,I626738,I626764,I626772,I626789,I626806,I626823,I626840,I626690,I626871,I626888,I626905,I626922,I626687,I626678,I626967,I626681,I626675,I627012,I627029,I627046,I626684,I627077,I627094,I627111,I627137,I627145,I626672,I626696,I627190,I627207,I627224,I626693,I627282,I627308,I627316,I627333,I627350,I627376,I627384,I627410,I627418,I627435,I627452,I627469,I627509,I627517,I627534,I627551,I627568,I627599,I627616,I627642,I627650,I627681,I627712,I627729,I627760,I627860,I627886,I627894,I627911,I627928,I627954,I627962,I627988,I627996,I628013,I628030,I628047,I628087,I628095,I628112,I628129,I628146,I628177,I628194,I628220,I628228,I628259,I628290,I628307,I628338,I628438,I628464,I628472,I628489,I628506,I628532,I628540,I628566,I628574,I628591,I628608,I628625,I628665,I628673,I628690,I628707,I628724,I628755,I628772,I628798,I628806,I628837,I628868,I628885,I628916,I629016,I958009,I629042,I629050,I629067,I957985,I958000,I629084,I958012,I629110,I629118,I957997,I957988,I629144,I629152,I629169,I629186,I629203,I629243,I629251,I629268,I629285,I629302,I629333,I958003,I957994,I629350,I958006,I629376,I629384,I629415,I629446,I629463,I629494,I957991,I629594,I1218306,I629620,I629628,I629645,I1218309,I1218318,I629662,I1218321,I629688,I629696,I1218330,I1218312,I629722,I629730,I629747,I629764,I629781,I629577,I629821,I629829,I629846,I629863,I629880,I629580,I629911,I1218327,I629928,I1218324,I629954,I629962,I629562,I629993,I629571,I630024,I630041,I629583,I630072,I1218315,I629574,I629565,I629568,I629586,I630172,I1285388,I630198,I630206,I630223,I1285412,I1285394,I630240,I1285400,I630266,I630274,I1285406,I1285391,I630300,I630308,I630325,I630342,I630359,I630155,I1285403,I630399,I630407,I630424,I630441,I630458,I630158,I630489,I1285409,I1285397,I630506,I630532,I630540,I630140,I630571,I630149,I630602,I630619,I630161,I630650,I630152,I630143,I630146,I630164,I630750,I1215586,I630776,I630784,I630801,I1215589,I1215598,I630818,I1215601,I630844,I630852,I1215610,I1215592,I630878,I630886,I630903,I630920,I630937,I630977,I630985,I631002,I631019,I631036,I631067,I1215607,I631084,I1215604,I631110,I631118,I631149,I631180,I631197,I631228,I1215595,I631328,I1163006,I631354,I631362,I631379,I1162988,I1163000,I631396,I1163003,I631422,I631430,I1162997,I1162994,I631456,I631464,I631481,I631498,I631515,I631311,I1163012,I631555,I631563,I631580,I631597,I631614,I631314,I631645,I1162991,I631662,I631688,I631696,I631296,I631727,I631305,I631758,I631775,I631317,I631806,I1163009,I631308,I631299,I631302,I631320,I631906,I631932,I631940,I631957,I631974,I632000,I632008,I632034,I632042,I632059,I632076,I632093,I631889,I632133,I632141,I632158,I632175,I632192,I631892,I632223,I632240,I632266,I632274,I631874,I632305,I631883,I632336,I632353,I631895,I632384,I631886,I631877,I631880,I631898,I632484,I632510,I632518,I632535,I632552,I632578,I632586,I632612,I632620,I632637,I632654,I632671,I632467,I632711,I632719,I632736,I632753,I632770,I632470,I632801,I632818,I632844,I632852,I632452,I632883,I632461,I632914,I632931,I632473,I632962,I632464,I632455,I632458,I632476,I633062,I633088,I633096,I633113,I633130,I633156,I633164,I633190,I633198,I633215,I633232,I633249,I633289,I633297,I633314,I633331,I633348,I633379,I633396,I633422,I633430,I633461,I633492,I633509,I633540,I633640,I947027,I633666,I633674,I633691,I947003,I947018,I633708,I947030,I633734,I633742,I947015,I947006,I633768,I633776,I633793,I633810,I633827,I633867,I633875,I633892,I633909,I633926,I633957,I947021,I947012,I633974,I947024,I634000,I634008,I634039,I634070,I634087,I634118,I947009,I634218,I1059544,I634244,I634252,I634269,I1059526,I1059538,I634286,I1059541,I634312,I634320,I1059535,I1059532,I634346,I634354,I634371,I634388,I634405,I634201,I1059550,I634445,I634453,I634470,I634487,I634504,I634204,I634535,I1059529,I634552,I634578,I634586,I634186,I634617,I634195,I634648,I634665,I634207,I634696,I1059547,I634198,I634189,I634192,I634210,I634796,I634822,I634830,I634847,I634864,I634890,I634898,I634924,I634932,I634949,I634966,I634983,I635023,I635031,I635048,I635065,I635082,I635113,I635130,I635156,I635164,I635195,I635226,I635243,I635274,I635374,I812803,I635400,I635408,I635425,I812791,I812809,I635442,I812806,I635468,I635476,I812797,I812794,I635502,I635510,I635527,I635544,I635561,I812788,I635601,I635609,I635626,I635643,I635660,I635691,I635708,I635734,I635742,I635773,I635804,I635821,I635852,I812800,I635952,I799628,I635978,I635986,I636003,I799616,I799634,I636020,I799631,I636046,I636054,I799622,I799619,I636080,I636088,I636105,I636122,I636139,I635935,I799613,I636179,I636187,I636204,I636221,I636238,I635938,I636269,I636286,I636312,I636320,I635920,I636351,I635929,I636382,I636399,I635941,I636430,I799625,I635932,I635923,I635926,I635944,I636530,I1107518,I636556,I636564,I636581,I1107500,I1107512,I636598,I1107515,I636624,I636632,I1107509,I1107506,I636658,I636666,I636683,I636700,I636717,I636513,I1107524,I636757,I636765,I636782,I636799,I636816,I636516,I636847,I1107503,I636864,I636890,I636898,I636498,I636929,I636507,I636960,I636977,I636519,I637008,I1107521,I636510,I636501,I636504,I636522,I637108,I1284810,I637134,I637142,I637159,I1284834,I1284816,I637176,I1284822,I637202,I637210,I1284828,I1284813,I637236,I637244,I637261,I637278,I637295,I1284825,I637335,I637343,I637360,I637377,I637394,I637425,I1284831,I1284819,I637442,I637468,I637476,I637507,I637538,I637555,I637586,I637686,I975451,I637712,I637720,I637737,I975427,I975442,I637754,I975454,I637780,I637788,I975439,I975430,I637814,I637822,I637839,I637856,I637873,I637669,I637913,I637921,I637938,I637955,I637972,I637672,I638003,I975445,I975436,I638020,I975448,I638046,I638054,I637654,I638085,I637663,I638116,I638133,I637675,I638164,I975433,I637666,I637657,I637660,I637678,I638264,I1153758,I638290,I638298,I638315,I1153740,I1153752,I638332,I1153755,I638358,I638366,I1153749,I1153746,I638392,I638400,I638417,I638434,I638451,I1153764,I638491,I638499,I638516,I638533,I638550,I638581,I1153743,I638598,I638624,I638632,I638663,I638694,I638711,I638742,I1153761,I638842,I638868,I638876,I638893,I638910,I638936,I638944,I638970,I638978,I638995,I639012,I639029,I639069,I639077,I639094,I639111,I639128,I639159,I639176,I639202,I639210,I639241,I639272,I639289,I639320,I639420,I794885,I639446,I639454,I639471,I794873,I794891,I639488,I794888,I639514,I639522,I794879,I794876,I639548,I639556,I639573,I639590,I639607,I794870,I639647,I639655,I639672,I639689,I639706,I639737,I639754,I639780,I639788,I639819,I639850,I639867,I639898,I794882,I639998,I640024,I640032,I640049,I640066,I640092,I640100,I640126,I640134,I640151,I640168,I640185,I639981,I640225,I640233,I640250,I640267,I640284,I639984,I640315,I640332,I640358,I640366,I639966,I640397,I639975,I640428,I640445,I639987,I640476,I639978,I639969,I639972,I639990,I640576,I1326164,I640602,I640610,I640627,I1326149,I1326137,I640644,I1326152,I640670,I640678,I1326155,I640704,I640712,I640729,I640746,I640763,I640559,I1326143,I640803,I640811,I640828,I640845,I640862,I640562,I640893,I1326140,I1326146,I640910,I1326161,I640936,I640944,I640544,I640975,I640553,I641006,I641023,I640565,I641054,I1326158,I640556,I640547,I640550,I640568,I641154,I1018001,I641180,I641188,I641205,I1017998,I1018016,I641222,I1018013,I641248,I641256,I1017995,I641282,I641290,I641307,I641324,I641341,I1018007,I641381,I641389,I641406,I641423,I641440,I641471,I1018010,I641488,I641514,I641522,I641553,I641584,I641601,I641632,I1018004,I641732,I641758,I641766,I641783,I641800,I641826,I641834,I641860,I641868,I641885,I641902,I641919,I641715,I641959,I641967,I641984,I642001,I642018,I641718,I642049,I642066,I642092,I642100,I641700,I642131,I641709,I642162,I642179,I641721,I642210,I641712,I641703,I641706,I641724,I642310,I642336,I642344,I642361,I642378,I642404,I642412,I642438,I642446,I642463,I642480,I642497,I642537,I642545,I642562,I642579,I642596,I642627,I642644,I642670,I642678,I642709,I642740,I642757,I642788,I642888,I642914,I642922,I642939,I642956,I642982,I642990,I643016,I643024,I643041,I643058,I643075,I642871,I643115,I643123,I643140,I643157,I643174,I642874,I643205,I643222,I643248,I643256,I642856,I643287,I642865,I643318,I643335,I642877,I643366,I642868,I642859,I642862,I642880,I643466,I643492,I643500,I643517,I643534,I643560,I643568,I643594,I643602,I643619,I643636,I643653,I643693,I643701,I643718,I643735,I643752,I643783,I643800,I643826,I643834,I643865,I643896,I643913,I643944,I644044,I1251490,I644070,I644078,I644095,I1251493,I1251502,I644112,I1251505,I644138,I644146,I1251514,I1251496,I644172,I644180,I644197,I644214,I644231,I644027,I644271,I644279,I644296,I644313,I644330,I644030,I644361,I1251511,I644378,I1251508,I644404,I644412,I644012,I644443,I644021,I644474,I644491,I644033,I644522,I1251499,I644024,I644015,I644018,I644036,I644622,I644648,I644656,I644673,I644690,I644716,I644724,I644750,I644758,I644775,I644792,I644809,I644849,I644857,I644874,I644891,I644908,I644939,I644956,I644982,I644990,I645021,I645052,I645069,I645100,I645200,I1337469,I645226,I645234,I645251,I1337454,I1337442,I645268,I1337457,I645294,I645302,I1337460,I645328,I645336,I645353,I645370,I645387,I645183,I1337448,I645427,I645435,I645452,I645469,I645486,I645186,I645517,I1337445,I1337451,I645534,I1337466,I645560,I645568,I645168,I645599,I645177,I645630,I645647,I645189,I645678,I1337463,I645180,I645171,I645174,I645192,I645778,I1348774,I645804,I645812,I645829,I1348759,I1348747,I645846,I1348762,I645872,I645880,I1348765,I645906,I645914,I645931,I645948,I645965,I645761,I1348753,I646005,I646013,I646030,I646047,I646064,I645764,I646095,I1348750,I1348756,I646112,I1348771,I646138,I646146,I645746,I646177,I645755,I646208,I646225,I645767,I646256,I1348768,I645758,I645749,I645752,I645770,I646356,I1269204,I646382,I646390,I646407,I1269228,I1269210,I646424,I1269216,I646450,I646458,I1269222,I1269207,I646484,I646492,I646509,I646526,I646543,I646339,I1269219,I646583,I646591,I646608,I646625,I646642,I646342,I646673,I1269225,I1269213,I646690,I646716,I646724,I646324,I646755,I646333,I646786,I646803,I646345,I646834,I646336,I646327,I646330,I646348,I646934,I646960,I646968,I646985,I647002,I647028,I647036,I647062,I647070,I647087,I647104,I647121,I646917,I647161,I647169,I647186,I647203,I647220,I646920,I647251,I647268,I647294,I647302,I646902,I647333,I646911,I647364,I647381,I646923,I647412,I646914,I646905,I646908,I646926,I647512,I647538,I647546,I647563,I647580,I647606,I647614,I647640,I647648,I647665,I647682,I647699,I647739,I647747,I647764,I647781,I647798,I647829,I647846,I647872,I647880,I647911,I647942,I647959,I647990,I648090,I1367814,I648116,I648124,I648141,I1367799,I1367787,I648158,I1367802,I648184,I648192,I1367805,I648218,I648226,I648243,I648260,I648277,I1367793,I648317,I648325,I648342,I648359,I648376,I648407,I1367790,I1367796,I648424,I1367811,I648450,I648458,I648489,I648520,I648537,I648568,I1367808,I648668,I648694,I648702,I648719,I648736,I648762,I648770,I648796,I648804,I648821,I648838,I648855,I648895,I648903,I648920,I648937,I648954,I648985,I649002,I649028,I649036,I649067,I649098,I649115,I649146,I649246,I649272,I649280,I649297,I649314,I649340,I649348,I649374,I649382,I649399,I649416,I649433,I649473,I649481,I649498,I649515,I649532,I649563,I649580,I649606,I649614,I649645,I649676,I649693,I649724,I649824,I919895,I649850,I649858,I649875,I919871,I919886,I649892,I919898,I649918,I649926,I919883,I919874,I649952,I649960,I649977,I649994,I650011,I649807,I650051,I650059,I650076,I650093,I650110,I649810,I650141,I919889,I919880,I650158,I919892,I650184,I650192,I649792,I650223,I649801,I650254,I650271,I649813,I650302,I919877,I649804,I649795,I649798,I649816,I650402,I1079196,I650428,I650436,I650453,I1079178,I1079190,I650470,I1079193,I650496,I650504,I1079187,I1079184,I650530,I650538,I650555,I650572,I650589,I650385,I1079202,I650629,I650637,I650654,I650671,I650688,I650388,I650719,I1079181,I650736,I650762,I650770,I650370,I650801,I650379,I650832,I650849,I650391,I650880,I1079199,I650382,I650373,I650376,I650394,I650980,I651006,I651014,I651031,I651048,I651074,I651082,I651108,I651116,I651133,I651150,I651167,I651207,I651215,I651232,I651249,I651266,I651297,I651314,I651340,I651348,I651379,I651410,I651427,I651458,I651558,I651584,I651592,I651609,I651626,I651652,I651660,I651686,I651694,I651711,I651728,I651745,I651541,I651785,I651793,I651810,I651827,I651844,I651544,I651875,I651892,I651918,I651926,I651526,I651957,I651535,I651988,I652005,I651547,I652036,I651538,I651529,I651532,I651550,I652136,I652162,I652170,I652187,I652204,I652230,I652238,I652264,I652272,I652289,I652306,I652323,I652363,I652371,I652388,I652405,I652422,I652453,I652470,I652496,I652504,I652535,I652566,I652583,I652614,I652714,I652740,I652748,I652765,I652782,I652808,I652816,I652842,I652850,I652867,I652884,I652901,I652941,I652949,I652966,I652983,I653000,I653031,I653048,I653074,I653082,I653113,I653144,I653161,I653192,I653292,I653318,I653326,I653343,I653360,I653386,I653394,I653420,I653428,I653445,I653462,I653479,I653519,I653527,I653544,I653561,I653578,I653609,I653626,I653652,I653660,I653691,I653722,I653739,I653770,I653870,I833883,I653896,I653904,I653921,I833871,I833889,I653938,I833886,I653964,I653972,I833877,I833874,I653998,I654006,I654023,I654040,I654057,I653853,I833868,I654097,I654105,I654122,I654139,I654156,I653856,I654187,I654204,I654230,I654238,I653838,I654269,I653847,I654300,I654317,I653859,I654348,I833880,I653850,I653841,I653844,I653862,I654448,I654474,I654482,I654499,I654516,I654542,I654550,I654576,I654584,I654601,I654618,I654635,I654431,I654675,I654683,I654700,I654717,I654734,I654434,I654765,I654782,I654808,I654816,I654416,I654847,I654425,I654878,I654895,I654437,I654926,I654428,I654419,I654422,I654440,I655026,I655052,I655060,I655077,I655094,I655120,I655128,I655154,I655162,I655179,I655196,I655213,I655253,I655261,I655278,I655295,I655312,I655343,I655360,I655386,I655394,I655425,I655456,I655473,I655504,I655604,I655630,I655638,I655655,I655672,I655698,I655706,I655732,I655740,I655757,I655774,I655791,I655587,I655831,I655839,I655856,I655873,I655890,I655590,I655921,I655938,I655964,I655972,I655572,I656003,I655581,I656034,I656051,I655593,I656082,I655584,I655575,I655578,I655596,I656182,I1311289,I656208,I656216,I656233,I1311274,I1311262,I656250,I1311277,I656276,I656284,I1311280,I656310,I656318,I656335,I656352,I656369,I656165,I1311268,I656409,I656417,I656434,I656451,I656468,I656168,I656499,I1311265,I1311271,I656516,I1311286,I656542,I656550,I656150,I656581,I656159,I656612,I656629,I656171,I656660,I1311283,I656162,I656153,I656156,I656174,I656760,I656786,I656794,I656811,I656828,I656854,I656862,I656888,I656896,I656913,I656930,I656947,I656987,I656995,I657012,I657029,I657046,I657077,I657094,I657120,I657128,I657159,I657190,I657207,I657238,I657338,I657364,I657372,I657389,I657406,I657432,I657440,I657466,I657474,I657491,I657508,I657525,I657565,I657573,I657590,I657607,I657624,I657655,I657672,I657698,I657706,I657737,I657768,I657785,I657816,I657916,I931523,I657942,I657950,I657967,I931499,I931514,I657984,I931526,I658010,I658018,I931511,I931502,I658044,I658052,I658069,I658086,I658103,I657899,I658143,I658151,I658168,I658185,I658202,I657902,I658233,I931517,I931508,I658250,I931520,I658276,I658284,I657884,I658315,I657893,I658346,I658363,I657905,I658394,I931505,I657896,I657887,I657890,I657908,I658494,I856544,I658520,I658528,I658545,I856532,I856550,I658562,I856547,I658588,I658596,I856538,I856535,I658622,I658630,I658647,I658664,I658681,I658477,I856529,I658721,I658729,I658746,I658763,I658780,I658480,I658811,I658828,I658854,I658862,I658462,I658893,I658471,I658924,I658941,I658483,I658972,I856541,I658474,I658465,I658468,I658486,I659072,I659098,I659106,I659123,I659140,I659166,I659174,I659200,I659208,I659225,I659242,I659259,I659055,I659299,I659307,I659324,I659341,I659358,I659058,I659389,I659406,I659432,I659440,I659040,I659471,I659049,I659502,I659519,I659061,I659550,I659052,I659043,I659046,I659064,I659650,I659676,I659684,I659701,I659718,I659744,I659752,I659778,I659786,I659803,I659820,I659837,I659633,I659877,I659885,I659902,I659919,I659936,I659636,I659967,I659984,I660010,I660018,I659618,I660049,I659627,I660080,I660097,I659639,I660128,I659630,I659621,I659624,I659642,I660228,I994831,I660254,I660262,I660279,I994807,I994822,I660296,I994834,I660322,I660330,I994819,I994810,I660356,I660364,I660381,I660398,I660415,I660211,I660455,I660463,I660480,I660497,I660514,I660214,I660545,I994825,I994816,I660562,I994828,I660588,I660596,I660196,I660627,I660205,I660658,I660675,I660217,I660706,I994813,I660208,I660199,I660202,I660220,I660806,I660832,I660840,I660857,I660874,I660900,I660908,I660934,I660942,I660959,I660976,I660993,I661033,I661041,I661058,I661075,I661092,I661123,I661140,I661166,I661174,I661205,I661236,I661253,I661284,I661384,I661410,I661418,I661435,I661452,I661478,I661486,I661512,I661520,I661537,I661554,I661571,I661367,I661611,I661619,I661636,I661653,I661670,I661370,I661701,I661718,I661744,I661752,I661352,I661783,I661361,I661814,I661831,I661373,I661862,I661364,I661355,I661358,I661376,I661962,I834937,I661988,I661996,I662013,I834925,I834943,I662030,I834940,I662056,I662064,I834931,I834928,I662090,I662098,I662115,I662132,I662149,I661945,I834922,I662189,I662197,I662214,I662231,I662248,I661948,I662279,I662296,I662322,I662330,I661930,I662361,I661939,I662392,I662409,I661951,I662440,I834934,I661942,I661933,I661936,I661954,I662540,I1173410,I662566,I662574,I662591,I1173392,I1173404,I662608,I1173407,I662634,I662642,I1173401,I1173398,I662668,I662676,I662693,I662710,I662727,I662523,I1173416,I662767,I662775,I662792,I662809,I662826,I662526,I662857,I1173395,I662874,I662900,I662908,I662508,I662939,I662517,I662970,I662987,I662529,I663018,I1173413,I662520,I662511,I662514,I662532,I663118,I790669,I663144,I663152,I663169,I790657,I790675,I663186,I790672,I663212,I663220,I790663,I790660,I663246,I663254,I663271,I663288,I663305,I790654,I663345,I663353,I663370,I663387,I663404,I663435,I663452,I663478,I663486,I663517,I663548,I663565,I663596,I790666,I663696,I1242242,I663722,I663730,I663747,I1242245,I1242254,I663764,I1242257,I663790,I663798,I1242266,I1242248,I663824,I663832,I663849,I663866,I663883,I663923,I663931,I663948,I663965,I663982,I664013,I1242263,I664030,I1242260,I664056,I664064,I664095,I664126,I664143,I664174,I1242251,I664274,I1202888,I664300,I664308,I664325,I1202870,I1202882,I664342,I1202885,I664368,I664376,I1202879,I1202876,I664402,I664410,I664427,I664444,I664461,I1202894,I664501,I664509,I664526,I664543,I664560,I664591,I1202873,I664608,I664634,I664642,I664673,I664704,I664721,I664752,I1202891,I664852,I664878,I664886,I664903,I664920,I664946,I664954,I664980,I664988,I665005,I665022,I665039,I664835,I665079,I665087,I665104,I665121,I665138,I664838,I665169,I665186,I665212,I665220,I664820,I665251,I664829,I665282,I665299,I664841,I665330,I664832,I664823,I664826,I664844,I665430,I1053905,I665456,I665464,I665481,I1053902,I1053920,I665498,I1053917,I665524,I665532,I1053899,I665558,I665566,I665583,I665600,I665617,I1053911,I665657,I665665,I665682,I665699,I665716,I665747,I1053914,I665764,I665790,I665798,I665829,I665860,I665877,I665908,I1053908,I666008,I1289434,I666034,I666042,I666059,I1289458,I1289440,I666076,I1289446,I666102,I666110,I1289452,I1289437,I666136,I666144,I666161,I666178,I666195,I665991,I1289449,I666235,I666243,I666260,I666277,I666294,I665994,I666325,I1289455,I1289443,I666342,I666368,I666376,I665976,I666407,I665985,I666438,I666455,I665997,I666486,I665988,I665979,I665982,I666000,I666586,I666612,I666620,I666637,I666654,I666680,I666688,I666714,I666722,I666739,I666756,I666773,I666569,I666813,I666821,I666838,I666855,I666872,I666572,I666903,I666920,I666946,I666954,I666554,I666985,I666563,I667016,I667033,I666575,I667064,I666566,I666557,I666560,I666578,I667164,I667190,I667198,I667215,I667232,I667258,I667266,I667292,I667300,I667317,I667334,I667351,I667391,I667399,I667416,I667433,I667450,I667481,I667498,I667524,I667532,I667563,I667594,I667611,I667642,I667742,I1162428,I667768,I667776,I667793,I1162410,I1162422,I667810,I1162425,I667836,I667844,I1162419,I1162416,I667870,I667878,I667895,I667912,I667929,I667725,I1162434,I667969,I667977,I667994,I668011,I668028,I667728,I668059,I1162413,I668076,I668102,I668110,I667710,I668141,I667719,I668172,I668189,I667731,I668220,I1162431,I667722,I667713,I667716,I667734,I668320,I929585,I668346,I668354,I668371,I929561,I929576,I668388,I929588,I668414,I668422,I929573,I929564,I668448,I668456,I668473,I668490,I668507,I668303,I668547,I668555,I668572,I668589,I668606,I668306,I668637,I929579,I929570,I668654,I929582,I668680,I668688,I668288,I668719,I668297,I668750,I668767,I668309,I668798,I929567,I668300,I668291,I668294,I668312,I668898,I668924,I668932,I668949,I668966,I668992,I669000,I669026,I669034,I669051,I669068,I669085,I669125,I669133,I669150,I669167,I669184,I669215,I669232,I669258,I669266,I669297,I669328,I669345,I669376,I669476,I824924,I669502,I669510,I669527,I824912,I824930,I669544,I824927,I669570,I669578,I824918,I824915,I669604,I669612,I669629,I669646,I669663,I824909,I669703,I669711,I669728,I669745,I669762,I669793,I669810,I669836,I669844,I669875,I669906,I669923,I669954,I824921,I670054,I670080,I670088,I670105,I670122,I670148,I670156,I670182,I670190,I670207,I670224,I670241,I670037,I670281,I670289,I670306,I670323,I670340,I670040,I670371,I670388,I670414,I670422,I670022,I670453,I670031,I670484,I670501,I670043,I670532,I670034,I670025,I670028,I670046,I670632,I670658,I670666,I670683,I670700,I670726,I670734,I670760,I670768,I670785,I670802,I670819,I670859,I670867,I670884,I670901,I670918,I670949,I670966,I670992,I671000,I671031,I671062,I671079,I671110,I671210,I1150868,I671236,I671244,I671261,I1150850,I1150862,I671278,I1150865,I671304,I671312,I1150859,I1150856,I671338,I671346,I671363,I671380,I671397,I1150874,I671437,I671445,I671462,I671479,I671496,I671527,I1150853,I671544,I671570,I671578,I671609,I671640,I671657,I671688,I1150871,I671788,I949611,I671814,I671822,I671839,I949587,I949602,I671856,I949614,I671882,I671890,I949599,I949590,I671916,I671924,I671941,I671958,I671975,I672015,I672023,I672040,I672057,I672074,I672105,I949605,I949596,I672122,I949608,I672148,I672156,I672187,I672218,I672235,I672266,I949593,I672366,I944443,I672392,I672400,I672417,I944419,I944434,I672434,I944446,I672460,I672468,I944431,I944422,I672494,I672502,I672519,I672536,I672553,I672593,I672601,I672618,I672635,I672652,I672683,I944437,I944428,I672700,I944440,I672726,I672734,I672765,I672796,I672813,I672844,I944425,I672944,I672970,I672978,I672995,I673012,I673038,I673046,I673072,I673080,I673097,I673114,I673131,I672927,I673171,I673179,I673196,I673213,I673230,I672930,I673261,I673278,I673304,I673312,I672912,I673343,I672921,I673374,I673391,I672933,I673422,I672924,I672915,I672918,I672936,I673522,I1000645,I673548,I673556,I673573,I1000621,I1000636,I673590,I1000648,I673616,I673624,I1000633,I1000624,I673650,I673658,I673675,I673692,I673709,I673505,I673749,I673757,I673774,I673791,I673808,I673508,I673839,I1000639,I1000630,I673856,I1000642,I673882,I673890,I673490,I673921,I673499,I673952,I673969,I673511,I674000,I1000627,I673502,I673493,I673496,I673514,I674100,I1314264,I674126,I674134,I674151,I1314249,I1314237,I674168,I1314252,I674194,I674202,I1314255,I674228,I674236,I674253,I674270,I674287,I1314243,I674327,I674335,I674352,I674369,I674386,I674417,I1314240,I1314246,I674434,I1314261,I674460,I674468,I674499,I674530,I674547,I674578,I1314258,I674678,I674704,I674712,I674729,I674746,I674772,I674780,I674806,I674814,I674831,I674848,I674865,I674905,I674913,I674930,I674947,I674964,I674995,I675012,I675038,I675046,I675077,I675108,I675125,I675156,I675256,I1135262,I675282,I675290,I675307,I1135244,I1135256,I675324,I1135259,I675350,I675358,I1135253,I1135250,I675384,I675392,I675409,I675426,I675443,I675239,I1135268,I675483,I675491,I675508,I675525,I675542,I675242,I675573,I1135247,I675590,I675616,I675624,I675224,I675655,I675233,I675686,I675703,I675245,I675734,I1135265,I675236,I675227,I675230,I675248,I675834,I981265,I675860,I675868,I675885,I981241,I981256,I675902,I981268,I675928,I675936,I981253,I981244,I675962,I675970,I675987,I676004,I676021,I675817,I676061,I676069,I676086,I676103,I676120,I675820,I676151,I981259,I981250,I676168,I981262,I676194,I676202,I675802,I676233,I675811,I676264,I676281,I675823,I676312,I981247,I675814,I675805,I675808,I675826,I676412,I676438,I676446,I676463,I676480,I676506,I676514,I676540,I676548,I676565,I676582,I676599,I676395,I676639,I676647,I676664,I676681,I676698,I676398,I676729,I676746,I676772,I676780,I676380,I676811,I676389,I676842,I676859,I676401,I676890,I676392,I676383,I676386,I676404,I676990,I1335089,I677016,I677024,I677041,I1335074,I1335062,I677058,I1335077,I677084,I677092,I1335080,I677118,I677126,I677143,I677160,I677177,I1335068,I677217,I677225,I677242,I677259,I677276,I677307,I1335065,I1335071,I677324,I1335086,I677350,I677358,I677389,I677420,I677437,I677468,I1335083,I677568,I853382,I677594,I677602,I677619,I853370,I853388,I677636,I853385,I677662,I677670,I853376,I853373,I677696,I677704,I677721,I677738,I677755,I677551,I853367,I677795,I677803,I677820,I677837,I677854,I677554,I677885,I677902,I677928,I677936,I677536,I677967,I677545,I677998,I678015,I677557,I678046,I853379,I677548,I677539,I677542,I677560,I678146,I1182080,I678172,I678180,I678197,I1182062,I1182074,I678214,I1182077,I678240,I678248,I1182071,I1182068,I678274,I678282,I678299,I678316,I678333,I678129,I1182086,I678373,I678381,I678398,I678415,I678432,I678132,I678463,I1182065,I678480,I678506,I678514,I678114,I678545,I678123,I678576,I678593,I678135,I678624,I1182083,I678126,I678117,I678120,I678138,I678724,I1153180,I678750,I678758,I678775,I1153162,I1153174,I678792,I1153177,I678818,I678826,I1153171,I1153168,I678852,I678860,I678877,I678894,I678911,I1153186,I678951,I678959,I678976,I678993,I679010,I679041,I1153165,I679058,I679084,I679092,I679123,I679154,I679171,I679202,I1153183,I679302,I679328,I679336,I679353,I679370,I679396,I679404,I679430,I679438,I679455,I679472,I679489,I679285,I679529,I679537,I679554,I679571,I679588,I679288,I679619,I679636,I679662,I679670,I679270,I679701,I679279,I679732,I679749,I679291,I679780,I679282,I679273,I679276,I679294,I679880,I679906,I679914,I679931,I679948,I679974,I679982,I680008,I680016,I680033,I680050,I680067,I680107,I680115,I680132,I680149,I680166,I680197,I680214,I680240,I680248,I680279,I680310,I680327,I680358,I680458,I680484,I680492,I680509,I680526,I680552,I680560,I680586,I680594,I680611,I680628,I680645,I680441,I680685,I680693,I680710,I680727,I680744,I680444,I680775,I680792,I680818,I680826,I680426,I680857,I680435,I680888,I680905,I680447,I680936,I680438,I680429,I680432,I680450,I681036,I681062,I681070,I681087,I681104,I681130,I681138,I681164,I681172,I681189,I681206,I681223,I681019,I681263,I681271,I681288,I681305,I681322,I681022,I681353,I681370,I681396,I681404,I681004,I681435,I681013,I681466,I681483,I681025,I681514,I681016,I681007,I681010,I681028,I681614,I681640,I681648,I681665,I681682,I681708,I681716,I681742,I681750,I681767,I681784,I681801,I681597,I681841,I681849,I681866,I681883,I681900,I681600,I681931,I681948,I681974,I681982,I681582,I682013,I681591,I682044,I682061,I681603,I682092,I681594,I681585,I681588,I681606,I682192,I682218,I682226,I682243,I682260,I682286,I682294,I682320,I682328,I682345,I682362,I682379,I682419,I682427,I682444,I682461,I682478,I682509,I682526,I682552,I682560,I682591,I682622,I682639,I682670,I682770,I1268048,I682796,I682804,I682821,I1268072,I1268054,I682838,I1268060,I682864,I682872,I1268066,I1268051,I682898,I682906,I682923,I682940,I682957,I1268063,I682997,I683005,I683022,I683039,I683056,I683087,I1268069,I1268057,I683104,I683130,I683138,I683169,I683200,I683217,I683248,I683348,I683374,I683382,I683399,I683416,I683442,I683450,I683476,I683484,I683501,I683518,I683535,I683575,I683583,I683600,I683617,I683634,I683665,I683682,I683708,I683716,I683747,I683778,I683795,I683826,I683926,I1095380,I683952,I683960,I683977,I1095362,I1095374,I683994,I1095377,I684020,I684028,I1095371,I1095368,I684054,I684062,I684079,I684096,I684113,I1095386,I684153,I684161,I684178,I684195,I684212,I684243,I1095365,I684260,I684286,I684294,I684325,I684356,I684373,I684404,I1095383,I684504,I684530,I684538,I684555,I684572,I684598,I684606,I684632,I684640,I684657,I684674,I684691,I684487,I684731,I684739,I684756,I684773,I684790,I684490,I684821,I684838,I684864,I684872,I684472,I684903,I684481,I684934,I684951,I684493,I684982,I684484,I684475,I684478,I684496,I685082,I958655,I685108,I685116,I685133,I958631,I958646,I685150,I958658,I685176,I685184,I958643,I958634,I685210,I685218,I685235,I685252,I685269,I685309,I685317,I685334,I685351,I685368,I685399,I958649,I958640,I685416,I958652,I685442,I685450,I685481,I685512,I685529,I685560,I958637,I685660,I685686,I685694,I685711,I685728,I685754,I685762,I685788,I685796,I685813,I685830,I685847,I685887,I685895,I685912,I685929,I685946,I685977,I685994,I686020,I686028,I686059,I686090,I686107,I686138,I686238,I1212866,I686264,I686272,I686289,I1212869,I1212878,I686306,I1212881,I686332,I686340,I1212890,I1212872,I686366,I686374,I686391,I686408,I686425,I686465,I686473,I686490,I686507,I686524,I686555,I1212887,I686572,I1212884,I686598,I686606,I686637,I686668,I686685,I686716,I1212875,I686816,I686842,I686850,I686867,I686884,I686910,I686918,I686944,I686952,I686969,I686986,I687003,I687043,I687051,I687068,I687085,I687102,I687133,I687150,I687176,I687184,I687215,I687246,I687263,I687294,I687394,I687420,I687428,I687445,I687462,I687488,I687496,I687522,I687530,I687547,I687564,I687581,I687621,I687629,I687646,I687663,I687680,I687711,I687728,I687754,I687762,I687793,I687824,I687841,I687872,I687972,I687998,I688006,I688023,I688040,I688066,I688074,I688100,I688108,I688125,I688142,I688159,I688199,I688207,I688224,I688241,I688258,I688289,I688306,I688332,I688340,I688371,I688402,I688419,I688450,I688550,I688576,I688584,I688601,I688618,I688644,I688652,I688678,I688686,I688703,I688720,I688737,I688533,I688777,I688785,I688802,I688819,I688836,I688536,I688867,I688884,I688910,I688918,I688518,I688949,I688527,I688980,I688997,I688539,I689028,I688530,I688521,I688524,I688542,I689128,I689154,I689162,I689179,I689196,I689222,I689230,I689256,I689264,I689281,I689298,I689315,I689355,I689363,I689380,I689397,I689414,I689445,I689462,I689488,I689496,I689527,I689558,I689575,I689606,I689706,I1226466,I689732,I689740,I689757,I1226469,I1226478,I689774,I1226481,I689800,I689808,I1226490,I1226472,I689834,I689842,I689859,I689876,I689893,I689933,I689941,I689958,I689975,I689992,I690023,I1226487,I690040,I1226484,I690066,I690074,I690105,I690136,I690153,I690184,I1226475,I690284,I1035953,I690310,I690318,I690335,I1035950,I1035968,I690352,I1035965,I690378,I690386,I1035947,I690412,I690420,I690437,I690454,I690471,I690267,I1035959,I690511,I690519,I690536,I690553,I690570,I690270,I690601,I1035962,I690618,I690644,I690652,I690252,I690683,I690261,I690714,I690731,I690273,I690762,I1035956,I690264,I690255,I690258,I690276,I690862,I941859,I690888,I690896,I690913,I941835,I941850,I690930,I941862,I690956,I690964,I941847,I941838,I690990,I690998,I691015,I691032,I691049,I690845,I691089,I691097,I691114,I691131,I691148,I690848,I691179,I941853,I941844,I691196,I941856,I691222,I691230,I690830,I691261,I690839,I691292,I691309,I690851,I691340,I941841,I690842,I690833,I690836,I690854,I691440,I691466,I691474,I691491,I691508,I691534,I691542,I691568,I691576,I691593,I691610,I691627,I691667,I691675,I691692,I691709,I691726,I691757,I691774,I691800,I691808,I691839,I691870,I691887,I691918,I692018,I692044,I692052,I692069,I692086,I692112,I692120,I692146,I692154,I692171,I692188,I692205,I692001,I692245,I692253,I692270,I692287,I692304,I692004,I692335,I692352,I692378,I692386,I691986,I692417,I691995,I692448,I692465,I692007,I692496,I691998,I691989,I691992,I692010,I692596,I1332114,I692622,I692630,I692647,I1332099,I1332087,I692664,I1332102,I692690,I692698,I1332105,I692724,I692732,I692749,I692766,I692783,I692579,I1332093,I692823,I692831,I692848,I692865,I692882,I692582,I692913,I1332090,I1332096,I692930,I1332111,I692956,I692964,I692564,I692995,I692573,I693026,I693043,I692585,I693074,I1332108,I692576,I692567,I692570,I692588,I693174,I1058393,I693200,I693208,I693225,I1058390,I1058408,I693242,I1058405,I693268,I693276,I1058387,I693302,I693310,I693327,I693344,I693361,I693157,I1058399,I693401,I693409,I693426,I693443,I693460,I693160,I693491,I1058402,I693508,I693534,I693542,I693142,I693573,I693151,I693604,I693621,I693163,I693652,I1058396,I693154,I693145,I693148,I693166,I693752,I693778,I693786,I693803,I693820,I693846,I693854,I693880,I693888,I693905,I693922,I693939,I693735,I693979,I693987,I694004,I694021,I694038,I693738,I694069,I694086,I694112,I694120,I693720,I694151,I693729,I694182,I694199,I693741,I694230,I693732,I693723,I693726,I693744,I694330,I826505,I694356,I694364,I694381,I826493,I826511,I694398,I826508,I694424,I694432,I826499,I826496,I694458,I694466,I694483,I694500,I694517,I694313,I826490,I694557,I694565,I694582,I694599,I694616,I694316,I694647,I694664,I694690,I694698,I694298,I694729,I694307,I694760,I694777,I694319,I694808,I826502,I694310,I694301,I694304,I694322,I694908,I694934,I694942,I694959,I694976,I695002,I695010,I695036,I695044,I695061,I695078,I695095,I695135,I695143,I695160,I695177,I695194,I695225,I695242,I695268,I695276,I695307,I695338,I695355,I695386,I695486,I936691,I695512,I695520,I695537,I936667,I936682,I695554,I936694,I695580,I695588,I936679,I936670,I695614,I695622,I695639,I695656,I695673,I695469,I695713,I695721,I695738,I695755,I695772,I695472,I695803,I936685,I936676,I695820,I936688,I695846,I695854,I695454,I695885,I695463,I695916,I695933,I695475,I695964,I936673,I695466,I695457,I695460,I695478,I696064,I1197108,I696090,I696098,I696115,I1197090,I1197102,I696132,I1197105,I696158,I696166,I1197099,I1197096,I696192,I696200,I696217,I696234,I696251,I1197114,I696291,I696299,I696316,I696333,I696350,I696381,I1197093,I696398,I696424,I696432,I696463,I696494,I696511,I696542,I1197111,I696642,I1105784,I696668,I696676,I696693,I1105766,I1105778,I696710,I1105781,I696736,I696744,I1105775,I1105772,I696770,I696778,I696795,I696812,I696829,I1105790,I696869,I696877,I696894,I696911,I696928,I696959,I1105769,I696976,I697002,I697010,I697041,I697072,I697089,I697120,I1105787,I697220,I697246,I697254,I697271,I697288,I697314,I697322,I697348,I697356,I697373,I697390,I697407,I697447,I697455,I697472,I697489,I697506,I697537,I697554,I697580,I697588,I697619,I697650,I697667,I697698,I697798,I1207426,I697824,I697832,I697849,I1207429,I1207438,I697866,I1207441,I697892,I697900,I1207450,I1207432,I697926,I697934,I697951,I697968,I697985,I697781,I698025,I698033,I698050,I698067,I698084,I697784,I698115,I1207447,I698132,I1207444,I698158,I698166,I697766,I698197,I697775,I698228,I698245,I697787,I698276,I1207435,I697778,I697769,I697772,I697790,I698376,I1041002,I698402,I698410,I698427,I1040999,I1041017,I698444,I1041014,I698470,I698478,I1040996,I698504,I698512,I698529,I698546,I698563,I1041008,I698603,I698611,I698628,I698645,I698662,I698693,I1041011,I698710,I698736,I698744,I698775,I698806,I698823,I698854,I1041005,I698954,I698980,I698988,I699005,I699022,I699048,I699056,I699082,I699090,I699107,I699124,I699141,I698937,I699181,I699189,I699206,I699223,I699240,I698940,I699271,I699288,I699314,I699322,I698922,I699353,I698931,I699384,I699401,I698943,I699432,I698934,I698925,I698928,I698946,I699532,I999353,I699558,I699566,I699583,I999329,I999344,I699600,I999356,I699626,I699634,I999341,I999332,I699660,I699668,I699685,I699702,I699719,I699515,I699759,I699767,I699784,I699801,I699818,I699518,I699849,I999347,I999338,I699866,I999350,I699892,I699900,I699500,I699931,I699509,I699962,I699979,I699521,I700010,I999335,I699512,I699503,I699506,I699524,I700110,I700136,I700144,I700161,I700178,I700204,I700212,I700238,I700246,I700263,I700280,I700297,I700093,I700337,I700345,I700362,I700379,I700396,I700096,I700427,I700444,I700470,I700478,I700078,I700509,I700087,I700540,I700557,I700099,I700588,I700090,I700081,I700084,I700102,I700688,I700714,I700722,I700739,I700756,I700782,I700790,I700816,I700824,I700841,I700858,I700875,I700671,I700915,I700923,I700940,I700957,I700974,I700674,I701005,I701022,I701048,I701056,I700656,I701087,I700665,I701118,I701135,I700677,I701166,I700668,I700659,I700662,I700680,I701266,I1358889,I701292,I701300,I701317,I1358874,I1358862,I701334,I1358877,I701360,I701368,I1358880,I701394,I701402,I701419,I701436,I701453,I701249,I1358868,I701493,I701501,I701518,I701535,I701552,I701252,I701583,I1358865,I1358871,I701600,I1358886,I701626,I701634,I701234,I701665,I701243,I701696,I701713,I701255,I701744,I1358883,I701246,I701237,I701240,I701258,I701844,I701870,I701878,I701895,I701912,I701938,I701946,I701972,I701980,I701997,I702014,I702031,I701827,I702071,I702079,I702096,I702113,I702130,I701830,I702161,I702178,I702204,I702212,I701812,I702243,I701821,I702274,I702291,I701833,I702322,I701824,I701815,I701818,I701836,I702422,I781183,I702448,I702456,I702473,I781171,I781189,I702490,I781186,I702516,I702524,I781177,I781174,I702550,I702558,I702575,I702592,I702609,I702405,I781168,I702649,I702657,I702674,I702691,I702708,I702408,I702739,I702756,I702782,I702790,I702390,I702821,I702399,I702852,I702869,I702411,I702900,I781180,I702402,I702393,I702396,I702414,I703000,I703026,I703034,I703051,I703068,I703094,I703102,I703128,I703136,I703153,I703170,I703187,I702983,I703227,I703235,I703252,I703269,I703286,I702986,I703317,I703334,I703360,I703368,I702968,I703399,I702977,I703430,I703447,I702989,I703478,I702980,I702971,I702974,I702992,I703578,I786980,I703604,I703612,I703629,I786968,I786986,I703646,I786983,I703672,I703680,I786974,I786971,I703706,I703714,I703731,I703748,I703765,I703561,I786965,I703805,I703813,I703830,I703847,I703864,I703564,I703895,I703912,I703938,I703946,I703546,I703977,I703555,I704008,I704025,I703567,I704056,I786977,I703558,I703549,I703552,I703570,I704156,I704182,I704190,I704207,I704224,I704250,I704258,I704284,I704292,I704309,I704326,I704343,I704139,I704383,I704391,I704408,I704425,I704442,I704142,I704473,I704490,I704516,I704524,I704124,I704555,I704133,I704586,I704603,I704145,I704634,I704136,I704127,I704130,I704148,I704734,I704760,I704768,I704785,I704802,I704828,I704836,I704862,I704870,I704887,I704904,I704921,I704961,I704969,I704986,I705003,I705020,I705051,I705068,I705094,I705102,I705133,I705164,I705181,I705212,I705312,I1320809,I705338,I705346,I705363,I1320794,I1320782,I705380,I1320797,I705406,I705414,I1320800,I705440,I705448,I705465,I705482,I705499,I1320788,I705539,I705547,I705564,I705581,I705598,I705629,I1320785,I1320791,I705646,I1320806,I705672,I705680,I705711,I705742,I705759,I705790,I1320803,I705890,I705916,I705924,I705941,I705958,I705984,I705992,I706018,I706026,I706043,I706060,I706077,I706117,I706125,I706142,I706159,I706176,I706207,I706224,I706250,I706258,I706289,I706320,I706337,I706368,I706468,I706494,I706502,I706519,I706536,I706562,I706570,I706596,I706604,I706621,I706638,I706655,I706695,I706703,I706720,I706737,I706754,I706785,I706802,I706828,I706836,I706867,I706898,I706915,I706946,I707046,I1188438,I707072,I707080,I707097,I1188420,I1188432,I707114,I1188435,I707140,I707148,I1188429,I1188426,I707174,I707182,I707199,I707216,I707233,I1188444,I707273,I707281,I707298,I707315,I707332,I707363,I1188423,I707380,I707406,I707414,I707445,I707476,I707493,I707524,I1188441,I707624,I707650,I707658,I707675,I707692,I707718,I707726,I707752,I707760,I707777,I707794,I707811,I707607,I707851,I707859,I707876,I707893,I707910,I707610,I707941,I707958,I707984,I707992,I707592,I708023,I707601,I708054,I708071,I707613,I708102,I707604,I707595,I707598,I707616,I708202,I1056710,I708228,I708236,I708253,I1056707,I1056725,I708270,I1056722,I708296,I708304,I1056704,I708330,I708338,I708355,I708372,I708389,I708185,I1056716,I708429,I708437,I708454,I708471,I708488,I708188,I708519,I1056719,I708536,I708562,I708570,I708170,I708601,I708179,I708632,I708649,I708191,I708680,I1056713,I708182,I708173,I708176,I708194,I708780,I779602,I708806,I708814,I708831,I779590,I779608,I708848,I779605,I708874,I708882,I779596,I779593,I708908,I708916,I708933,I708950,I708967,I708763,I779587,I709007,I709015,I709032,I709049,I709066,I708766,I709097,I709114,I709140,I709148,I708748,I709179,I708757,I709210,I709227,I708769,I709258,I779599,I708760,I708751,I708754,I708772,I709358,I1057832,I709384,I709392,I709409,I1057829,I1057847,I709426,I1057844,I709452,I709460,I1057826,I709486,I709494,I709511,I709528,I709545,I709341,I1057838,I709585,I709593,I709610,I709627,I709644,I709344,I709675,I1057841,I709692,I709718,I709726,I709326,I709757,I709335,I709788,I709805,I709347,I709836,I1057835,I709338,I709329,I709332,I709350,I709936,I807533,I709962,I709970,I709987,I807521,I807539,I710004,I807536,I710030,I710038,I807527,I807524,I710064,I710072,I710089,I710106,I710123,I709919,I807518,I710163,I710171,I710188,I710205,I710222,I709922,I710253,I710270,I710296,I710304,I709904,I710335,I709913,I710366,I710383,I709925,I710414,I807530,I709916,I709907,I709910,I709928,I710514,I964469,I710540,I710548,I710565,I964445,I964460,I710582,I964472,I710608,I710616,I964457,I964448,I710642,I710650,I710667,I710684,I710701,I710741,I710749,I710766,I710783,I710800,I710831,I964463,I964454,I710848,I964466,I710874,I710882,I710913,I710944,I710961,I710992,I964451,I711092,I711118,I711126,I711143,I711160,I711186,I711194,I711220,I711228,I711245,I711262,I711279,I711319,I711327,I711344,I711361,I711378,I711409,I711426,I711452,I711460,I711491,I711522,I711539,I711570,I711670,I711696,I711704,I711721,I711738,I711764,I711772,I711798,I711806,I711823,I711840,I711857,I711653,I711897,I711905,I711922,I711939,I711956,I711656,I711987,I712004,I712030,I712038,I711638,I712069,I711647,I712100,I712117,I711659,I712148,I711650,I711641,I711644,I711662,I712248,I1368409,I712274,I712282,I712299,I1368394,I1368382,I712316,I1368397,I712342,I712350,I1368400,I712376,I712384,I712401,I712418,I712435,I1368388,I712475,I712483,I712500,I712517,I712534,I712565,I1368385,I1368391,I712582,I1368406,I712608,I712616,I712647,I712678,I712695,I712726,I1368403,I712826,I712852,I712860,I712877,I712894,I712920,I712928,I712954,I712962,I712979,I712996,I713013,I712809,I713053,I713061,I713078,I713095,I713112,I712812,I713143,I713160,I713186,I713194,I712794,I713225,I712803,I713256,I713273,I712815,I713304,I712806,I712797,I712800,I712818,I713404,I1304239,I713430,I713438,I713455,I1304227,I1304245,I713472,I1304236,I713498,I713506,I1304251,I1304248,I713532,I713540,I713557,I713574,I713591,I1304230,I713631,I713639,I713656,I713673,I713690,I713721,I1304224,I713738,I1304233,I713764,I713772,I713803,I713834,I713851,I713882,I1304242,I713982,I831248,I714008,I714016,I714033,I831236,I831254,I714050,I831251,I714076,I714084,I831242,I831239,I714110,I714118,I714135,I714152,I714169,I831233,I714209,I714217,I714234,I714251,I714268,I714299,I714316,I714342,I714350,I714381,I714412,I714429,I714460,I831245,I714560,I1010147,I714586,I714594,I714611,I1010144,I1010162,I714628,I1010159,I714654,I714662,I1010141,I714688,I714696,I714713,I714730,I714747,I1010153,I714787,I714795,I714812,I714829,I714846,I714877,I1010156,I714894,I714920,I714928,I714959,I714990,I715007,I715038,I1010150,I715138,I1245506,I715164,I715172,I715189,I1245509,I1245518,I715206,I1245521,I715232,I715240,I1245530,I1245512,I715266,I715274,I715291,I715308,I715325,I715365,I715373,I715390,I715407,I715424,I715455,I1245527,I715472,I1245524,I715498,I715506,I715537,I715568,I715585,I715616,I1245515,I715716,I1029782,I715742,I715750,I715767,I1029779,I1029797,I715784,I1029794,I715810,I715818,I1029776,I715844,I715852,I715869,I715886,I715903,I1029788,I715943,I715951,I715968,I715985,I716002,I716033,I1029791,I716050,I716076,I716084,I716115,I716146,I716163,I716194,I1029785,I716294,I1071682,I716320,I716328,I716345,I1071664,I1071676,I716362,I1071679,I716388,I716396,I1071673,I1071670,I716422,I716430,I716447,I716464,I716481,I1071688,I716521,I716529,I716546,I716563,I716580,I716611,I1071667,I716628,I716654,I716662,I716693,I716724,I716741,I716772,I1071685,I716872,I1372574,I716898,I716906,I716923,I1372559,I1372547,I716940,I1372562,I716966,I716974,I1372565,I717000,I717008,I717025,I717042,I717059,I716855,I1372553,I717099,I717107,I717124,I717141,I717158,I716858,I717189,I1372550,I1372556,I717206,I1372571,I717232,I717240,I716840,I717271,I716849,I717302,I717319,I716861,I717350,I1372568,I716852,I716843,I716846,I716864,I717450,I717476,I717484,I717501,I717518,I717544,I717552,I717578,I717586,I717603,I717620,I717637,I717433,I717677,I717685,I717702,I717719,I717736,I717436,I717767,I717784,I717810,I717818,I717418,I717849,I717427,I717880,I717897,I717439,I717928,I717430,I717421,I717424,I717442,I718028,I985787,I718054,I718062,I718079,I985763,I985778,I718096,I985790,I718122,I718130,I985775,I985766,I718156,I718164,I718181,I718198,I718215,I718255,I718263,I718280,I718297,I718314,I718345,I985781,I985772,I718362,I985784,I718388,I718396,I718427,I718458,I718475,I718506,I985769,I718606,I718632,I718640,I718657,I718674,I718700,I718708,I718734,I718742,I718759,I718776,I718793,I718589,I718833,I718841,I718858,I718875,I718892,I718592,I718923,I718940,I718966,I718974,I718574,I719005,I718583,I719036,I719053,I718595,I719084,I718586,I718577,I718580,I718598,I719184,I719210,I719218,I719235,I719252,I719278,I719286,I719312,I719320,I719337,I719354,I719371,I719167,I719411,I719419,I719436,I719453,I719470,I719170,I719501,I719518,I719544,I719552,I719152,I719583,I719161,I719614,I719631,I719173,I719662,I719164,I719155,I719158,I719176,I719762,I719788,I719796,I719813,I719830,I719856,I719864,I719890,I719898,I719915,I719932,I719949,I719745,I719989,I719997,I720014,I720031,I720048,I719748,I720079,I720096,I720122,I720130,I719730,I720161,I719739,I720192,I720209,I719751,I720240,I719742,I719733,I719736,I719754,I720340,I720366,I720374,I720391,I720408,I720434,I720442,I720468,I720476,I720493,I720510,I720527,I720567,I720575,I720592,I720609,I720626,I720657,I720674,I720700,I720708,I720739,I720770,I720787,I720818,I720918,I720944,I720952,I720969,I720986,I721012,I721020,I721046,I721054,I721071,I721088,I721105,I720901,I721145,I721153,I721170,I721187,I721204,I720904,I721235,I721252,I721278,I721286,I720886,I721317,I720895,I721348,I721365,I720907,I721396,I720898,I720889,I720892,I720910,I721496,I1265736,I721522,I721530,I721547,I1265760,I1265742,I721564,I1265748,I721590,I721598,I1265754,I1265739,I721624,I721632,I721649,I721666,I721683,I721479,I1265751,I721723,I721731,I721748,I721765,I721782,I721482,I721813,I1265757,I1265745,I721830,I721856,I721864,I721464,I721895,I721473,I721926,I721943,I721485,I721974,I721476,I721467,I721470,I721488,I722074,I722100,I722108,I722125,I722142,I722168,I722176,I722202,I722210,I722227,I722244,I722261,I722301,I722309,I722326,I722343,I722360,I722391,I722408,I722434,I722442,I722473,I722504,I722521,I722552,I722652,I722678,I722686,I722703,I722720,I722746,I722754,I722780,I722788,I722805,I722822,I722839,I722635,I722879,I722887,I722904,I722921,I722938,I722638,I722969,I722986,I723012,I723020,I722620,I723051,I722629,I723082,I723099,I722641,I723130,I722632,I722623,I722626,I722644,I723230,I1092490,I723256,I723264,I723281,I1092472,I1092484,I723298,I1092487,I723324,I723332,I1092481,I1092478,I723358,I723366,I723383,I723400,I723417,I723213,I1092496,I723457,I723465,I723482,I723499,I723516,I723216,I723547,I1092475,I723564,I723590,I723598,I723198,I723629,I723207,I723660,I723677,I723219,I723708,I1092493,I723210,I723201,I723204,I723222,I723808,I723834,I723842,I723859,I723876,I723902,I723910,I723936,I723944,I723961,I723978,I723995,I724035,I724043,I724060,I724077,I724094,I724125,I724142,I724168,I724176,I724207,I724238,I724255,I724286,I724386,I1268626,I724412,I724420,I724437,I1268650,I1268632,I724454,I1268638,I724480,I724488,I1268644,I1268629,I724514,I724522,I724539,I724556,I724573,I724369,I1268641,I724613,I724621,I724638,I724655,I724672,I724372,I724703,I1268647,I1268635,I724720,I724746,I724754,I724354,I724785,I724363,I724816,I724833,I724375,I724864,I724366,I724357,I724360,I724378,I724964,I724990,I724998,I725015,I725032,I725058,I725066,I725092,I725100,I725117,I725134,I725151,I725191,I725199,I725216,I725233,I725250,I725281,I725298,I725324,I725332,I725363,I725394,I725411,I725442,I725542,I725568,I725576,I725593,I725610,I725636,I725644,I725670,I725678,I725695,I725712,I725729,I725769,I725777,I725794,I725811,I725828,I725859,I725876,I725902,I725910,I725941,I725972,I725989,I726020,I726120,I726146,I726154,I726171,I726188,I726214,I726222,I726248,I726256,I726273,I726290,I726307,I726103,I726347,I726355,I726372,I726389,I726406,I726106,I726437,I726454,I726480,I726488,I726088,I726519,I726097,I726550,I726567,I726109,I726598,I726100,I726091,I726094,I726112,I726698,I957363,I726724,I726732,I726749,I957339,I957354,I726766,I957366,I726792,I726800,I957351,I957342,I726826,I726834,I726851,I726868,I726885,I726681,I726925,I726933,I726950,I726967,I726984,I726684,I727015,I957357,I957348,I727032,I957360,I727058,I727066,I726666,I727097,I726675,I727128,I727145,I726687,I727176,I957345,I726678,I726669,I726672,I726690,I727276,I727302,I727310,I727327,I727344,I727370,I727378,I727404,I727412,I727429,I727446,I727463,I727259,I727503,I727511,I727528,I727545,I727562,I727262,I727593,I727610,I727636,I727644,I727244,I727675,I727253,I727706,I727723,I727265,I727754,I727256,I727247,I727250,I727268,I727854,I885657,I727880,I727888,I727905,I885633,I885648,I727922,I885660,I727948,I727956,I885645,I885636,I727982,I727990,I728007,I728024,I728041,I727837,I728081,I728089,I728106,I728123,I728140,I727840,I728171,I885651,I885642,I728188,I885654,I728214,I728222,I727822,I728253,I727831,I728284,I728301,I727843,I728332,I885639,I727834,I727825,I727828,I727846,I728432,I728458,I728466,I728483,I728500,I728526,I728534,I728560,I728568,I728585,I728602,I728619,I728659,I728667,I728684,I728701,I728718,I728749,I728766,I728792,I728800,I728831,I728862,I728879,I728910,I729010,I729036,I729044,I729061,I729078,I729104,I729112,I729138,I729146,I729163,I729180,I729197,I729237,I729245,I729262,I729279,I729296,I729327,I729344,I729370,I729378,I729409,I729440,I729457,I729488,I729588,I1225378,I729614,I729622,I729639,I1225381,I1225390,I729656,I1225393,I729682,I729690,I1225402,I1225384,I729716,I729724,I729741,I729758,I729775,I729571,I729815,I729823,I729840,I729857,I729874,I729574,I729905,I1225399,I729922,I1225396,I729948,I729956,I729556,I729987,I729565,I730018,I730035,I729577,I730066,I1225387,I729568,I729559,I729562,I729580,I730166,I1146822,I730192,I730200,I730217,I1146804,I1146816,I730234,I1146819,I730260,I730268,I1146813,I1146810,I730294,I730302,I730319,I730336,I730353,I730149,I1146828,I730393,I730401,I730418,I730435,I730452,I730152,I730483,I1146807,I730500,I730526,I730534,I730134,I730565,I730143,I730596,I730613,I730155,I730644,I1146825,I730146,I730137,I730140,I730158,I730744,I1172832,I730770,I730778,I730795,I1172814,I1172826,I730812,I1172829,I730838,I730846,I1172823,I1172820,I730872,I730880,I730897,I730914,I730931,I730727,I1172838,I730971,I730979,I730996,I731013,I731030,I730730,I731061,I1172817,I731078,I731104,I731112,I730712,I731143,I730721,I731174,I731191,I730733,I731222,I1172835,I730724,I730715,I730718,I730736,I731322,I731348,I731356,I731373,I731390,I731416,I731424,I731450,I731458,I731475,I731492,I731509,I731305,I731549,I731557,I731574,I731591,I731608,I731308,I731639,I731656,I731682,I731690,I731290,I731721,I731299,I731752,I731769,I731311,I731800,I731302,I731293,I731296,I731314,I731900,I1024733,I731926,I731934,I731951,I1024730,I1024748,I731968,I1024745,I731994,I732002,I1024727,I732028,I732036,I732053,I732070,I732087,I1024739,I732127,I732135,I732152,I732169,I732186,I732217,I1024742,I732234,I732260,I732268,I732299,I732330,I732347,I732378,I1024736,I732478,I845477,I732504,I732512,I732529,I845465,I845483,I732546,I845480,I732572,I732580,I845471,I845468,I732606,I732614,I732631,I732648,I732665,I845462,I732705,I732713,I732730,I732747,I732764,I732795,I732812,I732838,I732846,I732877,I732908,I732925,I732956,I845474,I733056,I1142198,I733082,I733090,I733107,I1142180,I1142192,I733124,I1142195,I733150,I733158,I1142189,I1142186,I733184,I733192,I733209,I733226,I733243,I733039,I1142204,I733283,I733291,I733308,I733325,I733342,I733042,I733373,I1142183,I733390,I733416,I733424,I733024,I733455,I733033,I733486,I733503,I733045,I733534,I1142201,I733036,I733027,I733030,I733048,I733634,I1309504,I733660,I733668,I733685,I1309489,I1309477,I733702,I1309492,I733728,I733736,I1309495,I733762,I733770,I733787,I733804,I733821,I733617,I1309483,I733861,I733869,I733886,I733903,I733920,I733620,I733951,I1309480,I1309486,I733968,I1309501,I733994,I734002,I733602,I734033,I733611,I734064,I734081,I733623,I734112,I1309498,I733614,I733605,I733608,I733626,I734212,I734238,I734246,I734263,I734280,I734306,I734314,I734340,I734348,I734365,I734382,I734399,I734439,I734447,I734464,I734481,I734498,I734529,I734546,I734572,I734580,I734611,I734642,I734659,I734690,I734790,I734816,I734824,I734841,I734858,I734884,I734892,I734918,I734926,I734943,I734960,I734977,I735017,I735025,I735042,I735059,I735076,I735107,I735124,I735150,I735158,I735189,I735220,I735237,I735268,I735368,I1229186,I735394,I735402,I735419,I1229189,I1229198,I735436,I1229201,I735462,I735470,I1229210,I1229192,I735496,I735504,I735521,I735538,I735555,I735595,I735603,I735620,I735637,I735654,I735685,I1229207,I735702,I1229204,I735728,I735736,I735767,I735798,I735815,I735846,I1229195,I735946,I735972,I735980,I735997,I736014,I736040,I736048,I736074,I736082,I736099,I736116,I736133,I736173,I736181,I736198,I736215,I736232,I736263,I736280,I736306,I736314,I736345,I736376,I736393,I736424,I736524,I736550,I736558,I736575,I736592,I736618,I736626,I736652,I736660,I736677,I736694,I736711,I736751,I736759,I736776,I736793,I736810,I736841,I736858,I736884,I736892,I736923,I736954,I736971,I737002,I737102,I940567,I737128,I737136,I737153,I940543,I940558,I737170,I940570,I737196,I737204,I940555,I940546,I737230,I737238,I737255,I737272,I737289,I737329,I737337,I737354,I737371,I737388,I737419,I940561,I940552,I737436,I940564,I737462,I737470,I737501,I737532,I737549,I737580,I940549,I737680,I737706,I737714,I737731,I737748,I737774,I737782,I737808,I737816,I737833,I737850,I737867,I737663,I737907,I737915,I737932,I737949,I737966,I737666,I737997,I738014,I738040,I738048,I737648,I738079,I737657,I738110,I738127,I737669,I738158,I737660,I737651,I737654,I737672,I738258,I738284,I738292,I738309,I738326,I738352,I738360,I738386,I738394,I738411,I738428,I738445,I738241,I738485,I738493,I738510,I738527,I738544,I738244,I738575,I738592,I738618,I738626,I738226,I738657,I738235,I738688,I738705,I738247,I738736,I738238,I738229,I738232,I738250,I738836,I841788,I738862,I738870,I738887,I841776,I841794,I738904,I841791,I738930,I738938,I841782,I841779,I738964,I738972,I738989,I739006,I739023,I841773,I739063,I739071,I739088,I739105,I739122,I739153,I739170,I739196,I739204,I739235,I739266,I739283,I739314,I841785,I739414,I739440,I739448,I739465,I739482,I739508,I739516,I739542,I739550,I739567,I739584,I739601,I739641,I739649,I739666,I739683,I739700,I739731,I739748,I739774,I739782,I739813,I739844,I739861,I739892,I739992,I740018,I740026,I740043,I740060,I740086,I740094,I740120,I740128,I740145,I740162,I740179,I739975,I740219,I740227,I740244,I740261,I740278,I739978,I740309,I740326,I740352,I740360,I739960,I740391,I739969,I740422,I740439,I739981,I740470,I739972,I739963,I739966,I739984,I740570,I1382689,I740596,I740604,I740621,I1382674,I1382662,I740638,I1382677,I740664,I740672,I1382680,I740698,I740706,I740723,I740740,I740757,I1382668,I740797,I740805,I740822,I740839,I740856,I740887,I1382665,I1382671,I740904,I1382686,I740930,I740938,I740969,I741000,I741017,I741048,I1382683,I741148,I933461,I741174,I741182,I741199,I933437,I933452,I741216,I933464,I741242,I741250,I933449,I933440,I741276,I741284,I741301,I741318,I741335,I741131,I741375,I741383,I741400,I741417,I741434,I741134,I741465,I933455,I933446,I741482,I933458,I741508,I741516,I741116,I741547,I741125,I741578,I741595,I741137,I741626,I933443,I741128,I741119,I741122,I741140,I741726,I741752,I741760,I741777,I741794,I741820,I741828,I741854,I741862,I741879,I741896,I741913,I741709,I741953,I741961,I741978,I741995,I742012,I741712,I742043,I742060,I742086,I742094,I741694,I742125,I741703,I742156,I742173,I741715,I742204,I741706,I741697,I741700,I741718,I742304,I742330,I742338,I742355,I742372,I742398,I742406,I742432,I742440,I742457,I742474,I742491,I742287,I742531,I742539,I742556,I742573,I742590,I742290,I742621,I742638,I742664,I742672,I742272,I742703,I742281,I742734,I742751,I742293,I742782,I742284,I742275,I742278,I742296,I742882,I1156070,I742908,I742916,I742933,I1156052,I1156064,I742950,I1156067,I742976,I742984,I1156061,I1156058,I743010,I743018,I743035,I743052,I743069,I742865,I1156076,I743109,I743117,I743134,I743151,I743168,I742868,I743199,I1156055,I743216,I743242,I743250,I742850,I743281,I742859,I743312,I743329,I742871,I743360,I1156073,I742862,I742853,I742856,I742874,I743460,I743486,I743494,I743511,I743528,I743554,I743562,I743588,I743596,I743613,I743630,I743647,I743687,I743695,I743712,I743729,I743746,I743777,I743794,I743820,I743828,I743859,I743890,I743907,I743938,I744038,I744064,I744072,I744089,I744106,I744132,I744140,I744166,I744174,I744191,I744208,I744225,I744265,I744273,I744290,I744307,I744324,I744355,I744372,I744398,I744406,I744437,I744468,I744485,I744516,I744616,I1351749,I744642,I744650,I744667,I1351734,I1351722,I744684,I1351737,I744710,I744718,I1351740,I744744,I744752,I744769,I744786,I744803,I744599,I1351728,I744843,I744851,I744868,I744885,I744902,I744602,I744933,I1351725,I1351731,I744950,I1351746,I744976,I744984,I744584,I745015,I744593,I745046,I745063,I744605,I745094,I1351743,I744596,I744587,I744590,I744608,I745194,I745220,I745228,I745245,I745262,I745288,I745296,I745322,I745330,I745347,I745364,I745381,I745421,I745429,I745446,I745463,I745480,I745511,I745528,I745554,I745562,I745593,I745624,I745641,I745672,I745772,I745798,I745806,I745823,I745840,I745866,I745874,I745900,I745908,I745925,I745942,I745959,I745999,I746007,I746024,I746041,I746058,I746089,I746106,I746132,I746140,I746171,I746202,I746219,I746250,I746350,I1189594,I746376,I746384,I746401,I1189576,I1189588,I746418,I1189591,I746444,I746452,I1189585,I1189582,I746478,I746486,I746503,I746520,I746537,I746333,I1189600,I746577,I746585,I746602,I746619,I746636,I746336,I746667,I1189579,I746684,I746710,I746718,I746318,I746749,I746327,I746780,I746797,I746339,I746828,I1189597,I746330,I746321,I746324,I746342,I746928,I1069370,I746954,I746962,I746979,I1069352,I1069364,I746996,I1069367,I747022,I747030,I1069361,I1069358,I747056,I747064,I747081,I747098,I747115,I1069376,I747155,I747163,I747180,I747197,I747214,I747245,I1069355,I747262,I747288,I747296,I747327,I747358,I747375,I747406,I1069373,I747506,I795939,I747532,I747540,I747557,I795927,I795945,I747574,I795942,I747600,I747608,I795933,I795930,I747634,I747642,I747659,I747676,I747693,I795924,I747733,I747741,I747758,I747775,I747792,I747823,I747840,I747866,I747874,I747905,I747936,I747953,I747984,I795936,I748084,I1102894,I748110,I748118,I748135,I1102876,I1102888,I748152,I1102891,I748178,I748186,I1102885,I1102882,I748212,I748220,I748237,I748254,I748271,I748067,I1102900,I748311,I748319,I748336,I748353,I748370,I748070,I748401,I1102879,I748418,I748444,I748452,I748052,I748483,I748061,I748514,I748531,I748073,I748562,I1102897,I748064,I748055,I748058,I748076,I748662,I748688,I748696,I748713,I748730,I748756,I748764,I748790,I748798,I748815,I748832,I748849,I748645,I748889,I748897,I748914,I748931,I748948,I748648,I748979,I748996,I749022,I749030,I748630,I749061,I748639,I749092,I749109,I748651,I749140,I748642,I748633,I748636,I748654,I749240,I1110986,I749266,I749274,I749291,I1110968,I1110980,I749308,I1110983,I749334,I749342,I1110977,I1110974,I749368,I749376,I749393,I749410,I749427,I1110992,I749467,I749475,I749492,I749509,I749526,I749557,I1110971,I749574,I749600,I749608,I749639,I749670,I749687,I749718,I1110989,I749818,I749844,I749852,I749869,I749886,I749912,I749920,I749946,I749954,I749971,I749988,I750005,I750045,I750053,I750070,I750087,I750104,I750135,I750152,I750178,I750186,I750217,I750248,I750265,I750296,I750396,I750422,I750430,I750447,I750464,I750490,I750498,I750524,I750532,I750549,I750566,I750583,I750623,I750631,I750648,I750665,I750682,I750713,I750730,I750756,I750764,I750795,I750826,I750843,I750874,I750974,I751000,I751008,I751025,I751042,I751068,I751076,I751102,I751110,I751127,I751144,I751161,I750957,I751201,I751209,I751226,I751243,I751260,I750960,I751291,I751308,I751334,I751342,I750942,I751373,I750951,I751404,I751421,I750963,I751452,I750954,I750945,I750948,I750966,I751552,I751578,I751586,I751603,I751620,I751646,I751654,I751680,I751688,I751705,I751722,I751739,I751535,I751779,I751787,I751804,I751821,I751838,I751538,I751869,I751886,I751912,I751920,I751520,I751951,I751529,I751982,I751999,I751541,I752030,I751532,I751523,I751526,I751544,I752130,I752156,I752164,I752181,I752198,I752224,I752232,I752258,I752266,I752283,I752300,I752317,I752357,I752365,I752382,I752399,I752416,I752447,I752464,I752490,I752498,I752529,I752560,I752577,I752608,I752708,I752734,I752742,I752759,I752776,I752802,I752810,I752836,I752844,I752861,I752878,I752895,I752935,I752943,I752960,I752977,I752994,I753025,I753042,I753068,I753076,I753107,I753138,I753155,I753186,I753286,I1193062,I753312,I753320,I753337,I1193044,I1193056,I753354,I1193059,I753380,I753388,I1193053,I1193050,I753414,I753422,I753439,I753456,I753473,I1193068,I753513,I753521,I753538,I753555,I753572,I753603,I1193047,I753620,I753646,I753654,I753685,I753716,I753733,I753764,I1193065,I753864,I753890,I753898,I753915,I753932,I753958,I753966,I753992,I754000,I754017,I754034,I754051,I754091,I754099,I754116,I754133,I754150,I754181,I754198,I754224,I754232,I754263,I754294,I754311,I754342,I754442,I754468,I754476,I754493,I754510,I754536,I754544,I754570,I754578,I754595,I754612,I754629,I754425,I754669,I754677,I754694,I754711,I754728,I754428,I754759,I754776,I754802,I754810,I754410,I754841,I754419,I754872,I754889,I754431,I754920,I754422,I754413,I754416,I754434,I755020,I1090178,I755046,I755054,I755071,I1090160,I1090172,I755088,I1090175,I755114,I755122,I1090169,I1090166,I755148,I755156,I755173,I755190,I755207,I755003,I1090184,I755247,I755255,I755272,I755289,I755306,I755006,I755337,I1090163,I755354,I755380,I755388,I754988,I755419,I754997,I755450,I755467,I755009,I755498,I1090181,I755000,I754991,I754994,I755012,I755598,I755624,I755632,I755649,I755666,I755692,I755700,I755726,I755734,I755751,I755768,I755785,I755825,I755833,I755850,I755867,I755884,I755915,I755932,I755958,I755966,I755997,I756028,I756045,I756076,I756176,I1388639,I756202,I756210,I756227,I1388624,I1388612,I756244,I1388627,I756270,I756278,I1388630,I756304,I756312,I756329,I756346,I756363,I756159,I1388618,I756403,I756411,I756428,I756445,I756462,I756162,I756493,I1388615,I1388621,I756510,I1388636,I756536,I756544,I756144,I756575,I756153,I756606,I756623,I756165,I756654,I1388633,I756156,I756147,I756150,I756168,I756754,I1065902,I756780,I756788,I756805,I1065884,I1065896,I756822,I1065899,I756848,I756856,I1065893,I1065890,I756882,I756890,I756907,I756924,I756941,I756737,I1065908,I756981,I756989,I757006,I757023,I757040,I756740,I757071,I1065887,I757088,I757114,I757122,I756722,I757153,I756731,I757184,I757201,I756743,I757232,I1065905,I756734,I756725,I756728,I756746,I757332,I757358,I757366,I757383,I757400,I757426,I757434,I757460,I757468,I757485,I757502,I757519,I757559,I757567,I757584,I757601,I757618,I757649,I757666,I757692,I757700,I757731,I757762,I757779,I757810,I757910,I757936,I757944,I757961,I757978,I758004,I758012,I758038,I758046,I758063,I758080,I758097,I758137,I758145,I758162,I758179,I758196,I758227,I758244,I758270,I758278,I758309,I758340,I758357,I758388,I758488,I1335684,I758514,I758522,I758539,I1335669,I1335657,I758556,I1335672,I758582,I758590,I1335675,I758616,I758624,I758641,I758658,I758675,I758471,I1335663,I758715,I758723,I758740,I758757,I758774,I758474,I758805,I1335660,I1335666,I758822,I1335681,I758848,I758856,I758456,I758887,I758465,I758918,I758935,I758477,I758966,I1335678,I758468,I758459,I758462,I758480,I759066,I1021367,I759092,I759100,I759117,I1021364,I1021382,I759134,I1021379,I759160,I759168,I1021361,I759194,I759202,I759219,I759236,I759253,I1021373,I759293,I759301,I759318,I759335,I759352,I759383,I1021376,I759400,I759426,I759434,I759465,I759496,I759513,I759544,I1021370,I759644,I1271516,I759670,I759678,I759695,I1271540,I1271522,I759712,I1271528,I759738,I759746,I1271534,I1271519,I759772,I759780,I759797,I759814,I759831,I1271531,I759871,I759879,I759896,I759913,I759930,I759961,I1271537,I1271525,I759978,I760004,I760012,I760043,I760074,I760091,I760122,I760222,I1145088,I760248,I760256,I760273,I1145070,I1145082,I760290,I1145085,I760316,I760324,I1145079,I1145076,I760350,I760358,I760375,I760392,I760409,I1145094,I760449,I760457,I760474,I760491,I760508,I760539,I1145073,I760556,I760582,I760590,I760621,I760652,I760669,I760700,I1145091,I760800,I760826,I760834,I760851,I760868,I760894,I760902,I760928,I760936,I760953,I760970,I760987,I761027,I761035,I761052,I761069,I761086,I761117,I761134,I761160,I761168,I761199,I761230,I761247,I761278,I761378,I761404,I761412,I761429,I761446,I761472,I761480,I761506,I761514,I761531,I761548,I761565,I761605,I761613,I761630,I761647,I761664,I761695,I761712,I761738,I761746,I761777,I761808,I761825,I761856,I761956,I800155,I761982,I761990,I762007,I800143,I800161,I762024,I800158,I762050,I762058,I800149,I800146,I762084,I762092,I762109,I762126,I762143,I761939,I800140,I762183,I762191,I762208,I762225,I762242,I761942,I762273,I762290,I762316,I762324,I761924,I762355,I761933,I762386,I762403,I761945,I762434,I800152,I761936,I761927,I761930,I761948,I762534,I836518,I762560,I762568,I762585,I836506,I836524,I762602,I836521,I762628,I762636,I836512,I836509,I762662,I762670,I762687,I762704,I762721,I836503,I762761,I762769,I762786,I762803,I762820,I762851,I762868,I762894,I762902,I762933,I762964,I762981,I763012,I836515,I763112,I763138,I763146,I763163,I763180,I763206,I763214,I763240,I763248,I763265,I763282,I763299,I763095,I763339,I763347,I763364,I763381,I763398,I763098,I763429,I763446,I763472,I763480,I763080,I763511,I763089,I763542,I763559,I763101,I763590,I763092,I763083,I763086,I763104,I763690,I763716,I763724,I763741,I763758,I763784,I763792,I763818,I763826,I763843,I763860,I763877,I763673,I763917,I763925,I763942,I763959,I763976,I763676,I764007,I764024,I764050,I764058,I763658,I764089,I763667,I764120,I764137,I763679,I764168,I763670,I763661,I763664,I763682,I764268,I764294,I764302,I764319,I764336,I764362,I764370,I764396,I764404,I764421,I764438,I764455,I764251,I764495,I764503,I764520,I764537,I764554,I764254,I764585,I764602,I764628,I764636,I764236,I764667,I764245,I764698,I764715,I764257,I764746,I764248,I764239,I764242,I764260,I764846,I986433,I764872,I764880,I764897,I986409,I986424,I764914,I986436,I764940,I764948,I986421,I986412,I764974,I764982,I764999,I765016,I765033,I765073,I765081,I765098,I765115,I765132,I765163,I986427,I986418,I765180,I986430,I765206,I765214,I765245,I765276,I765293,I765324,I986415,I765424,I765450,I765458,I765475,I765492,I765518,I765526,I765552,I765560,I765577,I765594,I765611,I765651,I765659,I765676,I765693,I765710,I765741,I765758,I765784,I765792,I765823,I765854,I765871,I765902,I766002,I878678,I766028,I766036,I766053,I878666,I878684,I766070,I878681,I766096,I766104,I878672,I878669,I766130,I766138,I766155,I766172,I766189,I765985,I878663,I766229,I766237,I766254,I766271,I766288,I765988,I766319,I766336,I766362,I766370,I765970,I766401,I765979,I766432,I766449,I765991,I766480,I878675,I765982,I765973,I765976,I765994,I766580,I1007105,I766606,I766614,I766631,I1007081,I1007096,I766648,I1007108,I766674,I766682,I1007093,I1007084,I766708,I766716,I766733,I766750,I766767,I766563,I766807,I766815,I766832,I766849,I766866,I766566,I766897,I1007099,I1007090,I766914,I1007102,I766940,I766948,I766548,I766979,I766557,I767010,I767027,I766569,I767058,I1007087,I766560,I766551,I766554,I766572,I767158,I767184,I767192,I767209,I767226,I767252,I767260,I767286,I767294,I767311,I767328,I767345,I767141,I767385,I767393,I767410,I767427,I767444,I767144,I767475,I767492,I767518,I767526,I767126,I767557,I767135,I767588,I767605,I767147,I767636,I767138,I767129,I767132,I767150,I767736,I767762,I767770,I767787,I767804,I767830,I767838,I767864,I767872,I767889,I767906,I767923,I767719,I767963,I767971,I767988,I768005,I768022,I767722,I768053,I768070,I768096,I768104,I767704,I768135,I767713,I768166,I768183,I767725,I768214,I767716,I767707,I767710,I767728,I768314,I1068214,I768340,I768348,I768365,I1068196,I1068208,I768382,I1068211,I768408,I768416,I1068205,I1068202,I768442,I768450,I768467,I768484,I768501,I768297,I1068220,I768541,I768549,I768566,I768583,I768600,I768300,I768631,I1068199,I768648,I768674,I768682,I768282,I768713,I768291,I768744,I768761,I768303,I768792,I1068217,I768294,I768285,I768288,I768306,I768892,I1049978,I768918,I768926,I768943,I1049975,I1049993,I768960,I1049990,I768986,I768994,I1049972,I769020,I769028,I769045,I769062,I769079,I1049984,I769119,I769127,I769144,I769161,I769178,I769209,I1049987,I769226,I769252,I769260,I769291,I769322,I769339,I769370,I1049981,I769470,I769496,I769504,I769521,I769538,I769564,I769572,I769598,I769606,I769623,I769640,I769657,I769697,I769705,I769722,I769739,I769756,I769787,I769804,I769830,I769838,I769869,I769900,I769917,I769948,I770048,I872354,I770074,I770082,I770099,I872342,I872360,I770116,I872357,I770142,I770150,I872348,I872345,I770176,I770184,I770201,I770218,I770235,I770031,I872339,I770275,I770283,I770300,I770317,I770334,I770034,I770365,I770382,I770408,I770416,I770016,I770447,I770025,I770478,I770495,I770037,I770526,I872351,I770028,I770019,I770022,I770040,I770626,I770652,I770660,I770677,I770694,I770720,I770728,I770754,I770762,I770779,I770796,I770813,I770853,I770861,I770878,I770895,I770912,I770943,I770960,I770986,I770994,I771025,I771056,I771073,I771104,I771204,I771230,I771238,I771255,I771272,I771298,I771306,I771332,I771340,I771357,I771374,I771391,I771431,I771439,I771456,I771473,I771490,I771521,I771538,I771564,I771572,I771603,I771634,I771651,I771682,I771782,I771808,I771816,I771833,I771850,I771876,I771884,I771910,I771918,I771935,I771952,I771969,I771765,I772009,I772017,I772034,I772051,I772068,I771768,I772099,I772116,I772142,I772150,I771750,I772181,I771759,I772212,I772229,I771771,I772260,I771762,I771753,I771756,I771774,I772360,I879732,I772386,I772394,I772411,I879720,I879738,I772428,I879735,I772454,I772462,I879726,I879723,I772488,I772496,I772513,I772530,I772547,I772343,I879717,I772587,I772595,I772612,I772629,I772646,I772346,I772677,I772694,I772720,I772728,I772328,I772759,I772337,I772790,I772807,I772349,I772838,I879729,I772340,I772331,I772334,I772352,I772938,I813330,I772964,I772972,I772989,I813318,I813336,I773006,I813333,I773032,I773040,I813324,I813321,I773066,I773074,I773091,I773108,I773125,I772921,I813315,I773165,I773173,I773190,I773207,I773224,I772924,I773255,I773272,I773298,I773306,I772906,I773337,I772915,I773368,I773385,I772927,I773416,I813327,I772918,I772909,I772912,I772930,I773516,I1288856,I773542,I773550,I773567,I1288880,I1288862,I773584,I1288868,I773610,I773618,I1288874,I1288859,I773644,I773652,I773669,I773686,I773703,I773499,I1288871,I773743,I773751,I773768,I773785,I773802,I773502,I773833,I1288877,I1288865,I773850,I773876,I773884,I773484,I773915,I773493,I773946,I773963,I773505,I773994,I773496,I773487,I773490,I773508,I774094,I774120,I774128,I774145,I774162,I774188,I774196,I774222,I774230,I774247,I774264,I774281,I774077,I774321,I774329,I774346,I774363,I774380,I774080,I774411,I774428,I774454,I774462,I774062,I774493,I774071,I774524,I774541,I774083,I774572,I774074,I774065,I774068,I774086,I774672,I1037636,I774698,I774706,I774723,I1037633,I1037651,I774740,I1037648,I774766,I774774,I1037630,I774800,I774808,I774825,I774842,I774859,I1037642,I774899,I774907,I774924,I774941,I774958,I774989,I1037645,I775006,I775032,I775040,I775071,I775102,I775119,I775150,I1037639,I775250,I775276,I775284,I775301,I775318,I775344,I775352,I775378,I775386,I775403,I775420,I775437,I775477,I775485,I775502,I775519,I775536,I775567,I775584,I775610,I775618,I775649,I775680,I775697,I775728,I775828,I1014635,I775854,I775862,I775879,I1014632,I1014650,I775896,I1014647,I775922,I775930,I1014629,I775956,I775964,I775981,I775998,I776015,I775811,I1014641,I776055,I776063,I776080,I776097,I776114,I775814,I776145,I1014644,I776162,I776188,I776196,I775796,I776227,I775805,I776258,I776275,I775817,I776306,I1014638,I775808,I775799,I775802,I775820,I776406,I776432,I776440,I776457,I776474,I776500,I776508,I776534,I776542,I776559,I776576,I776593,I776633,I776641,I776658,I776675,I776692,I776723,I776740,I776766,I776774,I776805,I776836,I776853,I776884,I776981,I1042127,I777007,I777015,I777032,I1042136,I1042124,I777049,I1042121,I777075,I776970,I777106,I777114,I1042118,I777131,I777157,I777165,I776973,I777205,I776964,I776955,I777241,I1042139,I1042130,I777258,I1042133,I777284,I777292,I777309,I776958,I777340,I777357,I777374,I776967,I777405,I776952,I777436,I777453,I776961,I777508,I777534,I777542,I777559,I777576,I777602,I777497,I777633,I777641,I777658,I777684,I777692,I777500,I777732,I777491,I777482,I777768,I777785,I777811,I777819,I777836,I777485,I777867,I777884,I777901,I777494,I777932,I777479,I777963,I777980,I777488,I778035,I778061,I778069,I778086,I778103,I778129,I778160,I778168,I778185,I778211,I778219,I778259,I778295,I778312,I778338,I778346,I778363,I778394,I778411,I778428,I778459,I778490,I778507,I778562,I778588,I778596,I778613,I778630,I778656,I778687,I778695,I778712,I778738,I778746,I778786,I778822,I778839,I778865,I778873,I778890,I778921,I778938,I778955,I778986,I779017,I779034,I779089,I779115,I779123,I779140,I779157,I779183,I779078,I779214,I779222,I779239,I779265,I779273,I779081,I779313,I779072,I779063,I779349,I779366,I779392,I779400,I779417,I779066,I779448,I779465,I779482,I779075,I779513,I779060,I779544,I779561,I779069,I779616,I779642,I779650,I779667,I779684,I779710,I779741,I779749,I779766,I779792,I779800,I779840,I779876,I779893,I779919,I779927,I779944,I779975,I779992,I780009,I780040,I780071,I780088,I780143,I1306517,I780169,I780177,I780194,I1306514,I1306523,I780211,I1306502,I780237,I780132,I1306505,I780268,I780276,I1306520,I780293,I780319,I780327,I780135,I1306526,I780367,I780126,I780117,I780403,I1306508,I1306529,I780420,I1306511,I780446,I780454,I780471,I780120,I780502,I780519,I780536,I780129,I780567,I780114,I780598,I780615,I780123,I780670,I780696,I780704,I780721,I780738,I780764,I780659,I780795,I780803,I780820,I780846,I780854,I780662,I780894,I780653,I780644,I780930,I780947,I780973,I780981,I780998,I780647,I781029,I781046,I781063,I780656,I781094,I780641,I781125,I781142,I780650,I781197,I1391007,I781223,I781231,I781248,I1391004,I1391013,I781265,I1390992,I781291,I1390995,I781322,I781330,I1391010,I781347,I781373,I781381,I1391016,I781421,I781457,I1390998,I1391019,I781474,I1391001,I781500,I781508,I781525,I781556,I781573,I781590,I781621,I781652,I781669,I781724,I1216142,I781750,I781758,I781775,I1216148,I1216130,I781792,I1216139,I781818,I1216145,I781849,I781857,I1216133,I781874,I781900,I781908,I1216151,I781948,I781984,I1216136,I782001,I1216154,I782027,I782035,I782052,I782083,I782100,I782117,I782148,I782179,I782196,I782251,I950236,I782277,I782285,I782302,I950251,I950233,I782319,I782345,I950242,I782376,I782384,I950260,I782401,I782427,I782435,I950257,I782475,I782511,I950254,I950245,I782528,I950239,I782554,I782562,I782579,I782610,I950248,I782627,I782644,I782675,I782706,I782723,I782778,I782804,I782812,I782829,I782846,I782872,I782903,I782911,I782928,I782954,I782962,I783002,I783038,I783055,I783081,I783089,I783106,I783137,I783154,I783171,I783202,I783233,I783250,I783305,I783331,I783339,I783356,I783373,I783399,I783430,I783438,I783455,I783481,I783489,I783529,I783565,I783582,I783608,I783616,I783633,I783664,I783681,I783698,I783729,I783760,I783777,I783832,I1361257,I783858,I783866,I783883,I1361254,I1361263,I783900,I1361242,I783926,I1361245,I783957,I783965,I1361260,I783982,I784008,I784016,I1361266,I784056,I784092,I1361248,I1361269,I784109,I1361251,I784135,I784143,I784160,I784191,I784208,I784225,I784256,I784287,I784304,I784359,I1330317,I784385,I784393,I784410,I1330314,I1330323,I784427,I1330302,I784453,I784348,I1330305,I784484,I784492,I1330320,I784509,I784535,I784543,I784351,I1330326,I784583,I784342,I784333,I784619,I1330308,I1330329,I784636,I1330311,I784662,I784670,I784687,I784336,I784718,I784735,I784752,I784345,I784783,I784330,I784814,I784831,I784339,I784886,I1238990,I784912,I784920,I784937,I1238996,I1238978,I784954,I1238987,I784980,I784875,I1238993,I785011,I785019,I1238981,I785036,I785062,I785070,I784878,I1238999,I785110,I784869,I784860,I785146,I1238984,I785163,I1239002,I785189,I785197,I785214,I784863,I785245,I785262,I785279,I784872,I785310,I784857,I785341,I785358,I784866,I785413,I785439,I785447,I785464,I785481,I785507,I785538,I785546,I785563,I785589,I785597,I785637,I785673,I785690,I785716,I785724,I785741,I785772,I785789,I785806,I785837,I785868,I785885,I785940,I785966,I785974,I785991,I786008,I786034,I785929,I786065,I786073,I786090,I786116,I786124,I785932,I786164,I785923,I785914,I786200,I786217,I786243,I786251,I786268,I785917,I786299,I786316,I786333,I785926,I786364,I785911,I786395,I786412,I785920,I786467,I786493,I786501,I786518,I786535,I786561,I786592,I786600,I786617,I786643,I786651,I786691,I786727,I786744,I786770,I786778,I786795,I786826,I786843,I786860,I786891,I786922,I786939,I786994,I1349357,I787020,I787028,I787045,I1349354,I1349363,I787062,I1349342,I787088,I1349345,I787119,I787127,I1349360,I787144,I787170,I787178,I1349366,I787218,I787254,I1349348,I1349369,I787271,I1349351,I787297,I787305,I787322,I787353,I787370,I787387,I787418,I787449,I787466,I787521,I1236814,I787547,I787555,I787572,I1236820,I1236802,I787589,I1236811,I787615,I787510,I1236817,I787646,I787654,I1236805,I787671,I787697,I787705,I787513,I1236823,I787745,I787504,I787495,I787781,I1236808,I787798,I1236826,I787824,I787832,I787849,I787498,I787880,I787897,I787914,I787507,I787945,I787492,I787976,I787993,I787501,I788048,I788074,I788082,I788099,I788116,I788142,I788037,I788173,I788181,I788198,I788224,I788232,I788040,I788272,I788031,I788022,I788308,I788325,I788351,I788359,I788376,I788025,I788407,I788424,I788441,I788034,I788472,I788019,I788503,I788520,I788028,I788575,I1246062,I788601,I788609,I788626,I1246068,I1246050,I788643,I1246059,I788669,I788564,I1246065,I788700,I788708,I1246053,I788725,I788751,I788759,I788567,I1246071,I788799,I788558,I788549,I788835,I1246056,I788852,I1246074,I788878,I788886,I788903,I788552,I788934,I788951,I788968,I788561,I788999,I788546,I789030,I789047,I788555,I789102,I1304791,I789128,I789136,I789153,I1304785,I1304803,I789170,I1304788,I789196,I789091,I1304809,I789227,I789235,I1304794,I789252,I789278,I789286,I789094,I1304806,I789326,I789085,I789076,I789362,I1304797,I1304812,I789379,I1304800,I789405,I789413,I789430,I789079,I789461,I789478,I789495,I789088,I789526,I789073,I789557,I789574,I789082,I789629,I789655,I789663,I789680,I789697,I789723,I789618,I789754,I789762,I789779,I789805,I789813,I789621,I789853,I789612,I789603,I789889,I789906,I789932,I789940,I789957,I789606,I789988,I790005,I790022,I789615,I790053,I789600,I790084,I790101,I789609,I790156,I790182,I790190,I790207,I790224,I790250,I790145,I790281,I790289,I790306,I790332,I790340,I790148,I790380,I790139,I790130,I790416,I790433,I790459,I790467,I790484,I790133,I790515,I790532,I790549,I790142,I790580,I790127,I790611,I790628,I790136,I790683,I790709,I790717,I790734,I790751,I790777,I790808,I790816,I790833,I790859,I790867,I790907,I790943,I790960,I790986,I790994,I791011,I791042,I791059,I791076,I791107,I791138,I791155,I791210,I791236,I791244,I791261,I791278,I791304,I791335,I791343,I791360,I791386,I791394,I791434,I791470,I791487,I791513,I791521,I791538,I791569,I791586,I791603,I791634,I791665,I791682,I791737,I928918,I791763,I791771,I791788,I928933,I928915,I791805,I791831,I791726,I928924,I791862,I791870,I928942,I791887,I791913,I791921,I791729,I928939,I791961,I791720,I791711,I791997,I928936,I928927,I792014,I928921,I792040,I792048,I792065,I791714,I792096,I928930,I792113,I792130,I791723,I792161,I791708,I792192,I792209,I791717,I792264,I792290,I792298,I792315,I792332,I792358,I792389,I792397,I792414,I792440,I792448,I792488,I792524,I792541,I792567,I792575,I792592,I792623,I792640,I792657,I792688,I792719,I792736,I792791,I792817,I792825,I792842,I792859,I792885,I792916,I792924,I792941,I792967,I792975,I793015,I793051,I793068,I793094,I793102,I793119,I793150,I793167,I793184,I793215,I793246,I793263,I793318,I793344,I793352,I793369,I793386,I793412,I793443,I793451,I793468,I793494,I793502,I793542,I793578,I793595,I793621,I793629,I793646,I793677,I793694,I793711,I793742,I793773,I793790,I793845,I793871,I793879,I793896,I793913,I793939,I793834,I793970,I793978,I793995,I794021,I794029,I793837,I794069,I793828,I793819,I794105,I794122,I794148,I794156,I794173,I793822,I794204,I794221,I794238,I793831,I794269,I793816,I794300,I794317,I793825,I794372,I794398,I794406,I794423,I794440,I794466,I794497,I794505,I794522,I794548,I794556,I794596,I794632,I794649,I794675,I794683,I794700,I794731,I794748,I794765,I794796,I794827,I794844,I794899,I794925,I794933,I794950,I794967,I794993,I795024,I795032,I795049,I795075,I795083,I795123,I795159,I795176,I795202,I795210,I795227,I795258,I795275,I795292,I795323,I795354,I795371,I795426,I795452,I795460,I795477,I795494,I795520,I795415,I795551,I795559,I795576,I795602,I795610,I795418,I795650,I795409,I795400,I795686,I795703,I795729,I795737,I795754,I795403,I795785,I795802,I795819,I795412,I795850,I795397,I795881,I795898,I795406,I795953,I1178612,I795979,I795987,I796004,I1178594,I796021,I1178600,I796047,I1178597,I796078,I796086,I1178606,I796103,I796129,I796137,I1178618,I796177,I796213,I1178609,I1178603,I796230,I796256,I796264,I796281,I796312,I1178615,I796329,I796346,I796377,I796408,I796425,I796480,I796506,I796514,I796531,I796548,I796574,I796605,I796613,I796630,I796656,I796664,I796704,I796740,I796757,I796783,I796791,I796808,I796839,I796856,I796873,I796904,I796935,I796952,I797007,I1215054,I797033,I797041,I797058,I1215060,I1215042,I797075,I1215051,I797101,I796996,I1215057,I797132,I797140,I1215045,I797157,I797183,I797191,I796999,I1215063,I797231,I796990,I796981,I797267,I1215048,I797284,I1215066,I797310,I797318,I797335,I796984,I797366,I797383,I797400,I796993,I797431,I796978,I797462,I797479,I796987,I797534,I797560,I797568,I797585,I797602,I797628,I797659,I797667,I797684,I797710,I797718,I797758,I797794,I797811,I797837,I797845,I797862,I797893,I797910,I797927,I797958,I797989,I798006,I798061,I995456,I798087,I798095,I798112,I995471,I995453,I798129,I798155,I995462,I798186,I798194,I995480,I798211,I798237,I798245,I995477,I798285,I798321,I995474,I995465,I798338,I995459,I798364,I798372,I798389,I798420,I995468,I798437,I798454,I798485,I798516,I798533,I798588,I798614,I798622,I798639,I798656,I798682,I798713,I798721,I798738,I798764,I798772,I798812,I798848,I798865,I798891,I798899,I798916,I798947,I798964,I798981,I799012,I799043,I799060,I799115,I1027541,I799141,I799149,I799166,I1027550,I1027538,I799183,I1027535,I799209,I799104,I799240,I799248,I1027532,I799265,I799291,I799299,I799107,I799339,I799098,I799089,I799375,I1027553,I1027544,I799392,I1027547,I799418,I799426,I799443,I799092,I799474,I799491,I799508,I799101,I799539,I799086,I799570,I799587,I799095,I799642,I799668,I799676,I799693,I799710,I799736,I799767,I799775,I799792,I799818,I799826,I799866,I799902,I799919,I799945,I799953,I799970,I800001,I800018,I800035,I800066,I800097,I800114,I800169,I1104628,I800195,I800203,I800220,I1104610,I800237,I1104616,I800263,I1104613,I800294,I800302,I1104622,I800319,I800345,I800353,I1104634,I800393,I800429,I1104625,I1104619,I800446,I800472,I800480,I800497,I800528,I1104631,I800545,I800562,I800593,I800624,I800641,I800696,I999978,I800722,I800730,I800747,I999993,I999975,I800764,I800790,I999984,I800821,I800829,I1000002,I800846,I800872,I800880,I999999,I800920,I800956,I999996,I999987,I800973,I999981,I800999,I801007,I801024,I801055,I999990,I801072,I801089,I801120,I801151,I801168,I801223,I801249,I801257,I801274,I801291,I801317,I801348,I801356,I801373,I801399,I801407,I801447,I801483,I801500,I801526,I801534,I801551,I801582,I801599,I801616,I801647,I801678,I801695,I801750,I801776,I801784,I801801,I801818,I801844,I801739,I801875,I801883,I801900,I801926,I801934,I801742,I801974,I801733,I801724,I802010,I802027,I802053,I802061,I802078,I801727,I802109,I802126,I802143,I801736,I802174,I801721,I802205,I802222,I801730,I802277,I802303,I802311,I802328,I802345,I802371,I802266,I802402,I802410,I802427,I802453,I802461,I802269,I802501,I802260,I802251,I802537,I802554,I802580,I802588,I802605,I802254,I802636,I802653,I802670,I802263,I802701,I802248,I802732,I802749,I802257,I802804,I802830,I802838,I802855,I802872,I802898,I802793,I802929,I802937,I802954,I802980,I802988,I802796,I803028,I802787,I802778,I803064,I803081,I803107,I803115,I803132,I802781,I803163,I803180,I803197,I802790,I803228,I802775,I803259,I803276,I802784,I803331,I803357,I803365,I803382,I803399,I803425,I803320,I803456,I803464,I803481,I803507,I803515,I803323,I803555,I803314,I803305,I803591,I803608,I803634,I803642,I803659,I803308,I803690,I803707,I803724,I803317,I803755,I803302,I803786,I803803,I803311,I803858,I803884,I803892,I803909,I803926,I803952,I803847,I803983,I803991,I804008,I804034,I804042,I803850,I804082,I803841,I803832,I804118,I804135,I804161,I804169,I804186,I803835,I804217,I804234,I804251,I803844,I804282,I803829,I804313,I804330,I803838,I804385,I1279048,I804411,I804419,I804436,I1279030,I1279033,I804453,I1279045,I804479,I1279054,I804510,I804518,I1279039,I804535,I804561,I804569,I1279051,I804609,I804645,I1279042,I1279036,I804662,I804688,I804696,I804713,I804744,I804761,I804778,I804809,I804840,I804857,I804912,I1272690,I804938,I804946,I804963,I1272672,I1272675,I804980,I1272687,I805006,I1272696,I805037,I805045,I1272681,I805062,I805088,I805096,I1272693,I805136,I805172,I1272684,I1272678,I805189,I805215,I805223,I805240,I805271,I805288,I805305,I805336,I805367,I805384,I805439,I805465,I805473,I805490,I805507,I805533,I805564,I805572,I805589,I805615,I805623,I805663,I805699,I805716,I805742,I805750,I805767,I805798,I805815,I805832,I805863,I805894,I805911,I805966,I805992,I806000,I806017,I806034,I806060,I805955,I806091,I806099,I806116,I806142,I806150,I805958,I806190,I805949,I805940,I806226,I806243,I806269,I806277,I806294,I805943,I806325,I806342,I806359,I805952,I806390,I805937,I806421,I806438,I805946,I806493,I806519,I806527,I806544,I806561,I806587,I806482,I806618,I806626,I806643,I806669,I806677,I806485,I806717,I806476,I806467,I806753,I806770,I806796,I806804,I806821,I806470,I806852,I806869,I806886,I806479,I806917,I806464,I806948,I806965,I806473,I807020,I807046,I807054,I807071,I807088,I807114,I807145,I807153,I807170,I807196,I807204,I807244,I807280,I807297,I807323,I807331,I807348,I807379,I807396,I807413,I807444,I807475,I807492,I807547,I1339242,I807573,I807581,I807598,I1339239,I1339248,I807615,I1339227,I807641,I1339230,I807672,I807680,I1339245,I807697,I807723,I807731,I1339251,I807771,I807807,I1339233,I1339254,I807824,I1339236,I807850,I807858,I807875,I807906,I807923,I807940,I807971,I808002,I808019,I808074,I808100,I808108,I808125,I808142,I808168,I808063,I808199,I808207,I808224,I808250,I808258,I808066,I808298,I808057,I808048,I808334,I808351,I808377,I808385,I808402,I808051,I808433,I808450,I808467,I808060,I808498,I808045,I808529,I808546,I808054,I808601,I1127170,I808627,I808635,I808652,I1127152,I808669,I1127158,I808695,I808590,I1127155,I808726,I808734,I1127164,I808751,I808777,I808785,I808593,I1127176,I808825,I808584,I808575,I808861,I1127167,I1127161,I808878,I808904,I808912,I808929,I808578,I808960,I1127173,I808977,I808994,I808587,I809025,I808572,I809056,I809073,I808581,I809128,I809154,I809162,I809179,I809196,I809222,I809253,I809261,I809278,I809304,I809312,I809352,I809388,I809405,I809431,I809439,I809456,I809487,I809504,I809521,I809552,I809583,I809600,I809655,I809681,I809689,I809706,I809723,I809749,I809644,I809780,I809788,I809805,I809831,I809839,I809647,I809879,I809638,I809629,I809915,I809932,I809958,I809966,I809983,I809632,I810014,I810031,I810048,I809641,I810079,I809626,I810110,I810127,I809635,I810182,I810208,I810216,I810233,I810250,I810276,I810307,I810315,I810332,I810358,I810366,I810406,I810442,I810459,I810485,I810493,I810510,I810541,I810558,I810575,I810606,I810637,I810654,I810709,I810735,I810743,I810760,I810777,I810803,I810698,I810834,I810842,I810859,I810885,I810893,I810701,I810933,I810692,I810683,I810969,I810986,I811012,I811020,I811037,I810686,I811068,I811085,I811102,I810695,I811133,I810680,I811164,I811181,I810689,I811236,I811262,I811270,I811287,I811304,I811330,I811361,I811369,I811386,I811412,I811420,I811460,I811496,I811513,I811539,I811547,I811564,I811595,I811612,I811629,I811660,I811691,I811708,I811763,I811789,I811797,I811814,I811831,I811857,I811888,I811896,I811913,I811939,I811947,I811987,I812023,I812040,I812066,I812074,I812091,I812122,I812139,I812156,I812187,I812218,I812235,I812290,I1112142,I812316,I812324,I812341,I1112124,I812358,I1112130,I812384,I1112127,I812415,I812423,I1112136,I812440,I812466,I812474,I1112148,I812514,I812550,I1112139,I1112133,I812567,I812593,I812601,I812618,I812649,I1112145,I812666,I812683,I812714,I812745,I812762,I812817,I812843,I812851,I812868,I812885,I812911,I812942,I812950,I812967,I812993,I813001,I813041,I813077,I813094,I813120,I813128,I813145,I813176,I813193,I813210,I813241,I813272,I813289,I813344,I813370,I813378,I813395,I813412,I813438,I813469,I813477,I813494,I813520,I813528,I813568,I813604,I813621,I813647,I813655,I813672,I813703,I813720,I813737,I813768,I813799,I813816,I813871,I1160116,I813897,I813905,I813922,I1160098,I813939,I1160104,I813965,I813860,I1160101,I813996,I814004,I1160110,I814021,I814047,I814055,I813863,I1160122,I814095,I813854,I813845,I814131,I1160113,I1160107,I814148,I814174,I814182,I814199,I813848,I814230,I1160119,I814247,I814264,I813857,I814295,I813842,I814326,I814343,I813851,I814398,I814424,I814432,I814449,I814466,I814492,I814523,I814531,I814548,I814574,I814582,I814622,I814658,I814675,I814701,I814709,I814726,I814757,I814774,I814791,I814822,I814853,I814870,I814925,I1100004,I814951,I814959,I814976,I1099986,I814993,I1099992,I815019,I1099989,I815050,I815058,I1099998,I815075,I815101,I815109,I1100010,I815149,I815185,I1100001,I1099995,I815202,I815228,I815236,I815253,I815284,I1100007,I815301,I815318,I815349,I815380,I815397,I815452,I815478,I815486,I815503,I815520,I815546,I815441,I815577,I815585,I815602,I815628,I815636,I815444,I815676,I815435,I815426,I815712,I815729,I815755,I815763,I815780,I815429,I815811,I815828,I815845,I815438,I815876,I815423,I815907,I815924,I815432,I815979,I816005,I816013,I816030,I816047,I816073,I816104,I816112,I816129,I816155,I816163,I816203,I816239,I816256,I816282,I816290,I816307,I816338,I816355,I816372,I816403,I816434,I816451,I816506,I816532,I816540,I816557,I816574,I816600,I816631,I816639,I816656,I816682,I816690,I816730,I816766,I816783,I816809,I816817,I816834,I816865,I816882,I816899,I816930,I816961,I816978,I817033,I817059,I817067,I817084,I817101,I817127,I817022,I817158,I817166,I817183,I817209,I817217,I817025,I817257,I817016,I817007,I817293,I817310,I817336,I817344,I817361,I817010,I817392,I817409,I817426,I817019,I817457,I817004,I817488,I817505,I817013,I817560,I817586,I817594,I817611,I817628,I817654,I817549,I817685,I817693,I817710,I817736,I817744,I817552,I817784,I817543,I817534,I817820,I817837,I817863,I817871,I817888,I817537,I817919,I817936,I817953,I817546,I817984,I817531,I818015,I818032,I817540,I818087,I818113,I818121,I818138,I818155,I818181,I818076,I818212,I818220,I818237,I818263,I818271,I818079,I818311,I818070,I818061,I818347,I818364,I818390,I818398,I818415,I818064,I818446,I818463,I818480,I818073,I818511,I818058,I818542,I818559,I818067,I818614,I818640,I818648,I818665,I818682,I818708,I818739,I818747,I818764,I818790,I818798,I818838,I818874,I818891,I818917,I818925,I818942,I818973,I818990,I819007,I819038,I819069,I819086,I819141,I819167,I819175,I819192,I819209,I819235,I819266,I819274,I819291,I819317,I819325,I819365,I819401,I819418,I819444,I819452,I819469,I819500,I819517,I819534,I819565,I819596,I819613,I819668,I819694,I819702,I819719,I819736,I819762,I819793,I819801,I819818,I819844,I819852,I819892,I819928,I819945,I819971,I819979,I819996,I820027,I820044,I820061,I820092,I820123,I820140,I820195,I820221,I820229,I820246,I820263,I820289,I820320,I820328,I820345,I820371,I820379,I820419,I820455,I820472,I820498,I820506,I820523,I820554,I820571,I820588,I820619,I820650,I820667,I820722,I820748,I820756,I820773,I820790,I820816,I820711,I820847,I820855,I820872,I820898,I820906,I820714,I820946,I820705,I820696,I820982,I820999,I821025,I821033,I821050,I820699,I821081,I821098,I821115,I820708,I821146,I820693,I821177,I821194,I820702,I821249,I821275,I821283,I821300,I821317,I821343,I821238,I821374,I821382,I821399,I821425,I821433,I821241,I821473,I821232,I821223,I821509,I821526,I821552,I821560,I821577,I821226,I821608,I821625,I821642,I821235,I821673,I821220,I821704,I821721,I821229,I821776,I897910,I821802,I821810,I821827,I897925,I897907,I821844,I821870,I821765,I897916,I821901,I821909,I897934,I821926,I821952,I821960,I821768,I897931,I822000,I821759,I821750,I822036,I897928,I897919,I822053,I897913,I822079,I822087,I822104,I821753,I822135,I897922,I822152,I822169,I821762,I822200,I821747,I822231,I822248,I821756,I822303,I822329,I822337,I822354,I822371,I822397,I822428,I822436,I822453,I822479,I822487,I822527,I822563,I822580,I822606,I822614,I822631,I822662,I822679,I822696,I822727,I822758,I822775,I822830,I822856,I822864,I822881,I822898,I822924,I822819,I822955,I822963,I822980,I823006,I823014,I822822,I823054,I822813,I822804,I823090,I823107,I823133,I823141,I823158,I822807,I823189,I823206,I823223,I822816,I823254,I822801,I823285,I823302,I822810,I823357,I1282516,I823383,I823391,I823408,I1282498,I1282501,I823425,I1282513,I823451,I823346,I1282522,I823482,I823490,I1282507,I823507,I823533,I823541,I823349,I1282519,I823581,I823340,I823331,I823617,I1282510,I1282504,I823634,I823660,I823668,I823685,I823334,I823716,I823733,I823750,I823343,I823781,I823328,I823812,I823829,I823337,I823884,I823910,I823918,I823935,I823952,I823978,I824009,I824017,I824034,I824060,I824068,I824108,I824144,I824161,I824187,I824195,I824212,I824243,I824260,I824277,I824308,I824339,I824356,I824411,I1136996,I824437,I824445,I824462,I1136978,I824479,I1136984,I824505,I824400,I1136981,I824536,I824544,I1136990,I824561,I824587,I824595,I824403,I1137002,I824635,I824394,I824385,I824671,I1136993,I1136987,I824688,I824714,I824722,I824739,I824388,I824770,I1136999,I824787,I824804,I824397,I824835,I824382,I824866,I824883,I824391,I824938,I948298,I824964,I824972,I824989,I948313,I948295,I825006,I825032,I948304,I825063,I825071,I948322,I825088,I825114,I825122,I948319,I825162,I825198,I948316,I948307,I825215,I948301,I825241,I825249,I825266,I825297,I948310,I825314,I825331,I825362,I825393,I825410,I825465,I1324367,I825491,I825499,I825516,I1324364,I1324373,I825533,I1324352,I825559,I825454,I1324355,I825590,I825598,I1324370,I825615,I825641,I825649,I825457,I1324376,I825689,I825448,I825439,I825725,I1324358,I1324379,I825742,I1324361,I825768,I825776,I825793,I825442,I825824,I825841,I825858,I825451,I825889,I825436,I825920,I825937,I825445,I825992,I1047737,I826018,I826026,I826043,I1047746,I1047734,I826060,I1047731,I826086,I825981,I826117,I826125,I1047728,I826142,I826168,I826176,I825984,I826216,I825975,I825966,I826252,I1047749,I1047740,I826269,I1047743,I826295,I826303,I826320,I825969,I826351,I826368,I826385,I825978,I826416,I825963,I826447,I826464,I825972,I826519,I826545,I826553,I826570,I826587,I826613,I826644,I826652,I826669,I826695,I826703,I826743,I826779,I826796,I826822,I826830,I826847,I826878,I826895,I826912,I826943,I826974,I826991,I827046,I1163584,I827072,I827080,I827097,I1163566,I827114,I1163572,I827140,I827035,I1163569,I827171,I827179,I1163578,I827196,I827222,I827230,I827038,I1163590,I827270,I827029,I827020,I827306,I1163581,I1163575,I827323,I827349,I827357,I827374,I827023,I827405,I1163587,I827422,I827439,I827032,I827470,I827017,I827501,I827518,I827026,I827573,I827599,I827607,I827624,I827641,I827667,I827562,I827698,I827706,I827723,I827749,I827757,I827565,I827797,I827556,I827547,I827833,I827850,I827876,I827884,I827901,I827550,I827932,I827949,I827966,I827559,I827997,I827544,I828028,I828045,I827553,I828100,I980598,I828126,I828134,I828151,I980613,I980595,I828168,I828194,I980604,I828225,I828233,I980622,I828250,I828276,I828284,I980619,I828324,I828360,I980616,I980607,I828377,I980601,I828403,I828411,I828428,I828459,I980610,I828476,I828493,I828524,I828555,I828572,I828627,I828653,I828661,I828678,I828695,I828721,I828616,I828752,I828760,I828777,I828803,I828811,I828619,I828851,I828610,I828601,I828887,I828904,I828930,I828938,I828955,I828604,I828986,I829003,I829020,I828613,I829051,I828598,I829082,I829099,I828607,I829154,I1143354,I829180,I829188,I829205,I1143336,I829222,I1143342,I829248,I1143339,I829279,I829287,I1143348,I829304,I829330,I829338,I1143360,I829378,I829414,I1143351,I1143345,I829431,I829457,I829465,I829482,I829513,I1143357,I829530,I829547,I829578,I829609,I829626,I829681,I1070526,I829707,I829715,I829732,I1070508,I829749,I1070514,I829775,I1070511,I829806,I829814,I1070520,I829831,I829857,I829865,I1070532,I829905,I829941,I1070523,I1070517,I829958,I829984,I829992,I830009,I830040,I1070529,I830057,I830074,I830105,I830136,I830153,I830208,I1284250,I830234,I830242,I830259,I1284232,I1284235,I830276,I1284247,I830302,I830197,I1284256,I830333,I830341,I1284241,I830358,I830384,I830392,I830200,I1284253,I830432,I830191,I830182,I830468,I1284244,I1284238,I830485,I830511,I830519,I830536,I830185,I830567,I830584,I830601,I830194,I830632,I830179,I830663,I830680,I830188,I830735,I1064746,I830761,I830769,I830786,I1064728,I830803,I1064734,I830829,I830724,I1064731,I830860,I830868,I1064740,I830885,I830911,I830919,I830727,I1064752,I830959,I830718,I830709,I830995,I1064743,I1064737,I831012,I831038,I831046,I831063,I830712,I831094,I1064749,I831111,I831128,I830721,I831159,I830706,I831190,I831207,I830715,I831262,I831288,I831296,I831313,I831330,I831356,I831387,I831395,I831412,I831438,I831446,I831486,I831522,I831539,I831565,I831573,I831590,I831621,I831638,I831655,I831686,I831717,I831734,I831789,I898556,I831815,I831823,I831840,I898571,I898553,I831857,I831883,I831778,I898562,I831914,I831922,I898580,I831939,I831965,I831973,I831781,I898577,I832013,I831772,I831763,I832049,I898574,I898565,I832066,I898559,I832092,I832100,I832117,I831766,I832148,I898568,I832165,I832182,I831775,I832213,I831760,I832244,I832261,I831769,I832316,I832342,I832350,I832367,I832384,I832410,I832441,I832449,I832466,I832492,I832500,I832540,I832576,I832593,I832619,I832627,I832644,I832675,I832692,I832709,I832740,I832771,I832788,I832843,I832869,I832877,I832894,I832911,I832937,I832968,I832976,I832993,I833019,I833027,I833067,I833103,I833120,I833146,I833154,I833171,I833202,I833219,I833236,I833267,I833298,I833315,I833370,I1315442,I833396,I833404,I833421,I1315439,I1315448,I833438,I1315427,I833464,I1315430,I833495,I833503,I1315445,I833520,I833546,I833554,I1315451,I833594,I833630,I1315433,I1315454,I833647,I1315436,I833673,I833681,I833698,I833729,I833746,I833763,I833794,I833825,I833842,I833897,I1354117,I833923,I833931,I833948,I1354114,I1354123,I833965,I1354102,I833991,I1354105,I834022,I834030,I1354120,I834047,I834073,I834081,I1354126,I834121,I834157,I1354108,I1354129,I834174,I1354111,I834200,I834208,I834225,I834256,I834273,I834290,I834321,I834352,I834369,I834424,I834450,I834458,I834475,I834492,I834518,I834549,I834557,I834574,I834600,I834608,I834648,I834684,I834701,I834727,I834735,I834752,I834783,I834800,I834817,I834848,I834879,I834896,I834951,I1264020,I834977,I834985,I835002,I1264002,I1264005,I835019,I1264017,I835045,I1264026,I835076,I835084,I1264011,I835101,I835127,I835135,I1264023,I835175,I835211,I1264014,I1264008,I835228,I835254,I835262,I835279,I835310,I835327,I835344,I835375,I835406,I835423,I835478,I835504,I835512,I835529,I835546,I835572,I835467,I835603,I835611,I835628,I835654,I835662,I835470,I835702,I835461,I835452,I835738,I835755,I835781,I835789,I835806,I835455,I835837,I835854,I835871,I835464,I835902,I835449,I835933,I835950,I835458,I836005,I1035395,I836031,I836039,I836056,I1035404,I1035392,I836073,I1035389,I836099,I836130,I836138,I1035386,I836155,I836181,I836189,I836229,I836265,I1035407,I1035398,I836282,I1035401,I836308,I836316,I836333,I836364,I836381,I836398,I836429,I836460,I836477,I836532,I836558,I836566,I836583,I836600,I836626,I836657,I836665,I836682,I836708,I836716,I836756,I836792,I836809,I836835,I836843,I836860,I836891,I836908,I836925,I836956,I836987,I837004,I837059,I921166,I837085,I837093,I837110,I921181,I921163,I837127,I837153,I837048,I921172,I837184,I837192,I921190,I837209,I837235,I837243,I837051,I921187,I837283,I837042,I837033,I837319,I921184,I921175,I837336,I921169,I837362,I837370,I837387,I837036,I837418,I921178,I837435,I837452,I837045,I837483,I837030,I837514,I837531,I837039,I837586,I837612,I837620,I837637,I837654,I837680,I837575,I837711,I837719,I837736,I837762,I837770,I837578,I837810,I837569,I837560,I837846,I837863,I837889,I837897,I837914,I837563,I837945,I837962,I837979,I837572,I838010,I837557,I838041,I838058,I837566,I838113,I838139,I838147,I838164,I838181,I838207,I838238,I838246,I838263,I838289,I838297,I838337,I838373,I838390,I838416,I838424,I838441,I838472,I838489,I838506,I838537,I838568,I838585,I838640,I838666,I838674,I838691,I838708,I838734,I838765,I838773,I838790,I838816,I838824,I838864,I838900,I838917,I838943,I838951,I838968,I838999,I839016,I839033,I839064,I839095,I839112,I839167,I1392197,I839193,I839201,I839218,I1392194,I1392203,I839235,I1392182,I839261,I839156,I1392185,I839292,I839300,I1392200,I839317,I839343,I839351,I839159,I1392206,I839391,I839150,I839141,I839427,I1392188,I1392209,I839444,I1392191,I839470,I839478,I839495,I839144,I839526,I839543,I839560,I839153,I839591,I839138,I839622,I839639,I839147,I839694,I839720,I839728,I839745,I839762,I839788,I839819,I839827,I839844,I839870,I839878,I839918,I839954,I839971,I839997,I840005,I840022,I840053,I840070,I840087,I840118,I840149,I840166,I840221,I840247,I840255,I840272,I840289,I840315,I840210,I840346,I840354,I840371,I840397,I840405,I840213,I840445,I840204,I840195,I840481,I840498,I840524,I840532,I840549,I840198,I840580,I840597,I840614,I840207,I840645,I840192,I840676,I840693,I840201,I840748,I1350547,I840774,I840782,I840799,I1350544,I1350553,I840816,I1350532,I840842,I840737,I1350535,I840873,I840881,I1350550,I840898,I840924,I840932,I840740,I1350556,I840972,I840731,I840722,I841008,I1350538,I1350559,I841025,I1350541,I841051,I841059,I841076,I840725,I841107,I841124,I841141,I840734,I841172,I840719,I841203,I841220,I840728,I841275,I841301,I841309,I841326,I841343,I841369,I841400,I841408,I841425,I841451,I841459,I841499,I841535,I841552,I841578,I841586,I841603,I841634,I841651,I841668,I841699,I841730,I841747,I841802,I841828,I841836,I841853,I841870,I841896,I841927,I841935,I841952,I841978,I841986,I842026,I842062,I842079,I842105,I842113,I842130,I842161,I842178,I842195,I842226,I842257,I842274,I842329,I1219406,I842355,I842363,I842380,I1219412,I1219394,I842397,I1219403,I842423,I1219409,I842454,I842462,I1219397,I842479,I842505,I842513,I1219415,I842553,I842589,I1219400,I842606,I1219418,I842632,I842640,I842657,I842688,I842705,I842722,I842753,I842784,I842801,I842856,I842882,I842890,I842907,I842924,I842950,I842981,I842989,I843006,I843032,I843040,I843080,I843116,I843133,I843159,I843167,I843184,I843215,I843232,I843249,I843280,I843311,I843328,I843383,I843409,I843417,I843434,I843451,I843477,I843508,I843516,I843533,I843559,I843567,I843607,I843643,I843660,I843686,I843694,I843711,I843742,I843759,I843776,I843807,I843838,I843855,I843910,I1049420,I843936,I843944,I843961,I1049429,I1049417,I843978,I1049414,I844004,I844035,I844043,I1049411,I844060,I844086,I844094,I844134,I844170,I1049432,I1049423,I844187,I1049426,I844213,I844221,I844238,I844269,I844286,I844303,I844334,I844365,I844382,I844437,I844463,I844471,I844488,I844505,I844531,I844426,I844562,I844570,I844587,I844613,I844621,I844429,I844661,I844420,I844411,I844697,I844714,I844740,I844748,I844765,I844414,I844796,I844813,I844830,I844423,I844861,I844408,I844892,I844909,I844417,I844964,I844990,I844998,I845015,I845032,I845058,I845089,I845097,I845114,I845140,I845148,I845188,I845224,I845241,I845267,I845275,I845292,I845323,I845340,I845357,I845388,I845419,I845436,I845491,I845517,I845525,I845542,I845559,I845585,I845616,I845624,I845641,I845667,I845675,I845715,I845751,I845768,I845794,I845802,I845819,I845850,I845867,I845884,I845915,I845946,I845963,I846018,I1279626,I846044,I846052,I846069,I1279608,I1279611,I846086,I1279623,I846112,I846007,I1279632,I846143,I846151,I1279617,I846168,I846194,I846202,I846010,I1279629,I846242,I846001,I845992,I846278,I1279620,I1279614,I846295,I846321,I846329,I846346,I845995,I846377,I846394,I846411,I846004,I846442,I845989,I846473,I846490,I845998,I846545,I846571,I846579,I846596,I846613,I846639,I846670,I846678,I846695,I846721,I846729,I846769,I846805,I846822,I846848,I846856,I846873,I846904,I846921,I846938,I846969,I847000,I847017,I847072,I847098,I847106,I847123,I847140,I847166,I847197,I847205,I847222,I847248,I847256,I847296,I847332,I847349,I847375,I847383,I847400,I847431,I847448,I847465,I847496,I847527,I847544,I847599,I847625,I847633,I847650,I847667,I847693,I847724,I847732,I847749,I847775,I847783,I847823,I847859,I847876,I847902,I847910,I847927,I847958,I847975,I847992,I848023,I848054,I848071,I848126,I848152,I848160,I848177,I848194,I848220,I848115,I848251,I848259,I848276,I848302,I848310,I848118,I848350,I848109,I848100,I848386,I848403,I848429,I848437,I848454,I848103,I848485,I848502,I848519,I848112,I848550,I848097,I848581,I848598,I848106,I848653,I848679,I848687,I848704,I848721,I848747,I848642,I848778,I848786,I848803,I848829,I848837,I848645,I848877,I848636,I848627,I848913,I848930,I848956,I848964,I848981,I848630,I849012,I849029,I849046,I848639,I849077,I848624,I849108,I849125,I848633,I849180,I1204622,I849206,I849214,I849231,I1204604,I849248,I1204610,I849274,I1204607,I849305,I849313,I1204616,I849330,I849356,I849364,I1204628,I849404,I849440,I1204619,I1204613,I849457,I849483,I849491,I849508,I849539,I1204625,I849556,I849573,I849604,I849635,I849652,I849707,I849733,I849741,I849758,I849775,I849801,I849696,I849832,I849840,I849857,I849883,I849891,I849699,I849931,I849690,I849681,I849967,I849984,I850010,I850018,I850035,I849684,I850066,I850083,I850100,I849693,I850131,I849678,I850162,I850179,I849687,I850234,I850260,I850268,I850285,I850302,I850328,I850359,I850367,I850384,I850410,I850418,I850458,I850494,I850511,I850537,I850545,I850562,I850593,I850610,I850627,I850658,I850689,I850706,I850761,I850787,I850795,I850812,I850829,I850855,I850886,I850894,I850911,I850937,I850945,I850985,I851021,I851038,I851064,I851072,I851089,I851120,I851137,I851154,I851185,I851216,I851233,I851288,I1265176,I851314,I851322,I851339,I1265158,I1265161,I851356,I1265173,I851382,I1265182,I851413,I851421,I1265167,I851438,I851464,I851472,I1265179,I851512,I851548,I1265170,I1265164,I851565,I851591,I851599,I851616,I851647,I851664,I851681,I851712,I851743,I851760,I851815,I851841,I851849,I851866,I851883,I851909,I851940,I851948,I851965,I851991,I851999,I852039,I852075,I852092,I852118,I852126,I852143,I852174,I852191,I852208,I852239,I852270,I852287,I852342,I852368,I852376,I852393,I852410,I852436,I852467,I852475,I852492,I852518,I852526,I852566,I852602,I852619,I852645,I852653,I852670,I852701,I852718,I852735,I852766,I852797,I852814,I852869,I1075150,I852895,I852903,I852920,I1075132,I852937,I1075138,I852963,I1075135,I852994,I853002,I1075144,I853019,I853045,I853053,I1075156,I853093,I853129,I1075147,I1075141,I853146,I853172,I853180,I853197,I853228,I1075153,I853245,I853262,I853293,I853324,I853341,I853396,I853422,I853430,I853447,I853464,I853490,I853521,I853529,I853546,I853572,I853580,I853620,I853656,I853673,I853699,I853707,I853724,I853755,I853772,I853789,I853820,I853851,I853868,I853923,I853949,I853957,I853974,I853991,I854017,I854048,I854056,I854073,I854099,I854107,I854147,I854183,I854200,I854226,I854234,I854251,I854282,I854299,I854316,I854347,I854378,I854395,I854450,I1380892,I854476,I854484,I854501,I1380889,I1380898,I854518,I1380877,I854544,I1380880,I854575,I854583,I1380895,I854600,I854626,I854634,I1380901,I854674,I854710,I1380883,I1380904,I854727,I1380886,I854753,I854761,I854778,I854809,I854826,I854843,I854874,I854905,I854922,I854977,I855003,I855011,I855028,I855045,I855071,I854966,I855102,I855110,I855127,I855153,I855161,I854969,I855201,I854960,I854951,I855237,I855254,I855280,I855288,I855305,I854954,I855336,I855353,I855370,I854963,I855401,I854948,I855432,I855449,I854957,I855504,I855530,I855538,I855555,I855572,I855598,I855629,I855637,I855654,I855680,I855688,I855728,I855764,I855781,I855807,I855815,I855832,I855863,I855880,I855897,I855928,I855959,I855976,I856031,I1183236,I856057,I856065,I856082,I1183218,I856099,I1183224,I856125,I1183221,I856156,I856164,I1183230,I856181,I856207,I856215,I1183242,I856255,I856291,I1183233,I1183227,I856308,I856334,I856342,I856359,I856390,I1183239,I856407,I856424,I856455,I856486,I856503,I856558,I856584,I856592,I856609,I856626,I856652,I856683,I856691,I856708,I856734,I856742,I856782,I856818,I856835,I856861,I856869,I856886,I856917,I856934,I856951,I856982,I857013,I857030,I857085,I978014,I857111,I857119,I857136,I978029,I978011,I857153,I857179,I857074,I978020,I857210,I857218,I978038,I857235,I857261,I857269,I857077,I978035,I857309,I857068,I857059,I857345,I978032,I978023,I857362,I978017,I857388,I857396,I857413,I857062,I857444,I978026,I857461,I857478,I857071,I857509,I857056,I857540,I857557,I857065,I857612,I997394,I857638,I857646,I857663,I997409,I997391,I857680,I857706,I857601,I997400,I857737,I857745,I997418,I857762,I857788,I857796,I857604,I997415,I857836,I857595,I857586,I857872,I997412,I997403,I857889,I997397,I857915,I857923,I857940,I857589,I857971,I997406,I857988,I858005,I857598,I858036,I857583,I858067,I858084,I857592,I858139,I1015199,I858165,I858173,I858190,I1015208,I1015196,I858207,I1015193,I858233,I858128,I858264,I858272,I1015190,I858289,I858315,I858323,I858131,I858363,I858122,I858113,I858399,I1015211,I1015202,I858416,I1015205,I858442,I858450,I858467,I858116,I858498,I858515,I858532,I858125,I858563,I858110,I858594,I858611,I858119,I858666,I858692,I858700,I858717,I858734,I858760,I858791,I858799,I858816,I858842,I858850,I858890,I858926,I858943,I858969,I858977,I858994,I859025,I859042,I859059,I859090,I859121,I859138,I859193,I890804,I859219,I859227,I859244,I890819,I890801,I859261,I859287,I859182,I890810,I859318,I859326,I890828,I859343,I859369,I859377,I859185,I890825,I859417,I859176,I859167,I859453,I890822,I890813,I859470,I890807,I859496,I859504,I859521,I859170,I859552,I890816,I859569,I859586,I859179,I859617,I859164,I859648,I859665,I859173,I859720,I859746,I859754,I859771,I859788,I859814,I859845,I859853,I859870,I859896,I859904,I859944,I859980,I859997,I860023,I860031,I860048,I860079,I860096,I860113,I860144,I860175,I860192,I860247,I860273,I860281,I860298,I860315,I860341,I860236,I860372,I860380,I860397,I860423,I860431,I860239,I860471,I860230,I860221,I860507,I860524,I860550,I860558,I860575,I860224,I860606,I860623,I860640,I860233,I860671,I860218,I860702,I860719,I860227,I860774,I923104,I860800,I860808,I860825,I923119,I923101,I860842,I860868,I923110,I860899,I860907,I923128,I860924,I860950,I860958,I923125,I860998,I861034,I923122,I923113,I861051,I923107,I861077,I861085,I861102,I861133,I923116,I861150,I861167,I861198,I861229,I861246,I861301,I861327,I861335,I861352,I861369,I861395,I861290,I861426,I861434,I861451,I861477,I861485,I861293,I861525,I861284,I861275,I861561,I861578,I861604,I861612,I861629,I861278,I861660,I861677,I861694,I861287,I861725,I861272,I861756,I861773,I861281,I861828,I1142776,I861854,I861862,I861879,I1142758,I861896,I1142764,I861922,I1142761,I861953,I861961,I1142770,I861978,I862004,I862012,I1142782,I862052,I862088,I1142773,I1142767,I862105,I862131,I862139,I862156,I862187,I1142779,I862204,I862221,I862252,I862283,I862300,I862355,I1028663,I862381,I862389,I862406,I1028672,I1028660,I862423,I1028657,I862449,I862344,I862480,I862488,I1028654,I862505,I862531,I862539,I862347,I862579,I862338,I862329,I862615,I1028675,I1028666,I862632,I1028669,I862658,I862666,I862683,I862332,I862714,I862731,I862748,I862341,I862779,I862326,I862810,I862827,I862335,I862882,I862908,I862916,I862933,I862950,I862976,I862871,I863007,I863015,I863032,I863058,I863066,I862874,I863106,I862865,I862856,I863142,I863159,I863185,I863193,I863210,I862859,I863241,I863258,I863275,I862868,I863306,I862853,I863337,I863354,I862862,I863409,I863435,I863443,I863460,I863477,I863503,I863534,I863542,I863559,I863585,I863593,I863633,I863669,I863686,I863712,I863720,I863737,I863768,I863785,I863802,I863833,I863864,I863881,I863936,I1301986,I863962,I863970,I863987,I1301980,I1301998,I864004,I1301983,I864030,I1302004,I864061,I864069,I1301989,I864086,I864112,I864120,I1302001,I864160,I864196,I1301992,I1302007,I864213,I1301995,I864239,I864247,I864264,I864295,I864312,I864329,I864360,I864391,I864408,I864463,I1249326,I864489,I864497,I864514,I1249332,I1249314,I864531,I1249323,I864557,I1249329,I864588,I864596,I1249317,I864613,I864639,I864647,I1249335,I864687,I864723,I1249320,I864740,I1249338,I864766,I864774,I864791,I864822,I864839,I864856,I864887,I864918,I864935,I864990,I865016,I865024,I865041,I865058,I865084,I865115,I865123,I865140,I865166,I865174,I865214,I865250,I865267,I865293,I865301,I865318,I865349,I865366,I865383,I865414,I865445,I865462,I865517,I1193640,I865543,I865551,I865568,I1193622,I865585,I1193628,I865611,I865506,I1193625,I865642,I865650,I1193634,I865667,I865693,I865701,I865509,I1193646,I865741,I865500,I865491,I865777,I1193637,I1193631,I865794,I865820,I865828,I865845,I865494,I865876,I1193643,I865893,I865910,I865503,I865941,I865488,I865972,I865989,I865497,I866044,I866070,I866078,I866095,I866112,I866138,I866169,I866177,I866194,I866220,I866228,I866268,I866304,I866321,I866347,I866355,I866372,I866403,I866420,I866437,I866468,I866499,I866516,I866571,I1131216,I866597,I866605,I866622,I1131198,I866639,I1131204,I866665,I1131201,I866696,I866704,I1131210,I866721,I866747,I866755,I1131222,I866795,I866831,I1131213,I1131207,I866848,I866874,I866882,I866899,I866930,I1131219,I866947,I866964,I866995,I867026,I867043,I867098,I867124,I867132,I867149,I867166,I867192,I867223,I867231,I867248,I867274,I867282,I867322,I867358,I867375,I867401,I867409,I867426,I867457,I867474,I867491,I867522,I867553,I867570,I867625,I867651,I867659,I867676,I867693,I867719,I867614,I867750,I867758,I867775,I867801,I867809,I867617,I867849,I867608,I867599,I867885,I867902,I867928,I867936,I867953,I867602,I867984,I868001,I868018,I867611,I868049,I867596,I868080,I868097,I867605,I868152,I868178,I868186,I868203,I868220,I868246,I868141,I868277,I868285,I868302,I868328,I868336,I868144,I868376,I868135,I868126,I868412,I868429,I868455,I868463,I868480,I868129,I868511,I868528,I868545,I868138,I868576,I868123,I868607,I868624,I868132,I868679,I1371372,I868705,I868713,I868730,I1371369,I1371378,I868747,I1371357,I868773,I868668,I1371360,I868804,I868812,I1371375,I868829,I868855,I868863,I868671,I1371381,I868903,I868662,I868653,I868939,I1371363,I1371384,I868956,I1371366,I868982,I868990,I869007,I868656,I869038,I869055,I869072,I868665,I869103,I868650,I869134,I869151,I868659,I869206,I869232,I869240,I869257,I869274,I869300,I869195,I869331,I869339,I869356,I869382,I869390,I869198,I869430,I869189,I869180,I869466,I869483,I869509,I869517,I869534,I869183,I869565,I869582,I869599,I869192,I869630,I869177,I869661,I869678,I869186,I869733,I869759,I869767,I869784,I869801,I869827,I869722,I869858,I869866,I869883,I869909,I869917,I869725,I869957,I869716,I869707,I869993,I870010,I870036,I870044,I870061,I869710,I870092,I870109,I870126,I869719,I870157,I869704,I870188,I870205,I869713,I870260,I870286,I870294,I870311,I870328,I870354,I870385,I870393,I870410,I870436,I870444,I870484,I870520,I870537,I870563,I870571,I870588,I870619,I870636,I870653,I870684,I870715,I870732,I870787,I870813,I870821,I870838,I870855,I870881,I870912,I870920,I870937,I870963,I870971,I871011,I871047,I871064,I871090,I871098,I871115,I871146,I871163,I871180,I871211,I871242,I871259,I871314,I1055591,I871340,I871348,I871365,I1055600,I1055588,I871382,I1055585,I871408,I871303,I871439,I871447,I1055582,I871464,I871490,I871498,I871306,I871538,I871297,I871288,I871574,I1055603,I1055594,I871591,I1055597,I871617,I871625,I871642,I871291,I871673,I871690,I871707,I871300,I871738,I871285,I871769,I871786,I871294,I871841,I871867,I871875,I871892,I871909,I871935,I871966,I871974,I871991,I872017,I872025,I872065,I872101,I872118,I872144,I872152,I872169,I872200,I872217,I872234,I872265,I872296,I872313,I872368,I872394,I872402,I872419,I872436,I872462,I872493,I872501,I872518,I872544,I872552,I872592,I872628,I872645,I872671,I872679,I872696,I872727,I872744,I872761,I872792,I872823,I872840,I872895,I872921,I872929,I872946,I872963,I872989,I873020,I873028,I873045,I873071,I873079,I873119,I873155,I873172,I873198,I873206,I873223,I873254,I873271,I873288,I873319,I873350,I873367,I873422,I962510,I873448,I873456,I873473,I962525,I962507,I873490,I873516,I873411,I962516,I873547,I873555,I962534,I873572,I873598,I873606,I873414,I962531,I873646,I873405,I873396,I873682,I962528,I962519,I873699,I962513,I873725,I873733,I873750,I873399,I873781,I962522,I873798,I873815,I873408,I873846,I873393,I873877,I873894,I873402,I873949,I1361852,I873975,I873983,I874000,I1361849,I1361858,I874017,I1361837,I874043,I1361840,I874074,I874082,I1361855,I874099,I874125,I874133,I1361861,I874173,I874209,I1361843,I1361864,I874226,I1361846,I874252,I874260,I874277,I874308,I874325,I874342,I874373,I874404,I874421,I874476,I874502,I874510,I874527,I874544,I874570,I874601,I874609,I874626,I874652,I874660,I874700,I874736,I874753,I874779,I874787,I874804,I874835,I874852,I874869,I874900,I874931,I874948,I875003,I875029,I875037,I875054,I875071,I875097,I875128,I875136,I875153,I875179,I875187,I875227,I875263,I875280,I875306,I875314,I875331,I875362,I875379,I875396,I875427,I875458,I875475,I875530,I875556,I875564,I875581,I875598,I875624,I875655,I875663,I875680,I875706,I875714,I875754,I875790,I875807,I875833,I875841,I875858,I875889,I875906,I875923,I875954,I875985,I876002,I876057,I876083,I876091,I876108,I876125,I876151,I876182,I876190,I876207,I876233,I876241,I876281,I876317,I876334,I876360,I876368,I876385,I876416,I876433,I876450,I876481,I876512,I876529,I876584,I876610,I876618,I876635,I876652,I876678,I876573,I876709,I876717,I876734,I876760,I876768,I876576,I876808,I876567,I876558,I876844,I876861,I876887,I876895,I876912,I876561,I876943,I876960,I876977,I876570,I877008,I876555,I877039,I877056,I876564,I877111,I877137,I877145,I877162,I877179,I877205,I877236,I877244,I877261,I877287,I877295,I877335,I877371,I877388,I877414,I877422,I877439,I877470,I877487,I877504,I877535,I877566,I877583,I877638,I877664,I877672,I877689,I877706,I877732,I877763,I877771,I877788,I877814,I877822,I877862,I877898,I877915,I877941,I877949,I877966,I877997,I878014,I878031,I878062,I878093,I878110,I878165,I1128326,I878191,I878199,I878216,I1128308,I878233,I1128314,I878259,I1128311,I878290,I878298,I1128320,I878315,I878341,I878349,I1128332,I878389,I878425,I1128323,I1128317,I878442,I878468,I878476,I878493,I878524,I1128329,I878541,I878558,I878589,I878620,I878637,I878692,I1093646,I878718,I878726,I878743,I1093628,I878760,I1093634,I878786,I1093631,I878817,I878825,I1093640,I878842,I878868,I878876,I1093652,I878916,I878952,I1093643,I1093637,I878969,I878995,I879003,I879020,I879051,I1093649,I879068,I879085,I879116,I879147,I879164,I879219,I879245,I879253,I879270,I879287,I879313,I879344,I879352,I879369,I879395,I879403,I879443,I879479,I879496,I879522,I879530,I879547,I879578,I879595,I879612,I879643,I879674,I879691,I879746,I879772,I879780,I879797,I879814,I879840,I879871,I879879,I879896,I879922,I879930,I879970,I880006,I880023,I880049,I880057,I880074,I880105,I880122,I880139,I880170,I880201,I880218,I880273,I1121390,I880299,I880307,I880324,I1121372,I880341,I1121378,I880367,I880262,I1121375,I880398,I880406,I1121384,I880423,I880449,I880457,I880265,I1121396,I880497,I880256,I880247,I880533,I1121387,I1121381,I880550,I880576,I880584,I880601,I880250,I880632,I1121393,I880649,I880666,I880259,I880697,I880244,I880728,I880745,I880253,I880800,I1285984,I880826,I880834,I880851,I1285966,I1285969,I880868,I1285981,I880894,I880789,I1285990,I880925,I880933,I1285975,I880950,I880976,I880984,I880792,I1285987,I881024,I880783,I880774,I881060,I1285978,I1285972,I881077,I881103,I881111,I881128,I880777,I881159,I881176,I881193,I880786,I881224,I880771,I881255,I881272,I880780,I881327,I881353,I881361,I881378,I881395,I881421,I881452,I881460,I881477,I881503,I881511,I881551,I881587,I881604,I881630,I881638,I881655,I881686,I881703,I881720,I881751,I881782,I881799,I881854,I881880,I881888,I881905,I881922,I881948,I881979,I881987,I882004,I882030,I882038,I882078,I882114,I882131,I882157,I882165,I882182,I882213,I882230,I882247,I882278,I882309,I882326,I882381,I1072260,I882407,I882415,I882432,I1072242,I882449,I1072248,I882475,I882370,I1072245,I882506,I882514,I1072254,I882531,I882557,I882565,I882373,I1072266,I882605,I882364,I882355,I882641,I1072257,I1072251,I882658,I882684,I882692,I882709,I882358,I882740,I1072263,I882757,I882774,I882367,I882805,I882352,I882836,I882853,I882361,I882908,I1277314,I882934,I882942,I882959,I1277296,I1277299,I882976,I1277311,I883002,I882897,I1277320,I883033,I883041,I1277305,I883058,I883084,I883092,I882900,I1277317,I883132,I882891,I882882,I883168,I1277308,I1277302,I883185,I883211,I883219,I883236,I882885,I883267,I883284,I883301,I882894,I883332,I882879,I883363,I883380,I882888,I883435,I1331507,I883461,I883469,I883486,I1331504,I1331513,I883503,I1331492,I883529,I883424,I1331495,I883560,I883568,I1331510,I883585,I883611,I883619,I883427,I1331516,I883659,I883418,I883409,I883695,I1331498,I1331519,I883712,I1331501,I883738,I883746,I883763,I883412,I883794,I883811,I883828,I883421,I883859,I883406,I883890,I883907,I883415,I883962,I883988,I883996,I884013,I884030,I884056,I884087,I884095,I884112,I884138,I884146,I884186,I884222,I884239,I884265,I884273,I884290,I884321,I884338,I884355,I884386,I884417,I884434,I884489,I884515,I884523,I884540,I884557,I884583,I884614,I884622,I884639,I884665,I884673,I884713,I884749,I884766,I884792,I884800,I884817,I884848,I884865,I884882,I884913,I884944,I884961,I885022,I885048,I885065,I885073,I885090,I885107,I885124,I885141,I885158,I885189,I885206,I885237,I885254,I885271,I885302,I885342,I885350,I885367,I885384,I885401,I885432,I885449,I885466,I885492,I885514,I885531,I885562,I885607,I885668,I885694,I885711,I885719,I885736,I885753,I885770,I885787,I885804,I885835,I885852,I885883,I885900,I885917,I885948,I885988,I885996,I886013,I886030,I886047,I886078,I886095,I886112,I886138,I886160,I886177,I886208,I886253,I886314,I886340,I886357,I886365,I886382,I886399,I886416,I886433,I886450,I886481,I886498,I886529,I886546,I886563,I886594,I886634,I886642,I886659,I886676,I886693,I886724,I886741,I886758,I886784,I886806,I886823,I886854,I886899,I886960,I886986,I887003,I887011,I887028,I887045,I887062,I887079,I887096,I887127,I887144,I887175,I887192,I887209,I887240,I887280,I887288,I887305,I887322,I887339,I887370,I887387,I887404,I887430,I887452,I887469,I887500,I887545,I887606,I1357672,I887632,I1357696,I887649,I887657,I887674,I1357678,I887691,I1357687,I887708,I887725,I1357693,I887742,I887592,I887773,I887790,I887595,I887821,I887838,I1357690,I887855,I887571,I887886,I887583,I887926,I887934,I887951,I887968,I1357684,I887985,I887598,I888016,I1357675,I888033,I1357699,I888050,I1357681,I888076,I887586,I888098,I888115,I887580,I888146,I887574,I887577,I888191,I887589,I888252,I888278,I888295,I888303,I888320,I888337,I888354,I888371,I888388,I888238,I888419,I888436,I888241,I888467,I888484,I888501,I888217,I888532,I888229,I888572,I888580,I888597,I888614,I888631,I888244,I888662,I888679,I888696,I888722,I888232,I888744,I888761,I888226,I888792,I888220,I888223,I888837,I888235,I888898,I888924,I888941,I888949,I888966,I888983,I889000,I889017,I889034,I889065,I889082,I889113,I889130,I889147,I889178,I889218,I889226,I889243,I889260,I889277,I889308,I889325,I889342,I889368,I889390,I889407,I889438,I889483,I889544,I889570,I889587,I889595,I889612,I889629,I889646,I889663,I889680,I889530,I889711,I889728,I889533,I889759,I889776,I889793,I889509,I889824,I889521,I889864,I889872,I889889,I889906,I889923,I889536,I889954,I889971,I889988,I890014,I889524,I890036,I890053,I889518,I890084,I889512,I889515,I890129,I889527,I890190,I1133528,I890216,I1133510,I890233,I890241,I890258,I1133519,I890275,I1133531,I890292,I1133513,I890309,I1133522,I890326,I890357,I890374,I890405,I890422,I1133534,I890439,I890470,I890510,I890518,I890535,I890552,I890569,I890600,I1133516,I890617,I1133525,I890634,I890660,I890682,I890699,I890730,I890775,I890836,I890862,I890879,I890887,I890904,I890921,I890938,I890955,I890972,I891003,I891020,I891051,I891068,I891085,I891116,I891156,I891164,I891181,I891198,I891215,I891246,I891263,I891280,I891306,I891328,I891345,I891376,I891421,I891482,I891508,I891525,I891533,I891550,I891567,I891584,I891601,I891618,I891649,I891666,I891697,I891714,I891731,I891762,I891802,I891810,I891827,I891844,I891861,I891892,I891909,I891926,I891952,I891974,I891991,I892022,I892067,I892128,I892154,I892171,I892179,I892196,I892213,I892230,I892247,I892264,I892295,I892312,I892343,I892360,I892377,I892408,I892448,I892456,I892473,I892490,I892507,I892538,I892555,I892572,I892598,I892620,I892637,I892668,I892713,I892774,I892800,I892817,I892825,I892842,I892859,I892876,I892893,I892910,I892760,I892941,I892958,I892763,I892989,I893006,I893023,I892739,I893054,I892751,I893094,I893102,I893119,I893136,I893153,I892766,I893184,I893201,I893218,I893244,I892754,I893266,I893283,I892748,I893314,I892742,I892745,I893359,I892757,I893420,I893446,I893463,I893471,I893488,I893505,I893522,I893539,I893556,I893406,I893587,I893604,I893409,I893635,I893652,I893669,I893385,I893700,I893397,I893740,I893748,I893765,I893782,I893799,I893412,I893830,I893847,I893864,I893890,I893400,I893912,I893929,I893394,I893960,I893388,I893391,I894005,I893403,I894066,I894092,I894109,I894117,I894134,I894151,I894168,I894185,I894202,I894233,I894250,I894281,I894298,I894315,I894346,I894386,I894394,I894411,I894428,I894445,I894476,I894493,I894510,I894536,I894558,I894575,I894606,I894651,I894712,I1185548,I894738,I1185530,I894755,I894763,I894780,I1185539,I894797,I1185551,I894814,I1185533,I894831,I1185542,I894848,I894879,I894896,I894927,I894944,I1185554,I894961,I894992,I895032,I895040,I895057,I895074,I895091,I895122,I1185536,I895139,I1185545,I895156,I895182,I895204,I895221,I895252,I895297,I895358,I1033703,I895384,I1033706,I895401,I895409,I895426,I895443,I1033715,I895460,I1033724,I895477,I1033712,I895494,I895344,I895525,I895542,I895347,I895573,I895590,I1033718,I895607,I895323,I895638,I895335,I895678,I895686,I895703,I895720,I1033709,I895737,I895350,I895768,I1033721,I895785,I895802,I895828,I895338,I895850,I895867,I895332,I895898,I895326,I895329,I895943,I895341,I896004,I896030,I896047,I896055,I896072,I896089,I896106,I896123,I896140,I896171,I896188,I896219,I896236,I896253,I896284,I896324,I896332,I896349,I896366,I896383,I896414,I896431,I896448,I896474,I896496,I896513,I896544,I896589,I896650,I896676,I896693,I896701,I896718,I896735,I896752,I896769,I896786,I896636,I896817,I896834,I896639,I896865,I896882,I896899,I896615,I896930,I896627,I896970,I896978,I896995,I897012,I897029,I896642,I897060,I897077,I897094,I897120,I896630,I897142,I897159,I896624,I897190,I896618,I896621,I897235,I896633,I897296,I897322,I897339,I897347,I897364,I897381,I897398,I897415,I897432,I897463,I897480,I897511,I897528,I897545,I897576,I897616,I897624,I897641,I897658,I897675,I897706,I897723,I897740,I897766,I897788,I897805,I897836,I897881,I897942,I897968,I897985,I897993,I898010,I898027,I898044,I898061,I898078,I898109,I898126,I898157,I898174,I898191,I898222,I898262,I898270,I898287,I898304,I898321,I898352,I898369,I898386,I898412,I898434,I898451,I898482,I898527,I898588,I1173988,I898614,I1173970,I898631,I898639,I898656,I1173979,I898673,I1173991,I898690,I1173973,I898707,I1173982,I898724,I898755,I898772,I898803,I898820,I1173994,I898837,I898868,I898908,I898916,I898933,I898950,I898967,I898998,I1173976,I899015,I1173985,I899032,I899058,I899080,I899097,I899128,I899173,I899234,I899260,I899277,I899285,I899302,I899319,I899336,I899353,I899370,I899401,I899418,I899449,I899466,I899483,I899514,I899554,I899562,I899579,I899596,I899613,I899644,I899661,I899678,I899704,I899726,I899743,I899774,I899819,I899880,I899906,I899923,I899931,I899948,I899965,I899982,I899999,I900016,I900047,I900064,I900095,I900112,I900129,I900160,I900200,I900208,I900225,I900242,I900259,I900290,I900307,I900324,I900350,I900372,I900389,I900420,I900465,I900526,I1220500,I900552,I1220506,I900569,I900577,I900594,I1220503,I900611,I1220482,I900628,I1220485,I900645,I1220491,I900662,I900512,I900693,I900710,I900515,I900741,I900758,I900775,I900491,I900806,I900503,I900846,I900854,I900871,I900888,I1220494,I900905,I900518,I900936,I900953,I1220488,I900970,I1220497,I900996,I900506,I901018,I901035,I900500,I901066,I900494,I900497,I901111,I900509,I901172,I901198,I901215,I901223,I901240,I901257,I901274,I901291,I901308,I901339,I901356,I901387,I901404,I901421,I901452,I901492,I901500,I901517,I901534,I901551,I901582,I901599,I901616,I901642,I901664,I901681,I901712,I901757,I901818,I901844,I901861,I901869,I901886,I901903,I901920,I901937,I901954,I901985,I902002,I902033,I902050,I902067,I902098,I902138,I902146,I902163,I902180,I902197,I902228,I902245,I902262,I902288,I902310,I902327,I902358,I902403,I902464,I902490,I902507,I902515,I902532,I902549,I902566,I902583,I902600,I902450,I902631,I902648,I902453,I902679,I902696,I902713,I902429,I902744,I902441,I902784,I902792,I902809,I902826,I902843,I902456,I902874,I902891,I902908,I902934,I902444,I902956,I902973,I902438,I903004,I902432,I902435,I903049,I902447,I903110,I903136,I903153,I903161,I903178,I903195,I903212,I903229,I903246,I903277,I903294,I903325,I903342,I903359,I903390,I903430,I903438,I903455,I903472,I903489,I903520,I903537,I903554,I903580,I903602,I903619,I903650,I903695,I903756,I1171676,I903782,I1171658,I903799,I903807,I903824,I1171667,I903841,I1171679,I903858,I1171661,I903875,I1171670,I903892,I903923,I903940,I903971,I903988,I1171682,I904005,I904036,I904076,I904084,I904101,I904118,I904135,I904166,I1171664,I904183,I1171673,I904200,I904226,I904248,I904265,I904296,I904341,I904402,I904428,I904445,I904453,I904470,I904487,I904504,I904521,I904538,I904569,I904586,I904617,I904634,I904651,I904682,I904722,I904730,I904747,I904764,I904781,I904812,I904829,I904846,I904872,I904894,I904911,I904942,I904987,I905048,I905074,I905091,I905099,I905116,I905133,I905150,I905167,I905184,I905215,I905232,I905263,I905280,I905297,I905328,I905368,I905376,I905393,I905410,I905427,I905458,I905475,I905492,I905518,I905540,I905557,I905588,I905633,I905694,I905720,I905737,I905745,I905762,I905779,I905796,I905813,I905830,I905861,I905878,I905909,I905926,I905943,I905974,I906014,I906022,I906039,I906056,I906073,I906104,I906121,I906138,I906164,I906186,I906203,I906234,I906279,I906340,I1102316,I906366,I1102298,I906383,I906391,I906408,I1102307,I906425,I1102319,I906442,I1102301,I906459,I1102310,I906476,I906326,I906507,I906524,I906329,I906555,I906572,I1102322,I906589,I906305,I906620,I906317,I906660,I906668,I906685,I906702,I906719,I906332,I906750,I1102304,I906767,I1102313,I906784,I906810,I906320,I906832,I906849,I906314,I906880,I906308,I906311,I906925,I906323,I906986,I907012,I907029,I907037,I907054,I907071,I907088,I907105,I907122,I907153,I907170,I907201,I907218,I907235,I907266,I907306,I907314,I907331,I907348,I907365,I907396,I907413,I907430,I907456,I907478,I907495,I907526,I907571,I907632,I907658,I907675,I907683,I907700,I907717,I907734,I907751,I907768,I907799,I907816,I907847,I907864,I907881,I907912,I907952,I907960,I907977,I907994,I908011,I908042,I908059,I908076,I908102,I908124,I908141,I908172,I908217,I908278,I1066480,I908304,I1066462,I908321,I908329,I908346,I1066471,I908363,I1066483,I908380,I1066465,I908397,I1066474,I908414,I908264,I908445,I908462,I908267,I908493,I908510,I1066486,I908527,I908243,I908558,I908255,I908598,I908606,I908623,I908640,I908657,I908270,I908688,I1066468,I908705,I1066477,I908722,I908748,I908258,I908770,I908787,I908252,I908818,I908246,I908249,I908863,I908261,I908924,I908950,I908967,I908975,I908992,I909009,I909026,I909043,I909060,I909091,I909108,I909139,I909156,I909173,I909204,I909244,I909252,I909269,I909286,I909303,I909334,I909351,I909368,I909394,I909416,I909433,I909464,I909509,I909570,I1318997,I909596,I1319021,I909613,I909621,I909638,I1319003,I909655,I1319012,I909672,I909689,I1319018,I909706,I909737,I909754,I909785,I909802,I1319015,I909819,I909850,I909890,I909898,I909915,I909932,I1319009,I909949,I909980,I1319000,I909997,I1319024,I910014,I1319006,I910040,I910062,I910079,I910110,I910155,I910216,I1023044,I910242,I1023047,I910259,I910267,I910284,I910301,I1023056,I910318,I1023065,I910335,I1023053,I910352,I910383,I910400,I910431,I910448,I1023059,I910465,I910496,I910536,I910544,I910561,I910578,I1023050,I910595,I910626,I1023062,I910643,I910660,I910686,I910708,I910725,I910756,I910801,I910862,I910888,I910905,I910913,I910930,I910947,I910964,I910981,I910998,I911029,I911046,I911077,I911094,I911111,I911142,I911182,I911190,I911207,I911224,I911241,I911272,I911289,I911306,I911332,I911354,I911371,I911402,I911447,I911508,I911534,I911551,I911559,I911576,I911593,I911610,I911627,I911644,I911675,I911692,I911723,I911740,I911757,I911788,I911828,I911836,I911853,I911870,I911887,I911918,I911935,I911952,I911978,I912000,I912017,I912048,I912093,I912154,I912180,I912197,I912205,I912222,I912239,I912256,I912273,I912290,I912321,I912338,I912369,I912386,I912403,I912434,I912474,I912482,I912499,I912516,I912533,I912564,I912581,I912598,I912624,I912646,I912663,I912694,I912739,I912800,I912826,I912843,I912851,I912868,I912885,I912902,I912919,I912936,I912967,I912984,I913015,I913032,I913049,I913080,I913120,I913128,I913145,I913162,I913179,I913210,I913227,I913244,I913270,I913292,I913309,I913340,I913385,I913446,I913472,I913489,I913497,I913514,I913531,I913548,I913565,I913582,I913613,I913630,I913661,I913678,I913695,I913726,I913766,I913774,I913791,I913808,I913825,I913856,I913873,I913890,I913916,I913938,I913955,I913986,I914031,I914092,I914118,I914135,I914143,I914160,I914177,I914194,I914211,I914228,I914259,I914276,I914307,I914324,I914341,I914372,I914412,I914420,I914437,I914454,I914471,I914502,I914519,I914536,I914562,I914584,I914601,I914632,I914677,I914738,I914764,I914781,I914789,I914806,I914823,I914840,I914857,I914874,I914905,I914922,I914953,I914970,I914987,I915018,I915058,I915066,I915083,I915100,I915117,I915148,I915165,I915182,I915208,I915230,I915247,I915278,I915323,I915384,I915410,I915427,I915435,I915452,I915469,I915486,I915503,I915520,I915551,I915568,I915599,I915616,I915633,I915664,I915704,I915712,I915729,I915746,I915763,I915794,I915811,I915828,I915854,I915876,I915893,I915924,I915969,I916030,I916056,I916073,I916081,I916098,I916115,I916132,I916149,I916166,I916197,I916214,I916245,I916262,I916279,I916310,I916350,I916358,I916375,I916392,I916409,I916440,I916457,I916474,I916500,I916522,I916539,I916570,I916615,I916676,I916702,I916719,I916727,I916744,I916761,I916778,I916795,I916812,I916843,I916860,I916891,I916908,I916925,I916956,I916996,I917004,I917021,I917038,I917055,I917086,I917103,I917120,I917146,I917168,I917185,I917216,I917261,I917322,I917348,I917365,I917373,I917390,I917407,I917424,I917441,I917458,I917489,I917506,I917537,I917554,I917571,I917602,I917642,I917650,I917667,I917684,I917701,I917732,I917749,I917766,I917792,I917814,I917831,I917862,I917907,I917968,I917994,I918011,I918019,I918036,I918053,I918070,I918087,I918104,I917954,I918135,I918152,I917957,I918183,I918200,I918217,I917933,I918248,I917945,I918288,I918296,I918313,I918330,I918347,I917960,I918378,I918395,I918412,I918438,I917948,I918460,I918477,I917942,I918508,I917936,I917939,I918553,I917951,I918614,I918640,I918657,I918665,I918682,I918699,I918716,I918733,I918750,I918600,I918781,I918798,I918603,I918829,I918846,I918863,I918579,I918894,I918591,I918934,I918942,I918959,I918976,I918993,I918606,I919024,I919041,I919058,I919084,I918594,I919106,I919123,I918588,I919154,I918582,I918585,I919199,I918597,I919260,I1081508,I919286,I1081490,I919303,I919311,I919328,I1081499,I919345,I1081511,I919362,I1081493,I919379,I1081502,I919396,I919427,I919444,I919475,I919492,I1081514,I919509,I919540,I919580,I919588,I919605,I919622,I919639,I919670,I1081496,I919687,I1081505,I919704,I919730,I919752,I919769,I919800,I919845,I919906,I919932,I919949,I919957,I919974,I919991,I920008,I920025,I920042,I920073,I920090,I920121,I920138,I920155,I920186,I920226,I920234,I920251,I920268,I920285,I920316,I920333,I920350,I920376,I920398,I920415,I920446,I920491,I920552,I920578,I920595,I920603,I920620,I920637,I920654,I920671,I920688,I920719,I920736,I920767,I920784,I920801,I920832,I920872,I920880,I920897,I920914,I920931,I920962,I920979,I920996,I921022,I921044,I921061,I921092,I921137,I921198,I921224,I921241,I921249,I921266,I921283,I921300,I921317,I921334,I921365,I921382,I921413,I921430,I921447,I921478,I921518,I921526,I921543,I921560,I921577,I921608,I921625,I921642,I921668,I921690,I921707,I921738,I921783,I921844,I921870,I921887,I921895,I921912,I921929,I921946,I921963,I921980,I922011,I922028,I922059,I922076,I922093,I922124,I922164,I922172,I922189,I922206,I922223,I922254,I922271,I922288,I922314,I922336,I922353,I922384,I922429,I922490,I1115610,I922516,I1115592,I922533,I922541,I922558,I1115601,I922575,I1115613,I922592,I1115595,I922609,I1115604,I922626,I922657,I922674,I922705,I922722,I1115616,I922739,I922770,I922810,I922818,I922835,I922852,I922869,I922900,I1115598,I922917,I1115607,I922934,I922960,I922982,I922999,I923030,I923075,I923136,I1146244,I923162,I1146226,I923179,I923187,I923204,I1146235,I923221,I1146247,I923238,I1146229,I923255,I1146238,I923272,I923303,I923320,I923351,I923368,I1146250,I923385,I923416,I923456,I923464,I923481,I923498,I923515,I923546,I1146232,I923563,I1146241,I923580,I923606,I923628,I923645,I923676,I923721,I923782,I923808,I923825,I923833,I923850,I923867,I923884,I923901,I923918,I923949,I923966,I923997,I924014,I924031,I924062,I924102,I924110,I924127,I924144,I924161,I924192,I924209,I924226,I924252,I924274,I924291,I924322,I924367,I924428,I924454,I924471,I924479,I924496,I924513,I924530,I924547,I924564,I924414,I924595,I924612,I924417,I924643,I924660,I924677,I924393,I924708,I924405,I924748,I924756,I924773,I924790,I924807,I924420,I924838,I924855,I924872,I924898,I924408,I924920,I924937,I924402,I924968,I924396,I924399,I925013,I924411,I925074,I925100,I925117,I925125,I925142,I925159,I925176,I925193,I925210,I925241,I925258,I925289,I925306,I925323,I925354,I925394,I925402,I925419,I925436,I925453,I925484,I925501,I925518,I925544,I925566,I925583,I925614,I925659,I925720,I925746,I925763,I925771,I925788,I925805,I925822,I925839,I925856,I925887,I925904,I925935,I925952,I925969,I926000,I926040,I926048,I926065,I926082,I926099,I926130,I926147,I926164,I926190,I926212,I926229,I926260,I926305,I926366,I926392,I926409,I926417,I926434,I926451,I926468,I926485,I926502,I926533,I926550,I926581,I926598,I926615,I926646,I926686,I926694,I926711,I926728,I926745,I926776,I926793,I926810,I926836,I926858,I926875,I926906,I926951,I927012,I1317212,I927038,I1317236,I927055,I927063,I927080,I1317218,I927097,I1317227,I927114,I927131,I1317233,I927148,I926998,I927179,I927196,I927001,I927227,I927244,I1317230,I927261,I926977,I927292,I926989,I927332,I927340,I927357,I927374,I1317224,I927391,I927004,I927422,I1317215,I927439,I1317239,I927456,I1317221,I927482,I926992,I927504,I927521,I926986,I927552,I926980,I926983,I927597,I926995,I927658,I1219956,I927684,I1219962,I927701,I927709,I927726,I1219959,I927743,I1219938,I927760,I1219941,I927777,I1219947,I927794,I927644,I927825,I927842,I927647,I927873,I927890,I927907,I927623,I927938,I927635,I927978,I927986,I928003,I928020,I1219950,I928037,I927650,I928068,I928085,I1219944,I928102,I1219953,I928128,I927638,I928150,I928167,I927632,I928198,I927626,I927629,I928243,I927641,I928304,I928330,I928347,I928355,I928372,I928389,I928406,I928423,I928440,I928290,I928471,I928488,I928293,I928519,I928536,I928553,I928269,I928584,I928281,I928624,I928632,I928649,I928666,I928683,I928296,I928714,I928731,I928748,I928774,I928284,I928796,I928813,I928278,I928844,I928272,I928275,I928889,I928287,I928950,I1294645,I928976,I1294639,I928993,I929001,I929018,I1294648,I929035,I1294660,I929052,I1294642,I929069,I929086,I929117,I929134,I929165,I929182,I1294636,I929199,I929230,I929270,I929278,I929295,I929312,I1294657,I929329,I929360,I1294651,I929377,I929394,I1294654,I929420,I929442,I929459,I929490,I929535,I929596,I929622,I929639,I929647,I929664,I929681,I929698,I929715,I929732,I929763,I929780,I929811,I929828,I929845,I929876,I929916,I929924,I929941,I929958,I929975,I930006,I930023,I930040,I930066,I930088,I930105,I930136,I930181,I930242,I930268,I930285,I930293,I930310,I930327,I930344,I930361,I930378,I930228,I930409,I930426,I930231,I930457,I930474,I930491,I930207,I930522,I930219,I930562,I930570,I930587,I930604,I930621,I930234,I930652,I930669,I930686,I930712,I930222,I930734,I930751,I930216,I930782,I930210,I930213,I930827,I930225,I930888,I930914,I930931,I930939,I930956,I930973,I930990,I931007,I931024,I930874,I931055,I931072,I930877,I931103,I931120,I931137,I930853,I931168,I930865,I931208,I931216,I931233,I931250,I931267,I930880,I931298,I931315,I931332,I931358,I930868,I931380,I931397,I930862,I931428,I930856,I930859,I931473,I930871,I931534,I931560,I931577,I931585,I931602,I931619,I931636,I931653,I931670,I931701,I931718,I931749,I931766,I931783,I931814,I931854,I931862,I931879,I931896,I931913,I931944,I931961,I931978,I932004,I932026,I932043,I932074,I932119,I932180,I1139308,I932206,I1139290,I932223,I932231,I932248,I1139299,I932265,I1139311,I932282,I1139293,I932299,I1139302,I932316,I932347,I932364,I932395,I932412,I1139314,I932429,I932460,I932500,I932508,I932525,I932542,I932559,I932590,I1139296,I932607,I1139305,I932624,I932650,I932672,I932689,I932720,I932765,I932826,I932852,I932869,I932877,I932894,I932911,I932928,I932945,I932962,I932812,I932993,I933010,I932815,I933041,I933058,I933075,I932791,I933106,I932803,I933146,I933154,I933171,I933188,I933205,I932818,I933236,I933253,I933270,I933296,I932806,I933318,I933335,I932800,I933366,I932794,I932797,I933411,I932809,I933472,I933498,I933515,I933523,I933540,I933557,I933574,I933591,I933608,I933639,I933656,I933687,I933704,I933721,I933752,I933792,I933800,I933817,I933834,I933851,I933882,I933899,I933916,I933942,I933964,I933981,I934012,I934057,I934118,I1316617,I934144,I1316641,I934161,I934169,I934186,I1316623,I934203,I1316632,I934220,I934237,I1316638,I934254,I934285,I934302,I934333,I934350,I1316635,I934367,I934398,I934438,I934446,I934463,I934480,I1316629,I934497,I934528,I1316620,I934545,I1316644,I934562,I1316626,I934588,I934610,I934627,I934658,I934703,I934764,I934790,I934807,I934815,I934832,I934849,I934866,I934883,I934900,I934931,I934948,I934979,I934996,I935013,I935044,I935084,I935092,I935109,I935126,I935143,I935174,I935191,I935208,I935234,I935256,I935273,I935304,I935349,I935410,I935436,I935453,I935461,I935478,I935495,I935512,I935529,I935546,I935577,I935594,I935625,I935642,I935659,I935690,I935730,I935738,I935755,I935772,I935789,I935820,I935837,I935854,I935880,I935902,I935919,I935950,I935995,I936056,I936082,I936099,I936107,I936124,I936141,I936158,I936175,I936192,I936223,I936240,I936271,I936288,I936305,I936336,I936376,I936384,I936401,I936418,I936435,I936466,I936483,I936500,I936526,I936548,I936565,I936596,I936641,I936702,I936728,I936745,I936753,I936770,I936787,I936804,I936821,I936838,I936869,I936886,I936917,I936934,I936951,I936982,I937022,I937030,I937047,I937064,I937081,I937112,I937129,I937146,I937172,I937194,I937211,I937242,I937287,I937348,I1214516,I937374,I1214522,I937391,I937399,I937416,I1214519,I937433,I1214498,I937450,I1214501,I937467,I1214507,I937484,I937515,I937532,I937563,I937580,I937597,I937628,I937668,I937676,I937693,I937710,I1214510,I937727,I937758,I937775,I1214504,I937792,I1214513,I937818,I937840,I937857,I937888,I937933,I937994,I938020,I938037,I938045,I938062,I938079,I938096,I938113,I938130,I938161,I938178,I938209,I938226,I938243,I938274,I938314,I938322,I938339,I938356,I938373,I938404,I938421,I938438,I938464,I938486,I938503,I938534,I938579,I938640,I938666,I938683,I938691,I938708,I938725,I938742,I938759,I938776,I938807,I938824,I938855,I938872,I938889,I938920,I938960,I938968,I938985,I939002,I939019,I939050,I939067,I939084,I939110,I939132,I939149,I939180,I939225,I939286,I939312,I939329,I939337,I939354,I939371,I939388,I939405,I939422,I939453,I939470,I939501,I939518,I939535,I939566,I939606,I939614,I939631,I939648,I939665,I939696,I939713,I939730,I939756,I939778,I939795,I939826,I939871,I939932,I939958,I939975,I939983,I940000,I940017,I940034,I940051,I940068,I940099,I940116,I940147,I940164,I940181,I940212,I940252,I940260,I940277,I940294,I940311,I940342,I940359,I940376,I940402,I940424,I940441,I940472,I940517,I940578,I1368977,I940604,I1369001,I940621,I940629,I940646,I1368983,I940663,I1368992,I940680,I940697,I1368998,I940714,I940745,I940762,I940793,I940810,I1368995,I940827,I940858,I940898,I940906,I940923,I940940,I1368989,I940957,I940988,I1368980,I941005,I1369004,I941022,I1368986,I941048,I941070,I941087,I941118,I941163,I941224,I941250,I941267,I941275,I941292,I941309,I941326,I941343,I941360,I941391,I941408,I941439,I941456,I941473,I941504,I941544,I941552,I941569,I941586,I941603,I941634,I941651,I941668,I941694,I941716,I941733,I941764,I941809,I941870,I941896,I941913,I941921,I941938,I941955,I941972,I941989,I942006,I942037,I942054,I942085,I942102,I942119,I942150,I942190,I942198,I942215,I942232,I942249,I942280,I942297,I942314,I942340,I942362,I942379,I942410,I942455,I942516,I942542,I942559,I942567,I942584,I942601,I942618,I942635,I942652,I942502,I942683,I942700,I942505,I942731,I942748,I942765,I942481,I942796,I942493,I942836,I942844,I942861,I942878,I942895,I942508,I942926,I942943,I942960,I942986,I942496,I943008,I943025,I942490,I943056,I942484,I942487,I943101,I942499,I943162,I943188,I943205,I943213,I943230,I943247,I943264,I943281,I943298,I943329,I943346,I943377,I943394,I943411,I943442,I943482,I943490,I943507,I943524,I943541,I943572,I943589,I943606,I943632,I943654,I943671,I943702,I943747,I943808,I943834,I943851,I943859,I943876,I943893,I943910,I943927,I943944,I943975,I943992,I944023,I944040,I944057,I944088,I944128,I944136,I944153,I944170,I944187,I944218,I944235,I944252,I944278,I944300,I944317,I944348,I944393,I944454,I944480,I944497,I944505,I944522,I944539,I944556,I944573,I944590,I944621,I944638,I944669,I944686,I944703,I944734,I944774,I944782,I944799,I944816,I944833,I944864,I944881,I944898,I944924,I944946,I944963,I944994,I945039,I945100,I945126,I945143,I945151,I945168,I945185,I945202,I945219,I945236,I945086,I945267,I945284,I945089,I945315,I945332,I945349,I945065,I945380,I945077,I945420,I945428,I945445,I945462,I945479,I945092,I945510,I945527,I945544,I945570,I945080,I945592,I945609,I945074,I945640,I945068,I945071,I945685,I945083,I945746,I945772,I945789,I945797,I945814,I945831,I945848,I945865,I945882,I945913,I945930,I945961,I945978,I945995,I946026,I946066,I946074,I946091,I946108,I946125,I946156,I946173,I946190,I946216,I946238,I946255,I946286,I946331,I946392,I946418,I946435,I946443,I946460,I946477,I946494,I946511,I946528,I946559,I946576,I946607,I946624,I946641,I946672,I946712,I946720,I946737,I946754,I946771,I946802,I946819,I946836,I946862,I946884,I946901,I946932,I946977,I947038,I1276727,I947064,I1276721,I947081,I947089,I947106,I1276730,I947123,I1276742,I947140,I1276724,I947157,I947174,I947205,I947222,I947253,I947270,I1276718,I947287,I947318,I947358,I947366,I947383,I947400,I1276739,I947417,I947448,I1276733,I947465,I947482,I1276736,I947508,I947530,I947547,I947578,I947623,I947684,I947710,I947727,I947735,I947752,I947769,I947786,I947803,I947820,I947851,I947868,I947899,I947916,I947933,I947964,I948004,I948012,I948029,I948046,I948063,I948094,I948111,I948128,I948154,I948176,I948193,I948224,I948269,I948330,I948356,I948373,I948381,I948398,I948415,I948432,I948449,I948466,I948497,I948514,I948545,I948562,I948579,I948610,I948650,I948658,I948675,I948692,I948709,I948740,I948757,I948774,I948800,I948822,I948839,I948870,I948915,I948976,I949002,I949019,I949027,I949044,I949061,I949078,I949095,I949112,I949143,I949160,I949191,I949208,I949225,I949256,I949296,I949304,I949321,I949338,I949355,I949386,I949403,I949420,I949446,I949468,I949485,I949516,I949561,I949622,I1077462,I949648,I1077444,I949665,I949673,I949690,I1077453,I949707,I1077465,I949724,I1077447,I949741,I1077456,I949758,I949789,I949806,I949837,I949854,I1077468,I949871,I949902,I949942,I949950,I949967,I949984,I950001,I950032,I1077450,I950049,I1077459,I950066,I950092,I950114,I950131,I950162,I950207,I950268,I950294,I950311,I950319,I950336,I950353,I950370,I950387,I950404,I950435,I950452,I950483,I950500,I950517,I950548,I950588,I950596,I950613,I950630,I950647,I950678,I950695,I950712,I950738,I950760,I950777,I950808,I950853,I950914,I950940,I950957,I950965,I950982,I950999,I951016,I951033,I951050,I950900,I951081,I951098,I950903,I951129,I951146,I951163,I950879,I951194,I950891,I951234,I951242,I951259,I951276,I951293,I950906,I951324,I951341,I951358,I951384,I950894,I951406,I951423,I950888,I951454,I950882,I950885,I951499,I950897,I951560,I1042679,I951586,I1042682,I951603,I951611,I951628,I951645,I1042691,I951662,I1042700,I951679,I1042688,I951696,I951546,I951727,I951744,I951549,I951775,I951792,I1042694,I951809,I951525,I951840,I951537,I951880,I951888,I951905,I951922,I1042685,I951939,I951552,I951970,I1042697,I951987,I952004,I952030,I951540,I952052,I952069,I951534,I952100,I951528,I951531,I952145,I951543,I952206,I1333277,I952232,I1333301,I952249,I952257,I952274,I1333283,I952291,I1333292,I952308,I952325,I1333298,I952342,I952373,I952390,I952421,I952438,I1333295,I952455,I952486,I952526,I952534,I952551,I952568,I1333289,I952585,I952616,I1333280,I952633,I1333304,I952650,I1333286,I952676,I952698,I952715,I952746,I952791,I952852,I952878,I952895,I952903,I952920,I952937,I952954,I952971,I952988,I952838,I953019,I953036,I952841,I953067,I953084,I953101,I952817,I953132,I952829,I953172,I953180,I953197,I953214,I953231,I952844,I953262,I953279,I953296,I953322,I952832,I953344,I953361,I952826,I953392,I952820,I952823,I953437,I952835,I953498,I953524,I953541,I953549,I953566,I953583,I953600,I953617,I953634,I953665,I953682,I953713,I953730,I953747,I953778,I953818,I953826,I953843,I953860,I953877,I953908,I953925,I953942,I953968,I953990,I954007,I954038,I954083,I954144,I954170,I954187,I954195,I954212,I954229,I954246,I954263,I954280,I954130,I954311,I954328,I954133,I954359,I954376,I954393,I954109,I954424,I954121,I954464,I954472,I954489,I954506,I954523,I954136,I954554,I954571,I954588,I954614,I954124,I954636,I954653,I954118,I954684,I954112,I954115,I954729,I954127,I954790,I954816,I954833,I954841,I954858,I954875,I954892,I954909,I954926,I954957,I954974,I955005,I955022,I955039,I955070,I955110,I955118,I955135,I955152,I955169,I955200,I955217,I955234,I955260,I955282,I955299,I955330,I955375,I955436,I1323757,I955462,I1323781,I955479,I955487,I955504,I1323763,I955521,I1323772,I955538,I955555,I1323778,I955572,I955603,I955620,I955651,I955668,I1323775,I955685,I955716,I955756,I955764,I955781,I955798,I1323769,I955815,I955846,I1323760,I955863,I1323784,I955880,I1323766,I955906,I955928,I955945,I955976,I956021,I956082,I956108,I956125,I956133,I956150,I956167,I956184,I956201,I956218,I956249,I956266,I956297,I956314,I956331,I956362,I956402,I956410,I956427,I956444,I956461,I956492,I956509,I956526,I956552,I956574,I956591,I956622,I956667,I956728,I956754,I956771,I956779,I956796,I956813,I956830,I956847,I956864,I956895,I956912,I956943,I956960,I956977,I957008,I957048,I957056,I957073,I957090,I957107,I957138,I957155,I957172,I957198,I957220,I957237,I957268,I957313,I957374,I957400,I957417,I957425,I957442,I957459,I957476,I957493,I957510,I957541,I957558,I957589,I957606,I957623,I957654,I957694,I957702,I957719,I957736,I957753,I957784,I957801,I957818,I957844,I957866,I957883,I957914,I957959,I958020,I958046,I958063,I958071,I958088,I958105,I958122,I958139,I958156,I958187,I958204,I958235,I958252,I958269,I958300,I958340,I958348,I958365,I958382,I958399,I958430,I958447,I958464,I958490,I958512,I958529,I958560,I958605,I958666,I958692,I958709,I958717,I958734,I958751,I958768,I958785,I958802,I958833,I958850,I958881,I958898,I958915,I958946,I958986,I958994,I959011,I959028,I959045,I959076,I959093,I959110,I959136,I959158,I959175,I959206,I959251,I959312,I959338,I959355,I959363,I959380,I959397,I959414,I959431,I959448,I959479,I959496,I959527,I959544,I959561,I959592,I959632,I959640,I959657,I959674,I959691,I959722,I959739,I959756,I959782,I959804,I959821,I959852,I959897,I959958,I959984,I960001,I960009,I960026,I960043,I960060,I960077,I960094,I959944,I960125,I960142,I959947,I960173,I960190,I960207,I959923,I960238,I959935,I960278,I960286,I960303,I960320,I960337,I959950,I960368,I960385,I960402,I960428,I959938,I960450,I960467,I959932,I960498,I959926,I959929,I960543,I959941,I960604,I1376117,I960630,I1376141,I960647,I960655,I960672,I1376123,I960689,I1376132,I960706,I960723,I1376138,I960740,I960590,I960771,I960788,I960593,I960819,I960836,I1376135,I960853,I960569,I960884,I960581,I960924,I960932,I960949,I960966,I1376129,I960983,I960596,I961014,I1376120,I961031,I1376144,I961048,I1376126,I961074,I960584,I961096,I961113,I960578,I961144,I960572,I960575,I961189,I960587,I961250,I961276,I961293,I961301,I961318,I961335,I961352,I961369,I961386,I961417,I961434,I961465,I961482,I961499,I961530,I961570,I961578,I961595,I961612,I961629,I961660,I961677,I961694,I961720,I961742,I961759,I961790,I961835,I961896,I1338037,I961922,I1338061,I961939,I961947,I961964,I1338043,I961981,I1338052,I961998,I962015,I1338058,I962032,I961882,I962063,I962080,I961885,I962111,I962128,I1338055,I962145,I961861,I962176,I961873,I962216,I962224,I962241,I962258,I1338049,I962275,I961888,I962306,I1338040,I962323,I1338064,I962340,I1338046,I962366,I961876,I962388,I962405,I961870,I962436,I961864,I961867,I962481,I961879,I962542,I962568,I962585,I962593,I962610,I962627,I962644,I962661,I962678,I962709,I962726,I962757,I962774,I962791,I962822,I962862,I962870,I962887,I962904,I962921,I962952,I962969,I962986,I963012,I963034,I963051,I963082,I963127,I963188,I963214,I963231,I963239,I963256,I963273,I963290,I963307,I963324,I963355,I963372,I963403,I963420,I963437,I963468,I963508,I963516,I963533,I963550,I963567,I963598,I963615,I963632,I963658,I963680,I963697,I963728,I963773,I963834,I1305361,I963860,I1305358,I963877,I963885,I963902,I1305355,I963919,I1305346,I963936,I1305367,I963953,I963970,I964001,I964018,I964049,I964066,I1305370,I964083,I964114,I964154,I964162,I964179,I964196,I1305349,I964213,I964244,I1305352,I964261,I1305373,I964278,I1305364,I964304,I964326,I964343,I964374,I964419,I964480,I964506,I964523,I964531,I964548,I964565,I964582,I964599,I964616,I964647,I964664,I964695,I964712,I964729,I964760,I964800,I964808,I964825,I964842,I964859,I964890,I964907,I964924,I964950,I964972,I964989,I965020,I965065,I965126,I965152,I965169,I965177,I965194,I965211,I965228,I965245,I965262,I965293,I965310,I965341,I965358,I965375,I965406,I965446,I965454,I965471,I965488,I965505,I965536,I965553,I965570,I965596,I965618,I965635,I965666,I965711,I965772,I1221044,I965798,I1221050,I965815,I965823,I965840,I1221047,I965857,I1221026,I965874,I1221029,I965891,I1221035,I965908,I965939,I965956,I965987,I966004,I966021,I966052,I966092,I966100,I966117,I966134,I1221038,I966151,I966182,I966199,I1221032,I966216,I1221041,I966242,I966264,I966281,I966312,I966357,I966418,I966444,I966461,I966469,I966486,I966503,I966520,I966537,I966554,I966585,I966602,I966633,I966650,I966667,I966698,I966738,I966746,I966763,I966780,I966797,I966828,I966845,I966862,I966888,I966910,I966927,I966958,I967003,I967064,I967090,I967107,I967115,I967132,I967149,I967166,I967183,I967200,I967231,I967248,I967279,I967296,I967313,I967344,I967384,I967392,I967409,I967426,I967443,I967474,I967491,I967508,I967534,I967556,I967573,I967604,I967649,I967710,I967736,I967753,I967761,I967778,I967795,I967812,I967829,I967846,I967877,I967894,I967925,I967942,I967959,I967990,I968030,I968038,I968055,I968072,I968089,I968120,I968137,I968154,I968180,I968202,I968219,I968250,I968295,I968356,I1203466,I968382,I1203448,I968399,I968407,I968424,I1203457,I968441,I1203469,I968458,I1203451,I968475,I1203460,I968492,I968523,I968540,I968571,I968588,I1203472,I968605,I968636,I968676,I968684,I968701,I968718,I968735,I968766,I1203454,I968783,I1203463,I968800,I968826,I968848,I968865,I968896,I968941,I969002,I969028,I969045,I969053,I969070,I969087,I969104,I969121,I969138,I968988,I969169,I969186,I968991,I969217,I969234,I969251,I968967,I969282,I968979,I969322,I969330,I969347,I969364,I969381,I968994,I969412,I969429,I969446,I969472,I968982,I969494,I969511,I968976,I969542,I968970,I968973,I969587,I968985,I969648,I969674,I969691,I969699,I969716,I969733,I969750,I969767,I969784,I969634,I969815,I969832,I969637,I969863,I969880,I969897,I969613,I969928,I969625,I969968,I969976,I969993,I970010,I970027,I969640,I970058,I970075,I970092,I970118,I969628,I970140,I970157,I969622,I970188,I969616,I969619,I970233,I969631,I970294,I970320,I970337,I970345,I970362,I970379,I970396,I970413,I970430,I970461,I970478,I970509,I970526,I970543,I970574,I970614,I970622,I970639,I970656,I970673,I970704,I970721,I970738,I970764,I970786,I970803,I970834,I970879,I970940,I970966,I970983,I970991,I971008,I971025,I971042,I971059,I971076,I970926,I971107,I971124,I970929,I971155,I971172,I971189,I970905,I971220,I970917,I971260,I971268,I971285,I971302,I971319,I970932,I971350,I971367,I971384,I971410,I970920,I971432,I971449,I970914,I971480,I970908,I970911,I971525,I970923,I971586,I971612,I971629,I971637,I971654,I971671,I971688,I971705,I971722,I971572,I971753,I971770,I971575,I971801,I971818,I971835,I971551,I971866,I971563,I971906,I971914,I971931,I971948,I971965,I971578,I971996,I972013,I972030,I972056,I971566,I972078,I972095,I971560,I972126,I971554,I971557,I972171,I971569,I972232,I972258,I972275,I972283,I972300,I972317,I972334,I972351,I972368,I972399,I972416,I972447,I972464,I972481,I972512,I972552,I972560,I972577,I972594,I972611,I972642,I972659,I972676,I972702,I972724,I972741,I972772,I972817,I972878,I972904,I972921,I972929,I972946,I972963,I972980,I972997,I973014,I973045,I973062,I973093,I973110,I973127,I973158,I973198,I973206,I973223,I973240,I973257,I973288,I973305,I973322,I973348,I973370,I973387,I973418,I973463,I973524,I1026410,I973550,I1026413,I973567,I973575,I973592,I973609,I1026422,I973626,I1026431,I973643,I1026419,I973660,I973691,I973708,I973739,I973756,I1026425,I973773,I973804,I973844,I973852,I973869,I973886,I1026416,I973903,I973934,I1026428,I973951,I973968,I973994,I974016,I974033,I974064,I974109,I974170,I974196,I974213,I974221,I974238,I974255,I974272,I974289,I974306,I974337,I974354,I974385,I974402,I974419,I974450,I974490,I974498,I974515,I974532,I974549,I974580,I974597,I974614,I974640,I974662,I974679,I974710,I974755,I974816,I974842,I974859,I974867,I974884,I974901,I974918,I974935,I974952,I974802,I974983,I975000,I974805,I975031,I975048,I975065,I974781,I975096,I974793,I975136,I975144,I975161,I975178,I975195,I974808,I975226,I975243,I975260,I975286,I974796,I975308,I975325,I974790,I975356,I974784,I974787,I975401,I974799,I975462,I975488,I975505,I975513,I975530,I975547,I975564,I975581,I975598,I975629,I975646,I975677,I975694,I975711,I975742,I975782,I975790,I975807,I975824,I975841,I975872,I975889,I975906,I975932,I975954,I975971,I976002,I976047,I976108,I976134,I976151,I976159,I976176,I976193,I976210,I976227,I976244,I976275,I976292,I976323,I976340,I976357,I976388,I976428,I976436,I976453,I976470,I976487,I976518,I976535,I976552,I976578,I976600,I976617,I976648,I976693,I976754,I976780,I976797,I976805,I976822,I976839,I976856,I976873,I976890,I976921,I976938,I976969,I976986,I977003,I977034,I977074,I977082,I977099,I977116,I977133,I977164,I977181,I977198,I977224,I977246,I977263,I977294,I977339,I977400,I977426,I977443,I977451,I977468,I977485,I977502,I977519,I977536,I977567,I977584,I977615,I977632,I977649,I977680,I977720,I977728,I977745,I977762,I977779,I977810,I977827,I977844,I977870,I977892,I977909,I977940,I977985,I978046,I978072,I978089,I978097,I978114,I978131,I978148,I978165,I978182,I978213,I978230,I978261,I978278,I978295,I978326,I978366,I978374,I978391,I978408,I978425,I978456,I978473,I978490,I978516,I978538,I978555,I978586,I978631,I978692,I1156648,I978718,I1156630,I978735,I978743,I978760,I1156639,I978777,I1156651,I978794,I1156633,I978811,I1156642,I978828,I978859,I978876,I978907,I978924,I1156654,I978941,I978972,I979012,I979020,I979037,I979054,I979071,I979102,I1156636,I979119,I1156645,I979136,I979162,I979184,I979201,I979232,I979277,I979338,I979364,I979381,I979389,I979406,I979423,I979440,I979457,I979474,I979324,I979505,I979522,I979327,I979553,I979570,I979587,I979303,I979618,I979315,I979658,I979666,I979683,I979700,I979717,I979330,I979748,I979765,I979782,I979808,I979318,I979830,I979847,I979312,I979878,I979306,I979309,I979923,I979321,I979984,I1388017,I980010,I1388041,I980027,I980035,I980052,I1388023,I980069,I1388032,I980086,I980103,I1388038,I980120,I979970,I980151,I980168,I979973,I980199,I980216,I1388035,I980233,I979949,I980264,I979961,I980304,I980312,I980329,I980346,I1388029,I980363,I979976,I980394,I1388020,I980411,I1388044,I980428,I1388026,I980454,I979964,I980476,I980493,I979958,I980524,I979952,I979955,I980569,I979967,I980630,I980656,I980673,I980681,I980698,I980715,I980732,I980749,I980766,I980797,I980814,I980845,I980862,I980879,I980910,I980950,I980958,I980975,I980992,I981009,I981040,I981057,I981074,I981100,I981122,I981139,I981170,I981215,I981276,I981302,I981319,I981327,I981344,I981361,I981378,I981395,I981412,I981443,I981460,I981491,I981508,I981525,I981556,I981596,I981604,I981621,I981638,I981655,I981686,I981703,I981720,I981746,I981768,I981785,I981816,I981861,I981922,I981948,I981965,I981973,I981990,I982007,I982024,I982041,I982058,I981908,I982089,I982106,I981911,I982137,I982154,I982171,I981887,I982202,I981899,I982242,I982250,I982267,I982284,I982301,I981914,I982332,I982349,I982366,I982392,I981902,I982414,I982431,I981896,I982462,I981890,I981893,I982507,I981905,I982568,I982594,I982611,I982619,I982636,I982653,I982670,I982687,I982704,I982554,I982735,I982752,I982557,I982783,I982800,I982817,I982533,I982848,I982545,I982888,I982896,I982913,I982930,I982947,I982560,I982978,I982995,I983012,I983038,I982548,I983060,I983077,I982542,I983108,I982536,I982539,I983153,I982551,I983214,I1212340,I983240,I1212346,I983257,I983265,I983282,I1212343,I983299,I1212322,I983316,I1212325,I983333,I1212331,I983350,I983381,I983398,I983429,I983446,I983463,I983494,I983534,I983542,I983559,I983576,I1212334,I983593,I983624,I983641,I1212328,I983658,I1212337,I983684,I983706,I983723,I983754,I983799,I983860,I983886,I983903,I983911,I983928,I983945,I983962,I983979,I983996,I984027,I984044,I984075,I984092,I984109,I984140,I984180,I984188,I984205,I984222,I984239,I984270,I984287,I984304,I984330,I984352,I984369,I984400,I984445,I984506,I984532,I984549,I984557,I984574,I984591,I984608,I984625,I984642,I984673,I984690,I984721,I984738,I984755,I984786,I984826,I984834,I984851,I984868,I984885,I984916,I984933,I984950,I984976,I984998,I985015,I985046,I985091,I985152,I985178,I985195,I985203,I985220,I985237,I985254,I985271,I985288,I985319,I985336,I985367,I985384,I985401,I985432,I985472,I985480,I985497,I985514,I985531,I985562,I985579,I985596,I985622,I985644,I985661,I985692,I985737,I985798,I985824,I985841,I985849,I985866,I985883,I985900,I985917,I985934,I985965,I985982,I986013,I986030,I986047,I986078,I986118,I986126,I986143,I986160,I986177,I986208,I986225,I986242,I986268,I986290,I986307,I986338,I986383,I986444,I1109252,I986470,I1109234,I986487,I986495,I986512,I1109243,I986529,I1109255,I986546,I1109237,I986563,I1109246,I986580,I986611,I986628,I986659,I986676,I1109258,I986693,I986724,I986764,I986772,I986789,I986806,I986823,I986854,I1109240,I986871,I1109249,I986888,I986914,I986936,I986953,I986984,I987029,I987090,I987116,I987133,I987141,I987158,I987175,I987192,I987209,I987226,I987076,I987257,I987274,I987079,I987305,I987322,I987339,I987055,I987370,I987067,I987410,I987418,I987435,I987452,I987469,I987082,I987500,I987517,I987534,I987560,I987070,I987582,I987599,I987064,I987630,I987058,I987061,I987675,I987073,I987736,I987762,I987779,I987787,I987804,I987821,I987838,I987855,I987872,I987722,I987903,I987920,I987725,I987951,I987968,I987985,I987701,I988016,I987713,I988056,I988064,I988081,I988098,I988115,I987728,I988146,I988163,I988180,I988206,I987716,I988228,I988245,I987710,I988276,I987704,I987707,I988321,I987719,I988382,I988408,I988425,I988433,I988450,I988467,I988484,I988501,I988518,I988368,I988549,I988566,I988371,I988597,I988614,I988631,I988347,I988662,I988359,I988702,I988710,I988727,I988744,I988761,I988374,I988792,I988809,I988826,I988852,I988362,I988874,I988891,I988356,I988922,I988350,I988353,I988967,I988365,I989028,I989054,I989071,I989079,I989096,I989113,I989130,I989147,I989164,I989014,I989195,I989212,I989017,I989243,I989260,I989277,I988993,I989308,I989005,I989348,I989356,I989373,I989390,I989407,I989020,I989438,I989455,I989472,I989498,I989008,I989520,I989537,I989002,I989568,I988996,I988999,I989613,I989011,I989674,I989700,I989717,I989725,I989742,I989759,I989776,I989793,I989810,I989660,I989841,I989858,I989663,I989889,I989906,I989923,I989639,I989954,I989651,I989994,I990002,I990019,I990036,I990053,I989666,I990084,I990101,I990118,I990144,I989654,I990166,I990183,I989648,I990214,I989642,I989645,I990259,I989657,I990320,I990346,I990363,I990371,I990388,I990405,I990422,I990439,I990456,I990306,I990487,I990504,I990309,I990535,I990552,I990569,I990285,I990600,I990297,I990640,I990648,I990665,I990682,I990699,I990312,I990730,I990747,I990764,I990790,I990300,I990812,I990829,I990294,I990860,I990288,I990291,I990905,I990303,I990966,I990992,I991009,I991017,I991034,I991051,I991068,I991085,I991102,I991133,I991150,I991181,I991198,I991215,I991246,I991286,I991294,I991311,I991328,I991345,I991376,I991393,I991410,I991436,I991458,I991475,I991506,I991551,I991612,I991638,I991655,I991663,I991680,I991697,I991714,I991731,I991748,I991779,I991796,I991827,I991844,I991861,I991892,I991932,I991940,I991957,I991974,I991991,I992022,I992039,I992056,I992082,I992104,I992121,I992152,I992197,I992258,I992284,I992301,I992309,I992326,I992343,I992360,I992377,I992394,I992425,I992442,I992473,I992490,I992507,I992538,I992578,I992586,I992603,I992620,I992637,I992668,I992685,I992702,I992728,I992750,I992767,I992798,I992843,I992904,I1191906,I992930,I1191888,I992947,I992955,I992972,I1191897,I992989,I1191909,I993006,I1191891,I993023,I1191900,I993040,I992890,I993071,I993088,I992893,I993119,I993136,I1191912,I993153,I992869,I993184,I992881,I993224,I993232,I993249,I993266,I993283,I992896,I993314,I1191894,I993331,I1191903,I993348,I993374,I992884,I993396,I993413,I992878,I993444,I992872,I992875,I993489,I992887,I993550,I993576,I993593,I993601,I993618,I993635,I993652,I993669,I993686,I993536,I993717,I993734,I993539,I993765,I993782,I993799,I993515,I993830,I993527,I993870,I993878,I993895,I993912,I993929,I993542,I993960,I993977,I993994,I994020,I993530,I994042,I994059,I993524,I994090,I993518,I993521,I994135,I993533,I994196,I994222,I994239,I994247,I994264,I994281,I994298,I994315,I994332,I994182,I994363,I994380,I994185,I994411,I994428,I994445,I994161,I994476,I994173,I994516,I994524,I994541,I994558,I994575,I994188,I994606,I994623,I994640,I994666,I994176,I994688,I994705,I994170,I994736,I994164,I994167,I994781,I994179,I994842,I1073994,I994868,I1073976,I994885,I994893,I994910,I1073985,I994927,I1073997,I994944,I1073979,I994961,I1073988,I994978,I995009,I995026,I995057,I995074,I1074000,I995091,I995122,I995162,I995170,I995187,I995204,I995221,I995252,I1073982,I995269,I1073991,I995286,I995312,I995334,I995351,I995382,I995427,I995488,I995514,I995531,I995539,I995556,I995573,I995590,I995607,I995624,I995655,I995672,I995703,I995720,I995737,I995768,I995808,I995816,I995833,I995850,I995867,I995898,I995915,I995932,I995958,I995980,I995997,I996028,I996073,I996134,I996160,I996177,I996185,I996202,I996219,I996236,I996253,I996270,I996301,I996318,I996349,I996366,I996383,I996414,I996454,I996462,I996479,I996496,I996513,I996544,I996561,I996578,I996604,I996626,I996643,I996674,I996719,I996780,I1085554,I996806,I1085536,I996823,I996831,I996848,I1085545,I996865,I1085557,I996882,I1085539,I996899,I1085548,I996916,I996766,I996947,I996964,I996769,I996995,I997012,I1085560,I997029,I996745,I997060,I996757,I997100,I997108,I997125,I997142,I997159,I996772,I997190,I1085542,I997207,I1085551,I997224,I997250,I996760,I997272,I997289,I996754,I997320,I996748,I996751,I997365,I996763,I997426,I997452,I997469,I997477,I997494,I997511,I997528,I997545,I997562,I997593,I997610,I997641,I997658,I997675,I997706,I997746,I997754,I997771,I997788,I997805,I997836,I997853,I997870,I997896,I997918,I997935,I997966,I998011,I998072,I1393967,I998098,I1393991,I998115,I998123,I998140,I1393973,I998157,I1393982,I998174,I998191,I1393988,I998208,I998239,I998256,I998287,I998304,I1393985,I998321,I998352,I998392,I998400,I998417,I998434,I1393979,I998451,I998482,I1393970,I998499,I1393994,I998516,I1393976,I998542,I998564,I998581,I998612,I998657,I998718,I998744,I998761,I998769,I998786,I998803,I998820,I998837,I998854,I998704,I998885,I998902,I998707,I998933,I998950,I998967,I998683,I998998,I998695,I999038,I999046,I999063,I999080,I999097,I998710,I999128,I999145,I999162,I999188,I998698,I999210,I999227,I998692,I999258,I998686,I998689,I999303,I998701,I999364,I1175722,I999390,I1175704,I999407,I999415,I999432,I1175713,I999449,I1175725,I999466,I1175707,I999483,I1175716,I999500,I999531,I999548,I999579,I999596,I1175728,I999613,I999644,I999684,I999692,I999709,I999726,I999743,I999774,I1175710,I999791,I1175719,I999808,I999834,I999856,I999873,I999904,I999949,I1000010,I1000036,I1000053,I1000061,I1000078,I1000095,I1000112,I1000129,I1000146,I1000177,I1000194,I1000225,I1000242,I1000259,I1000290,I1000330,I1000338,I1000355,I1000372,I1000389,I1000420,I1000437,I1000454,I1000480,I1000502,I1000519,I1000550,I1000595,I1000656,I1000682,I1000699,I1000707,I1000724,I1000741,I1000758,I1000775,I1000792,I1000823,I1000840,I1000871,I1000888,I1000905,I1000936,I1000976,I1000984,I1001001,I1001018,I1001035,I1001066,I1001083,I1001100,I1001126,I1001148,I1001165,I1001196,I1001241,I1001302,I1199420,I1001328,I1199402,I1001345,I1001353,I1001370,I1199411,I1001387,I1199423,I1001404,I1199405,I1001421,I1199414,I1001438,I1001288,I1001469,I1001486,I1001291,I1001517,I1001534,I1199426,I1001551,I1001267,I1001582,I1001279,I1001622,I1001630,I1001647,I1001664,I1001681,I1001294,I1001712,I1199408,I1001729,I1199417,I1001746,I1001772,I1001282,I1001794,I1001811,I1001276,I1001842,I1001270,I1001273,I1001887,I1001285,I1001948,I1381472,I1001974,I1381496,I1001991,I1001999,I1002016,I1381478,I1002033,I1381487,I1002050,I1002067,I1381493,I1002084,I1002115,I1002132,I1002163,I1002180,I1381490,I1002197,I1002228,I1002268,I1002276,I1002293,I1002310,I1381484,I1002327,I1002358,I1381475,I1002375,I1381499,I1002392,I1381481,I1002418,I1002440,I1002457,I1002488,I1002533,I1002594,I1083820,I1002620,I1083802,I1002637,I1002645,I1002662,I1083811,I1002679,I1083823,I1002696,I1083805,I1002713,I1083814,I1002730,I1002761,I1002778,I1002809,I1002826,I1083826,I1002843,I1002874,I1002914,I1002922,I1002939,I1002956,I1002973,I1003004,I1083808,I1003021,I1083817,I1003038,I1003064,I1003086,I1003103,I1003134,I1003179,I1003240,I1366597,I1003266,I1366621,I1003283,I1003291,I1003308,I1366603,I1003325,I1366612,I1003342,I1003359,I1366618,I1003376,I1003407,I1003424,I1003455,I1003472,I1366615,I1003489,I1003520,I1003560,I1003568,I1003585,I1003602,I1366609,I1003619,I1003650,I1366600,I1003667,I1366624,I1003684,I1366606,I1003710,I1003732,I1003749,I1003780,I1003825,I1003886,I1003912,I1003929,I1003937,I1003954,I1003971,I1003988,I1004005,I1004022,I1004053,I1004070,I1004101,I1004118,I1004135,I1004166,I1004206,I1004214,I1004231,I1004248,I1004265,I1004296,I1004313,I1004330,I1004356,I1004378,I1004395,I1004426,I1004471,I1004532,I1243348,I1004558,I1243354,I1004575,I1004583,I1004600,I1243351,I1004617,I1243330,I1004634,I1243333,I1004651,I1243339,I1004668,I1004699,I1004716,I1004747,I1004764,I1004781,I1004812,I1004852,I1004860,I1004877,I1004894,I1243342,I1004911,I1004942,I1004959,I1243336,I1004976,I1243345,I1005002,I1005024,I1005041,I1005072,I1005117,I1005178,I1005204,I1005221,I1005229,I1005246,I1005263,I1005280,I1005297,I1005314,I1005164,I1005345,I1005362,I1005167,I1005393,I1005410,I1005427,I1005143,I1005458,I1005155,I1005498,I1005506,I1005523,I1005540,I1005557,I1005170,I1005588,I1005605,I1005622,I1005648,I1005158,I1005670,I1005687,I1005152,I1005718,I1005146,I1005149,I1005763,I1005161,I1005824,I1005850,I1005867,I1005875,I1005892,I1005909,I1005926,I1005943,I1005960,I1005991,I1006008,I1006039,I1006056,I1006073,I1006104,I1006144,I1006152,I1006169,I1006186,I1006203,I1006234,I1006251,I1006268,I1006294,I1006316,I1006333,I1006364,I1006409,I1006470,I1006496,I1006513,I1006521,I1006538,I1006555,I1006572,I1006589,I1006606,I1006456,I1006637,I1006654,I1006459,I1006685,I1006702,I1006719,I1006435,I1006750,I1006447,I1006790,I1006798,I1006815,I1006832,I1006849,I1006462,I1006880,I1006897,I1006914,I1006940,I1006450,I1006962,I1006979,I1006444,I1007010,I1006438,I1006441,I1007055,I1006453,I1007116,I1007142,I1007159,I1007167,I1007184,I1007201,I1007218,I1007235,I1007252,I1007283,I1007300,I1007331,I1007348,I1007365,I1007396,I1007436,I1007444,I1007461,I1007478,I1007495,I1007526,I1007543,I1007560,I1007586,I1007608,I1007625,I1007656,I1007701,I1007762,I1007788,I1007805,I1007813,I1007830,I1007847,I1007864,I1007881,I1007898,I1007929,I1007946,I1007977,I1007994,I1008011,I1008042,I1008082,I1008090,I1008107,I1008124,I1008141,I1008172,I1008189,I1008206,I1008232,I1008254,I1008271,I1008302,I1008347,I1008408,I1008434,I1008451,I1008459,I1008476,I1008493,I1008510,I1008527,I1008544,I1008575,I1008592,I1008623,I1008640,I1008657,I1008688,I1008728,I1008736,I1008753,I1008770,I1008787,I1008818,I1008835,I1008852,I1008878,I1008900,I1008917,I1008948,I1008993,I1009048,I1009074,I1009091,I1009040,I1009113,I1009139,I1009147,I1009164,I1009181,I1009198,I1009215,I1009232,I1009249,I1009022,I1009280,I1009025,I1009311,I1009328,I1009345,I1009362,I1009034,I1009393,I1009037,I1009031,I1009438,I1009455,I1009472,I1009498,I1009506,I1009019,I1009537,I1009554,I1009028,I1009609,I1009635,I1009652,I1009601,I1009674,I1009700,I1009708,I1009725,I1009742,I1009759,I1009776,I1009793,I1009810,I1009583,I1009841,I1009586,I1009872,I1009889,I1009906,I1009923,I1009595,I1009954,I1009598,I1009592,I1009999,I1010016,I1010033,I1010059,I1010067,I1009580,I1010098,I1010115,I1009589,I1010170,I1010196,I1010213,I1010235,I1010261,I1010269,I1010286,I1010303,I1010320,I1010337,I1010354,I1010371,I1010402,I1010433,I1010450,I1010467,I1010484,I1010515,I1010560,I1010577,I1010594,I1010620,I1010628,I1010659,I1010676,I1010731,I1182655,I1010757,I1010774,I1010723,I1010796,I1182646,I1010822,I1010830,I1182643,I1010847,I1010864,I1182652,I1010881,I1182661,I1010898,I1010915,I1182640,I1010932,I1010705,I1010963,I1010708,I1010994,I1182649,I1011011,I1011028,I1011045,I1010717,I1011076,I1010720,I1010714,I1011121,I1182664,I1011138,I1011155,I1182658,I1011181,I1011189,I1010702,I1011220,I1011237,I1010711,I1011292,I1011318,I1011335,I1011284,I1011357,I1011383,I1011391,I1011408,I1011425,I1011442,I1011459,I1011476,I1011493,I1011266,I1011524,I1011269,I1011555,I1011572,I1011589,I1011606,I1011278,I1011637,I1011281,I1011275,I1011682,I1011699,I1011716,I1011742,I1011750,I1011263,I1011781,I1011798,I1011272,I1011853,I1011879,I1011896,I1011918,I1011944,I1011952,I1011969,I1011986,I1012003,I1012020,I1012037,I1012054,I1012085,I1012116,I1012133,I1012150,I1012167,I1012198,I1012243,I1012260,I1012277,I1012303,I1012311,I1012342,I1012359,I1012414,I1292905,I1012440,I1012457,I1012406,I1012479,I1292902,I1012505,I1012513,I1292908,I1012530,I1012547,I1292917,I1012564,I1292911,I1012581,I1012598,I1292923,I1012615,I1012388,I1012646,I1012391,I1012677,I1292920,I1012694,I1012711,I1012728,I1012400,I1012759,I1012403,I1012397,I1012804,I1292914,I1012821,I1292926,I1012838,I1012864,I1012872,I1012385,I1012903,I1012920,I1012394,I1012975,I1013001,I1013018,I1013040,I1013066,I1013074,I1013091,I1013108,I1013125,I1013142,I1013159,I1013176,I1013207,I1013238,I1013255,I1013272,I1013289,I1013320,I1013365,I1013382,I1013399,I1013425,I1013433,I1013464,I1013481,I1013536,I1013562,I1013579,I1013601,I1013627,I1013635,I1013652,I1013669,I1013686,I1013703,I1013720,I1013737,I1013768,I1013799,I1013816,I1013833,I1013850,I1013881,I1013926,I1013943,I1013960,I1013986,I1013994,I1014025,I1014042,I1014097,I1014123,I1014140,I1014162,I1014188,I1014196,I1014213,I1014230,I1014247,I1014264,I1014281,I1014298,I1014329,I1014360,I1014377,I1014394,I1014411,I1014442,I1014487,I1014504,I1014521,I1014547,I1014555,I1014586,I1014603,I1014658,I1014684,I1014701,I1014723,I1014749,I1014757,I1014774,I1014791,I1014808,I1014825,I1014842,I1014859,I1014890,I1014921,I1014938,I1014955,I1014972,I1015003,I1015048,I1015065,I1015082,I1015108,I1015116,I1015147,I1015164,I1015219,I1308897,I1015245,I1015262,I1015284,I1308891,I1015310,I1015318,I1308882,I1015335,I1015352,I1308909,I1015369,I1308894,I1308903,I1015386,I1015403,I1308888,I1015420,I1015451,I1015482,I1308906,I1015499,I1015516,I1015533,I1015564,I1015609,I1308900,I1015626,I1015643,I1308885,I1015669,I1015677,I1015708,I1015725,I1015780,I1015806,I1015823,I1015772,I1015845,I1015871,I1015879,I1015896,I1015913,I1015930,I1015947,I1015964,I1015981,I1015754,I1016012,I1015757,I1016043,I1016060,I1016077,I1016094,I1015766,I1016125,I1015769,I1015763,I1016170,I1016187,I1016204,I1016230,I1016238,I1015751,I1016269,I1016286,I1015760,I1016341,I1016367,I1016384,I1016406,I1016432,I1016440,I1016457,I1016474,I1016491,I1016508,I1016525,I1016542,I1016573,I1016604,I1016621,I1016638,I1016655,I1016686,I1016731,I1016748,I1016765,I1016791,I1016799,I1016830,I1016847,I1016902,I1016928,I1016945,I1016894,I1016967,I1016993,I1017001,I1017018,I1017035,I1017052,I1017069,I1017086,I1017103,I1016876,I1017134,I1016879,I1017165,I1017182,I1017199,I1017216,I1016888,I1017247,I1016891,I1016885,I1017292,I1017309,I1017326,I1017352,I1017360,I1016873,I1017391,I1017408,I1016882,I1017463,I1068789,I1017489,I1017506,I1017455,I1017528,I1068780,I1017554,I1017562,I1068777,I1017579,I1017596,I1068786,I1017613,I1068795,I1017630,I1017647,I1068774,I1017664,I1017437,I1017695,I1017440,I1017726,I1068783,I1017743,I1017760,I1017777,I1017449,I1017808,I1017452,I1017446,I1017853,I1068798,I1017870,I1017887,I1068792,I1017913,I1017921,I1017434,I1017952,I1017969,I1017443,I1018024,I1018050,I1018067,I1018089,I1018115,I1018123,I1018140,I1018157,I1018174,I1018191,I1018208,I1018225,I1018256,I1018287,I1018304,I1018321,I1018338,I1018369,I1018414,I1018431,I1018448,I1018474,I1018482,I1018513,I1018530,I1018585,I1018611,I1018628,I1018577,I1018650,I1018676,I1018684,I1018701,I1018718,I1018735,I1018752,I1018769,I1018786,I1018559,I1018817,I1018562,I1018848,I1018865,I1018882,I1018899,I1018571,I1018930,I1018574,I1018568,I1018975,I1018992,I1019009,I1019035,I1019043,I1018556,I1019074,I1019091,I1018565,I1019146,I1019172,I1019189,I1019211,I1019237,I1019245,I1019262,I1019279,I1019296,I1019313,I1019330,I1019347,I1019378,I1019409,I1019426,I1019443,I1019460,I1019491,I1019536,I1019553,I1019570,I1019596,I1019604,I1019635,I1019652,I1019707,I1067055,I1019733,I1019750,I1019772,I1067046,I1019798,I1019806,I1067043,I1019823,I1019840,I1067052,I1019857,I1067061,I1019874,I1019891,I1067040,I1019908,I1019939,I1019970,I1067049,I1019987,I1020004,I1020021,I1020052,I1020097,I1067064,I1020114,I1020131,I1067058,I1020157,I1020165,I1020196,I1020213,I1020268,I1020294,I1020311,I1020333,I1020359,I1020367,I1020384,I1020401,I1020418,I1020435,I1020452,I1020469,I1020500,I1020531,I1020548,I1020565,I1020582,I1020613,I1020658,I1020675,I1020692,I1020718,I1020726,I1020757,I1020774,I1020829,I1020855,I1020872,I1020821,I1020894,I1020920,I1020928,I1020945,I1020962,I1020979,I1020996,I1021013,I1021030,I1020803,I1021061,I1020806,I1021092,I1021109,I1021126,I1021143,I1020815,I1021174,I1020818,I1020812,I1021219,I1021236,I1021253,I1021279,I1021287,I1020800,I1021318,I1021335,I1020809,I1021390,I1021416,I1021433,I1021455,I1021481,I1021489,I1021506,I1021523,I1021540,I1021557,I1021574,I1021591,I1021622,I1021653,I1021670,I1021687,I1021704,I1021735,I1021780,I1021797,I1021814,I1021840,I1021848,I1021879,I1021896,I1021951,I1021977,I1021994,I1022016,I1022042,I1022050,I1022067,I1022084,I1022101,I1022118,I1022135,I1022152,I1022183,I1022214,I1022231,I1022248,I1022265,I1022296,I1022341,I1022358,I1022375,I1022401,I1022409,I1022440,I1022457,I1022512,I1345787,I1022538,I1022555,I1022504,I1022577,I1345781,I1022603,I1022611,I1345772,I1022628,I1022645,I1345799,I1022662,I1345784,I1345793,I1022679,I1022696,I1345778,I1022713,I1022486,I1022744,I1022489,I1022775,I1345796,I1022792,I1022809,I1022826,I1022498,I1022857,I1022501,I1022495,I1022902,I1345790,I1022919,I1022936,I1345775,I1022962,I1022970,I1022483,I1023001,I1023018,I1022492,I1023073,I1222120,I1023099,I1023116,I1023138,I1222126,I1023164,I1023172,I1222135,I1023189,I1023206,I1222114,I1023223,I1222117,I1023240,I1023257,I1222129,I1023274,I1023305,I1023336,I1222123,I1023353,I1023370,I1023387,I1023418,I1023463,I1222138,I1023480,I1023497,I1222132,I1023523,I1023531,I1023562,I1023579,I1023634,I1023660,I1023677,I1023699,I1023725,I1023733,I1023750,I1023767,I1023784,I1023801,I1023818,I1023835,I1023866,I1023897,I1023914,I1023931,I1023948,I1023979,I1024024,I1024041,I1024058,I1024084,I1024092,I1024123,I1024140,I1024195,I1024221,I1024238,I1024260,I1024286,I1024294,I1024311,I1024328,I1024345,I1024362,I1024379,I1024396,I1024427,I1024458,I1024475,I1024492,I1024509,I1024540,I1024585,I1024602,I1024619,I1024645,I1024653,I1024684,I1024701,I1024756,I1024782,I1024799,I1024821,I1024847,I1024855,I1024872,I1024889,I1024906,I1024923,I1024940,I1024957,I1024988,I1025019,I1025036,I1025053,I1025070,I1025101,I1025146,I1025163,I1025180,I1025206,I1025214,I1025245,I1025262,I1025317,I1230280,I1025343,I1025360,I1025382,I1230286,I1025408,I1025416,I1230295,I1025433,I1025450,I1230274,I1025467,I1230277,I1025484,I1025501,I1230289,I1025518,I1025549,I1025580,I1230283,I1025597,I1025614,I1025631,I1025662,I1025707,I1230298,I1025724,I1025741,I1230292,I1025767,I1025775,I1025806,I1025823,I1025878,I1025904,I1025921,I1025870,I1025943,I1025969,I1025977,I1025994,I1026011,I1026028,I1026045,I1026062,I1026079,I1025852,I1026110,I1025855,I1026141,I1026158,I1026175,I1026192,I1025864,I1026223,I1025867,I1025861,I1026268,I1026285,I1026302,I1026328,I1026336,I1025849,I1026367,I1026384,I1025858,I1026439,I1026465,I1026482,I1026504,I1026530,I1026538,I1026555,I1026572,I1026589,I1026606,I1026623,I1026640,I1026671,I1026702,I1026719,I1026736,I1026753,I1026784,I1026829,I1026846,I1026863,I1026889,I1026897,I1026928,I1026945,I1027000,I1027026,I1027043,I1027065,I1027091,I1027099,I1027116,I1027133,I1027150,I1027167,I1027184,I1027201,I1027232,I1027263,I1027280,I1027297,I1027314,I1027345,I1027390,I1027407,I1027424,I1027450,I1027458,I1027489,I1027506,I1027561,I1027587,I1027604,I1027626,I1027652,I1027660,I1027677,I1027694,I1027711,I1027728,I1027745,I1027762,I1027793,I1027824,I1027841,I1027858,I1027875,I1027906,I1027951,I1027968,I1027985,I1028011,I1028019,I1028050,I1028067,I1028122,I1233544,I1028148,I1028165,I1028187,I1233550,I1028213,I1028221,I1233559,I1028238,I1028255,I1233538,I1028272,I1233541,I1028289,I1028306,I1233553,I1028323,I1028354,I1028385,I1233547,I1028402,I1028419,I1028436,I1028467,I1028512,I1233562,I1028529,I1028546,I1233556,I1028572,I1028580,I1028611,I1028628,I1028683,I1028709,I1028726,I1028748,I1028774,I1028782,I1028799,I1028816,I1028833,I1028850,I1028867,I1028884,I1028915,I1028946,I1028963,I1028980,I1028997,I1029028,I1029073,I1029090,I1029107,I1029133,I1029141,I1029172,I1029189,I1029244,I1029270,I1029287,I1029309,I1029335,I1029343,I1029360,I1029377,I1029394,I1029411,I1029428,I1029445,I1029476,I1029507,I1029524,I1029541,I1029558,I1029589,I1029634,I1029651,I1029668,I1029694,I1029702,I1029733,I1029750,I1029805,I1029831,I1029848,I1029870,I1029896,I1029904,I1029921,I1029938,I1029955,I1029972,I1029989,I1030006,I1030037,I1030068,I1030085,I1030102,I1030119,I1030150,I1030195,I1030212,I1030229,I1030255,I1030263,I1030294,I1030311,I1030366,I1030392,I1030409,I1030431,I1030457,I1030465,I1030482,I1030499,I1030516,I1030533,I1030550,I1030567,I1030598,I1030629,I1030646,I1030663,I1030680,I1030711,I1030756,I1030773,I1030790,I1030816,I1030824,I1030855,I1030872,I1030927,I1030953,I1030970,I1030992,I1031018,I1031026,I1031043,I1031060,I1031077,I1031094,I1031111,I1031128,I1031159,I1031190,I1031207,I1031224,I1031241,I1031272,I1031317,I1031334,I1031351,I1031377,I1031385,I1031416,I1031433,I1031488,I1181499,I1031514,I1031531,I1031553,I1181490,I1031579,I1031587,I1181487,I1031604,I1031621,I1181496,I1031638,I1181505,I1031655,I1031672,I1181484,I1031689,I1031720,I1031751,I1181493,I1031768,I1031785,I1031802,I1031833,I1031878,I1181508,I1031895,I1031912,I1181502,I1031938,I1031946,I1031977,I1031994,I1032049,I1090753,I1032075,I1032092,I1032041,I1032114,I1090744,I1032140,I1032148,I1090741,I1032165,I1032182,I1090750,I1032199,I1090759,I1032216,I1032233,I1090738,I1032250,I1032023,I1032281,I1032026,I1032312,I1090747,I1032329,I1032346,I1032363,I1032035,I1032394,I1032038,I1032032,I1032439,I1090762,I1032456,I1032473,I1090756,I1032499,I1032507,I1032020,I1032538,I1032555,I1032029,I1032610,I1032636,I1032653,I1032602,I1032675,I1032701,I1032709,I1032726,I1032743,I1032760,I1032777,I1032794,I1032811,I1032584,I1032842,I1032587,I1032873,I1032890,I1032907,I1032924,I1032596,I1032955,I1032599,I1032593,I1033000,I1033017,I1033034,I1033060,I1033068,I1032581,I1033099,I1033116,I1032590,I1033171,I1033197,I1033214,I1033236,I1033262,I1033270,I1033287,I1033304,I1033321,I1033338,I1033355,I1033372,I1033403,I1033434,I1033451,I1033468,I1033485,I1033516,I1033561,I1033578,I1033595,I1033621,I1033629,I1033660,I1033677,I1033732,I1033758,I1033775,I1033797,I1033823,I1033831,I1033848,I1033865,I1033882,I1033899,I1033916,I1033933,I1033964,I1033995,I1034012,I1034029,I1034046,I1034077,I1034122,I1034139,I1034156,I1034182,I1034190,I1034221,I1034238,I1034293,I1034319,I1034336,I1034285,I1034358,I1034384,I1034392,I1034409,I1034426,I1034443,I1034460,I1034477,I1034494,I1034267,I1034525,I1034270,I1034556,I1034573,I1034590,I1034607,I1034279,I1034638,I1034282,I1034276,I1034683,I1034700,I1034717,I1034743,I1034751,I1034264,I1034782,I1034799,I1034273,I1034854,I1034880,I1034897,I1034846,I1034919,I1034945,I1034953,I1034970,I1034987,I1035004,I1035021,I1035038,I1035055,I1034828,I1035086,I1034831,I1035117,I1035134,I1035151,I1035168,I1034840,I1035199,I1034843,I1034837,I1035244,I1035261,I1035278,I1035304,I1035312,I1034825,I1035343,I1035360,I1034834,I1035415,I1035441,I1035458,I1035480,I1035506,I1035514,I1035531,I1035548,I1035565,I1035582,I1035599,I1035616,I1035647,I1035678,I1035695,I1035712,I1035729,I1035760,I1035805,I1035822,I1035839,I1035865,I1035873,I1035904,I1035921,I1035976,I1036002,I1036019,I1036041,I1036067,I1036075,I1036092,I1036109,I1036126,I1036143,I1036160,I1036177,I1036208,I1036239,I1036256,I1036273,I1036290,I1036321,I1036366,I1036383,I1036400,I1036426,I1036434,I1036465,I1036482,I1036537,I1036563,I1036580,I1036602,I1036628,I1036636,I1036653,I1036670,I1036687,I1036704,I1036721,I1036738,I1036769,I1036800,I1036817,I1036834,I1036851,I1036882,I1036927,I1036944,I1036961,I1036987,I1036995,I1037026,I1037043,I1037098,I1195949,I1037124,I1037141,I1037163,I1195940,I1037189,I1037197,I1195937,I1037214,I1037231,I1195946,I1037248,I1195955,I1037265,I1037282,I1195934,I1037299,I1037330,I1037361,I1195943,I1037378,I1037395,I1037412,I1037443,I1037488,I1195958,I1037505,I1037522,I1195952,I1037548,I1037556,I1037587,I1037604,I1037659,I1197683,I1037685,I1037702,I1037724,I1197674,I1037750,I1037758,I1197671,I1037775,I1037792,I1197680,I1037809,I1197689,I1037826,I1037843,I1197668,I1037860,I1037891,I1037922,I1197677,I1037939,I1037956,I1037973,I1038004,I1038049,I1197692,I1038066,I1038083,I1197686,I1038109,I1038117,I1038148,I1038165,I1038220,I1038246,I1038263,I1038212,I1038285,I1038311,I1038319,I1038336,I1038353,I1038370,I1038387,I1038404,I1038421,I1038194,I1038452,I1038197,I1038483,I1038500,I1038517,I1038534,I1038206,I1038565,I1038209,I1038203,I1038610,I1038627,I1038644,I1038670,I1038678,I1038191,I1038709,I1038726,I1038200,I1038781,I1038807,I1038824,I1038773,I1038846,I1038872,I1038880,I1038897,I1038914,I1038931,I1038948,I1038965,I1038982,I1038755,I1039013,I1038758,I1039044,I1039061,I1039078,I1039095,I1038767,I1039126,I1038770,I1038764,I1039171,I1039188,I1039205,I1039231,I1039239,I1038752,I1039270,I1039287,I1038761,I1039342,I1039368,I1039385,I1039407,I1039433,I1039441,I1039458,I1039475,I1039492,I1039509,I1039526,I1039543,I1039574,I1039605,I1039622,I1039639,I1039656,I1039687,I1039732,I1039749,I1039766,I1039792,I1039800,I1039831,I1039848,I1039903,I1039929,I1039946,I1039968,I1039994,I1040002,I1040019,I1040036,I1040053,I1040070,I1040087,I1040104,I1040135,I1040166,I1040183,I1040200,I1040217,I1040248,I1040293,I1040310,I1040327,I1040353,I1040361,I1040392,I1040409,I1040464,I1040490,I1040507,I1040456,I1040529,I1040555,I1040563,I1040580,I1040597,I1040614,I1040631,I1040648,I1040665,I1040438,I1040696,I1040441,I1040727,I1040744,I1040761,I1040778,I1040450,I1040809,I1040453,I1040447,I1040854,I1040871,I1040888,I1040914,I1040922,I1040435,I1040953,I1040970,I1040444,I1041025,I1041051,I1041068,I1041090,I1041116,I1041124,I1041141,I1041158,I1041175,I1041192,I1041209,I1041226,I1041257,I1041288,I1041305,I1041322,I1041339,I1041370,I1041415,I1041432,I1041449,I1041475,I1041483,I1041514,I1041531,I1041586,I1180343,I1041612,I1041629,I1041651,I1180334,I1041677,I1041685,I1180331,I1041702,I1041719,I1180340,I1041736,I1180349,I1041753,I1041770,I1180328,I1041787,I1041818,I1041849,I1180337,I1041866,I1041883,I1041900,I1041931,I1041976,I1180352,I1041993,I1042010,I1180346,I1042036,I1042044,I1042075,I1042092,I1042147,I1042173,I1042190,I1042212,I1042238,I1042246,I1042263,I1042280,I1042297,I1042314,I1042331,I1042348,I1042379,I1042410,I1042427,I1042444,I1042461,I1042492,I1042537,I1042554,I1042571,I1042597,I1042605,I1042636,I1042653,I1042708,I1042734,I1042751,I1042773,I1042799,I1042807,I1042824,I1042841,I1042858,I1042875,I1042892,I1042909,I1042940,I1042971,I1042988,I1043005,I1043022,I1043053,I1043098,I1043115,I1043132,I1043158,I1043166,I1043197,I1043214,I1043269,I1248232,I1043295,I1043312,I1043334,I1248238,I1043360,I1043368,I1248247,I1043385,I1043402,I1248226,I1043419,I1248229,I1043436,I1043453,I1248241,I1043470,I1043501,I1043532,I1248235,I1043549,I1043566,I1043583,I1043614,I1043659,I1248250,I1043676,I1043693,I1248244,I1043719,I1043727,I1043758,I1043775,I1043830,I1043856,I1043873,I1043895,I1043921,I1043929,I1043946,I1043963,I1043980,I1043997,I1044014,I1044031,I1044062,I1044093,I1044110,I1044127,I1044144,I1044175,I1044220,I1044237,I1044254,I1044280,I1044288,I1044319,I1044336,I1044391,I1044417,I1044434,I1044383,I1044456,I1044482,I1044490,I1044507,I1044524,I1044541,I1044558,I1044575,I1044592,I1044365,I1044623,I1044368,I1044654,I1044671,I1044688,I1044705,I1044377,I1044736,I1044380,I1044374,I1044781,I1044798,I1044815,I1044841,I1044849,I1044362,I1044880,I1044897,I1044371,I1044952,I1044978,I1044995,I1045017,I1045043,I1045051,I1045068,I1045085,I1045102,I1045119,I1045136,I1045153,I1045184,I1045215,I1045232,I1045249,I1045266,I1045297,I1045342,I1045359,I1045376,I1045402,I1045410,I1045441,I1045458,I1045513,I1045539,I1045556,I1045578,I1045604,I1045612,I1045629,I1045646,I1045663,I1045680,I1045697,I1045714,I1045745,I1045776,I1045793,I1045810,I1045827,I1045858,I1045903,I1045920,I1045937,I1045963,I1045971,I1046002,I1046019,I1046074,I1385057,I1046100,I1046117,I1046066,I1046139,I1385051,I1046165,I1046173,I1385042,I1046190,I1046207,I1385069,I1046224,I1385054,I1385063,I1046241,I1046258,I1385048,I1046275,I1046048,I1046306,I1046051,I1046337,I1385066,I1046354,I1046371,I1046388,I1046060,I1046419,I1046063,I1046057,I1046464,I1385060,I1046481,I1046498,I1385045,I1046524,I1046532,I1046045,I1046563,I1046580,I1046054,I1046635,I1046661,I1046678,I1046627,I1046700,I1046726,I1046734,I1046751,I1046768,I1046785,I1046802,I1046819,I1046836,I1046609,I1046867,I1046612,I1046898,I1046915,I1046932,I1046949,I1046621,I1046980,I1046624,I1046618,I1047025,I1047042,I1047059,I1047085,I1047093,I1046606,I1047124,I1047141,I1046615,I1047196,I1047222,I1047239,I1047261,I1047287,I1047295,I1047312,I1047329,I1047346,I1047363,I1047380,I1047397,I1047428,I1047459,I1047476,I1047493,I1047510,I1047541,I1047586,I1047603,I1047620,I1047646,I1047654,I1047685,I1047702,I1047757,I1047783,I1047800,I1047822,I1047848,I1047856,I1047873,I1047890,I1047907,I1047924,I1047941,I1047958,I1047989,I1048020,I1048037,I1048054,I1048071,I1048102,I1048147,I1048164,I1048181,I1048207,I1048215,I1048246,I1048263,I1048318,I1048344,I1048361,I1048383,I1048409,I1048417,I1048434,I1048451,I1048468,I1048485,I1048502,I1048519,I1048550,I1048581,I1048598,I1048615,I1048632,I1048663,I1048708,I1048725,I1048742,I1048768,I1048776,I1048807,I1048824,I1048879,I1048905,I1048922,I1048944,I1048970,I1048978,I1048995,I1049012,I1049029,I1049046,I1049063,I1049080,I1049111,I1049142,I1049159,I1049176,I1049193,I1049224,I1049269,I1049286,I1049303,I1049329,I1049337,I1049368,I1049385,I1049440,I1049466,I1049483,I1049505,I1049531,I1049539,I1049556,I1049573,I1049590,I1049607,I1049624,I1049641,I1049672,I1049703,I1049720,I1049737,I1049754,I1049785,I1049830,I1049847,I1049864,I1049890,I1049898,I1049929,I1049946,I1050001,I1050027,I1050044,I1050066,I1050092,I1050100,I1050117,I1050134,I1050151,I1050168,I1050185,I1050202,I1050233,I1050264,I1050281,I1050298,I1050315,I1050346,I1050391,I1050408,I1050425,I1050451,I1050459,I1050490,I1050507,I1050562,I1050588,I1050605,I1050627,I1050653,I1050661,I1050678,I1050695,I1050712,I1050729,I1050746,I1050763,I1050794,I1050825,I1050842,I1050859,I1050876,I1050907,I1050952,I1050969,I1050986,I1051012,I1051020,I1051051,I1051068,I1051123,I1075725,I1051149,I1051166,I1051115,I1051188,I1075716,I1051214,I1051222,I1075713,I1051239,I1051256,I1075722,I1051273,I1075731,I1051290,I1051307,I1075710,I1051324,I1051097,I1051355,I1051100,I1051386,I1075719,I1051403,I1051420,I1051437,I1051109,I1051468,I1051112,I1051106,I1051513,I1075734,I1051530,I1051547,I1075728,I1051573,I1051581,I1051094,I1051612,I1051629,I1051103,I1051684,I1323177,I1051710,I1051727,I1051749,I1323171,I1051775,I1051783,I1323162,I1051800,I1051817,I1323189,I1051834,I1323174,I1323183,I1051851,I1051868,I1323168,I1051885,I1051916,I1051947,I1323186,I1051964,I1051981,I1051998,I1052029,I1052074,I1323180,I1052091,I1052108,I1323165,I1052134,I1052142,I1052173,I1052190,I1052245,I1332697,I1052271,I1052288,I1052310,I1332691,I1052336,I1052344,I1332682,I1052361,I1052378,I1332709,I1052395,I1332694,I1332703,I1052412,I1052429,I1332688,I1052446,I1052477,I1052508,I1332706,I1052525,I1052542,I1052559,I1052590,I1052635,I1332700,I1052652,I1052669,I1332685,I1052695,I1052703,I1052734,I1052751,I1052806,I1052832,I1052849,I1052798,I1052871,I1052897,I1052905,I1052922,I1052939,I1052956,I1052973,I1052990,I1053007,I1052780,I1053038,I1052783,I1053069,I1053086,I1053103,I1053120,I1052792,I1053151,I1052795,I1052789,I1053196,I1053213,I1053230,I1053256,I1053264,I1052777,I1053295,I1053312,I1052786,I1053367,I1063009,I1053393,I1053410,I1053359,I1053432,I1063000,I1053458,I1053466,I1062997,I1053483,I1053500,I1063006,I1053517,I1063015,I1053534,I1053551,I1062994,I1053568,I1053341,I1053599,I1053344,I1053630,I1063003,I1053647,I1053664,I1053681,I1053353,I1053712,I1053356,I1053350,I1053757,I1063018,I1053774,I1053791,I1063012,I1053817,I1053825,I1053338,I1053856,I1053873,I1053347,I1053928,I1210696,I1053954,I1053971,I1053993,I1210702,I1054019,I1054027,I1210711,I1054044,I1054061,I1210690,I1054078,I1210693,I1054095,I1054112,I1210705,I1054129,I1054160,I1054191,I1210699,I1054208,I1054225,I1054242,I1054273,I1054318,I1210714,I1054335,I1054352,I1210708,I1054378,I1054386,I1054417,I1054434,I1054489,I1054515,I1054532,I1054481,I1054554,I1054580,I1054588,I1054605,I1054622,I1054639,I1054656,I1054673,I1054690,I1054463,I1054721,I1054466,I1054752,I1054769,I1054786,I1054803,I1054475,I1054834,I1054478,I1054472,I1054879,I1054896,I1054913,I1054939,I1054947,I1054460,I1054978,I1054995,I1054469,I1055050,I1055076,I1055093,I1055115,I1055141,I1055149,I1055166,I1055183,I1055200,I1055217,I1055234,I1055251,I1055282,I1055313,I1055330,I1055347,I1055364,I1055395,I1055440,I1055457,I1055474,I1055500,I1055508,I1055539,I1055556,I1055611,I1055637,I1055654,I1055676,I1055702,I1055710,I1055727,I1055744,I1055761,I1055778,I1055795,I1055812,I1055843,I1055874,I1055891,I1055908,I1055925,I1055956,I1056001,I1056018,I1056035,I1056061,I1056069,I1056100,I1056117,I1056172,I1056198,I1056215,I1056237,I1056263,I1056271,I1056288,I1056305,I1056322,I1056339,I1056356,I1056373,I1056404,I1056435,I1056452,I1056469,I1056486,I1056517,I1056562,I1056579,I1056596,I1056622,I1056630,I1056661,I1056678,I1056733,I1137571,I1056759,I1056776,I1056798,I1137562,I1056824,I1056832,I1137559,I1056849,I1056866,I1137568,I1056883,I1137577,I1056900,I1056917,I1137556,I1056934,I1056965,I1056996,I1137565,I1057013,I1057030,I1057047,I1057078,I1057123,I1137580,I1057140,I1057157,I1137574,I1057183,I1057191,I1057222,I1057239,I1057294,I1057320,I1057337,I1057359,I1057385,I1057393,I1057410,I1057427,I1057444,I1057461,I1057478,I1057495,I1057526,I1057557,I1057574,I1057591,I1057608,I1057639,I1057684,I1057701,I1057718,I1057744,I1057752,I1057783,I1057800,I1057855,I1057881,I1057898,I1057920,I1057946,I1057954,I1057971,I1057988,I1058005,I1058022,I1058039,I1058056,I1058087,I1058118,I1058135,I1058152,I1058169,I1058200,I1058245,I1058262,I1058279,I1058305,I1058313,I1058344,I1058361,I1058416,I1058442,I1058459,I1058481,I1058507,I1058515,I1058532,I1058549,I1058566,I1058583,I1058600,I1058617,I1058648,I1058679,I1058696,I1058713,I1058730,I1058761,I1058806,I1058823,I1058840,I1058866,I1058874,I1058905,I1058922,I1058980,I1059006,I1059014,I1059054,I1059062,I1059079,I1059096,I1059136,I1059158,I1059175,I1059201,I1059209,I1059226,I1059243,I1059260,I1059277,I1059322,I1059353,I1059370,I1059396,I1059404,I1059435,I1059452,I1059469,I1059486,I1059558,I1059584,I1059592,I1059632,I1059640,I1059657,I1059674,I1059714,I1059736,I1059753,I1059779,I1059787,I1059804,I1059821,I1059838,I1059855,I1059900,I1059931,I1059948,I1059974,I1059982,I1060013,I1060030,I1060047,I1060064,I1060136,I1060162,I1060170,I1060210,I1060218,I1060235,I1060252,I1060292,I1060314,I1060331,I1060357,I1060365,I1060382,I1060399,I1060416,I1060433,I1060478,I1060509,I1060526,I1060552,I1060560,I1060591,I1060608,I1060625,I1060642,I1060714,I1060740,I1060748,I1060788,I1060796,I1060813,I1060830,I1060870,I1060892,I1060909,I1060935,I1060943,I1060960,I1060977,I1060994,I1061011,I1061056,I1061087,I1061104,I1061130,I1061138,I1061169,I1061186,I1061203,I1061220,I1061292,I1061318,I1061326,I1061366,I1061374,I1061391,I1061408,I1061448,I1061470,I1061487,I1061513,I1061521,I1061538,I1061555,I1061572,I1061589,I1061634,I1061665,I1061682,I1061708,I1061716,I1061747,I1061764,I1061781,I1061798,I1061870,I1061896,I1061904,I1061944,I1061952,I1061969,I1061986,I1062026,I1062048,I1062065,I1062091,I1062099,I1062116,I1062133,I1062150,I1062167,I1062212,I1062243,I1062260,I1062286,I1062294,I1062325,I1062342,I1062359,I1062376,I1062448,I1062474,I1062482,I1062522,I1062530,I1062547,I1062564,I1062604,I1062626,I1062643,I1062669,I1062677,I1062694,I1062711,I1062728,I1062745,I1062790,I1062821,I1062838,I1062864,I1062872,I1062903,I1062920,I1062937,I1062954,I1063026,I1063052,I1063060,I1063100,I1063108,I1063125,I1063142,I1063182,I1063204,I1063221,I1063247,I1063255,I1063272,I1063289,I1063306,I1063323,I1063368,I1063399,I1063416,I1063442,I1063450,I1063481,I1063498,I1063515,I1063532,I1063604,I1063630,I1063638,I1063678,I1063686,I1063703,I1063720,I1063760,I1063782,I1063799,I1063825,I1063833,I1063850,I1063867,I1063884,I1063901,I1063946,I1063977,I1063994,I1064020,I1064028,I1064059,I1064076,I1064093,I1064110,I1064182,I1064208,I1064216,I1064256,I1064264,I1064281,I1064298,I1064338,I1064360,I1064377,I1064403,I1064411,I1064428,I1064445,I1064462,I1064479,I1064524,I1064555,I1064572,I1064598,I1064606,I1064637,I1064654,I1064671,I1064688,I1064760,I1064786,I1064794,I1064834,I1064842,I1064859,I1064876,I1064916,I1064938,I1064955,I1064981,I1064989,I1065006,I1065023,I1065040,I1065057,I1065102,I1065133,I1065150,I1065176,I1065184,I1065215,I1065232,I1065249,I1065266,I1065338,I1065364,I1065372,I1065412,I1065420,I1065437,I1065454,I1065494,I1065516,I1065533,I1065559,I1065567,I1065584,I1065601,I1065618,I1065635,I1065680,I1065711,I1065728,I1065754,I1065762,I1065793,I1065810,I1065827,I1065844,I1065916,I1065942,I1065950,I1065990,I1065998,I1066015,I1066032,I1066072,I1066094,I1066111,I1066137,I1066145,I1066162,I1066179,I1066196,I1066213,I1066258,I1066289,I1066306,I1066332,I1066340,I1066371,I1066388,I1066405,I1066422,I1066494,I1066520,I1066528,I1066568,I1066576,I1066593,I1066610,I1066650,I1066672,I1066689,I1066715,I1066723,I1066740,I1066757,I1066774,I1066791,I1066836,I1066867,I1066884,I1066910,I1066918,I1066949,I1066966,I1066983,I1067000,I1067072,I1067098,I1067106,I1067146,I1067154,I1067171,I1067188,I1067228,I1067250,I1067267,I1067293,I1067301,I1067318,I1067335,I1067352,I1067369,I1067414,I1067445,I1067462,I1067488,I1067496,I1067527,I1067544,I1067561,I1067578,I1067650,I1067676,I1067684,I1067724,I1067732,I1067749,I1067766,I1067806,I1067828,I1067845,I1067871,I1067879,I1067896,I1067913,I1067930,I1067947,I1067992,I1068023,I1068040,I1068066,I1068074,I1068105,I1068122,I1068139,I1068156,I1068228,I1068254,I1068262,I1068302,I1068310,I1068327,I1068344,I1068384,I1068406,I1068423,I1068449,I1068457,I1068474,I1068491,I1068508,I1068525,I1068570,I1068601,I1068618,I1068644,I1068652,I1068683,I1068700,I1068717,I1068734,I1068806,I1068832,I1068840,I1068880,I1068888,I1068905,I1068922,I1068962,I1068984,I1069001,I1069027,I1069035,I1069052,I1069069,I1069086,I1069103,I1069148,I1069179,I1069196,I1069222,I1069230,I1069261,I1069278,I1069295,I1069312,I1069384,I1069410,I1069418,I1069458,I1069466,I1069483,I1069500,I1069540,I1069562,I1069579,I1069605,I1069613,I1069630,I1069647,I1069664,I1069681,I1069726,I1069757,I1069774,I1069800,I1069808,I1069839,I1069856,I1069873,I1069890,I1069962,I1228119,I1069988,I1069996,I1228113,I1228098,I1070036,I1070044,I1228104,I1070061,I1228116,I1070078,I1070118,I1070140,I1070157,I1070183,I1070191,I1070208,I1228122,I1070225,I1228110,I1070242,I1070259,I1070304,I1228101,I1070335,I1070352,I1228107,I1070378,I1070386,I1070417,I1070434,I1070451,I1070468,I1070540,I1070566,I1070574,I1070614,I1070622,I1070639,I1070656,I1070696,I1070718,I1070735,I1070761,I1070769,I1070786,I1070803,I1070820,I1070837,I1070882,I1070913,I1070930,I1070956,I1070964,I1070995,I1071012,I1071029,I1071046,I1071118,I1329139,I1071144,I1071152,I1329121,I1329112,I1071192,I1071200,I1329127,I1071217,I1329115,I1071234,I1071274,I1071296,I1329124,I1071313,I1071339,I1071347,I1071364,I1329133,I1071381,I1071398,I1071415,I1071460,I1329136,I1071491,I1071508,I1329130,I1329118,I1071534,I1071542,I1071573,I1071590,I1071607,I1071624,I1071696,I1071722,I1071730,I1071770,I1071778,I1071795,I1071812,I1071852,I1071874,I1071891,I1071917,I1071925,I1071942,I1071959,I1071976,I1071993,I1072038,I1072069,I1072086,I1072112,I1072120,I1072151,I1072168,I1072185,I1072202,I1072274,I1072300,I1072308,I1072348,I1072356,I1072373,I1072390,I1072430,I1072452,I1072469,I1072495,I1072503,I1072520,I1072537,I1072554,I1072571,I1072616,I1072647,I1072664,I1072690,I1072698,I1072729,I1072746,I1072763,I1072780,I1072852,I1256512,I1072878,I1072886,I1256494,I1256503,I1072926,I1072934,I1256488,I1072951,I1256500,I1072968,I1073008,I1073030,I1256491,I1073047,I1073073,I1073081,I1073098,I1073115,I1073132,I1073149,I1073194,I1256509,I1073225,I1073242,I1256497,I1256506,I1073268,I1073276,I1073307,I1073324,I1073341,I1073358,I1073430,I1073456,I1073464,I1073504,I1073512,I1073529,I1073546,I1073586,I1073608,I1073625,I1073651,I1073659,I1073676,I1073693,I1073710,I1073727,I1073772,I1073803,I1073820,I1073846,I1073854,I1073885,I1073902,I1073919,I1073936,I1074008,I1074034,I1074042,I1074082,I1074090,I1074107,I1074124,I1074164,I1074186,I1074203,I1074229,I1074237,I1074254,I1074271,I1074288,I1074305,I1074350,I1074381,I1074398,I1074424,I1074432,I1074463,I1074480,I1074497,I1074514,I1074586,I1074612,I1074620,I1074660,I1074668,I1074685,I1074702,I1074742,I1074764,I1074781,I1074807,I1074815,I1074832,I1074849,I1074866,I1074883,I1074928,I1074959,I1074976,I1075002,I1075010,I1075041,I1075058,I1075075,I1075092,I1075164,I1075190,I1075198,I1075238,I1075246,I1075263,I1075280,I1075320,I1075342,I1075359,I1075385,I1075393,I1075410,I1075427,I1075444,I1075461,I1075506,I1075537,I1075554,I1075580,I1075588,I1075619,I1075636,I1075653,I1075670,I1075742,I1379714,I1075768,I1075776,I1379696,I1379687,I1075816,I1075824,I1379702,I1075841,I1379690,I1075858,I1075898,I1075920,I1379699,I1075937,I1075963,I1075971,I1075988,I1379708,I1076005,I1076022,I1076039,I1076084,I1379711,I1076115,I1076132,I1379705,I1379693,I1076158,I1076166,I1076197,I1076214,I1076231,I1076248,I1076320,I1076346,I1076354,I1076394,I1076402,I1076419,I1076436,I1076476,I1076498,I1076515,I1076541,I1076549,I1076566,I1076583,I1076600,I1076617,I1076662,I1076693,I1076710,I1076736,I1076744,I1076775,I1076792,I1076809,I1076826,I1076898,I1076924,I1076932,I1076972,I1076980,I1076997,I1077014,I1077054,I1077076,I1077093,I1077119,I1077127,I1077144,I1077161,I1077178,I1077195,I1077240,I1077271,I1077288,I1077314,I1077322,I1077353,I1077370,I1077387,I1077404,I1077476,I1077502,I1077510,I1077550,I1077558,I1077575,I1077592,I1077632,I1077654,I1077671,I1077697,I1077705,I1077722,I1077739,I1077756,I1077773,I1077818,I1077849,I1077866,I1077892,I1077900,I1077931,I1077948,I1077965,I1077982,I1078054,I1078080,I1078088,I1078128,I1078136,I1078153,I1078170,I1078210,I1078232,I1078249,I1078275,I1078283,I1078300,I1078317,I1078334,I1078351,I1078396,I1078427,I1078444,I1078470,I1078478,I1078509,I1078526,I1078543,I1078560,I1078632,I1257668,I1078658,I1078666,I1257650,I1257659,I1078706,I1078714,I1257644,I1078731,I1257656,I1078748,I1078788,I1078810,I1257647,I1078827,I1078853,I1078861,I1078878,I1078895,I1078912,I1078929,I1078974,I1257665,I1079005,I1079022,I1257653,I1257662,I1079048,I1079056,I1079087,I1079104,I1079121,I1079138,I1079210,I1079236,I1079244,I1079284,I1079292,I1079309,I1079326,I1079366,I1079388,I1079405,I1079431,I1079439,I1079456,I1079473,I1079490,I1079507,I1079552,I1079583,I1079600,I1079626,I1079634,I1079665,I1079682,I1079699,I1079716,I1079788,I1079814,I1079822,I1079862,I1079870,I1079887,I1079904,I1079944,I1079966,I1079983,I1080009,I1080017,I1080034,I1080051,I1080068,I1080085,I1080130,I1080161,I1080178,I1080204,I1080212,I1080243,I1080260,I1080277,I1080294,I1080366,I1342229,I1080392,I1080400,I1342211,I1342202,I1080440,I1080448,I1342217,I1080465,I1342205,I1080482,I1080522,I1080544,I1342214,I1080561,I1080587,I1080595,I1080612,I1342223,I1080629,I1080646,I1080663,I1080708,I1342226,I1080739,I1080756,I1342220,I1342208,I1080782,I1080790,I1080821,I1080838,I1080855,I1080872,I1080944,I1080970,I1080978,I1081018,I1081026,I1081043,I1081060,I1081100,I1081122,I1081139,I1081165,I1081173,I1081190,I1081207,I1081224,I1081241,I1081286,I1081317,I1081334,I1081360,I1081368,I1081399,I1081416,I1081433,I1081450,I1081522,I1081548,I1081556,I1081596,I1081604,I1081621,I1081638,I1081678,I1081700,I1081717,I1081743,I1081751,I1081768,I1081785,I1081802,I1081819,I1081864,I1081895,I1081912,I1081938,I1081946,I1081977,I1081994,I1082011,I1082028,I1082100,I1276164,I1082126,I1082134,I1276146,I1276155,I1082174,I1082182,I1276140,I1082199,I1276152,I1082216,I1082256,I1082278,I1276143,I1082295,I1082321,I1082329,I1082346,I1082363,I1082380,I1082397,I1082442,I1276161,I1082473,I1082490,I1276149,I1276158,I1082516,I1082524,I1082555,I1082572,I1082589,I1082606,I1082678,I1082704,I1082712,I1082752,I1082760,I1082777,I1082794,I1082834,I1082856,I1082873,I1082899,I1082907,I1082924,I1082941,I1082958,I1082975,I1083020,I1083051,I1083068,I1083094,I1083102,I1083133,I1083150,I1083167,I1083184,I1083256,I1083282,I1083290,I1083330,I1083338,I1083355,I1083372,I1083412,I1083434,I1083451,I1083477,I1083485,I1083502,I1083519,I1083536,I1083553,I1083598,I1083629,I1083646,I1083672,I1083680,I1083711,I1083728,I1083745,I1083762,I1083834,I1083860,I1083868,I1083908,I1083916,I1083933,I1083950,I1083990,I1084012,I1084029,I1084055,I1084063,I1084080,I1084097,I1084114,I1084131,I1084176,I1084207,I1084224,I1084250,I1084258,I1084289,I1084306,I1084323,I1084340,I1084412,I1393399,I1084438,I1084446,I1393381,I1393372,I1084486,I1084494,I1393387,I1084511,I1393375,I1084528,I1084568,I1084590,I1393384,I1084607,I1084633,I1084641,I1084658,I1393393,I1084675,I1084692,I1084709,I1084754,I1393396,I1084785,I1084802,I1393390,I1393378,I1084828,I1084836,I1084867,I1084884,I1084901,I1084918,I1084990,I1085016,I1085024,I1084973,I1085064,I1085072,I1085089,I1085106,I1084961,I1085146,I1084982,I1085168,I1085185,I1085211,I1085219,I1085236,I1085253,I1085270,I1085287,I1084958,I1084979,I1085332,I1084970,I1085363,I1085380,I1085406,I1085414,I1084976,I1085445,I1085462,I1085479,I1085496,I1084967,I1084964,I1085568,I1085594,I1085602,I1085642,I1085650,I1085667,I1085684,I1085724,I1085746,I1085763,I1085789,I1085797,I1085814,I1085831,I1085848,I1085865,I1085910,I1085941,I1085958,I1085984,I1085992,I1086023,I1086040,I1086057,I1086074,I1086146,I1227031,I1086172,I1086180,I1227025,I1227010,I1086220,I1086228,I1227016,I1086245,I1227028,I1086262,I1086302,I1086324,I1086341,I1086367,I1086375,I1086392,I1227034,I1086409,I1227022,I1086426,I1086443,I1086488,I1227013,I1086519,I1086536,I1227019,I1086562,I1086570,I1086601,I1086618,I1086635,I1086652,I1086724,I1261714,I1086750,I1086758,I1261696,I1261705,I1086798,I1086806,I1261690,I1086823,I1261702,I1086840,I1086880,I1086902,I1261693,I1086919,I1086945,I1086953,I1086970,I1086987,I1087004,I1087021,I1087066,I1261711,I1087097,I1087114,I1261699,I1261708,I1087140,I1087148,I1087179,I1087196,I1087213,I1087230,I1087302,I1087328,I1087336,I1087285,I1087376,I1087384,I1087401,I1087418,I1087273,I1087458,I1087294,I1087480,I1087497,I1087523,I1087531,I1087548,I1087565,I1087582,I1087599,I1087270,I1087291,I1087644,I1087282,I1087675,I1087692,I1087718,I1087726,I1087288,I1087757,I1087774,I1087791,I1087808,I1087279,I1087276,I1087880,I1358294,I1087906,I1087914,I1358276,I1087863,I1358267,I1087954,I1087962,I1358282,I1087979,I1358270,I1087996,I1087851,I1088036,I1087872,I1088058,I1358279,I1088075,I1088101,I1088109,I1088126,I1358288,I1088143,I1088160,I1088177,I1087848,I1087869,I1088222,I1358291,I1087860,I1088253,I1088270,I1358285,I1358273,I1088296,I1088304,I1087866,I1088335,I1088352,I1088369,I1088386,I1087857,I1087854,I1088458,I1088484,I1088492,I1088532,I1088540,I1088557,I1088574,I1088614,I1088636,I1088653,I1088679,I1088687,I1088704,I1088721,I1088738,I1088755,I1088800,I1088831,I1088848,I1088874,I1088882,I1088913,I1088930,I1088947,I1088964,I1089036,I1089062,I1089070,I1089019,I1089110,I1089118,I1089135,I1089152,I1089007,I1089192,I1089028,I1089214,I1089231,I1089257,I1089265,I1089282,I1089299,I1089316,I1089333,I1089004,I1089025,I1089378,I1089016,I1089409,I1089426,I1089452,I1089460,I1089022,I1089491,I1089508,I1089525,I1089542,I1089013,I1089010,I1089614,I1089640,I1089648,I1089688,I1089696,I1089713,I1089730,I1089770,I1089792,I1089809,I1089835,I1089843,I1089860,I1089877,I1089894,I1089911,I1089956,I1089987,I1090004,I1090030,I1090038,I1090069,I1090086,I1090103,I1090120,I1090192,I1090218,I1090226,I1090266,I1090274,I1090291,I1090308,I1090348,I1090370,I1090387,I1090413,I1090421,I1090438,I1090455,I1090472,I1090489,I1090534,I1090565,I1090582,I1090608,I1090616,I1090647,I1090664,I1090681,I1090698,I1090770,I1240087,I1090796,I1090804,I1240081,I1240066,I1090844,I1090852,I1240072,I1090869,I1240084,I1090886,I1090926,I1090948,I1090965,I1090991,I1090999,I1091016,I1240090,I1091033,I1240078,I1091050,I1091067,I1091112,I1240069,I1091143,I1091160,I1240075,I1091186,I1091194,I1091225,I1091242,I1091259,I1091276,I1091348,I1091374,I1091382,I1091422,I1091430,I1091447,I1091464,I1091504,I1091526,I1091543,I1091569,I1091577,I1091594,I1091611,I1091628,I1091645,I1091690,I1091721,I1091738,I1091764,I1091772,I1091803,I1091820,I1091837,I1091854,I1091926,I1091952,I1091960,I1092000,I1092008,I1092025,I1092042,I1092082,I1092104,I1092121,I1092147,I1092155,I1092172,I1092189,I1092206,I1092223,I1092268,I1092299,I1092316,I1092342,I1092350,I1092381,I1092398,I1092415,I1092432,I1092504,I1310694,I1092530,I1092538,I1310676,I1310667,I1092578,I1092586,I1310682,I1092603,I1310670,I1092620,I1092660,I1092682,I1310679,I1092699,I1092725,I1092733,I1092750,I1310688,I1092767,I1092784,I1092801,I1092846,I1310691,I1092877,I1092894,I1310685,I1310673,I1092920,I1092928,I1092959,I1092976,I1092993,I1093010,I1093082,I1093108,I1093116,I1093156,I1093164,I1093181,I1093198,I1093238,I1093260,I1093277,I1093303,I1093311,I1093328,I1093345,I1093362,I1093379,I1093424,I1093455,I1093472,I1093498,I1093506,I1093537,I1093554,I1093571,I1093588,I1093660,I1093686,I1093694,I1093734,I1093742,I1093759,I1093776,I1093816,I1093838,I1093855,I1093881,I1093889,I1093906,I1093923,I1093940,I1093957,I1094002,I1094033,I1094050,I1094076,I1094084,I1094115,I1094132,I1094149,I1094166,I1094238,I1094264,I1094272,I1094221,I1094312,I1094320,I1094337,I1094354,I1094209,I1094394,I1094230,I1094416,I1094433,I1094459,I1094467,I1094484,I1094501,I1094518,I1094535,I1094206,I1094227,I1094580,I1094218,I1094611,I1094628,I1094654,I1094662,I1094224,I1094693,I1094710,I1094727,I1094744,I1094215,I1094212,I1094816,I1094842,I1094850,I1094799,I1094890,I1094898,I1094915,I1094932,I1094787,I1094972,I1094808,I1094994,I1095011,I1095037,I1095045,I1095062,I1095079,I1095096,I1095113,I1094784,I1094805,I1095158,I1094796,I1095189,I1095206,I1095232,I1095240,I1094802,I1095271,I1095288,I1095305,I1095322,I1094793,I1094790,I1095394,I1275008,I1095420,I1095428,I1274990,I1274999,I1095468,I1095476,I1274984,I1095493,I1274996,I1095510,I1095550,I1095572,I1274987,I1095589,I1095615,I1095623,I1095640,I1095657,I1095674,I1095691,I1095736,I1275005,I1095767,I1095784,I1274993,I1275002,I1095810,I1095818,I1095849,I1095866,I1095883,I1095900,I1095972,I1233015,I1095998,I1096006,I1233009,I1232994,I1096046,I1096054,I1233000,I1096071,I1233012,I1096088,I1096128,I1096150,I1096167,I1096193,I1096201,I1096218,I1233018,I1096235,I1233006,I1096252,I1096269,I1096314,I1232997,I1096345,I1096362,I1233003,I1096388,I1096396,I1096427,I1096444,I1096461,I1096478,I1096550,I1096576,I1096584,I1096624,I1096632,I1096649,I1096666,I1096706,I1096728,I1096745,I1096771,I1096779,I1096796,I1096813,I1096830,I1096847,I1096892,I1096923,I1096940,I1096966,I1096974,I1097005,I1097022,I1097039,I1097056,I1097128,I1097154,I1097162,I1097202,I1097210,I1097227,I1097244,I1097284,I1097306,I1097323,I1097349,I1097357,I1097374,I1097391,I1097408,I1097425,I1097470,I1097501,I1097518,I1097544,I1097552,I1097583,I1097600,I1097617,I1097634,I1097706,I1097732,I1097740,I1097780,I1097788,I1097805,I1097822,I1097862,I1097884,I1097901,I1097927,I1097935,I1097952,I1097969,I1097986,I1098003,I1098048,I1098079,I1098096,I1098122,I1098130,I1098161,I1098178,I1098195,I1098212,I1098284,I1098310,I1098318,I1098358,I1098366,I1098383,I1098400,I1098440,I1098462,I1098479,I1098505,I1098513,I1098530,I1098547,I1098564,I1098581,I1098626,I1098657,I1098674,I1098700,I1098708,I1098739,I1098756,I1098773,I1098790,I1098862,I1098888,I1098896,I1098936,I1098944,I1098961,I1098978,I1099018,I1099040,I1099057,I1099083,I1099091,I1099108,I1099125,I1099142,I1099159,I1099204,I1099235,I1099252,I1099278,I1099286,I1099317,I1099334,I1099351,I1099368,I1099440,I1099466,I1099474,I1099514,I1099522,I1099539,I1099556,I1099596,I1099618,I1099635,I1099661,I1099669,I1099686,I1099703,I1099720,I1099737,I1099782,I1099813,I1099830,I1099856,I1099864,I1099895,I1099912,I1099929,I1099946,I1100018,I1100044,I1100052,I1100092,I1100100,I1100117,I1100134,I1100174,I1100196,I1100213,I1100239,I1100247,I1100264,I1100281,I1100298,I1100315,I1100360,I1100391,I1100408,I1100434,I1100442,I1100473,I1100490,I1100507,I1100524,I1100596,I1100622,I1100630,I1100579,I1100670,I1100678,I1100695,I1100712,I1100567,I1100752,I1100588,I1100774,I1100791,I1100817,I1100825,I1100842,I1100859,I1100876,I1100893,I1100564,I1100585,I1100938,I1100576,I1100969,I1100986,I1101012,I1101020,I1100582,I1101051,I1101068,I1101085,I1101102,I1100573,I1100570,I1101174,I1101200,I1101208,I1101248,I1101256,I1101273,I1101290,I1101330,I1101352,I1101369,I1101395,I1101403,I1101420,I1101437,I1101454,I1101471,I1101516,I1101547,I1101564,I1101590,I1101598,I1101629,I1101646,I1101663,I1101680,I1101752,I1101778,I1101786,I1101826,I1101834,I1101851,I1101868,I1101908,I1101930,I1101947,I1101973,I1101981,I1101998,I1102015,I1102032,I1102049,I1102094,I1102125,I1102142,I1102168,I1102176,I1102207,I1102224,I1102241,I1102258,I1102330,I1102356,I1102364,I1102404,I1102412,I1102429,I1102446,I1102486,I1102508,I1102525,I1102551,I1102559,I1102576,I1102593,I1102610,I1102627,I1102672,I1102703,I1102720,I1102746,I1102754,I1102785,I1102802,I1102819,I1102836,I1102908,I1102934,I1102942,I1102982,I1102990,I1103007,I1103024,I1103064,I1103086,I1103103,I1103129,I1103137,I1103154,I1103171,I1103188,I1103205,I1103250,I1103281,I1103298,I1103324,I1103332,I1103363,I1103380,I1103397,I1103414,I1103486,I1103512,I1103520,I1103469,I1103560,I1103568,I1103585,I1103602,I1103457,I1103642,I1103478,I1103664,I1103681,I1103707,I1103715,I1103732,I1103749,I1103766,I1103783,I1103454,I1103475,I1103828,I1103466,I1103859,I1103876,I1103902,I1103910,I1103472,I1103941,I1103958,I1103975,I1103992,I1103463,I1103460,I1104064,I1104090,I1104098,I1104047,I1104138,I1104146,I1104163,I1104180,I1104035,I1104220,I1104056,I1104242,I1104259,I1104285,I1104293,I1104310,I1104327,I1104344,I1104361,I1104032,I1104053,I1104406,I1104044,I1104437,I1104454,I1104480,I1104488,I1104050,I1104519,I1104536,I1104553,I1104570,I1104041,I1104038,I1104642,I1291192,I1104668,I1104676,I1291174,I1291183,I1104716,I1104724,I1291168,I1104741,I1291180,I1104758,I1104798,I1104820,I1291171,I1104837,I1104863,I1104871,I1104888,I1104905,I1104922,I1104939,I1104984,I1291189,I1105015,I1105032,I1291177,I1291186,I1105058,I1105066,I1105097,I1105114,I1105131,I1105148,I1105220,I1105246,I1105254,I1105203,I1105294,I1105302,I1105319,I1105336,I1105191,I1105376,I1105212,I1105398,I1105415,I1105441,I1105449,I1105466,I1105483,I1105500,I1105517,I1105188,I1105209,I1105562,I1105200,I1105593,I1105610,I1105636,I1105644,I1105206,I1105675,I1105692,I1105709,I1105726,I1105197,I1105194,I1105798,I1105824,I1105832,I1105872,I1105880,I1105897,I1105914,I1105954,I1105976,I1105993,I1106019,I1106027,I1106044,I1106061,I1106078,I1106095,I1106140,I1106171,I1106188,I1106214,I1106222,I1106253,I1106270,I1106287,I1106304,I1106376,I1106402,I1106410,I1106450,I1106458,I1106475,I1106492,I1106532,I1106554,I1106571,I1106597,I1106605,I1106622,I1106639,I1106656,I1106673,I1106718,I1106749,I1106766,I1106792,I1106800,I1106831,I1106848,I1106865,I1106882,I1106954,I1106980,I1106988,I1107028,I1107036,I1107053,I1107070,I1107110,I1107132,I1107149,I1107175,I1107183,I1107200,I1107217,I1107234,I1107251,I1107296,I1107327,I1107344,I1107370,I1107378,I1107409,I1107426,I1107443,I1107460,I1107532,I1240631,I1107558,I1107566,I1240625,I1240610,I1107606,I1107614,I1240616,I1107631,I1240628,I1107648,I1107688,I1107710,I1107727,I1107753,I1107761,I1107778,I1240634,I1107795,I1240622,I1107812,I1107829,I1107874,I1240613,I1107905,I1107922,I1240619,I1107948,I1107956,I1107987,I1108004,I1108021,I1108038,I1108110,I1108136,I1108144,I1108184,I1108192,I1108209,I1108226,I1108266,I1108288,I1108305,I1108331,I1108339,I1108356,I1108373,I1108390,I1108407,I1108452,I1108483,I1108500,I1108526,I1108534,I1108565,I1108582,I1108599,I1108616,I1108688,I1108714,I1108722,I1108762,I1108770,I1108787,I1108804,I1108844,I1108866,I1108883,I1108909,I1108917,I1108934,I1108951,I1108968,I1108985,I1109030,I1109061,I1109078,I1109104,I1109112,I1109143,I1109160,I1109177,I1109194,I1109266,I1109292,I1109300,I1109340,I1109348,I1109365,I1109382,I1109422,I1109444,I1109461,I1109487,I1109495,I1109512,I1109529,I1109546,I1109563,I1109608,I1109639,I1109656,I1109682,I1109690,I1109721,I1109738,I1109755,I1109772,I1109844,I1109870,I1109878,I1109918,I1109926,I1109943,I1109960,I1110000,I1110022,I1110039,I1110065,I1110073,I1110090,I1110107,I1110124,I1110141,I1110186,I1110217,I1110234,I1110260,I1110268,I1110299,I1110316,I1110333,I1110350,I1110422,I1338659,I1110448,I1110456,I1338641,I1338632,I1110496,I1110504,I1338647,I1110521,I1338635,I1110538,I1110578,I1110600,I1338644,I1110617,I1110643,I1110651,I1110668,I1338653,I1110685,I1110702,I1110719,I1110764,I1338656,I1110795,I1110812,I1338650,I1338638,I1110838,I1110846,I1110877,I1110894,I1110911,I1110928,I1111000,I1324974,I1111026,I1111034,I1324956,I1324947,I1111074,I1111082,I1324962,I1111099,I1324950,I1111116,I1111156,I1111178,I1324959,I1111195,I1111221,I1111229,I1111246,I1324968,I1111263,I1111280,I1111297,I1111342,I1324971,I1111373,I1111390,I1324965,I1324953,I1111416,I1111424,I1111455,I1111472,I1111489,I1111506,I1111578,I1236279,I1111604,I1111612,I1236273,I1111561,I1236258,I1111652,I1111660,I1236264,I1111677,I1236276,I1111694,I1111549,I1111734,I1111570,I1111756,I1111773,I1111799,I1111807,I1111824,I1236282,I1111841,I1236270,I1111858,I1111875,I1111546,I1111567,I1111920,I1236261,I1111558,I1111951,I1111968,I1236267,I1111994,I1112002,I1111564,I1112033,I1112050,I1112067,I1112084,I1111555,I1111552,I1112156,I1112182,I1112190,I1112230,I1112238,I1112255,I1112272,I1112312,I1112334,I1112351,I1112377,I1112385,I1112402,I1112419,I1112436,I1112453,I1112498,I1112529,I1112546,I1112572,I1112580,I1112611,I1112628,I1112645,I1112662,I1112734,I1112760,I1112768,I1112808,I1112816,I1112833,I1112850,I1112890,I1112912,I1112929,I1112955,I1112963,I1112980,I1112997,I1113014,I1113031,I1113076,I1113107,I1113124,I1113150,I1113158,I1113189,I1113206,I1113223,I1113240,I1113312,I1113338,I1113346,I1113386,I1113394,I1113411,I1113428,I1113468,I1113490,I1113507,I1113533,I1113541,I1113558,I1113575,I1113592,I1113609,I1113654,I1113685,I1113702,I1113728,I1113736,I1113767,I1113784,I1113801,I1113818,I1113890,I1254778,I1113916,I1113924,I1254760,I1113873,I1254769,I1113964,I1113972,I1254754,I1113989,I1254766,I1114006,I1113861,I1114046,I1113882,I1114068,I1254757,I1114085,I1114111,I1114119,I1114136,I1114153,I1114170,I1114187,I1113858,I1113879,I1114232,I1254775,I1113870,I1114263,I1114280,I1254763,I1254772,I1114306,I1114314,I1113876,I1114345,I1114362,I1114379,I1114396,I1113867,I1113864,I1114468,I1114494,I1114502,I1114542,I1114550,I1114567,I1114584,I1114624,I1114646,I1114663,I1114689,I1114697,I1114714,I1114731,I1114748,I1114765,I1114810,I1114841,I1114858,I1114884,I1114892,I1114923,I1114940,I1114957,I1114974,I1115046,I1115072,I1115080,I1115120,I1115128,I1115145,I1115162,I1115202,I1115224,I1115241,I1115267,I1115275,I1115292,I1115309,I1115326,I1115343,I1115388,I1115419,I1115436,I1115462,I1115470,I1115501,I1115518,I1115535,I1115552,I1115624,I1115650,I1115658,I1115698,I1115706,I1115723,I1115740,I1115780,I1115802,I1115819,I1115845,I1115853,I1115870,I1115887,I1115904,I1115921,I1115966,I1115997,I1116014,I1116040,I1116048,I1116079,I1116096,I1116113,I1116130,I1116202,I1116228,I1116236,I1116276,I1116284,I1116301,I1116318,I1116358,I1116380,I1116397,I1116423,I1116431,I1116448,I1116465,I1116482,I1116499,I1116544,I1116575,I1116592,I1116618,I1116626,I1116657,I1116674,I1116691,I1116708,I1116780,I1116806,I1116814,I1116854,I1116862,I1116879,I1116896,I1116936,I1116958,I1116975,I1117001,I1117009,I1117026,I1117043,I1117060,I1117077,I1117122,I1117153,I1117170,I1117196,I1117204,I1117235,I1117252,I1117269,I1117286,I1117358,I1117384,I1117392,I1117341,I1117432,I1117440,I1117457,I1117474,I1117329,I1117514,I1117350,I1117536,I1117553,I1117579,I1117587,I1117604,I1117621,I1117638,I1117655,I1117326,I1117347,I1117700,I1117338,I1117731,I1117748,I1117774,I1117782,I1117344,I1117813,I1117830,I1117847,I1117864,I1117335,I1117332,I1117936,I1117962,I1117970,I1118010,I1118018,I1118035,I1118052,I1118092,I1118114,I1118131,I1118157,I1118165,I1118182,I1118199,I1118216,I1118233,I1118278,I1118309,I1118326,I1118352,I1118360,I1118391,I1118408,I1118425,I1118442,I1118514,I1118540,I1118548,I1118588,I1118596,I1118613,I1118630,I1118670,I1118692,I1118709,I1118735,I1118743,I1118760,I1118777,I1118794,I1118811,I1118856,I1118887,I1118904,I1118930,I1118938,I1118969,I1118986,I1119003,I1119020,I1119092,I1119118,I1119126,I1119166,I1119174,I1119191,I1119208,I1119248,I1119270,I1119287,I1119313,I1119321,I1119338,I1119355,I1119372,I1119389,I1119434,I1119465,I1119482,I1119508,I1119516,I1119547,I1119564,I1119581,I1119598,I1119670,I1119696,I1119704,I1119744,I1119752,I1119769,I1119786,I1119826,I1119848,I1119865,I1119891,I1119899,I1119916,I1119933,I1119950,I1119967,I1120012,I1120043,I1120060,I1120086,I1120094,I1120125,I1120142,I1120159,I1120176,I1120248,I1120274,I1120282,I1120322,I1120330,I1120347,I1120364,I1120404,I1120426,I1120443,I1120469,I1120477,I1120494,I1120511,I1120528,I1120545,I1120590,I1120621,I1120638,I1120664,I1120672,I1120703,I1120720,I1120737,I1120754,I1120826,I1355914,I1120852,I1120860,I1355896,I1355887,I1120900,I1120908,I1355902,I1120925,I1355890,I1120942,I1120982,I1121004,I1355899,I1121021,I1121047,I1121055,I1121072,I1355908,I1121089,I1121106,I1121123,I1121168,I1355911,I1121199,I1121216,I1355905,I1355893,I1121242,I1121250,I1121281,I1121298,I1121315,I1121332,I1121404,I1121430,I1121438,I1121478,I1121486,I1121503,I1121520,I1121560,I1121582,I1121599,I1121625,I1121633,I1121650,I1121667,I1121684,I1121701,I1121746,I1121777,I1121794,I1121820,I1121828,I1121859,I1121876,I1121893,I1121910,I1121982,I1122008,I1122016,I1122056,I1122064,I1122081,I1122098,I1122138,I1122160,I1122177,I1122203,I1122211,I1122228,I1122245,I1122262,I1122279,I1122324,I1122355,I1122372,I1122398,I1122406,I1122437,I1122454,I1122471,I1122488,I1122560,I1394589,I1122586,I1122594,I1394571,I1394562,I1122634,I1122642,I1394577,I1122659,I1394565,I1122676,I1122716,I1122738,I1394574,I1122755,I1122781,I1122789,I1122806,I1394583,I1122823,I1122840,I1122857,I1122902,I1394586,I1122933,I1122950,I1394580,I1394568,I1122976,I1122984,I1123015,I1123032,I1123049,I1123066,I1123138,I1123164,I1123172,I1123212,I1123220,I1123237,I1123254,I1123294,I1123316,I1123333,I1123359,I1123367,I1123384,I1123401,I1123418,I1123435,I1123480,I1123511,I1123528,I1123554,I1123562,I1123593,I1123610,I1123627,I1123644,I1123716,I1123742,I1123750,I1123790,I1123798,I1123815,I1123832,I1123872,I1123894,I1123911,I1123937,I1123945,I1123962,I1123979,I1123996,I1124013,I1124058,I1124089,I1124106,I1124132,I1124140,I1124171,I1124188,I1124205,I1124222,I1124294,I1124320,I1124328,I1124368,I1124376,I1124393,I1124410,I1124450,I1124472,I1124489,I1124515,I1124523,I1124540,I1124557,I1124574,I1124591,I1124636,I1124667,I1124684,I1124710,I1124718,I1124749,I1124766,I1124783,I1124800,I1124872,I1124898,I1124906,I1124855,I1124946,I1124954,I1124971,I1124988,I1124843,I1125028,I1124864,I1125050,I1125067,I1125093,I1125101,I1125118,I1125135,I1125152,I1125169,I1124840,I1124861,I1125214,I1124852,I1125245,I1125262,I1125288,I1125296,I1124858,I1125327,I1125344,I1125361,I1125378,I1124849,I1124846,I1125450,I1125476,I1125484,I1125524,I1125532,I1125549,I1125566,I1125606,I1125628,I1125645,I1125671,I1125679,I1125696,I1125713,I1125730,I1125747,I1125792,I1125823,I1125840,I1125866,I1125874,I1125905,I1125922,I1125939,I1125956,I1126028,I1126054,I1126062,I1126102,I1126110,I1126127,I1126144,I1126184,I1126206,I1126223,I1126249,I1126257,I1126274,I1126291,I1126308,I1126325,I1126370,I1126401,I1126418,I1126444,I1126452,I1126483,I1126500,I1126517,I1126534,I1126606,I1126632,I1126640,I1126680,I1126688,I1126705,I1126722,I1126762,I1126784,I1126801,I1126827,I1126835,I1126852,I1126869,I1126886,I1126903,I1126948,I1126979,I1126996,I1127022,I1127030,I1127061,I1127078,I1127095,I1127112,I1127184,I1127210,I1127218,I1127258,I1127266,I1127283,I1127300,I1127340,I1127362,I1127379,I1127405,I1127413,I1127430,I1127447,I1127464,I1127481,I1127526,I1127557,I1127574,I1127600,I1127608,I1127639,I1127656,I1127673,I1127690,I1127762,I1377334,I1127788,I1127796,I1377316,I1127745,I1377307,I1127836,I1127844,I1377322,I1127861,I1377310,I1127878,I1127733,I1127918,I1127754,I1127940,I1377319,I1127957,I1127983,I1127991,I1128008,I1377328,I1128025,I1128042,I1128059,I1127730,I1127751,I1128104,I1377331,I1127742,I1128135,I1128152,I1377325,I1377313,I1128178,I1128186,I1127748,I1128217,I1128234,I1128251,I1128268,I1127739,I1127736,I1128340,I1128366,I1128374,I1128414,I1128422,I1128439,I1128456,I1128496,I1128518,I1128535,I1128561,I1128569,I1128586,I1128603,I1128620,I1128637,I1128682,I1128713,I1128730,I1128756,I1128764,I1128795,I1128812,I1128829,I1128846,I1128918,I1364839,I1128944,I1128952,I1364821,I1364812,I1128992,I1129000,I1364827,I1129017,I1364815,I1129034,I1129074,I1129096,I1364824,I1129113,I1129139,I1129147,I1129164,I1364833,I1129181,I1129198,I1129215,I1129260,I1364836,I1129291,I1129308,I1364830,I1364818,I1129334,I1129342,I1129373,I1129390,I1129407,I1129424,I1129496,I1129522,I1129530,I1129570,I1129578,I1129595,I1129612,I1129652,I1129674,I1129691,I1129717,I1129725,I1129742,I1129759,I1129776,I1129793,I1129838,I1129869,I1129886,I1129912,I1129920,I1129951,I1129968,I1129985,I1130002,I1130074,I1130100,I1130108,I1130148,I1130156,I1130173,I1130190,I1130230,I1130252,I1130269,I1130295,I1130303,I1130320,I1130337,I1130354,I1130371,I1130416,I1130447,I1130464,I1130490,I1130498,I1130529,I1130546,I1130563,I1130580,I1130652,I1130678,I1130686,I1130726,I1130734,I1130751,I1130768,I1130808,I1130830,I1130847,I1130873,I1130881,I1130898,I1130915,I1130932,I1130949,I1130994,I1131025,I1131042,I1131068,I1131076,I1131107,I1131124,I1131141,I1131158,I1131230,I1259402,I1131256,I1131264,I1259384,I1259393,I1131304,I1131312,I1259378,I1131329,I1259390,I1131346,I1131386,I1131408,I1259381,I1131425,I1131451,I1131459,I1131476,I1131493,I1131510,I1131527,I1131572,I1259399,I1131603,I1131620,I1259387,I1259396,I1131646,I1131654,I1131685,I1131702,I1131719,I1131736,I1131808,I1131834,I1131842,I1131882,I1131890,I1131907,I1131924,I1131964,I1131986,I1132003,I1132029,I1132037,I1132054,I1132071,I1132088,I1132105,I1132150,I1132181,I1132198,I1132224,I1132232,I1132263,I1132280,I1132297,I1132314,I1132386,I1132412,I1132420,I1132460,I1132468,I1132485,I1132502,I1132542,I1132564,I1132581,I1132607,I1132615,I1132632,I1132649,I1132666,I1132683,I1132728,I1132759,I1132776,I1132802,I1132810,I1132841,I1132858,I1132875,I1132892,I1132964,I1132990,I1132998,I1133038,I1133046,I1133063,I1133080,I1133120,I1133142,I1133159,I1133185,I1133193,I1133210,I1133227,I1133244,I1133261,I1133306,I1133337,I1133354,I1133380,I1133388,I1133419,I1133436,I1133453,I1133470,I1133542,I1133568,I1133576,I1133616,I1133624,I1133641,I1133658,I1133698,I1133720,I1133737,I1133763,I1133771,I1133788,I1133805,I1133822,I1133839,I1133884,I1133915,I1133932,I1133958,I1133966,I1133997,I1134014,I1134031,I1134048,I1134120,I1134146,I1134154,I1134103,I1134194,I1134202,I1134219,I1134236,I1134091,I1134276,I1134112,I1134298,I1134315,I1134341,I1134349,I1134366,I1134383,I1134400,I1134417,I1134088,I1134109,I1134462,I1134100,I1134493,I1134510,I1134536,I1134544,I1134106,I1134575,I1134592,I1134609,I1134626,I1134097,I1134094,I1134698,I1266338,I1134724,I1134732,I1266320,I1266329,I1134772,I1134780,I1266314,I1134797,I1266326,I1134814,I1134854,I1134876,I1266317,I1134893,I1134919,I1134927,I1134944,I1134961,I1134978,I1134995,I1135040,I1266335,I1135071,I1135088,I1266323,I1266332,I1135114,I1135122,I1135153,I1135170,I1135187,I1135204,I1135276,I1135302,I1135310,I1135350,I1135358,I1135375,I1135392,I1135432,I1135454,I1135471,I1135497,I1135505,I1135522,I1135539,I1135556,I1135573,I1135618,I1135649,I1135666,I1135692,I1135700,I1135731,I1135748,I1135765,I1135782,I1135854,I1135880,I1135888,I1135837,I1135928,I1135936,I1135953,I1135970,I1135825,I1136010,I1135846,I1136032,I1136049,I1136075,I1136083,I1136100,I1136117,I1136134,I1136151,I1135822,I1135843,I1136196,I1135834,I1136227,I1136244,I1136270,I1136278,I1135840,I1136309,I1136326,I1136343,I1136360,I1135831,I1135828,I1136432,I1136458,I1136466,I1136506,I1136514,I1136531,I1136548,I1136588,I1136610,I1136627,I1136653,I1136661,I1136678,I1136695,I1136712,I1136729,I1136774,I1136805,I1136822,I1136848,I1136856,I1136887,I1136904,I1136921,I1136938,I1137010,I1137036,I1137044,I1137084,I1137092,I1137109,I1137126,I1137166,I1137188,I1137205,I1137231,I1137239,I1137256,I1137273,I1137290,I1137307,I1137352,I1137383,I1137400,I1137426,I1137434,I1137465,I1137482,I1137499,I1137516,I1137588,I1137614,I1137622,I1137662,I1137670,I1137687,I1137704,I1137744,I1137766,I1137783,I1137809,I1137817,I1137834,I1137851,I1137868,I1137885,I1137930,I1137961,I1137978,I1138004,I1138012,I1138043,I1138060,I1138077,I1138094,I1138166,I1138192,I1138200,I1138240,I1138248,I1138265,I1138282,I1138322,I1138344,I1138361,I1138387,I1138395,I1138412,I1138429,I1138446,I1138463,I1138508,I1138539,I1138556,I1138582,I1138590,I1138621,I1138638,I1138655,I1138672,I1138744,I1138770,I1138778,I1138818,I1138826,I1138843,I1138860,I1138900,I1138922,I1138939,I1138965,I1138973,I1138990,I1139007,I1139024,I1139041,I1139086,I1139117,I1139134,I1139160,I1139168,I1139199,I1139216,I1139233,I1139250,I1139322,I1139348,I1139356,I1139396,I1139404,I1139421,I1139438,I1139478,I1139500,I1139517,I1139543,I1139551,I1139568,I1139585,I1139602,I1139619,I1139664,I1139695,I1139712,I1139738,I1139746,I1139777,I1139794,I1139811,I1139828,I1139900,I1139926,I1139934,I1139974,I1139982,I1139999,I1140016,I1140056,I1140078,I1140095,I1140121,I1140129,I1140146,I1140163,I1140180,I1140197,I1140242,I1140273,I1140290,I1140316,I1140324,I1140355,I1140372,I1140389,I1140406,I1140478,I1140504,I1140512,I1140461,I1140552,I1140560,I1140577,I1140594,I1140449,I1140634,I1140470,I1140656,I1140673,I1140699,I1140707,I1140724,I1140741,I1140758,I1140775,I1140446,I1140467,I1140820,I1140458,I1140851,I1140868,I1140894,I1140902,I1140464,I1140933,I1140950,I1140967,I1140984,I1140455,I1140452,I1141056,I1141082,I1141090,I1141130,I1141138,I1141155,I1141172,I1141212,I1141234,I1141251,I1141277,I1141285,I1141302,I1141319,I1141336,I1141353,I1141398,I1141429,I1141446,I1141472,I1141480,I1141511,I1141528,I1141545,I1141562,I1141634,I1141660,I1141668,I1141617,I1141708,I1141716,I1141733,I1141750,I1141605,I1141790,I1141626,I1141812,I1141829,I1141855,I1141863,I1141880,I1141897,I1141914,I1141931,I1141602,I1141623,I1141976,I1141614,I1142007,I1142024,I1142050,I1142058,I1141620,I1142089,I1142106,I1142123,I1142140,I1141611,I1141608,I1142212,I1142238,I1142246,I1142286,I1142294,I1142311,I1142328,I1142368,I1142390,I1142407,I1142433,I1142441,I1142458,I1142475,I1142492,I1142509,I1142554,I1142585,I1142602,I1142628,I1142636,I1142667,I1142684,I1142701,I1142718,I1142790,I1142816,I1142824,I1142864,I1142872,I1142889,I1142906,I1142946,I1142968,I1142985,I1143011,I1143019,I1143036,I1143053,I1143070,I1143087,I1143132,I1143163,I1143180,I1143206,I1143214,I1143245,I1143262,I1143279,I1143296,I1143368,I1143394,I1143402,I1143442,I1143450,I1143467,I1143484,I1143524,I1143546,I1143563,I1143589,I1143597,I1143614,I1143631,I1143648,I1143665,I1143710,I1143741,I1143758,I1143784,I1143792,I1143823,I1143840,I1143857,I1143874,I1143946,I1143972,I1143980,I1144020,I1144028,I1144045,I1144062,I1144102,I1144124,I1144141,I1144167,I1144175,I1144192,I1144209,I1144226,I1144243,I1144288,I1144319,I1144336,I1144362,I1144370,I1144401,I1144418,I1144435,I1144452,I1144524,I1144550,I1144558,I1144507,I1144598,I1144606,I1144623,I1144640,I1144495,I1144680,I1144516,I1144702,I1144719,I1144745,I1144753,I1144770,I1144787,I1144804,I1144821,I1144492,I1144513,I1144866,I1144504,I1144897,I1144914,I1144940,I1144948,I1144510,I1144979,I1144996,I1145013,I1145030,I1144501,I1144498,I1145102,I1224311,I1145128,I1145136,I1224305,I1224290,I1145176,I1145184,I1224296,I1145201,I1224308,I1145218,I1145258,I1145280,I1145297,I1145323,I1145331,I1145348,I1224314,I1145365,I1224302,I1145382,I1145399,I1145444,I1224293,I1145475,I1145492,I1224299,I1145518,I1145526,I1145557,I1145574,I1145591,I1145608,I1145680,I1145706,I1145714,I1145754,I1145762,I1145779,I1145796,I1145836,I1145858,I1145875,I1145901,I1145909,I1145926,I1145943,I1145960,I1145977,I1146022,I1146053,I1146070,I1146096,I1146104,I1146135,I1146152,I1146169,I1146186,I1146258,I1146284,I1146292,I1146332,I1146340,I1146357,I1146374,I1146414,I1146436,I1146453,I1146479,I1146487,I1146504,I1146521,I1146538,I1146555,I1146600,I1146631,I1146648,I1146674,I1146682,I1146713,I1146730,I1146747,I1146764,I1146836,I1146862,I1146870,I1146910,I1146918,I1146935,I1146952,I1146992,I1147014,I1147031,I1147057,I1147065,I1147082,I1147099,I1147116,I1147133,I1147178,I1147209,I1147226,I1147252,I1147260,I1147291,I1147308,I1147325,I1147342,I1147414,I1147440,I1147448,I1147488,I1147496,I1147513,I1147530,I1147570,I1147592,I1147609,I1147635,I1147643,I1147660,I1147677,I1147694,I1147711,I1147756,I1147787,I1147804,I1147830,I1147838,I1147869,I1147886,I1147903,I1147920,I1147992,I1148018,I1148026,I1147975,I1148066,I1148074,I1148091,I1148108,I1147963,I1148148,I1147984,I1148170,I1148187,I1148213,I1148221,I1148238,I1148255,I1148272,I1148289,I1147960,I1147981,I1148334,I1147972,I1148365,I1148382,I1148408,I1148416,I1147978,I1148447,I1148464,I1148481,I1148498,I1147969,I1147966,I1148570,I1148596,I1148604,I1148644,I1148652,I1148669,I1148686,I1148726,I1148748,I1148765,I1148791,I1148799,I1148816,I1148833,I1148850,I1148867,I1148912,I1148943,I1148960,I1148986,I1148994,I1149025,I1149042,I1149059,I1149076,I1149148,I1149174,I1149182,I1149222,I1149230,I1149247,I1149264,I1149304,I1149326,I1149343,I1149369,I1149377,I1149394,I1149411,I1149428,I1149445,I1149490,I1149521,I1149538,I1149564,I1149572,I1149603,I1149620,I1149637,I1149654,I1149726,I1149752,I1149760,I1149800,I1149808,I1149825,I1149842,I1149882,I1149904,I1149921,I1149947,I1149955,I1149972,I1149989,I1150006,I1150023,I1150068,I1150099,I1150116,I1150142,I1150150,I1150181,I1150198,I1150215,I1150232,I1150304,I1150330,I1150338,I1150378,I1150386,I1150403,I1150420,I1150460,I1150482,I1150499,I1150525,I1150533,I1150550,I1150567,I1150584,I1150601,I1150646,I1150677,I1150694,I1150720,I1150728,I1150759,I1150776,I1150793,I1150810,I1150882,I1150908,I1150916,I1150956,I1150964,I1150981,I1150998,I1151038,I1151060,I1151077,I1151103,I1151111,I1151128,I1151145,I1151162,I1151179,I1151224,I1151255,I1151272,I1151298,I1151306,I1151337,I1151354,I1151371,I1151388,I1151460,I1151486,I1151494,I1151534,I1151542,I1151559,I1151576,I1151616,I1151638,I1151655,I1151681,I1151689,I1151706,I1151723,I1151740,I1151757,I1151802,I1151833,I1151850,I1151876,I1151884,I1151915,I1151932,I1151949,I1151966,I1152038,I1152064,I1152072,I1152112,I1152120,I1152137,I1152154,I1152194,I1152216,I1152233,I1152259,I1152267,I1152284,I1152301,I1152318,I1152335,I1152380,I1152411,I1152428,I1152454,I1152462,I1152493,I1152510,I1152527,I1152544,I1152616,I1152642,I1152650,I1152599,I1152690,I1152698,I1152715,I1152732,I1152587,I1152772,I1152608,I1152794,I1152811,I1152837,I1152845,I1152862,I1152879,I1152896,I1152913,I1152584,I1152605,I1152958,I1152596,I1152989,I1153006,I1153032,I1153040,I1152602,I1153071,I1153088,I1153105,I1153122,I1152593,I1152590,I1153194,I1218871,I1153220,I1153228,I1218865,I1218850,I1153268,I1153276,I1218856,I1153293,I1218868,I1153310,I1153350,I1153372,I1153389,I1153415,I1153423,I1153440,I1218874,I1153457,I1218862,I1153474,I1153491,I1153536,I1218853,I1153567,I1153584,I1218859,I1153610,I1153618,I1153649,I1153666,I1153683,I1153700,I1153772,I1153798,I1153806,I1153846,I1153854,I1153871,I1153888,I1153928,I1153950,I1153967,I1153993,I1154001,I1154018,I1154035,I1154052,I1154069,I1154114,I1154145,I1154162,I1154188,I1154196,I1154227,I1154244,I1154261,I1154278,I1154350,I1154376,I1154384,I1154424,I1154432,I1154449,I1154466,I1154506,I1154528,I1154545,I1154571,I1154579,I1154596,I1154613,I1154630,I1154647,I1154692,I1154723,I1154740,I1154766,I1154774,I1154805,I1154822,I1154839,I1154856,I1154928,I1346989,I1154954,I1154962,I1346971,I1154911,I1346962,I1155002,I1155010,I1346977,I1155027,I1346965,I1155044,I1154899,I1155084,I1154920,I1155106,I1346974,I1155123,I1155149,I1155157,I1155174,I1346983,I1155191,I1155208,I1155225,I1154896,I1154917,I1155270,I1346986,I1154908,I1155301,I1155318,I1346980,I1346968,I1155344,I1155352,I1154914,I1155383,I1155400,I1155417,I1155434,I1154905,I1154902,I1155506,I1155532,I1155540,I1155580,I1155588,I1155605,I1155622,I1155662,I1155684,I1155701,I1155727,I1155735,I1155752,I1155769,I1155786,I1155803,I1155848,I1155879,I1155896,I1155922,I1155930,I1155961,I1155978,I1155995,I1156012,I1156084,I1156110,I1156118,I1156158,I1156166,I1156183,I1156200,I1156240,I1156262,I1156279,I1156305,I1156313,I1156330,I1156347,I1156364,I1156381,I1156426,I1156457,I1156474,I1156500,I1156508,I1156539,I1156556,I1156573,I1156590,I1156662,I1156688,I1156696,I1156736,I1156744,I1156761,I1156778,I1156818,I1156840,I1156857,I1156883,I1156891,I1156908,I1156925,I1156942,I1156959,I1157004,I1157035,I1157052,I1157078,I1157086,I1157117,I1157134,I1157151,I1157168,I1157240,I1157266,I1157274,I1157314,I1157322,I1157339,I1157356,I1157396,I1157418,I1157435,I1157461,I1157469,I1157486,I1157503,I1157520,I1157537,I1157582,I1157613,I1157630,I1157656,I1157664,I1157695,I1157712,I1157729,I1157746,I1157818,I1157844,I1157852,I1157892,I1157900,I1157917,I1157934,I1157974,I1157996,I1158013,I1158039,I1158047,I1158064,I1158081,I1158098,I1158115,I1158160,I1158191,I1158208,I1158234,I1158242,I1158273,I1158290,I1158307,I1158324,I1158396,I1248791,I1158422,I1158430,I1248785,I1248770,I1158470,I1158478,I1248776,I1158495,I1248788,I1158512,I1158552,I1158574,I1158591,I1158617,I1158625,I1158642,I1248794,I1158659,I1248782,I1158676,I1158693,I1158738,I1248773,I1158769,I1158786,I1248779,I1158812,I1158820,I1158851,I1158868,I1158885,I1158902,I1158974,I1159000,I1159008,I1158957,I1159048,I1159056,I1159073,I1159090,I1158945,I1159130,I1158966,I1159152,I1159169,I1159195,I1159203,I1159220,I1159237,I1159254,I1159271,I1158942,I1158963,I1159316,I1158954,I1159347,I1159364,I1159390,I1159398,I1158960,I1159429,I1159446,I1159463,I1159480,I1158951,I1158948,I1159552,I1159578,I1159586,I1159535,I1159626,I1159634,I1159651,I1159668,I1159523,I1159708,I1159544,I1159730,I1159747,I1159773,I1159781,I1159798,I1159815,I1159832,I1159849,I1159520,I1159541,I1159894,I1159532,I1159925,I1159942,I1159968,I1159976,I1159538,I1160007,I1160024,I1160041,I1160058,I1159529,I1159526,I1160130,I1160156,I1160164,I1160204,I1160212,I1160229,I1160246,I1160286,I1160308,I1160325,I1160351,I1160359,I1160376,I1160393,I1160410,I1160427,I1160472,I1160503,I1160520,I1160546,I1160554,I1160585,I1160602,I1160619,I1160636,I1160708,I1160734,I1160742,I1160782,I1160790,I1160807,I1160824,I1160864,I1160886,I1160903,I1160929,I1160937,I1160954,I1160971,I1160988,I1161005,I1161050,I1161081,I1161098,I1161124,I1161132,I1161163,I1161180,I1161197,I1161214,I1161286,I1161312,I1161320,I1161269,I1161360,I1161368,I1161385,I1161402,I1161257,I1161442,I1161278,I1161464,I1161481,I1161507,I1161515,I1161532,I1161549,I1161566,I1161583,I1161254,I1161275,I1161628,I1161266,I1161659,I1161676,I1161702,I1161710,I1161272,I1161741,I1161758,I1161775,I1161792,I1161263,I1161260,I1161864,I1161890,I1161898,I1161938,I1161946,I1161963,I1161980,I1162020,I1162042,I1162059,I1162085,I1162093,I1162110,I1162127,I1162144,I1162161,I1162206,I1162237,I1162254,I1162280,I1162288,I1162319,I1162336,I1162353,I1162370,I1162442,I1162468,I1162476,I1162516,I1162524,I1162541,I1162558,I1162598,I1162620,I1162637,I1162663,I1162671,I1162688,I1162705,I1162722,I1162739,I1162784,I1162815,I1162832,I1162858,I1162866,I1162897,I1162914,I1162931,I1162948,I1163020,I1163046,I1163054,I1163094,I1163102,I1163119,I1163136,I1163176,I1163198,I1163215,I1163241,I1163249,I1163266,I1163283,I1163300,I1163317,I1163362,I1163393,I1163410,I1163436,I1163444,I1163475,I1163492,I1163509,I1163526,I1163598,I1232471,I1163624,I1163632,I1232465,I1232450,I1163672,I1163680,I1232456,I1163697,I1232468,I1163714,I1163754,I1163776,I1163793,I1163819,I1163827,I1163844,I1232474,I1163861,I1232462,I1163878,I1163895,I1163940,I1232453,I1163971,I1163988,I1232459,I1164014,I1164022,I1164053,I1164070,I1164087,I1164104,I1164176,I1164202,I1164210,I1164250,I1164258,I1164275,I1164292,I1164332,I1164354,I1164371,I1164397,I1164405,I1164422,I1164439,I1164456,I1164473,I1164518,I1164549,I1164566,I1164592,I1164600,I1164631,I1164648,I1164665,I1164682,I1164754,I1299736,I1164780,I1164788,I1299763,I1299745,I1164828,I1164836,I1299754,I1164853,I1299757,I1164870,I1164910,I1164932,I1299751,I1164949,I1164975,I1164983,I1165000,I1299739,I1165017,I1299742,I1165034,I1165051,I1165096,I1299760,I1165127,I1165144,I1299748,I1165170,I1165178,I1165209,I1165226,I1165243,I1165260,I1165332,I1165358,I1165366,I1165406,I1165414,I1165431,I1165448,I1165488,I1165510,I1165527,I1165553,I1165561,I1165578,I1165595,I1165612,I1165629,I1165674,I1165705,I1165722,I1165748,I1165756,I1165787,I1165804,I1165821,I1165838,I1165910,I1165936,I1165944,I1165984,I1165992,I1166009,I1166026,I1166066,I1166088,I1166105,I1166131,I1166139,I1166156,I1166173,I1166190,I1166207,I1166252,I1166283,I1166300,I1166326,I1166334,I1166365,I1166382,I1166399,I1166416,I1166488,I1166514,I1166522,I1166562,I1166570,I1166587,I1166604,I1166644,I1166666,I1166683,I1166709,I1166717,I1166734,I1166751,I1166768,I1166785,I1166830,I1166861,I1166878,I1166904,I1166912,I1166943,I1166960,I1166977,I1166994,I1167066,I1167092,I1167100,I1167140,I1167148,I1167165,I1167182,I1167222,I1167244,I1167261,I1167287,I1167295,I1167312,I1167329,I1167346,I1167363,I1167408,I1167439,I1167456,I1167482,I1167490,I1167521,I1167538,I1167555,I1167572,I1167644,I1167670,I1167678,I1167718,I1167726,I1167743,I1167760,I1167800,I1167822,I1167839,I1167865,I1167873,I1167890,I1167907,I1167924,I1167941,I1167986,I1168017,I1168034,I1168060,I1168068,I1168099,I1168116,I1168133,I1168150,I1168222,I1168248,I1168256,I1168296,I1168304,I1168321,I1168338,I1168378,I1168400,I1168417,I1168443,I1168451,I1168468,I1168485,I1168502,I1168519,I1168564,I1168595,I1168612,I1168638,I1168646,I1168677,I1168694,I1168711,I1168728,I1168800,I1168826,I1168834,I1168874,I1168882,I1168899,I1168916,I1168956,I1168978,I1168995,I1169021,I1169029,I1169046,I1169063,I1169080,I1169097,I1169142,I1169173,I1169190,I1169216,I1169224,I1169255,I1169272,I1169289,I1169306,I1169378,I1169404,I1169412,I1169452,I1169460,I1169477,I1169494,I1169534,I1169556,I1169573,I1169599,I1169607,I1169624,I1169641,I1169658,I1169675,I1169720,I1169751,I1169768,I1169794,I1169802,I1169833,I1169850,I1169867,I1169884,I1169956,I1169982,I1169990,I1170030,I1170038,I1170055,I1170072,I1170112,I1170134,I1170151,I1170177,I1170185,I1170202,I1170219,I1170236,I1170253,I1170298,I1170329,I1170346,I1170372,I1170380,I1170411,I1170428,I1170445,I1170462,I1170534,I1170560,I1170568,I1170608,I1170616,I1170633,I1170650,I1170690,I1170712,I1170729,I1170755,I1170763,I1170780,I1170797,I1170814,I1170831,I1170876,I1170907,I1170924,I1170950,I1170958,I1170989,I1171006,I1171023,I1171040,I1171112,I1171138,I1171146,I1171186,I1171194,I1171211,I1171228,I1171268,I1171290,I1171307,I1171333,I1171341,I1171358,I1171375,I1171392,I1171409,I1171454,I1171485,I1171502,I1171528,I1171536,I1171567,I1171584,I1171601,I1171618,I1171690,I1171716,I1171724,I1171764,I1171772,I1171789,I1171806,I1171846,I1171868,I1171885,I1171911,I1171919,I1171936,I1171953,I1171970,I1171987,I1172032,I1172063,I1172080,I1172106,I1172114,I1172145,I1172162,I1172179,I1172196,I1172268,I1344014,I1172294,I1172302,I1343996,I1172251,I1343987,I1172342,I1172350,I1344002,I1172367,I1343990,I1172384,I1172239,I1172424,I1172260,I1172446,I1343999,I1172463,I1172489,I1172497,I1172514,I1344008,I1172531,I1172548,I1172565,I1172236,I1172257,I1172610,I1344011,I1172248,I1172641,I1172658,I1344005,I1343993,I1172684,I1172692,I1172254,I1172723,I1172740,I1172757,I1172774,I1172245,I1172242,I1172846,I1172872,I1172880,I1172920,I1172928,I1172945,I1172962,I1173002,I1173024,I1173041,I1173067,I1173075,I1173092,I1173109,I1173126,I1173143,I1173188,I1173219,I1173236,I1173262,I1173270,I1173301,I1173318,I1173335,I1173352,I1173424,I1173450,I1173458,I1173498,I1173506,I1173523,I1173540,I1173580,I1173602,I1173619,I1173645,I1173653,I1173670,I1173687,I1173704,I1173721,I1173766,I1173797,I1173814,I1173840,I1173848,I1173879,I1173896,I1173913,I1173930,I1174002,I1174028,I1174036,I1174076,I1174084,I1174101,I1174118,I1174158,I1174180,I1174197,I1174223,I1174231,I1174248,I1174265,I1174282,I1174299,I1174344,I1174375,I1174392,I1174418,I1174426,I1174457,I1174474,I1174491,I1174508,I1174580,I1252055,I1174606,I1174614,I1252049,I1174563,I1252034,I1174654,I1174662,I1252040,I1174679,I1252052,I1174696,I1174551,I1174736,I1174572,I1174758,I1174775,I1174801,I1174809,I1174826,I1252058,I1174843,I1252046,I1174860,I1174877,I1174548,I1174569,I1174922,I1252037,I1174560,I1174953,I1174970,I1252043,I1174996,I1175004,I1174566,I1175035,I1175052,I1175069,I1175086,I1174557,I1174554,I1175158,I1175184,I1175192,I1175232,I1175240,I1175257,I1175274,I1175314,I1175336,I1175353,I1175379,I1175387,I1175404,I1175421,I1175438,I1175455,I1175500,I1175531,I1175548,I1175574,I1175582,I1175613,I1175630,I1175647,I1175664,I1175736,I1175762,I1175770,I1175810,I1175818,I1175835,I1175852,I1175892,I1175914,I1175931,I1175957,I1175965,I1175982,I1175999,I1176016,I1176033,I1176078,I1176109,I1176126,I1176152,I1176160,I1176191,I1176208,I1176225,I1176242,I1176314,I1176340,I1176348,I1176297,I1176388,I1176396,I1176413,I1176430,I1176285,I1176470,I1176306,I1176492,I1176509,I1176535,I1176543,I1176560,I1176577,I1176594,I1176611,I1176282,I1176303,I1176656,I1176294,I1176687,I1176704,I1176730,I1176738,I1176300,I1176769,I1176786,I1176803,I1176820,I1176291,I1176288,I1176892,I1176918,I1176926,I1176966,I1176974,I1176991,I1177008,I1177048,I1177070,I1177087,I1177113,I1177121,I1177138,I1177155,I1177172,I1177189,I1177234,I1177265,I1177282,I1177308,I1177316,I1177347,I1177364,I1177381,I1177398,I1177470,I1177496,I1177504,I1177544,I1177552,I1177569,I1177586,I1177626,I1177648,I1177665,I1177691,I1177699,I1177716,I1177733,I1177750,I1177767,I1177812,I1177843,I1177860,I1177886,I1177894,I1177925,I1177942,I1177959,I1177976,I1178048,I1178074,I1178082,I1178122,I1178130,I1178147,I1178164,I1178204,I1178226,I1178243,I1178269,I1178277,I1178294,I1178311,I1178328,I1178345,I1178390,I1178421,I1178438,I1178464,I1178472,I1178503,I1178520,I1178537,I1178554,I1178626,I1178652,I1178660,I1178700,I1178708,I1178725,I1178742,I1178782,I1178804,I1178821,I1178847,I1178855,I1178872,I1178889,I1178906,I1178923,I1178968,I1178999,I1179016,I1179042,I1179050,I1179081,I1179098,I1179115,I1179132,I1179204,I1179230,I1179238,I1179278,I1179286,I1179303,I1179320,I1179360,I1179382,I1179399,I1179425,I1179433,I1179450,I1179467,I1179484,I1179501,I1179546,I1179577,I1179594,I1179620,I1179628,I1179659,I1179676,I1179693,I1179710,I1179782,I1179808,I1179816,I1179856,I1179864,I1179881,I1179898,I1179938,I1179960,I1179977,I1180003,I1180011,I1180028,I1180045,I1180062,I1180079,I1180124,I1180155,I1180172,I1180198,I1180206,I1180237,I1180254,I1180271,I1180288,I1180360,I1180386,I1180394,I1180434,I1180442,I1180459,I1180476,I1180516,I1180538,I1180555,I1180581,I1180589,I1180606,I1180623,I1180640,I1180657,I1180702,I1180733,I1180750,I1180776,I1180784,I1180815,I1180832,I1180849,I1180866,I1180938,I1180964,I1180972,I1180921,I1181012,I1181020,I1181037,I1181054,I1180909,I1181094,I1180930,I1181116,I1181133,I1181159,I1181167,I1181184,I1181201,I1181218,I1181235,I1180906,I1180927,I1181280,I1180918,I1181311,I1181328,I1181354,I1181362,I1180924,I1181393,I1181410,I1181427,I1181444,I1180915,I1180912,I1181516,I1181542,I1181550,I1181590,I1181598,I1181615,I1181632,I1181672,I1181694,I1181711,I1181737,I1181745,I1181762,I1181779,I1181796,I1181813,I1181858,I1181889,I1181906,I1181932,I1181940,I1181971,I1181988,I1182005,I1182022,I1182094,I1182120,I1182128,I1182168,I1182176,I1182193,I1182210,I1182250,I1182272,I1182289,I1182315,I1182323,I1182340,I1182357,I1182374,I1182391,I1182436,I1182467,I1182484,I1182510,I1182518,I1182549,I1182566,I1182583,I1182600,I1182672,I1182698,I1182706,I1182746,I1182754,I1182771,I1182788,I1182828,I1182850,I1182867,I1182893,I1182901,I1182918,I1182935,I1182952,I1182969,I1183014,I1183045,I1183062,I1183088,I1183096,I1183127,I1183144,I1183161,I1183178,I1183250,I1183276,I1183284,I1183324,I1183332,I1183349,I1183366,I1183406,I1183428,I1183445,I1183471,I1183479,I1183496,I1183513,I1183530,I1183547,I1183592,I1183623,I1183640,I1183666,I1183674,I1183705,I1183722,I1183739,I1183756,I1183828,I1183854,I1183862,I1183902,I1183910,I1183927,I1183944,I1183984,I1184006,I1184023,I1184049,I1184057,I1184074,I1184091,I1184108,I1184125,I1184170,I1184201,I1184218,I1184244,I1184252,I1184283,I1184300,I1184317,I1184334,I1184406,I1184432,I1184440,I1184480,I1184488,I1184505,I1184522,I1184562,I1184584,I1184601,I1184627,I1184635,I1184652,I1184669,I1184686,I1184703,I1184748,I1184779,I1184796,I1184822,I1184830,I1184861,I1184878,I1184895,I1184912,I1184984,I1185010,I1185018,I1185058,I1185066,I1185083,I1185100,I1185140,I1185162,I1185179,I1185205,I1185213,I1185230,I1185247,I1185264,I1185281,I1185326,I1185357,I1185374,I1185400,I1185408,I1185439,I1185456,I1185473,I1185490,I1185562,I1185588,I1185596,I1185636,I1185644,I1185661,I1185678,I1185718,I1185740,I1185757,I1185783,I1185791,I1185808,I1185825,I1185842,I1185859,I1185904,I1185935,I1185952,I1185978,I1185986,I1186017,I1186034,I1186051,I1186068,I1186140,I1186166,I1186174,I1186123,I1186214,I1186222,I1186239,I1186256,I1186111,I1186296,I1186132,I1186318,I1186335,I1186361,I1186369,I1186386,I1186403,I1186420,I1186437,I1186108,I1186129,I1186482,I1186120,I1186513,I1186530,I1186556,I1186564,I1186126,I1186595,I1186612,I1186629,I1186646,I1186117,I1186114,I1186718,I1307719,I1186744,I1186752,I1307701,I1307692,I1186792,I1186800,I1307707,I1186817,I1307695,I1186834,I1186874,I1186896,I1307704,I1186913,I1186939,I1186947,I1186964,I1307713,I1186981,I1186998,I1187015,I1187060,I1307716,I1187091,I1187108,I1307710,I1307698,I1187134,I1187142,I1187173,I1187190,I1187207,I1187224,I1187296,I1187322,I1187330,I1187279,I1187370,I1187378,I1187395,I1187412,I1187267,I1187452,I1187288,I1187474,I1187491,I1187517,I1187525,I1187542,I1187559,I1187576,I1187593,I1187264,I1187285,I1187638,I1187276,I1187669,I1187686,I1187712,I1187720,I1187282,I1187751,I1187768,I1187785,I1187802,I1187273,I1187270,I1187874,I1187900,I1187908,I1187857,I1187948,I1187956,I1187973,I1187990,I1187845,I1188030,I1187866,I1188052,I1188069,I1188095,I1188103,I1188120,I1188137,I1188154,I1188171,I1187842,I1187863,I1188216,I1187854,I1188247,I1188264,I1188290,I1188298,I1187860,I1188329,I1188346,I1188363,I1188380,I1187851,I1187848,I1188452,I1235191,I1188478,I1188486,I1235185,I1235170,I1188526,I1188534,I1235176,I1188551,I1235188,I1188568,I1188608,I1188630,I1188647,I1188673,I1188681,I1188698,I1235194,I1188715,I1235182,I1188732,I1188749,I1188794,I1235173,I1188825,I1188842,I1235179,I1188868,I1188876,I1188907,I1188924,I1188941,I1188958,I1189030,I1189056,I1189064,I1189104,I1189112,I1189129,I1189146,I1189186,I1189208,I1189225,I1189251,I1189259,I1189276,I1189293,I1189310,I1189327,I1189372,I1189403,I1189420,I1189446,I1189454,I1189485,I1189502,I1189519,I1189536,I1189608,I1189634,I1189642,I1189682,I1189690,I1189707,I1189724,I1189764,I1189786,I1189803,I1189829,I1189837,I1189854,I1189871,I1189888,I1189905,I1189950,I1189981,I1189998,I1190024,I1190032,I1190063,I1190080,I1190097,I1190114,I1190186,I1190212,I1190220,I1190260,I1190268,I1190285,I1190302,I1190342,I1190364,I1190381,I1190407,I1190415,I1190432,I1190449,I1190466,I1190483,I1190528,I1190559,I1190576,I1190602,I1190610,I1190641,I1190658,I1190675,I1190692,I1190764,I1190790,I1190798,I1190838,I1190846,I1190863,I1190880,I1190920,I1190942,I1190959,I1190985,I1190993,I1191010,I1191027,I1191044,I1191061,I1191106,I1191137,I1191154,I1191180,I1191188,I1191219,I1191236,I1191253,I1191270,I1191342,I1247159,I1191368,I1191376,I1247153,I1191325,I1247138,I1191416,I1191424,I1247144,I1191441,I1247156,I1191458,I1191313,I1191498,I1191334,I1191520,I1191537,I1191563,I1191571,I1191588,I1247162,I1191605,I1247150,I1191622,I1191639,I1191310,I1191331,I1191684,I1247141,I1191322,I1191715,I1191732,I1247147,I1191758,I1191766,I1191328,I1191797,I1191814,I1191831,I1191848,I1191319,I1191316,I1191920,I1191946,I1191954,I1191994,I1192002,I1192019,I1192036,I1192076,I1192098,I1192115,I1192141,I1192149,I1192166,I1192183,I1192200,I1192217,I1192262,I1192293,I1192310,I1192336,I1192344,I1192375,I1192392,I1192409,I1192426,I1192498,I1192524,I1192532,I1192572,I1192580,I1192597,I1192614,I1192654,I1192676,I1192693,I1192719,I1192727,I1192744,I1192761,I1192778,I1192795,I1192840,I1192871,I1192888,I1192914,I1192922,I1192953,I1192970,I1192987,I1193004,I1193076,I1193102,I1193110,I1193150,I1193158,I1193175,I1193192,I1193232,I1193254,I1193271,I1193297,I1193305,I1193322,I1193339,I1193356,I1193373,I1193418,I1193449,I1193466,I1193492,I1193500,I1193531,I1193548,I1193565,I1193582,I1193654,I1193680,I1193688,I1193728,I1193736,I1193753,I1193770,I1193810,I1193832,I1193849,I1193875,I1193883,I1193900,I1193917,I1193934,I1193951,I1193996,I1194027,I1194044,I1194070,I1194078,I1194109,I1194126,I1194143,I1194160,I1194232,I1194258,I1194266,I1194215,I1194306,I1194314,I1194331,I1194348,I1194203,I1194388,I1194224,I1194410,I1194427,I1194453,I1194461,I1194478,I1194495,I1194512,I1194529,I1194200,I1194221,I1194574,I1194212,I1194605,I1194622,I1194648,I1194656,I1194218,I1194687,I1194704,I1194721,I1194738,I1194209,I1194206,I1194810,I1194836,I1194844,I1194884,I1194892,I1194909,I1194926,I1194966,I1194988,I1195005,I1195031,I1195039,I1195056,I1195073,I1195090,I1195107,I1195152,I1195183,I1195200,I1195226,I1195234,I1195265,I1195282,I1195299,I1195316,I1195388,I1277898,I1195414,I1195422,I1277880,I1277889,I1195462,I1195470,I1277874,I1195487,I1277886,I1195504,I1195544,I1195566,I1277877,I1195583,I1195609,I1195617,I1195634,I1195651,I1195668,I1195685,I1195730,I1277895,I1195761,I1195778,I1277883,I1277892,I1195804,I1195812,I1195843,I1195860,I1195877,I1195894,I1195966,I1195992,I1196000,I1196040,I1196048,I1196065,I1196082,I1196122,I1196144,I1196161,I1196187,I1196195,I1196212,I1196229,I1196246,I1196263,I1196308,I1196339,I1196356,I1196382,I1196390,I1196421,I1196438,I1196455,I1196472,I1196544,I1196570,I1196578,I1196527,I1196618,I1196626,I1196643,I1196660,I1196515,I1196700,I1196536,I1196722,I1196739,I1196765,I1196773,I1196790,I1196807,I1196824,I1196841,I1196512,I1196533,I1196886,I1196524,I1196917,I1196934,I1196960,I1196968,I1196530,I1196999,I1197016,I1197033,I1197050,I1196521,I1196518,I1197122,I1197148,I1197156,I1197196,I1197204,I1197221,I1197238,I1197278,I1197300,I1197317,I1197343,I1197351,I1197368,I1197385,I1197402,I1197419,I1197464,I1197495,I1197512,I1197538,I1197546,I1197577,I1197594,I1197611,I1197628,I1197700,I1197726,I1197734,I1197774,I1197782,I1197799,I1197816,I1197856,I1197878,I1197895,I1197921,I1197929,I1197946,I1197963,I1197980,I1197997,I1198042,I1198073,I1198090,I1198116,I1198124,I1198155,I1198172,I1198189,I1198206,I1198278,I1250423,I1198304,I1198312,I1250417,I1250402,I1198352,I1198360,I1250408,I1198377,I1250420,I1198394,I1198434,I1198456,I1198473,I1198499,I1198507,I1198524,I1250426,I1198541,I1250414,I1198558,I1198575,I1198620,I1250405,I1198651,I1198668,I1250411,I1198694,I1198702,I1198733,I1198750,I1198767,I1198784,I1198856,I1198882,I1198890,I1198930,I1198938,I1198955,I1198972,I1199012,I1199034,I1199051,I1199077,I1199085,I1199102,I1199119,I1199136,I1199153,I1199198,I1199229,I1199246,I1199272,I1199280,I1199311,I1199328,I1199345,I1199362,I1199434,I1199460,I1199468,I1199508,I1199516,I1199533,I1199550,I1199590,I1199612,I1199629,I1199655,I1199663,I1199680,I1199697,I1199714,I1199731,I1199776,I1199807,I1199824,I1199850,I1199858,I1199889,I1199906,I1199923,I1199940,I1200012,I1346394,I1200038,I1200046,I1346376,I1346367,I1200086,I1200094,I1346382,I1200111,I1346370,I1200128,I1200168,I1200190,I1346379,I1200207,I1200233,I1200241,I1200258,I1346388,I1200275,I1200292,I1200309,I1200354,I1346391,I1200385,I1200402,I1346385,I1346373,I1200428,I1200436,I1200467,I1200484,I1200501,I1200518,I1200590,I1200616,I1200624,I1200664,I1200672,I1200689,I1200706,I1200746,I1200768,I1200785,I1200811,I1200819,I1200836,I1200853,I1200870,I1200887,I1200932,I1200963,I1200980,I1201006,I1201014,I1201045,I1201062,I1201079,I1201096,I1201168,I1210167,I1201194,I1201202,I1210161,I1210146,I1201242,I1201250,I1210152,I1201267,I1210164,I1201284,I1201324,I1201346,I1201363,I1201389,I1201397,I1201414,I1210170,I1201431,I1210158,I1201448,I1201465,I1201510,I1210149,I1201541,I1201558,I1210155,I1201584,I1201592,I1201623,I1201640,I1201657,I1201674,I1201746,I1201772,I1201780,I1201820,I1201828,I1201845,I1201862,I1201902,I1201924,I1201941,I1201967,I1201975,I1201992,I1202009,I1202026,I1202043,I1202088,I1202119,I1202136,I1202162,I1202170,I1202201,I1202218,I1202235,I1202252,I1202324,I1202350,I1202358,I1202307,I1202398,I1202406,I1202423,I1202440,I1202295,I1202480,I1202316,I1202502,I1202519,I1202545,I1202553,I1202570,I1202587,I1202604,I1202621,I1202292,I1202313,I1202666,I1202304,I1202697,I1202714,I1202740,I1202748,I1202310,I1202779,I1202796,I1202813,I1202830,I1202301,I1202298,I1202902,I1202928,I1202936,I1202976,I1202984,I1203001,I1203018,I1203058,I1203080,I1203097,I1203123,I1203131,I1203148,I1203165,I1203182,I1203199,I1203244,I1203275,I1203292,I1203318,I1203326,I1203357,I1203374,I1203391,I1203408,I1203480,I1203506,I1203514,I1203554,I1203562,I1203579,I1203596,I1203636,I1203658,I1203675,I1203701,I1203709,I1203726,I1203743,I1203760,I1203777,I1203822,I1203853,I1203870,I1203896,I1203904,I1203935,I1203952,I1203969,I1203986,I1204058,I1204084,I1204092,I1204132,I1204140,I1204157,I1204174,I1204214,I1204236,I1204253,I1204279,I1204287,I1204304,I1204321,I1204338,I1204355,I1204400,I1204431,I1204448,I1204474,I1204482,I1204513,I1204530,I1204547,I1204564,I1204636,I1204662,I1204670,I1204710,I1204718,I1204735,I1204752,I1204792,I1204814,I1204831,I1204857,I1204865,I1204882,I1204899,I1204916,I1204933,I1204978,I1205009,I1205026,I1205052,I1205060,I1205091,I1205108,I1205125,I1205142,I1205214,I1253143,I1205240,I1205248,I1253137,I1205197,I1253122,I1205288,I1205296,I1253128,I1205313,I1253140,I1205330,I1205185,I1205370,I1205206,I1205392,I1205409,I1205435,I1205443,I1205460,I1253146,I1205477,I1253134,I1205494,I1205511,I1205182,I1205203,I1205556,I1253125,I1205194,I1205587,I1205604,I1253131,I1205630,I1205638,I1205200,I1205669,I1205686,I1205703,I1205720,I1205191,I1205188,I1205792,I1205818,I1205826,I1205866,I1205874,I1205891,I1205908,I1205948,I1205970,I1205987,I1206013,I1206021,I1206038,I1206055,I1206072,I1206089,I1206134,I1206165,I1206182,I1206208,I1206216,I1206247,I1206264,I1206281,I1206298,I1206370,I1206396,I1206404,I1206430,I1206447,I1206469,I1206486,I1206503,I1206520,I1206537,I1206568,I1206585,I1206602,I1206619,I1206664,I1206681,I1206698,I1206757,I1206783,I1206791,I1206808,I1206825,I1206856,I1206914,I1316049,I1206940,I1206948,I1316034,I1316028,I1206974,I1206991,I1207013,I1316022,I1207030,I1316043,I1207047,I1316031,I1207064,I1207081,I1207112,I1316040,I1207129,I1316046,I1207146,I1316037,I1207163,I1207208,I1316025,I1207225,I1207242,I1207301,I1207327,I1207335,I1207352,I1207369,I1207400,I1207458,I1207484,I1207492,I1207518,I1207535,I1207557,I1207574,I1207591,I1207608,I1207625,I1207656,I1207673,I1207690,I1207707,I1207752,I1207769,I1207786,I1207845,I1207871,I1207879,I1207896,I1207913,I1207944,I1208002,I1369599,I1208028,I1208036,I1369584,I1369578,I1208062,I1208079,I1208101,I1369572,I1208118,I1369593,I1208135,I1369581,I1208152,I1208169,I1208200,I1369590,I1208217,I1369596,I1208234,I1369587,I1208251,I1208296,I1369575,I1208313,I1208330,I1208389,I1208415,I1208423,I1208440,I1208457,I1208488,I1208546,I1208572,I1208580,I1208606,I1208623,I1208645,I1208662,I1208679,I1208696,I1208713,I1208744,I1208761,I1208778,I1208795,I1208840,I1208857,I1208874,I1208933,I1208959,I1208967,I1208984,I1209001,I1209032,I1209090,I1209116,I1209124,I1209150,I1209167,I1209189,I1209206,I1209223,I1209240,I1209257,I1209288,I1209305,I1209322,I1209339,I1209384,I1209401,I1209418,I1209477,I1209503,I1209511,I1209528,I1209545,I1209576,I1209634,I1209660,I1209668,I1209694,I1209711,I1209733,I1209750,I1209767,I1209784,I1209801,I1209832,I1209849,I1209866,I1209883,I1209928,I1209945,I1209962,I1210021,I1210047,I1210055,I1210072,I1210089,I1210120,I1210178,I1210204,I1210212,I1210238,I1210255,I1210277,I1210294,I1210311,I1210328,I1210345,I1210376,I1210393,I1210410,I1210427,I1210472,I1210489,I1210506,I1210565,I1210591,I1210599,I1210616,I1210633,I1210664,I1210722,I1210748,I1210756,I1210782,I1210799,I1210821,I1210838,I1210855,I1210872,I1210889,I1210920,I1210937,I1210954,I1210971,I1211016,I1211033,I1211050,I1211109,I1211135,I1211143,I1211160,I1211177,I1211208,I1211266,I1211292,I1211300,I1211326,I1211343,I1211258,I1211365,I1211382,I1211399,I1211416,I1211433,I1211237,I1211464,I1211481,I1211498,I1211515,I1211240,I1211255,I1211560,I1211577,I1211594,I1211252,I1211249,I1211246,I1211653,I1211679,I1211687,I1211704,I1211721,I1211234,I1211752,I1211243,I1211810,I1211836,I1211844,I1211870,I1211887,I1211909,I1211926,I1211943,I1211960,I1211977,I1212008,I1212025,I1212042,I1212059,I1212104,I1212121,I1212138,I1212197,I1212223,I1212231,I1212248,I1212265,I1212296,I1212354,I1212380,I1212388,I1212414,I1212431,I1212453,I1212470,I1212487,I1212504,I1212521,I1212552,I1212569,I1212586,I1212603,I1212648,I1212665,I1212682,I1212741,I1212767,I1212775,I1212792,I1212809,I1212840,I1212898,I1212924,I1212932,I1212958,I1212975,I1212997,I1213014,I1213031,I1213048,I1213065,I1213096,I1213113,I1213130,I1213147,I1213192,I1213209,I1213226,I1213285,I1213311,I1213319,I1213336,I1213353,I1213384,I1213442,I1213468,I1213476,I1213502,I1213519,I1213541,I1213558,I1213575,I1213592,I1213609,I1213640,I1213657,I1213674,I1213691,I1213736,I1213753,I1213770,I1213829,I1213855,I1213863,I1213880,I1213897,I1213928,I1213986,I1352344,I1214012,I1214020,I1352329,I1352323,I1214046,I1214063,I1214085,I1352317,I1214102,I1352338,I1214119,I1352326,I1214136,I1214153,I1214184,I1352335,I1214201,I1352341,I1214218,I1352332,I1214235,I1214280,I1352320,I1214297,I1214314,I1214373,I1214399,I1214407,I1214424,I1214441,I1214472,I1214530,I1214556,I1214564,I1214590,I1214607,I1214629,I1214646,I1214663,I1214680,I1214697,I1214728,I1214745,I1214762,I1214779,I1214824,I1214841,I1214858,I1214917,I1214943,I1214951,I1214968,I1214985,I1215016,I1215074,I1215100,I1215108,I1215134,I1215151,I1215173,I1215190,I1215207,I1215224,I1215241,I1215272,I1215289,I1215306,I1215323,I1215368,I1215385,I1215402,I1215461,I1215487,I1215495,I1215512,I1215529,I1215560,I1215618,I1215644,I1215652,I1215678,I1215695,I1215717,I1215734,I1215751,I1215768,I1215785,I1215816,I1215833,I1215850,I1215867,I1215912,I1215929,I1215946,I1216005,I1216031,I1216039,I1216056,I1216073,I1216104,I1216162,I1216188,I1216196,I1216222,I1216239,I1216261,I1216278,I1216295,I1216312,I1216329,I1216360,I1216377,I1216394,I1216411,I1216456,I1216473,I1216490,I1216549,I1216575,I1216583,I1216600,I1216617,I1216648,I1216706,I1216732,I1216740,I1216766,I1216783,I1216698,I1216805,I1216822,I1216839,I1216856,I1216873,I1216677,I1216904,I1216921,I1216938,I1216955,I1216680,I1216695,I1217000,I1217017,I1217034,I1216692,I1216689,I1216686,I1217093,I1217119,I1217127,I1217144,I1217161,I1216674,I1217192,I1216683,I1217250,I1217276,I1217284,I1217310,I1217327,I1217349,I1217366,I1217383,I1217400,I1217417,I1217448,I1217465,I1217482,I1217499,I1217544,I1217561,I1217578,I1217637,I1217663,I1217671,I1217688,I1217705,I1217736,I1217794,I1294067,I1217820,I1217828,I1294076,I1294079,I1217854,I1217871,I1217893,I1294073,I1217910,I1294070,I1217927,I1294064,I1217944,I1217961,I1217992,I1294061,I1218009,I1294058,I1218026,I1218043,I1218088,I1218105,I1218122,I1218181,I1294082,I1218207,I1218215,I1218232,I1218249,I1218280,I1218338,I1305934,I1218364,I1218372,I1305919,I1305913,I1218398,I1218415,I1218437,I1305907,I1218454,I1305928,I1218471,I1305916,I1218488,I1218505,I1218536,I1305925,I1218553,I1305931,I1218570,I1305922,I1218587,I1218632,I1305910,I1218649,I1218666,I1218725,I1218751,I1218759,I1218776,I1218793,I1218824,I1218882,I1218908,I1218916,I1218942,I1218959,I1218981,I1218998,I1219015,I1219032,I1219049,I1219080,I1219097,I1219114,I1219131,I1219176,I1219193,I1219210,I1219269,I1219295,I1219303,I1219320,I1219337,I1219368,I1219426,I1219452,I1219460,I1219486,I1219503,I1219525,I1219542,I1219559,I1219576,I1219593,I1219624,I1219641,I1219658,I1219675,I1219720,I1219737,I1219754,I1219813,I1219839,I1219847,I1219864,I1219881,I1219912,I1219970,I1219996,I1220004,I1220030,I1220047,I1220069,I1220086,I1220103,I1220120,I1220137,I1220168,I1220185,I1220202,I1220219,I1220264,I1220281,I1220298,I1220357,I1220383,I1220391,I1220408,I1220425,I1220456,I1220514,I1270369,I1220540,I1220548,I1270378,I1270381,I1220574,I1220591,I1220613,I1270375,I1220630,I1270372,I1220647,I1270366,I1220664,I1220681,I1220712,I1270363,I1220729,I1270360,I1220746,I1220763,I1220808,I1220825,I1220842,I1220901,I1270384,I1220927,I1220935,I1220952,I1220969,I1221000,I1221058,I1221084,I1221092,I1221118,I1221135,I1221157,I1221174,I1221191,I1221208,I1221225,I1221256,I1221273,I1221290,I1221307,I1221352,I1221369,I1221386,I1221445,I1221471,I1221479,I1221496,I1221513,I1221544,I1221602,I1221628,I1221636,I1221662,I1221679,I1221701,I1221718,I1221735,I1221752,I1221769,I1221800,I1221817,I1221834,I1221851,I1221896,I1221913,I1221930,I1221989,I1222015,I1222023,I1222040,I1222057,I1222088,I1222146,I1222172,I1222180,I1222206,I1222223,I1222245,I1222262,I1222279,I1222296,I1222313,I1222344,I1222361,I1222378,I1222395,I1222440,I1222457,I1222474,I1222533,I1222559,I1222567,I1222584,I1222601,I1222632,I1222690,I1222716,I1222724,I1222750,I1222767,I1222789,I1222806,I1222823,I1222840,I1222857,I1222888,I1222905,I1222922,I1222939,I1222984,I1223001,I1223018,I1223077,I1223103,I1223111,I1223128,I1223145,I1223176,I1223234,I1223260,I1223268,I1223294,I1223311,I1223333,I1223350,I1223367,I1223384,I1223401,I1223432,I1223449,I1223466,I1223483,I1223528,I1223545,I1223562,I1223621,I1223647,I1223655,I1223672,I1223689,I1223720,I1223778,I1223804,I1223812,I1223838,I1223855,I1223877,I1223894,I1223911,I1223928,I1223945,I1223976,I1223993,I1224010,I1224027,I1224072,I1224089,I1224106,I1224165,I1224191,I1224199,I1224216,I1224233,I1224264,I1224322,I1224348,I1224356,I1224382,I1224399,I1224421,I1224438,I1224455,I1224472,I1224489,I1224520,I1224537,I1224554,I1224571,I1224616,I1224633,I1224650,I1224709,I1224735,I1224743,I1224760,I1224777,I1224808,I1224866,I1224892,I1224900,I1224926,I1224943,I1224858,I1224965,I1224982,I1224999,I1225016,I1225033,I1224837,I1225064,I1225081,I1225098,I1225115,I1224840,I1224855,I1225160,I1225177,I1225194,I1224852,I1224849,I1224846,I1225253,I1225279,I1225287,I1225304,I1225321,I1224834,I1225352,I1224843,I1225410,I1225436,I1225444,I1225470,I1225487,I1225509,I1225526,I1225543,I1225560,I1225577,I1225608,I1225625,I1225642,I1225659,I1225704,I1225721,I1225738,I1225797,I1225823,I1225831,I1225848,I1225865,I1225896,I1225954,I1225980,I1225988,I1226014,I1226031,I1226053,I1226070,I1226087,I1226104,I1226121,I1226152,I1226169,I1226186,I1226203,I1226248,I1226265,I1226282,I1226341,I1226367,I1226375,I1226392,I1226409,I1226440,I1226498,I1226524,I1226532,I1226558,I1226575,I1226597,I1226614,I1226631,I1226648,I1226665,I1226696,I1226713,I1226730,I1226747,I1226792,I1226809,I1226826,I1226885,I1226911,I1226919,I1226936,I1226953,I1226984,I1227042,I1227068,I1227076,I1227102,I1227119,I1227141,I1227158,I1227175,I1227192,I1227209,I1227240,I1227257,I1227274,I1227291,I1227336,I1227353,I1227370,I1227429,I1227455,I1227463,I1227480,I1227497,I1227528,I1227586,I1227612,I1227620,I1227646,I1227663,I1227685,I1227702,I1227719,I1227736,I1227753,I1227784,I1227801,I1227818,I1227835,I1227880,I1227897,I1227914,I1227973,I1227999,I1228007,I1228024,I1228041,I1228072,I1228130,I1228156,I1228164,I1228190,I1228207,I1228229,I1228246,I1228263,I1228280,I1228297,I1228328,I1228345,I1228362,I1228379,I1228424,I1228441,I1228458,I1228517,I1228543,I1228551,I1228568,I1228585,I1228616,I1228674,I1228700,I1228708,I1228734,I1228751,I1228773,I1228790,I1228807,I1228824,I1228841,I1228872,I1228889,I1228906,I1228923,I1228968,I1228985,I1229002,I1229061,I1229087,I1229095,I1229112,I1229129,I1229160,I1229218,I1229244,I1229252,I1229278,I1229295,I1229317,I1229334,I1229351,I1229368,I1229385,I1229416,I1229433,I1229450,I1229467,I1229512,I1229529,I1229546,I1229605,I1229631,I1229639,I1229656,I1229673,I1229704,I1229762,I1229788,I1229796,I1229822,I1229839,I1229861,I1229878,I1229895,I1229912,I1229929,I1229960,I1229977,I1229994,I1230011,I1230056,I1230073,I1230090,I1230149,I1230175,I1230183,I1230200,I1230217,I1230248,I1230306,I1230332,I1230340,I1230366,I1230383,I1230405,I1230422,I1230439,I1230456,I1230473,I1230504,I1230521,I1230538,I1230555,I1230600,I1230617,I1230634,I1230693,I1230719,I1230727,I1230744,I1230761,I1230792,I1230850,I1230876,I1230884,I1230910,I1230927,I1230949,I1230966,I1230983,I1231000,I1231017,I1231048,I1231065,I1231082,I1231099,I1231144,I1231161,I1231178,I1231237,I1231263,I1231271,I1231288,I1231305,I1231336,I1231394,I1231420,I1231428,I1231454,I1231471,I1231493,I1231510,I1231527,I1231544,I1231561,I1231592,I1231609,I1231626,I1231643,I1231688,I1231705,I1231722,I1231781,I1231807,I1231815,I1231832,I1231849,I1231880,I1231938,I1231964,I1231972,I1231998,I1232015,I1232037,I1232054,I1232071,I1232088,I1232105,I1232136,I1232153,I1232170,I1232187,I1232232,I1232249,I1232266,I1232325,I1232351,I1232359,I1232376,I1232393,I1232424,I1232482,I1232508,I1232516,I1232542,I1232559,I1232581,I1232598,I1232615,I1232632,I1232649,I1232680,I1232697,I1232714,I1232731,I1232776,I1232793,I1232810,I1232869,I1232895,I1232903,I1232920,I1232937,I1232968,I1233026,I1233052,I1233060,I1233086,I1233103,I1233125,I1233142,I1233159,I1233176,I1233193,I1233224,I1233241,I1233258,I1233275,I1233320,I1233337,I1233354,I1233413,I1233439,I1233447,I1233464,I1233481,I1233512,I1233570,I1233596,I1233604,I1233630,I1233647,I1233669,I1233686,I1233703,I1233720,I1233737,I1233768,I1233785,I1233802,I1233819,I1233864,I1233881,I1233898,I1233957,I1233983,I1233991,I1234008,I1234025,I1234056,I1234114,I1234140,I1234148,I1234174,I1234191,I1234213,I1234230,I1234247,I1234264,I1234281,I1234312,I1234329,I1234346,I1234363,I1234408,I1234425,I1234442,I1234501,I1234527,I1234535,I1234552,I1234569,I1234600,I1234658,I1234684,I1234692,I1234718,I1234735,I1234757,I1234774,I1234791,I1234808,I1234825,I1234856,I1234873,I1234890,I1234907,I1234952,I1234969,I1234986,I1235045,I1235071,I1235079,I1235096,I1235113,I1235144,I1235202,I1235228,I1235236,I1235262,I1235279,I1235301,I1235318,I1235335,I1235352,I1235369,I1235400,I1235417,I1235434,I1235451,I1235496,I1235513,I1235530,I1235589,I1235615,I1235623,I1235640,I1235657,I1235688,I1235746,I1235772,I1235780,I1235806,I1235823,I1235845,I1235862,I1235879,I1235896,I1235913,I1235944,I1235961,I1235978,I1235995,I1236040,I1236057,I1236074,I1236133,I1236159,I1236167,I1236184,I1236201,I1236232,I1236290,I1236316,I1236324,I1236350,I1236367,I1236389,I1236406,I1236423,I1236440,I1236457,I1236488,I1236505,I1236522,I1236539,I1236584,I1236601,I1236618,I1236677,I1236703,I1236711,I1236728,I1236745,I1236776,I1236834,I1236860,I1236868,I1236894,I1236911,I1236933,I1236950,I1236967,I1236984,I1237001,I1237032,I1237049,I1237066,I1237083,I1237128,I1237145,I1237162,I1237221,I1237247,I1237255,I1237272,I1237289,I1237320,I1237378,I1237404,I1237412,I1237438,I1237455,I1237477,I1237494,I1237511,I1237528,I1237545,I1237576,I1237593,I1237610,I1237627,I1237672,I1237689,I1237706,I1237765,I1237791,I1237799,I1237816,I1237833,I1237864,I1237922,I1237948,I1237956,I1237982,I1237999,I1238021,I1238038,I1238055,I1238072,I1238089,I1238120,I1238137,I1238154,I1238171,I1238216,I1238233,I1238250,I1238309,I1238335,I1238343,I1238360,I1238377,I1238408,I1238466,I1238492,I1238500,I1238526,I1238543,I1238565,I1238582,I1238599,I1238616,I1238633,I1238664,I1238681,I1238698,I1238715,I1238760,I1238777,I1238794,I1238853,I1238879,I1238887,I1238904,I1238921,I1238952,I1239010,I1239036,I1239044,I1239070,I1239087,I1239109,I1239126,I1239143,I1239160,I1239177,I1239208,I1239225,I1239242,I1239259,I1239304,I1239321,I1239338,I1239397,I1239423,I1239431,I1239448,I1239465,I1239496,I1239554,I1239580,I1239588,I1239614,I1239631,I1239546,I1239653,I1239670,I1239687,I1239704,I1239721,I1239525,I1239752,I1239769,I1239786,I1239803,I1239528,I1239543,I1239848,I1239865,I1239882,I1239540,I1239537,I1239534,I1239941,I1239967,I1239975,I1239992,I1240009,I1239522,I1240040,I1239531,I1240098,I1240124,I1240132,I1240158,I1240175,I1240197,I1240214,I1240231,I1240248,I1240265,I1240296,I1240313,I1240330,I1240347,I1240392,I1240409,I1240426,I1240485,I1240511,I1240519,I1240536,I1240553,I1240584,I1240642,I1240668,I1240676,I1240702,I1240719,I1240741,I1240758,I1240775,I1240792,I1240809,I1240840,I1240857,I1240874,I1240891,I1240936,I1240953,I1240970,I1241029,I1241055,I1241063,I1241080,I1241097,I1241128,I1241186,I1241212,I1241220,I1241246,I1241263,I1241285,I1241302,I1241319,I1241336,I1241353,I1241384,I1241401,I1241418,I1241435,I1241480,I1241497,I1241514,I1241573,I1241599,I1241607,I1241624,I1241641,I1241672,I1241730,I1241756,I1241764,I1241790,I1241807,I1241829,I1241846,I1241863,I1241880,I1241897,I1241928,I1241945,I1241962,I1241979,I1242024,I1242041,I1242058,I1242117,I1242143,I1242151,I1242168,I1242185,I1242216,I1242274,I1242300,I1242308,I1242334,I1242351,I1242373,I1242390,I1242407,I1242424,I1242441,I1242472,I1242489,I1242506,I1242523,I1242568,I1242585,I1242602,I1242661,I1242687,I1242695,I1242712,I1242729,I1242760,I1242818,I1242844,I1242852,I1242878,I1242895,I1242917,I1242934,I1242951,I1242968,I1242985,I1243016,I1243033,I1243050,I1243067,I1243112,I1243129,I1243146,I1243205,I1243231,I1243239,I1243256,I1243273,I1243304,I1243362,I1243388,I1243396,I1243422,I1243439,I1243461,I1243478,I1243495,I1243512,I1243529,I1243560,I1243577,I1243594,I1243611,I1243656,I1243673,I1243690,I1243749,I1243775,I1243783,I1243800,I1243817,I1243848,I1243906,I1243932,I1243940,I1243966,I1243983,I1244005,I1244022,I1244039,I1244056,I1244073,I1244104,I1244121,I1244138,I1244155,I1244200,I1244217,I1244234,I1244293,I1244319,I1244327,I1244344,I1244361,I1244392,I1244450,I1244476,I1244484,I1244510,I1244527,I1244549,I1244566,I1244583,I1244600,I1244617,I1244648,I1244665,I1244682,I1244699,I1244744,I1244761,I1244778,I1244837,I1244863,I1244871,I1244888,I1244905,I1244936,I1244994,I1245020,I1245028,I1245054,I1245071,I1245093,I1245110,I1245127,I1245144,I1245161,I1245192,I1245209,I1245226,I1245243,I1245288,I1245305,I1245322,I1245381,I1245407,I1245415,I1245432,I1245449,I1245480,I1245538,I1245564,I1245572,I1245598,I1245615,I1245637,I1245654,I1245671,I1245688,I1245705,I1245736,I1245753,I1245770,I1245787,I1245832,I1245849,I1245866,I1245925,I1245951,I1245959,I1245976,I1245993,I1246024,I1246082,I1246108,I1246116,I1246142,I1246159,I1246181,I1246198,I1246215,I1246232,I1246249,I1246280,I1246297,I1246314,I1246331,I1246376,I1246393,I1246410,I1246469,I1246495,I1246503,I1246520,I1246537,I1246568,I1246626,I1246652,I1246660,I1246686,I1246703,I1246725,I1246742,I1246759,I1246776,I1246793,I1246824,I1246841,I1246858,I1246875,I1246920,I1246937,I1246954,I1247013,I1247039,I1247047,I1247064,I1247081,I1247112,I1247170,I1247196,I1247204,I1247230,I1247247,I1247269,I1247286,I1247303,I1247320,I1247337,I1247368,I1247385,I1247402,I1247419,I1247464,I1247481,I1247498,I1247557,I1247583,I1247591,I1247608,I1247625,I1247656,I1247714,I1247740,I1247748,I1247774,I1247791,I1247813,I1247830,I1247847,I1247864,I1247881,I1247912,I1247929,I1247946,I1247963,I1248008,I1248025,I1248042,I1248101,I1248127,I1248135,I1248152,I1248169,I1248200,I1248258,I1248284,I1248292,I1248318,I1248335,I1248357,I1248374,I1248391,I1248408,I1248425,I1248456,I1248473,I1248490,I1248507,I1248552,I1248569,I1248586,I1248645,I1248671,I1248679,I1248696,I1248713,I1248744,I1248802,I1248828,I1248836,I1248862,I1248879,I1248901,I1248918,I1248935,I1248952,I1248969,I1249000,I1249017,I1249034,I1249051,I1249096,I1249113,I1249130,I1249189,I1249215,I1249223,I1249240,I1249257,I1249288,I1249346,I1249372,I1249380,I1249406,I1249423,I1249445,I1249462,I1249479,I1249496,I1249513,I1249544,I1249561,I1249578,I1249595,I1249640,I1249657,I1249674,I1249733,I1249759,I1249767,I1249784,I1249801,I1249832,I1249890,I1249916,I1249924,I1249950,I1249967,I1249989,I1250006,I1250023,I1250040,I1250057,I1250088,I1250105,I1250122,I1250139,I1250184,I1250201,I1250218,I1250277,I1250303,I1250311,I1250328,I1250345,I1250376,I1250434,I1250460,I1250468,I1250494,I1250511,I1250533,I1250550,I1250567,I1250584,I1250601,I1250632,I1250649,I1250666,I1250683,I1250728,I1250745,I1250762,I1250821,I1250847,I1250855,I1250872,I1250889,I1250920,I1250978,I1251004,I1251012,I1251038,I1251055,I1251077,I1251094,I1251111,I1251128,I1251145,I1251176,I1251193,I1251210,I1251227,I1251272,I1251289,I1251306,I1251365,I1251391,I1251399,I1251416,I1251433,I1251464,I1251522,I1251548,I1251556,I1251582,I1251599,I1251621,I1251638,I1251655,I1251672,I1251689,I1251720,I1251737,I1251754,I1251771,I1251816,I1251833,I1251850,I1251909,I1251935,I1251943,I1251960,I1251977,I1252008,I1252066,I1252092,I1252100,I1252126,I1252143,I1252165,I1252182,I1252199,I1252216,I1252233,I1252264,I1252281,I1252298,I1252315,I1252360,I1252377,I1252394,I1252453,I1252479,I1252487,I1252504,I1252521,I1252552,I1252610,I1252636,I1252644,I1252670,I1252687,I1252709,I1252726,I1252743,I1252760,I1252777,I1252808,I1252825,I1252842,I1252859,I1252904,I1252921,I1252938,I1252997,I1253023,I1253031,I1253048,I1253065,I1253096,I1253154,I1253180,I1253188,I1253214,I1253231,I1253253,I1253270,I1253287,I1253304,I1253321,I1253352,I1253369,I1253386,I1253403,I1253448,I1253465,I1253482,I1253541,I1253567,I1253575,I1253592,I1253609,I1253640,I1253698,I1253724,I1253732,I1253758,I1253775,I1253797,I1253814,I1253831,I1253848,I1253865,I1253896,I1253913,I1253930,I1253947,I1253992,I1254009,I1254026,I1254085,I1254111,I1254119,I1254136,I1254153,I1254184,I1254242,I1254268,I1254276,I1254302,I1254319,I1254341,I1254358,I1254375,I1254392,I1254409,I1254440,I1254457,I1254474,I1254491,I1254536,I1254553,I1254570,I1254629,I1254655,I1254663,I1254680,I1254697,I1254728,I1254786,I1254812,I1254820,I1254837,I1254863,I1254871,I1254888,I1254905,I1254922,I1254939,I1254970,I1254987,I1255004,I1255035,I1255052,I1255092,I1255100,I1255131,I1255148,I1255165,I1255182,I1255213,I1255244,I1255270,I1255292,I1255364,I1255390,I1255398,I1255415,I1255441,I1255449,I1255466,I1255483,I1255500,I1255517,I1255548,I1255565,I1255582,I1255613,I1255630,I1255670,I1255678,I1255709,I1255726,I1255743,I1255760,I1255791,I1255822,I1255848,I1255870,I1255942,I1255968,I1255976,I1255993,I1256019,I1256027,I1256044,I1256061,I1256078,I1256095,I1256126,I1256143,I1256160,I1256191,I1256208,I1256248,I1256256,I1256287,I1256304,I1256321,I1256338,I1256369,I1256400,I1256426,I1256448,I1256520,I1256546,I1256554,I1256571,I1256597,I1256605,I1256622,I1256639,I1256656,I1256673,I1256704,I1256721,I1256738,I1256769,I1256786,I1256826,I1256834,I1256865,I1256882,I1256899,I1256916,I1256947,I1256978,I1257004,I1257026,I1257098,I1257124,I1257132,I1257149,I1257175,I1257183,I1257200,I1257217,I1257234,I1257251,I1257282,I1257299,I1257316,I1257347,I1257364,I1257404,I1257412,I1257443,I1257460,I1257477,I1257494,I1257525,I1257556,I1257582,I1257604,I1257676,I1257702,I1257710,I1257727,I1257753,I1257761,I1257778,I1257795,I1257812,I1257829,I1257860,I1257877,I1257894,I1257925,I1257942,I1257982,I1257990,I1258021,I1258038,I1258055,I1258072,I1258103,I1258134,I1258160,I1258182,I1258254,I1258280,I1258288,I1258305,I1258331,I1258339,I1258356,I1258373,I1258390,I1258407,I1258438,I1258455,I1258472,I1258503,I1258520,I1258560,I1258568,I1258599,I1258616,I1258633,I1258650,I1258681,I1258712,I1258738,I1258760,I1258832,I1258858,I1258866,I1258883,I1258909,I1258917,I1258934,I1258951,I1258968,I1258985,I1259016,I1259033,I1259050,I1259081,I1259098,I1259138,I1259146,I1259177,I1259194,I1259211,I1259228,I1259259,I1259290,I1259316,I1259338,I1259410,I1259436,I1259444,I1259461,I1259487,I1259495,I1259512,I1259529,I1259546,I1259563,I1259594,I1259611,I1259628,I1259659,I1259676,I1259716,I1259724,I1259755,I1259772,I1259789,I1259806,I1259837,I1259868,I1259894,I1259916,I1259988,I1260014,I1260022,I1260039,I1260065,I1260073,I1260090,I1260107,I1260124,I1260141,I1260172,I1260189,I1260206,I1260237,I1260254,I1260294,I1260302,I1260333,I1260350,I1260367,I1260384,I1260415,I1260446,I1260472,I1260494,I1260566,I1297510,I1260592,I1260600,I1297504,I1260617,I1297519,I1260643,I1260651,I1260668,I1297495,I1260685,I1297492,I1260702,I1260719,I1297498,I1260750,I1260767,I1297507,I1260784,I1260815,I1297501,I1260832,I1260872,I1260880,I1260911,I1297516,I1260928,I1260945,I1260962,I1260993,I1261024,I1297513,I1261050,I1261072,I1261144,I1261170,I1261178,I1261195,I1261221,I1261229,I1261246,I1261263,I1261280,I1261297,I1261328,I1261345,I1261362,I1261393,I1261410,I1261450,I1261458,I1261489,I1261506,I1261523,I1261540,I1261571,I1261602,I1261628,I1261650,I1261722,I1261748,I1261756,I1261773,I1261799,I1261807,I1261824,I1261841,I1261858,I1261875,I1261906,I1261923,I1261940,I1261971,I1261988,I1262028,I1262036,I1262067,I1262084,I1262101,I1262118,I1262149,I1262180,I1262206,I1262228,I1262300,I1262326,I1262334,I1262351,I1262377,I1262385,I1262402,I1262419,I1262436,I1262453,I1262484,I1262501,I1262518,I1262549,I1262566,I1262606,I1262614,I1262645,I1262662,I1262679,I1262696,I1262727,I1262758,I1262784,I1262806,I1262878,I1262904,I1262912,I1262929,I1262955,I1262963,I1262980,I1262997,I1263014,I1263031,I1263062,I1263079,I1263096,I1263127,I1263144,I1263184,I1263192,I1263223,I1263240,I1263257,I1263274,I1263305,I1263336,I1263362,I1263384,I1263456,I1263482,I1263490,I1263507,I1263533,I1263541,I1263558,I1263575,I1263592,I1263609,I1263640,I1263657,I1263674,I1263705,I1263722,I1263762,I1263770,I1263801,I1263818,I1263835,I1263852,I1263883,I1263914,I1263940,I1263962,I1264034,I1264060,I1264068,I1264085,I1264111,I1264119,I1264136,I1264153,I1264170,I1264187,I1264218,I1264235,I1264252,I1264283,I1264300,I1264340,I1264348,I1264379,I1264396,I1264413,I1264430,I1264461,I1264492,I1264518,I1264540,I1264612,I1264638,I1264646,I1264663,I1264689,I1264697,I1264714,I1264731,I1264748,I1264765,I1264796,I1264813,I1264830,I1264861,I1264878,I1264918,I1264926,I1264957,I1264974,I1264991,I1265008,I1265039,I1265070,I1265096,I1265118,I1265190,I1265216,I1265224,I1265241,I1265267,I1265275,I1265292,I1265309,I1265326,I1265343,I1265374,I1265391,I1265408,I1265439,I1265456,I1265496,I1265504,I1265535,I1265552,I1265569,I1265586,I1265617,I1265648,I1265674,I1265696,I1265768,I1265794,I1265802,I1265819,I1265845,I1265853,I1265870,I1265887,I1265904,I1265921,I1265952,I1265969,I1265986,I1266017,I1266034,I1266074,I1266082,I1266113,I1266130,I1266147,I1266164,I1266195,I1266226,I1266252,I1266274,I1266346,I1266372,I1266380,I1266397,I1266423,I1266431,I1266448,I1266465,I1266482,I1266499,I1266530,I1266547,I1266564,I1266595,I1266612,I1266652,I1266660,I1266691,I1266708,I1266725,I1266742,I1266773,I1266804,I1266830,I1266852,I1266924,I1266950,I1266958,I1266975,I1267001,I1267009,I1267026,I1267043,I1267060,I1267077,I1267108,I1267125,I1267142,I1267173,I1267190,I1267230,I1267238,I1267269,I1267286,I1267303,I1267320,I1267351,I1267382,I1267408,I1267430,I1267502,I1267528,I1267536,I1267553,I1267579,I1267587,I1267604,I1267621,I1267638,I1267655,I1267686,I1267703,I1267720,I1267751,I1267768,I1267808,I1267816,I1267847,I1267864,I1267881,I1267898,I1267929,I1267960,I1267986,I1268008,I1268080,I1268106,I1268114,I1268131,I1268157,I1268165,I1268182,I1268199,I1268216,I1268233,I1268264,I1268281,I1268298,I1268329,I1268346,I1268386,I1268394,I1268425,I1268442,I1268459,I1268476,I1268507,I1268538,I1268564,I1268586,I1268658,I1268684,I1268692,I1268709,I1268735,I1268743,I1268760,I1268777,I1268794,I1268811,I1268842,I1268859,I1268876,I1268907,I1268924,I1268964,I1268972,I1269003,I1269020,I1269037,I1269054,I1269085,I1269116,I1269142,I1269164,I1269236,I1269262,I1269270,I1269287,I1269313,I1269321,I1269338,I1269355,I1269372,I1269389,I1269420,I1269437,I1269454,I1269485,I1269502,I1269542,I1269550,I1269581,I1269598,I1269615,I1269632,I1269663,I1269694,I1269720,I1269742,I1269814,I1269840,I1269848,I1269865,I1269891,I1269899,I1269916,I1269933,I1269950,I1269967,I1269998,I1270015,I1270032,I1270063,I1270080,I1270120,I1270128,I1270159,I1270176,I1270193,I1270210,I1270241,I1270272,I1270298,I1270320,I1270392,I1270418,I1270426,I1270443,I1270469,I1270477,I1270494,I1270511,I1270528,I1270545,I1270576,I1270593,I1270610,I1270641,I1270658,I1270698,I1270706,I1270737,I1270754,I1270771,I1270788,I1270819,I1270850,I1270876,I1270898,I1270970,I1270996,I1271004,I1271021,I1271047,I1271055,I1271072,I1271089,I1271106,I1271123,I1270962,I1271154,I1271171,I1271188,I1270941,I1271219,I1271236,I1270947,I1271276,I1271284,I1270956,I1271315,I1271332,I1271349,I1271366,I1270959,I1271397,I1270938,I1271428,I1271454,I1270953,I1271476,I1270950,I1270944,I1271548,I1271574,I1271582,I1271599,I1271625,I1271633,I1271650,I1271667,I1271684,I1271701,I1271732,I1271749,I1271766,I1271797,I1271814,I1271854,I1271862,I1271893,I1271910,I1271927,I1271944,I1271975,I1272006,I1272032,I1272054,I1272126,I1317831,I1272152,I1272160,I1317822,I1272177,I1317807,I1272203,I1272211,I1272228,I1317810,I1272245,I1317819,I1272262,I1272279,I1317816,I1272310,I1317828,I1272327,I1272344,I1272375,I1317813,I1272392,I1272432,I1272440,I1272471,I1317834,I1272488,I1272505,I1272522,I1272553,I1272584,I1317825,I1272610,I1272632,I1272704,I1272730,I1272738,I1272755,I1272781,I1272789,I1272806,I1272823,I1272840,I1272857,I1272888,I1272905,I1272922,I1272953,I1272970,I1273010,I1273018,I1273049,I1273066,I1273083,I1273100,I1273131,I1273162,I1273188,I1273210,I1273282,I1273308,I1273316,I1273333,I1273359,I1273367,I1273384,I1273401,I1273418,I1273435,I1273274,I1273466,I1273483,I1273500,I1273253,I1273531,I1273548,I1273259,I1273588,I1273596,I1273268,I1273627,I1273644,I1273661,I1273678,I1273271,I1273709,I1273250,I1273740,I1273766,I1273265,I1273788,I1273262,I1273256,I1273860,I1273886,I1273894,I1273911,I1273937,I1273945,I1273962,I1273979,I1273996,I1274013,I1274044,I1274061,I1274078,I1274109,I1274126,I1274166,I1274174,I1274205,I1274222,I1274239,I1274256,I1274287,I1274318,I1274344,I1274366,I1274438,I1274464,I1274472,I1274489,I1274515,I1274523,I1274540,I1274557,I1274574,I1274591,I1274622,I1274639,I1274656,I1274687,I1274704,I1274744,I1274752,I1274783,I1274800,I1274817,I1274834,I1274865,I1274896,I1274922,I1274944,I1275016,I1275042,I1275050,I1275067,I1275093,I1275101,I1275118,I1275135,I1275152,I1275169,I1275200,I1275217,I1275234,I1275265,I1275282,I1275322,I1275330,I1275361,I1275378,I1275395,I1275412,I1275443,I1275474,I1275500,I1275522,I1275594,I1275620,I1275628,I1275645,I1275671,I1275679,I1275696,I1275713,I1275730,I1275747,I1275778,I1275795,I1275812,I1275843,I1275860,I1275900,I1275908,I1275939,I1275956,I1275973,I1275990,I1276021,I1276052,I1276078,I1276100,I1276172,I1276198,I1276206,I1276223,I1276249,I1276257,I1276274,I1276291,I1276308,I1276325,I1276356,I1276373,I1276390,I1276421,I1276438,I1276478,I1276486,I1276517,I1276534,I1276551,I1276568,I1276599,I1276630,I1276656,I1276678,I1276750,I1276776,I1276784,I1276801,I1276827,I1276835,I1276852,I1276869,I1276886,I1276903,I1276934,I1276951,I1276968,I1276999,I1277016,I1277056,I1277064,I1277095,I1277112,I1277129,I1277146,I1277177,I1277208,I1277234,I1277256,I1277328,I1277354,I1277362,I1277379,I1277405,I1277413,I1277430,I1277447,I1277464,I1277481,I1277512,I1277529,I1277546,I1277577,I1277594,I1277634,I1277642,I1277673,I1277690,I1277707,I1277724,I1277755,I1277786,I1277812,I1277834,I1277906,I1277932,I1277940,I1277957,I1277983,I1277991,I1278008,I1278025,I1278042,I1278059,I1278090,I1278107,I1278124,I1278155,I1278172,I1278212,I1278220,I1278251,I1278268,I1278285,I1278302,I1278333,I1278364,I1278390,I1278412,I1278484,I1278510,I1278518,I1278535,I1278561,I1278569,I1278586,I1278603,I1278620,I1278637,I1278668,I1278685,I1278702,I1278733,I1278750,I1278790,I1278798,I1278829,I1278846,I1278863,I1278880,I1278911,I1278942,I1278968,I1278990,I1279062,I1279088,I1279096,I1279113,I1279139,I1279147,I1279164,I1279181,I1279198,I1279215,I1279246,I1279263,I1279280,I1279311,I1279328,I1279368,I1279376,I1279407,I1279424,I1279441,I1279458,I1279489,I1279520,I1279546,I1279568,I1279640,I1279666,I1279674,I1279691,I1279717,I1279725,I1279742,I1279759,I1279776,I1279793,I1279824,I1279841,I1279858,I1279889,I1279906,I1279946,I1279954,I1279985,I1280002,I1280019,I1280036,I1280067,I1280098,I1280124,I1280146,I1280218,I1328541,I1280244,I1280252,I1328532,I1280269,I1328517,I1280295,I1280303,I1280320,I1328520,I1280337,I1328529,I1280354,I1280371,I1328526,I1280402,I1328538,I1280419,I1280436,I1280467,I1328523,I1280484,I1280524,I1280532,I1280563,I1328544,I1280580,I1280597,I1280614,I1280645,I1280676,I1328535,I1280702,I1280724,I1280796,I1280822,I1280830,I1280847,I1280873,I1280881,I1280898,I1280915,I1280932,I1280949,I1280980,I1280997,I1281014,I1281045,I1281062,I1281102,I1281110,I1281141,I1281158,I1281175,I1281192,I1281223,I1281254,I1281280,I1281302,I1281374,I1281400,I1281408,I1281425,I1281451,I1281459,I1281476,I1281493,I1281510,I1281527,I1281558,I1281575,I1281592,I1281623,I1281640,I1281680,I1281688,I1281719,I1281736,I1281753,I1281770,I1281801,I1281832,I1281858,I1281880,I1281952,I1281978,I1281986,I1282003,I1282029,I1282037,I1282054,I1282071,I1282088,I1282105,I1282136,I1282153,I1282170,I1282201,I1282218,I1282258,I1282266,I1282297,I1282314,I1282331,I1282348,I1282379,I1282410,I1282436,I1282458,I1282530,I1282556,I1282564,I1282581,I1282607,I1282615,I1282632,I1282649,I1282666,I1282683,I1282714,I1282731,I1282748,I1282779,I1282796,I1282836,I1282844,I1282875,I1282892,I1282909,I1282926,I1282957,I1282988,I1283014,I1283036,I1283108,I1283134,I1283142,I1283159,I1283185,I1283193,I1283210,I1283227,I1283244,I1283261,I1283292,I1283309,I1283326,I1283357,I1283374,I1283414,I1283422,I1283453,I1283470,I1283487,I1283504,I1283535,I1283566,I1283592,I1283614,I1283686,I1283712,I1283720,I1283737,I1283763,I1283771,I1283788,I1283805,I1283822,I1283839,I1283870,I1283887,I1283904,I1283935,I1283952,I1283992,I1284000,I1284031,I1284048,I1284065,I1284082,I1284113,I1284144,I1284170,I1284192,I1284264,I1374356,I1284290,I1284298,I1374347,I1284315,I1374332,I1284341,I1284349,I1284366,I1374335,I1284383,I1374344,I1284400,I1284417,I1374341,I1284448,I1374353,I1284465,I1284482,I1284513,I1374338,I1284530,I1284570,I1284578,I1284609,I1374359,I1284626,I1284643,I1284660,I1284691,I1284722,I1374350,I1284748,I1284770,I1284842,I1284868,I1284876,I1284893,I1284919,I1284927,I1284944,I1284961,I1284978,I1284995,I1285026,I1285043,I1285060,I1285091,I1285108,I1285148,I1285156,I1285187,I1285204,I1285221,I1285238,I1285269,I1285300,I1285326,I1285348,I1285420,I1285446,I1285454,I1285471,I1285497,I1285505,I1285522,I1285539,I1285556,I1285573,I1285604,I1285621,I1285638,I1285669,I1285686,I1285726,I1285734,I1285765,I1285782,I1285799,I1285816,I1285847,I1285878,I1285904,I1285926,I1285998,I1286024,I1286032,I1286049,I1286075,I1286083,I1286100,I1286117,I1286134,I1286151,I1286182,I1286199,I1286216,I1286247,I1286264,I1286304,I1286312,I1286343,I1286360,I1286377,I1286394,I1286425,I1286456,I1286482,I1286504,I1286576,I1286602,I1286610,I1286627,I1286653,I1286661,I1286678,I1286695,I1286712,I1286729,I1286760,I1286777,I1286794,I1286825,I1286842,I1286882,I1286890,I1286921,I1286938,I1286955,I1286972,I1287003,I1287034,I1287060,I1287082,I1287154,I1287180,I1287188,I1287205,I1287231,I1287239,I1287256,I1287273,I1287290,I1287307,I1287338,I1287355,I1287372,I1287403,I1287420,I1287460,I1287468,I1287499,I1287516,I1287533,I1287550,I1287581,I1287612,I1287638,I1287660,I1287732,I1287758,I1287766,I1287783,I1287809,I1287817,I1287834,I1287851,I1287868,I1287885,I1287916,I1287933,I1287950,I1287981,I1287998,I1288038,I1288046,I1288077,I1288094,I1288111,I1288128,I1288159,I1288190,I1288216,I1288238,I1288310,I1288336,I1288344,I1288361,I1288387,I1288395,I1288412,I1288429,I1288446,I1288463,I1288494,I1288511,I1288528,I1288559,I1288576,I1288616,I1288624,I1288655,I1288672,I1288689,I1288706,I1288737,I1288768,I1288794,I1288816,I1288888,I1288914,I1288922,I1288939,I1288965,I1288973,I1288990,I1289007,I1289024,I1289041,I1289072,I1289089,I1289106,I1289137,I1289154,I1289194,I1289202,I1289233,I1289250,I1289267,I1289284,I1289315,I1289346,I1289372,I1289394,I1289466,I1289492,I1289500,I1289517,I1289543,I1289551,I1289568,I1289585,I1289602,I1289619,I1289650,I1289667,I1289684,I1289715,I1289732,I1289772,I1289780,I1289811,I1289828,I1289845,I1289862,I1289893,I1289924,I1289950,I1289972,I1290044,I1290070,I1290078,I1290095,I1290121,I1290129,I1290146,I1290163,I1290180,I1290197,I1290228,I1290245,I1290262,I1290293,I1290310,I1290350,I1290358,I1290389,I1290406,I1290423,I1290440,I1290471,I1290502,I1290528,I1290550,I1290622,I1298071,I1290648,I1290656,I1298065,I1290673,I1298080,I1290699,I1290707,I1290724,I1298056,I1290741,I1298053,I1290758,I1290775,I1298059,I1290806,I1290823,I1298068,I1290840,I1290871,I1298062,I1290888,I1290928,I1290936,I1290967,I1298077,I1290984,I1291001,I1291018,I1291049,I1291080,I1298074,I1291106,I1291128,I1291200,I1291226,I1291234,I1291251,I1291277,I1291285,I1291302,I1291319,I1291336,I1291353,I1291384,I1291401,I1291418,I1291449,I1291466,I1291506,I1291514,I1291545,I1291562,I1291579,I1291596,I1291627,I1291658,I1291684,I1291706,I1291778,I1291804,I1291812,I1291829,I1291855,I1291863,I1291880,I1291897,I1291914,I1291931,I1291962,I1291979,I1291996,I1292027,I1292044,I1292084,I1292092,I1292123,I1292140,I1292157,I1292174,I1292205,I1292236,I1292262,I1292284,I1292356,I1292382,I1292390,I1292407,I1292433,I1292441,I1292458,I1292475,I1292492,I1292509,I1292540,I1292557,I1292574,I1292605,I1292622,I1292662,I1292670,I1292701,I1292718,I1292735,I1292752,I1292783,I1292814,I1292840,I1292862,I1292934,I1333896,I1292960,I1292968,I1333887,I1292985,I1333872,I1293011,I1293019,I1293036,I1333875,I1293053,I1333884,I1293070,I1293087,I1333881,I1293118,I1333893,I1293135,I1293152,I1293183,I1333878,I1293200,I1293240,I1293248,I1293279,I1333899,I1293296,I1293313,I1293330,I1293361,I1293392,I1333890,I1293418,I1293440,I1293512,I1293538,I1293546,I1293563,I1293589,I1293597,I1293614,I1293631,I1293648,I1293665,I1293504,I1293696,I1293713,I1293730,I1293483,I1293761,I1293778,I1293489,I1293818,I1293826,I1293498,I1293857,I1293874,I1293891,I1293908,I1293501,I1293939,I1293480,I1293970,I1293996,I1293495,I1294018,I1293492,I1293486,I1294090,I1294116,I1294124,I1294141,I1294167,I1294175,I1294192,I1294209,I1294226,I1294243,I1294274,I1294291,I1294308,I1294339,I1294356,I1294396,I1294404,I1294435,I1294452,I1294469,I1294486,I1294517,I1294548,I1294574,I1294596,I1294668,I1294694,I1294702,I1294719,I1294745,I1294753,I1294770,I1294787,I1294804,I1294821,I1294852,I1294869,I1294886,I1294917,I1294934,I1294974,I1294982,I1295013,I1295030,I1295047,I1295064,I1295095,I1295126,I1295152,I1295174,I1295246,I1326756,I1295272,I1295280,I1326747,I1295297,I1326732,I1295323,I1295331,I1295348,I1326735,I1295365,I1326744,I1295382,I1295399,I1326741,I1295430,I1326753,I1295447,I1295464,I1295495,I1326738,I1295512,I1295552,I1295560,I1295591,I1326759,I1295608,I1295625,I1295642,I1295673,I1295704,I1326750,I1295730,I1295752,I1295824,I1295850,I1295858,I1295875,I1295901,I1295909,I1295926,I1295943,I1295960,I1295977,I1296008,I1296025,I1296042,I1296073,I1296090,I1296130,I1296138,I1296169,I1296186,I1296203,I1296220,I1296251,I1296282,I1296308,I1296330,I1296405,I1296431,I1296439,I1296456,I1296482,I1296490,I1296507,I1296524,I1296555,I1296586,I1296603,I1296620,I1296637,I1296654,I1296685,I1296744,I1296761,I1296787,I1296809,I1296835,I1296843,I1296860,I1296891,I1296966,I1296992,I1297000,I1297017,I1297043,I1297051,I1297068,I1297085,I1297116,I1297147,I1297164,I1297181,I1297198,I1297215,I1297246,I1297305,I1297322,I1297348,I1297370,I1297396,I1297404,I1297421,I1297452,I1297527,I1297553,I1297561,I1297578,I1297604,I1297612,I1297629,I1297646,I1297677,I1297708,I1297725,I1297742,I1297759,I1297776,I1297807,I1297866,I1297883,I1297909,I1297931,I1297957,I1297965,I1297982,I1298013,I1298088,I1298114,I1298122,I1298139,I1298165,I1298173,I1298190,I1298207,I1298238,I1298269,I1298286,I1298303,I1298320,I1298337,I1298368,I1298427,I1298444,I1298470,I1298492,I1298518,I1298526,I1298543,I1298574,I1298649,I1298675,I1298683,I1298700,I1298726,I1298734,I1298751,I1298768,I1298799,I1298830,I1298847,I1298864,I1298881,I1298898,I1298929,I1298988,I1299005,I1299031,I1299053,I1299079,I1299087,I1299104,I1299135,I1299210,I1325557,I1299236,I1299244,I1325551,I1299261,I1325569,I1299287,I1299295,I1299312,I1325554,I1325545,I1299329,I1299360,I1325560,I1299391,I1325563,I1299408,I1325566,I1299425,I1299442,I1325548,I1299459,I1299490,I1299549,I1325542,I1299566,I1299592,I1299614,I1299640,I1299648,I1299665,I1299696,I1299771,I1299797,I1299805,I1299822,I1299848,I1299856,I1299873,I1299890,I1299921,I1299952,I1299969,I1299986,I1300003,I1300020,I1300051,I1300110,I1300127,I1300153,I1300175,I1300201,I1300209,I1300226,I1300257,I1300332,I1300358,I1300366,I1300383,I1300409,I1300417,I1300434,I1300451,I1300482,I1300513,I1300530,I1300547,I1300564,I1300581,I1300612,I1300671,I1300688,I1300714,I1300736,I1300762,I1300770,I1300787,I1300818,I1300893,I1341622,I1300919,I1300927,I1341616,I1300944,I1341634,I1300970,I1300978,I1300995,I1341619,I1341610,I1301012,I1301043,I1341625,I1301074,I1341628,I1301091,I1341631,I1301108,I1301125,I1341613,I1301142,I1301173,I1301232,I1341607,I1301249,I1301275,I1301297,I1301323,I1301331,I1301348,I1301379,I1301454,I1301480,I1301488,I1301505,I1301531,I1301539,I1301556,I1301573,I1301604,I1301635,I1301652,I1301669,I1301686,I1301703,I1301734,I1301793,I1301810,I1301836,I1301858,I1301884,I1301892,I1301909,I1301940,I1302015,I1302041,I1302049,I1302066,I1302092,I1302100,I1302117,I1302134,I1302165,I1302196,I1302213,I1302230,I1302247,I1302264,I1302295,I1302354,I1302371,I1302397,I1302419,I1302445,I1302453,I1302470,I1302501,I1302576,I1302602,I1302610,I1302627,I1302653,I1302661,I1302678,I1302695,I1302726,I1302757,I1302774,I1302791,I1302808,I1302825,I1302856,I1302915,I1302932,I1302958,I1302980,I1303006,I1303014,I1303031,I1303062,I1303137,I1303163,I1303171,I1303188,I1303214,I1303222,I1303239,I1303256,I1303287,I1303318,I1303335,I1303352,I1303369,I1303386,I1303417,I1303476,I1303493,I1303519,I1303541,I1303567,I1303575,I1303592,I1303623,I1303698,I1339837,I1303724,I1303732,I1339831,I1303749,I1339849,I1303775,I1303783,I1303800,I1339834,I1339825,I1303817,I1303848,I1339840,I1303879,I1339843,I1303896,I1339846,I1303913,I1303930,I1339828,I1303947,I1303978,I1304037,I1339822,I1304054,I1304080,I1304102,I1304128,I1304136,I1304153,I1304184,I1304259,I1304285,I1304293,I1304310,I1304336,I1304344,I1304361,I1304378,I1304409,I1304440,I1304457,I1304474,I1304491,I1304508,I1304539,I1304598,I1304615,I1304641,I1304663,I1304689,I1304697,I1304714,I1304745,I1304820,I1304846,I1304854,I1304871,I1304897,I1304905,I1304922,I1304939,I1304970,I1305001,I1305018,I1305035,I1305052,I1305069,I1305100,I1305159,I1305176,I1305202,I1305224,I1305250,I1305258,I1305275,I1305306,I1305381,I1305407,I1305415,I1305432,I1305458,I1305466,I1305483,I1305500,I1305531,I1305562,I1305579,I1305596,I1305613,I1305630,I1305661,I1305720,I1305737,I1305763,I1305785,I1305811,I1305819,I1305836,I1305867,I1305942,I1305968,I1305985,I1305993,I1306038,I1306055,I1306072,I1306089,I1306106,I1306123,I1306140,I1306171,I1306188,I1306233,I1306250,I1306267,I1306298,I1306324,I1306332,I1306363,I1306380,I1306397,I1306423,I1306431,I1306448,I1306537,I1306563,I1306580,I1306588,I1306633,I1306650,I1306667,I1306684,I1306701,I1306718,I1306735,I1306766,I1306783,I1306828,I1306845,I1306862,I1306893,I1306919,I1306927,I1306958,I1306975,I1306992,I1307018,I1307026,I1307043,I1307132,I1307158,I1307175,I1307183,I1307228,I1307245,I1307262,I1307279,I1307296,I1307313,I1307330,I1307361,I1307378,I1307423,I1307440,I1307457,I1307488,I1307514,I1307522,I1307553,I1307570,I1307587,I1307613,I1307621,I1307638,I1307727,I1307753,I1307770,I1307778,I1307823,I1307840,I1307857,I1307874,I1307891,I1307908,I1307925,I1307956,I1307973,I1308018,I1308035,I1308052,I1308083,I1308109,I1308117,I1308148,I1308165,I1308182,I1308208,I1308216,I1308233,I1308322,I1308348,I1308365,I1308373,I1308418,I1308435,I1308452,I1308469,I1308486,I1308503,I1308520,I1308551,I1308568,I1308613,I1308630,I1308647,I1308678,I1308704,I1308712,I1308743,I1308760,I1308777,I1308803,I1308811,I1308828,I1308917,I1308943,I1308960,I1308968,I1309013,I1309030,I1309047,I1309064,I1309081,I1309098,I1309115,I1309146,I1309163,I1309208,I1309225,I1309242,I1309273,I1309299,I1309307,I1309338,I1309355,I1309372,I1309398,I1309406,I1309423,I1309512,I1309538,I1309555,I1309563,I1309608,I1309625,I1309642,I1309659,I1309676,I1309693,I1309710,I1309741,I1309758,I1309803,I1309820,I1309837,I1309868,I1309894,I1309902,I1309933,I1309950,I1309967,I1309993,I1310001,I1310018,I1310107,I1310133,I1310150,I1310158,I1310203,I1310220,I1310237,I1310254,I1310271,I1310288,I1310305,I1310336,I1310353,I1310398,I1310415,I1310432,I1310463,I1310489,I1310497,I1310528,I1310545,I1310562,I1310588,I1310596,I1310613,I1310702,I1310728,I1310745,I1310753,I1310798,I1310815,I1310832,I1310849,I1310866,I1310883,I1310900,I1310931,I1310948,I1310993,I1311010,I1311027,I1311058,I1311084,I1311092,I1311123,I1311140,I1311157,I1311183,I1311191,I1311208,I1311297,I1311323,I1311340,I1311348,I1311393,I1311410,I1311427,I1311444,I1311461,I1311478,I1311495,I1311526,I1311543,I1311588,I1311605,I1311622,I1311653,I1311679,I1311687,I1311718,I1311735,I1311752,I1311778,I1311786,I1311803,I1311892,I1311918,I1311935,I1311943,I1311988,I1312005,I1312022,I1312039,I1312056,I1312073,I1312090,I1312121,I1312138,I1312183,I1312200,I1312217,I1312248,I1312274,I1312282,I1312313,I1312330,I1312347,I1312373,I1312381,I1312398,I1312487,I1312513,I1312530,I1312538,I1312583,I1312600,I1312617,I1312634,I1312651,I1312668,I1312685,I1312716,I1312733,I1312778,I1312795,I1312812,I1312843,I1312869,I1312877,I1312908,I1312925,I1312942,I1312968,I1312976,I1312993,I1313082,I1313108,I1313125,I1313133,I1313178,I1313195,I1313212,I1313229,I1313246,I1313263,I1313280,I1313311,I1313328,I1313373,I1313390,I1313407,I1313438,I1313464,I1313472,I1313503,I1313520,I1313537,I1313563,I1313571,I1313588,I1313677,I1313703,I1313720,I1313728,I1313773,I1313790,I1313807,I1313824,I1313841,I1313858,I1313875,I1313906,I1313923,I1313968,I1313985,I1314002,I1314033,I1314059,I1314067,I1314098,I1314115,I1314132,I1314158,I1314166,I1314183,I1314272,I1314298,I1314315,I1314323,I1314368,I1314385,I1314402,I1314419,I1314436,I1314453,I1314470,I1314501,I1314518,I1314563,I1314580,I1314597,I1314628,I1314654,I1314662,I1314693,I1314710,I1314727,I1314753,I1314761,I1314778,I1314867,I1314893,I1314910,I1314918,I1314963,I1314980,I1314997,I1315014,I1315031,I1315048,I1315065,I1315096,I1315113,I1315158,I1315175,I1315192,I1315223,I1315249,I1315257,I1315288,I1315305,I1315322,I1315348,I1315356,I1315373,I1315462,I1315488,I1315505,I1315513,I1315558,I1315575,I1315592,I1315609,I1315626,I1315643,I1315660,I1315691,I1315708,I1315753,I1315770,I1315787,I1315818,I1315844,I1315852,I1315883,I1315900,I1315917,I1315943,I1315951,I1315968,I1316057,I1316083,I1316100,I1316108,I1316153,I1316170,I1316187,I1316204,I1316221,I1316238,I1316255,I1316286,I1316303,I1316348,I1316365,I1316382,I1316413,I1316439,I1316447,I1316478,I1316495,I1316512,I1316538,I1316546,I1316563,I1316652,I1316678,I1316695,I1316703,I1316748,I1316765,I1316782,I1316799,I1316816,I1316833,I1316850,I1316881,I1316898,I1316943,I1316960,I1316977,I1317008,I1317034,I1317042,I1317073,I1317090,I1317107,I1317133,I1317141,I1317158,I1317247,I1317273,I1317290,I1317298,I1317343,I1317360,I1317377,I1317394,I1317411,I1317428,I1317445,I1317476,I1317493,I1317538,I1317555,I1317572,I1317603,I1317629,I1317637,I1317668,I1317685,I1317702,I1317728,I1317736,I1317753,I1317842,I1317868,I1317885,I1317893,I1317938,I1317955,I1317972,I1317989,I1318006,I1318023,I1318040,I1318071,I1318088,I1318133,I1318150,I1318167,I1318198,I1318224,I1318232,I1318263,I1318280,I1318297,I1318323,I1318331,I1318348,I1318437,I1318463,I1318480,I1318488,I1318533,I1318550,I1318567,I1318584,I1318601,I1318618,I1318635,I1318666,I1318683,I1318728,I1318745,I1318762,I1318793,I1318819,I1318827,I1318858,I1318875,I1318892,I1318918,I1318926,I1318943,I1319032,I1319058,I1319075,I1319083,I1319128,I1319145,I1319162,I1319179,I1319196,I1319213,I1319230,I1319261,I1319278,I1319323,I1319340,I1319357,I1319388,I1319414,I1319422,I1319453,I1319470,I1319487,I1319513,I1319521,I1319538,I1319627,I1319653,I1319670,I1319678,I1319723,I1319740,I1319757,I1319774,I1319791,I1319808,I1319825,I1319856,I1319873,I1319918,I1319935,I1319952,I1319983,I1320009,I1320017,I1320048,I1320065,I1320082,I1320108,I1320116,I1320133,I1320222,I1320248,I1320265,I1320273,I1320318,I1320335,I1320352,I1320369,I1320386,I1320403,I1320420,I1320451,I1320468,I1320513,I1320530,I1320547,I1320578,I1320604,I1320612,I1320643,I1320660,I1320677,I1320703,I1320711,I1320728,I1320817,I1320843,I1320860,I1320868,I1320913,I1320930,I1320947,I1320964,I1320981,I1320998,I1321015,I1321046,I1321063,I1321108,I1321125,I1321142,I1321173,I1321199,I1321207,I1321238,I1321255,I1321272,I1321298,I1321306,I1321323,I1321412,I1321438,I1321455,I1321463,I1321508,I1321525,I1321542,I1321559,I1321576,I1321593,I1321610,I1321641,I1321658,I1321703,I1321720,I1321737,I1321768,I1321794,I1321802,I1321833,I1321850,I1321867,I1321893,I1321901,I1321918,I1322007,I1322033,I1322050,I1322058,I1322103,I1322120,I1322137,I1322154,I1322171,I1322188,I1322205,I1322236,I1322253,I1322298,I1322315,I1322332,I1322363,I1322389,I1322397,I1322428,I1322445,I1322462,I1322488,I1322496,I1322513,I1322602,I1322628,I1322645,I1322653,I1322698,I1322715,I1322732,I1322749,I1322766,I1322783,I1322800,I1322831,I1322848,I1322893,I1322910,I1322927,I1322958,I1322984,I1322992,I1323023,I1323040,I1323057,I1323083,I1323091,I1323108,I1323197,I1323223,I1323240,I1323248,I1323293,I1323310,I1323327,I1323344,I1323361,I1323378,I1323395,I1323426,I1323443,I1323488,I1323505,I1323522,I1323553,I1323579,I1323587,I1323618,I1323635,I1323652,I1323678,I1323686,I1323703,I1323792,I1323818,I1323835,I1323843,I1323888,I1323905,I1323922,I1323939,I1323956,I1323973,I1323990,I1324021,I1324038,I1324083,I1324100,I1324117,I1324148,I1324174,I1324182,I1324213,I1324230,I1324247,I1324273,I1324281,I1324298,I1324387,I1324413,I1324430,I1324438,I1324483,I1324500,I1324517,I1324534,I1324551,I1324568,I1324585,I1324616,I1324633,I1324678,I1324695,I1324712,I1324743,I1324769,I1324777,I1324808,I1324825,I1324842,I1324868,I1324876,I1324893,I1324982,I1325008,I1325025,I1325033,I1325078,I1325095,I1325112,I1325129,I1325146,I1325163,I1325180,I1325211,I1325228,I1325273,I1325290,I1325307,I1325338,I1325364,I1325372,I1325403,I1325420,I1325437,I1325463,I1325471,I1325488,I1325577,I1325603,I1325620,I1325628,I1325673,I1325690,I1325707,I1325724,I1325741,I1325758,I1325775,I1325806,I1325823,I1325868,I1325885,I1325902,I1325933,I1325959,I1325967,I1325998,I1326015,I1326032,I1326058,I1326066,I1326083,I1326172,I1326198,I1326215,I1326223,I1326268,I1326285,I1326302,I1326319,I1326336,I1326353,I1326370,I1326401,I1326418,I1326463,I1326480,I1326497,I1326528,I1326554,I1326562,I1326593,I1326610,I1326627,I1326653,I1326661,I1326678,I1326767,I1326793,I1326810,I1326818,I1326863,I1326880,I1326897,I1326914,I1326931,I1326948,I1326965,I1326996,I1327013,I1327058,I1327075,I1327092,I1327123,I1327149,I1327157,I1327188,I1327205,I1327222,I1327248,I1327256,I1327273,I1327362,I1327388,I1327405,I1327413,I1327458,I1327475,I1327492,I1327509,I1327526,I1327543,I1327560,I1327591,I1327608,I1327653,I1327670,I1327687,I1327718,I1327744,I1327752,I1327783,I1327800,I1327817,I1327843,I1327851,I1327868,I1327957,I1327983,I1328000,I1328008,I1328053,I1328070,I1328087,I1328104,I1328121,I1328138,I1328155,I1328186,I1328203,I1328248,I1328265,I1328282,I1328313,I1328339,I1328347,I1328378,I1328395,I1328412,I1328438,I1328446,I1328463,I1328552,I1328578,I1328595,I1328603,I1328648,I1328665,I1328682,I1328699,I1328716,I1328733,I1328750,I1328781,I1328798,I1328843,I1328860,I1328877,I1328908,I1328934,I1328942,I1328973,I1328990,I1329007,I1329033,I1329041,I1329058,I1329147,I1329173,I1329190,I1329198,I1329243,I1329260,I1329277,I1329294,I1329311,I1329328,I1329345,I1329376,I1329393,I1329438,I1329455,I1329472,I1329503,I1329529,I1329537,I1329568,I1329585,I1329602,I1329628,I1329636,I1329653,I1329742,I1329768,I1329785,I1329793,I1329838,I1329855,I1329872,I1329889,I1329906,I1329923,I1329940,I1329971,I1329988,I1330033,I1330050,I1330067,I1330098,I1330124,I1330132,I1330163,I1330180,I1330197,I1330223,I1330231,I1330248,I1330337,I1330363,I1330380,I1330388,I1330433,I1330450,I1330467,I1330484,I1330501,I1330518,I1330535,I1330566,I1330583,I1330628,I1330645,I1330662,I1330693,I1330719,I1330727,I1330758,I1330775,I1330792,I1330818,I1330826,I1330843,I1330932,I1330958,I1330975,I1330983,I1331028,I1331045,I1331062,I1331079,I1331096,I1331113,I1331130,I1331161,I1331178,I1331223,I1331240,I1331257,I1331288,I1331314,I1331322,I1331353,I1331370,I1331387,I1331413,I1331421,I1331438,I1331527,I1331553,I1331570,I1331578,I1331623,I1331640,I1331657,I1331674,I1331691,I1331708,I1331725,I1331756,I1331773,I1331818,I1331835,I1331852,I1331883,I1331909,I1331917,I1331948,I1331965,I1331982,I1332008,I1332016,I1332033,I1332122,I1332148,I1332165,I1332173,I1332218,I1332235,I1332252,I1332269,I1332286,I1332303,I1332320,I1332351,I1332368,I1332413,I1332430,I1332447,I1332478,I1332504,I1332512,I1332543,I1332560,I1332577,I1332603,I1332611,I1332628,I1332717,I1332743,I1332760,I1332768,I1332813,I1332830,I1332847,I1332864,I1332881,I1332898,I1332915,I1332946,I1332963,I1333008,I1333025,I1333042,I1333073,I1333099,I1333107,I1333138,I1333155,I1333172,I1333198,I1333206,I1333223,I1333312,I1333338,I1333355,I1333363,I1333408,I1333425,I1333442,I1333459,I1333476,I1333493,I1333510,I1333541,I1333558,I1333603,I1333620,I1333637,I1333668,I1333694,I1333702,I1333733,I1333750,I1333767,I1333793,I1333801,I1333818,I1333907,I1333933,I1333950,I1333958,I1334003,I1334020,I1334037,I1334054,I1334071,I1334088,I1334105,I1334136,I1334153,I1334198,I1334215,I1334232,I1334263,I1334289,I1334297,I1334328,I1334345,I1334362,I1334388,I1334396,I1334413,I1334502,I1334528,I1334545,I1334553,I1334598,I1334615,I1334632,I1334649,I1334666,I1334683,I1334700,I1334731,I1334748,I1334793,I1334810,I1334827,I1334858,I1334884,I1334892,I1334923,I1334940,I1334957,I1334983,I1334991,I1335008,I1335097,I1335123,I1335140,I1335148,I1335193,I1335210,I1335227,I1335244,I1335261,I1335278,I1335295,I1335326,I1335343,I1335388,I1335405,I1335422,I1335453,I1335479,I1335487,I1335518,I1335535,I1335552,I1335578,I1335586,I1335603,I1335692,I1335718,I1335735,I1335743,I1335788,I1335805,I1335822,I1335839,I1335856,I1335873,I1335890,I1335921,I1335938,I1335983,I1336000,I1336017,I1336048,I1336074,I1336082,I1336113,I1336130,I1336147,I1336173,I1336181,I1336198,I1336287,I1336313,I1336330,I1336338,I1336383,I1336400,I1336417,I1336434,I1336451,I1336468,I1336485,I1336516,I1336533,I1336578,I1336595,I1336612,I1336643,I1336669,I1336677,I1336708,I1336725,I1336742,I1336768,I1336776,I1336793,I1336882,I1336908,I1336925,I1336933,I1336978,I1336995,I1337012,I1337029,I1337046,I1337063,I1337080,I1337111,I1337128,I1337173,I1337190,I1337207,I1337238,I1337264,I1337272,I1337303,I1337320,I1337337,I1337363,I1337371,I1337388,I1337477,I1337503,I1337520,I1337528,I1337573,I1337590,I1337607,I1337624,I1337641,I1337658,I1337675,I1337706,I1337723,I1337768,I1337785,I1337802,I1337833,I1337859,I1337867,I1337898,I1337915,I1337932,I1337958,I1337966,I1337983,I1338072,I1338098,I1338115,I1338123,I1338168,I1338185,I1338202,I1338219,I1338236,I1338253,I1338270,I1338301,I1338318,I1338363,I1338380,I1338397,I1338428,I1338454,I1338462,I1338493,I1338510,I1338527,I1338553,I1338561,I1338578,I1338667,I1338693,I1338710,I1338718,I1338763,I1338780,I1338797,I1338814,I1338831,I1338848,I1338865,I1338896,I1338913,I1338958,I1338975,I1338992,I1339023,I1339049,I1339057,I1339088,I1339105,I1339122,I1339148,I1339156,I1339173,I1339262,I1339288,I1339305,I1339313,I1339358,I1339375,I1339392,I1339409,I1339426,I1339443,I1339460,I1339491,I1339508,I1339553,I1339570,I1339587,I1339618,I1339644,I1339652,I1339683,I1339700,I1339717,I1339743,I1339751,I1339768,I1339857,I1339883,I1339900,I1339908,I1339953,I1339970,I1339987,I1340004,I1340021,I1340038,I1340055,I1340086,I1340103,I1340148,I1340165,I1340182,I1340213,I1340239,I1340247,I1340278,I1340295,I1340312,I1340338,I1340346,I1340363,I1340452,I1340478,I1340495,I1340503,I1340548,I1340565,I1340582,I1340599,I1340616,I1340633,I1340650,I1340681,I1340698,I1340743,I1340760,I1340777,I1340808,I1340834,I1340842,I1340873,I1340890,I1340907,I1340933,I1340941,I1340958,I1341047,I1341073,I1341090,I1341098,I1341143,I1341160,I1341177,I1341194,I1341211,I1341228,I1341245,I1341276,I1341293,I1341338,I1341355,I1341372,I1341403,I1341429,I1341437,I1341468,I1341485,I1341502,I1341528,I1341536,I1341553,I1341642,I1341668,I1341685,I1341693,I1341738,I1341755,I1341772,I1341789,I1341806,I1341823,I1341840,I1341871,I1341888,I1341933,I1341950,I1341967,I1341998,I1342024,I1342032,I1342063,I1342080,I1342097,I1342123,I1342131,I1342148,I1342237,I1342263,I1342280,I1342288,I1342333,I1342350,I1342367,I1342384,I1342401,I1342418,I1342435,I1342466,I1342483,I1342528,I1342545,I1342562,I1342593,I1342619,I1342627,I1342658,I1342675,I1342692,I1342718,I1342726,I1342743,I1342832,I1342858,I1342875,I1342883,I1342928,I1342945,I1342962,I1342979,I1342996,I1343013,I1343030,I1343061,I1343078,I1343123,I1343140,I1343157,I1343188,I1343214,I1343222,I1343253,I1343270,I1343287,I1343313,I1343321,I1343338,I1343427,I1343453,I1343470,I1343478,I1343523,I1343540,I1343557,I1343574,I1343591,I1343608,I1343625,I1343656,I1343673,I1343718,I1343735,I1343752,I1343783,I1343809,I1343817,I1343848,I1343865,I1343882,I1343908,I1343916,I1343933,I1344022,I1344048,I1344065,I1344073,I1344118,I1344135,I1344152,I1344169,I1344186,I1344203,I1344220,I1344251,I1344268,I1344313,I1344330,I1344347,I1344378,I1344404,I1344412,I1344443,I1344460,I1344477,I1344503,I1344511,I1344528,I1344617,I1344643,I1344660,I1344668,I1344713,I1344730,I1344747,I1344764,I1344781,I1344798,I1344815,I1344846,I1344863,I1344908,I1344925,I1344942,I1344973,I1344999,I1345007,I1345038,I1345055,I1345072,I1345098,I1345106,I1345123,I1345212,I1345238,I1345255,I1345263,I1345308,I1345325,I1345342,I1345359,I1345376,I1345393,I1345410,I1345441,I1345458,I1345503,I1345520,I1345537,I1345568,I1345594,I1345602,I1345633,I1345650,I1345667,I1345693,I1345701,I1345718,I1345807,I1345833,I1345850,I1345858,I1345903,I1345920,I1345937,I1345954,I1345971,I1345988,I1346005,I1346036,I1346053,I1346098,I1346115,I1346132,I1346163,I1346189,I1346197,I1346228,I1346245,I1346262,I1346288,I1346296,I1346313,I1346402,I1346428,I1346445,I1346453,I1346498,I1346515,I1346532,I1346549,I1346566,I1346583,I1346600,I1346631,I1346648,I1346693,I1346710,I1346727,I1346758,I1346784,I1346792,I1346823,I1346840,I1346857,I1346883,I1346891,I1346908,I1346997,I1347023,I1347040,I1347048,I1347093,I1347110,I1347127,I1347144,I1347161,I1347178,I1347195,I1347226,I1347243,I1347288,I1347305,I1347322,I1347353,I1347379,I1347387,I1347418,I1347435,I1347452,I1347478,I1347486,I1347503,I1347592,I1347618,I1347635,I1347643,I1347688,I1347705,I1347722,I1347739,I1347756,I1347773,I1347790,I1347821,I1347838,I1347883,I1347900,I1347917,I1347948,I1347974,I1347982,I1348013,I1348030,I1348047,I1348073,I1348081,I1348098,I1348187,I1348213,I1348230,I1348238,I1348283,I1348300,I1348317,I1348334,I1348351,I1348368,I1348385,I1348416,I1348433,I1348478,I1348495,I1348512,I1348543,I1348569,I1348577,I1348608,I1348625,I1348642,I1348668,I1348676,I1348693,I1348782,I1348808,I1348825,I1348833,I1348878,I1348895,I1348912,I1348929,I1348946,I1348963,I1348980,I1349011,I1349028,I1349073,I1349090,I1349107,I1349138,I1349164,I1349172,I1349203,I1349220,I1349237,I1349263,I1349271,I1349288,I1349377,I1349403,I1349420,I1349428,I1349473,I1349490,I1349507,I1349524,I1349541,I1349558,I1349575,I1349606,I1349623,I1349668,I1349685,I1349702,I1349733,I1349759,I1349767,I1349798,I1349815,I1349832,I1349858,I1349866,I1349883,I1349972,I1349998,I1350015,I1350023,I1350068,I1350085,I1350102,I1350119,I1350136,I1350153,I1350170,I1350201,I1350218,I1350263,I1350280,I1350297,I1350328,I1350354,I1350362,I1350393,I1350410,I1350427,I1350453,I1350461,I1350478,I1350567,I1350593,I1350610,I1350618,I1350663,I1350680,I1350697,I1350714,I1350731,I1350748,I1350765,I1350796,I1350813,I1350858,I1350875,I1350892,I1350923,I1350949,I1350957,I1350988,I1351005,I1351022,I1351048,I1351056,I1351073,I1351162,I1351188,I1351205,I1351213,I1351258,I1351275,I1351292,I1351309,I1351326,I1351343,I1351360,I1351391,I1351408,I1351453,I1351470,I1351487,I1351518,I1351544,I1351552,I1351583,I1351600,I1351617,I1351643,I1351651,I1351668,I1351757,I1351783,I1351800,I1351808,I1351853,I1351870,I1351887,I1351904,I1351921,I1351938,I1351955,I1351986,I1352003,I1352048,I1352065,I1352082,I1352113,I1352139,I1352147,I1352178,I1352195,I1352212,I1352238,I1352246,I1352263,I1352352,I1352378,I1352395,I1352403,I1352448,I1352465,I1352482,I1352499,I1352516,I1352533,I1352550,I1352581,I1352598,I1352643,I1352660,I1352677,I1352708,I1352734,I1352742,I1352773,I1352790,I1352807,I1352833,I1352841,I1352858,I1352947,I1352973,I1352990,I1352998,I1353043,I1353060,I1353077,I1353094,I1353111,I1353128,I1353145,I1353176,I1353193,I1353238,I1353255,I1353272,I1353303,I1353329,I1353337,I1353368,I1353385,I1353402,I1353428,I1353436,I1353453,I1353542,I1353568,I1353585,I1353593,I1353638,I1353655,I1353672,I1353689,I1353706,I1353723,I1353740,I1353771,I1353788,I1353833,I1353850,I1353867,I1353898,I1353924,I1353932,I1353963,I1353980,I1353997,I1354023,I1354031,I1354048,I1354137,I1354163,I1354180,I1354188,I1354233,I1354250,I1354267,I1354284,I1354301,I1354318,I1354335,I1354366,I1354383,I1354428,I1354445,I1354462,I1354493,I1354519,I1354527,I1354558,I1354575,I1354592,I1354618,I1354626,I1354643,I1354732,I1354758,I1354775,I1354783,I1354828,I1354845,I1354862,I1354879,I1354896,I1354913,I1354930,I1354961,I1354978,I1355023,I1355040,I1355057,I1355088,I1355114,I1355122,I1355153,I1355170,I1355187,I1355213,I1355221,I1355238,I1355327,I1355353,I1355370,I1355378,I1355423,I1355440,I1355457,I1355474,I1355491,I1355508,I1355525,I1355556,I1355573,I1355618,I1355635,I1355652,I1355683,I1355709,I1355717,I1355748,I1355765,I1355782,I1355808,I1355816,I1355833,I1355922,I1355948,I1355965,I1355973,I1356018,I1356035,I1356052,I1356069,I1356086,I1356103,I1356120,I1356151,I1356168,I1356213,I1356230,I1356247,I1356278,I1356304,I1356312,I1356343,I1356360,I1356377,I1356403,I1356411,I1356428,I1356517,I1356543,I1356560,I1356568,I1356613,I1356630,I1356647,I1356664,I1356681,I1356698,I1356715,I1356746,I1356763,I1356808,I1356825,I1356842,I1356873,I1356899,I1356907,I1356938,I1356955,I1356972,I1356998,I1357006,I1357023,I1357112,I1357138,I1357155,I1357163,I1357208,I1357225,I1357242,I1357259,I1357276,I1357293,I1357310,I1357341,I1357358,I1357403,I1357420,I1357437,I1357468,I1357494,I1357502,I1357533,I1357550,I1357567,I1357593,I1357601,I1357618,I1357707,I1357733,I1357750,I1357758,I1357803,I1357820,I1357837,I1357854,I1357871,I1357888,I1357905,I1357936,I1357953,I1357998,I1358015,I1358032,I1358063,I1358089,I1358097,I1358128,I1358145,I1358162,I1358188,I1358196,I1358213,I1358302,I1358328,I1358345,I1358353,I1358398,I1358415,I1358432,I1358449,I1358466,I1358483,I1358500,I1358531,I1358548,I1358593,I1358610,I1358627,I1358658,I1358684,I1358692,I1358723,I1358740,I1358757,I1358783,I1358791,I1358808,I1358897,I1358923,I1358940,I1358948,I1358993,I1359010,I1359027,I1359044,I1359061,I1359078,I1359095,I1359126,I1359143,I1359188,I1359205,I1359222,I1359253,I1359279,I1359287,I1359318,I1359335,I1359352,I1359378,I1359386,I1359403,I1359492,I1359518,I1359535,I1359543,I1359588,I1359605,I1359622,I1359639,I1359656,I1359673,I1359690,I1359721,I1359738,I1359783,I1359800,I1359817,I1359848,I1359874,I1359882,I1359913,I1359930,I1359947,I1359973,I1359981,I1359998,I1360087,I1360113,I1360130,I1360138,I1360183,I1360200,I1360217,I1360234,I1360251,I1360268,I1360285,I1360316,I1360333,I1360378,I1360395,I1360412,I1360443,I1360469,I1360477,I1360508,I1360525,I1360542,I1360568,I1360576,I1360593,I1360682,I1360708,I1360725,I1360733,I1360778,I1360795,I1360812,I1360829,I1360846,I1360863,I1360880,I1360911,I1360928,I1360973,I1360990,I1361007,I1361038,I1361064,I1361072,I1361103,I1361120,I1361137,I1361163,I1361171,I1361188,I1361277,I1361303,I1361320,I1361328,I1361373,I1361390,I1361407,I1361424,I1361441,I1361458,I1361475,I1361506,I1361523,I1361568,I1361585,I1361602,I1361633,I1361659,I1361667,I1361698,I1361715,I1361732,I1361758,I1361766,I1361783,I1361872,I1361898,I1361915,I1361923,I1361968,I1361985,I1362002,I1362019,I1362036,I1362053,I1362070,I1362101,I1362118,I1362163,I1362180,I1362197,I1362228,I1362254,I1362262,I1362293,I1362310,I1362327,I1362353,I1362361,I1362378,I1362467,I1362493,I1362510,I1362518,I1362563,I1362580,I1362597,I1362614,I1362631,I1362648,I1362665,I1362696,I1362713,I1362758,I1362775,I1362792,I1362823,I1362849,I1362857,I1362888,I1362905,I1362922,I1362948,I1362956,I1362973,I1363062,I1363088,I1363105,I1363113,I1363158,I1363175,I1363192,I1363209,I1363226,I1363243,I1363260,I1363291,I1363308,I1363353,I1363370,I1363387,I1363418,I1363444,I1363452,I1363483,I1363500,I1363517,I1363543,I1363551,I1363568,I1363657,I1363683,I1363700,I1363708,I1363753,I1363770,I1363787,I1363804,I1363821,I1363838,I1363855,I1363886,I1363903,I1363948,I1363965,I1363982,I1364013,I1364039,I1364047,I1364078,I1364095,I1364112,I1364138,I1364146,I1364163,I1364252,I1364278,I1364295,I1364303,I1364348,I1364365,I1364382,I1364399,I1364416,I1364433,I1364450,I1364481,I1364498,I1364543,I1364560,I1364577,I1364608,I1364634,I1364642,I1364673,I1364690,I1364707,I1364733,I1364741,I1364758,I1364847,I1364873,I1364890,I1364898,I1364943,I1364960,I1364977,I1364994,I1365011,I1365028,I1365045,I1365076,I1365093,I1365138,I1365155,I1365172,I1365203,I1365229,I1365237,I1365268,I1365285,I1365302,I1365328,I1365336,I1365353,I1365442,I1365468,I1365485,I1365493,I1365538,I1365555,I1365572,I1365589,I1365606,I1365623,I1365640,I1365671,I1365688,I1365733,I1365750,I1365767,I1365798,I1365824,I1365832,I1365863,I1365880,I1365897,I1365923,I1365931,I1365948,I1366037,I1366063,I1366080,I1366088,I1366133,I1366150,I1366167,I1366184,I1366201,I1366218,I1366235,I1366266,I1366283,I1366328,I1366345,I1366362,I1366393,I1366419,I1366427,I1366458,I1366475,I1366492,I1366518,I1366526,I1366543,I1366632,I1366658,I1366675,I1366683,I1366728,I1366745,I1366762,I1366779,I1366796,I1366813,I1366830,I1366861,I1366878,I1366923,I1366940,I1366957,I1366988,I1367014,I1367022,I1367053,I1367070,I1367087,I1367113,I1367121,I1367138,I1367227,I1367253,I1367270,I1367278,I1367323,I1367340,I1367357,I1367374,I1367391,I1367408,I1367425,I1367456,I1367473,I1367518,I1367535,I1367552,I1367583,I1367609,I1367617,I1367648,I1367665,I1367682,I1367708,I1367716,I1367733,I1367822,I1367848,I1367865,I1367873,I1367918,I1367935,I1367952,I1367969,I1367986,I1368003,I1368020,I1368051,I1368068,I1368113,I1368130,I1368147,I1368178,I1368204,I1368212,I1368243,I1368260,I1368277,I1368303,I1368311,I1368328,I1368417,I1368443,I1368460,I1368468,I1368513,I1368530,I1368547,I1368564,I1368581,I1368598,I1368615,I1368646,I1368663,I1368708,I1368725,I1368742,I1368773,I1368799,I1368807,I1368838,I1368855,I1368872,I1368898,I1368906,I1368923,I1369012,I1369038,I1369055,I1369063,I1369108,I1369125,I1369142,I1369159,I1369176,I1369193,I1369210,I1369241,I1369258,I1369303,I1369320,I1369337,I1369368,I1369394,I1369402,I1369433,I1369450,I1369467,I1369493,I1369501,I1369518,I1369607,I1369633,I1369650,I1369658,I1369703,I1369720,I1369737,I1369754,I1369771,I1369788,I1369805,I1369836,I1369853,I1369898,I1369915,I1369932,I1369963,I1369989,I1369997,I1370028,I1370045,I1370062,I1370088,I1370096,I1370113,I1370202,I1370228,I1370245,I1370253,I1370298,I1370315,I1370332,I1370349,I1370366,I1370383,I1370400,I1370431,I1370448,I1370493,I1370510,I1370527,I1370558,I1370584,I1370592,I1370623,I1370640,I1370657,I1370683,I1370691,I1370708,I1370797,I1370823,I1370840,I1370848,I1370893,I1370910,I1370927,I1370944,I1370961,I1370978,I1370995,I1371026,I1371043,I1371088,I1371105,I1371122,I1371153,I1371179,I1371187,I1371218,I1371235,I1371252,I1371278,I1371286,I1371303,I1371392,I1371418,I1371435,I1371443,I1371488,I1371505,I1371522,I1371539,I1371556,I1371573,I1371590,I1371621,I1371638,I1371683,I1371700,I1371717,I1371748,I1371774,I1371782,I1371813,I1371830,I1371847,I1371873,I1371881,I1371898,I1371987,I1372013,I1372030,I1372038,I1372083,I1372100,I1372117,I1372134,I1372151,I1372168,I1372185,I1372216,I1372233,I1372278,I1372295,I1372312,I1372343,I1372369,I1372377,I1372408,I1372425,I1372442,I1372468,I1372476,I1372493,I1372582,I1372608,I1372625,I1372633,I1372678,I1372695,I1372712,I1372729,I1372746,I1372763,I1372780,I1372811,I1372828,I1372873,I1372890,I1372907,I1372938,I1372964,I1372972,I1373003,I1373020,I1373037,I1373063,I1373071,I1373088,I1373177,I1373203,I1373220,I1373228,I1373273,I1373290,I1373307,I1373324,I1373341,I1373358,I1373375,I1373406,I1373423,I1373468,I1373485,I1373502,I1373533,I1373559,I1373567,I1373598,I1373615,I1373632,I1373658,I1373666,I1373683,I1373772,I1373798,I1373815,I1373823,I1373868,I1373885,I1373902,I1373919,I1373936,I1373953,I1373970,I1374001,I1374018,I1374063,I1374080,I1374097,I1374128,I1374154,I1374162,I1374193,I1374210,I1374227,I1374253,I1374261,I1374278,I1374367,I1374393,I1374410,I1374418,I1374463,I1374480,I1374497,I1374514,I1374531,I1374548,I1374565,I1374596,I1374613,I1374658,I1374675,I1374692,I1374723,I1374749,I1374757,I1374788,I1374805,I1374822,I1374848,I1374856,I1374873,I1374962,I1374988,I1375005,I1375013,I1375058,I1375075,I1375092,I1375109,I1375126,I1375143,I1375160,I1375191,I1375208,I1375253,I1375270,I1375287,I1375318,I1375344,I1375352,I1375383,I1375400,I1375417,I1375443,I1375451,I1375468,I1375557,I1375583,I1375600,I1375608,I1375653,I1375670,I1375687,I1375704,I1375721,I1375738,I1375755,I1375786,I1375803,I1375848,I1375865,I1375882,I1375913,I1375939,I1375947,I1375978,I1375995,I1376012,I1376038,I1376046,I1376063,I1376152,I1376178,I1376195,I1376203,I1376248,I1376265,I1376282,I1376299,I1376316,I1376333,I1376350,I1376381,I1376398,I1376443,I1376460,I1376477,I1376508,I1376534,I1376542,I1376573,I1376590,I1376607,I1376633,I1376641,I1376658,I1376747,I1376773,I1376790,I1376798,I1376843,I1376860,I1376877,I1376894,I1376911,I1376928,I1376945,I1376976,I1376993,I1377038,I1377055,I1377072,I1377103,I1377129,I1377137,I1377168,I1377185,I1377202,I1377228,I1377236,I1377253,I1377342,I1377368,I1377385,I1377393,I1377438,I1377455,I1377472,I1377489,I1377506,I1377523,I1377540,I1377571,I1377588,I1377633,I1377650,I1377667,I1377698,I1377724,I1377732,I1377763,I1377780,I1377797,I1377823,I1377831,I1377848,I1377937,I1377963,I1377980,I1377988,I1378033,I1378050,I1378067,I1378084,I1378101,I1378118,I1378135,I1378166,I1378183,I1378228,I1378245,I1378262,I1378293,I1378319,I1378327,I1378358,I1378375,I1378392,I1378418,I1378426,I1378443,I1378532,I1378558,I1378575,I1378583,I1378628,I1378645,I1378662,I1378679,I1378696,I1378713,I1378730,I1378761,I1378778,I1378823,I1378840,I1378857,I1378888,I1378914,I1378922,I1378953,I1378970,I1378987,I1379013,I1379021,I1379038,I1379127,I1379153,I1379170,I1379178,I1379223,I1379240,I1379257,I1379274,I1379291,I1379308,I1379325,I1379356,I1379373,I1379418,I1379435,I1379452,I1379483,I1379509,I1379517,I1379548,I1379565,I1379582,I1379608,I1379616,I1379633,I1379722,I1379748,I1379765,I1379773,I1379818,I1379835,I1379852,I1379869,I1379886,I1379903,I1379920,I1379951,I1379968,I1380013,I1380030,I1380047,I1380078,I1380104,I1380112,I1380143,I1380160,I1380177,I1380203,I1380211,I1380228,I1380317,I1380343,I1380360,I1380368,I1380413,I1380430,I1380447,I1380464,I1380481,I1380498,I1380515,I1380546,I1380563,I1380608,I1380625,I1380642,I1380673,I1380699,I1380707,I1380738,I1380755,I1380772,I1380798,I1380806,I1380823,I1380912,I1380938,I1380955,I1380963,I1381008,I1381025,I1381042,I1381059,I1381076,I1381093,I1381110,I1381141,I1381158,I1381203,I1381220,I1381237,I1381268,I1381294,I1381302,I1381333,I1381350,I1381367,I1381393,I1381401,I1381418,I1381507,I1381533,I1381550,I1381558,I1381603,I1381620,I1381637,I1381654,I1381671,I1381688,I1381705,I1381736,I1381753,I1381798,I1381815,I1381832,I1381863,I1381889,I1381897,I1381928,I1381945,I1381962,I1381988,I1381996,I1382013,I1382102,I1382128,I1382145,I1382153,I1382198,I1382215,I1382232,I1382249,I1382266,I1382283,I1382300,I1382331,I1382348,I1382393,I1382410,I1382427,I1382458,I1382484,I1382492,I1382523,I1382540,I1382557,I1382583,I1382591,I1382608,I1382697,I1382723,I1382740,I1382748,I1382793,I1382810,I1382827,I1382844,I1382861,I1382878,I1382895,I1382926,I1382943,I1382988,I1383005,I1383022,I1383053,I1383079,I1383087,I1383118,I1383135,I1383152,I1383178,I1383186,I1383203,I1383292,I1383318,I1383335,I1383343,I1383388,I1383405,I1383422,I1383439,I1383456,I1383473,I1383490,I1383521,I1383538,I1383583,I1383600,I1383617,I1383648,I1383674,I1383682,I1383713,I1383730,I1383747,I1383773,I1383781,I1383798,I1383887,I1383913,I1383930,I1383938,I1383983,I1384000,I1384017,I1384034,I1384051,I1384068,I1384085,I1384116,I1384133,I1384178,I1384195,I1384212,I1384243,I1384269,I1384277,I1384308,I1384325,I1384342,I1384368,I1384376,I1384393,I1384482,I1384508,I1384525,I1384533,I1384578,I1384595,I1384612,I1384629,I1384646,I1384663,I1384680,I1384711,I1384728,I1384773,I1384790,I1384807,I1384838,I1384864,I1384872,I1384903,I1384920,I1384937,I1384963,I1384971,I1384988,I1385077,I1385103,I1385120,I1385128,I1385173,I1385190,I1385207,I1385224,I1385241,I1385258,I1385275,I1385306,I1385323,I1385368,I1385385,I1385402,I1385433,I1385459,I1385467,I1385498,I1385515,I1385532,I1385558,I1385566,I1385583,I1385672,I1385698,I1385715,I1385723,I1385768,I1385785,I1385802,I1385819,I1385836,I1385853,I1385870,I1385901,I1385918,I1385963,I1385980,I1385997,I1386028,I1386054,I1386062,I1386093,I1386110,I1386127,I1386153,I1386161,I1386178,I1386267,I1386293,I1386310,I1386318,I1386363,I1386380,I1386397,I1386414,I1386431,I1386448,I1386465,I1386496,I1386513,I1386558,I1386575,I1386592,I1386623,I1386649,I1386657,I1386688,I1386705,I1386722,I1386748,I1386756,I1386773,I1386862,I1386888,I1386905,I1386913,I1386958,I1386975,I1386992,I1387009,I1387026,I1387043,I1387060,I1387091,I1387108,I1387153,I1387170,I1387187,I1387218,I1387244,I1387252,I1387283,I1387300,I1387317,I1387343,I1387351,I1387368,I1387457,I1387483,I1387500,I1387508,I1387553,I1387570,I1387587,I1387604,I1387621,I1387638,I1387655,I1387686,I1387703,I1387748,I1387765,I1387782,I1387813,I1387839,I1387847,I1387878,I1387895,I1387912,I1387938,I1387946,I1387963,I1388052,I1388078,I1388095,I1388103,I1388148,I1388165,I1388182,I1388199,I1388216,I1388233,I1388250,I1388281,I1388298,I1388343,I1388360,I1388377,I1388408,I1388434,I1388442,I1388473,I1388490,I1388507,I1388533,I1388541,I1388558,I1388647,I1388673,I1388690,I1388698,I1388743,I1388760,I1388777,I1388794,I1388811,I1388828,I1388845,I1388876,I1388893,I1388938,I1388955,I1388972,I1389003,I1389029,I1389037,I1389068,I1389085,I1389102,I1389128,I1389136,I1389153,I1389242,I1389268,I1389285,I1389293,I1389338,I1389355,I1389372,I1389389,I1389406,I1389423,I1389440,I1389471,I1389488,I1389533,I1389550,I1389567,I1389598,I1389624,I1389632,I1389663,I1389680,I1389697,I1389723,I1389731,I1389748,I1389837,I1389863,I1389880,I1389888,I1389933,I1389950,I1389967,I1389984,I1390001,I1390018,I1390035,I1390066,I1390083,I1390128,I1390145,I1390162,I1390193,I1390219,I1390227,I1390258,I1390275,I1390292,I1390318,I1390326,I1390343,I1390432,I1390458,I1390475,I1390483,I1390528,I1390545,I1390562,I1390579,I1390596,I1390613,I1390630,I1390661,I1390678,I1390723,I1390740,I1390757,I1390788,I1390814,I1390822,I1390853,I1390870,I1390887,I1390913,I1390921,I1390938,I1391027,I1391053,I1391070,I1391078,I1391123,I1391140,I1391157,I1391174,I1391191,I1391208,I1391225,I1391256,I1391273,I1391318,I1391335,I1391352,I1391383,I1391409,I1391417,I1391448,I1391465,I1391482,I1391508,I1391516,I1391533,I1391622,I1391648,I1391665,I1391673,I1391718,I1391735,I1391752,I1391769,I1391786,I1391803,I1391820,I1391851,I1391868,I1391913,I1391930,I1391947,I1391978,I1392004,I1392012,I1392043,I1392060,I1392077,I1392103,I1392111,I1392128,I1392217,I1392243,I1392260,I1392268,I1392313,I1392330,I1392347,I1392364,I1392381,I1392398,I1392415,I1392446,I1392463,I1392508,I1392525,I1392542,I1392573,I1392599,I1392607,I1392638,I1392655,I1392672,I1392698,I1392706,I1392723,I1392812,I1392838,I1392855,I1392863,I1392908,I1392925,I1392942,I1392959,I1392976,I1392993,I1393010,I1393041,I1393058,I1393103,I1393120,I1393137,I1393168,I1393194,I1393202,I1393233,I1393250,I1393267,I1393293,I1393301,I1393318,I1393407,I1393433,I1393450,I1393458,I1393503,I1393520,I1393537,I1393554,I1393571,I1393588,I1393605,I1393636,I1393653,I1393698,I1393715,I1393732,I1393763,I1393789,I1393797,I1393828,I1393845,I1393862,I1393888,I1393896,I1393913,I1394002,I1394028,I1394045,I1394053,I1394098,I1394115,I1394132,I1394149,I1394166,I1394183,I1394200,I1394231,I1394248,I1394293,I1394310,I1394327,I1394358,I1394384,I1394392,I1394423,I1394440,I1394457,I1394483,I1394491,I1394508,I1394597,I1394623,I1394640,I1394648,I1394693,I1394710,I1394727,I1394744,I1394761,I1394778,I1394795,I1394826,I1394843,I1394888,I1394905,I1394922,I1394953,I1394979,I1394987,I1395018,I1395035,I1395052,I1395078,I1395086,I1395103,I1395192,I1395218,I1395235,I1395243,I1395288,I1395305,I1395322,I1395339,I1395356,I1395373,I1395390,I1395421,I1395438,I1395483,I1395500,I1395517,I1395548,I1395574,I1395582,I1395613,I1395630,I1395647,I1395673,I1395681,I1395698,I1395787,I1395813,I1395830,I1395838,I1395883,I1395900,I1395917,I1395934,I1395951,I1395968,I1395985,I1396016,I1396033,I1396078,I1396095,I1396112,I1396143,I1396169,I1396177,I1396208,I1396225,I1396242,I1396268,I1396276,I1396293;
not I_0 (I2546,I2514);
DFFARX1 I_1 (I208543,I2507,I2546,I2572,);
nand I_2 (I2580,I2572,I208543);
not I_3 (I2597,I2580);
DFFARX1 I_4 (I2597,I2507,I2546,I2538,);
DFFARX1 I_5 (I208549,I2507,I2546,I2637,);
not I_6 (I2645,I2637);
not I_7 (I2662,I208558);
not I_8 (I2679,I208552);
nand I_9 (I2696,I2645,I2679);
nor I_10 (I2713,I2696,I208558);
DFFARX1 I_11 (I2713,I2507,I2546,I2517,);
nor I_12 (I2744,I208552,I208558);
nand I_13 (I2761,I2637,I2744);
nor I_14 (I2778,I208555,I208561);
nor I_15 (I2520,I2696,I208555);
not I_16 (I2809,I208555);
not I_17 (I2826,I208564);
nand I_18 (I2843,I2826,I208540);
nand I_19 (I2860,I2662,I2843);
not I_20 (I2877,I2860);
nor I_21 (I2894,I208564,I208561);
nor I_22 (I2529,I2877,I2894);
nor I_23 (I2925,I208546,I208564);
and I_24 (I2942,I2925,I2778);
nor I_25 (I2959,I2860,I2942);
DFFARX1 I_26 (I2959,I2507,I2546,I2535,);
nor I_27 (I2990,I2580,I2942);
DFFARX1 I_28 (I2990,I2507,I2546,I2532,);
nor I_29 (I3021,I208546,I208540);
DFFARX1 I_30 (I3021,I2507,I2546,I3047,);
nor I_31 (I3055,I3047,I208552);
nand I_32 (I3072,I3055,I2662);
nand I_33 (I2526,I3072,I2761);
nand I_34 (I2523,I3055,I2809);
not I_35 (I3141,I2514);
DFFARX1 I_36 (I775242,I2507,I3141,I3167,);
nand I_37 (I3175,I3167,I775221);
not I_38 (I3192,I3175);
DFFARX1 I_39 (I3192,I2507,I3141,I3133,);
DFFARX1 I_40 (I775230,I2507,I3141,I3232,);
not I_41 (I3240,I3232);
not I_42 (I3257,I775236);
not I_43 (I3274,I775233);
nand I_44 (I3291,I3240,I3274);
nor I_45 (I3308,I3291,I775236);
DFFARX1 I_46 (I3308,I2507,I3141,I3112,);
nor I_47 (I3339,I775233,I775236);
nand I_48 (I3356,I3232,I3339);
nor I_49 (I3373,I775224,I775218);
nor I_50 (I3115,I3291,I775224);
not I_51 (I3404,I775224);
not I_52 (I3421,I775239);
nand I_53 (I3438,I3421,I775221);
nand I_54 (I3455,I3257,I3438);
not I_55 (I3472,I3455);
nor I_56 (I3489,I775239,I775218);
nor I_57 (I3124,I3472,I3489);
nor I_58 (I3520,I775227,I775239);
and I_59 (I3537,I3520,I3373);
nor I_60 (I3554,I3455,I3537);
DFFARX1 I_61 (I3554,I2507,I3141,I3130,);
nor I_62 (I3585,I3175,I3537);
DFFARX1 I_63 (I3585,I2507,I3141,I3127,);
nor I_64 (I3616,I775227,I775218);
DFFARX1 I_65 (I3616,I2507,I3141,I3642,);
nor I_66 (I3650,I3642,I775233);
nand I_67 (I3667,I3650,I3257);
nand I_68 (I3121,I3667,I3356);
nand I_69 (I3118,I3650,I3404);
not I_70 (I3736,I2514);
DFFARX1 I_71 (I740562,I2507,I3736,I3762,);
nand I_72 (I3770,I3762,I740541);
not I_73 (I3787,I3770);
DFFARX1 I_74 (I3787,I2507,I3736,I3728,);
DFFARX1 I_75 (I740550,I2507,I3736,I3827,);
not I_76 (I3835,I3827);
not I_77 (I3852,I740556);
not I_78 (I3869,I740553);
nand I_79 (I3886,I3835,I3869);
nor I_80 (I3903,I3886,I740556);
DFFARX1 I_81 (I3903,I2507,I3736,I3707,);
nor I_82 (I3934,I740553,I740556);
nand I_83 (I3951,I3827,I3934);
nor I_84 (I3968,I740544,I740538);
nor I_85 (I3710,I3886,I740544);
not I_86 (I3999,I740544);
not I_87 (I4016,I740559);
nand I_88 (I4033,I4016,I740541);
nand I_89 (I4050,I3852,I4033);
not I_90 (I4067,I4050);
nor I_91 (I4084,I740559,I740538);
nor I_92 (I3719,I4067,I4084);
nor I_93 (I4115,I740547,I740559);
and I_94 (I4132,I4115,I3968);
nor I_95 (I4149,I4050,I4132);
DFFARX1 I_96 (I4149,I2507,I3736,I3725,);
nor I_97 (I4180,I3770,I4132);
DFFARX1 I_98 (I4180,I2507,I3736,I3722,);
nor I_99 (I4211,I740547,I740538);
DFFARX1 I_100 (I4211,I2507,I3736,I4237,);
nor I_101 (I4245,I4237,I740553);
nand I_102 (I4262,I4245,I3852);
nand I_103 (I3716,I4262,I3951);
nand I_104 (I3713,I4245,I3999);
not I_105 (I4331,I2514);
DFFARX1 I_106 (I696634,I2507,I4331,I4357,);
nand I_107 (I4365,I4357,I696613);
not I_108 (I4382,I4365);
DFFARX1 I_109 (I4382,I2507,I4331,I4323,);
DFFARX1 I_110 (I696622,I2507,I4331,I4422,);
not I_111 (I4430,I4422);
not I_112 (I4447,I696628);
not I_113 (I4464,I696625);
nand I_114 (I4481,I4430,I4464);
nor I_115 (I4498,I4481,I696628);
DFFARX1 I_116 (I4498,I2507,I4331,I4302,);
nor I_117 (I4529,I696625,I696628);
nand I_118 (I4546,I4422,I4529);
nor I_119 (I4563,I696616,I696610);
nor I_120 (I4305,I4481,I696616);
not I_121 (I4594,I696616);
not I_122 (I4611,I696631);
nand I_123 (I4628,I4611,I696613);
nand I_124 (I4645,I4447,I4628);
not I_125 (I4662,I4645);
nor I_126 (I4679,I696631,I696610);
nor I_127 (I4314,I4662,I4679);
nor I_128 (I4710,I696619,I696631);
and I_129 (I4727,I4710,I4563);
nor I_130 (I4744,I4645,I4727);
DFFARX1 I_131 (I4744,I2507,I4331,I4320,);
nor I_132 (I4775,I4365,I4727);
DFFARX1 I_133 (I4775,I2507,I4331,I4317,);
nor I_134 (I4806,I696619,I696610);
DFFARX1 I_135 (I4806,I2507,I4331,I4832,);
nor I_136 (I4840,I4832,I696625);
nand I_137 (I4857,I4840,I4447);
nand I_138 (I4311,I4857,I4546);
nand I_139 (I4308,I4840,I4594);
not I_140 (I4926,I2514);
DFFARX1 I_141 (I765416,I2507,I4926,I4952,);
nand I_142 (I4960,I4952,I765395);
not I_143 (I4977,I4960);
DFFARX1 I_144 (I4977,I2507,I4926,I4918,);
DFFARX1 I_145 (I765404,I2507,I4926,I5017,);
not I_146 (I5025,I5017);
not I_147 (I5042,I765410);
not I_148 (I5059,I765407);
nand I_149 (I5076,I5025,I5059);
nor I_150 (I5093,I5076,I765410);
DFFARX1 I_151 (I5093,I2507,I4926,I4897,);
nor I_152 (I5124,I765407,I765410);
nand I_153 (I5141,I5017,I5124);
nor I_154 (I5158,I765398,I765392);
nor I_155 (I4900,I5076,I765398);
not I_156 (I5189,I765398);
not I_157 (I5206,I765413);
nand I_158 (I5223,I5206,I765395);
nand I_159 (I5240,I5042,I5223);
not I_160 (I5257,I5240);
nor I_161 (I5274,I765413,I765392);
nor I_162 (I4909,I5257,I5274);
nor I_163 (I5305,I765401,I765413);
and I_164 (I5322,I5305,I5158);
nor I_165 (I5339,I5240,I5322);
DFFARX1 I_166 (I5339,I2507,I4926,I4915,);
nor I_167 (I5370,I4960,I5322);
DFFARX1 I_168 (I5370,I2507,I4926,I4912,);
nor I_169 (I5401,I765401,I765392);
DFFARX1 I_170 (I5401,I2507,I4926,I5427,);
nor I_171 (I5435,I5427,I765407);
nand I_172 (I5452,I5435,I5042);
nand I_173 (I4906,I5452,I5141);
nand I_174 (I4903,I5435,I5189);
not I_175 (I5521,I2514);
DFFARX1 I_176 (I1043246,I2507,I5521,I5547,);
nand I_177 (I5555,I5547,I1043258);
not I_178 (I5572,I5555);
DFFARX1 I_179 (I5572,I2507,I5521,I5513,);
DFFARX1 I_180 (I1043243,I2507,I5521,I5612,);
not I_181 (I5620,I5612);
not I_182 (I5637,I1043246);
not I_183 (I5654,I1043240);
nand I_184 (I5671,I5620,I5654);
nor I_185 (I5688,I5671,I1043246);
DFFARX1 I_186 (I5688,I2507,I5521,I5492,);
nor I_187 (I5719,I1043240,I1043246);
nand I_188 (I5736,I5612,I5719);
nor I_189 (I5753,I1043249,I1043243);
nor I_190 (I5495,I5671,I1043249);
not I_191 (I5784,I1043249);
not I_192 (I5801,I1043255);
nand I_193 (I5818,I5801,I1043240);
nand I_194 (I5835,I5637,I5818);
not I_195 (I5852,I5835);
nor I_196 (I5869,I1043255,I1043243);
nor I_197 (I5504,I5852,I5869);
nor I_198 (I5900,I1043252,I1043255);
and I_199 (I5917,I5900,I5753);
nor I_200 (I5934,I5835,I5917);
DFFARX1 I_201 (I5934,I2507,I5521,I5510,);
nor I_202 (I5965,I5555,I5917);
DFFARX1 I_203 (I5965,I2507,I5521,I5507,);
nor I_204 (I5996,I1043252,I1043261);
DFFARX1 I_205 (I5996,I2507,I5521,I6022,);
nor I_206 (I6030,I6022,I1043240);
nand I_207 (I6047,I6030,I5637);
nand I_208 (I5501,I6047,I5736);
nand I_209 (I5498,I6030,I5784);
not I_210 (I6116,I2514);
DFFARX1 I_211 (I48548,I2507,I6116,I6142,);
nand I_212 (I6150,I6142,I48539);
not I_213 (I6167,I6150);
DFFARX1 I_214 (I6167,I2507,I6116,I6108,);
DFFARX1 I_215 (I48560,I2507,I6116,I6207,);
not I_216 (I6215,I6207);
not I_217 (I6232,I48536);
not I_218 (I6249,I48536);
nand I_219 (I6266,I6215,I6249);
nor I_220 (I6283,I6266,I48536);
DFFARX1 I_221 (I6283,I2507,I6116,I6087,);
nor I_222 (I6314,I48536,I48536);
nand I_223 (I6331,I6207,I6314);
nor I_224 (I6348,I48545,I48539);
nor I_225 (I6090,I6266,I48545);
not I_226 (I6379,I48545);
not I_227 (I6396,I48557);
nand I_228 (I6413,I6396,I48554);
nand I_229 (I6430,I6232,I6413);
not I_230 (I6447,I6430);
nor I_231 (I6464,I48557,I48539);
nor I_232 (I6099,I6447,I6464);
nor I_233 (I6495,I48551,I48557);
and I_234 (I6512,I6495,I6348);
nor I_235 (I6529,I6430,I6512);
DFFARX1 I_236 (I6529,I2507,I6116,I6105,);
nor I_237 (I6560,I6150,I6512);
DFFARX1 I_238 (I6560,I2507,I6116,I6102,);
nor I_239 (I6591,I48551,I48542);
DFFARX1 I_240 (I6591,I2507,I6116,I6617,);
nor I_241 (I6625,I6617,I48536);
nand I_242 (I6642,I6625,I6232);
nand I_243 (I6096,I6642,I6331);
nand I_244 (I6093,I6625,I6379);
not I_245 (I6711,I2514);
DFFARX1 I_246 (I359294,I2507,I6711,I6737,);
nand I_247 (I6745,I6737,I359285);
not I_248 (I6762,I6745);
DFFARX1 I_249 (I6762,I2507,I6711,I6703,);
DFFARX1 I_250 (I359288,I2507,I6711,I6802,);
not I_251 (I6810,I6802);
not I_252 (I6827,I359282);
not I_253 (I6844,I359291);
nand I_254 (I6861,I6810,I6844);
nor I_255 (I6878,I6861,I359282);
DFFARX1 I_256 (I6878,I2507,I6711,I6682,);
nor I_257 (I6909,I359291,I359282);
nand I_258 (I6926,I6802,I6909);
nor I_259 (I6943,I359279,I359297);
nor I_260 (I6685,I6861,I359279);
not I_261 (I6974,I359279);
not I_262 (I6991,I359279);
nand I_263 (I7008,I6991,I359303);
nand I_264 (I7025,I6827,I7008);
not I_265 (I7042,I7025);
nor I_266 (I7059,I359279,I359297);
nor I_267 (I6694,I7042,I7059);
nor I_268 (I7090,I359300,I359279);
and I_269 (I7107,I7090,I6943);
nor I_270 (I7124,I7025,I7107);
DFFARX1 I_271 (I7124,I2507,I6711,I6700,);
nor I_272 (I7155,I6745,I7107);
DFFARX1 I_273 (I7155,I2507,I6711,I6697,);
nor I_274 (I7186,I359300,I359306);
DFFARX1 I_275 (I7186,I2507,I6711,I7212,);
nor I_276 (I7220,I7212,I359291);
nand I_277 (I7237,I7220,I6827);
nand I_278 (I6691,I7237,I6926);
nand I_279 (I6688,I7220,I6974);
not I_280 (I7306,I2514);
DFFARX1 I_281 (I273393,I2507,I7306,I7332,);
nand I_282 (I7340,I7332,I273384);
not I_283 (I7357,I7340);
DFFARX1 I_284 (I7357,I2507,I7306,I7298,);
DFFARX1 I_285 (I273387,I2507,I7306,I7397,);
not I_286 (I7405,I7397);
not I_287 (I7422,I273381);
not I_288 (I7439,I273390);
nand I_289 (I7456,I7405,I7439);
nor I_290 (I7473,I7456,I273381);
DFFARX1 I_291 (I7473,I2507,I7306,I7277,);
nor I_292 (I7504,I273390,I273381);
nand I_293 (I7521,I7397,I7504);
nor I_294 (I7538,I273378,I273396);
nor I_295 (I7280,I7456,I273378);
not I_296 (I7569,I273378);
not I_297 (I7586,I273378);
nand I_298 (I7603,I7586,I273402);
nand I_299 (I7620,I7422,I7603);
not I_300 (I7637,I7620);
nor I_301 (I7654,I273378,I273396);
nor I_302 (I7289,I7637,I7654);
nor I_303 (I7685,I273399,I273378);
and I_304 (I7702,I7685,I7538);
nor I_305 (I7719,I7620,I7702);
DFFARX1 I_306 (I7719,I2507,I7306,I7295,);
nor I_307 (I7750,I7340,I7702);
DFFARX1 I_308 (I7750,I2507,I7306,I7292,);
nor I_309 (I7781,I273399,I273405);
DFFARX1 I_310 (I7781,I2507,I7306,I7807,);
nor I_311 (I7815,I7807,I273390);
nand I_312 (I7832,I7815,I7422);
nand I_313 (I7286,I7832,I7521);
nand I_314 (I7283,I7815,I7569);
not I_315 (I7901,I2514);
DFFARX1 I_316 (I854430,I2507,I7901,I7927,);
nand I_317 (I7935,I7927,I854421);
not I_318 (I7952,I7935);
DFFARX1 I_319 (I7952,I2507,I7901,I7893,);
DFFARX1 I_320 (I854427,I2507,I7901,I7992,);
not I_321 (I8000,I7992);
not I_322 (I8017,I854421);
not I_323 (I8034,I854433);
nand I_324 (I8051,I8000,I8034);
nor I_325 (I8068,I8051,I854421);
DFFARX1 I_326 (I8068,I2507,I7901,I7872,);
nor I_327 (I8099,I854433,I854421);
nand I_328 (I8116,I7992,I8099);
nor I_329 (I8133,I854442,I854439);
nor I_330 (I7875,I8051,I854442);
not I_331 (I8164,I854442);
not I_332 (I8181,I854427);
nand I_333 (I8198,I8181,I854424);
nand I_334 (I8215,I8017,I8198);
not I_335 (I8232,I8215);
nor I_336 (I8249,I854427,I854439);
nor I_337 (I7884,I8232,I8249);
nor I_338 (I8280,I854424,I854427);
and I_339 (I8297,I8280,I8133);
nor I_340 (I8314,I8215,I8297);
DFFARX1 I_341 (I8314,I2507,I7901,I7890,);
nor I_342 (I8345,I7935,I8297);
DFFARX1 I_343 (I8345,I2507,I7901,I7887,);
nor I_344 (I8376,I854424,I854436);
DFFARX1 I_345 (I8376,I2507,I7901,I8402,);
nor I_346 (I8410,I8402,I854433);
nand I_347 (I8427,I8410,I8017);
nand I_348 (I7881,I8427,I8116);
nand I_349 (I7878,I8410,I8164);
not I_350 (I8496,I2514);
DFFARX1 I_351 (I604133,I2507,I8496,I8522,);
nand I_352 (I8530,I8522,I604151);
not I_353 (I8547,I8530);
DFFARX1 I_354 (I8547,I2507,I8496,I8488,);
DFFARX1 I_355 (I604145,I2507,I8496,I8587,);
not I_356 (I8595,I8587);
not I_357 (I8612,I604136);
not I_358 (I8629,I604133);
nand I_359 (I8646,I8595,I8629);
nor I_360 (I8663,I8646,I604136);
DFFARX1 I_361 (I8663,I2507,I8496,I8467,);
nor I_362 (I8694,I604133,I604136);
nand I_363 (I8711,I8587,I8694);
nor I_364 (I8728,I604142,I604130);
nor I_365 (I8470,I8646,I604142);
not I_366 (I8759,I604142);
not I_367 (I8776,I604148);
nand I_368 (I8793,I8776,I604154);
nand I_369 (I8810,I8612,I8793);
not I_370 (I8827,I8810);
nor I_371 (I8844,I604148,I604130);
nor I_372 (I8479,I8827,I8844);
nor I_373 (I8875,I604130,I604148);
and I_374 (I8892,I8875,I8728);
nor I_375 (I8909,I8810,I8892);
DFFARX1 I_376 (I8909,I2507,I8496,I8485,);
nor I_377 (I8940,I8530,I8892);
DFFARX1 I_378 (I8940,I2507,I8496,I8482,);
nor I_379 (I8971,I604130,I604139);
DFFARX1 I_380 (I8971,I2507,I8496,I8997,);
nor I_381 (I9005,I8997,I604133);
nand I_382 (I9022,I9005,I8612);
nand I_383 (I8476,I9022,I8711);
nand I_384 (I8473,I9005,I8759);
not I_385 (I9091,I2514);
DFFARX1 I_386 (I600665,I2507,I9091,I9117,);
nand I_387 (I9125,I9117,I600683);
not I_388 (I9142,I9125);
DFFARX1 I_389 (I9142,I2507,I9091,I9083,);
DFFARX1 I_390 (I600677,I2507,I9091,I9182,);
not I_391 (I9190,I9182);
not I_392 (I9207,I600668);
not I_393 (I9224,I600665);
nand I_394 (I9241,I9190,I9224);
nor I_395 (I9258,I9241,I600668);
DFFARX1 I_396 (I9258,I2507,I9091,I9062,);
nor I_397 (I9289,I600665,I600668);
nand I_398 (I9306,I9182,I9289);
nor I_399 (I9323,I600674,I600662);
nor I_400 (I9065,I9241,I600674);
not I_401 (I9354,I600674);
not I_402 (I9371,I600680);
nand I_403 (I9388,I9371,I600686);
nand I_404 (I9405,I9207,I9388);
not I_405 (I9422,I9405);
nor I_406 (I9439,I600680,I600662);
nor I_407 (I9074,I9422,I9439);
nor I_408 (I9470,I600662,I600680);
and I_409 (I9487,I9470,I9323);
nor I_410 (I9504,I9405,I9487);
DFFARX1 I_411 (I9504,I2507,I9091,I9080,);
nor I_412 (I9535,I9125,I9487);
DFFARX1 I_413 (I9535,I2507,I9091,I9077,);
nor I_414 (I9566,I600662,I600671);
DFFARX1 I_415 (I9566,I2507,I9091,I9592,);
nor I_416 (I9600,I9592,I600665);
nand I_417 (I9617,I9600,I9207);
nand I_418 (I9071,I9617,I9306);
nand I_419 (I9068,I9600,I9354);
not I_420 (I9686,I2514);
DFFARX1 I_421 (I624363,I2507,I9686,I9712,);
nand I_422 (I9720,I9712,I624381);
not I_423 (I9737,I9720);
DFFARX1 I_424 (I9737,I2507,I9686,I9678,);
DFFARX1 I_425 (I624375,I2507,I9686,I9777,);
not I_426 (I9785,I9777);
not I_427 (I9802,I624366);
not I_428 (I9819,I624363);
nand I_429 (I9836,I9785,I9819);
nor I_430 (I9853,I9836,I624366);
DFFARX1 I_431 (I9853,I2507,I9686,I9657,);
nor I_432 (I9884,I624363,I624366);
nand I_433 (I9901,I9777,I9884);
nor I_434 (I9918,I624372,I624360);
nor I_435 (I9660,I9836,I624372);
not I_436 (I9949,I624372);
not I_437 (I9966,I624378);
nand I_438 (I9983,I9966,I624384);
nand I_439 (I10000,I9802,I9983);
not I_440 (I10017,I10000);
nor I_441 (I10034,I624378,I624360);
nor I_442 (I9669,I10017,I10034);
nor I_443 (I10065,I624360,I624378);
and I_444 (I10082,I10065,I9918);
nor I_445 (I10099,I10000,I10082);
DFFARX1 I_446 (I10099,I2507,I9686,I9675,);
nor I_447 (I10130,I9720,I10082);
DFFARX1 I_448 (I10130,I2507,I9686,I9672,);
nor I_449 (I10161,I624360,I624369);
DFFARX1 I_450 (I10161,I2507,I9686,I10187,);
nor I_451 (I10195,I10187,I624363);
nand I_452 (I10212,I10195,I9802);
nand I_453 (I9666,I10212,I9901);
nand I_454 (I9663,I10195,I9949);
not I_455 (I10281,I2514);
DFFARX1 I_456 (I60669,I2507,I10281,I10307,);
nand I_457 (I10315,I10307,I60660);
not I_458 (I10332,I10315);
DFFARX1 I_459 (I10332,I2507,I10281,I10273,);
DFFARX1 I_460 (I60681,I2507,I10281,I10372,);
not I_461 (I10380,I10372);
not I_462 (I10397,I60657);
not I_463 (I10414,I60657);
nand I_464 (I10431,I10380,I10414);
nor I_465 (I10448,I10431,I60657);
DFFARX1 I_466 (I10448,I2507,I10281,I10252,);
nor I_467 (I10479,I60657,I60657);
nand I_468 (I10496,I10372,I10479);
nor I_469 (I10513,I60666,I60660);
nor I_470 (I10255,I10431,I60666);
not I_471 (I10544,I60666);
not I_472 (I10561,I60678);
nand I_473 (I10578,I10561,I60675);
nand I_474 (I10595,I10397,I10578);
not I_475 (I10612,I10595);
nor I_476 (I10629,I60678,I60660);
nor I_477 (I10264,I10612,I10629);
nor I_478 (I10660,I60672,I60678);
and I_479 (I10677,I10660,I10513);
nor I_480 (I10694,I10595,I10677);
DFFARX1 I_481 (I10694,I2507,I10281,I10270,);
nor I_482 (I10725,I10315,I10677);
DFFARX1 I_483 (I10725,I2507,I10281,I10267,);
nor I_484 (I10756,I60672,I60663);
DFFARX1 I_485 (I10756,I2507,I10281,I10782,);
nor I_486 (I10790,I10782,I60657);
nand I_487 (I10807,I10790,I10397);
nand I_488 (I10261,I10807,I10496);
nand I_489 (I10258,I10790,I10544);
not I_490 (I10876,I2514);
DFFARX1 I_491 (I904388,I2507,I10876,I10902,);
nand I_492 (I10910,I10902,I904379);
not I_493 (I10927,I10910);
DFFARX1 I_494 (I10927,I2507,I10876,I10868,);
DFFARX1 I_495 (I904382,I2507,I10876,I10967,);
not I_496 (I10975,I10967);
not I_497 (I10992,I904394);
not I_498 (I11009,I904373);
nand I_499 (I11026,I10975,I11009);
nor I_500 (I11043,I11026,I904394);
DFFARX1 I_501 (I11043,I2507,I10876,I10847,);
nor I_502 (I11074,I904373,I904394);
nand I_503 (I11091,I10967,I11074);
nor I_504 (I11108,I904385,I904391);
nor I_505 (I10850,I11026,I904385);
not I_506 (I11139,I904385);
not I_507 (I11156,I904376);
nand I_508 (I11173,I11156,I904367);
nand I_509 (I11190,I10992,I11173);
not I_510 (I11207,I11190);
nor I_511 (I11224,I904376,I904391);
nor I_512 (I10859,I11207,I11224);
nor I_513 (I11255,I904367,I904376);
and I_514 (I11272,I11255,I11108);
nor I_515 (I11289,I11190,I11272);
DFFARX1 I_516 (I11289,I2507,I10876,I10865,);
nor I_517 (I11320,I10910,I11272);
DFFARX1 I_518 (I11320,I2507,I10876,I10862,);
nor I_519 (I11351,I904367,I904370);
DFFARX1 I_520 (I11351,I2507,I10876,I11377,);
nor I_521 (I11385,I11377,I904373);
nand I_522 (I11402,I11385,I10992);
nand I_523 (I10856,I11402,I11091);
nand I_524 (I10853,I11385,I11139);
not I_525 (I11471,I2514);
DFFARX1 I_526 (I383780,I2507,I11471,I11497,);
nand I_527 (I11505,I11497,I383762);
not I_528 (I11522,I11505);
DFFARX1 I_529 (I11522,I2507,I11471,I11463,);
DFFARX1 I_530 (I383774,I2507,I11471,I11562,);
not I_531 (I11570,I11562);
not I_532 (I11587,I383759);
not I_533 (I11604,I383768);
nand I_534 (I11621,I11570,I11604);
nor I_535 (I11638,I11621,I383759);
DFFARX1 I_536 (I11638,I2507,I11471,I11442,);
nor I_537 (I11669,I383768,I383759);
nand I_538 (I11686,I11562,I11669);
nor I_539 (I11703,I383765,I383786);
nor I_540 (I11445,I11621,I383765);
not I_541 (I11734,I383765);
not I_542 (I11751,I383777);
nand I_543 (I11768,I11751,I383783);
nand I_544 (I11785,I11587,I11768);
not I_545 (I11802,I11785);
nor I_546 (I11819,I383777,I383786);
nor I_547 (I11454,I11802,I11819);
nor I_548 (I11850,I383759,I383777);
and I_549 (I11867,I11850,I11703);
nor I_550 (I11884,I11785,I11867);
DFFARX1 I_551 (I11884,I2507,I11471,I11460,);
nor I_552 (I11915,I11505,I11867);
DFFARX1 I_553 (I11915,I2507,I11471,I11457,);
nor I_554 (I11946,I383759,I383771);
DFFARX1 I_555 (I11946,I2507,I11471,I11972,);
nor I_556 (I11980,I11972,I383768);
nand I_557 (I11997,I11980,I11587);
nand I_558 (I11451,I11997,I11686);
nand I_559 (I11448,I11980,I11734);
not I_560 (I12066,I2514);
DFFARX1 I_561 (I2308,I2507,I12066,I12092,);
nand I_562 (I12100,I12092,I2500);
not I_563 (I12117,I12100);
DFFARX1 I_564 (I12117,I2507,I12066,I12058,);
DFFARX1 I_565 (I1660,I2507,I12066,I12157,);
not I_566 (I12165,I12157);
not I_567 (I12182,I2316);
not I_568 (I12199,I1812);
nand I_569 (I12216,I12165,I12199);
nor I_570 (I12233,I12216,I2316);
DFFARX1 I_571 (I12233,I2507,I12066,I12037,);
nor I_572 (I12264,I1812,I2316);
nand I_573 (I12281,I12157,I12264);
nor I_574 (I12298,I1444,I1468);
nor I_575 (I12040,I12216,I1444);
not I_576 (I12329,I1444);
not I_577 (I12346,I2052);
nand I_578 (I12363,I12346,I1364);
nand I_579 (I12380,I12182,I12363);
not I_580 (I12397,I12380);
nor I_581 (I12414,I2052,I1468);
nor I_582 (I12049,I12397,I12414);
nor I_583 (I12445,I2300,I2052);
and I_584 (I12462,I12445,I12298);
nor I_585 (I12479,I12380,I12462);
DFFARX1 I_586 (I12479,I2507,I12066,I12055,);
nor I_587 (I12510,I12100,I12462);
DFFARX1 I_588 (I12510,I2507,I12066,I12052,);
nor I_589 (I12541,I2300,I1924);
DFFARX1 I_590 (I12541,I2507,I12066,I12567,);
nor I_591 (I12575,I12567,I1812);
nand I_592 (I12592,I12575,I12182);
nand I_593 (I12046,I12592,I12281);
nand I_594 (I12043,I12575,I12329);
not I_595 (I12661,I2514);
DFFARX1 I_596 (I903096,I2507,I12661,I12687,);
nand I_597 (I12695,I12687,I903087);
not I_598 (I12712,I12695);
DFFARX1 I_599 (I12712,I2507,I12661,I12653,);
DFFARX1 I_600 (I903090,I2507,I12661,I12752,);
not I_601 (I12760,I12752);
not I_602 (I12777,I903102);
not I_603 (I12794,I903081);
nand I_604 (I12811,I12760,I12794);
nor I_605 (I12828,I12811,I903102);
DFFARX1 I_606 (I12828,I2507,I12661,I12632,);
nor I_607 (I12859,I903081,I903102);
nand I_608 (I12876,I12752,I12859);
nor I_609 (I12893,I903093,I903099);
nor I_610 (I12635,I12811,I903093);
not I_611 (I12924,I903093);
not I_612 (I12941,I903084);
nand I_613 (I12958,I12941,I903075);
nand I_614 (I12975,I12777,I12958);
not I_615 (I12992,I12975);
nor I_616 (I13009,I903084,I903099);
nor I_617 (I12644,I12992,I13009);
nor I_618 (I13040,I903075,I903084);
and I_619 (I13057,I13040,I12893);
nor I_620 (I13074,I12975,I13057);
DFFARX1 I_621 (I13074,I2507,I12661,I12650,);
nor I_622 (I13105,I12695,I13057);
DFFARX1 I_623 (I13105,I2507,I12661,I12647,);
nor I_624 (I13136,I903075,I903078);
DFFARX1 I_625 (I13136,I2507,I12661,I13162,);
nor I_626 (I13170,I13162,I903081);
nand I_627 (I13187,I13170,I12777);
nand I_628 (I12641,I13187,I12876);
nand I_629 (I12638,I13170,I12924);
not I_630 (I13259,I2514);
DFFARX1 I_631 (I224016,I2507,I13259,I13285,);
DFFARX1 I_632 (I13285,I2507,I13259,I13302,);
not I_633 (I13310,I13302);
nand I_634 (I13327,I224034,I224019);
and I_635 (I13344,I13327,I224022);
DFFARX1 I_636 (I13344,I2507,I13259,I13370,);
DFFARX1 I_637 (I13370,I2507,I13259,I13251,);
DFFARX1 I_638 (I13370,I2507,I13259,I13242,);
DFFARX1 I_639 (I224010,I2507,I13259,I13415,);
nand I_640 (I13423,I13415,I224013);
not I_641 (I13440,I13423);
nor I_642 (I13239,I13285,I13440);
DFFARX1 I_643 (I224025,I2507,I13259,I13480,);
not I_644 (I13488,I13480);
nor I_645 (I13245,I13488,I13310);
nand I_646 (I13233,I13488,I13423);
nand I_647 (I13533,I224031,I224028);
and I_648 (I13550,I13533,I224013);
DFFARX1 I_649 (I13550,I2507,I13259,I13576,);
nor I_650 (I13584,I13576,I13285);
DFFARX1 I_651 (I13584,I2507,I13259,I13227,);
not I_652 (I13615,I13576);
nor I_653 (I13632,I224010,I224028);
not I_654 (I13649,I13632);
nor I_655 (I13666,I13423,I13649);
nor I_656 (I13683,I13615,I13666);
DFFARX1 I_657 (I13683,I2507,I13259,I13248,);
nor I_658 (I13714,I13576,I13649);
nor I_659 (I13236,I13440,I13714);
nor I_660 (I13230,I13576,I13632);
not I_661 (I13786,I2514);
DFFARX1 I_662 (I1039880,I2507,I13786,I13812,);
DFFARX1 I_663 (I13812,I2507,I13786,I13829,);
not I_664 (I13837,I13829);
nand I_665 (I13854,I1039874,I1039895);
and I_666 (I13871,I13854,I1039880);
DFFARX1 I_667 (I13871,I2507,I13786,I13897,);
DFFARX1 I_668 (I13897,I2507,I13786,I13778,);
DFFARX1 I_669 (I13897,I2507,I13786,I13769,);
DFFARX1 I_670 (I1039877,I2507,I13786,I13942,);
nand I_671 (I13950,I13942,I1039886);
not I_672 (I13967,I13950);
nor I_673 (I13766,I13812,I13967);
DFFARX1 I_674 (I1039874,I2507,I13786,I14007,);
not I_675 (I14015,I14007);
nor I_676 (I13772,I14015,I13837);
nand I_677 (I13760,I14015,I13950);
nand I_678 (I14060,I1039877,I1039892);
and I_679 (I14077,I14060,I1039883);
DFFARX1 I_680 (I14077,I2507,I13786,I14103,);
nor I_681 (I14111,I14103,I13812);
DFFARX1 I_682 (I14111,I2507,I13786,I13754,);
not I_683 (I14142,I14103);
nor I_684 (I14159,I1039889,I1039892);
not I_685 (I14176,I14159);
nor I_686 (I14193,I13950,I14176);
nor I_687 (I14210,I14142,I14193);
DFFARX1 I_688 (I14210,I2507,I13786,I13775,);
nor I_689 (I14241,I14103,I14176);
nor I_690 (I13763,I13967,I14241);
nor I_691 (I13757,I14103,I14159);
not I_692 (I14313,I2514);
DFFARX1 I_693 (I859700,I2507,I14313,I14339,);
DFFARX1 I_694 (I14339,I2507,I14313,I14356,);
not I_695 (I14364,I14356);
nand I_696 (I14381,I859691,I859712);
and I_697 (I14398,I14381,I859694);
DFFARX1 I_698 (I14398,I2507,I14313,I14424,);
DFFARX1 I_699 (I14424,I2507,I14313,I14305,);
DFFARX1 I_700 (I14424,I2507,I14313,I14296,);
DFFARX1 I_701 (I859694,I2507,I14313,I14469,);
nand I_702 (I14477,I14469,I859709);
not I_703 (I14494,I14477);
nor I_704 (I14293,I14339,I14494);
DFFARX1 I_705 (I859703,I2507,I14313,I14534,);
not I_706 (I14542,I14534);
nor I_707 (I14299,I14542,I14364);
nand I_708 (I14287,I14542,I14477);
nand I_709 (I14587,I859697,I859706);
and I_710 (I14604,I14587,I859691);
DFFARX1 I_711 (I14604,I2507,I14313,I14630,);
nor I_712 (I14638,I14630,I14339);
DFFARX1 I_713 (I14638,I2507,I14313,I14281,);
not I_714 (I14669,I14630);
nor I_715 (I14686,I859697,I859706);
not I_716 (I14703,I14686);
nor I_717 (I14720,I14477,I14703);
nor I_718 (I14737,I14669,I14720);
DFFARX1 I_719 (I14737,I2507,I14313,I14302,);
nor I_720 (I14768,I14630,I14703);
nor I_721 (I14290,I14494,I14768);
nor I_722 (I14284,I14630,I14686);
not I_723 (I14840,I2514);
DFFARX1 I_724 (I53282,I2507,I14840,I14866,);
DFFARX1 I_725 (I14866,I2507,I14840,I14883,);
not I_726 (I14891,I14883);
nand I_727 (I14908,I53282,I53297);
and I_728 (I14925,I14908,I53300);
DFFARX1 I_729 (I14925,I2507,I14840,I14951,);
DFFARX1 I_730 (I14951,I2507,I14840,I14832,);
DFFARX1 I_731 (I14951,I2507,I14840,I14823,);
DFFARX1 I_732 (I53294,I2507,I14840,I14996,);
nand I_733 (I15004,I14996,I53303);
not I_734 (I15021,I15004);
nor I_735 (I14820,I14866,I15021);
DFFARX1 I_736 (I53279,I2507,I14840,I15061,);
not I_737 (I15069,I15061);
nor I_738 (I14826,I15069,I14891);
nand I_739 (I14814,I15069,I15004);
nand I_740 (I15114,I53279,I53285);
and I_741 (I15131,I15114,I53288);
DFFARX1 I_742 (I15131,I2507,I14840,I15157,);
nor I_743 (I15165,I15157,I14866);
DFFARX1 I_744 (I15165,I2507,I14840,I14808,);
not I_745 (I15196,I15157);
nor I_746 (I15213,I53291,I53285);
not I_747 (I15230,I15213);
nor I_748 (I15247,I15004,I15230);
nor I_749 (I15264,I15196,I15247);
DFFARX1 I_750 (I15264,I2507,I14840,I14829,);
nor I_751 (I15295,I15157,I15230);
nor I_752 (I14817,I15021,I15295);
nor I_753 (I14811,I15157,I15213);
not I_754 (I15367,I2514);
DFFARX1 I_755 (I1136424,I2507,I15367,I15393,);
DFFARX1 I_756 (I15393,I2507,I15367,I15410,);
not I_757 (I15418,I15410);
nand I_758 (I15435,I1136412,I1136403);
and I_759 (I15452,I15435,I1136400);
DFFARX1 I_760 (I15452,I2507,I15367,I15478,);
DFFARX1 I_761 (I15478,I2507,I15367,I15359,);
DFFARX1 I_762 (I15478,I2507,I15367,I15350,);
DFFARX1 I_763 (I1136406,I2507,I15367,I15523,);
nand I_764 (I15531,I15523,I1136418);
not I_765 (I15548,I15531);
nor I_766 (I15347,I15393,I15548);
DFFARX1 I_767 (I1136415,I2507,I15367,I15588,);
not I_768 (I15596,I15588);
nor I_769 (I15353,I15596,I15418);
nand I_770 (I15341,I15596,I15531);
nand I_771 (I15641,I1136409,I1136403);
and I_772 (I15658,I15641,I1136421);
DFFARX1 I_773 (I15658,I2507,I15367,I15684,);
nor I_774 (I15692,I15684,I15393);
DFFARX1 I_775 (I15692,I2507,I15367,I15335,);
not I_776 (I15723,I15684);
nor I_777 (I15740,I1136400,I1136403);
not I_778 (I15757,I15740);
nor I_779 (I15774,I15531,I15757);
nor I_780 (I15791,I15723,I15774);
DFFARX1 I_781 (I15791,I2507,I15367,I15356,);
nor I_782 (I15822,I15684,I15757);
nor I_783 (I15344,I15548,I15822);
nor I_784 (I15338,I15684,I15740);
not I_785 (I15894,I2514);
DFFARX1 I_786 (I205571,I2507,I15894,I15920,);
DFFARX1 I_787 (I15920,I2507,I15894,I15937,);
not I_788 (I15945,I15937);
nand I_789 (I15962,I205589,I205574);
and I_790 (I15979,I15962,I205577);
DFFARX1 I_791 (I15979,I2507,I15894,I16005,);
DFFARX1 I_792 (I16005,I2507,I15894,I15886,);
DFFARX1 I_793 (I16005,I2507,I15894,I15877,);
DFFARX1 I_794 (I205565,I2507,I15894,I16050,);
nand I_795 (I16058,I16050,I205568);
not I_796 (I16075,I16058);
nor I_797 (I15874,I15920,I16075);
DFFARX1 I_798 (I205580,I2507,I15894,I16115,);
not I_799 (I16123,I16115);
nor I_800 (I15880,I16123,I15945);
nand I_801 (I15868,I16123,I16058);
nand I_802 (I16168,I205586,I205583);
and I_803 (I16185,I16168,I205568);
DFFARX1 I_804 (I16185,I2507,I15894,I16211,);
nor I_805 (I16219,I16211,I15920);
DFFARX1 I_806 (I16219,I2507,I15894,I15862,);
not I_807 (I16250,I16211);
nor I_808 (I16267,I205565,I205583);
not I_809 (I16284,I16267);
nor I_810 (I16301,I16058,I16284);
nor I_811 (I16318,I16250,I16301);
DFFARX1 I_812 (I16318,I2507,I15894,I15883,);
nor I_813 (I16349,I16211,I16284);
nor I_814 (I15871,I16075,I16349);
nor I_815 (I15865,I16211,I16267);
not I_816 (I16421,I2514);
DFFARX1 I_817 (I649220,I2507,I16421,I16447,);
DFFARX1 I_818 (I16447,I2507,I16421,I16464,);
not I_819 (I16472,I16464);
nand I_820 (I16489,I649235,I649238);
and I_821 (I16506,I16489,I649217);
DFFARX1 I_822 (I16506,I2507,I16421,I16532,);
DFFARX1 I_823 (I16532,I2507,I16421,I16413,);
DFFARX1 I_824 (I16532,I2507,I16421,I16404,);
DFFARX1 I_825 (I649223,I2507,I16421,I16577,);
nand I_826 (I16585,I16577,I649229);
not I_827 (I16602,I16585);
nor I_828 (I16401,I16447,I16602);
DFFARX1 I_829 (I649217,I2507,I16421,I16642,);
not I_830 (I16650,I16642);
nor I_831 (I16407,I16650,I16472);
nand I_832 (I16395,I16650,I16585);
nand I_833 (I16695,I649232,I649214);
and I_834 (I16712,I16695,I649226);
DFFARX1 I_835 (I16712,I2507,I16421,I16738,);
nor I_836 (I16746,I16738,I16447);
DFFARX1 I_837 (I16746,I2507,I16421,I16389,);
not I_838 (I16777,I16738);
nor I_839 (I16794,I649214,I649214);
not I_840 (I16811,I16794);
nor I_841 (I16828,I16585,I16811);
nor I_842 (I16845,I16777,I16828);
DFFARX1 I_843 (I16845,I2507,I16421,I16410,);
nor I_844 (I16876,I16738,I16811);
nor I_845 (I16398,I16602,I16876);
nor I_846 (I16392,I16738,I16794);
not I_847 (I16948,I2514);
DFFARX1 I_848 (I818594,I2507,I16948,I16974,);
DFFARX1 I_849 (I16974,I2507,I16948,I16991,);
not I_850 (I16999,I16991);
nand I_851 (I17016,I818585,I818606);
and I_852 (I17033,I17016,I818588);
DFFARX1 I_853 (I17033,I2507,I16948,I17059,);
DFFARX1 I_854 (I17059,I2507,I16948,I16940,);
DFFARX1 I_855 (I17059,I2507,I16948,I16931,);
DFFARX1 I_856 (I818588,I2507,I16948,I17104,);
nand I_857 (I17112,I17104,I818603);
not I_858 (I17129,I17112);
nor I_859 (I16928,I16974,I17129);
DFFARX1 I_860 (I818597,I2507,I16948,I17169,);
not I_861 (I17177,I17169);
nor I_862 (I16934,I17177,I16999);
nand I_863 (I16922,I17177,I17112);
nand I_864 (I17222,I818591,I818600);
and I_865 (I17239,I17222,I818585);
DFFARX1 I_866 (I17239,I2507,I16948,I17265,);
nor I_867 (I17273,I17265,I16974);
DFFARX1 I_868 (I17273,I2507,I16948,I16916,);
not I_869 (I17304,I17265);
nor I_870 (I17321,I818591,I818600);
not I_871 (I17338,I17321);
nor I_872 (I17355,I17112,I17338);
nor I_873 (I17372,I17304,I17355);
DFFARX1 I_874 (I17372,I2507,I16948,I16937,);
nor I_875 (I17403,I17265,I17338);
nor I_876 (I16925,I17129,I17403);
nor I_877 (I16919,I17265,I17321);
not I_878 (I17475,I2514);
DFFARX1 I_879 (I853903,I2507,I17475,I17501,);
DFFARX1 I_880 (I17501,I2507,I17475,I17518,);
not I_881 (I17526,I17518);
nand I_882 (I17543,I853894,I853915);
and I_883 (I17560,I17543,I853897);
DFFARX1 I_884 (I17560,I2507,I17475,I17586,);
DFFARX1 I_885 (I17586,I2507,I17475,I17467,);
DFFARX1 I_886 (I17586,I2507,I17475,I17458,);
DFFARX1 I_887 (I853897,I2507,I17475,I17631,);
nand I_888 (I17639,I17631,I853912);
not I_889 (I17656,I17639);
nor I_890 (I17455,I17501,I17656);
DFFARX1 I_891 (I853906,I2507,I17475,I17696,);
not I_892 (I17704,I17696);
nor I_893 (I17461,I17704,I17526);
nand I_894 (I17449,I17704,I17639);
nand I_895 (I17749,I853900,I853909);
and I_896 (I17766,I17749,I853894);
DFFARX1 I_897 (I17766,I2507,I17475,I17792,);
nor I_898 (I17800,I17792,I17501);
DFFARX1 I_899 (I17800,I2507,I17475,I17443,);
not I_900 (I17831,I17792);
nor I_901 (I17848,I853900,I853909);
not I_902 (I17865,I17848);
nor I_903 (I17882,I17639,I17865);
nor I_904 (I17899,I17831,I17882);
DFFARX1 I_905 (I17899,I2507,I17475,I17464,);
nor I_906 (I17930,I17792,I17865);
nor I_907 (I17452,I17656,I17930);
nor I_908 (I17446,I17792,I17848);
not I_909 (I18002,I2514);
DFFARX1 I_910 (I375643,I2507,I18002,I18028,);
DFFARX1 I_911 (I18028,I2507,I18002,I18045,);
not I_912 (I18053,I18045);
nand I_913 (I18070,I375640,I375634);
and I_914 (I18087,I18070,I375628);
DFFARX1 I_915 (I18087,I2507,I18002,I18113,);
DFFARX1 I_916 (I18113,I2507,I18002,I17994,);
DFFARX1 I_917 (I18113,I2507,I18002,I17985,);
DFFARX1 I_918 (I375616,I2507,I18002,I18158,);
nand I_919 (I18166,I18158,I375625);
not I_920 (I18183,I18166);
nor I_921 (I17982,I18028,I18183);
DFFARX1 I_922 (I375622,I2507,I18002,I18223,);
not I_923 (I18231,I18223);
nor I_924 (I17988,I18231,I18053);
nand I_925 (I17976,I18231,I18166);
nand I_926 (I18276,I375619,I375637);
and I_927 (I18293,I18276,I375616);
DFFARX1 I_928 (I18293,I2507,I18002,I18319,);
nor I_929 (I18327,I18319,I18028);
DFFARX1 I_930 (I18327,I2507,I18002,I17970,);
not I_931 (I18358,I18319);
nor I_932 (I18375,I375631,I375637);
not I_933 (I18392,I18375);
nor I_934 (I18409,I18166,I18392);
nor I_935 (I18426,I18358,I18409);
DFFARX1 I_936 (I18426,I2507,I18002,I17991,);
nor I_937 (I18457,I18319,I18392);
nor I_938 (I17979,I18183,I18457);
nor I_939 (I17973,I18319,I18375);
not I_940 (I18529,I2514);
DFFARX1 I_941 (I493103,I2507,I18529,I18555,);
DFFARX1 I_942 (I18555,I2507,I18529,I18572,);
not I_943 (I18580,I18572);
nand I_944 (I18597,I493103,I493106);
and I_945 (I18614,I18597,I493127);
DFFARX1 I_946 (I18614,I2507,I18529,I18640,);
DFFARX1 I_947 (I18640,I2507,I18529,I18521,);
DFFARX1 I_948 (I18640,I2507,I18529,I18512,);
DFFARX1 I_949 (I493115,I2507,I18529,I18685,);
nand I_950 (I18693,I18685,I493118);
not I_951 (I18710,I18693);
nor I_952 (I18509,I18555,I18710);
DFFARX1 I_953 (I493124,I2507,I18529,I18750,);
not I_954 (I18758,I18750);
nor I_955 (I18515,I18758,I18580);
nand I_956 (I18503,I18758,I18693);
nand I_957 (I18803,I493121,I493109);
and I_958 (I18820,I18803,I493112);
DFFARX1 I_959 (I18820,I2507,I18529,I18846,);
nor I_960 (I18854,I18846,I18555);
DFFARX1 I_961 (I18854,I2507,I18529,I18497,);
not I_962 (I18885,I18846);
nor I_963 (I18902,I493130,I493109);
not I_964 (I18919,I18902);
nor I_965 (I18936,I18693,I18919);
nor I_966 (I18953,I18885,I18936);
DFFARX1 I_967 (I18953,I2507,I18529,I18518,);
nor I_968 (I18984,I18846,I18919);
nor I_969 (I18506,I18710,I18984);
nor I_970 (I18500,I18846,I18902);
not I_971 (I19056,I2514);
DFFARX1 I_972 (I252325,I2507,I19056,I19082,);
DFFARX1 I_973 (I19082,I2507,I19056,I19099,);
not I_974 (I19107,I19099);
nand I_975 (I19124,I252322,I252316);
and I_976 (I19141,I19124,I252310);
DFFARX1 I_977 (I19141,I2507,I19056,I19167,);
DFFARX1 I_978 (I19167,I2507,I19056,I19048,);
DFFARX1 I_979 (I19167,I2507,I19056,I19039,);
DFFARX1 I_980 (I252298,I2507,I19056,I19212,);
nand I_981 (I19220,I19212,I252307);
not I_982 (I19237,I19220);
nor I_983 (I19036,I19082,I19237);
DFFARX1 I_984 (I252304,I2507,I19056,I19277,);
not I_985 (I19285,I19277);
nor I_986 (I19042,I19285,I19107);
nand I_987 (I19030,I19285,I19220);
nand I_988 (I19330,I252301,I252319);
and I_989 (I19347,I19330,I252298);
DFFARX1 I_990 (I19347,I2507,I19056,I19373,);
nor I_991 (I19381,I19373,I19082);
DFFARX1 I_992 (I19381,I2507,I19056,I19024,);
not I_993 (I19412,I19373);
nor I_994 (I19429,I252313,I252319);
not I_995 (I19446,I19429);
nor I_996 (I19463,I19220,I19446);
nor I_997 (I19480,I19412,I19463);
DFFARX1 I_998 (I19480,I2507,I19056,I19045,);
nor I_999 (I19511,I19373,I19446);
nor I_1000 (I19033,I19237,I19511);
nor I_1001 (I19027,I19373,I19429);
not I_1002 (I19583,I2514);
DFFARX1 I_1003 (I351928,I2507,I19583,I19609,);
DFFARX1 I_1004 (I19609,I2507,I19583,I19626,);
not I_1005 (I19634,I19626);
nand I_1006 (I19651,I351925,I351919);
and I_1007 (I19668,I19651,I351913);
DFFARX1 I_1008 (I19668,I2507,I19583,I19694,);
DFFARX1 I_1009 (I19694,I2507,I19583,I19575,);
DFFARX1 I_1010 (I19694,I2507,I19583,I19566,);
DFFARX1 I_1011 (I351901,I2507,I19583,I19739,);
nand I_1012 (I19747,I19739,I351910);
not I_1013 (I19764,I19747);
nor I_1014 (I19563,I19609,I19764);
DFFARX1 I_1015 (I351907,I2507,I19583,I19804,);
not I_1016 (I19812,I19804);
nor I_1017 (I19569,I19812,I19634);
nand I_1018 (I19557,I19812,I19747);
nand I_1019 (I19857,I351904,I351922);
and I_1020 (I19874,I19857,I351901);
DFFARX1 I_1021 (I19874,I2507,I19583,I19900,);
nor I_1022 (I19908,I19900,I19609);
DFFARX1 I_1023 (I19908,I2507,I19583,I19551,);
not I_1024 (I19939,I19900);
nor I_1025 (I19956,I351916,I351922);
not I_1026 (I19973,I19956);
nor I_1027 (I19990,I19747,I19973);
nor I_1028 (I20007,I19939,I19990);
DFFARX1 I_1029 (I20007,I2507,I19583,I19572,);
nor I_1030 (I20038,I19900,I19973);
nor I_1031 (I19560,I19764,I20038);
nor I_1032 (I19554,I19900,I19956);
not I_1033 (I20110,I2514);
DFFARX1 I_1034 (I354563,I2507,I20110,I20136,);
DFFARX1 I_1035 (I20136,I2507,I20110,I20153,);
not I_1036 (I20161,I20153);
nand I_1037 (I20178,I354560,I354554);
and I_1038 (I20195,I20178,I354548);
DFFARX1 I_1039 (I20195,I2507,I20110,I20221,);
DFFARX1 I_1040 (I20221,I2507,I20110,I20102,);
DFFARX1 I_1041 (I20221,I2507,I20110,I20093,);
DFFARX1 I_1042 (I354536,I2507,I20110,I20266,);
nand I_1043 (I20274,I20266,I354545);
not I_1044 (I20291,I20274);
nor I_1045 (I20090,I20136,I20291);
DFFARX1 I_1046 (I354542,I2507,I20110,I20331,);
not I_1047 (I20339,I20331);
nor I_1048 (I20096,I20339,I20161);
nand I_1049 (I20084,I20339,I20274);
nand I_1050 (I20384,I354539,I354557);
and I_1051 (I20401,I20384,I354536);
DFFARX1 I_1052 (I20401,I2507,I20110,I20427,);
nor I_1053 (I20435,I20427,I20136);
DFFARX1 I_1054 (I20435,I2507,I20110,I20078,);
not I_1055 (I20466,I20427);
nor I_1056 (I20483,I354551,I354557);
not I_1057 (I20500,I20483);
nor I_1058 (I20517,I20274,I20500);
nor I_1059 (I20534,I20466,I20517);
DFFARX1 I_1060 (I20534,I2507,I20110,I20099,);
nor I_1061 (I20565,I20427,I20500);
nor I_1062 (I20087,I20291,I20565);
nor I_1063 (I20081,I20427,I20483);
not I_1064 (I20637,I2514);
DFFARX1 I_1065 (I90172,I2507,I20637,I20663,);
DFFARX1 I_1066 (I20663,I2507,I20637,I20680,);
not I_1067 (I20688,I20680);
nand I_1068 (I20705,I90172,I90187);
and I_1069 (I20722,I20705,I90190);
DFFARX1 I_1070 (I20722,I2507,I20637,I20748,);
DFFARX1 I_1071 (I20748,I2507,I20637,I20629,);
DFFARX1 I_1072 (I20748,I2507,I20637,I20620,);
DFFARX1 I_1073 (I90184,I2507,I20637,I20793,);
nand I_1074 (I20801,I20793,I90193);
not I_1075 (I20818,I20801);
nor I_1076 (I20617,I20663,I20818);
DFFARX1 I_1077 (I90169,I2507,I20637,I20858,);
not I_1078 (I20866,I20858);
nor I_1079 (I20623,I20866,I20688);
nand I_1080 (I20611,I20866,I20801);
nand I_1081 (I20911,I90169,I90175);
and I_1082 (I20928,I20911,I90178);
DFFARX1 I_1083 (I20928,I2507,I20637,I20954,);
nor I_1084 (I20962,I20954,I20663);
DFFARX1 I_1085 (I20962,I2507,I20637,I20605,);
not I_1086 (I20993,I20954);
nor I_1087 (I21010,I90181,I90175);
not I_1088 (I21027,I21010);
nor I_1089 (I21044,I20801,I21027);
nor I_1090 (I21061,I20993,I21044);
DFFARX1 I_1091 (I21061,I2507,I20637,I20626,);
nor I_1092 (I21092,I20954,I21027);
nor I_1093 (I20614,I20818,I21092);
nor I_1094 (I20608,I20954,I21010);
not I_1095 (I21164,I2514);
DFFARX1 I_1096 (I1300882,I2507,I21164,I21190,);
DFFARX1 I_1097 (I21190,I2507,I21164,I21207,);
not I_1098 (I21215,I21207);
nand I_1099 (I21232,I1300873,I1300879);
and I_1100 (I21249,I21232,I1300858);
DFFARX1 I_1101 (I21249,I2507,I21164,I21275,);
DFFARX1 I_1102 (I21275,I2507,I21164,I21156,);
DFFARX1 I_1103 (I21275,I2507,I21164,I21147,);
DFFARX1 I_1104 (I1300876,I2507,I21164,I21320,);
nand I_1105 (I21328,I21320,I1300858);
not I_1106 (I21345,I21328);
nor I_1107 (I21144,I21190,I21345);
DFFARX1 I_1108 (I1300870,I2507,I21164,I21385,);
not I_1109 (I21393,I21385);
nor I_1110 (I21150,I21393,I21215);
nand I_1111 (I21138,I21393,I21328);
nand I_1112 (I21438,I1300864,I1300885);
and I_1113 (I21455,I21438,I1300867);
DFFARX1 I_1114 (I21455,I2507,I21164,I21481,);
nor I_1115 (I21489,I21481,I21190);
DFFARX1 I_1116 (I21489,I2507,I21164,I21132,);
not I_1117 (I21520,I21481);
nor I_1118 (I21537,I1300861,I1300885);
not I_1119 (I21554,I21537);
nor I_1120 (I21571,I21328,I21554);
nor I_1121 (I21588,I21520,I21571);
DFFARX1 I_1122 (I21588,I2507,I21164,I21153,);
nor I_1123 (I21619,I21481,I21554);
nor I_1124 (I21141,I21345,I21619);
nor I_1125 (I21135,I21481,I21537);
not I_1126 (I21691,I2514);
DFFARX1 I_1127 (I671184,I2507,I21691,I21717,);
DFFARX1 I_1128 (I21717,I2507,I21691,I21734,);
not I_1129 (I21742,I21734);
nand I_1130 (I21759,I671199,I671202);
and I_1131 (I21776,I21759,I671181);
DFFARX1 I_1132 (I21776,I2507,I21691,I21802,);
DFFARX1 I_1133 (I21802,I2507,I21691,I21683,);
DFFARX1 I_1134 (I21802,I2507,I21691,I21674,);
DFFARX1 I_1135 (I671187,I2507,I21691,I21847,);
nand I_1136 (I21855,I21847,I671193);
not I_1137 (I21872,I21855);
nor I_1138 (I21671,I21717,I21872);
DFFARX1 I_1139 (I671181,I2507,I21691,I21912,);
not I_1140 (I21920,I21912);
nor I_1141 (I21677,I21920,I21742);
nand I_1142 (I21665,I21920,I21855);
nand I_1143 (I21965,I671196,I671178);
and I_1144 (I21982,I21965,I671190);
DFFARX1 I_1145 (I21982,I2507,I21691,I22008,);
nor I_1146 (I22016,I22008,I21717);
DFFARX1 I_1147 (I22016,I2507,I21691,I21659,);
not I_1148 (I22047,I22008);
nor I_1149 (I22064,I671178,I671178);
not I_1150 (I22081,I22064);
nor I_1151 (I22098,I21855,I22081);
nor I_1152 (I22115,I22047,I22098);
DFFARX1 I_1153 (I22115,I2507,I21691,I21680,);
nor I_1154 (I22146,I22008,I22081);
nor I_1155 (I21668,I21872,I22146);
nor I_1156 (I21662,I22008,I22064);
not I_1157 (I22218,I2514);
DFFARX1 I_1158 (I749214,I2507,I22218,I22244,);
DFFARX1 I_1159 (I22244,I2507,I22218,I22261,);
not I_1160 (I22269,I22261);
nand I_1161 (I22286,I749229,I749232);
and I_1162 (I22303,I22286,I749211);
DFFARX1 I_1163 (I22303,I2507,I22218,I22329,);
DFFARX1 I_1164 (I22329,I2507,I22218,I22210,);
DFFARX1 I_1165 (I22329,I2507,I22218,I22201,);
DFFARX1 I_1166 (I749217,I2507,I22218,I22374,);
nand I_1167 (I22382,I22374,I749223);
not I_1168 (I22399,I22382);
nor I_1169 (I22198,I22244,I22399);
DFFARX1 I_1170 (I749211,I2507,I22218,I22439,);
not I_1171 (I22447,I22439);
nor I_1172 (I22204,I22447,I22269);
nand I_1173 (I22192,I22447,I22382);
nand I_1174 (I22492,I749226,I749208);
and I_1175 (I22509,I22492,I749220);
DFFARX1 I_1176 (I22509,I2507,I22218,I22535,);
nor I_1177 (I22543,I22535,I22244);
DFFARX1 I_1178 (I22543,I2507,I22218,I22186,);
not I_1179 (I22574,I22535);
nor I_1180 (I22591,I749208,I749208);
not I_1181 (I22608,I22591);
nor I_1182 (I22625,I22382,I22608);
nor I_1183 (I22642,I22574,I22625);
DFFARX1 I_1184 (I22642,I2507,I22218,I22207,);
nor I_1185 (I22673,I22535,I22608);
nor I_1186 (I22195,I22399,I22673);
nor I_1187 (I22189,I22535,I22591);
not I_1188 (I22745,I2514);
DFFARX1 I_1189 (I1157810,I2507,I22745,I22771,);
DFFARX1 I_1190 (I22771,I2507,I22745,I22788,);
not I_1191 (I22796,I22788);
nand I_1192 (I22813,I1157798,I1157789);
and I_1193 (I22830,I22813,I1157786);
DFFARX1 I_1194 (I22830,I2507,I22745,I22856,);
DFFARX1 I_1195 (I22856,I2507,I22745,I22737,);
DFFARX1 I_1196 (I22856,I2507,I22745,I22728,);
DFFARX1 I_1197 (I1157792,I2507,I22745,I22901,);
nand I_1198 (I22909,I22901,I1157804);
not I_1199 (I22926,I22909);
nor I_1200 (I22725,I22771,I22926);
DFFARX1 I_1201 (I1157801,I2507,I22745,I22966,);
not I_1202 (I22974,I22966);
nor I_1203 (I22731,I22974,I22796);
nand I_1204 (I22719,I22974,I22909);
nand I_1205 (I23019,I1157795,I1157789);
and I_1206 (I23036,I23019,I1157807);
DFFARX1 I_1207 (I23036,I2507,I22745,I23062,);
nor I_1208 (I23070,I23062,I22771);
DFFARX1 I_1209 (I23070,I2507,I22745,I22713,);
not I_1210 (I23101,I23062);
nor I_1211 (I23118,I1157786,I1157789);
not I_1212 (I23135,I23118);
nor I_1213 (I23152,I22909,I23135);
nor I_1214 (I23169,I23101,I23152);
DFFARX1 I_1215 (I23169,I2507,I22745,I22734,);
nor I_1216 (I23200,I23062,I23135);
nor I_1217 (I22722,I22926,I23200);
nor I_1218 (I22716,I23062,I23118);
not I_1219 (I23272,I2514);
DFFARX1 I_1220 (I771178,I2507,I23272,I23298,);
DFFARX1 I_1221 (I23298,I2507,I23272,I23315,);
not I_1222 (I23323,I23315);
nand I_1223 (I23340,I771193,I771196);
and I_1224 (I23357,I23340,I771175);
DFFARX1 I_1225 (I23357,I2507,I23272,I23383,);
DFFARX1 I_1226 (I23383,I2507,I23272,I23264,);
DFFARX1 I_1227 (I23383,I2507,I23272,I23255,);
DFFARX1 I_1228 (I771181,I2507,I23272,I23428,);
nand I_1229 (I23436,I23428,I771187);
not I_1230 (I23453,I23436);
nor I_1231 (I23252,I23298,I23453);
DFFARX1 I_1232 (I771175,I2507,I23272,I23493,);
not I_1233 (I23501,I23493);
nor I_1234 (I23258,I23501,I23323);
nand I_1235 (I23246,I23501,I23436);
nand I_1236 (I23546,I771190,I771172);
and I_1237 (I23563,I23546,I771184);
DFFARX1 I_1238 (I23563,I2507,I23272,I23589,);
nor I_1239 (I23597,I23589,I23298);
DFFARX1 I_1240 (I23597,I2507,I23272,I23240,);
not I_1241 (I23628,I23589);
nor I_1242 (I23645,I771172,I771172);
not I_1243 (I23662,I23645);
nor I_1244 (I23679,I23436,I23662);
nor I_1245 (I23696,I23628,I23679);
DFFARX1 I_1246 (I23696,I2507,I23272,I23261,);
nor I_1247 (I23727,I23589,I23662);
nor I_1248 (I23249,I23453,I23727);
nor I_1249 (I23243,I23589,I23645);
not I_1250 (I23799,I2514);
DFFARX1 I_1251 (I444143,I2507,I23799,I23825,);
DFFARX1 I_1252 (I23825,I2507,I23799,I23842,);
not I_1253 (I23850,I23842);
nand I_1254 (I23867,I444143,I444146);
and I_1255 (I23884,I23867,I444167);
DFFARX1 I_1256 (I23884,I2507,I23799,I23910,);
DFFARX1 I_1257 (I23910,I2507,I23799,I23791,);
DFFARX1 I_1258 (I23910,I2507,I23799,I23782,);
DFFARX1 I_1259 (I444155,I2507,I23799,I23955,);
nand I_1260 (I23963,I23955,I444158);
not I_1261 (I23980,I23963);
nor I_1262 (I23779,I23825,I23980);
DFFARX1 I_1263 (I444164,I2507,I23799,I24020,);
not I_1264 (I24028,I24020);
nor I_1265 (I23785,I24028,I23850);
nand I_1266 (I23773,I24028,I23963);
nand I_1267 (I24073,I444161,I444149);
and I_1268 (I24090,I24073,I444152);
DFFARX1 I_1269 (I24090,I2507,I23799,I24116,);
nor I_1270 (I24124,I24116,I23825);
DFFARX1 I_1271 (I24124,I2507,I23799,I23767,);
not I_1272 (I24155,I24116);
nor I_1273 (I24172,I444170,I444149);
not I_1274 (I24189,I24172);
nor I_1275 (I24206,I23963,I24189);
nor I_1276 (I24223,I24155,I24206);
DFFARX1 I_1277 (I24223,I2507,I23799,I23788,);
nor I_1278 (I24254,I24116,I24189);
nor I_1279 (I23776,I23980,I24254);
nor I_1280 (I23770,I24116,I24172);
not I_1281 (I24326,I2514);
DFFARX1 I_1282 (I610503,I2507,I24326,I24352,);
DFFARX1 I_1283 (I24352,I2507,I24326,I24369,);
not I_1284 (I24377,I24369);
nand I_1285 (I24394,I610488,I610506);
and I_1286 (I24411,I24394,I610500);
DFFARX1 I_1287 (I24411,I2507,I24326,I24437,);
DFFARX1 I_1288 (I24437,I2507,I24326,I24318,);
DFFARX1 I_1289 (I24437,I2507,I24326,I24309,);
DFFARX1 I_1290 (I610497,I2507,I24326,I24482,);
nand I_1291 (I24490,I24482,I610488);
not I_1292 (I24507,I24490);
nor I_1293 (I24306,I24352,I24507);
DFFARX1 I_1294 (I610491,I2507,I24326,I24547,);
not I_1295 (I24555,I24547);
nor I_1296 (I24312,I24555,I24377);
nand I_1297 (I24300,I24555,I24490);
nand I_1298 (I24600,I610512,I610494);
and I_1299 (I24617,I24600,I610509);
DFFARX1 I_1300 (I24617,I2507,I24326,I24643,);
nor I_1301 (I24651,I24643,I24352);
DFFARX1 I_1302 (I24651,I2507,I24326,I24294,);
not I_1303 (I24682,I24643);
nor I_1304 (I24699,I610491,I610494);
not I_1305 (I24716,I24699);
nor I_1306 (I24733,I24490,I24716);
nor I_1307 (I24750,I24682,I24733);
DFFARX1 I_1308 (I24750,I2507,I24326,I24315,);
nor I_1309 (I24781,I24643,I24716);
nor I_1310 (I24303,I24507,I24781);
nor I_1311 (I24297,I24643,I24699);
not I_1312 (I24853,I2514);
DFFARX1 I_1313 (I1109836,I2507,I24853,I24879,);
DFFARX1 I_1314 (I24879,I2507,I24853,I24896,);
not I_1315 (I24904,I24896);
nand I_1316 (I24921,I1109824,I1109815);
and I_1317 (I24938,I24921,I1109812);
DFFARX1 I_1318 (I24938,I2507,I24853,I24964,);
DFFARX1 I_1319 (I24964,I2507,I24853,I24845,);
DFFARX1 I_1320 (I24964,I2507,I24853,I24836,);
DFFARX1 I_1321 (I1109818,I2507,I24853,I25009,);
nand I_1322 (I25017,I25009,I1109830);
not I_1323 (I25034,I25017);
nor I_1324 (I24833,I24879,I25034);
DFFARX1 I_1325 (I1109827,I2507,I24853,I25074,);
not I_1326 (I25082,I25074);
nor I_1327 (I24839,I25082,I24904);
nand I_1328 (I24827,I25082,I25017);
nand I_1329 (I25127,I1109821,I1109815);
and I_1330 (I25144,I25127,I1109833);
DFFARX1 I_1331 (I25144,I2507,I24853,I25170,);
nor I_1332 (I25178,I25170,I24879);
DFFARX1 I_1333 (I25178,I2507,I24853,I24821,);
not I_1334 (I25209,I25170);
nor I_1335 (I25226,I1109812,I1109815);
not I_1336 (I25243,I25226);
nor I_1337 (I25260,I25017,I25243);
nor I_1338 (I25277,I25209,I25260);
DFFARX1 I_1339 (I25277,I2507,I24853,I24842,);
nor I_1340 (I25308,I25170,I25243);
nor I_1341 (I24830,I25034,I25308);
nor I_1342 (I24824,I25170,I25226);
not I_1343 (I25380,I2514);
DFFARX1 I_1344 (I113360,I2507,I25380,I25406,);
DFFARX1 I_1345 (I25406,I2507,I25380,I25423,);
not I_1346 (I25431,I25423);
nand I_1347 (I25448,I113360,I113375);
and I_1348 (I25465,I25448,I113378);
DFFARX1 I_1349 (I25465,I2507,I25380,I25491,);
DFFARX1 I_1350 (I25491,I2507,I25380,I25372,);
DFFARX1 I_1351 (I25491,I2507,I25380,I25363,);
DFFARX1 I_1352 (I113372,I2507,I25380,I25536,);
nand I_1353 (I25544,I25536,I113381);
not I_1354 (I25561,I25544);
nor I_1355 (I25360,I25406,I25561);
DFFARX1 I_1356 (I113357,I2507,I25380,I25601,);
not I_1357 (I25609,I25601);
nor I_1358 (I25366,I25609,I25431);
nand I_1359 (I25354,I25609,I25544);
nand I_1360 (I25654,I113357,I113363);
and I_1361 (I25671,I25654,I113366);
DFFARX1 I_1362 (I25671,I2507,I25380,I25697,);
nor I_1363 (I25705,I25697,I25406);
DFFARX1 I_1364 (I25705,I2507,I25380,I25348,);
not I_1365 (I25736,I25697);
nor I_1366 (I25753,I113369,I113363);
not I_1367 (I25770,I25753);
nor I_1368 (I25787,I25544,I25770);
nor I_1369 (I25804,I25736,I25787);
DFFARX1 I_1370 (I25804,I2507,I25380,I25369,);
nor I_1371 (I25835,I25697,I25770);
nor I_1372 (I25357,I25561,I25835);
nor I_1373 (I25351,I25697,I25753);
not I_1374 (I25907,I2514);
DFFARX1 I_1375 (I972867,I2507,I25907,I25933,);
DFFARX1 I_1376 (I25933,I2507,I25907,I25950,);
not I_1377 (I25958,I25950);
nand I_1378 (I25975,I972843,I972870);
and I_1379 (I25992,I25975,I972855);
DFFARX1 I_1380 (I25992,I2507,I25907,I26018,);
DFFARX1 I_1381 (I26018,I2507,I25907,I25899,);
DFFARX1 I_1382 (I26018,I2507,I25907,I25890,);
DFFARX1 I_1383 (I972861,I2507,I25907,I26063,);
nand I_1384 (I26071,I26063,I972846);
not I_1385 (I26088,I26071);
nor I_1386 (I25887,I25933,I26088);
DFFARX1 I_1387 (I972864,I2507,I25907,I26128,);
not I_1388 (I26136,I26128);
nor I_1389 (I25893,I26136,I25958);
nand I_1390 (I25881,I26136,I26071);
nand I_1391 (I26181,I972849,I972852);
and I_1392 (I26198,I26181,I972843);
DFFARX1 I_1393 (I26198,I2507,I25907,I26224,);
nor I_1394 (I26232,I26224,I25933);
DFFARX1 I_1395 (I26232,I2507,I25907,I25875,);
not I_1396 (I26263,I26224);
nor I_1397 (I26280,I972858,I972852);
not I_1398 (I26297,I26280);
nor I_1399 (I26314,I26071,I26297);
nor I_1400 (I26331,I26263,I26314);
DFFARX1 I_1401 (I26331,I2507,I25907,I25896,);
nor I_1402 (I26362,I26224,I26297);
nor I_1403 (I25884,I26088,I26362);
nor I_1404 (I25878,I26224,I26280);
not I_1405 (I26434,I2514);
DFFARX1 I_1406 (I143105,I2507,I26434,I26460,);
DFFARX1 I_1407 (I26460,I2507,I26434,I26477,);
not I_1408 (I26485,I26477);
nand I_1409 (I26502,I143108,I143090);
and I_1410 (I26519,I26502,I143096);
DFFARX1 I_1411 (I26519,I2507,I26434,I26545,);
DFFARX1 I_1412 (I26545,I2507,I26434,I26426,);
DFFARX1 I_1413 (I26545,I2507,I26434,I26417,);
DFFARX1 I_1414 (I143099,I2507,I26434,I26590,);
nand I_1415 (I26598,I26590,I143090);
not I_1416 (I26615,I26598);
nor I_1417 (I26414,I26460,I26615);
DFFARX1 I_1418 (I143111,I2507,I26434,I26655,);
not I_1419 (I26663,I26655);
nor I_1420 (I26420,I26663,I26485);
nand I_1421 (I26408,I26663,I26598);
nand I_1422 (I26708,I143114,I143102);
and I_1423 (I26725,I26708,I143093);
DFFARX1 I_1424 (I26725,I2507,I26434,I26751,);
nor I_1425 (I26759,I26751,I26460);
DFFARX1 I_1426 (I26759,I2507,I26434,I26402,);
not I_1427 (I26790,I26751);
nor I_1428 (I26807,I143117,I143102);
not I_1429 (I26824,I26807);
nor I_1430 (I26841,I26598,I26824);
nor I_1431 (I26858,I26790,I26841);
DFFARX1 I_1432 (I26858,I2507,I26434,I26423,);
nor I_1433 (I26889,I26751,I26824);
nor I_1434 (I26411,I26615,I26889);
nor I_1435 (I26405,I26751,I26807);
not I_1436 (I26961,I2514);
DFFARX1 I_1437 (I728984,I2507,I26961,I26987,);
DFFARX1 I_1438 (I26987,I2507,I26961,I27004,);
not I_1439 (I27012,I27004);
nand I_1440 (I27029,I728999,I729002);
and I_1441 (I27046,I27029,I728981);
DFFARX1 I_1442 (I27046,I2507,I26961,I27072,);
DFFARX1 I_1443 (I27072,I2507,I26961,I26953,);
DFFARX1 I_1444 (I27072,I2507,I26961,I26944,);
DFFARX1 I_1445 (I728987,I2507,I26961,I27117,);
nand I_1446 (I27125,I27117,I728993);
not I_1447 (I27142,I27125);
nor I_1448 (I26941,I26987,I27142);
DFFARX1 I_1449 (I728981,I2507,I26961,I27182,);
not I_1450 (I27190,I27182);
nor I_1451 (I26947,I27190,I27012);
nand I_1452 (I26935,I27190,I27125);
nand I_1453 (I27235,I728996,I728978);
and I_1454 (I27252,I27235,I728990);
DFFARX1 I_1455 (I27252,I2507,I26961,I27278,);
nor I_1456 (I27286,I27278,I26987);
DFFARX1 I_1457 (I27286,I2507,I26961,I26929,);
not I_1458 (I27317,I27278);
nor I_1459 (I27334,I728978,I728978);
not I_1460 (I27351,I27334);
nor I_1461 (I27368,I27125,I27351);
nor I_1462 (I27385,I27317,I27368);
DFFARX1 I_1463 (I27385,I2507,I26961,I26950,);
nor I_1464 (I27416,I27278,I27351);
nor I_1465 (I26938,I27142,I27416);
nor I_1466 (I26932,I27278,I27334);
not I_1467 (I27488,I2514);
DFFARX1 I_1468 (I336645,I2507,I27488,I27514,);
DFFARX1 I_1469 (I27514,I2507,I27488,I27531,);
not I_1470 (I27539,I27531);
nand I_1471 (I27556,I336642,I336636);
and I_1472 (I27573,I27556,I336630);
DFFARX1 I_1473 (I27573,I2507,I27488,I27599,);
DFFARX1 I_1474 (I27599,I2507,I27488,I27480,);
DFFARX1 I_1475 (I27599,I2507,I27488,I27471,);
DFFARX1 I_1476 (I336618,I2507,I27488,I27644,);
nand I_1477 (I27652,I27644,I336627);
not I_1478 (I27669,I27652);
nor I_1479 (I27468,I27514,I27669);
DFFARX1 I_1480 (I336624,I2507,I27488,I27709,);
not I_1481 (I27717,I27709);
nor I_1482 (I27474,I27717,I27539);
nand I_1483 (I27462,I27717,I27652);
nand I_1484 (I27762,I336621,I336639);
and I_1485 (I27779,I27762,I336618);
DFFARX1 I_1486 (I27779,I2507,I27488,I27805,);
nor I_1487 (I27813,I27805,I27514);
DFFARX1 I_1488 (I27813,I2507,I27488,I27456,);
not I_1489 (I27844,I27805);
nor I_1490 (I27861,I336633,I336639);
not I_1491 (I27878,I27861);
nor I_1492 (I27895,I27652,I27878);
nor I_1493 (I27912,I27844,I27895);
DFFARX1 I_1494 (I27912,I2507,I27488,I27477,);
nor I_1495 (I27943,I27805,I27878);
nor I_1496 (I27465,I27669,I27943);
nor I_1497 (I27459,I27805,I27861);
not I_1498 (I28015,I2514);
DFFARX1 I_1499 (I557327,I2507,I28015,I28041,);
DFFARX1 I_1500 (I28041,I2507,I28015,I28058,);
not I_1501 (I28066,I28058);
nand I_1502 (I28083,I557312,I557330);
and I_1503 (I28100,I28083,I557324);
DFFARX1 I_1504 (I28100,I2507,I28015,I28126,);
DFFARX1 I_1505 (I28126,I2507,I28015,I28007,);
DFFARX1 I_1506 (I28126,I2507,I28015,I27998,);
DFFARX1 I_1507 (I557321,I2507,I28015,I28171,);
nand I_1508 (I28179,I28171,I557312);
not I_1509 (I28196,I28179);
nor I_1510 (I27995,I28041,I28196);
DFFARX1 I_1511 (I557315,I2507,I28015,I28236,);
not I_1512 (I28244,I28236);
nor I_1513 (I28001,I28244,I28066);
nand I_1514 (I27989,I28244,I28179);
nand I_1515 (I28289,I557336,I557318);
and I_1516 (I28306,I28289,I557333);
DFFARX1 I_1517 (I28306,I2507,I28015,I28332,);
nor I_1518 (I28340,I28332,I28041);
DFFARX1 I_1519 (I28340,I2507,I28015,I27983,);
not I_1520 (I28371,I28332);
nor I_1521 (I28388,I557315,I557318);
not I_1522 (I28405,I28388);
nor I_1523 (I28422,I28179,I28405);
nor I_1524 (I28439,I28371,I28422);
DFFARX1 I_1525 (I28439,I2507,I28015,I28004,);
nor I_1526 (I28470,I28332,I28405);
nor I_1527 (I27992,I28196,I28470);
nor I_1528 (I27986,I28332,I28388);
not I_1529 (I28542,I2514);
DFFARX1 I_1530 (I1024172,I2507,I28542,I28568,);
DFFARX1 I_1531 (I28568,I2507,I28542,I28585,);
not I_1532 (I28593,I28585);
nand I_1533 (I28610,I1024166,I1024187);
and I_1534 (I28627,I28610,I1024172);
DFFARX1 I_1535 (I28627,I2507,I28542,I28653,);
DFFARX1 I_1536 (I28653,I2507,I28542,I28534,);
DFFARX1 I_1537 (I28653,I2507,I28542,I28525,);
DFFARX1 I_1538 (I1024169,I2507,I28542,I28698,);
nand I_1539 (I28706,I28698,I1024178);
not I_1540 (I28723,I28706);
nor I_1541 (I28522,I28568,I28723);
DFFARX1 I_1542 (I1024166,I2507,I28542,I28763,);
not I_1543 (I28771,I28763);
nor I_1544 (I28528,I28771,I28593);
nand I_1545 (I28516,I28771,I28706);
nand I_1546 (I28816,I1024169,I1024184);
and I_1547 (I28833,I28816,I1024175);
DFFARX1 I_1548 (I28833,I2507,I28542,I28859,);
nor I_1549 (I28867,I28859,I28568);
DFFARX1 I_1550 (I28867,I2507,I28542,I28510,);
not I_1551 (I28898,I28859);
nor I_1552 (I28915,I1024181,I1024184);
not I_1553 (I28932,I28915);
nor I_1554 (I28949,I28706,I28932);
nor I_1555 (I28966,I28898,I28949);
DFFARX1 I_1556 (I28966,I2507,I28542,I28531,);
nor I_1557 (I28997,I28859,I28932);
nor I_1558 (I28519,I28723,I28997);
nor I_1559 (I28513,I28859,I28915);
not I_1560 (I29069,I2514);
DFFARX1 I_1561 (I804892,I2507,I29069,I29095,);
DFFARX1 I_1562 (I29095,I2507,I29069,I29112,);
not I_1563 (I29120,I29112);
nand I_1564 (I29137,I804883,I804904);
and I_1565 (I29154,I29137,I804886);
DFFARX1 I_1566 (I29154,I2507,I29069,I29180,);
DFFARX1 I_1567 (I29180,I2507,I29069,I29061,);
DFFARX1 I_1568 (I29180,I2507,I29069,I29052,);
DFFARX1 I_1569 (I804886,I2507,I29069,I29225,);
nand I_1570 (I29233,I29225,I804901);
not I_1571 (I29250,I29233);
nor I_1572 (I29049,I29095,I29250);
DFFARX1 I_1573 (I804895,I2507,I29069,I29290,);
not I_1574 (I29298,I29290);
nor I_1575 (I29055,I29298,I29120);
nand I_1576 (I29043,I29298,I29233);
nand I_1577 (I29343,I804889,I804898);
and I_1578 (I29360,I29343,I804883);
DFFARX1 I_1579 (I29360,I2507,I29069,I29386,);
nor I_1580 (I29394,I29386,I29095);
DFFARX1 I_1581 (I29394,I2507,I29069,I29037,);
not I_1582 (I29425,I29386);
nor I_1583 (I29442,I804889,I804898);
not I_1584 (I29459,I29442);
nor I_1585 (I29476,I29233,I29459);
nor I_1586 (I29493,I29425,I29476);
DFFARX1 I_1587 (I29493,I2507,I29069,I29058,);
nor I_1588 (I29524,I29386,I29459);
nor I_1589 (I29046,I29250,I29524);
nor I_1590 (I29040,I29386,I29442);
not I_1591 (I29596,I2514);
DFFARX1 I_1592 (I1119662,I2507,I29596,I29622,);
DFFARX1 I_1593 (I29622,I2507,I29596,I29639,);
not I_1594 (I29647,I29639);
nand I_1595 (I29664,I1119650,I1119641);
and I_1596 (I29681,I29664,I1119638);
DFFARX1 I_1597 (I29681,I2507,I29596,I29707,);
DFFARX1 I_1598 (I29707,I2507,I29596,I29588,);
DFFARX1 I_1599 (I29707,I2507,I29596,I29579,);
DFFARX1 I_1600 (I1119644,I2507,I29596,I29752,);
nand I_1601 (I29760,I29752,I1119656);
not I_1602 (I29777,I29760);
nor I_1603 (I29576,I29622,I29777);
DFFARX1 I_1604 (I1119653,I2507,I29596,I29817,);
not I_1605 (I29825,I29817);
nor I_1606 (I29582,I29825,I29647);
nand I_1607 (I29570,I29825,I29760);
nand I_1608 (I29870,I1119647,I1119641);
and I_1609 (I29887,I29870,I1119659);
DFFARX1 I_1610 (I29887,I2507,I29596,I29913,);
nor I_1611 (I29921,I29913,I29622);
DFFARX1 I_1612 (I29921,I2507,I29596,I29564,);
not I_1613 (I29952,I29913);
nor I_1614 (I29969,I1119638,I1119641);
not I_1615 (I29986,I29969);
nor I_1616 (I30003,I29760,I29986);
nor I_1617 (I30020,I29952,I30003);
DFFARX1 I_1618 (I30020,I2507,I29596,I29585,);
nor I_1619 (I30051,I29913,I29986);
nor I_1620 (I29573,I29777,I30051);
nor I_1621 (I29567,I29913,I29969);
not I_1622 (I30123,I2514);
DFFARX1 I_1623 (I724938,I2507,I30123,I30149,);
DFFARX1 I_1624 (I30149,I2507,I30123,I30166,);
not I_1625 (I30174,I30166);
nand I_1626 (I30191,I724953,I724956);
and I_1627 (I30208,I30191,I724935);
DFFARX1 I_1628 (I30208,I2507,I30123,I30234,);
DFFARX1 I_1629 (I30234,I2507,I30123,I30115,);
DFFARX1 I_1630 (I30234,I2507,I30123,I30106,);
DFFARX1 I_1631 (I724941,I2507,I30123,I30279,);
nand I_1632 (I30287,I30279,I724947);
not I_1633 (I30304,I30287);
nor I_1634 (I30103,I30149,I30304);
DFFARX1 I_1635 (I724935,I2507,I30123,I30344,);
not I_1636 (I30352,I30344);
nor I_1637 (I30109,I30352,I30174);
nand I_1638 (I30097,I30352,I30287);
nand I_1639 (I30397,I724950,I724932);
and I_1640 (I30414,I30397,I724944);
DFFARX1 I_1641 (I30414,I2507,I30123,I30440,);
nor I_1642 (I30448,I30440,I30149);
DFFARX1 I_1643 (I30448,I2507,I30123,I30091,);
not I_1644 (I30479,I30440);
nor I_1645 (I30496,I724932,I724932);
not I_1646 (I30513,I30496);
nor I_1647 (I30530,I30287,I30513);
nor I_1648 (I30547,I30479,I30530);
DFFARX1 I_1649 (I30547,I2507,I30123,I30112,);
nor I_1650 (I30578,I30440,I30513);
nor I_1651 (I30100,I30304,I30578);
nor I_1652 (I30094,I30440,I30496);
not I_1653 (I30650,I2514);
DFFARX1 I_1654 (I395183,I2507,I30650,I30676,);
DFFARX1 I_1655 (I30676,I2507,I30650,I30693,);
not I_1656 (I30701,I30693);
nand I_1657 (I30718,I395183,I395186);
and I_1658 (I30735,I30718,I395207);
DFFARX1 I_1659 (I30735,I2507,I30650,I30761,);
DFFARX1 I_1660 (I30761,I2507,I30650,I30642,);
DFFARX1 I_1661 (I30761,I2507,I30650,I30633,);
DFFARX1 I_1662 (I395195,I2507,I30650,I30806,);
nand I_1663 (I30814,I30806,I395198);
not I_1664 (I30831,I30814);
nor I_1665 (I30630,I30676,I30831);
DFFARX1 I_1666 (I395204,I2507,I30650,I30871,);
not I_1667 (I30879,I30871);
nor I_1668 (I30636,I30879,I30701);
nand I_1669 (I30624,I30879,I30814);
nand I_1670 (I30924,I395201,I395189);
and I_1671 (I30941,I30924,I395192);
DFFARX1 I_1672 (I30941,I2507,I30650,I30967,);
nor I_1673 (I30975,I30967,I30676);
DFFARX1 I_1674 (I30975,I2507,I30650,I30618,);
not I_1675 (I31006,I30967);
nor I_1676 (I31023,I395210,I395189);
not I_1677 (I31040,I31023);
nor I_1678 (I31057,I30814,I31040);
nor I_1679 (I31074,I31006,I31057);
DFFARX1 I_1680 (I31074,I2507,I30650,I30639,);
nor I_1681 (I31105,I30967,I31040);
nor I_1682 (I30627,I30831,I31105);
nor I_1683 (I30621,I30967,I31023);
not I_1684 (I31177,I2514);
DFFARX1 I_1685 (I561951,I2507,I31177,I31203,);
DFFARX1 I_1686 (I31203,I2507,I31177,I31220,);
not I_1687 (I31228,I31220);
nand I_1688 (I31245,I561936,I561954);
and I_1689 (I31262,I31245,I561948);
DFFARX1 I_1690 (I31262,I2507,I31177,I31288,);
DFFARX1 I_1691 (I31288,I2507,I31177,I31169,);
DFFARX1 I_1692 (I31288,I2507,I31177,I31160,);
DFFARX1 I_1693 (I561945,I2507,I31177,I31333,);
nand I_1694 (I31341,I31333,I561936);
not I_1695 (I31358,I31341);
nor I_1696 (I31157,I31203,I31358);
DFFARX1 I_1697 (I561939,I2507,I31177,I31398,);
not I_1698 (I31406,I31398);
nor I_1699 (I31163,I31406,I31228);
nand I_1700 (I31151,I31406,I31341);
nand I_1701 (I31451,I561960,I561942);
and I_1702 (I31468,I31451,I561957);
DFFARX1 I_1703 (I31468,I2507,I31177,I31494,);
nor I_1704 (I31502,I31494,I31203);
DFFARX1 I_1705 (I31502,I2507,I31177,I31145,);
not I_1706 (I31533,I31494);
nor I_1707 (I31550,I561939,I561942);
not I_1708 (I31567,I31550);
nor I_1709 (I31584,I31341,I31567);
nor I_1710 (I31601,I31533,I31584);
DFFARX1 I_1711 (I31601,I2507,I31177,I31166,);
nor I_1712 (I31632,I31494,I31567);
nor I_1713 (I31154,I31358,I31632);
nor I_1714 (I31148,I31494,I31550);
not I_1715 (I31704,I2514);
DFFARX1 I_1716 (I1132378,I2507,I31704,I31730,);
DFFARX1 I_1717 (I31730,I2507,I31704,I31747,);
not I_1718 (I31755,I31747);
nand I_1719 (I31772,I1132366,I1132357);
and I_1720 (I31789,I31772,I1132354);
DFFARX1 I_1721 (I31789,I2507,I31704,I31815,);
DFFARX1 I_1722 (I31815,I2507,I31704,I31696,);
DFFARX1 I_1723 (I31815,I2507,I31704,I31687,);
DFFARX1 I_1724 (I1132360,I2507,I31704,I31860,);
nand I_1725 (I31868,I31860,I1132372);
not I_1726 (I31885,I31868);
nor I_1727 (I31684,I31730,I31885);
DFFARX1 I_1728 (I1132369,I2507,I31704,I31925,);
not I_1729 (I31933,I31925);
nor I_1730 (I31690,I31933,I31755);
nand I_1731 (I31678,I31933,I31868);
nand I_1732 (I31978,I1132363,I1132357);
and I_1733 (I31995,I31978,I1132375);
DFFARX1 I_1734 (I31995,I2507,I31704,I32021,);
nor I_1735 (I32029,I32021,I31730);
DFFARX1 I_1736 (I32029,I2507,I31704,I31672,);
not I_1737 (I32060,I32021);
nor I_1738 (I32077,I1132354,I1132357);
not I_1739 (I32094,I32077);
nor I_1740 (I32111,I31868,I32094);
nor I_1741 (I32128,I32060,I32111);
DFFARX1 I_1742 (I32128,I2507,I31704,I31693,);
nor I_1743 (I32159,I32021,I32094);
nor I_1744 (I31681,I31885,I32159);
nor I_1745 (I31675,I32021,I32077);
not I_1746 (I32231,I2514);
DFFARX1 I_1747 (I725516,I2507,I32231,I32257,);
DFFARX1 I_1748 (I32257,I2507,I32231,I32274,);
not I_1749 (I32282,I32274);
nand I_1750 (I32299,I725531,I725534);
and I_1751 (I32316,I32299,I725513);
DFFARX1 I_1752 (I32316,I2507,I32231,I32342,);
DFFARX1 I_1753 (I32342,I2507,I32231,I32223,);
DFFARX1 I_1754 (I32342,I2507,I32231,I32214,);
DFFARX1 I_1755 (I725519,I2507,I32231,I32387,);
nand I_1756 (I32395,I32387,I725525);
not I_1757 (I32412,I32395);
nor I_1758 (I32211,I32257,I32412);
DFFARX1 I_1759 (I725513,I2507,I32231,I32452,);
not I_1760 (I32460,I32452);
nor I_1761 (I32217,I32460,I32282);
nand I_1762 (I32205,I32460,I32395);
nand I_1763 (I32505,I725528,I725510);
and I_1764 (I32522,I32505,I725522);
DFFARX1 I_1765 (I32522,I2507,I32231,I32548,);
nor I_1766 (I32556,I32548,I32257);
DFFARX1 I_1767 (I32556,I2507,I32231,I32199,);
not I_1768 (I32587,I32548);
nor I_1769 (I32604,I725510,I725510);
not I_1770 (I32621,I32604);
nor I_1771 (I32638,I32395,I32621);
nor I_1772 (I32655,I32587,I32638);
DFFARX1 I_1773 (I32655,I2507,I32231,I32220,);
nor I_1774 (I32686,I32548,I32621);
nor I_1775 (I32208,I32412,I32686);
nor I_1776 (I32202,I32548,I32604);
not I_1777 (I32758,I2514);
DFFARX1 I_1778 (I302390,I2507,I32758,I32784,);
DFFARX1 I_1779 (I32784,I2507,I32758,I32801,);
not I_1780 (I32809,I32801);
nand I_1781 (I32826,I302387,I302381);
and I_1782 (I32843,I32826,I302375);
DFFARX1 I_1783 (I32843,I2507,I32758,I32869,);
DFFARX1 I_1784 (I32869,I2507,I32758,I32750,);
DFFARX1 I_1785 (I32869,I2507,I32758,I32741,);
DFFARX1 I_1786 (I302363,I2507,I32758,I32914,);
nand I_1787 (I32922,I32914,I302372);
not I_1788 (I32939,I32922);
nor I_1789 (I32738,I32784,I32939);
DFFARX1 I_1790 (I302369,I2507,I32758,I32979,);
not I_1791 (I32987,I32979);
nor I_1792 (I32744,I32987,I32809);
nand I_1793 (I32732,I32987,I32922);
nand I_1794 (I33032,I302366,I302384);
and I_1795 (I33049,I33032,I302363);
DFFARX1 I_1796 (I33049,I2507,I32758,I33075,);
nor I_1797 (I33083,I33075,I32784);
DFFARX1 I_1798 (I33083,I2507,I32758,I32726,);
not I_1799 (I33114,I33075);
nor I_1800 (I33131,I302378,I302384);
not I_1801 (I33148,I33131);
nor I_1802 (I33165,I32922,I33148);
nor I_1803 (I33182,I33114,I33165);
DFFARX1 I_1804 (I33182,I2507,I32758,I32747,);
nor I_1805 (I33213,I33075,I33148);
nor I_1806 (I32735,I32939,I33213);
nor I_1807 (I32729,I33075,I33131);
not I_1808 (I33285,I2514);
DFFARX1 I_1809 (I315565,I2507,I33285,I33311,);
DFFARX1 I_1810 (I33311,I2507,I33285,I33328,);
not I_1811 (I33336,I33328);
nand I_1812 (I33353,I315562,I315556);
and I_1813 (I33370,I33353,I315550);
DFFARX1 I_1814 (I33370,I2507,I33285,I33396,);
DFFARX1 I_1815 (I33396,I2507,I33285,I33277,);
DFFARX1 I_1816 (I33396,I2507,I33285,I33268,);
DFFARX1 I_1817 (I315538,I2507,I33285,I33441,);
nand I_1818 (I33449,I33441,I315547);
not I_1819 (I33466,I33449);
nor I_1820 (I33265,I33311,I33466);
DFFARX1 I_1821 (I315544,I2507,I33285,I33506,);
not I_1822 (I33514,I33506);
nor I_1823 (I33271,I33514,I33336);
nand I_1824 (I33259,I33514,I33449);
nand I_1825 (I33559,I315541,I315559);
and I_1826 (I33576,I33559,I315538);
DFFARX1 I_1827 (I33576,I2507,I33285,I33602,);
nor I_1828 (I33610,I33602,I33311);
DFFARX1 I_1829 (I33610,I2507,I33285,I33253,);
not I_1830 (I33641,I33602);
nor I_1831 (I33658,I315553,I315559);
not I_1832 (I33675,I33658);
nor I_1833 (I33692,I33449,I33675);
nor I_1834 (I33709,I33641,I33692);
DFFARX1 I_1835 (I33709,I2507,I33285,I33274,);
nor I_1836 (I33740,I33602,I33675);
nor I_1837 (I33262,I33466,I33740);
nor I_1838 (I33256,I33602,I33658);
not I_1839 (I33812,I2514);
DFFARX1 I_1840 (I1280779,I2507,I33812,I33838,);
DFFARX1 I_1841 (I33838,I2507,I33812,I33855,);
not I_1842 (I33863,I33855);
nand I_1843 (I33880,I1280782,I1280776);
and I_1844 (I33897,I33880,I1280785);
DFFARX1 I_1845 (I33897,I2507,I33812,I33923,);
DFFARX1 I_1846 (I33923,I2507,I33812,I33804,);
DFFARX1 I_1847 (I33923,I2507,I33812,I33795,);
DFFARX1 I_1848 (I1280773,I2507,I33812,I33968,);
nand I_1849 (I33976,I33968,I1280788);
not I_1850 (I33993,I33976);
nor I_1851 (I33792,I33838,I33993);
DFFARX1 I_1852 (I1280764,I2507,I33812,I34033,);
not I_1853 (I34041,I34033);
nor I_1854 (I33798,I34041,I33863);
nand I_1855 (I33786,I34041,I33976);
nand I_1856 (I34086,I1280767,I1280767);
and I_1857 (I34103,I34086,I1280764);
DFFARX1 I_1858 (I34103,I2507,I33812,I34129,);
nor I_1859 (I34137,I34129,I33838);
DFFARX1 I_1860 (I34137,I2507,I33812,I33780,);
not I_1861 (I34168,I34129);
nor I_1862 (I34185,I1280770,I1280767);
not I_1863 (I34202,I34185);
nor I_1864 (I34219,I33976,I34202);
nor I_1865 (I34236,I34168,I34219);
DFFARX1 I_1866 (I34236,I2507,I33812,I33801,);
nor I_1867 (I34267,I34129,I34202);
nor I_1868 (I33789,I33993,I34267);
nor I_1869 (I33783,I34129,I34185);
not I_1870 (I34339,I2514);
DFFARX1 I_1871 (I1264595,I2507,I34339,I34365,);
DFFARX1 I_1872 (I34365,I2507,I34339,I34382,);
not I_1873 (I34390,I34382);
nand I_1874 (I34407,I1264598,I1264592);
and I_1875 (I34424,I34407,I1264601);
DFFARX1 I_1876 (I34424,I2507,I34339,I34450,);
DFFARX1 I_1877 (I34450,I2507,I34339,I34331,);
DFFARX1 I_1878 (I34450,I2507,I34339,I34322,);
DFFARX1 I_1879 (I1264589,I2507,I34339,I34495,);
nand I_1880 (I34503,I34495,I1264604);
not I_1881 (I34520,I34503);
nor I_1882 (I34319,I34365,I34520);
DFFARX1 I_1883 (I1264580,I2507,I34339,I34560,);
not I_1884 (I34568,I34560);
nor I_1885 (I34325,I34568,I34390);
nand I_1886 (I34313,I34568,I34503);
nand I_1887 (I34613,I1264583,I1264583);
and I_1888 (I34630,I34613,I1264580);
DFFARX1 I_1889 (I34630,I2507,I34339,I34656,);
nor I_1890 (I34664,I34656,I34365);
DFFARX1 I_1891 (I34664,I2507,I34339,I34307,);
not I_1892 (I34695,I34656);
nor I_1893 (I34712,I1264586,I1264583);
not I_1894 (I34729,I34712);
nor I_1895 (I34746,I34503,I34729);
nor I_1896 (I34763,I34695,I34746);
DFFARX1 I_1897 (I34763,I2507,I34339,I34328,);
nor I_1898 (I34794,I34656,I34729);
nor I_1899 (I34316,I34520,I34794);
nor I_1900 (I34310,I34656,I34712);
not I_1901 (I34866,I2514);
DFFARX1 I_1902 (I1026977,I2507,I34866,I34892,);
DFFARX1 I_1903 (I34892,I2507,I34866,I34909,);
not I_1904 (I34917,I34909);
nand I_1905 (I34934,I1026971,I1026992);
and I_1906 (I34951,I34934,I1026977);
DFFARX1 I_1907 (I34951,I2507,I34866,I34977,);
DFFARX1 I_1908 (I34977,I2507,I34866,I34858,);
DFFARX1 I_1909 (I34977,I2507,I34866,I34849,);
DFFARX1 I_1910 (I1026974,I2507,I34866,I35022,);
nand I_1911 (I35030,I35022,I1026983);
not I_1912 (I35047,I35030);
nor I_1913 (I34846,I34892,I35047);
DFFARX1 I_1914 (I1026971,I2507,I34866,I35087,);
not I_1915 (I35095,I35087);
nor I_1916 (I34852,I35095,I34917);
nand I_1917 (I34840,I35095,I35030);
nand I_1918 (I35140,I1026974,I1026989);
and I_1919 (I35157,I35140,I1026980);
DFFARX1 I_1920 (I35157,I2507,I34866,I35183,);
nor I_1921 (I35191,I35183,I34892);
DFFARX1 I_1922 (I35191,I2507,I34866,I34834,);
not I_1923 (I35222,I35183);
nor I_1924 (I35239,I1026986,I1026989);
not I_1925 (I35256,I35239);
nor I_1926 (I35273,I35030,I35256);
nor I_1927 (I35290,I35222,I35273);
DFFARX1 I_1928 (I35290,I2507,I34866,I34855,);
nor I_1929 (I35321,I35183,I35256);
nor I_1930 (I34843,I35047,I35321);
nor I_1931 (I34837,I35183,I35239);
not I_1932 (I35393,I2514);
DFFARX1 I_1933 (I897285,I2507,I35393,I35419,);
DFFARX1 I_1934 (I35419,I2507,I35393,I35436,);
not I_1935 (I35444,I35436);
nand I_1936 (I35461,I897261,I897288);
and I_1937 (I35478,I35461,I897273);
DFFARX1 I_1938 (I35478,I2507,I35393,I35504,);
DFFARX1 I_1939 (I35504,I2507,I35393,I35385,);
DFFARX1 I_1940 (I35504,I2507,I35393,I35376,);
DFFARX1 I_1941 (I897279,I2507,I35393,I35549,);
nand I_1942 (I35557,I35549,I897264);
not I_1943 (I35574,I35557);
nor I_1944 (I35373,I35419,I35574);
DFFARX1 I_1945 (I897282,I2507,I35393,I35614,);
not I_1946 (I35622,I35614);
nor I_1947 (I35379,I35622,I35444);
nand I_1948 (I35367,I35622,I35557);
nand I_1949 (I35667,I897267,I897270);
and I_1950 (I35684,I35667,I897261);
DFFARX1 I_1951 (I35684,I2507,I35393,I35710,);
nor I_1952 (I35718,I35710,I35419);
DFFARX1 I_1953 (I35718,I2507,I35393,I35361,);
not I_1954 (I35749,I35710);
nor I_1955 (I35766,I897276,I897270);
not I_1956 (I35783,I35766);
nor I_1957 (I35800,I35557,I35783);
nor I_1958 (I35817,I35749,I35800);
DFFARX1 I_1959 (I35817,I2507,I35393,I35382,);
nor I_1960 (I35848,I35710,I35783);
nor I_1961 (I35370,I35574,I35848);
nor I_1962 (I35364,I35710,I35766);
not I_1963 (I35920,I2514);
DFFARX1 I_1964 (I901807,I2507,I35920,I35946,);
DFFARX1 I_1965 (I35946,I2507,I35920,I35963,);
not I_1966 (I35971,I35963);
nand I_1967 (I35988,I901783,I901810);
and I_1968 (I36005,I35988,I901795);
DFFARX1 I_1969 (I36005,I2507,I35920,I36031,);
DFFARX1 I_1970 (I36031,I2507,I35920,I35912,);
DFFARX1 I_1971 (I36031,I2507,I35920,I35903,);
DFFARX1 I_1972 (I901801,I2507,I35920,I36076,);
nand I_1973 (I36084,I36076,I901786);
not I_1974 (I36101,I36084);
nor I_1975 (I35900,I35946,I36101);
DFFARX1 I_1976 (I901804,I2507,I35920,I36141,);
not I_1977 (I36149,I36141);
nor I_1978 (I35906,I36149,I35971);
nand I_1979 (I35894,I36149,I36084);
nand I_1980 (I36194,I901789,I901792);
and I_1981 (I36211,I36194,I901783);
DFFARX1 I_1982 (I36211,I2507,I35920,I36237,);
nor I_1983 (I36245,I36237,I35946);
DFFARX1 I_1984 (I36245,I2507,I35920,I35888,);
not I_1985 (I36276,I36237);
nor I_1986 (I36293,I901798,I901792);
not I_1987 (I36310,I36293);
nor I_1988 (I36327,I36084,I36310);
nor I_1989 (I36344,I36276,I36327);
DFFARX1 I_1990 (I36344,I2507,I35920,I35909,);
nor I_1991 (I36375,I36237,I36310);
nor I_1992 (I35897,I36101,I36375);
nor I_1993 (I35891,I36237,I36293);
not I_1994 (I36447,I2514);
DFFARX1 I_1995 (I866024,I2507,I36447,I36473,);
DFFARX1 I_1996 (I36473,I2507,I36447,I36490,);
not I_1997 (I36498,I36490);
nand I_1998 (I36515,I866015,I866036);
and I_1999 (I36532,I36515,I866018);
DFFARX1 I_2000 (I36532,I2507,I36447,I36558,);
DFFARX1 I_2001 (I36558,I2507,I36447,I36439,);
DFFARX1 I_2002 (I36558,I2507,I36447,I36430,);
DFFARX1 I_2003 (I866018,I2507,I36447,I36603,);
nand I_2004 (I36611,I36603,I866033);
not I_2005 (I36628,I36611);
nor I_2006 (I36427,I36473,I36628);
DFFARX1 I_2007 (I866027,I2507,I36447,I36668,);
not I_2008 (I36676,I36668);
nor I_2009 (I36433,I36676,I36498);
nand I_2010 (I36421,I36676,I36611);
nand I_2011 (I36721,I866021,I866030);
and I_2012 (I36738,I36721,I866015);
DFFARX1 I_2013 (I36738,I2507,I36447,I36764,);
nor I_2014 (I36772,I36764,I36473);
DFFARX1 I_2015 (I36772,I2507,I36447,I36415,);
not I_2016 (I36803,I36764);
nor I_2017 (I36820,I866021,I866030);
not I_2018 (I36837,I36820);
nor I_2019 (I36854,I36611,I36837);
nor I_2020 (I36871,I36803,I36854);
DFFARX1 I_2021 (I36871,I2507,I36447,I36436,);
nor I_2022 (I36902,I36764,I36837);
nor I_2023 (I36424,I36628,I36902);
nor I_2024 (I36418,I36764,I36820);
not I_2025 (I36974,I2514);
DFFARX1 I_2026 (I1299199,I2507,I36974,I37000,);
DFFARX1 I_2027 (I37000,I2507,I36974,I37017,);
not I_2028 (I37025,I37017);
nand I_2029 (I37042,I1299190,I1299196);
and I_2030 (I37059,I37042,I1299175);
DFFARX1 I_2031 (I37059,I2507,I36974,I37085,);
DFFARX1 I_2032 (I37085,I2507,I36974,I36966,);
DFFARX1 I_2033 (I37085,I2507,I36974,I36957,);
DFFARX1 I_2034 (I1299193,I2507,I36974,I37130,);
nand I_2035 (I37138,I37130,I1299175);
not I_2036 (I37155,I37138);
nor I_2037 (I36954,I37000,I37155);
DFFARX1 I_2038 (I1299187,I2507,I36974,I37195,);
not I_2039 (I37203,I37195);
nor I_2040 (I36960,I37203,I37025);
nand I_2041 (I36948,I37203,I37138);
nand I_2042 (I37248,I1299181,I1299202);
and I_2043 (I37265,I37248,I1299184);
DFFARX1 I_2044 (I37265,I2507,I36974,I37291,);
nor I_2045 (I37299,I37291,I37000);
DFFARX1 I_2046 (I37299,I2507,I36974,I36942,);
not I_2047 (I37330,I37291);
nor I_2048 (I37347,I1299178,I1299202);
not I_2049 (I37364,I37347);
nor I_2050 (I37381,I37138,I37364);
nor I_2051 (I37398,I37330,I37381);
DFFARX1 I_2052 (I37398,I2507,I36974,I36963,);
nor I_2053 (I37429,I37291,I37364);
nor I_2054 (I36951,I37155,I37429);
nor I_2055 (I36945,I37291,I37347);
not I_2056 (I37501,I2514);
DFFARX1 I_2057 (I689680,I2507,I37501,I37527,);
DFFARX1 I_2058 (I37527,I2507,I37501,I37544,);
not I_2059 (I37552,I37544);
nand I_2060 (I37569,I689695,I689698);
and I_2061 (I37586,I37569,I689677);
DFFARX1 I_2062 (I37586,I2507,I37501,I37612,);
DFFARX1 I_2063 (I37612,I2507,I37501,I37493,);
DFFARX1 I_2064 (I37612,I2507,I37501,I37484,);
DFFARX1 I_2065 (I689683,I2507,I37501,I37657,);
nand I_2066 (I37665,I37657,I689689);
not I_2067 (I37682,I37665);
nor I_2068 (I37481,I37527,I37682);
DFFARX1 I_2069 (I689677,I2507,I37501,I37722,);
not I_2070 (I37730,I37722);
nor I_2071 (I37487,I37730,I37552);
nand I_2072 (I37475,I37730,I37665);
nand I_2073 (I37775,I689692,I689674);
and I_2074 (I37792,I37775,I689686);
DFFARX1 I_2075 (I37792,I2507,I37501,I37818,);
nor I_2076 (I37826,I37818,I37527);
DFFARX1 I_2077 (I37826,I2507,I37501,I37469,);
not I_2078 (I37857,I37818);
nor I_2079 (I37874,I689674,I689674);
not I_2080 (I37891,I37874);
nor I_2081 (I37908,I37665,I37891);
nor I_2082 (I37925,I37857,I37908);
DFFARX1 I_2083 (I37925,I2507,I37501,I37490,);
nor I_2084 (I37956,I37818,I37891);
nor I_2085 (I37478,I37682,I37956);
nor I_2086 (I37472,I37818,I37874);
not I_2087 (I38028,I2514);
DFFARX1 I_2088 (I503023,I2507,I38028,I38054,);
DFFARX1 I_2089 (I38054,I2507,I38028,I38071,);
not I_2090 (I38079,I38071);
nand I_2091 (I38096,I503029,I503017);
and I_2092 (I38113,I38096,I503014);
DFFARX1 I_2093 (I38113,I2507,I38028,I38139,);
DFFARX1 I_2094 (I38139,I2507,I38028,I38020,);
DFFARX1 I_2095 (I38139,I2507,I38028,I38011,);
DFFARX1 I_2096 (I503026,I2507,I38028,I38184,);
nand I_2097 (I38192,I38184,I503020);
not I_2098 (I38209,I38192);
nor I_2099 (I38008,I38054,I38209);
DFFARX1 I_2100 (I503038,I2507,I38028,I38249,);
not I_2101 (I38257,I38249);
nor I_2102 (I38014,I38257,I38079);
nand I_2103 (I38002,I38257,I38192);
nand I_2104 (I38302,I503032,I503035);
and I_2105 (I38319,I38302,I503017);
DFFARX1 I_2106 (I38319,I2507,I38028,I38345,);
nor I_2107 (I38353,I38345,I38054);
DFFARX1 I_2108 (I38353,I2507,I38028,I37996,);
not I_2109 (I38384,I38345);
nor I_2110 (I38401,I503014,I503035);
not I_2111 (I38418,I38401);
nor I_2112 (I38435,I38192,I38418);
nor I_2113 (I38452,I38384,I38435);
DFFARX1 I_2114 (I38452,I2507,I38028,I38017,);
nor I_2115 (I38483,I38345,I38418);
nor I_2116 (I38005,I38209,I38483);
nor I_2117 (I37999,I38345,I38401);
not I_2118 (I38555,I2514);
DFFARX1 I_2119 (I273932,I2507,I38555,I38581,);
DFFARX1 I_2120 (I38581,I2507,I38555,I38598,);
not I_2121 (I38606,I38598);
nand I_2122 (I38623,I273929,I273923);
and I_2123 (I38640,I38623,I273917);
DFFARX1 I_2124 (I38640,I2507,I38555,I38666,);
DFFARX1 I_2125 (I38666,I2507,I38555,I38547,);
DFFARX1 I_2126 (I38666,I2507,I38555,I38538,);
DFFARX1 I_2127 (I273905,I2507,I38555,I38711,);
nand I_2128 (I38719,I38711,I273914);
not I_2129 (I38736,I38719);
nor I_2130 (I38535,I38581,I38736);
DFFARX1 I_2131 (I273911,I2507,I38555,I38776,);
not I_2132 (I38784,I38776);
nor I_2133 (I38541,I38784,I38606);
nand I_2134 (I38529,I38784,I38719);
nand I_2135 (I38829,I273908,I273926);
and I_2136 (I38846,I38829,I273905);
DFFARX1 I_2137 (I38846,I2507,I38555,I38872,);
nor I_2138 (I38880,I38872,I38581);
DFFARX1 I_2139 (I38880,I2507,I38555,I38523,);
not I_2140 (I38911,I38872);
nor I_2141 (I38928,I273920,I273926);
not I_2142 (I38945,I38928);
nor I_2143 (I38962,I38719,I38945);
nor I_2144 (I38979,I38911,I38962);
DFFARX1 I_2145 (I38979,I2507,I38555,I38544,);
nor I_2146 (I39010,I38872,I38945);
nor I_2147 (I38532,I38736,I39010);
nor I_2148 (I38526,I38872,I38928);
not I_2149 (I39082,I2514);
DFFARX1 I_2150 (I148451,I2507,I39082,I39108,);
DFFARX1 I_2151 (I39108,I2507,I39082,I39125,);
not I_2152 (I39133,I39125);
nand I_2153 (I39150,I148469,I148454);
and I_2154 (I39167,I39150,I148457);
DFFARX1 I_2155 (I39167,I2507,I39082,I39193,);
DFFARX1 I_2156 (I39193,I2507,I39082,I39074,);
DFFARX1 I_2157 (I39193,I2507,I39082,I39065,);
DFFARX1 I_2158 (I148445,I2507,I39082,I39238,);
nand I_2159 (I39246,I39238,I148448);
not I_2160 (I39263,I39246);
nor I_2161 (I39062,I39108,I39263);
DFFARX1 I_2162 (I148460,I2507,I39082,I39303,);
not I_2163 (I39311,I39303);
nor I_2164 (I39068,I39311,I39133);
nand I_2165 (I39056,I39311,I39246);
nand I_2166 (I39356,I148466,I148463);
and I_2167 (I39373,I39356,I148448);
DFFARX1 I_2168 (I39373,I2507,I39082,I39399,);
nor I_2169 (I39407,I39399,I39108);
DFFARX1 I_2170 (I39407,I2507,I39082,I39050,);
not I_2171 (I39438,I39399);
nor I_2172 (I39455,I148445,I148463);
not I_2173 (I39472,I39455);
nor I_2174 (I39489,I39246,I39472);
nor I_2175 (I39506,I39438,I39489);
DFFARX1 I_2176 (I39506,I2507,I39082,I39071,);
nor I_2177 (I39537,I39399,I39472);
nor I_2178 (I39059,I39263,I39537);
nor I_2179 (I39053,I39399,I39455);
not I_2180 (I39609,I2514);
DFFARX1 I_2181 (I1130644,I2507,I39609,I39635,);
DFFARX1 I_2182 (I39635,I2507,I39609,I39652,);
not I_2183 (I39660,I39652);
nand I_2184 (I39677,I1130632,I1130623);
and I_2185 (I39694,I39677,I1130620);
DFFARX1 I_2186 (I39694,I2507,I39609,I39720,);
DFFARX1 I_2187 (I39720,I2507,I39609,I39601,);
DFFARX1 I_2188 (I39720,I2507,I39609,I39592,);
DFFARX1 I_2189 (I1130626,I2507,I39609,I39765,);
nand I_2190 (I39773,I39765,I1130638);
not I_2191 (I39790,I39773);
nor I_2192 (I39589,I39635,I39790);
DFFARX1 I_2193 (I1130635,I2507,I39609,I39830,);
not I_2194 (I39838,I39830);
nor I_2195 (I39595,I39838,I39660);
nand I_2196 (I39583,I39838,I39773);
nand I_2197 (I39883,I1130629,I1130623);
and I_2198 (I39900,I39883,I1130641);
DFFARX1 I_2199 (I39900,I2507,I39609,I39926,);
nor I_2200 (I39934,I39926,I39635);
DFFARX1 I_2201 (I39934,I2507,I39609,I39577,);
not I_2202 (I39965,I39926);
nor I_2203 (I39982,I1130620,I1130623);
not I_2204 (I39999,I39982);
nor I_2205 (I40016,I39773,I39999);
nor I_2206 (I40033,I39965,I40016);
DFFARX1 I_2207 (I40033,I2507,I39609,I39598,);
nor I_2208 (I40064,I39926,I39999);
nor I_2209 (I39586,I39790,I40064);
nor I_2210 (I39580,I39926,I39982);
not I_2211 (I40136,I2514);
DFFARX1 I_2212 (I514328,I2507,I40136,I40162,);
DFFARX1 I_2213 (I40162,I2507,I40136,I40179,);
not I_2214 (I40187,I40179);
nand I_2215 (I40204,I514334,I514322);
and I_2216 (I40221,I40204,I514319);
DFFARX1 I_2217 (I40221,I2507,I40136,I40247,);
DFFARX1 I_2218 (I40247,I2507,I40136,I40128,);
DFFARX1 I_2219 (I40247,I2507,I40136,I40119,);
DFFARX1 I_2220 (I514331,I2507,I40136,I40292,);
nand I_2221 (I40300,I40292,I514325);
not I_2222 (I40317,I40300);
nor I_2223 (I40116,I40162,I40317);
DFFARX1 I_2224 (I514343,I2507,I40136,I40357,);
not I_2225 (I40365,I40357);
nor I_2226 (I40122,I40365,I40187);
nand I_2227 (I40110,I40365,I40300);
nand I_2228 (I40410,I514337,I514340);
and I_2229 (I40427,I40410,I514322);
DFFARX1 I_2230 (I40427,I2507,I40136,I40453,);
nor I_2231 (I40461,I40453,I40162);
DFFARX1 I_2232 (I40461,I2507,I40136,I40104,);
not I_2233 (I40492,I40453);
nor I_2234 (I40509,I514319,I514340);
not I_2235 (I40526,I40509);
nor I_2236 (I40543,I40300,I40526);
nor I_2237 (I40560,I40492,I40543);
DFFARX1 I_2238 (I40560,I2507,I40136,I40125,);
nor I_2239 (I40591,I40453,I40526);
nor I_2240 (I40113,I40317,I40591);
nor I_2241 (I40107,I40453,I40509);
not I_2242 (I40663,I2514);
DFFARX1 I_2243 (I49593,I2507,I40663,I40689,);
DFFARX1 I_2244 (I40689,I2507,I40663,I40706,);
not I_2245 (I40714,I40706);
nand I_2246 (I40731,I49593,I49608);
and I_2247 (I40748,I40731,I49611);
DFFARX1 I_2248 (I40748,I2507,I40663,I40774,);
DFFARX1 I_2249 (I40774,I2507,I40663,I40655,);
DFFARX1 I_2250 (I40774,I2507,I40663,I40646,);
DFFARX1 I_2251 (I49605,I2507,I40663,I40819,);
nand I_2252 (I40827,I40819,I49614);
not I_2253 (I40844,I40827);
nor I_2254 (I40643,I40689,I40844);
DFFARX1 I_2255 (I49590,I2507,I40663,I40884,);
not I_2256 (I40892,I40884);
nor I_2257 (I40649,I40892,I40714);
nand I_2258 (I40637,I40892,I40827);
nand I_2259 (I40937,I49590,I49596);
and I_2260 (I40954,I40937,I49599);
DFFARX1 I_2261 (I40954,I2507,I40663,I40980,);
nor I_2262 (I40988,I40980,I40689);
DFFARX1 I_2263 (I40988,I2507,I40663,I40631,);
not I_2264 (I41019,I40980);
nor I_2265 (I41036,I49602,I49596);
not I_2266 (I41053,I41036);
nor I_2267 (I41070,I40827,I41053);
nor I_2268 (I41087,I41019,I41070);
DFFARX1 I_2269 (I41087,I2507,I40663,I40652,);
nor I_2270 (I41118,I40980,I41053);
nor I_2271 (I40640,I40844,I41118);
nor I_2272 (I40634,I40980,I41036);
not I_2273 (I41190,I2514);
DFFARX1 I_2274 (I1132956,I2507,I41190,I41216,);
DFFARX1 I_2275 (I41216,I2507,I41190,I41233,);
not I_2276 (I41241,I41233);
nand I_2277 (I41258,I1132944,I1132935);
and I_2278 (I41275,I41258,I1132932);
DFFARX1 I_2279 (I41275,I2507,I41190,I41301,);
DFFARX1 I_2280 (I41301,I2507,I41190,I41182,);
DFFARX1 I_2281 (I41301,I2507,I41190,I41173,);
DFFARX1 I_2282 (I1132938,I2507,I41190,I41346,);
nand I_2283 (I41354,I41346,I1132950);
not I_2284 (I41371,I41354);
nor I_2285 (I41170,I41216,I41371);
DFFARX1 I_2286 (I1132947,I2507,I41190,I41411,);
not I_2287 (I41419,I41411);
nor I_2288 (I41176,I41419,I41241);
nand I_2289 (I41164,I41419,I41354);
nand I_2290 (I41464,I1132941,I1132935);
and I_2291 (I41481,I41464,I1132953);
DFFARX1 I_2292 (I41481,I2507,I41190,I41507,);
nor I_2293 (I41515,I41507,I41216);
DFFARX1 I_2294 (I41515,I2507,I41190,I41158,);
not I_2295 (I41546,I41507);
nor I_2296 (I41563,I1132932,I1132935);
not I_2297 (I41580,I41563);
nor I_2298 (I41597,I41354,I41580);
nor I_2299 (I41614,I41546,I41597);
DFFARX1 I_2300 (I41614,I2507,I41190,I41179,);
nor I_2301 (I41645,I41507,I41580);
nor I_2302 (I41167,I41371,I41645);
nor I_2303 (I41161,I41507,I41563);
not I_2304 (I41717,I2514);
DFFARX1 I_2305 (I757306,I2507,I41717,I41743,);
DFFARX1 I_2306 (I41743,I2507,I41717,I41760,);
not I_2307 (I41768,I41760);
nand I_2308 (I41785,I757321,I757324);
and I_2309 (I41802,I41785,I757303);
DFFARX1 I_2310 (I41802,I2507,I41717,I41828,);
DFFARX1 I_2311 (I41828,I2507,I41717,I41709,);
DFFARX1 I_2312 (I41828,I2507,I41717,I41700,);
DFFARX1 I_2313 (I757309,I2507,I41717,I41873,);
nand I_2314 (I41881,I41873,I757315);
not I_2315 (I41898,I41881);
nor I_2316 (I41697,I41743,I41898);
DFFARX1 I_2317 (I757303,I2507,I41717,I41938,);
not I_2318 (I41946,I41938);
nor I_2319 (I41703,I41946,I41768);
nand I_2320 (I41691,I41946,I41881);
nand I_2321 (I41991,I757318,I757300);
and I_2322 (I42008,I41991,I757312);
DFFARX1 I_2323 (I42008,I2507,I41717,I42034,);
nor I_2324 (I42042,I42034,I41743);
DFFARX1 I_2325 (I42042,I2507,I41717,I41685,);
not I_2326 (I42073,I42034);
nor I_2327 (I42090,I757300,I757300);
not I_2328 (I42107,I42090);
nor I_2329 (I42124,I41881,I42107);
nor I_2330 (I42141,I42073,I42124);
DFFARX1 I_2331 (I42141,I2507,I41717,I41706,);
nor I_2332 (I42172,I42034,I42107);
nor I_2333 (I41694,I41898,I42172);
nor I_2334 (I41688,I42034,I42090);
not I_2335 (I42244,I2514);
DFFARX1 I_2336 (I168086,I2507,I42244,I42270,);
DFFARX1 I_2337 (I42270,I2507,I42244,I42287,);
not I_2338 (I42295,I42287);
nand I_2339 (I42312,I168104,I168089);
and I_2340 (I42329,I42312,I168092);
DFFARX1 I_2341 (I42329,I2507,I42244,I42355,);
DFFARX1 I_2342 (I42355,I2507,I42244,I42236,);
DFFARX1 I_2343 (I42355,I2507,I42244,I42227,);
DFFARX1 I_2344 (I168080,I2507,I42244,I42400,);
nand I_2345 (I42408,I42400,I168083);
not I_2346 (I42425,I42408);
nor I_2347 (I42224,I42270,I42425);
DFFARX1 I_2348 (I168095,I2507,I42244,I42465,);
not I_2349 (I42473,I42465);
nor I_2350 (I42230,I42473,I42295);
nand I_2351 (I42218,I42473,I42408);
nand I_2352 (I42518,I168101,I168098);
and I_2353 (I42535,I42518,I168083);
DFFARX1 I_2354 (I42535,I2507,I42244,I42561,);
nor I_2355 (I42569,I42561,I42270);
DFFARX1 I_2356 (I42569,I2507,I42244,I42212,);
not I_2357 (I42600,I42561);
nor I_2358 (I42617,I168080,I168098);
not I_2359 (I42634,I42617);
nor I_2360 (I42651,I42408,I42634);
nor I_2361 (I42668,I42600,I42651);
DFFARX1 I_2362 (I42668,I2507,I42244,I42233,);
nor I_2363 (I42699,I42561,I42634);
nor I_2364 (I42221,I42425,I42699);
nor I_2365 (I42215,I42561,I42617);
not I_2366 (I42771,I2514);
DFFARX1 I_2367 (I295012,I2507,I42771,I42797,);
DFFARX1 I_2368 (I42797,I2507,I42771,I42814,);
not I_2369 (I42822,I42814);
nand I_2370 (I42839,I295009,I295003);
and I_2371 (I42856,I42839,I294997);
DFFARX1 I_2372 (I42856,I2507,I42771,I42882,);
DFFARX1 I_2373 (I42882,I2507,I42771,I42763,);
DFFARX1 I_2374 (I42882,I2507,I42771,I42754,);
DFFARX1 I_2375 (I294985,I2507,I42771,I42927,);
nand I_2376 (I42935,I42927,I294994);
not I_2377 (I42952,I42935);
nor I_2378 (I42751,I42797,I42952);
DFFARX1 I_2379 (I294991,I2507,I42771,I42992,);
not I_2380 (I43000,I42992);
nor I_2381 (I42757,I43000,I42822);
nand I_2382 (I42745,I43000,I42935);
nand I_2383 (I43045,I294988,I295006);
and I_2384 (I43062,I43045,I294985);
DFFARX1 I_2385 (I43062,I2507,I42771,I43088,);
nor I_2386 (I43096,I43088,I42797);
DFFARX1 I_2387 (I43096,I2507,I42771,I42739,);
not I_2388 (I43127,I43088);
nor I_2389 (I43144,I295000,I295006);
not I_2390 (I43161,I43144);
nor I_2391 (I43178,I42935,I43161);
nor I_2392 (I43195,I43127,I43178);
DFFARX1 I_2393 (I43195,I2507,I42771,I42760,);
nor I_2394 (I43226,I43088,I43161);
nor I_2395 (I42748,I42952,I43226);
nor I_2396 (I42742,I43088,I43144);
not I_2397 (I43298,I2514);
DFFARX1 I_2398 (I564841,I2507,I43298,I43324,);
DFFARX1 I_2399 (I43324,I2507,I43298,I43341,);
not I_2400 (I43349,I43341);
nand I_2401 (I43366,I564826,I564844);
and I_2402 (I43383,I43366,I564838);
DFFARX1 I_2403 (I43383,I2507,I43298,I43409,);
DFFARX1 I_2404 (I43409,I2507,I43298,I43290,);
DFFARX1 I_2405 (I43409,I2507,I43298,I43281,);
DFFARX1 I_2406 (I564835,I2507,I43298,I43454,);
nand I_2407 (I43462,I43454,I564826);
not I_2408 (I43479,I43462);
nor I_2409 (I43278,I43324,I43479);
DFFARX1 I_2410 (I564829,I2507,I43298,I43519,);
not I_2411 (I43527,I43519);
nor I_2412 (I43284,I43527,I43349);
nand I_2413 (I43272,I43527,I43462);
nand I_2414 (I43572,I564850,I564832);
and I_2415 (I43589,I43572,I564847);
DFFARX1 I_2416 (I43589,I2507,I43298,I43615,);
nor I_2417 (I43623,I43615,I43324);
DFFARX1 I_2418 (I43623,I2507,I43298,I43266,);
not I_2419 (I43654,I43615);
nor I_2420 (I43671,I564829,I564832);
not I_2421 (I43688,I43671);
nor I_2422 (I43705,I43462,I43688);
nor I_2423 (I43722,I43654,I43705);
DFFARX1 I_2424 (I43722,I2507,I43298,I43287,);
nor I_2425 (I43753,I43615,I43688);
nor I_2426 (I43275,I43479,I43753);
nor I_2427 (I43269,I43615,I43671);
not I_2428 (I43825,I2514);
DFFARX1 I_2429 (I1131800,I2507,I43825,I43851,);
DFFARX1 I_2430 (I43851,I2507,I43825,I43868,);
not I_2431 (I43876,I43868);
nand I_2432 (I43893,I1131788,I1131779);
and I_2433 (I43910,I43893,I1131776);
DFFARX1 I_2434 (I43910,I2507,I43825,I43936,);
DFFARX1 I_2435 (I43936,I2507,I43825,I43817,);
DFFARX1 I_2436 (I43936,I2507,I43825,I43808,);
DFFARX1 I_2437 (I1131782,I2507,I43825,I43981,);
nand I_2438 (I43989,I43981,I1131794);
not I_2439 (I44006,I43989);
nor I_2440 (I43805,I43851,I44006);
DFFARX1 I_2441 (I1131791,I2507,I43825,I44046,);
not I_2442 (I44054,I44046);
nor I_2443 (I43811,I44054,I43876);
nand I_2444 (I43799,I44054,I43989);
nand I_2445 (I44099,I1131785,I1131779);
and I_2446 (I44116,I44099,I1131797);
DFFARX1 I_2447 (I44116,I2507,I43825,I44142,);
nor I_2448 (I44150,I44142,I43851);
DFFARX1 I_2449 (I44150,I2507,I43825,I43793,);
not I_2450 (I44181,I44142);
nor I_2451 (I44198,I1131776,I1131779);
not I_2452 (I44215,I44198);
nor I_2453 (I44232,I43989,I44215);
nor I_2454 (I44249,I44181,I44232);
DFFARX1 I_2455 (I44249,I2507,I43825,I43814,);
nor I_2456 (I44280,I44142,I44215);
nor I_2457 (I43802,I44006,I44280);
nor I_2458 (I43796,I44142,I44198);
not I_2459 (I44352,I2514);
DFFARX1 I_2460 (I679854,I2507,I44352,I44378,);
DFFARX1 I_2461 (I44378,I2507,I44352,I44395,);
not I_2462 (I44403,I44395);
nand I_2463 (I44420,I679869,I679872);
and I_2464 (I44437,I44420,I679851);
DFFARX1 I_2465 (I44437,I2507,I44352,I44463,);
DFFARX1 I_2466 (I44463,I2507,I44352,I44344,);
DFFARX1 I_2467 (I44463,I2507,I44352,I44335,);
DFFARX1 I_2468 (I679857,I2507,I44352,I44508,);
nand I_2469 (I44516,I44508,I679863);
not I_2470 (I44533,I44516);
nor I_2471 (I44332,I44378,I44533);
DFFARX1 I_2472 (I679851,I2507,I44352,I44573,);
not I_2473 (I44581,I44573);
nor I_2474 (I44338,I44581,I44403);
nand I_2475 (I44326,I44581,I44516);
nand I_2476 (I44626,I679866,I679848);
and I_2477 (I44643,I44626,I679860);
DFFARX1 I_2478 (I44643,I2507,I44352,I44669,);
nor I_2479 (I44677,I44669,I44378);
DFFARX1 I_2480 (I44677,I2507,I44352,I44320,);
not I_2481 (I44708,I44669);
nor I_2482 (I44725,I679848,I679848);
not I_2483 (I44742,I44725);
nor I_2484 (I44759,I44516,I44742);
nor I_2485 (I44776,I44708,I44759);
DFFARX1 I_2486 (I44776,I2507,I44352,I44341,);
nor I_2487 (I44807,I44669,I44742);
nor I_2488 (I44329,I44533,I44807);
nor I_2489 (I44323,I44669,I44725);
not I_2490 (I44879,I2514);
DFFARX1 I_2491 (I1013513,I2507,I44879,I44905,);
DFFARX1 I_2492 (I44905,I2507,I44879,I44922,);
not I_2493 (I44930,I44922);
nand I_2494 (I44947,I1013507,I1013528);
and I_2495 (I44964,I44947,I1013513);
DFFARX1 I_2496 (I44964,I2507,I44879,I44990,);
DFFARX1 I_2497 (I44990,I2507,I44879,I44871,);
DFFARX1 I_2498 (I44990,I2507,I44879,I44862,);
DFFARX1 I_2499 (I1013510,I2507,I44879,I45035,);
nand I_2500 (I45043,I45035,I1013519);
not I_2501 (I45060,I45043);
nor I_2502 (I44859,I44905,I45060);
DFFARX1 I_2503 (I1013507,I2507,I44879,I45100,);
not I_2504 (I45108,I45100);
nor I_2505 (I44865,I45108,I44930);
nand I_2506 (I44853,I45108,I45043);
nand I_2507 (I45153,I1013510,I1013525);
and I_2508 (I45170,I45153,I1013516);
DFFARX1 I_2509 (I45170,I2507,I44879,I45196,);
nor I_2510 (I45204,I45196,I44905);
DFFARX1 I_2511 (I45204,I2507,I44879,I44847,);
not I_2512 (I45235,I45196);
nor I_2513 (I45252,I1013522,I1013525);
not I_2514 (I45269,I45252);
nor I_2515 (I45286,I45043,I45269);
nor I_2516 (I45303,I45235,I45286);
DFFARX1 I_2517 (I45303,I2507,I44879,I44868,);
nor I_2518 (I45334,I45196,I45269);
nor I_2519 (I44856,I45060,I45334);
nor I_2520 (I44850,I45196,I45252);
not I_2521 (I45406,I2514);
DFFARX1 I_2522 (I655000,I2507,I45406,I45432,);
DFFARX1 I_2523 (I45432,I2507,I45406,I45449,);
not I_2524 (I45457,I45449);
nand I_2525 (I45474,I655015,I655018);
and I_2526 (I45491,I45474,I654997);
DFFARX1 I_2527 (I45491,I2507,I45406,I45517,);
DFFARX1 I_2528 (I45517,I2507,I45406,I45398,);
DFFARX1 I_2529 (I45517,I2507,I45406,I45389,);
DFFARX1 I_2530 (I655003,I2507,I45406,I45562,);
nand I_2531 (I45570,I45562,I655009);
not I_2532 (I45587,I45570);
nor I_2533 (I45386,I45432,I45587);
DFFARX1 I_2534 (I654997,I2507,I45406,I45627,);
not I_2535 (I45635,I45627);
nor I_2536 (I45392,I45635,I45457);
nand I_2537 (I45380,I45635,I45570);
nand I_2538 (I45680,I655012,I654994);
and I_2539 (I45697,I45680,I655006);
DFFARX1 I_2540 (I45697,I2507,I45406,I45723,);
nor I_2541 (I45731,I45723,I45432);
DFFARX1 I_2542 (I45731,I2507,I45406,I45374,);
not I_2543 (I45762,I45723);
nor I_2544 (I45779,I654994,I654994);
not I_2545 (I45796,I45779);
nor I_2546 (I45813,I45570,I45796);
nor I_2547 (I45830,I45762,I45813);
DFFARX1 I_2548 (I45830,I2507,I45406,I45395,);
nor I_2549 (I45861,I45723,I45796);
nor I_2550 (I45383,I45587,I45861);
nor I_2551 (I45377,I45723,I45779);
not I_2552 (I45933,I2514);
DFFARX1 I_2553 (I565997,I2507,I45933,I45959,);
DFFARX1 I_2554 (I45959,I2507,I45933,I45976,);
not I_2555 (I45984,I45976);
nand I_2556 (I46001,I565982,I566000);
and I_2557 (I46018,I46001,I565994);
DFFARX1 I_2558 (I46018,I2507,I45933,I46044,);
DFFARX1 I_2559 (I46044,I2507,I45933,I45925,);
DFFARX1 I_2560 (I46044,I2507,I45933,I45916,);
DFFARX1 I_2561 (I565991,I2507,I45933,I46089,);
nand I_2562 (I46097,I46089,I565982);
not I_2563 (I46114,I46097);
nor I_2564 (I45913,I45959,I46114);
DFFARX1 I_2565 (I565985,I2507,I45933,I46154,);
not I_2566 (I46162,I46154);
nor I_2567 (I45919,I46162,I45984);
nand I_2568 (I45907,I46162,I46097);
nand I_2569 (I46207,I566006,I565988);
and I_2570 (I46224,I46207,I566003);
DFFARX1 I_2571 (I46224,I2507,I45933,I46250,);
nor I_2572 (I46258,I46250,I45959);
DFFARX1 I_2573 (I46258,I2507,I45933,I45901,);
not I_2574 (I46289,I46250);
nor I_2575 (I46306,I565985,I565988);
not I_2576 (I46323,I46306);
nor I_2577 (I46340,I46097,I46323);
nor I_2578 (I46357,I46289,I46340);
DFFARX1 I_2579 (I46357,I2507,I45933,I45922,);
nor I_2580 (I46388,I46250,I46323);
nor I_2581 (I45910,I46114,I46388);
nor I_2582 (I45904,I46250,I46306);
not I_2583 (I46460,I2514);
DFFARX1 I_2584 (I415855,I2507,I46460,I46486,);
DFFARX1 I_2585 (I46486,I2507,I46460,I46503,);
not I_2586 (I46511,I46503);
nand I_2587 (I46528,I415855,I415858);
and I_2588 (I46545,I46528,I415879);
DFFARX1 I_2589 (I46545,I2507,I46460,I46571,);
DFFARX1 I_2590 (I46571,I2507,I46460,I46452,);
DFFARX1 I_2591 (I46571,I2507,I46460,I46443,);
DFFARX1 I_2592 (I415867,I2507,I46460,I46616,);
nand I_2593 (I46624,I46616,I415870);
not I_2594 (I46641,I46624);
nor I_2595 (I46440,I46486,I46641);
DFFARX1 I_2596 (I415876,I2507,I46460,I46681,);
not I_2597 (I46689,I46681);
nor I_2598 (I46446,I46689,I46511);
nand I_2599 (I46434,I46689,I46624);
nand I_2600 (I46734,I415873,I415861);
and I_2601 (I46751,I46734,I415864);
DFFARX1 I_2602 (I46751,I2507,I46460,I46777,);
nor I_2603 (I46785,I46777,I46486);
DFFARX1 I_2604 (I46785,I2507,I46460,I46428,);
not I_2605 (I46816,I46777);
nor I_2606 (I46833,I415882,I415861);
not I_2607 (I46850,I46833);
nor I_2608 (I46867,I46624,I46850);
nor I_2609 (I46884,I46816,I46867);
DFFARX1 I_2610 (I46884,I2507,I46460,I46449,);
nor I_2611 (I46915,I46777,I46850);
nor I_2612 (I46437,I46641,I46915);
nor I_2613 (I46431,I46777,I46833);
not I_2614 (I46987,I2514);
DFFARX1 I_2615 (I1076890,I2507,I46987,I47013,);
DFFARX1 I_2616 (I47013,I2507,I46987,I47030,);
not I_2617 (I47038,I47030);
nand I_2618 (I47055,I1076878,I1076869);
and I_2619 (I47072,I47055,I1076866);
DFFARX1 I_2620 (I47072,I2507,I46987,I47098,);
DFFARX1 I_2621 (I47098,I2507,I46987,I46979,);
DFFARX1 I_2622 (I47098,I2507,I46987,I46970,);
DFFARX1 I_2623 (I1076872,I2507,I46987,I47143,);
nand I_2624 (I47151,I47143,I1076884);
not I_2625 (I47168,I47151);
nor I_2626 (I46967,I47013,I47168);
DFFARX1 I_2627 (I1076881,I2507,I46987,I47208,);
not I_2628 (I47216,I47208);
nor I_2629 (I46973,I47216,I47038);
nand I_2630 (I46961,I47216,I47151);
nand I_2631 (I47261,I1076875,I1076869);
and I_2632 (I47278,I47261,I1076887);
DFFARX1 I_2633 (I47278,I2507,I46987,I47304,);
nor I_2634 (I47312,I47304,I47013);
DFFARX1 I_2635 (I47312,I2507,I46987,I46955,);
not I_2636 (I47343,I47304);
nor I_2637 (I47360,I1076866,I1076869);
not I_2638 (I47377,I47360);
nor I_2639 (I47394,I47151,I47377);
nor I_2640 (I47411,I47343,I47394);
DFFARX1 I_2641 (I47411,I2507,I46987,I46976,);
nor I_2642 (I47442,I47304,I47377);
nor I_2643 (I46964,I47168,I47442);
nor I_2644 (I46958,I47304,I47360);
not I_2645 (I47514,I2514);
DFFARX1 I_2646 (I140130,I2507,I47514,I47540,);
DFFARX1 I_2647 (I47540,I2507,I47514,I47557,);
not I_2648 (I47565,I47557);
nand I_2649 (I47582,I140133,I140115);
and I_2650 (I47599,I47582,I140121);
DFFARX1 I_2651 (I47599,I2507,I47514,I47625,);
DFFARX1 I_2652 (I47625,I2507,I47514,I47506,);
DFFARX1 I_2653 (I47625,I2507,I47514,I47497,);
DFFARX1 I_2654 (I140124,I2507,I47514,I47670,);
nand I_2655 (I47678,I47670,I140115);
not I_2656 (I47695,I47678);
nor I_2657 (I47494,I47540,I47695);
DFFARX1 I_2658 (I140136,I2507,I47514,I47735,);
not I_2659 (I47743,I47735);
nor I_2660 (I47500,I47743,I47565);
nand I_2661 (I47488,I47743,I47678);
nand I_2662 (I47788,I140139,I140127);
and I_2663 (I47805,I47788,I140118);
DFFARX1 I_2664 (I47805,I2507,I47514,I47831,);
nor I_2665 (I47839,I47831,I47540);
DFFARX1 I_2666 (I47839,I2507,I47514,I47482,);
not I_2667 (I47870,I47831);
nor I_2668 (I47887,I140142,I140127);
not I_2669 (I47904,I47887);
nor I_2670 (I47921,I47678,I47904);
nor I_2671 (I47938,I47870,I47921);
DFFARX1 I_2672 (I47938,I2507,I47514,I47503,);
nor I_2673 (I47969,I47831,I47904);
nor I_2674 (I47491,I47695,I47969);
nor I_2675 (I47485,I47831,I47887);
not I_2676 (I48041,I2514);
DFFARX1 I_2677 (I943151,I2507,I48041,I48067,);
DFFARX1 I_2678 (I48067,I2507,I48041,I48084,);
not I_2679 (I48092,I48084);
nand I_2680 (I48109,I943127,I943154);
and I_2681 (I48126,I48109,I943139);
DFFARX1 I_2682 (I48126,I2507,I48041,I48152,);
DFFARX1 I_2683 (I48152,I2507,I48041,I48033,);
DFFARX1 I_2684 (I48152,I2507,I48041,I48024,);
DFFARX1 I_2685 (I943145,I2507,I48041,I48197,);
nand I_2686 (I48205,I48197,I943130);
not I_2687 (I48222,I48205);
nor I_2688 (I48021,I48067,I48222);
DFFARX1 I_2689 (I943148,I2507,I48041,I48262,);
not I_2690 (I48270,I48262);
nor I_2691 (I48027,I48270,I48092);
nand I_2692 (I48015,I48270,I48205);
nand I_2693 (I48315,I943133,I943136);
and I_2694 (I48332,I48315,I943127);
DFFARX1 I_2695 (I48332,I2507,I48041,I48358,);
nor I_2696 (I48366,I48358,I48067);
DFFARX1 I_2697 (I48366,I2507,I48041,I48009,);
not I_2698 (I48397,I48358);
nor I_2699 (I48414,I943142,I943136);
not I_2700 (I48431,I48414);
nor I_2701 (I48448,I48205,I48431);
nor I_2702 (I48465,I48397,I48448);
DFFARX1 I_2703 (I48465,I2507,I48041,I48030,);
nor I_2704 (I48496,I48358,I48431);
nor I_2705 (I48018,I48222,I48496);
nor I_2706 (I48012,I48358,I48414);
not I_2707 (I48568,I2514);
DFFARX1 I_2708 (I611653,I2507,I48568,I48594,);
not I_2709 (I48602,I48594);
nand I_2710 (I48619,I611665,I611650);
and I_2711 (I48636,I48619,I611644);
DFFARX1 I_2712 (I48636,I2507,I48568,I48662,);
DFFARX1 I_2713 (I611659,I2507,I48568,I48679,);
and I_2714 (I48687,I48679,I611647);
nor I_2715 (I48704,I48662,I48687);
DFFARX1 I_2716 (I48704,I2507,I48568,I48536,);
nand I_2717 (I48735,I48679,I611647);
nand I_2718 (I48752,I48602,I48735);
not I_2719 (I48548,I48752);
DFFARX1 I_2720 (I611656,I2507,I48568,I48792,);
DFFARX1 I_2721 (I48792,I2507,I48568,I48557,);
nand I_2722 (I48814,I611662,I611668);
and I_2723 (I48831,I48814,I611644);
DFFARX1 I_2724 (I48831,I2507,I48568,I48857,);
DFFARX1 I_2725 (I48857,I2507,I48568,I48874,);
not I_2726 (I48560,I48874);
not I_2727 (I48896,I48857);
nand I_2728 (I48545,I48896,I48735);
nor I_2729 (I48927,I611647,I611668);
not I_2730 (I48944,I48927);
nor I_2731 (I48961,I48896,I48944);
nor I_2732 (I48978,I48602,I48961);
DFFARX1 I_2733 (I48978,I2507,I48568,I48554,);
nor I_2734 (I49009,I48662,I48944);
nor I_2735 (I48542,I48857,I49009);
nor I_2736 (I48551,I48792,I48927);
nor I_2737 (I48539,I48662,I48927);
not I_2738 (I49095,I2514);
DFFARX1 I_2739 (I757890,I2507,I49095,I49121,);
not I_2740 (I49129,I49121);
nand I_2741 (I49146,I757881,I757899);
and I_2742 (I49163,I49146,I757878);
DFFARX1 I_2743 (I49163,I2507,I49095,I49189,);
DFFARX1 I_2744 (I757881,I2507,I49095,I49206,);
and I_2745 (I49214,I49206,I757884);
nor I_2746 (I49231,I49189,I49214);
DFFARX1 I_2747 (I49231,I2507,I49095,I49063,);
nand I_2748 (I49262,I49206,I757884);
nand I_2749 (I49279,I49129,I49262);
not I_2750 (I49075,I49279);
DFFARX1 I_2751 (I757878,I2507,I49095,I49319,);
DFFARX1 I_2752 (I49319,I2507,I49095,I49084,);
nand I_2753 (I49341,I757896,I757887);
and I_2754 (I49358,I49341,I757902);
DFFARX1 I_2755 (I49358,I2507,I49095,I49384,);
DFFARX1 I_2756 (I49384,I2507,I49095,I49401,);
not I_2757 (I49087,I49401);
not I_2758 (I49423,I49384);
nand I_2759 (I49072,I49423,I49262);
nor I_2760 (I49454,I757893,I757887);
not I_2761 (I49471,I49454);
nor I_2762 (I49488,I49423,I49471);
nor I_2763 (I49505,I49129,I49488);
DFFARX1 I_2764 (I49505,I2507,I49095,I49081,);
nor I_2765 (I49536,I49189,I49471);
nor I_2766 (I49069,I49384,I49536);
nor I_2767 (I49078,I49319,I49454);
nor I_2768 (I49066,I49189,I49454);
not I_2769 (I49622,I2514);
DFFARX1 I_2770 (I1138718,I2507,I49622,I49648,);
not I_2771 (I49656,I49648);
nand I_2772 (I49673,I1138733,I1138712);
and I_2773 (I49690,I49673,I1138715);
DFFARX1 I_2774 (I49690,I2507,I49622,I49716,);
DFFARX1 I_2775 (I1138736,I2507,I49622,I49733,);
and I_2776 (I49741,I49733,I1138715);
nor I_2777 (I49758,I49716,I49741);
DFFARX1 I_2778 (I49758,I2507,I49622,I49590,);
nand I_2779 (I49789,I49733,I1138715);
nand I_2780 (I49806,I49656,I49789);
not I_2781 (I49602,I49806);
DFFARX1 I_2782 (I1138712,I2507,I49622,I49846,);
DFFARX1 I_2783 (I49846,I2507,I49622,I49611,);
nand I_2784 (I49868,I1138724,I1138721);
and I_2785 (I49885,I49868,I1138727);
DFFARX1 I_2786 (I49885,I2507,I49622,I49911,);
DFFARX1 I_2787 (I49911,I2507,I49622,I49928,);
not I_2788 (I49614,I49928);
not I_2789 (I49950,I49911);
nand I_2790 (I49599,I49950,I49789);
nor I_2791 (I49981,I1138730,I1138721);
not I_2792 (I49998,I49981);
nor I_2793 (I50015,I49950,I49998);
nor I_2794 (I50032,I49656,I50015);
DFFARX1 I_2795 (I50032,I2507,I49622,I49608,);
nor I_2796 (I50063,I49716,I49998);
nor I_2797 (I49596,I49911,I50063);
nor I_2798 (I49605,I49846,I49981);
nor I_2799 (I49593,I49716,I49981);
not I_2800 (I50149,I2514);
DFFARX1 I_2801 (I306079,I2507,I50149,I50175,);
not I_2802 (I50183,I50175);
nand I_2803 (I50200,I306061,I306076);
and I_2804 (I50217,I50200,I306052);
DFFARX1 I_2805 (I50217,I2507,I50149,I50243,);
DFFARX1 I_2806 (I306055,I2507,I50149,I50260,);
and I_2807 (I50268,I50260,I306070);
nor I_2808 (I50285,I50243,I50268);
DFFARX1 I_2809 (I50285,I2507,I50149,I50117,);
nand I_2810 (I50316,I50260,I306070);
nand I_2811 (I50333,I50183,I50316);
not I_2812 (I50129,I50333);
DFFARX1 I_2813 (I306073,I2507,I50149,I50373,);
DFFARX1 I_2814 (I50373,I2507,I50149,I50138,);
nand I_2815 (I50395,I306052,I306064);
and I_2816 (I50412,I50395,I306058);
DFFARX1 I_2817 (I50412,I2507,I50149,I50438,);
DFFARX1 I_2818 (I50438,I2507,I50149,I50455,);
not I_2819 (I50141,I50455);
not I_2820 (I50477,I50438);
nand I_2821 (I50126,I50477,I50316);
nor I_2822 (I50508,I306067,I306064);
not I_2823 (I50525,I50508);
nor I_2824 (I50542,I50477,I50525);
nor I_2825 (I50559,I50183,I50542);
DFFARX1 I_2826 (I50559,I2507,I50149,I50135,);
nor I_2827 (I50590,I50243,I50525);
nor I_2828 (I50123,I50438,I50590);
nor I_2829 (I50132,I50373,I50508);
nor I_2830 (I50120,I50243,I50508);
not I_2831 (I50676,I2514);
DFFARX1 I_2832 (I1286565,I2507,I50676,I50702,);
not I_2833 (I50710,I50702);
nand I_2834 (I50727,I1286568,I1286562);
and I_2835 (I50744,I50727,I1286559);
DFFARX1 I_2836 (I50744,I2507,I50676,I50770,);
DFFARX1 I_2837 (I1286544,I2507,I50676,I50787,);
and I_2838 (I50795,I50787,I1286553);
nor I_2839 (I50812,I50770,I50795);
DFFARX1 I_2840 (I50812,I2507,I50676,I50644,);
nand I_2841 (I50843,I50787,I1286553);
nand I_2842 (I50860,I50710,I50843);
not I_2843 (I50656,I50860);
DFFARX1 I_2844 (I1286544,I2507,I50676,I50900,);
DFFARX1 I_2845 (I50900,I2507,I50676,I50665,);
nand I_2846 (I50922,I1286547,I1286550);
and I_2847 (I50939,I50922,I1286556);
DFFARX1 I_2848 (I50939,I2507,I50676,I50965,);
DFFARX1 I_2849 (I50965,I2507,I50676,I50982,);
not I_2850 (I50668,I50982);
not I_2851 (I51004,I50965);
nand I_2852 (I50653,I51004,I50843);
nor I_2853 (I51035,I1286547,I1286550);
not I_2854 (I51052,I51035);
nor I_2855 (I51069,I51004,I51052);
nor I_2856 (I51086,I50710,I51069);
DFFARX1 I_2857 (I51086,I2507,I50676,I50662,);
nor I_2858 (I51117,I50770,I51052);
nor I_2859 (I50650,I50965,I51117);
nor I_2860 (I50659,I50900,I51035);
nor I_2861 (I50647,I50770,I51035);
not I_2862 (I51203,I2514);
DFFARX1 I_2863 (I1141030,I2507,I51203,I51229,);
not I_2864 (I51237,I51229);
nand I_2865 (I51254,I1141045,I1141024);
and I_2866 (I51271,I51254,I1141027);
DFFARX1 I_2867 (I51271,I2507,I51203,I51297,);
DFFARX1 I_2868 (I1141048,I2507,I51203,I51314,);
and I_2869 (I51322,I51314,I1141027);
nor I_2870 (I51339,I51297,I51322);
DFFARX1 I_2871 (I51339,I2507,I51203,I51171,);
nand I_2872 (I51370,I51314,I1141027);
nand I_2873 (I51387,I51237,I51370);
not I_2874 (I51183,I51387);
DFFARX1 I_2875 (I1141024,I2507,I51203,I51427,);
DFFARX1 I_2876 (I51427,I2507,I51203,I51192,);
nand I_2877 (I51449,I1141036,I1141033);
and I_2878 (I51466,I51449,I1141039);
DFFARX1 I_2879 (I51466,I2507,I51203,I51492,);
DFFARX1 I_2880 (I51492,I2507,I51203,I51509,);
not I_2881 (I51195,I51509);
not I_2882 (I51531,I51492);
nand I_2883 (I51180,I51531,I51370);
nor I_2884 (I51562,I1141042,I1141033);
not I_2885 (I51579,I51562);
nor I_2886 (I51596,I51531,I51579);
nor I_2887 (I51613,I51237,I51596);
DFFARX1 I_2888 (I51613,I2507,I51203,I51189,);
nor I_2889 (I51644,I51297,I51579);
nor I_2890 (I51177,I51492,I51644);
nor I_2891 (I51186,I51427,I51562);
nor I_2892 (I51174,I51297,I51562);
not I_2893 (I51730,I2514);
DFFARX1 I_2894 (I1118488,I2507,I51730,I51756,);
not I_2895 (I51764,I51756);
nand I_2896 (I51781,I1118503,I1118482);
and I_2897 (I51798,I51781,I1118485);
DFFARX1 I_2898 (I51798,I2507,I51730,I51824,);
DFFARX1 I_2899 (I1118506,I2507,I51730,I51841,);
and I_2900 (I51849,I51841,I1118485);
nor I_2901 (I51866,I51824,I51849);
DFFARX1 I_2902 (I51866,I2507,I51730,I51698,);
nand I_2903 (I51897,I51841,I1118485);
nand I_2904 (I51914,I51764,I51897);
not I_2905 (I51710,I51914);
DFFARX1 I_2906 (I1118482,I2507,I51730,I51954,);
DFFARX1 I_2907 (I51954,I2507,I51730,I51719,);
nand I_2908 (I51976,I1118494,I1118491);
and I_2909 (I51993,I51976,I1118497);
DFFARX1 I_2910 (I51993,I2507,I51730,I52019,);
DFFARX1 I_2911 (I52019,I2507,I51730,I52036,);
not I_2912 (I51722,I52036);
not I_2913 (I52058,I52019);
nand I_2914 (I51707,I52058,I51897);
nor I_2915 (I52089,I1118500,I1118491);
not I_2916 (I52106,I52089);
nor I_2917 (I52123,I52058,I52106);
nor I_2918 (I52140,I51764,I52123);
DFFARX1 I_2919 (I52140,I2507,I51730,I51716,);
nor I_2920 (I52171,I51824,I52106);
nor I_2921 (I51704,I52019,I52171);
nor I_2922 (I51713,I51954,I52089);
nor I_2923 (I51701,I51824,I52089);
not I_2924 (I52257,I2514);
DFFARX1 I_2925 (I991586,I2507,I52257,I52283,);
not I_2926 (I52291,I52283);
nand I_2927 (I52308,I991604,I991598);
and I_2928 (I52325,I52308,I991577);
DFFARX1 I_2929 (I52325,I2507,I52257,I52351,);
DFFARX1 I_2930 (I991595,I2507,I52257,I52368,);
and I_2931 (I52376,I52368,I991580);
nor I_2932 (I52393,I52351,I52376);
DFFARX1 I_2933 (I52393,I2507,I52257,I52225,);
nand I_2934 (I52424,I52368,I991580);
nand I_2935 (I52441,I52291,I52424);
not I_2936 (I52237,I52441);
DFFARX1 I_2937 (I991592,I2507,I52257,I52481,);
DFFARX1 I_2938 (I52481,I2507,I52257,I52246,);
nand I_2939 (I52503,I991601,I991589);
and I_2940 (I52520,I52503,I991583);
DFFARX1 I_2941 (I52520,I2507,I52257,I52546,);
DFFARX1 I_2942 (I52546,I2507,I52257,I52563,);
not I_2943 (I52249,I52563);
not I_2944 (I52585,I52546);
nand I_2945 (I52234,I52585,I52424);
nor I_2946 (I52616,I991577,I991589);
not I_2947 (I52633,I52616);
nor I_2948 (I52650,I52585,I52633);
nor I_2949 (I52667,I52291,I52650);
DFFARX1 I_2950 (I52667,I2507,I52257,I52243,);
nor I_2951 (I52698,I52351,I52633);
nor I_2952 (I52231,I52546,I52698);
nor I_2953 (I52240,I52481,I52616);
nor I_2954 (I52228,I52351,I52616);
not I_2955 (I52784,I2514);
DFFARX1 I_2956 (I1327934,I2507,I52784,I52810,);
not I_2957 (I52818,I52810);
nand I_2958 (I52835,I1327928,I1327949);
and I_2959 (I52852,I52835,I1327925);
DFFARX1 I_2960 (I52852,I2507,I52784,I52878,);
DFFARX1 I_2961 (I1327946,I2507,I52784,I52895,);
and I_2962 (I52903,I52895,I1327943);
nor I_2963 (I52920,I52878,I52903);
DFFARX1 I_2964 (I52920,I2507,I52784,I52752,);
nand I_2965 (I52951,I52895,I1327943);
nand I_2966 (I52968,I52818,I52951);
not I_2967 (I52764,I52968);
DFFARX1 I_2968 (I1327931,I2507,I52784,I53008,);
DFFARX1 I_2969 (I53008,I2507,I52784,I52773,);
nand I_2970 (I53030,I1327940,I1327937);
and I_2971 (I53047,I53030,I1327922);
DFFARX1 I_2972 (I53047,I2507,I52784,I53073,);
DFFARX1 I_2973 (I53073,I2507,I52784,I53090,);
not I_2974 (I52776,I53090);
not I_2975 (I53112,I53073);
nand I_2976 (I52761,I53112,I52951);
nor I_2977 (I53143,I1327922,I1327937);
not I_2978 (I53160,I53143);
nor I_2979 (I53177,I53112,I53160);
nor I_2980 (I53194,I52818,I53177);
DFFARX1 I_2981 (I53194,I2507,I52784,I52770,);
nor I_2982 (I53225,I52878,I53160);
nor I_2983 (I52758,I53073,I53225);
nor I_2984 (I52767,I53008,I53143);
nor I_2985 (I52755,I52878,I53143);
not I_2986 (I53311,I2514);
DFFARX1 I_2987 (I44344,I2507,I53311,I53337,);
not I_2988 (I53345,I53337);
nand I_2989 (I53362,I44332,I44338);
and I_2990 (I53379,I53362,I44341);
DFFARX1 I_2991 (I53379,I2507,I53311,I53405,);
DFFARX1 I_2992 (I44323,I2507,I53311,I53422,);
and I_2993 (I53430,I53422,I44329);
nor I_2994 (I53447,I53405,I53430);
DFFARX1 I_2995 (I53447,I2507,I53311,I53279,);
nand I_2996 (I53478,I53422,I44329);
nand I_2997 (I53495,I53345,I53478);
not I_2998 (I53291,I53495);
DFFARX1 I_2999 (I44323,I2507,I53311,I53535,);
DFFARX1 I_3000 (I53535,I2507,I53311,I53300,);
nand I_3001 (I53557,I44326,I44320);
and I_3002 (I53574,I53557,I44335);
DFFARX1 I_3003 (I53574,I2507,I53311,I53600,);
DFFARX1 I_3004 (I53600,I2507,I53311,I53617,);
not I_3005 (I53303,I53617);
not I_3006 (I53639,I53600);
nand I_3007 (I53288,I53639,I53478);
nor I_3008 (I53670,I44320,I44320);
not I_3009 (I53687,I53670);
nor I_3010 (I53704,I53639,I53687);
nor I_3011 (I53721,I53345,I53704);
DFFARX1 I_3012 (I53721,I2507,I53311,I53297,);
nor I_3013 (I53752,I53405,I53687);
nor I_3014 (I53285,I53600,I53752);
nor I_3015 (I53294,I53535,I53670);
nor I_3016 (I53282,I53405,I53670);
not I_3017 (I53838,I2514);
DFFARX1 I_3018 (I1030901,I2507,I53838,I53864,);
not I_3019 (I53872,I53864);
nand I_3020 (I53889,I1030898,I1030904);
and I_3021 (I53906,I53889,I1030901);
DFFARX1 I_3022 (I53906,I2507,I53838,I53932,);
DFFARX1 I_3023 (I1030904,I2507,I53838,I53949,);
and I_3024 (I53957,I53949,I1030898);
nor I_3025 (I53974,I53932,I53957);
DFFARX1 I_3026 (I53974,I2507,I53838,I53806,);
nand I_3027 (I54005,I53949,I1030898);
nand I_3028 (I54022,I53872,I54005);
not I_3029 (I53818,I54022);
DFFARX1 I_3030 (I1030907,I2507,I53838,I54062,);
DFFARX1 I_3031 (I54062,I2507,I53838,I53827,);
nand I_3032 (I54084,I1030910,I1030919);
and I_3033 (I54101,I54084,I1030913);
DFFARX1 I_3034 (I54101,I2507,I53838,I54127,);
DFFARX1 I_3035 (I54127,I2507,I53838,I54144,);
not I_3036 (I53830,I54144);
not I_3037 (I54166,I54127);
nand I_3038 (I53815,I54166,I54005);
nor I_3039 (I54197,I1030916,I1030919);
not I_3040 (I54214,I54197);
nor I_3041 (I54231,I54166,I54214);
nor I_3042 (I54248,I53872,I54231);
DFFARX1 I_3043 (I54248,I2507,I53838,I53824,);
nor I_3044 (I54279,I53932,I54214);
nor I_3045 (I53812,I54127,I54279);
nor I_3046 (I53821,I54062,I54197);
nor I_3047 (I53809,I53932,I54197);
not I_3048 (I54365,I2514);
DFFARX1 I_3049 (I669456,I2507,I54365,I54391,);
not I_3050 (I54399,I54391);
nand I_3051 (I54416,I669447,I669465);
and I_3052 (I54433,I54416,I669444);
DFFARX1 I_3053 (I54433,I2507,I54365,I54459,);
DFFARX1 I_3054 (I669447,I2507,I54365,I54476,);
and I_3055 (I54484,I54476,I669450);
nor I_3056 (I54501,I54459,I54484);
DFFARX1 I_3057 (I54501,I2507,I54365,I54333,);
nand I_3058 (I54532,I54476,I669450);
nand I_3059 (I54549,I54399,I54532);
not I_3060 (I54345,I54549);
DFFARX1 I_3061 (I669444,I2507,I54365,I54589,);
DFFARX1 I_3062 (I54589,I2507,I54365,I54354,);
nand I_3063 (I54611,I669462,I669453);
and I_3064 (I54628,I54611,I669468);
DFFARX1 I_3065 (I54628,I2507,I54365,I54654,);
DFFARX1 I_3066 (I54654,I2507,I54365,I54671,);
not I_3067 (I54357,I54671);
not I_3068 (I54693,I54654);
nand I_3069 (I54342,I54693,I54532);
nor I_3070 (I54724,I669459,I669453);
not I_3071 (I54741,I54724);
nor I_3072 (I54758,I54693,I54741);
nor I_3073 (I54775,I54399,I54758);
DFFARX1 I_3074 (I54775,I2507,I54365,I54351,);
nor I_3075 (I54806,I54459,I54741);
nor I_3076 (I54339,I54654,I54806);
nor I_3077 (I54348,I54589,I54724);
nor I_3078 (I54336,I54459,I54724);
not I_3079 (I54892,I2514);
DFFARX1 I_3080 (I883942,I2507,I54892,I54918,);
not I_3081 (I54926,I54918);
nand I_3082 (I54943,I883939,I883954);
and I_3083 (I54960,I54943,I883936);
DFFARX1 I_3084 (I54960,I2507,I54892,I54986,);
DFFARX1 I_3085 (I883933,I2507,I54892,I55003,);
and I_3086 (I55011,I55003,I883933);
nor I_3087 (I55028,I54986,I55011);
DFFARX1 I_3088 (I55028,I2507,I54892,I54860,);
nand I_3089 (I55059,I55003,I883933);
nand I_3090 (I55076,I54926,I55059);
not I_3091 (I54872,I55076);
DFFARX1 I_3092 (I883936,I2507,I54892,I55116,);
DFFARX1 I_3093 (I55116,I2507,I54892,I54881,);
nand I_3094 (I55138,I883948,I883939);
and I_3095 (I55155,I55138,I883951);
DFFARX1 I_3096 (I55155,I2507,I54892,I55181,);
DFFARX1 I_3097 (I55181,I2507,I54892,I55198,);
not I_3098 (I54884,I55198);
not I_3099 (I55220,I55181);
nand I_3100 (I54869,I55220,I55059);
nor I_3101 (I55251,I883945,I883939);
not I_3102 (I55268,I55251);
nor I_3103 (I55285,I55220,I55268);
nor I_3104 (I55302,I54926,I55285);
DFFARX1 I_3105 (I55302,I2507,I54892,I54878,);
nor I_3106 (I55333,I54986,I55268);
nor I_3107 (I54866,I55181,I55333);
nor I_3108 (I54875,I55116,I55251);
nor I_3109 (I54863,I54986,I55251);
not I_3110 (I55419,I2514);
DFFARX1 I_3111 (I536337,I2507,I55419,I55445,);
not I_3112 (I55453,I55445);
nand I_3113 (I55470,I536358,I536352);
and I_3114 (I55487,I55470,I536334);
DFFARX1 I_3115 (I55487,I2507,I55419,I55513,);
DFFARX1 I_3116 (I536337,I2507,I55419,I55530,);
and I_3117 (I55538,I55530,I536346);
nor I_3118 (I55555,I55513,I55538);
DFFARX1 I_3119 (I55555,I2507,I55419,I55387,);
nand I_3120 (I55586,I55530,I536346);
nand I_3121 (I55603,I55453,I55586);
not I_3122 (I55399,I55603);
DFFARX1 I_3123 (I536343,I2507,I55419,I55643,);
DFFARX1 I_3124 (I55643,I2507,I55419,I55408,);
nand I_3125 (I55665,I536349,I536340);
and I_3126 (I55682,I55665,I536334);
DFFARX1 I_3127 (I55682,I2507,I55419,I55708,);
DFFARX1 I_3128 (I55708,I2507,I55419,I55725,);
not I_3129 (I55411,I55725);
not I_3130 (I55747,I55708);
nand I_3131 (I55396,I55747,I55586);
nor I_3132 (I55778,I536355,I536340);
not I_3133 (I55795,I55778);
nor I_3134 (I55812,I55747,I55795);
nor I_3135 (I55829,I55453,I55812);
DFFARX1 I_3136 (I55829,I2507,I55419,I55405,);
nor I_3137 (I55860,I55513,I55795);
nor I_3138 (I55393,I55708,I55860);
nor I_3139 (I55402,I55643,I55778);
nor I_3140 (I55390,I55513,I55778);
not I_3141 (I55946,I2514);
DFFARX1 I_3142 (I219262,I2507,I55946,I55972,);
not I_3143 (I55980,I55972);
nand I_3144 (I55997,I219256,I219250);
and I_3145 (I56014,I55997,I219271);
DFFARX1 I_3146 (I56014,I2507,I55946,I56040,);
DFFARX1 I_3147 (I219268,I2507,I55946,I56057,);
and I_3148 (I56065,I56057,I219265);
nor I_3149 (I56082,I56040,I56065);
DFFARX1 I_3150 (I56082,I2507,I55946,I55914,);
nand I_3151 (I56113,I56057,I219265);
nand I_3152 (I56130,I55980,I56113);
not I_3153 (I55926,I56130);
DFFARX1 I_3154 (I219250,I2507,I55946,I56170,);
DFFARX1 I_3155 (I56170,I2507,I55946,I55935,);
nand I_3156 (I56192,I219253,I219253);
and I_3157 (I56209,I56192,I219274);
DFFARX1 I_3158 (I56209,I2507,I55946,I56235,);
DFFARX1 I_3159 (I56235,I2507,I55946,I56252,);
not I_3160 (I55938,I56252);
not I_3161 (I56274,I56235);
nand I_3162 (I55923,I56274,I56113);
nor I_3163 (I56305,I219259,I219253);
not I_3164 (I56322,I56305);
nor I_3165 (I56339,I56274,I56322);
nor I_3166 (I56356,I55980,I56339);
DFFARX1 I_3167 (I56356,I2507,I55946,I55932,);
nor I_3168 (I56387,I56040,I56322);
nor I_3169 (I55920,I56235,I56387);
nor I_3170 (I55929,I56170,I56305);
nor I_3171 (I55917,I56040,I56305);
not I_3172 (I56473,I2514);
DFFARX1 I_3173 (I819121,I2507,I56473,I56499,);
not I_3174 (I56507,I56499);
nand I_3175 (I56524,I819118,I819133);
and I_3176 (I56541,I56524,I819115);
DFFARX1 I_3177 (I56541,I2507,I56473,I56567,);
DFFARX1 I_3178 (I819112,I2507,I56473,I56584,);
and I_3179 (I56592,I56584,I819112);
nor I_3180 (I56609,I56567,I56592);
DFFARX1 I_3181 (I56609,I2507,I56473,I56441,);
nand I_3182 (I56640,I56584,I819112);
nand I_3183 (I56657,I56507,I56640);
not I_3184 (I56453,I56657);
DFFARX1 I_3185 (I819115,I2507,I56473,I56697,);
DFFARX1 I_3186 (I56697,I2507,I56473,I56462,);
nand I_3187 (I56719,I819127,I819118);
and I_3188 (I56736,I56719,I819130);
DFFARX1 I_3189 (I56736,I2507,I56473,I56762,);
DFFARX1 I_3190 (I56762,I2507,I56473,I56779,);
not I_3191 (I56465,I56779);
not I_3192 (I56801,I56762);
nand I_3193 (I56450,I56801,I56640);
nor I_3194 (I56832,I819124,I819118);
not I_3195 (I56849,I56832);
nor I_3196 (I56866,I56801,I56849);
nor I_3197 (I56883,I56507,I56866);
DFFARX1 I_3198 (I56883,I2507,I56473,I56459,);
nor I_3199 (I56914,I56567,I56849);
nor I_3200 (I56447,I56762,I56914);
nor I_3201 (I56456,I56697,I56832);
nor I_3202 (I56444,I56567,I56832);
not I_3203 (I57000,I2514);
DFFARX1 I_3204 (I713384,I2507,I57000,I57026,);
not I_3205 (I57034,I57026);
nand I_3206 (I57051,I713375,I713393);
and I_3207 (I57068,I57051,I713372);
DFFARX1 I_3208 (I57068,I2507,I57000,I57094,);
DFFARX1 I_3209 (I713375,I2507,I57000,I57111,);
and I_3210 (I57119,I57111,I713378);
nor I_3211 (I57136,I57094,I57119);
DFFARX1 I_3212 (I57136,I2507,I57000,I56968,);
nand I_3213 (I57167,I57111,I713378);
nand I_3214 (I57184,I57034,I57167);
not I_3215 (I56980,I57184);
DFFARX1 I_3216 (I713372,I2507,I57000,I57224,);
DFFARX1 I_3217 (I57224,I2507,I57000,I56989,);
nand I_3218 (I57246,I713390,I713381);
and I_3219 (I57263,I57246,I713396);
DFFARX1 I_3220 (I57263,I2507,I57000,I57289,);
DFFARX1 I_3221 (I57289,I2507,I57000,I57306,);
not I_3222 (I56992,I57306);
not I_3223 (I57328,I57289);
nand I_3224 (I56977,I57328,I57167);
nor I_3225 (I57359,I713387,I713381);
not I_3226 (I57376,I57359);
nor I_3227 (I57393,I57328,I57376);
nor I_3228 (I57410,I57034,I57393);
DFFARX1 I_3229 (I57410,I2507,I57000,I56986,);
nor I_3230 (I57441,I57094,I57376);
nor I_3231 (I56974,I57289,I57441);
nor I_3232 (I56983,I57224,I57359);
nor I_3233 (I56971,I57094,I57359);
not I_3234 (I57527,I2514);
DFFARX1 I_3235 (I832296,I2507,I57527,I57553,);
not I_3236 (I57561,I57553);
nand I_3237 (I57578,I832293,I832308);
and I_3238 (I57595,I57578,I832290);
DFFARX1 I_3239 (I57595,I2507,I57527,I57621,);
DFFARX1 I_3240 (I832287,I2507,I57527,I57638,);
and I_3241 (I57646,I57638,I832287);
nor I_3242 (I57663,I57621,I57646);
DFFARX1 I_3243 (I57663,I2507,I57527,I57495,);
nand I_3244 (I57694,I57638,I832287);
nand I_3245 (I57711,I57561,I57694);
not I_3246 (I57507,I57711);
DFFARX1 I_3247 (I832290,I2507,I57527,I57751,);
DFFARX1 I_3248 (I57751,I2507,I57527,I57516,);
nand I_3249 (I57773,I832302,I832293);
and I_3250 (I57790,I57773,I832305);
DFFARX1 I_3251 (I57790,I2507,I57527,I57816,);
DFFARX1 I_3252 (I57816,I2507,I57527,I57833,);
not I_3253 (I57519,I57833);
not I_3254 (I57855,I57816);
nand I_3255 (I57504,I57855,I57694);
nor I_3256 (I57886,I832299,I832293);
not I_3257 (I57903,I57886);
nor I_3258 (I57920,I57855,I57903);
nor I_3259 (I57937,I57561,I57920);
DFFARX1 I_3260 (I57937,I2507,I57527,I57513,);
nor I_3261 (I57968,I57621,I57903);
nor I_3262 (I57501,I57816,I57968);
nor I_3263 (I57510,I57751,I57886);
nor I_3264 (I57498,I57621,I57886);
not I_3265 (I58054,I2514);
DFFARX1 I_3266 (I457761,I2507,I58054,I58080,);
not I_3267 (I58088,I58080);
nand I_3268 (I58105,I457755,I457746);
and I_3269 (I58122,I58105,I457767);
DFFARX1 I_3270 (I58122,I2507,I58054,I58148,);
DFFARX1 I_3271 (I457749,I2507,I58054,I58165,);
and I_3272 (I58173,I58165,I457743);
nor I_3273 (I58190,I58148,I58173);
DFFARX1 I_3274 (I58190,I2507,I58054,I58022,);
nand I_3275 (I58221,I58165,I457743);
nand I_3276 (I58238,I58088,I58221);
not I_3277 (I58034,I58238);
DFFARX1 I_3278 (I457743,I2507,I58054,I58278,);
DFFARX1 I_3279 (I58278,I2507,I58054,I58043,);
nand I_3280 (I58300,I457770,I457752);
and I_3281 (I58317,I58300,I457758);
DFFARX1 I_3282 (I58317,I2507,I58054,I58343,);
DFFARX1 I_3283 (I58343,I2507,I58054,I58360,);
not I_3284 (I58046,I58360);
not I_3285 (I58382,I58343);
nand I_3286 (I58031,I58382,I58221);
nor I_3287 (I58413,I457764,I457752);
not I_3288 (I58430,I58413);
nor I_3289 (I58447,I58382,I58430);
nor I_3290 (I58464,I58088,I58447);
DFFARX1 I_3291 (I58464,I2507,I58054,I58040,);
nor I_3292 (I58495,I58148,I58430);
nor I_3293 (I58028,I58343,I58495);
nor I_3294 (I58037,I58278,I58413);
nor I_3295 (I58025,I58148,I58413);
not I_3296 (I58581,I2514);
DFFARX1 I_3297 (I846525,I2507,I58581,I58607,);
not I_3298 (I58615,I58607);
nand I_3299 (I58632,I846522,I846537);
and I_3300 (I58649,I58632,I846519);
DFFARX1 I_3301 (I58649,I2507,I58581,I58675,);
DFFARX1 I_3302 (I846516,I2507,I58581,I58692,);
and I_3303 (I58700,I58692,I846516);
nor I_3304 (I58717,I58675,I58700);
DFFARX1 I_3305 (I58717,I2507,I58581,I58549,);
nand I_3306 (I58748,I58692,I846516);
nand I_3307 (I58765,I58615,I58748);
not I_3308 (I58561,I58765);
DFFARX1 I_3309 (I846519,I2507,I58581,I58805,);
DFFARX1 I_3310 (I58805,I2507,I58581,I58570,);
nand I_3311 (I58827,I846531,I846522);
and I_3312 (I58844,I58827,I846534);
DFFARX1 I_3313 (I58844,I2507,I58581,I58870,);
DFFARX1 I_3314 (I58870,I2507,I58581,I58887,);
not I_3315 (I58573,I58887);
not I_3316 (I58909,I58870);
nand I_3317 (I58558,I58909,I58748);
nor I_3318 (I58940,I846528,I846522);
not I_3319 (I58957,I58940);
nor I_3320 (I58974,I58909,I58957);
nor I_3321 (I58991,I58615,I58974);
DFFARX1 I_3322 (I58991,I2507,I58581,I58567,);
nor I_3323 (I59022,I58675,I58957);
nor I_3324 (I58555,I58870,I59022);
nor I_3325 (I58564,I58805,I58940);
nor I_3326 (I58552,I58675,I58940);
not I_3327 (I59108,I2514);
DFFARX1 I_3328 (I877091,I2507,I59108,I59134,);
not I_3329 (I59142,I59134);
nand I_3330 (I59159,I877088,I877103);
and I_3331 (I59176,I59159,I877085);
DFFARX1 I_3332 (I59176,I2507,I59108,I59202,);
DFFARX1 I_3333 (I877082,I2507,I59108,I59219,);
and I_3334 (I59227,I59219,I877082);
nor I_3335 (I59244,I59202,I59227);
DFFARX1 I_3336 (I59244,I2507,I59108,I59076,);
nand I_3337 (I59275,I59219,I877082);
nand I_3338 (I59292,I59142,I59275);
not I_3339 (I59088,I59292);
DFFARX1 I_3340 (I877085,I2507,I59108,I59332,);
DFFARX1 I_3341 (I59332,I2507,I59108,I59097,);
nand I_3342 (I59354,I877097,I877088);
and I_3343 (I59371,I59354,I877100);
DFFARX1 I_3344 (I59371,I2507,I59108,I59397,);
DFFARX1 I_3345 (I59397,I2507,I59108,I59414,);
not I_3346 (I59100,I59414);
not I_3347 (I59436,I59397);
nand I_3348 (I59085,I59436,I59275);
nor I_3349 (I59467,I877094,I877088);
not I_3350 (I59484,I59467);
nor I_3351 (I59501,I59436,I59484);
nor I_3352 (I59518,I59142,I59501);
DFFARX1 I_3353 (I59518,I2507,I59108,I59094,);
nor I_3354 (I59549,I59202,I59484);
nor I_3355 (I59082,I59397,I59549);
nor I_3356 (I59091,I59332,I59467);
nor I_3357 (I59079,I59202,I59467);
not I_3358 (I59635,I2514);
DFFARX1 I_3359 (I360887,I2507,I59635,I59661,);
not I_3360 (I59669,I59661);
nand I_3361 (I59686,I360869,I360884);
and I_3362 (I59703,I59686,I360860);
DFFARX1 I_3363 (I59703,I2507,I59635,I59729,);
DFFARX1 I_3364 (I360863,I2507,I59635,I59746,);
and I_3365 (I59754,I59746,I360878);
nor I_3366 (I59771,I59729,I59754);
DFFARX1 I_3367 (I59771,I2507,I59635,I59603,);
nand I_3368 (I59802,I59746,I360878);
nand I_3369 (I59819,I59669,I59802);
not I_3370 (I59615,I59819);
DFFARX1 I_3371 (I360881,I2507,I59635,I59859,);
DFFARX1 I_3372 (I59859,I2507,I59635,I59624,);
nand I_3373 (I59881,I360860,I360872);
and I_3374 (I59898,I59881,I360866);
DFFARX1 I_3375 (I59898,I2507,I59635,I59924,);
DFFARX1 I_3376 (I59924,I2507,I59635,I59941,);
not I_3377 (I59627,I59941);
not I_3378 (I59963,I59924);
nand I_3379 (I59612,I59963,I59802);
nor I_3380 (I59994,I360875,I360872);
not I_3381 (I60011,I59994);
nor I_3382 (I60028,I59963,I60011);
nor I_3383 (I60045,I59669,I60028);
DFFARX1 I_3384 (I60045,I2507,I59635,I59621,);
nor I_3385 (I60076,I59729,I60011);
nor I_3386 (I59609,I59924,I60076);
nor I_3387 (I59618,I59859,I59994);
nor I_3388 (I59606,I59729,I59994);
not I_3389 (I60162,I2514);
DFFARX1 I_3390 (I592001,I2507,I60162,I60188,);
not I_3391 (I60196,I60188);
nand I_3392 (I60213,I592013,I591998);
and I_3393 (I60230,I60213,I591992);
DFFARX1 I_3394 (I60230,I2507,I60162,I60256,);
DFFARX1 I_3395 (I592007,I2507,I60162,I60273,);
and I_3396 (I60281,I60273,I591995);
nor I_3397 (I60298,I60256,I60281);
DFFARX1 I_3398 (I60298,I2507,I60162,I60130,);
nand I_3399 (I60329,I60273,I591995);
nand I_3400 (I60346,I60196,I60329);
not I_3401 (I60142,I60346);
DFFARX1 I_3402 (I592004,I2507,I60162,I60386,);
DFFARX1 I_3403 (I60386,I2507,I60162,I60151,);
nand I_3404 (I60408,I592010,I592016);
and I_3405 (I60425,I60408,I591992);
DFFARX1 I_3406 (I60425,I2507,I60162,I60451,);
DFFARX1 I_3407 (I60451,I2507,I60162,I60468,);
not I_3408 (I60154,I60468);
not I_3409 (I60490,I60451);
nand I_3410 (I60139,I60490,I60329);
nor I_3411 (I60521,I591995,I592016);
not I_3412 (I60538,I60521);
nor I_3413 (I60555,I60490,I60538);
nor I_3414 (I60572,I60196,I60555);
DFFARX1 I_3415 (I60572,I2507,I60162,I60148,);
nor I_3416 (I60603,I60256,I60538);
nor I_3417 (I60136,I60451,I60603);
nor I_3418 (I60145,I60386,I60521);
nor I_3419 (I60133,I60256,I60521);
not I_3420 (I60689,I2514);
DFFARX1 I_3421 (I339807,I2507,I60689,I60715,);
not I_3422 (I60723,I60715);
nand I_3423 (I60740,I339789,I339804);
and I_3424 (I60757,I60740,I339780);
DFFARX1 I_3425 (I60757,I2507,I60689,I60783,);
DFFARX1 I_3426 (I339783,I2507,I60689,I60800,);
and I_3427 (I60808,I60800,I339798);
nor I_3428 (I60825,I60783,I60808);
DFFARX1 I_3429 (I60825,I2507,I60689,I60657,);
nand I_3430 (I60856,I60800,I339798);
nand I_3431 (I60873,I60723,I60856);
not I_3432 (I60669,I60873);
DFFARX1 I_3433 (I339801,I2507,I60689,I60913,);
DFFARX1 I_3434 (I60913,I2507,I60689,I60678,);
nand I_3435 (I60935,I339780,I339792);
and I_3436 (I60952,I60935,I339786);
DFFARX1 I_3437 (I60952,I2507,I60689,I60978,);
DFFARX1 I_3438 (I60978,I2507,I60689,I60995,);
not I_3439 (I60681,I60995);
not I_3440 (I61017,I60978);
nand I_3441 (I60666,I61017,I60856);
nor I_3442 (I61048,I339795,I339792);
not I_3443 (I61065,I61048);
nor I_3444 (I61082,I61017,I61065);
nor I_3445 (I61099,I60723,I61082);
DFFARX1 I_3446 (I61099,I2507,I60689,I60675,);
nor I_3447 (I61130,I60783,I61065);
nor I_3448 (I60663,I60978,I61130);
nor I_3449 (I60672,I60913,I61048);
nor I_3450 (I60660,I60783,I61048);
not I_3451 (I61216,I2514);
DFFARX1 I_3452 (I12647,I2507,I61216,I61242,);
not I_3453 (I61250,I61242);
nand I_3454 (I61267,I12632,I12632);
and I_3455 (I61284,I61267,I12653);
DFFARX1 I_3456 (I61284,I2507,I61216,I61310,);
DFFARX1 I_3457 (I12635,I2507,I61216,I61327,);
and I_3458 (I61335,I61327,I12644);
nor I_3459 (I61352,I61310,I61335);
DFFARX1 I_3460 (I61352,I2507,I61216,I61184,);
nand I_3461 (I61383,I61327,I12644);
nand I_3462 (I61400,I61250,I61383);
not I_3463 (I61196,I61400);
DFFARX1 I_3464 (I12638,I2507,I61216,I61440,);
DFFARX1 I_3465 (I61440,I2507,I61216,I61205,);
nand I_3466 (I61462,I12641,I12650);
and I_3467 (I61479,I61462,I12635);
DFFARX1 I_3468 (I61479,I2507,I61216,I61505,);
DFFARX1 I_3469 (I61505,I2507,I61216,I61522,);
not I_3470 (I61208,I61522);
not I_3471 (I61544,I61505);
nand I_3472 (I61193,I61544,I61383);
nor I_3473 (I61575,I12638,I12650);
not I_3474 (I61592,I61575);
nor I_3475 (I61609,I61544,I61592);
nor I_3476 (I61626,I61250,I61609);
DFFARX1 I_3477 (I61626,I2507,I61216,I61202,);
nor I_3478 (I61657,I61310,I61592);
nor I_3479 (I61190,I61505,I61657);
nor I_3480 (I61199,I61440,I61575);
nor I_3481 (I61187,I61310,I61575);
not I_3482 (I61743,I2514);
DFFARX1 I_3483 (I715118,I2507,I61743,I61769,);
not I_3484 (I61777,I61769);
nand I_3485 (I61794,I715109,I715127);
and I_3486 (I61811,I61794,I715106);
DFFARX1 I_3487 (I61811,I2507,I61743,I61837,);
DFFARX1 I_3488 (I715109,I2507,I61743,I61854,);
and I_3489 (I61862,I61854,I715112);
nor I_3490 (I61879,I61837,I61862);
DFFARX1 I_3491 (I61879,I2507,I61743,I61711,);
nand I_3492 (I61910,I61854,I715112);
nand I_3493 (I61927,I61777,I61910);
not I_3494 (I61723,I61927);
DFFARX1 I_3495 (I715106,I2507,I61743,I61967,);
DFFARX1 I_3496 (I61967,I2507,I61743,I61732,);
nand I_3497 (I61989,I715124,I715115);
and I_3498 (I62006,I61989,I715130);
DFFARX1 I_3499 (I62006,I2507,I61743,I62032,);
DFFARX1 I_3500 (I62032,I2507,I61743,I62049,);
not I_3501 (I61735,I62049);
not I_3502 (I62071,I62032);
nand I_3503 (I61720,I62071,I61910);
nor I_3504 (I62102,I715121,I715115);
not I_3505 (I62119,I62102);
nor I_3506 (I62136,I62071,I62119);
nor I_3507 (I62153,I61777,I62136);
DFFARX1 I_3508 (I62153,I2507,I61743,I61729,);
nor I_3509 (I62184,I61837,I62119);
nor I_3510 (I61717,I62032,I62184);
nor I_3511 (I61726,I61967,I62102);
nor I_3512 (I61714,I61837,I62102);
not I_3513 (I62270,I2514);
DFFARX1 I_3514 (I196652,I2507,I62270,I62296,);
not I_3515 (I62304,I62296);
nand I_3516 (I62321,I196646,I196640);
and I_3517 (I62338,I62321,I196661);
DFFARX1 I_3518 (I62338,I2507,I62270,I62364,);
DFFARX1 I_3519 (I196658,I2507,I62270,I62381,);
and I_3520 (I62389,I62381,I196655);
nor I_3521 (I62406,I62364,I62389);
DFFARX1 I_3522 (I62406,I2507,I62270,I62238,);
nand I_3523 (I62437,I62381,I196655);
nand I_3524 (I62454,I62304,I62437);
not I_3525 (I62250,I62454);
DFFARX1 I_3526 (I196640,I2507,I62270,I62494,);
DFFARX1 I_3527 (I62494,I2507,I62270,I62259,);
nand I_3528 (I62516,I196643,I196643);
and I_3529 (I62533,I62516,I196664);
DFFARX1 I_3530 (I62533,I2507,I62270,I62559,);
DFFARX1 I_3531 (I62559,I2507,I62270,I62576,);
not I_3532 (I62262,I62576);
not I_3533 (I62598,I62559);
nand I_3534 (I62247,I62598,I62437);
nor I_3535 (I62629,I196649,I196643);
not I_3536 (I62646,I62629);
nor I_3537 (I62663,I62598,I62646);
nor I_3538 (I62680,I62304,I62663);
DFFARX1 I_3539 (I62680,I2507,I62270,I62256,);
nor I_3540 (I62711,I62364,I62646);
nor I_3541 (I62244,I62559,I62711);
nor I_3542 (I62253,I62494,I62629);
nor I_3543 (I62241,I62364,I62629);
not I_3544 (I62797,I2514);
DFFARX1 I_3545 (I1253672,I2507,I62797,I62823,);
not I_3546 (I62831,I62823);
nand I_3547 (I62848,I1253666,I1253687);
and I_3548 (I62865,I62848,I1253678);
DFFARX1 I_3549 (I62865,I2507,I62797,I62891,);
DFFARX1 I_3550 (I1253669,I2507,I62797,I62908,);
and I_3551 (I62916,I62908,I1253681);
nor I_3552 (I62933,I62891,I62916);
DFFARX1 I_3553 (I62933,I2507,I62797,I62765,);
nand I_3554 (I62964,I62908,I1253681);
nand I_3555 (I62981,I62831,I62964);
not I_3556 (I62777,I62981);
DFFARX1 I_3557 (I1253669,I2507,I62797,I63021,);
DFFARX1 I_3558 (I63021,I2507,I62797,I62786,);
nand I_3559 (I63043,I1253690,I1253675);
and I_3560 (I63060,I63043,I1253666);
DFFARX1 I_3561 (I63060,I2507,I62797,I63086,);
DFFARX1 I_3562 (I63086,I2507,I62797,I63103,);
not I_3563 (I62789,I63103);
not I_3564 (I63125,I63086);
nand I_3565 (I62774,I63125,I62964);
nor I_3566 (I63156,I1253684,I1253675);
not I_3567 (I63173,I63156);
nor I_3568 (I63190,I63125,I63173);
nor I_3569 (I63207,I62831,I63190);
DFFARX1 I_3570 (I63207,I2507,I62797,I62783,);
nor I_3571 (I63238,I62891,I63173);
nor I_3572 (I62771,I63086,I63238);
nor I_3573 (I62780,I63021,I63156);
nor I_3574 (I62768,I62891,I63156);
not I_3575 (I63324,I2514);
DFFARX1 I_3576 (I209742,I2507,I63324,I63350,);
not I_3577 (I63358,I63350);
nand I_3578 (I63375,I209736,I209730);
and I_3579 (I63392,I63375,I209751);
DFFARX1 I_3580 (I63392,I2507,I63324,I63418,);
DFFARX1 I_3581 (I209748,I2507,I63324,I63435,);
and I_3582 (I63443,I63435,I209745);
nor I_3583 (I63460,I63418,I63443);
DFFARX1 I_3584 (I63460,I2507,I63324,I63292,);
nand I_3585 (I63491,I63435,I209745);
nand I_3586 (I63508,I63358,I63491);
not I_3587 (I63304,I63508);
DFFARX1 I_3588 (I209730,I2507,I63324,I63548,);
DFFARX1 I_3589 (I63548,I2507,I63324,I63313,);
nand I_3590 (I63570,I209733,I209733);
and I_3591 (I63587,I63570,I209754);
DFFARX1 I_3592 (I63587,I2507,I63324,I63613,);
DFFARX1 I_3593 (I63613,I2507,I63324,I63630,);
not I_3594 (I63316,I63630);
not I_3595 (I63652,I63613);
nand I_3596 (I63301,I63652,I63491);
nor I_3597 (I63683,I209739,I209733);
not I_3598 (I63700,I63683);
nor I_3599 (I63717,I63652,I63700);
nor I_3600 (I63734,I63358,I63717);
DFFARX1 I_3601 (I63734,I2507,I63324,I63310,);
nor I_3602 (I63765,I63418,I63700);
nor I_3603 (I63298,I63613,I63765);
nor I_3604 (I63307,I63548,I63683);
nor I_3605 (I63295,I63418,I63683);
not I_3606 (I63851,I2514);
DFFARX1 I_3607 (I479521,I2507,I63851,I63877,);
not I_3608 (I63885,I63877);
nand I_3609 (I63902,I479515,I479506);
and I_3610 (I63919,I63902,I479527);
DFFARX1 I_3611 (I63919,I2507,I63851,I63945,);
DFFARX1 I_3612 (I479509,I2507,I63851,I63962,);
and I_3613 (I63970,I63962,I479503);
nor I_3614 (I63987,I63945,I63970);
DFFARX1 I_3615 (I63987,I2507,I63851,I63819,);
nand I_3616 (I64018,I63962,I479503);
nand I_3617 (I64035,I63885,I64018);
not I_3618 (I63831,I64035);
DFFARX1 I_3619 (I479503,I2507,I63851,I64075,);
DFFARX1 I_3620 (I64075,I2507,I63851,I63840,);
nand I_3621 (I64097,I479530,I479512);
and I_3622 (I64114,I64097,I479518);
DFFARX1 I_3623 (I64114,I2507,I63851,I64140,);
DFFARX1 I_3624 (I64140,I2507,I63851,I64157,);
not I_3625 (I63843,I64157);
not I_3626 (I64179,I64140);
nand I_3627 (I63828,I64179,I64018);
nor I_3628 (I64210,I479524,I479512);
not I_3629 (I64227,I64210);
nor I_3630 (I64244,I64179,I64227);
nor I_3631 (I64261,I63885,I64244);
DFFARX1 I_3632 (I64261,I2507,I63851,I63837,);
nor I_3633 (I64292,I63945,I64227);
nor I_3634 (I63825,I64140,I64292);
nor I_3635 (I63834,I64075,I64210);
nor I_3636 (I63822,I63945,I64210);
not I_3637 (I64378,I2514);
DFFARX1 I_3638 (I268135,I2507,I64378,I64404,);
not I_3639 (I64412,I64404);
nand I_3640 (I64429,I268117,I268132);
and I_3641 (I64446,I64429,I268108);
DFFARX1 I_3642 (I64446,I2507,I64378,I64472,);
DFFARX1 I_3643 (I268111,I2507,I64378,I64489,);
and I_3644 (I64497,I64489,I268126);
nor I_3645 (I64514,I64472,I64497);
DFFARX1 I_3646 (I64514,I2507,I64378,I64346,);
nand I_3647 (I64545,I64489,I268126);
nand I_3648 (I64562,I64412,I64545);
not I_3649 (I64358,I64562);
DFFARX1 I_3650 (I268129,I2507,I64378,I64602,);
DFFARX1 I_3651 (I64602,I2507,I64378,I64367,);
nand I_3652 (I64624,I268108,I268120);
and I_3653 (I64641,I64624,I268114);
DFFARX1 I_3654 (I64641,I2507,I64378,I64667,);
DFFARX1 I_3655 (I64667,I2507,I64378,I64684,);
not I_3656 (I64370,I64684);
not I_3657 (I64706,I64667);
nand I_3658 (I64355,I64706,I64545);
nor I_3659 (I64737,I268123,I268120);
not I_3660 (I64754,I64737);
nor I_3661 (I64771,I64706,I64754);
nor I_3662 (I64788,I64412,I64771);
DFFARX1 I_3663 (I64788,I2507,I64378,I64364,);
nor I_3664 (I64819,I64472,I64754);
nor I_3665 (I64352,I64667,I64819);
nor I_3666 (I64361,I64602,I64737);
nor I_3667 (I64349,I64472,I64737);
not I_3668 (I64905,I2514);
DFFARX1 I_3669 (I143706,I2507,I64905,I64931,);
not I_3670 (I64939,I64931);
nand I_3671 (I64956,I143703,I143685);
and I_3672 (I64973,I64956,I143691);
DFFARX1 I_3673 (I64973,I2507,I64905,I64999,);
DFFARX1 I_3674 (I143700,I2507,I64905,I65016,);
and I_3675 (I65024,I65016,I143694);
nor I_3676 (I65041,I64999,I65024);
DFFARX1 I_3677 (I65041,I2507,I64905,I64873,);
nand I_3678 (I65072,I65016,I143694);
nand I_3679 (I65089,I64939,I65072);
not I_3680 (I64885,I65089);
DFFARX1 I_3681 (I143709,I2507,I64905,I65129,);
DFFARX1 I_3682 (I65129,I2507,I64905,I64894,);
nand I_3683 (I65151,I143697,I143688);
and I_3684 (I65168,I65151,I143685);
DFFARX1 I_3685 (I65168,I2507,I64905,I65194,);
DFFARX1 I_3686 (I65194,I2507,I64905,I65211,);
not I_3687 (I64897,I65211);
not I_3688 (I65233,I65194);
nand I_3689 (I64882,I65233,I65072);
nor I_3690 (I65264,I143712,I143688);
not I_3691 (I65281,I65264);
nor I_3692 (I65298,I65233,I65281);
nor I_3693 (I65315,I64939,I65298);
DFFARX1 I_3694 (I65315,I2507,I64905,I64891,);
nor I_3695 (I65346,I64999,I65281);
nor I_3696 (I64879,I65194,I65346);
nor I_3697 (I64888,I65129,I65264);
nor I_3698 (I64876,I64999,I65264);
not I_3699 (I65432,I2514);
DFFARX1 I_3700 (I1290033,I2507,I65432,I65458,);
not I_3701 (I65466,I65458);
nand I_3702 (I65483,I1290036,I1290030);
and I_3703 (I65500,I65483,I1290027);
DFFARX1 I_3704 (I65500,I2507,I65432,I65526,);
DFFARX1 I_3705 (I1290012,I2507,I65432,I65543,);
and I_3706 (I65551,I65543,I1290021);
nor I_3707 (I65568,I65526,I65551);
DFFARX1 I_3708 (I65568,I2507,I65432,I65400,);
nand I_3709 (I65599,I65543,I1290021);
nand I_3710 (I65616,I65466,I65599);
not I_3711 (I65412,I65616);
DFFARX1 I_3712 (I1290012,I2507,I65432,I65656,);
DFFARX1 I_3713 (I65656,I2507,I65432,I65421,);
nand I_3714 (I65678,I1290015,I1290018);
and I_3715 (I65695,I65678,I1290024);
DFFARX1 I_3716 (I65695,I2507,I65432,I65721,);
DFFARX1 I_3717 (I65721,I2507,I65432,I65738,);
not I_3718 (I65424,I65738);
not I_3719 (I65760,I65721);
nand I_3720 (I65409,I65760,I65599);
nor I_3721 (I65791,I1290015,I1290018);
not I_3722 (I65808,I65791);
nor I_3723 (I65825,I65760,I65808);
nor I_3724 (I65842,I65466,I65825);
DFFARX1 I_3725 (I65842,I2507,I65432,I65418,);
nor I_3726 (I65873,I65526,I65808);
nor I_3727 (I65406,I65721,I65873);
nor I_3728 (I65415,I65656,I65791);
nor I_3729 (I65403,I65526,I65791);
not I_3730 (I65959,I2514);
DFFARX1 I_3731 (I181777,I2507,I65959,I65985,);
not I_3732 (I65993,I65985);
nand I_3733 (I66010,I181771,I181765);
and I_3734 (I66027,I66010,I181786);
DFFARX1 I_3735 (I66027,I2507,I65959,I66053,);
DFFARX1 I_3736 (I181783,I2507,I65959,I66070,);
and I_3737 (I66078,I66070,I181780);
nor I_3738 (I66095,I66053,I66078);
DFFARX1 I_3739 (I66095,I2507,I65959,I65927,);
nand I_3740 (I66126,I66070,I181780);
nand I_3741 (I66143,I65993,I66126);
not I_3742 (I65939,I66143);
DFFARX1 I_3743 (I181765,I2507,I65959,I66183,);
DFFARX1 I_3744 (I66183,I2507,I65959,I65948,);
nand I_3745 (I66205,I181768,I181768);
and I_3746 (I66222,I66205,I181789);
DFFARX1 I_3747 (I66222,I2507,I65959,I66248,);
DFFARX1 I_3748 (I66248,I2507,I65959,I66265,);
not I_3749 (I65951,I66265);
not I_3750 (I66287,I66248);
nand I_3751 (I65936,I66287,I66126);
nor I_3752 (I66318,I181774,I181768);
not I_3753 (I66335,I66318);
nor I_3754 (I66352,I66287,I66335);
nor I_3755 (I66369,I65993,I66352);
DFFARX1 I_3756 (I66369,I2507,I65959,I65945,);
nor I_3757 (I66400,I66053,I66335);
nor I_3758 (I65933,I66248,I66400);
nor I_3759 (I65942,I66183,I66318);
nor I_3760 (I65930,I66053,I66318);
not I_3761 (I66486,I2514);
DFFARX1 I_3762 (I399009,I2507,I66486,I66512,);
not I_3763 (I66520,I66512);
nand I_3764 (I66537,I399003,I398994);
and I_3765 (I66554,I66537,I399015);
DFFARX1 I_3766 (I66554,I2507,I66486,I66580,);
DFFARX1 I_3767 (I398997,I2507,I66486,I66597,);
and I_3768 (I66605,I66597,I398991);
nor I_3769 (I66622,I66580,I66605);
DFFARX1 I_3770 (I66622,I2507,I66486,I66454,);
nand I_3771 (I66653,I66597,I398991);
nand I_3772 (I66670,I66520,I66653);
not I_3773 (I66466,I66670);
DFFARX1 I_3774 (I398991,I2507,I66486,I66710,);
DFFARX1 I_3775 (I66710,I2507,I66486,I66475,);
nand I_3776 (I66732,I399018,I399000);
and I_3777 (I66749,I66732,I399006);
DFFARX1 I_3778 (I66749,I2507,I66486,I66775,);
DFFARX1 I_3779 (I66775,I2507,I66486,I66792,);
not I_3780 (I66478,I66792);
not I_3781 (I66814,I66775);
nand I_3782 (I66463,I66814,I66653);
nor I_3783 (I66845,I399012,I399000);
not I_3784 (I66862,I66845);
nor I_3785 (I66879,I66814,I66862);
nor I_3786 (I66896,I66520,I66879);
DFFARX1 I_3787 (I66896,I2507,I66486,I66472,);
nor I_3788 (I66927,I66580,I66862);
nor I_3789 (I66460,I66775,I66927);
nor I_3790 (I66469,I66710,I66845);
nor I_3791 (I66457,I66580,I66845);
not I_3792 (I67013,I2514);
DFFARX1 I_3793 (I907606,I2507,I67013,I67039,);
not I_3794 (I67047,I67039);
nand I_3795 (I67064,I907624,I907618);
and I_3796 (I67081,I67064,I907597);
DFFARX1 I_3797 (I67081,I2507,I67013,I67107,);
DFFARX1 I_3798 (I907615,I2507,I67013,I67124,);
and I_3799 (I67132,I67124,I907600);
nor I_3800 (I67149,I67107,I67132);
DFFARX1 I_3801 (I67149,I2507,I67013,I66981,);
nand I_3802 (I67180,I67124,I907600);
nand I_3803 (I67197,I67047,I67180);
not I_3804 (I66993,I67197);
DFFARX1 I_3805 (I907612,I2507,I67013,I67237,);
DFFARX1 I_3806 (I67237,I2507,I67013,I67002,);
nand I_3807 (I67259,I907621,I907609);
and I_3808 (I67276,I67259,I907603);
DFFARX1 I_3809 (I67276,I2507,I67013,I67302,);
DFFARX1 I_3810 (I67302,I2507,I67013,I67319,);
not I_3811 (I67005,I67319);
not I_3812 (I67341,I67302);
nand I_3813 (I66990,I67341,I67180);
nor I_3814 (I67372,I907597,I907609);
not I_3815 (I67389,I67372);
nor I_3816 (I67406,I67341,I67389);
nor I_3817 (I67423,I67047,I67406);
DFFARX1 I_3818 (I67423,I2507,I67013,I66999,);
nor I_3819 (I67454,I67107,I67389);
nor I_3820 (I66987,I67302,I67454);
nor I_3821 (I66996,I67237,I67372);
nor I_3822 (I66984,I67107,I67372);
not I_3823 (I67540,I2514);
DFFARX1 I_3824 (I685062,I2507,I67540,I67566,);
not I_3825 (I67574,I67566);
nand I_3826 (I67591,I685053,I685071);
and I_3827 (I67608,I67591,I685050);
DFFARX1 I_3828 (I67608,I2507,I67540,I67634,);
DFFARX1 I_3829 (I685053,I2507,I67540,I67651,);
and I_3830 (I67659,I67651,I685056);
nor I_3831 (I67676,I67634,I67659);
DFFARX1 I_3832 (I67676,I2507,I67540,I67508,);
nand I_3833 (I67707,I67651,I685056);
nand I_3834 (I67724,I67574,I67707);
not I_3835 (I67520,I67724);
DFFARX1 I_3836 (I685050,I2507,I67540,I67764,);
DFFARX1 I_3837 (I67764,I2507,I67540,I67529,);
nand I_3838 (I67786,I685068,I685059);
and I_3839 (I67803,I67786,I685074);
DFFARX1 I_3840 (I67803,I2507,I67540,I67829,);
DFFARX1 I_3841 (I67829,I2507,I67540,I67846,);
not I_3842 (I67532,I67846);
not I_3843 (I67868,I67829);
nand I_3844 (I67517,I67868,I67707);
nor I_3845 (I67899,I685065,I685059);
not I_3846 (I67916,I67899);
nor I_3847 (I67933,I67868,I67916);
nor I_3848 (I67950,I67574,I67933);
DFFARX1 I_3849 (I67950,I2507,I67540,I67526,);
nor I_3850 (I67981,I67634,I67916);
nor I_3851 (I67514,I67829,I67981);
nor I_3852 (I67523,I67764,I67899);
nor I_3853 (I67511,I67634,I67899);
not I_3854 (I68067,I2514);
DFFARX1 I_3855 (I144301,I2507,I68067,I68093,);
not I_3856 (I68101,I68093);
nand I_3857 (I68118,I144298,I144280);
and I_3858 (I68135,I68118,I144286);
DFFARX1 I_3859 (I68135,I2507,I68067,I68161,);
DFFARX1 I_3860 (I144295,I2507,I68067,I68178,);
and I_3861 (I68186,I68178,I144289);
nor I_3862 (I68203,I68161,I68186);
DFFARX1 I_3863 (I68203,I2507,I68067,I68035,);
nand I_3864 (I68234,I68178,I144289);
nand I_3865 (I68251,I68101,I68234);
not I_3866 (I68047,I68251);
DFFARX1 I_3867 (I144304,I2507,I68067,I68291,);
DFFARX1 I_3868 (I68291,I2507,I68067,I68056,);
nand I_3869 (I68313,I144292,I144283);
and I_3870 (I68330,I68313,I144280);
DFFARX1 I_3871 (I68330,I2507,I68067,I68356,);
DFFARX1 I_3872 (I68356,I2507,I68067,I68373,);
not I_3873 (I68059,I68373);
not I_3874 (I68395,I68356);
nand I_3875 (I68044,I68395,I68234);
nor I_3876 (I68426,I144307,I144283);
not I_3877 (I68443,I68426);
nor I_3878 (I68460,I68395,I68443);
nor I_3879 (I68477,I68101,I68460);
DFFARX1 I_3880 (I68477,I2507,I68067,I68053,);
nor I_3881 (I68508,I68161,I68443);
nor I_3882 (I68041,I68356,I68508);
nor I_3883 (I68050,I68291,I68426);
nor I_3884 (I68038,I68161,I68426);
not I_3885 (I68594,I2514);
DFFARX1 I_3886 (I476257,I2507,I68594,I68620,);
not I_3887 (I68628,I68620);
nand I_3888 (I68645,I476251,I476242);
and I_3889 (I68662,I68645,I476263);
DFFARX1 I_3890 (I68662,I2507,I68594,I68688,);
DFFARX1 I_3891 (I476245,I2507,I68594,I68705,);
and I_3892 (I68713,I68705,I476239);
nor I_3893 (I68730,I68688,I68713);
DFFARX1 I_3894 (I68730,I2507,I68594,I68562,);
nand I_3895 (I68761,I68705,I476239);
nand I_3896 (I68778,I68628,I68761);
not I_3897 (I68574,I68778);
DFFARX1 I_3898 (I476239,I2507,I68594,I68818,);
DFFARX1 I_3899 (I68818,I2507,I68594,I68583,);
nand I_3900 (I68840,I476266,I476248);
and I_3901 (I68857,I68840,I476254);
DFFARX1 I_3902 (I68857,I2507,I68594,I68883,);
DFFARX1 I_3903 (I68883,I2507,I68594,I68900,);
not I_3904 (I68586,I68900);
not I_3905 (I68922,I68883);
nand I_3906 (I68571,I68922,I68761);
nor I_3907 (I68953,I476260,I476248);
not I_3908 (I68970,I68953);
nor I_3909 (I68987,I68922,I68970);
nor I_3910 (I69004,I68628,I68987);
DFFARX1 I_3911 (I69004,I2507,I68594,I68580,);
nor I_3912 (I69035,I68688,I68970);
nor I_3913 (I68568,I68883,I69035);
nor I_3914 (I68577,I68818,I68953);
nor I_3915 (I68565,I68688,I68953);
not I_3916 (I69121,I2514);
DFFARX1 I_3917 (I1033145,I2507,I69121,I69147,);
not I_3918 (I69155,I69147);
nand I_3919 (I69172,I1033142,I1033148);
and I_3920 (I69189,I69172,I1033145);
DFFARX1 I_3921 (I69189,I2507,I69121,I69215,);
DFFARX1 I_3922 (I1033148,I2507,I69121,I69232,);
and I_3923 (I69240,I69232,I1033142);
nor I_3924 (I69257,I69215,I69240);
DFFARX1 I_3925 (I69257,I2507,I69121,I69089,);
nand I_3926 (I69288,I69232,I1033142);
nand I_3927 (I69305,I69155,I69288);
not I_3928 (I69101,I69305);
DFFARX1 I_3929 (I1033151,I2507,I69121,I69345,);
DFFARX1 I_3930 (I69345,I2507,I69121,I69110,);
nand I_3931 (I69367,I1033154,I1033163);
and I_3932 (I69384,I69367,I1033157);
DFFARX1 I_3933 (I69384,I2507,I69121,I69410,);
DFFARX1 I_3934 (I69410,I2507,I69121,I69427,);
not I_3935 (I69113,I69427);
not I_3936 (I69449,I69410);
nand I_3937 (I69098,I69449,I69288);
nor I_3938 (I69480,I1033160,I1033163);
not I_3939 (I69497,I69480);
nor I_3940 (I69514,I69449,I69497);
nor I_3941 (I69531,I69155,I69514);
DFFARX1 I_3942 (I69531,I2507,I69121,I69107,);
nor I_3943 (I69562,I69215,I69497);
nor I_3944 (I69095,I69410,I69562);
nor I_3945 (I69104,I69345,I69480);
nor I_3946 (I69092,I69215,I69480);
not I_3947 (I69648,I2514);
DFFARX1 I_3948 (I797514,I2507,I69648,I69674,);
not I_3949 (I69682,I69674);
nand I_3950 (I69699,I797511,I797526);
and I_3951 (I69716,I69699,I797508);
DFFARX1 I_3952 (I69716,I2507,I69648,I69742,);
DFFARX1 I_3953 (I797505,I2507,I69648,I69759,);
and I_3954 (I69767,I69759,I797505);
nor I_3955 (I69784,I69742,I69767);
DFFARX1 I_3956 (I69784,I2507,I69648,I69616,);
nand I_3957 (I69815,I69759,I797505);
nand I_3958 (I69832,I69682,I69815);
not I_3959 (I69628,I69832);
DFFARX1 I_3960 (I797508,I2507,I69648,I69872,);
DFFARX1 I_3961 (I69872,I2507,I69648,I69637,);
nand I_3962 (I69894,I797520,I797511);
and I_3963 (I69911,I69894,I797523);
DFFARX1 I_3964 (I69911,I2507,I69648,I69937,);
DFFARX1 I_3965 (I69937,I2507,I69648,I69954,);
not I_3966 (I69640,I69954);
not I_3967 (I69976,I69937);
nand I_3968 (I69625,I69976,I69815);
nor I_3969 (I70007,I797517,I797511);
not I_3970 (I70024,I70007);
nor I_3971 (I70041,I69976,I70024);
nor I_3972 (I70058,I69682,I70041);
DFFARX1 I_3973 (I70058,I2507,I69648,I69634,);
nor I_3974 (I70089,I69742,I70024);
nor I_3975 (I69622,I69937,I70089);
nor I_3976 (I69631,I69872,I70007);
nor I_3977 (I69619,I69742,I70007);
not I_3978 (I70175,I2514);
DFFARX1 I_3979 (I872875,I2507,I70175,I70201,);
not I_3980 (I70209,I70201);
nand I_3981 (I70226,I872872,I872887);
and I_3982 (I70243,I70226,I872869);
DFFARX1 I_3983 (I70243,I2507,I70175,I70269,);
DFFARX1 I_3984 (I872866,I2507,I70175,I70286,);
and I_3985 (I70294,I70286,I872866);
nor I_3986 (I70311,I70269,I70294);
DFFARX1 I_3987 (I70311,I2507,I70175,I70143,);
nand I_3988 (I70342,I70286,I872866);
nand I_3989 (I70359,I70209,I70342);
not I_3990 (I70155,I70359);
DFFARX1 I_3991 (I872869,I2507,I70175,I70399,);
DFFARX1 I_3992 (I70399,I2507,I70175,I70164,);
nand I_3993 (I70421,I872881,I872872);
and I_3994 (I70438,I70421,I872884);
DFFARX1 I_3995 (I70438,I2507,I70175,I70464,);
DFFARX1 I_3996 (I70464,I2507,I70175,I70481,);
not I_3997 (I70167,I70481);
not I_3998 (I70503,I70464);
nand I_3999 (I70152,I70503,I70342);
nor I_4000 (I70534,I872878,I872872);
not I_4001 (I70551,I70534);
nor I_4002 (I70568,I70503,I70551);
nor I_4003 (I70585,I70209,I70568);
DFFARX1 I_4004 (I70585,I2507,I70175,I70161,);
nor I_4005 (I70616,I70269,I70551);
nor I_4006 (I70149,I70464,I70616);
nor I_4007 (I70158,I70399,I70534);
nor I_4008 (I70146,I70269,I70534);
not I_4009 (I70702,I2514);
DFFARX1 I_4010 (I1287143,I2507,I70702,I70728,);
not I_4011 (I70736,I70728);
nand I_4012 (I70753,I1287146,I1287140);
and I_4013 (I70770,I70753,I1287137);
DFFARX1 I_4014 (I70770,I2507,I70702,I70796,);
DFFARX1 I_4015 (I1287122,I2507,I70702,I70813,);
and I_4016 (I70821,I70813,I1287131);
nor I_4017 (I70838,I70796,I70821);
DFFARX1 I_4018 (I70838,I2507,I70702,I70670,);
nand I_4019 (I70869,I70813,I1287131);
nand I_4020 (I70886,I70736,I70869);
not I_4021 (I70682,I70886);
DFFARX1 I_4022 (I1287122,I2507,I70702,I70926,);
DFFARX1 I_4023 (I70926,I2507,I70702,I70691,);
nand I_4024 (I70948,I1287125,I1287128);
and I_4025 (I70965,I70948,I1287134);
DFFARX1 I_4026 (I70965,I2507,I70702,I70991,);
DFFARX1 I_4027 (I70991,I2507,I70702,I71008,);
not I_4028 (I70694,I71008);
not I_4029 (I71030,I70991);
nand I_4030 (I70679,I71030,I70869);
nor I_4031 (I71061,I1287125,I1287128);
not I_4032 (I71078,I71061);
nor I_4033 (I71095,I71030,I71078);
nor I_4034 (I71112,I70736,I71095);
DFFARX1 I_4035 (I71112,I2507,I70702,I70688,);
nor I_4036 (I71143,I70796,I71078);
nor I_4037 (I70676,I70991,I71143);
nor I_4038 (I70685,I70926,I71061);
nor I_4039 (I70673,I70796,I71061);
not I_4040 (I71229,I2514);
DFFARX1 I_4041 (I21683,I2507,I71229,I71255,);
not I_4042 (I71263,I71255);
nand I_4043 (I71280,I21671,I21677);
and I_4044 (I71297,I71280,I21680);
DFFARX1 I_4045 (I71297,I2507,I71229,I71323,);
DFFARX1 I_4046 (I21662,I2507,I71229,I71340,);
and I_4047 (I71348,I71340,I21668);
nor I_4048 (I71365,I71323,I71348);
DFFARX1 I_4049 (I71365,I2507,I71229,I71197,);
nand I_4050 (I71396,I71340,I21668);
nand I_4051 (I71413,I71263,I71396);
not I_4052 (I71209,I71413);
DFFARX1 I_4053 (I21662,I2507,I71229,I71453,);
DFFARX1 I_4054 (I71453,I2507,I71229,I71218,);
nand I_4055 (I71475,I21665,I21659);
and I_4056 (I71492,I71475,I21674);
DFFARX1 I_4057 (I71492,I2507,I71229,I71518,);
DFFARX1 I_4058 (I71518,I2507,I71229,I71535,);
not I_4059 (I71221,I71535);
not I_4060 (I71557,I71518);
nand I_4061 (I71206,I71557,I71396);
nor I_4062 (I71588,I21659,I21659);
not I_4063 (I71605,I71588);
nor I_4064 (I71622,I71557,I71605);
nor I_4065 (I71639,I71263,I71622);
DFFARX1 I_4066 (I71639,I2507,I71229,I71215,);
nor I_4067 (I71670,I71323,I71605);
nor I_4068 (I71203,I71518,I71670);
nor I_4069 (I71212,I71453,I71588);
nor I_4070 (I71200,I71323,I71588);
not I_4071 (I71756,I2514);
DFFARX1 I_4072 (I1345189,I2507,I71756,I71782,);
not I_4073 (I71790,I71782);
nand I_4074 (I71807,I1345183,I1345204);
and I_4075 (I71824,I71807,I1345180);
DFFARX1 I_4076 (I71824,I2507,I71756,I71850,);
DFFARX1 I_4077 (I1345201,I2507,I71756,I71867,);
and I_4078 (I71875,I71867,I1345198);
nor I_4079 (I71892,I71850,I71875);
DFFARX1 I_4080 (I71892,I2507,I71756,I71724,);
nand I_4081 (I71923,I71867,I1345198);
nand I_4082 (I71940,I71790,I71923);
not I_4083 (I71736,I71940);
DFFARX1 I_4084 (I1345186,I2507,I71756,I71980,);
DFFARX1 I_4085 (I71980,I2507,I71756,I71745,);
nand I_4086 (I72002,I1345195,I1345192);
and I_4087 (I72019,I72002,I1345177);
DFFARX1 I_4088 (I72019,I2507,I71756,I72045,);
DFFARX1 I_4089 (I72045,I2507,I71756,I72062,);
not I_4090 (I71748,I72062);
not I_4091 (I72084,I72045);
nand I_4092 (I71733,I72084,I71923);
nor I_4093 (I72115,I1345177,I1345192);
not I_4094 (I72132,I72115);
nor I_4095 (I72149,I72084,I72132);
nor I_4096 (I72166,I71790,I72149);
DFFARX1 I_4097 (I72166,I2507,I71756,I71742,);
nor I_4098 (I72197,I71850,I72132);
nor I_4099 (I71730,I72045,I72197);
nor I_4100 (I71739,I71980,I72115);
nor I_4101 (I71727,I71850,I72115);
not I_4102 (I72283,I2514);
DFFARX1 I_4103 (I484961,I2507,I72283,I72309,);
not I_4104 (I72317,I72309);
nand I_4105 (I72334,I484955,I484946);
and I_4106 (I72351,I72334,I484967);
DFFARX1 I_4107 (I72351,I2507,I72283,I72377,);
DFFARX1 I_4108 (I484949,I2507,I72283,I72394,);
and I_4109 (I72402,I72394,I484943);
nor I_4110 (I72419,I72377,I72402);
DFFARX1 I_4111 (I72419,I2507,I72283,I72251,);
nand I_4112 (I72450,I72394,I484943);
nand I_4113 (I72467,I72317,I72450);
not I_4114 (I72263,I72467);
DFFARX1 I_4115 (I484943,I2507,I72283,I72507,);
DFFARX1 I_4116 (I72507,I2507,I72283,I72272,);
nand I_4117 (I72529,I484970,I484952);
and I_4118 (I72546,I72529,I484958);
DFFARX1 I_4119 (I72546,I2507,I72283,I72572,);
DFFARX1 I_4120 (I72572,I2507,I72283,I72589,);
not I_4121 (I72275,I72589);
not I_4122 (I72611,I72572);
nand I_4123 (I72260,I72611,I72450);
nor I_4124 (I72642,I484964,I484952);
not I_4125 (I72659,I72642);
nor I_4126 (I72676,I72611,I72659);
nor I_4127 (I72693,I72317,I72676);
DFFARX1 I_4128 (I72693,I2507,I72283,I72269,);
nor I_4129 (I72724,I72377,I72659);
nor I_4130 (I72257,I72572,I72724);
nor I_4131 (I72266,I72507,I72642);
nor I_4132 (I72254,I72377,I72642);
not I_4133 (I72810,I2514);
DFFARX1 I_4134 (I473537,I2507,I72810,I72836,);
not I_4135 (I72844,I72836);
nand I_4136 (I72861,I473531,I473522);
and I_4137 (I72878,I72861,I473543);
DFFARX1 I_4138 (I72878,I2507,I72810,I72904,);
DFFARX1 I_4139 (I473525,I2507,I72810,I72921,);
and I_4140 (I72929,I72921,I473519);
nor I_4141 (I72946,I72904,I72929);
DFFARX1 I_4142 (I72946,I2507,I72810,I72778,);
nand I_4143 (I72977,I72921,I473519);
nand I_4144 (I72994,I72844,I72977);
not I_4145 (I72790,I72994);
DFFARX1 I_4146 (I473519,I2507,I72810,I73034,);
DFFARX1 I_4147 (I73034,I2507,I72810,I72799,);
nand I_4148 (I73056,I473546,I473528);
and I_4149 (I73073,I73056,I473534);
DFFARX1 I_4150 (I73073,I2507,I72810,I73099,);
DFFARX1 I_4151 (I73099,I2507,I72810,I73116,);
not I_4152 (I72802,I73116);
not I_4153 (I73138,I73099);
nand I_4154 (I72787,I73138,I72977);
nor I_4155 (I73169,I473540,I473528);
not I_4156 (I73186,I73169);
nor I_4157 (I73203,I73138,I73186);
nor I_4158 (I73220,I72844,I73203);
DFFARX1 I_4159 (I73220,I2507,I72810,I72796,);
nor I_4160 (I73251,I72904,I73186);
nor I_4161 (I72784,I73099,I73251);
nor I_4162 (I72793,I73034,I73169);
nor I_4163 (I72781,I72904,I73169);
not I_4164 (I73337,I2514);
DFFARX1 I_4165 (I1243880,I2507,I73337,I73363,);
not I_4166 (I73371,I73363);
nand I_4167 (I73388,I1243874,I1243895);
and I_4168 (I73405,I73388,I1243886);
DFFARX1 I_4169 (I73405,I2507,I73337,I73431,);
DFFARX1 I_4170 (I1243877,I2507,I73337,I73448,);
and I_4171 (I73456,I73448,I1243889);
nor I_4172 (I73473,I73431,I73456);
DFFARX1 I_4173 (I73473,I2507,I73337,I73305,);
nand I_4174 (I73504,I73448,I1243889);
nand I_4175 (I73521,I73371,I73504);
not I_4176 (I73317,I73521);
DFFARX1 I_4177 (I1243877,I2507,I73337,I73561,);
DFFARX1 I_4178 (I73561,I2507,I73337,I73326,);
nand I_4179 (I73583,I1243898,I1243883);
and I_4180 (I73600,I73583,I1243874);
DFFARX1 I_4181 (I73600,I2507,I73337,I73626,);
DFFARX1 I_4182 (I73626,I2507,I73337,I73643,);
not I_4183 (I73329,I73643);
not I_4184 (I73665,I73626);
nand I_4185 (I73314,I73665,I73504);
nor I_4186 (I73696,I1243892,I1243883);
not I_4187 (I73713,I73696);
nor I_4188 (I73730,I73665,I73713);
nor I_4189 (I73747,I73371,I73730);
DFFARX1 I_4190 (I73747,I2507,I73337,I73323,);
nor I_4191 (I73778,I73431,I73713);
nor I_4192 (I73311,I73626,I73778);
nor I_4193 (I73320,I73561,I73696);
nor I_4194 (I73308,I73431,I73696);
not I_4195 (I73864,I2514);
DFFARX1 I_4196 (I280783,I2507,I73864,I73890,);
not I_4197 (I73898,I73890);
nand I_4198 (I73915,I280765,I280780);
and I_4199 (I73932,I73915,I280756);
DFFARX1 I_4200 (I73932,I2507,I73864,I73958,);
DFFARX1 I_4201 (I280759,I2507,I73864,I73975,);
and I_4202 (I73983,I73975,I280774);
nor I_4203 (I74000,I73958,I73983);
DFFARX1 I_4204 (I74000,I2507,I73864,I73832,);
nand I_4205 (I74031,I73975,I280774);
nand I_4206 (I74048,I73898,I74031);
not I_4207 (I73844,I74048);
DFFARX1 I_4208 (I280777,I2507,I73864,I74088,);
DFFARX1 I_4209 (I74088,I2507,I73864,I73853,);
nand I_4210 (I74110,I280756,I280768);
and I_4211 (I74127,I74110,I280762);
DFFARX1 I_4212 (I74127,I2507,I73864,I74153,);
DFFARX1 I_4213 (I74153,I2507,I73864,I74170,);
not I_4214 (I73856,I74170);
not I_4215 (I74192,I74153);
nand I_4216 (I73841,I74192,I74031);
nor I_4217 (I74223,I280771,I280768);
not I_4218 (I74240,I74223);
nor I_4219 (I74257,I74192,I74240);
nor I_4220 (I74274,I73898,I74257);
DFFARX1 I_4221 (I74274,I2507,I73864,I73850,);
nor I_4222 (I74305,I73958,I74240);
nor I_4223 (I73838,I74153,I74305);
nor I_4224 (I73847,I74088,I74223);
nor I_4225 (I73835,I73958,I74223);
not I_4226 (I74391,I2514);
DFFARX1 I_4227 (I254960,I2507,I74391,I74417,);
not I_4228 (I74425,I74417);
nand I_4229 (I74442,I254942,I254957);
and I_4230 (I74459,I74442,I254933);
DFFARX1 I_4231 (I74459,I2507,I74391,I74485,);
DFFARX1 I_4232 (I254936,I2507,I74391,I74502,);
and I_4233 (I74510,I74502,I254951);
nor I_4234 (I74527,I74485,I74510);
DFFARX1 I_4235 (I74527,I2507,I74391,I74359,);
nand I_4236 (I74558,I74502,I254951);
nand I_4237 (I74575,I74425,I74558);
not I_4238 (I74371,I74575);
DFFARX1 I_4239 (I254954,I2507,I74391,I74615,);
DFFARX1 I_4240 (I74615,I2507,I74391,I74380,);
nand I_4241 (I74637,I254933,I254945);
and I_4242 (I74654,I74637,I254939);
DFFARX1 I_4243 (I74654,I2507,I74391,I74680,);
DFFARX1 I_4244 (I74680,I2507,I74391,I74697,);
not I_4245 (I74383,I74697);
not I_4246 (I74719,I74680);
nand I_4247 (I74368,I74719,I74558);
nor I_4248 (I74750,I254948,I254945);
not I_4249 (I74767,I74750);
nor I_4250 (I74784,I74719,I74767);
nor I_4251 (I74801,I74425,I74784);
DFFARX1 I_4252 (I74801,I2507,I74391,I74377,);
nor I_4253 (I74832,I74485,I74767);
nor I_4254 (I74365,I74680,I74832);
nor I_4255 (I74374,I74615,I74750);
nor I_4256 (I74362,I74485,I74750);
not I_4257 (I74918,I2514);
DFFARX1 I_4258 (I835985,I2507,I74918,I74944,);
not I_4259 (I74952,I74944);
nand I_4260 (I74969,I835982,I835997);
and I_4261 (I74986,I74969,I835979);
DFFARX1 I_4262 (I74986,I2507,I74918,I75012,);
DFFARX1 I_4263 (I835976,I2507,I74918,I75029,);
and I_4264 (I75037,I75029,I835976);
nor I_4265 (I75054,I75012,I75037);
DFFARX1 I_4266 (I75054,I2507,I74918,I74886,);
nand I_4267 (I75085,I75029,I835976);
nand I_4268 (I75102,I74952,I75085);
not I_4269 (I74898,I75102);
DFFARX1 I_4270 (I835979,I2507,I74918,I75142,);
DFFARX1 I_4271 (I75142,I2507,I74918,I74907,);
nand I_4272 (I75164,I835991,I835982);
and I_4273 (I75181,I75164,I835994);
DFFARX1 I_4274 (I75181,I2507,I74918,I75207,);
DFFARX1 I_4275 (I75207,I2507,I74918,I75224,);
not I_4276 (I74910,I75224);
not I_4277 (I75246,I75207);
nand I_4278 (I74895,I75246,I75085);
nor I_4279 (I75277,I835988,I835982);
not I_4280 (I75294,I75277);
nor I_4281 (I75311,I75246,I75294);
nor I_4282 (I75328,I74952,I75311);
DFFARX1 I_4283 (I75328,I2507,I74918,I74904,);
nor I_4284 (I75359,I75012,I75294);
nor I_4285 (I74892,I75207,I75359);
nor I_4286 (I74901,I75142,I75277);
nor I_4287 (I74889,I75012,I75277);
not I_4288 (I75445,I2514);
DFFARX1 I_4289 (I223427,I2507,I75445,I75471,);
not I_4290 (I75479,I75471);
nand I_4291 (I75496,I223421,I223415);
and I_4292 (I75513,I75496,I223436);
DFFARX1 I_4293 (I75513,I2507,I75445,I75539,);
DFFARX1 I_4294 (I223433,I2507,I75445,I75556,);
and I_4295 (I75564,I75556,I223430);
nor I_4296 (I75581,I75539,I75564);
DFFARX1 I_4297 (I75581,I2507,I75445,I75413,);
nand I_4298 (I75612,I75556,I223430);
nand I_4299 (I75629,I75479,I75612);
not I_4300 (I75425,I75629);
DFFARX1 I_4301 (I223415,I2507,I75445,I75669,);
DFFARX1 I_4302 (I75669,I2507,I75445,I75434,);
nand I_4303 (I75691,I223418,I223418);
and I_4304 (I75708,I75691,I223439);
DFFARX1 I_4305 (I75708,I2507,I75445,I75734,);
DFFARX1 I_4306 (I75734,I2507,I75445,I75751,);
not I_4307 (I75437,I75751);
not I_4308 (I75773,I75734);
nand I_4309 (I75422,I75773,I75612);
nor I_4310 (I75804,I223424,I223418);
not I_4311 (I75821,I75804);
nor I_4312 (I75838,I75773,I75821);
nor I_4313 (I75855,I75479,I75838);
DFFARX1 I_4314 (I75855,I2507,I75445,I75431,);
nor I_4315 (I75886,I75539,I75821);
nor I_4316 (I75419,I75734,I75886);
nor I_4317 (I75428,I75669,I75804);
nor I_4318 (I75416,I75539,I75804);
not I_4319 (I75972,I2514);
DFFARX1 I_4320 (I1157214,I2507,I75972,I75998,);
not I_4321 (I76006,I75998);
nand I_4322 (I76023,I1157229,I1157208);
and I_4323 (I76040,I76023,I1157211);
DFFARX1 I_4324 (I76040,I2507,I75972,I76066,);
DFFARX1 I_4325 (I1157232,I2507,I75972,I76083,);
and I_4326 (I76091,I76083,I1157211);
nor I_4327 (I76108,I76066,I76091);
DFFARX1 I_4328 (I76108,I2507,I75972,I75940,);
nand I_4329 (I76139,I76083,I1157211);
nand I_4330 (I76156,I76006,I76139);
not I_4331 (I75952,I76156);
DFFARX1 I_4332 (I1157208,I2507,I75972,I76196,);
DFFARX1 I_4333 (I76196,I2507,I75972,I75961,);
nand I_4334 (I76218,I1157220,I1157217);
and I_4335 (I76235,I76218,I1157223);
DFFARX1 I_4336 (I76235,I2507,I75972,I76261,);
DFFARX1 I_4337 (I76261,I2507,I75972,I76278,);
not I_4338 (I75964,I76278);
not I_4339 (I76300,I76261);
nand I_4340 (I75949,I76300,I76139);
nor I_4341 (I76331,I1157226,I1157217);
not I_4342 (I76348,I76331);
nor I_4343 (I76365,I76300,I76348);
nor I_4344 (I76382,I76006,I76365);
DFFARX1 I_4345 (I76382,I2507,I75972,I75958,);
nor I_4346 (I76413,I76066,I76348);
nor I_4347 (I75946,I76261,I76413);
nor I_4348 (I75955,I76196,I76331);
nor I_4349 (I75943,I76066,I76331);
not I_4350 (I76499,I2514);
DFFARX1 I_4351 (I306606,I2507,I76499,I76525,);
not I_4352 (I76533,I76525);
nand I_4353 (I76550,I306588,I306603);
and I_4354 (I76567,I76550,I306579);
DFFARX1 I_4355 (I76567,I2507,I76499,I76593,);
DFFARX1 I_4356 (I306582,I2507,I76499,I76610,);
and I_4357 (I76618,I76610,I306597);
nor I_4358 (I76635,I76593,I76618);
DFFARX1 I_4359 (I76635,I2507,I76499,I76467,);
nand I_4360 (I76666,I76610,I306597);
nand I_4361 (I76683,I76533,I76666);
not I_4362 (I76479,I76683);
DFFARX1 I_4363 (I306600,I2507,I76499,I76723,);
DFFARX1 I_4364 (I76723,I2507,I76499,I76488,);
nand I_4365 (I76745,I306579,I306591);
and I_4366 (I76762,I76745,I306585);
DFFARX1 I_4367 (I76762,I2507,I76499,I76788,);
DFFARX1 I_4368 (I76788,I2507,I76499,I76805,);
not I_4369 (I76491,I76805);
not I_4370 (I76827,I76788);
nand I_4371 (I76476,I76827,I76666);
nor I_4372 (I76858,I306594,I306591);
not I_4373 (I76875,I76858);
nor I_4374 (I76892,I76827,I76875);
nor I_4375 (I76909,I76533,I76892);
DFFARX1 I_4376 (I76909,I2507,I76499,I76485,);
nor I_4377 (I76940,I76593,I76875);
nor I_4378 (I76473,I76788,I76940);
nor I_4379 (I76482,I76723,I76858);
nor I_4380 (I76470,I76593,I76858);
not I_4381 (I77026,I2514);
DFFARX1 I_4382 (I908898,I2507,I77026,I77052,);
not I_4383 (I77060,I77052);
nand I_4384 (I77077,I908916,I908910);
and I_4385 (I77094,I77077,I908889);
DFFARX1 I_4386 (I77094,I2507,I77026,I77120,);
DFFARX1 I_4387 (I908907,I2507,I77026,I77137,);
and I_4388 (I77145,I77137,I908892);
nor I_4389 (I77162,I77120,I77145);
DFFARX1 I_4390 (I77162,I2507,I77026,I76994,);
nand I_4391 (I77193,I77137,I908892);
nand I_4392 (I77210,I77060,I77193);
not I_4393 (I77006,I77210);
DFFARX1 I_4394 (I908904,I2507,I77026,I77250,);
DFFARX1 I_4395 (I77250,I2507,I77026,I77015,);
nand I_4396 (I77272,I908913,I908901);
and I_4397 (I77289,I77272,I908895);
DFFARX1 I_4398 (I77289,I2507,I77026,I77315,);
DFFARX1 I_4399 (I77315,I2507,I77026,I77332,);
not I_4400 (I77018,I77332);
not I_4401 (I77354,I77315);
nand I_4402 (I77003,I77354,I77193);
nor I_4403 (I77385,I908889,I908901);
not I_4404 (I77402,I77385);
nor I_4405 (I77419,I77354,I77402);
nor I_4406 (I77436,I77060,I77419);
DFFARX1 I_4407 (I77436,I2507,I77026,I77012,);
nor I_4408 (I77467,I77120,I77402);
nor I_4409 (I77000,I77315,I77467);
nor I_4410 (I77009,I77250,I77385);
nor I_4411 (I76997,I77120,I77385);
not I_4412 (I77553,I2514);
DFFARX1 I_4413 (I41182,I2507,I77553,I77579,);
not I_4414 (I77587,I77579);
nand I_4415 (I77604,I41170,I41176);
and I_4416 (I77621,I77604,I41179);
DFFARX1 I_4417 (I77621,I2507,I77553,I77647,);
DFFARX1 I_4418 (I41161,I2507,I77553,I77664,);
and I_4419 (I77672,I77664,I41167);
nor I_4420 (I77689,I77647,I77672);
DFFARX1 I_4421 (I77689,I2507,I77553,I77521,);
nand I_4422 (I77720,I77664,I41167);
nand I_4423 (I77737,I77587,I77720);
not I_4424 (I77533,I77737);
DFFARX1 I_4425 (I41161,I2507,I77553,I77777,);
DFFARX1 I_4426 (I77777,I2507,I77553,I77542,);
nand I_4427 (I77799,I41164,I41158);
and I_4428 (I77816,I77799,I41173);
DFFARX1 I_4429 (I77816,I2507,I77553,I77842,);
DFFARX1 I_4430 (I77842,I2507,I77553,I77859,);
not I_4431 (I77545,I77859);
not I_4432 (I77881,I77842);
nand I_4433 (I77530,I77881,I77720);
nor I_4434 (I77912,I41158,I41158);
not I_4435 (I77929,I77912);
nor I_4436 (I77946,I77881,I77929);
nor I_4437 (I77963,I77587,I77946);
DFFARX1 I_4438 (I77963,I2507,I77553,I77539,);
nor I_4439 (I77994,I77647,I77929);
nor I_4440 (I77527,I77842,I77994);
nor I_4441 (I77536,I77777,I77912);
nor I_4442 (I77524,I77647,I77912);
not I_4443 (I78080,I2514);
DFFARX1 I_4444 (I1095946,I2507,I78080,I78106,);
not I_4445 (I78114,I78106);
nand I_4446 (I78131,I1095961,I1095940);
and I_4447 (I78148,I78131,I1095943);
DFFARX1 I_4448 (I78148,I2507,I78080,I78174,);
DFFARX1 I_4449 (I1095964,I2507,I78080,I78191,);
and I_4450 (I78199,I78191,I1095943);
nor I_4451 (I78216,I78174,I78199);
DFFARX1 I_4452 (I78216,I2507,I78080,I78048,);
nand I_4453 (I78247,I78191,I1095943);
nand I_4454 (I78264,I78114,I78247);
not I_4455 (I78060,I78264);
DFFARX1 I_4456 (I1095940,I2507,I78080,I78304,);
DFFARX1 I_4457 (I78304,I2507,I78080,I78069,);
nand I_4458 (I78326,I1095952,I1095949);
and I_4459 (I78343,I78326,I1095955);
DFFARX1 I_4460 (I78343,I2507,I78080,I78369,);
DFFARX1 I_4461 (I78369,I2507,I78080,I78386,);
not I_4462 (I78072,I78386);
not I_4463 (I78408,I78369);
nand I_4464 (I78057,I78408,I78247);
nor I_4465 (I78439,I1095958,I1095949);
not I_4466 (I78456,I78439);
nor I_4467 (I78473,I78408,I78456);
nor I_4468 (I78490,I78114,I78473);
DFFARX1 I_4469 (I78490,I2507,I78080,I78066,);
nor I_4470 (I78521,I78174,I78456);
nor I_4471 (I78054,I78369,I78521);
nor I_4472 (I78063,I78304,I78439);
nor I_4473 (I78051,I78174,I78439);
not I_4474 (I78607,I2514);
DFFARX1 I_4475 (I5507,I2507,I78607,I78633,);
not I_4476 (I78641,I78633);
nand I_4477 (I78658,I5492,I5492);
and I_4478 (I78675,I78658,I5513);
DFFARX1 I_4479 (I78675,I2507,I78607,I78701,);
DFFARX1 I_4480 (I5495,I2507,I78607,I78718,);
and I_4481 (I78726,I78718,I5504);
nor I_4482 (I78743,I78701,I78726);
DFFARX1 I_4483 (I78743,I2507,I78607,I78575,);
nand I_4484 (I78774,I78718,I5504);
nand I_4485 (I78791,I78641,I78774);
not I_4486 (I78587,I78791);
DFFARX1 I_4487 (I5498,I2507,I78607,I78831,);
DFFARX1 I_4488 (I78831,I2507,I78607,I78596,);
nand I_4489 (I78853,I5501,I5510);
and I_4490 (I78870,I78853,I5495);
DFFARX1 I_4491 (I78870,I2507,I78607,I78896,);
DFFARX1 I_4492 (I78896,I2507,I78607,I78913,);
not I_4493 (I78599,I78913);
not I_4494 (I78935,I78896);
nand I_4495 (I78584,I78935,I78774);
nor I_4496 (I78966,I5498,I5510);
not I_4497 (I78983,I78966);
nor I_4498 (I79000,I78935,I78983);
nor I_4499 (I79017,I78641,I79000);
DFFARX1 I_4500 (I79017,I2507,I78607,I78593,);
nor I_4501 (I79048,I78701,I78983);
nor I_4502 (I78581,I78896,I79048);
nor I_4503 (I78590,I78831,I78966);
nor I_4504 (I78578,I78701,I78966);
not I_4505 (I79134,I2514);
DFFARX1 I_4506 (I529792,I2507,I79134,I79160,);
not I_4507 (I79168,I79160);
nand I_4508 (I79185,I529813,I529807);
and I_4509 (I79202,I79185,I529789);
DFFARX1 I_4510 (I79202,I2507,I79134,I79228,);
DFFARX1 I_4511 (I529792,I2507,I79134,I79245,);
and I_4512 (I79253,I79245,I529801);
nor I_4513 (I79270,I79228,I79253);
DFFARX1 I_4514 (I79270,I2507,I79134,I79102,);
nand I_4515 (I79301,I79245,I529801);
nand I_4516 (I79318,I79168,I79301);
not I_4517 (I79114,I79318);
DFFARX1 I_4518 (I529798,I2507,I79134,I79358,);
DFFARX1 I_4519 (I79358,I2507,I79134,I79123,);
nand I_4520 (I79380,I529804,I529795);
and I_4521 (I79397,I79380,I529789);
DFFARX1 I_4522 (I79397,I2507,I79134,I79423,);
DFFARX1 I_4523 (I79423,I2507,I79134,I79440,);
not I_4524 (I79126,I79440);
not I_4525 (I79462,I79423);
nand I_4526 (I79111,I79462,I79301);
nor I_4527 (I79493,I529810,I529795);
not I_4528 (I79510,I79493);
nor I_4529 (I79527,I79462,I79510);
nor I_4530 (I79544,I79168,I79527);
DFFARX1 I_4531 (I79544,I2507,I79134,I79120,);
nor I_4532 (I79575,I79228,I79510);
nor I_4533 (I79108,I79423,I79575);
nor I_4534 (I79117,I79358,I79493);
nor I_4535 (I79105,I79228,I79493);
not I_4536 (I79661,I2514);
DFFARX1 I_4537 (I1086120,I2507,I79661,I79687,);
not I_4538 (I79695,I79687);
nand I_4539 (I79712,I1086135,I1086114);
and I_4540 (I79729,I79712,I1086117);
DFFARX1 I_4541 (I79729,I2507,I79661,I79755,);
DFFARX1 I_4542 (I1086138,I2507,I79661,I79772,);
and I_4543 (I79780,I79772,I1086117);
nor I_4544 (I79797,I79755,I79780);
DFFARX1 I_4545 (I79797,I2507,I79661,I79629,);
nand I_4546 (I79828,I79772,I1086117);
nand I_4547 (I79845,I79695,I79828);
not I_4548 (I79641,I79845);
DFFARX1 I_4549 (I1086114,I2507,I79661,I79885,);
DFFARX1 I_4550 (I79885,I2507,I79661,I79650,);
nand I_4551 (I79907,I1086126,I1086123);
and I_4552 (I79924,I79907,I1086129);
DFFARX1 I_4553 (I79924,I2507,I79661,I79950,);
DFFARX1 I_4554 (I79950,I2507,I79661,I79967,);
not I_4555 (I79653,I79967);
not I_4556 (I79989,I79950);
nand I_4557 (I79638,I79989,I79828);
nor I_4558 (I80020,I1086132,I1086123);
not I_4559 (I80037,I80020);
nor I_4560 (I80054,I79989,I80037);
nor I_4561 (I80071,I79695,I80054);
DFFARX1 I_4562 (I80071,I2507,I79661,I79647,);
nor I_4563 (I80102,I79755,I80037);
nor I_4564 (I79635,I79950,I80102);
nor I_4565 (I79644,I79885,I80020);
nor I_4566 (I79632,I79755,I80020);
not I_4567 (I80188,I2514);
DFFARX1 I_4568 (I867078,I2507,I80188,I80214,);
not I_4569 (I80222,I80214);
nand I_4570 (I80239,I867075,I867090);
and I_4571 (I80256,I80239,I867072);
DFFARX1 I_4572 (I80256,I2507,I80188,I80282,);
DFFARX1 I_4573 (I867069,I2507,I80188,I80299,);
and I_4574 (I80307,I80299,I867069);
nor I_4575 (I80324,I80282,I80307);
DFFARX1 I_4576 (I80324,I2507,I80188,I80156,);
nand I_4577 (I80355,I80299,I867069);
nand I_4578 (I80372,I80222,I80355);
not I_4579 (I80168,I80372);
DFFARX1 I_4580 (I867072,I2507,I80188,I80412,);
DFFARX1 I_4581 (I80412,I2507,I80188,I80177,);
nand I_4582 (I80434,I867084,I867075);
and I_4583 (I80451,I80434,I867087);
DFFARX1 I_4584 (I80451,I2507,I80188,I80477,);
DFFARX1 I_4585 (I80477,I2507,I80188,I80494,);
not I_4586 (I80180,I80494);
not I_4587 (I80516,I80477);
nand I_4588 (I80165,I80516,I80355);
nor I_4589 (I80547,I867081,I867075);
not I_4590 (I80564,I80547);
nor I_4591 (I80581,I80516,I80564);
nor I_4592 (I80598,I80222,I80581);
DFFARX1 I_4593 (I80598,I2507,I80188,I80174,);
nor I_4594 (I80629,I80282,I80564);
nor I_4595 (I80162,I80477,I80629);
nor I_4596 (I80171,I80412,I80547);
nor I_4597 (I80159,I80282,I80547);
not I_4598 (I80715,I2514);
DFFARX1 I_4599 (I293958,I2507,I80715,I80741,);
not I_4600 (I80749,I80741);
nand I_4601 (I80766,I293940,I293955);
and I_4602 (I80783,I80766,I293931);
DFFARX1 I_4603 (I80783,I2507,I80715,I80809,);
DFFARX1 I_4604 (I293934,I2507,I80715,I80826,);
and I_4605 (I80834,I80826,I293949);
nor I_4606 (I80851,I80809,I80834);
DFFARX1 I_4607 (I80851,I2507,I80715,I80683,);
nand I_4608 (I80882,I80826,I293949);
nand I_4609 (I80899,I80749,I80882);
not I_4610 (I80695,I80899);
DFFARX1 I_4611 (I293952,I2507,I80715,I80939,);
DFFARX1 I_4612 (I80939,I2507,I80715,I80704,);
nand I_4613 (I80961,I293931,I293943);
and I_4614 (I80978,I80961,I293937);
DFFARX1 I_4615 (I80978,I2507,I80715,I81004,);
DFFARX1 I_4616 (I81004,I2507,I80715,I81021,);
not I_4617 (I80707,I81021);
not I_4618 (I81043,I81004);
nand I_4619 (I80692,I81043,I80882);
nor I_4620 (I81074,I293946,I293943);
not I_4621 (I81091,I81074);
nor I_4622 (I81108,I81043,I81091);
nor I_4623 (I81125,I80749,I81108);
DFFARX1 I_4624 (I81125,I2507,I80715,I80701,);
nor I_4625 (I81156,I80809,I81091);
nor I_4626 (I80689,I81004,I81156);
nor I_4627 (I80698,I80939,I81074);
nor I_4628 (I80686,I80809,I81074);
not I_4629 (I81242,I2514);
DFFARX1 I_4630 (I508967,I2507,I81242,I81268,);
not I_4631 (I81276,I81268);
nand I_4632 (I81293,I508988,I508982);
and I_4633 (I81310,I81293,I508964);
DFFARX1 I_4634 (I81310,I2507,I81242,I81336,);
DFFARX1 I_4635 (I508967,I2507,I81242,I81353,);
and I_4636 (I81361,I81353,I508976);
nor I_4637 (I81378,I81336,I81361);
DFFARX1 I_4638 (I81378,I2507,I81242,I81210,);
nand I_4639 (I81409,I81353,I508976);
nand I_4640 (I81426,I81276,I81409);
not I_4641 (I81222,I81426);
DFFARX1 I_4642 (I508973,I2507,I81242,I81466,);
DFFARX1 I_4643 (I81466,I2507,I81242,I81231,);
nand I_4644 (I81488,I508979,I508970);
and I_4645 (I81505,I81488,I508964);
DFFARX1 I_4646 (I81505,I2507,I81242,I81531,);
DFFARX1 I_4647 (I81531,I2507,I81242,I81548,);
not I_4648 (I81234,I81548);
not I_4649 (I81570,I81531);
nand I_4650 (I81219,I81570,I81409);
nor I_4651 (I81601,I508985,I508970);
not I_4652 (I81618,I81601);
nor I_4653 (I81635,I81570,I81618);
nor I_4654 (I81652,I81276,I81635);
DFFARX1 I_4655 (I81652,I2507,I81242,I81228,);
nor I_4656 (I81683,I81336,I81618);
nor I_4657 (I81216,I81531,I81683);
nor I_4658 (I81225,I81466,I81601);
nor I_4659 (I81213,I81336,I81601);
not I_4660 (I81769,I2514);
DFFARX1 I_4661 (I468097,I2507,I81769,I81795,);
not I_4662 (I81803,I81795);
nand I_4663 (I81820,I468091,I468082);
and I_4664 (I81837,I81820,I468103);
DFFARX1 I_4665 (I81837,I2507,I81769,I81863,);
DFFARX1 I_4666 (I468085,I2507,I81769,I81880,);
and I_4667 (I81888,I81880,I468079);
nor I_4668 (I81905,I81863,I81888);
DFFARX1 I_4669 (I81905,I2507,I81769,I81737,);
nand I_4670 (I81936,I81880,I468079);
nand I_4671 (I81953,I81803,I81936);
not I_4672 (I81749,I81953);
DFFARX1 I_4673 (I468079,I2507,I81769,I81993,);
DFFARX1 I_4674 (I81993,I2507,I81769,I81758,);
nand I_4675 (I82015,I468106,I468088);
and I_4676 (I82032,I82015,I468094);
DFFARX1 I_4677 (I82032,I2507,I81769,I82058,);
DFFARX1 I_4678 (I82058,I2507,I81769,I82075,);
not I_4679 (I81761,I82075);
not I_4680 (I82097,I82058);
nand I_4681 (I81746,I82097,I81936);
nor I_4682 (I82128,I468100,I468088);
not I_4683 (I82145,I82128);
nor I_4684 (I82162,I82097,I82145);
nor I_4685 (I82179,I81803,I82162);
DFFARX1 I_4686 (I82179,I2507,I81769,I81755,);
nor I_4687 (I82210,I81863,I82145);
nor I_4688 (I81743,I82058,I82210);
nor I_4689 (I81752,I81993,I82128);
nor I_4690 (I81740,I81863,I82128);
not I_4691 (I82296,I2514);
DFFARX1 I_4692 (I329794,I2507,I82296,I82322,);
not I_4693 (I82330,I82322);
nand I_4694 (I82347,I329776,I329791);
and I_4695 (I82364,I82347,I329767);
DFFARX1 I_4696 (I82364,I2507,I82296,I82390,);
DFFARX1 I_4697 (I329770,I2507,I82296,I82407,);
and I_4698 (I82415,I82407,I329785);
nor I_4699 (I82432,I82390,I82415);
DFFARX1 I_4700 (I82432,I2507,I82296,I82264,);
nand I_4701 (I82463,I82407,I329785);
nand I_4702 (I82480,I82330,I82463);
not I_4703 (I82276,I82480);
DFFARX1 I_4704 (I329788,I2507,I82296,I82520,);
DFFARX1 I_4705 (I82520,I2507,I82296,I82285,);
nand I_4706 (I82542,I329767,I329779);
and I_4707 (I82559,I82542,I329773);
DFFARX1 I_4708 (I82559,I2507,I82296,I82585,);
DFFARX1 I_4709 (I82585,I2507,I82296,I82602,);
not I_4710 (I82288,I82602);
not I_4711 (I82624,I82585);
nand I_4712 (I82273,I82624,I82463);
nor I_4713 (I82655,I329782,I329779);
not I_4714 (I82672,I82655);
nor I_4715 (I82689,I82624,I82672);
nor I_4716 (I82706,I82330,I82689);
DFFARX1 I_4717 (I82706,I2507,I82296,I82282,);
nor I_4718 (I82737,I82390,I82672);
nor I_4719 (I82270,I82585,I82737);
nor I_4720 (I82279,I82520,I82655);
nor I_4721 (I82267,I82390,I82655);
not I_4722 (I82823,I2514);
DFFARX1 I_4723 (I1164728,I2507,I82823,I82849,);
not I_4724 (I82857,I82849);
nand I_4725 (I82874,I1164743,I1164722);
and I_4726 (I82891,I82874,I1164725);
DFFARX1 I_4727 (I82891,I2507,I82823,I82917,);
DFFARX1 I_4728 (I1164746,I2507,I82823,I82934,);
and I_4729 (I82942,I82934,I1164725);
nor I_4730 (I82959,I82917,I82942);
DFFARX1 I_4731 (I82959,I2507,I82823,I82791,);
nand I_4732 (I82990,I82934,I1164725);
nand I_4733 (I83007,I82857,I82990);
not I_4734 (I82803,I83007);
DFFARX1 I_4735 (I1164722,I2507,I82823,I83047,);
DFFARX1 I_4736 (I83047,I2507,I82823,I82812,);
nand I_4737 (I83069,I1164734,I1164731);
and I_4738 (I83086,I83069,I1164737);
DFFARX1 I_4739 (I83086,I2507,I82823,I83112,);
DFFARX1 I_4740 (I83112,I2507,I82823,I83129,);
not I_4741 (I82815,I83129);
not I_4742 (I83151,I83112);
nand I_4743 (I82800,I83151,I82990);
nor I_4744 (I83182,I1164740,I1164731);
not I_4745 (I83199,I83182);
nor I_4746 (I83216,I83151,I83199);
nor I_4747 (I83233,I82857,I83216);
DFFARX1 I_4748 (I83233,I2507,I82823,I82809,);
nor I_4749 (I83264,I82917,I83199);
nor I_4750 (I82797,I83112,I83264);
nor I_4751 (I82806,I83047,I83182);
nor I_4752 (I82794,I82917,I83182);
not I_4753 (I83350,I2514);
DFFARX1 I_4754 (I760202,I2507,I83350,I83376,);
not I_4755 (I83384,I83376);
nand I_4756 (I83401,I760193,I760211);
and I_4757 (I83418,I83401,I760190);
DFFARX1 I_4758 (I83418,I2507,I83350,I83444,);
DFFARX1 I_4759 (I760193,I2507,I83350,I83461,);
and I_4760 (I83469,I83461,I760196);
nor I_4761 (I83486,I83444,I83469);
DFFARX1 I_4762 (I83486,I2507,I83350,I83318,);
nand I_4763 (I83517,I83461,I760196);
nand I_4764 (I83534,I83384,I83517);
not I_4765 (I83330,I83534);
DFFARX1 I_4766 (I760190,I2507,I83350,I83574,);
DFFARX1 I_4767 (I83574,I2507,I83350,I83339,);
nand I_4768 (I83596,I760208,I760199);
and I_4769 (I83613,I83596,I760214);
DFFARX1 I_4770 (I83613,I2507,I83350,I83639,);
DFFARX1 I_4771 (I83639,I2507,I83350,I83656,);
not I_4772 (I83342,I83656);
not I_4773 (I83678,I83639);
nand I_4774 (I83327,I83678,I83517);
nor I_4775 (I83709,I760205,I760199);
not I_4776 (I83726,I83709);
nor I_4777 (I83743,I83678,I83726);
nor I_4778 (I83760,I83384,I83743);
DFFARX1 I_4779 (I83760,I2507,I83350,I83336,);
nor I_4780 (I83791,I83444,I83726);
nor I_4781 (I83324,I83639,I83791);
nor I_4782 (I83333,I83574,I83709);
nor I_4783 (I83321,I83444,I83709);
not I_4784 (I83877,I2514);
DFFARX1 I_4785 (I191297,I2507,I83877,I83903,);
not I_4786 (I83911,I83903);
nand I_4787 (I83928,I191291,I191285);
and I_4788 (I83945,I83928,I191306);
DFFARX1 I_4789 (I83945,I2507,I83877,I83971,);
DFFARX1 I_4790 (I191303,I2507,I83877,I83988,);
and I_4791 (I83996,I83988,I191300);
nor I_4792 (I84013,I83971,I83996);
DFFARX1 I_4793 (I84013,I2507,I83877,I83845,);
nand I_4794 (I84044,I83988,I191300);
nand I_4795 (I84061,I83911,I84044);
not I_4796 (I83857,I84061);
DFFARX1 I_4797 (I191285,I2507,I83877,I84101,);
DFFARX1 I_4798 (I84101,I2507,I83877,I83866,);
nand I_4799 (I84123,I191288,I191288);
and I_4800 (I84140,I84123,I191309);
DFFARX1 I_4801 (I84140,I2507,I83877,I84166,);
DFFARX1 I_4802 (I84166,I2507,I83877,I84183,);
not I_4803 (I83869,I84183);
not I_4804 (I84205,I84166);
nand I_4805 (I83854,I84205,I84044);
nor I_4806 (I84236,I191294,I191288);
not I_4807 (I84253,I84236);
nor I_4808 (I84270,I84205,I84253);
nor I_4809 (I84287,I83911,I84270);
DFFARX1 I_4810 (I84287,I2507,I83877,I83863,);
nor I_4811 (I84318,I83971,I84253);
nor I_4812 (I83851,I84166,I84318);
nor I_4813 (I83860,I84101,I84236);
nor I_4814 (I83848,I83971,I84236);
not I_4815 (I84404,I2514);
DFFARX1 I_4816 (I1091900,I2507,I84404,I84430,);
not I_4817 (I84438,I84430);
nand I_4818 (I84455,I1091915,I1091894);
and I_4819 (I84472,I84455,I1091897);
DFFARX1 I_4820 (I84472,I2507,I84404,I84498,);
DFFARX1 I_4821 (I1091918,I2507,I84404,I84515,);
and I_4822 (I84523,I84515,I1091897);
nor I_4823 (I84540,I84498,I84523);
DFFARX1 I_4824 (I84540,I2507,I84404,I84372,);
nand I_4825 (I84571,I84515,I1091897);
nand I_4826 (I84588,I84438,I84571);
not I_4827 (I84384,I84588);
DFFARX1 I_4828 (I1091894,I2507,I84404,I84628,);
DFFARX1 I_4829 (I84628,I2507,I84404,I84393,);
nand I_4830 (I84650,I1091906,I1091903);
and I_4831 (I84667,I84650,I1091909);
DFFARX1 I_4832 (I84667,I2507,I84404,I84693,);
DFFARX1 I_4833 (I84693,I2507,I84404,I84710,);
not I_4834 (I84396,I84710);
not I_4835 (I84732,I84693);
nand I_4836 (I84381,I84732,I84571);
nor I_4837 (I84763,I1091912,I1091903);
not I_4838 (I84780,I84763);
nor I_4839 (I84797,I84732,I84780);
nor I_4840 (I84814,I84438,I84797);
DFFARX1 I_4841 (I84814,I2507,I84404,I84390,);
nor I_4842 (I84845,I84498,I84780);
nor I_4843 (I84378,I84693,I84845);
nor I_4844 (I84387,I84628,I84763);
nor I_4845 (I84375,I84498,I84763);
not I_4846 (I84931,I2514);
DFFARX1 I_4847 (I1278473,I2507,I84931,I84957,);
not I_4848 (I84965,I84957);
nand I_4849 (I84982,I1278476,I1278470);
and I_4850 (I84999,I84982,I1278467);
DFFARX1 I_4851 (I84999,I2507,I84931,I85025,);
DFFARX1 I_4852 (I1278452,I2507,I84931,I85042,);
and I_4853 (I85050,I85042,I1278461);
nor I_4854 (I85067,I85025,I85050);
DFFARX1 I_4855 (I85067,I2507,I84931,I84899,);
nand I_4856 (I85098,I85042,I1278461);
nand I_4857 (I85115,I84965,I85098);
not I_4858 (I84911,I85115);
DFFARX1 I_4859 (I1278452,I2507,I84931,I85155,);
DFFARX1 I_4860 (I85155,I2507,I84931,I84920,);
nand I_4861 (I85177,I1278455,I1278458);
and I_4862 (I85194,I85177,I1278464);
DFFARX1 I_4863 (I85194,I2507,I84931,I85220,);
DFFARX1 I_4864 (I85220,I2507,I84931,I85237,);
not I_4865 (I84923,I85237);
not I_4866 (I85259,I85220);
nand I_4867 (I84908,I85259,I85098);
nor I_4868 (I85290,I1278455,I1278458);
not I_4869 (I85307,I85290);
nor I_4870 (I85324,I85259,I85307);
nor I_4871 (I85341,I84965,I85324);
DFFARX1 I_4872 (I85341,I2507,I84931,I84917,);
nor I_4873 (I85372,I85025,I85307);
nor I_4874 (I84905,I85220,I85372);
nor I_4875 (I84914,I85155,I85290);
nor I_4876 (I84902,I85025,I85290);
not I_4877 (I85458,I2514);
DFFARX1 I_4878 (I390305,I2507,I85458,I85484,);
not I_4879 (I85492,I85484);
nand I_4880 (I85509,I390299,I390290);
and I_4881 (I85526,I85509,I390311);
DFFARX1 I_4882 (I85526,I2507,I85458,I85552,);
DFFARX1 I_4883 (I390293,I2507,I85458,I85569,);
and I_4884 (I85577,I85569,I390287);
nor I_4885 (I85594,I85552,I85577);
DFFARX1 I_4886 (I85594,I2507,I85458,I85426,);
nand I_4887 (I85625,I85569,I390287);
nand I_4888 (I85642,I85492,I85625);
not I_4889 (I85438,I85642);
DFFARX1 I_4890 (I390287,I2507,I85458,I85682,);
DFFARX1 I_4891 (I85682,I2507,I85458,I85447,);
nand I_4892 (I85704,I390314,I390296);
and I_4893 (I85721,I85704,I390302);
DFFARX1 I_4894 (I85721,I2507,I85458,I85747,);
DFFARX1 I_4895 (I85747,I2507,I85458,I85764,);
not I_4896 (I85450,I85764);
not I_4897 (I85786,I85747);
nand I_4898 (I85435,I85786,I85625);
nor I_4899 (I85817,I390308,I390296);
not I_4900 (I85834,I85817);
nor I_4901 (I85851,I85786,I85834);
nor I_4902 (I85868,I85492,I85851);
DFFARX1 I_4903 (I85868,I2507,I85458,I85444,);
nor I_4904 (I85899,I85552,I85834);
nor I_4905 (I85432,I85747,I85899);
nor I_4906 (I85441,I85682,I85817);
nor I_4907 (I85429,I85552,I85817);
not I_4908 (I85985,I2514);
DFFARX1 I_4909 (I607607,I2507,I85985,I86011,);
not I_4910 (I86019,I86011);
nand I_4911 (I86036,I607619,I607604);
and I_4912 (I86053,I86036,I607598);
DFFARX1 I_4913 (I86053,I2507,I85985,I86079,);
DFFARX1 I_4914 (I607613,I2507,I85985,I86096,);
and I_4915 (I86104,I86096,I607601);
nor I_4916 (I86121,I86079,I86104);
DFFARX1 I_4917 (I86121,I2507,I85985,I85953,);
nand I_4918 (I86152,I86096,I607601);
nand I_4919 (I86169,I86019,I86152);
not I_4920 (I85965,I86169);
DFFARX1 I_4921 (I607610,I2507,I85985,I86209,);
DFFARX1 I_4922 (I86209,I2507,I85985,I85974,);
nand I_4923 (I86231,I607616,I607622);
and I_4924 (I86248,I86231,I607598);
DFFARX1 I_4925 (I86248,I2507,I85985,I86274,);
DFFARX1 I_4926 (I86274,I2507,I85985,I86291,);
not I_4927 (I85977,I86291);
not I_4928 (I86313,I86274);
nand I_4929 (I85962,I86313,I86152);
nor I_4930 (I86344,I607601,I607622);
not I_4931 (I86361,I86344);
nor I_4932 (I86378,I86313,I86361);
nor I_4933 (I86395,I86019,I86378);
DFFARX1 I_4934 (I86395,I2507,I85985,I85971,);
nor I_4935 (I86426,I86079,I86361);
nor I_4936 (I85959,I86274,I86426);
nor I_4937 (I85968,I86209,I86344);
nor I_4938 (I85956,I86079,I86344);
not I_4939 (I86512,I2514);
DFFARX1 I_4940 (I1147388,I2507,I86512,I86538,);
not I_4941 (I86546,I86538);
nand I_4942 (I86563,I1147403,I1147382);
and I_4943 (I86580,I86563,I1147385);
DFFARX1 I_4944 (I86580,I2507,I86512,I86606,);
DFFARX1 I_4945 (I1147406,I2507,I86512,I86623,);
and I_4946 (I86631,I86623,I1147385);
nor I_4947 (I86648,I86606,I86631);
DFFARX1 I_4948 (I86648,I2507,I86512,I86480,);
nand I_4949 (I86679,I86623,I1147385);
nand I_4950 (I86696,I86546,I86679);
not I_4951 (I86492,I86696);
DFFARX1 I_4952 (I1147382,I2507,I86512,I86736,);
DFFARX1 I_4953 (I86736,I2507,I86512,I86501,);
nand I_4954 (I86758,I1147394,I1147391);
and I_4955 (I86775,I86758,I1147397);
DFFARX1 I_4956 (I86775,I2507,I86512,I86801,);
DFFARX1 I_4957 (I86801,I2507,I86512,I86818,);
not I_4958 (I86504,I86818);
not I_4959 (I86840,I86801);
nand I_4960 (I86489,I86840,I86679);
nor I_4961 (I86871,I1147400,I1147391);
not I_4962 (I86888,I86871);
nor I_4963 (I86905,I86840,I86888);
nor I_4964 (I86922,I86546,I86905);
DFFARX1 I_4965 (I86922,I2507,I86512,I86498,);
nor I_4966 (I86953,I86606,I86888);
nor I_4967 (I86486,I86801,I86953);
nor I_4968 (I86495,I86736,I86871);
nor I_4969 (I86483,I86606,I86871);
not I_4970 (I87039,I2514);
DFFARX1 I_4971 (I1151434,I2507,I87039,I87065,);
not I_4972 (I87073,I87065);
nand I_4973 (I87090,I1151449,I1151428);
and I_4974 (I87107,I87090,I1151431);
DFFARX1 I_4975 (I87107,I2507,I87039,I87133,);
DFFARX1 I_4976 (I1151452,I2507,I87039,I87150,);
and I_4977 (I87158,I87150,I1151431);
nor I_4978 (I87175,I87133,I87158);
DFFARX1 I_4979 (I87175,I2507,I87039,I87007,);
nand I_4980 (I87206,I87150,I1151431);
nand I_4981 (I87223,I87073,I87206);
not I_4982 (I87019,I87223);
DFFARX1 I_4983 (I1151428,I2507,I87039,I87263,);
DFFARX1 I_4984 (I87263,I2507,I87039,I87028,);
nand I_4985 (I87285,I1151440,I1151437);
and I_4986 (I87302,I87285,I1151443);
DFFARX1 I_4987 (I87302,I2507,I87039,I87328,);
DFFARX1 I_4988 (I87328,I2507,I87039,I87345,);
not I_4989 (I87031,I87345);
not I_4990 (I87367,I87328);
nand I_4991 (I87016,I87367,I87206);
nor I_4992 (I87398,I1151446,I1151437);
not I_4993 (I87415,I87398);
nor I_4994 (I87432,I87367,I87415);
nor I_4995 (I87449,I87073,I87432);
DFFARX1 I_4996 (I87449,I2507,I87039,I87025,);
nor I_4997 (I87480,I87133,I87415);
nor I_4998 (I87013,I87328,I87480);
nor I_4999 (I87022,I87263,I87398);
nor I_5000 (I87010,I87133,I87398);
not I_5001 (I87566,I2514);
DFFARX1 I_5002 (I1252584,I2507,I87566,I87592,);
not I_5003 (I87600,I87592);
nand I_5004 (I87617,I1252578,I1252599);
and I_5005 (I87634,I87617,I1252590);
DFFARX1 I_5006 (I87634,I2507,I87566,I87660,);
DFFARX1 I_5007 (I1252581,I2507,I87566,I87677,);
and I_5008 (I87685,I87677,I1252593);
nor I_5009 (I87702,I87660,I87685);
DFFARX1 I_5010 (I87702,I2507,I87566,I87534,);
nand I_5011 (I87733,I87677,I1252593);
nand I_5012 (I87750,I87600,I87733);
not I_5013 (I87546,I87750);
DFFARX1 I_5014 (I1252581,I2507,I87566,I87790,);
DFFARX1 I_5015 (I87790,I2507,I87566,I87555,);
nand I_5016 (I87812,I1252602,I1252587);
and I_5017 (I87829,I87812,I1252578);
DFFARX1 I_5018 (I87829,I2507,I87566,I87855,);
DFFARX1 I_5019 (I87855,I2507,I87566,I87872,);
not I_5020 (I87558,I87872);
not I_5021 (I87894,I87855);
nand I_5022 (I87543,I87894,I87733);
nor I_5023 (I87925,I1252596,I1252587);
not I_5024 (I87942,I87925);
nor I_5025 (I87959,I87894,I87942);
nor I_5026 (I87976,I87600,I87959);
DFFARX1 I_5027 (I87976,I2507,I87566,I87552,);
nor I_5028 (I88007,I87660,I87942);
nor I_5029 (I87540,I87855,I88007);
nor I_5030 (I87549,I87790,I87925);
nor I_5031 (I87537,I87660,I87925);
not I_5032 (I88093,I2514);
DFFARX1 I_5033 (I1336264,I2507,I88093,I88119,);
not I_5034 (I88127,I88119);
nand I_5035 (I88144,I1336258,I1336279);
and I_5036 (I88161,I88144,I1336255);
DFFARX1 I_5037 (I88161,I2507,I88093,I88187,);
DFFARX1 I_5038 (I1336276,I2507,I88093,I88204,);
and I_5039 (I88212,I88204,I1336273);
nor I_5040 (I88229,I88187,I88212);
DFFARX1 I_5041 (I88229,I2507,I88093,I88061,);
nand I_5042 (I88260,I88204,I1336273);
nand I_5043 (I88277,I88127,I88260);
not I_5044 (I88073,I88277);
DFFARX1 I_5045 (I1336261,I2507,I88093,I88317,);
DFFARX1 I_5046 (I88317,I2507,I88093,I88082,);
nand I_5047 (I88339,I1336270,I1336267);
and I_5048 (I88356,I88339,I1336252);
DFFARX1 I_5049 (I88356,I2507,I88093,I88382,);
DFFARX1 I_5050 (I88382,I2507,I88093,I88399,);
not I_5051 (I88085,I88399);
not I_5052 (I88421,I88382);
nand I_5053 (I88070,I88421,I88260);
nor I_5054 (I88452,I1336252,I1336267);
not I_5055 (I88469,I88452);
nor I_5056 (I88486,I88421,I88469);
nor I_5057 (I88503,I88127,I88486);
DFFARX1 I_5058 (I88503,I2507,I88093,I88079,);
nor I_5059 (I88534,I88187,I88469);
nor I_5060 (I88067,I88382,I88534);
nor I_5061 (I88076,I88317,I88452);
nor I_5062 (I88064,I88187,I88452);
not I_5063 (I88620,I2514);
DFFARX1 I_5064 (I533957,I2507,I88620,I88646,);
not I_5065 (I88654,I88646);
nand I_5066 (I88671,I533978,I533972);
and I_5067 (I88688,I88671,I533954);
DFFARX1 I_5068 (I88688,I2507,I88620,I88714,);
DFFARX1 I_5069 (I533957,I2507,I88620,I88731,);
and I_5070 (I88739,I88731,I533966);
nor I_5071 (I88756,I88714,I88739);
DFFARX1 I_5072 (I88756,I2507,I88620,I88588,);
nand I_5073 (I88787,I88731,I533966);
nand I_5074 (I88804,I88654,I88787);
not I_5075 (I88600,I88804);
DFFARX1 I_5076 (I533963,I2507,I88620,I88844,);
DFFARX1 I_5077 (I88844,I2507,I88620,I88609,);
nand I_5078 (I88866,I533969,I533960);
and I_5079 (I88883,I88866,I533954);
DFFARX1 I_5080 (I88883,I2507,I88620,I88909,);
DFFARX1 I_5081 (I88909,I2507,I88620,I88926,);
not I_5082 (I88612,I88926);
not I_5083 (I88948,I88909);
nand I_5084 (I88597,I88948,I88787);
nor I_5085 (I88979,I533975,I533960);
not I_5086 (I88996,I88979);
nor I_5087 (I89013,I88948,I88996);
nor I_5088 (I89030,I88654,I89013);
DFFARX1 I_5089 (I89030,I2507,I88620,I88606,);
nor I_5090 (I89061,I88714,I88996);
nor I_5091 (I88594,I88909,I89061);
nor I_5092 (I88603,I88844,I88979);
nor I_5093 (I88591,I88714,I88979);
not I_5094 (I89147,I2514);
DFFARX1 I_5095 (I663098,I2507,I89147,I89173,);
not I_5096 (I89181,I89173);
nand I_5097 (I89198,I663089,I663107);
and I_5098 (I89215,I89198,I663086);
DFFARX1 I_5099 (I89215,I2507,I89147,I89241,);
DFFARX1 I_5100 (I663089,I2507,I89147,I89258,);
and I_5101 (I89266,I89258,I663092);
nor I_5102 (I89283,I89241,I89266);
DFFARX1 I_5103 (I89283,I2507,I89147,I89115,);
nand I_5104 (I89314,I89258,I663092);
nand I_5105 (I89331,I89181,I89314);
not I_5106 (I89127,I89331);
DFFARX1 I_5107 (I663086,I2507,I89147,I89371,);
DFFARX1 I_5108 (I89371,I2507,I89147,I89136,);
nand I_5109 (I89393,I663104,I663095);
and I_5110 (I89410,I89393,I663110);
DFFARX1 I_5111 (I89410,I2507,I89147,I89436,);
DFFARX1 I_5112 (I89436,I2507,I89147,I89453,);
not I_5113 (I89139,I89453);
not I_5114 (I89475,I89436);
nand I_5115 (I89124,I89475,I89314);
nor I_5116 (I89506,I663101,I663095);
not I_5117 (I89523,I89506);
nor I_5118 (I89540,I89475,I89523);
nor I_5119 (I89557,I89181,I89540);
DFFARX1 I_5120 (I89557,I2507,I89147,I89133,);
nor I_5121 (I89588,I89241,I89523);
nor I_5122 (I89121,I89436,I89588);
nor I_5123 (I89130,I89371,I89506);
nor I_5124 (I89118,I89241,I89506);
not I_5125 (I89674,I2514);
DFFARX1 I_5126 (I467009,I2507,I89674,I89700,);
not I_5127 (I89708,I89700);
nand I_5128 (I89725,I467003,I466994);
and I_5129 (I89742,I89725,I467015);
DFFARX1 I_5130 (I89742,I2507,I89674,I89768,);
DFFARX1 I_5131 (I466997,I2507,I89674,I89785,);
and I_5132 (I89793,I89785,I466991);
nor I_5133 (I89810,I89768,I89793);
DFFARX1 I_5134 (I89810,I2507,I89674,I89642,);
nand I_5135 (I89841,I89785,I466991);
nand I_5136 (I89858,I89708,I89841);
not I_5137 (I89654,I89858);
DFFARX1 I_5138 (I466991,I2507,I89674,I89898,);
DFFARX1 I_5139 (I89898,I2507,I89674,I89663,);
nand I_5140 (I89920,I467018,I467000);
and I_5141 (I89937,I89920,I467006);
DFFARX1 I_5142 (I89937,I2507,I89674,I89963,);
DFFARX1 I_5143 (I89963,I2507,I89674,I89980,);
not I_5144 (I89666,I89980);
not I_5145 (I90002,I89963);
nand I_5146 (I89651,I90002,I89841);
nor I_5147 (I90033,I467012,I467000);
not I_5148 (I90050,I90033);
nor I_5149 (I90067,I90002,I90050);
nor I_5150 (I90084,I89708,I90067);
DFFARX1 I_5151 (I90084,I2507,I89674,I89660,);
nor I_5152 (I90115,I89768,I90050);
nor I_5153 (I89648,I89963,I90115);
nor I_5154 (I89657,I89898,I90033);
nor I_5155 (I89645,I89768,I90033);
not I_5156 (I90201,I2514);
DFFARX1 I_5157 (I38020,I2507,I90201,I90227,);
not I_5158 (I90235,I90227);
nand I_5159 (I90252,I38008,I38014);
and I_5160 (I90269,I90252,I38017);
DFFARX1 I_5161 (I90269,I2507,I90201,I90295,);
DFFARX1 I_5162 (I37999,I2507,I90201,I90312,);
and I_5163 (I90320,I90312,I38005);
nor I_5164 (I90337,I90295,I90320);
DFFARX1 I_5165 (I90337,I2507,I90201,I90169,);
nand I_5166 (I90368,I90312,I38005);
nand I_5167 (I90385,I90235,I90368);
not I_5168 (I90181,I90385);
DFFARX1 I_5169 (I37999,I2507,I90201,I90425,);
DFFARX1 I_5170 (I90425,I2507,I90201,I90190,);
nand I_5171 (I90447,I38002,I37996);
and I_5172 (I90464,I90447,I38011);
DFFARX1 I_5173 (I90464,I2507,I90201,I90490,);
DFFARX1 I_5174 (I90490,I2507,I90201,I90507,);
not I_5175 (I90193,I90507);
not I_5176 (I90529,I90490);
nand I_5177 (I90178,I90529,I90368);
nor I_5178 (I90560,I37996,I37996);
not I_5179 (I90577,I90560);
nor I_5180 (I90594,I90529,I90577);
nor I_5181 (I90611,I90235,I90594);
DFFARX1 I_5182 (I90611,I2507,I90201,I90187,);
nor I_5183 (I90642,I90295,I90577);
nor I_5184 (I90175,I90490,I90642);
nor I_5185 (I90184,I90425,I90560);
nor I_5186 (I90172,I90295,I90560);
not I_5187 (I90728,I2514);
DFFARX1 I_5188 (I905668,I2507,I90728,I90754,);
not I_5189 (I90762,I90754);
nand I_5190 (I90779,I905686,I905680);
and I_5191 (I90796,I90779,I905659);
DFFARX1 I_5192 (I90796,I2507,I90728,I90822,);
DFFARX1 I_5193 (I905677,I2507,I90728,I90839,);
and I_5194 (I90847,I90839,I905662);
nor I_5195 (I90864,I90822,I90847);
DFFARX1 I_5196 (I90864,I2507,I90728,I90696,);
nand I_5197 (I90895,I90839,I905662);
nand I_5198 (I90912,I90762,I90895);
not I_5199 (I90708,I90912);
DFFARX1 I_5200 (I905674,I2507,I90728,I90952,);
DFFARX1 I_5201 (I90952,I2507,I90728,I90717,);
nand I_5202 (I90974,I905683,I905671);
and I_5203 (I90991,I90974,I905665);
DFFARX1 I_5204 (I90991,I2507,I90728,I91017,);
DFFARX1 I_5205 (I91017,I2507,I90728,I91034,);
not I_5206 (I90720,I91034);
not I_5207 (I91056,I91017);
nand I_5208 (I90705,I91056,I90895);
nor I_5209 (I91087,I905659,I905671);
not I_5210 (I91104,I91087);
nor I_5211 (I91121,I91056,I91104);
nor I_5212 (I91138,I90762,I91121);
DFFARX1 I_5213 (I91138,I2507,I90728,I90714,);
nor I_5214 (I91169,I90822,I91104);
nor I_5215 (I90702,I91017,I91169);
nor I_5216 (I90711,I90952,I91087);
nor I_5217 (I90699,I90822,I91087);
not I_5218 (I91255,I2514);
DFFARX1 I_5219 (I1247688,I2507,I91255,I91281,);
not I_5220 (I91289,I91281);
nand I_5221 (I91306,I1247682,I1247703);
and I_5222 (I91323,I91306,I1247694);
DFFARX1 I_5223 (I91323,I2507,I91255,I91349,);
DFFARX1 I_5224 (I1247685,I2507,I91255,I91366,);
and I_5225 (I91374,I91366,I1247697);
nor I_5226 (I91391,I91349,I91374);
DFFARX1 I_5227 (I91391,I2507,I91255,I91223,);
nand I_5228 (I91422,I91366,I1247697);
nand I_5229 (I91439,I91289,I91422);
not I_5230 (I91235,I91439);
DFFARX1 I_5231 (I1247685,I2507,I91255,I91479,);
DFFARX1 I_5232 (I91479,I2507,I91255,I91244,);
nand I_5233 (I91501,I1247706,I1247691);
and I_5234 (I91518,I91501,I1247682);
DFFARX1 I_5235 (I91518,I2507,I91255,I91544,);
DFFARX1 I_5236 (I91544,I2507,I91255,I91561,);
not I_5237 (I91247,I91561);
not I_5238 (I91583,I91544);
nand I_5239 (I91232,I91583,I91422);
nor I_5240 (I91614,I1247700,I1247691);
not I_5241 (I91631,I91614);
nor I_5242 (I91648,I91583,I91631);
nor I_5243 (I91665,I91289,I91648);
DFFARX1 I_5244 (I91665,I2507,I91255,I91241,);
nor I_5245 (I91696,I91349,I91631);
nor I_5246 (I91229,I91544,I91696);
nor I_5247 (I91238,I91479,I91614);
nor I_5248 (I91226,I91349,I91614);
not I_5249 (I91782,I2514);
DFFARX1 I_5250 (I152622,I2507,I91782,I91808,);
not I_5251 (I91816,I91808);
nand I_5252 (I91833,I152616,I152610);
and I_5253 (I91850,I91833,I152631);
DFFARX1 I_5254 (I91850,I2507,I91782,I91876,);
DFFARX1 I_5255 (I152628,I2507,I91782,I91893,);
and I_5256 (I91901,I91893,I152625);
nor I_5257 (I91918,I91876,I91901);
DFFARX1 I_5258 (I91918,I2507,I91782,I91750,);
nand I_5259 (I91949,I91893,I152625);
nand I_5260 (I91966,I91816,I91949);
not I_5261 (I91762,I91966);
DFFARX1 I_5262 (I152610,I2507,I91782,I92006,);
DFFARX1 I_5263 (I92006,I2507,I91782,I91771,);
nand I_5264 (I92028,I152613,I152613);
and I_5265 (I92045,I92028,I152634);
DFFARX1 I_5266 (I92045,I2507,I91782,I92071,);
DFFARX1 I_5267 (I92071,I2507,I91782,I92088,);
not I_5268 (I91774,I92088);
not I_5269 (I92110,I92071);
nand I_5270 (I91759,I92110,I91949);
nor I_5271 (I92141,I152619,I152613);
not I_5272 (I92158,I92141);
nor I_5273 (I92175,I92110,I92158);
nor I_5274 (I92192,I91816,I92175);
DFFARX1 I_5275 (I92192,I2507,I91782,I91768,);
nor I_5276 (I92223,I91876,I92158);
nor I_5277 (I91756,I92071,I92223);
nor I_5278 (I91765,I92006,I92141);
nor I_5279 (I91753,I91876,I92141);
not I_5280 (I92309,I2514);
DFFARX1 I_5281 (I747486,I2507,I92309,I92335,);
not I_5282 (I92343,I92335);
nand I_5283 (I92360,I747477,I747495);
and I_5284 (I92377,I92360,I747474);
DFFARX1 I_5285 (I92377,I2507,I92309,I92403,);
DFFARX1 I_5286 (I747477,I2507,I92309,I92420,);
and I_5287 (I92428,I92420,I747480);
nor I_5288 (I92445,I92403,I92428);
DFFARX1 I_5289 (I92445,I2507,I92309,I92277,);
nand I_5290 (I92476,I92420,I747480);
nand I_5291 (I92493,I92343,I92476);
not I_5292 (I92289,I92493);
DFFARX1 I_5293 (I747474,I2507,I92309,I92533,);
DFFARX1 I_5294 (I92533,I2507,I92309,I92298,);
nand I_5295 (I92555,I747492,I747483);
and I_5296 (I92572,I92555,I747498);
DFFARX1 I_5297 (I92572,I2507,I92309,I92598,);
DFFARX1 I_5298 (I92598,I2507,I92309,I92615,);
not I_5299 (I92301,I92615);
not I_5300 (I92637,I92598);
nand I_5301 (I92286,I92637,I92476);
nor I_5302 (I92668,I747489,I747483);
not I_5303 (I92685,I92668);
nor I_5304 (I92702,I92637,I92685);
nor I_5305 (I92719,I92343,I92702);
DFFARX1 I_5306 (I92719,I2507,I92309,I92295,);
nor I_5307 (I92750,I92403,I92685);
nor I_5308 (I92283,I92598,I92750);
nor I_5309 (I92292,I92533,I92668);
nor I_5310 (I92280,I92403,I92668);
not I_5311 (I92836,I2514);
DFFARX1 I_5312 (I1234088,I2507,I92836,I92862,);
not I_5313 (I92870,I92862);
nand I_5314 (I92887,I1234082,I1234103);
and I_5315 (I92904,I92887,I1234094);
DFFARX1 I_5316 (I92904,I2507,I92836,I92930,);
DFFARX1 I_5317 (I1234085,I2507,I92836,I92947,);
and I_5318 (I92955,I92947,I1234097);
nor I_5319 (I92972,I92930,I92955);
DFFARX1 I_5320 (I92972,I2507,I92836,I92804,);
nand I_5321 (I93003,I92947,I1234097);
nand I_5322 (I93020,I92870,I93003);
not I_5323 (I92816,I93020);
DFFARX1 I_5324 (I1234085,I2507,I92836,I93060,);
DFFARX1 I_5325 (I93060,I2507,I92836,I92825,);
nand I_5326 (I93082,I1234106,I1234091);
and I_5327 (I93099,I93082,I1234082);
DFFARX1 I_5328 (I93099,I2507,I92836,I93125,);
DFFARX1 I_5329 (I93125,I2507,I92836,I93142,);
not I_5330 (I92828,I93142);
not I_5331 (I93164,I93125);
nand I_5332 (I92813,I93164,I93003);
nor I_5333 (I93195,I1234100,I1234091);
not I_5334 (I93212,I93195);
nor I_5335 (I93229,I93164,I93212);
nor I_5336 (I93246,I92870,I93229);
DFFARX1 I_5337 (I93246,I2507,I92836,I92822,);
nor I_5338 (I93277,I92930,I93212);
nor I_5339 (I92810,I93125,I93277);
nor I_5340 (I92819,I93060,I93195);
nor I_5341 (I92807,I92930,I93195);
not I_5342 (I93363,I2514);
DFFARX1 I_5343 (I246037,I2507,I93363,I93389,);
not I_5344 (I93397,I93389);
nand I_5345 (I93414,I246031,I246025);
and I_5346 (I93431,I93414,I246046);
DFFARX1 I_5347 (I93431,I2507,I93363,I93457,);
DFFARX1 I_5348 (I246043,I2507,I93363,I93474,);
and I_5349 (I93482,I93474,I246040);
nor I_5350 (I93499,I93457,I93482);
DFFARX1 I_5351 (I93499,I2507,I93363,I93331,);
nand I_5352 (I93530,I93474,I246040);
nand I_5353 (I93547,I93397,I93530);
not I_5354 (I93343,I93547);
DFFARX1 I_5355 (I246025,I2507,I93363,I93587,);
DFFARX1 I_5356 (I93587,I2507,I93363,I93352,);
nand I_5357 (I93609,I246028,I246028);
and I_5358 (I93626,I93609,I246049);
DFFARX1 I_5359 (I93626,I2507,I93363,I93652,);
DFFARX1 I_5360 (I93652,I2507,I93363,I93669,);
not I_5361 (I93355,I93669);
not I_5362 (I93691,I93652);
nand I_5363 (I93340,I93691,I93530);
nor I_5364 (I93722,I246034,I246028);
not I_5365 (I93739,I93722);
nor I_5366 (I93756,I93691,I93739);
nor I_5367 (I93773,I93397,I93756);
DFFARX1 I_5368 (I93773,I2507,I93363,I93349,);
nor I_5369 (I93804,I93457,I93739);
nor I_5370 (I93337,I93652,I93804);
nor I_5371 (I93346,I93587,I93722);
nor I_5372 (I93334,I93457,I93722);
not I_5373 (I93890,I2514);
DFFARX1 I_5374 (I895978,I2507,I93890,I93916,);
not I_5375 (I93924,I93916);
nand I_5376 (I93941,I895996,I895990);
and I_5377 (I93958,I93941,I895969);
DFFARX1 I_5378 (I93958,I2507,I93890,I93984,);
DFFARX1 I_5379 (I895987,I2507,I93890,I94001,);
and I_5380 (I94009,I94001,I895972);
nor I_5381 (I94026,I93984,I94009);
DFFARX1 I_5382 (I94026,I2507,I93890,I93858,);
nand I_5383 (I94057,I94001,I895972);
nand I_5384 (I94074,I93924,I94057);
not I_5385 (I93870,I94074);
DFFARX1 I_5386 (I895984,I2507,I93890,I94114,);
DFFARX1 I_5387 (I94114,I2507,I93890,I93879,);
nand I_5388 (I94136,I895993,I895981);
and I_5389 (I94153,I94136,I895975);
DFFARX1 I_5390 (I94153,I2507,I93890,I94179,);
DFFARX1 I_5391 (I94179,I2507,I93890,I94196,);
not I_5392 (I93882,I94196);
not I_5393 (I94218,I94179);
nand I_5394 (I93867,I94218,I94057);
nor I_5395 (I94249,I895969,I895981);
not I_5396 (I94266,I94249);
nor I_5397 (I94283,I94218,I94266);
nor I_5398 (I94300,I93924,I94283);
DFFARX1 I_5399 (I94300,I2507,I93890,I93876,);
nor I_5400 (I94331,I93984,I94266);
nor I_5401 (I93864,I94179,I94331);
nor I_5402 (I93873,I94114,I94249);
nor I_5403 (I93861,I93984,I94249);
not I_5404 (I94417,I2514);
DFFARX1 I_5405 (I955410,I2507,I94417,I94443,);
not I_5406 (I94451,I94443);
nand I_5407 (I94468,I955428,I955422);
and I_5408 (I94485,I94468,I955401);
DFFARX1 I_5409 (I94485,I2507,I94417,I94511,);
DFFARX1 I_5410 (I955419,I2507,I94417,I94528,);
and I_5411 (I94536,I94528,I955404);
nor I_5412 (I94553,I94511,I94536);
DFFARX1 I_5413 (I94553,I2507,I94417,I94385,);
nand I_5414 (I94584,I94528,I955404);
nand I_5415 (I94601,I94451,I94584);
not I_5416 (I94397,I94601);
DFFARX1 I_5417 (I955416,I2507,I94417,I94641,);
DFFARX1 I_5418 (I94641,I2507,I94417,I94406,);
nand I_5419 (I94663,I955425,I955413);
and I_5420 (I94680,I94663,I955407);
DFFARX1 I_5421 (I94680,I2507,I94417,I94706,);
DFFARX1 I_5422 (I94706,I2507,I94417,I94723,);
not I_5423 (I94409,I94723);
not I_5424 (I94745,I94706);
nand I_5425 (I94394,I94745,I94584);
nor I_5426 (I94776,I955401,I955413);
not I_5427 (I94793,I94776);
nor I_5428 (I94810,I94745,I94793);
nor I_5429 (I94827,I94451,I94810);
DFFARX1 I_5430 (I94827,I2507,I94417,I94403,);
nor I_5431 (I94858,I94511,I94793);
nor I_5432 (I94391,I94706,I94858);
nor I_5433 (I94400,I94641,I94776);
nor I_5434 (I94388,I94511,I94776);
not I_5435 (I94944,I2514);
DFFARX1 I_5436 (I553853,I2507,I94944,I94970,);
not I_5437 (I94978,I94970);
nand I_5438 (I94995,I553865,I553850);
and I_5439 (I95012,I94995,I553844);
DFFARX1 I_5440 (I95012,I2507,I94944,I95038,);
DFFARX1 I_5441 (I553859,I2507,I94944,I95055,);
and I_5442 (I95063,I95055,I553847);
nor I_5443 (I95080,I95038,I95063);
DFFARX1 I_5444 (I95080,I2507,I94944,I94912,);
nand I_5445 (I95111,I95055,I553847);
nand I_5446 (I95128,I94978,I95111);
not I_5447 (I94924,I95128);
DFFARX1 I_5448 (I553856,I2507,I94944,I95168,);
DFFARX1 I_5449 (I95168,I2507,I94944,I94933,);
nand I_5450 (I95190,I553862,I553868);
and I_5451 (I95207,I95190,I553844);
DFFARX1 I_5452 (I95207,I2507,I94944,I95233,);
DFFARX1 I_5453 (I95233,I2507,I94944,I95250,);
not I_5454 (I94936,I95250);
not I_5455 (I95272,I95233);
nand I_5456 (I94921,I95272,I95111);
nor I_5457 (I95303,I553847,I553868);
not I_5458 (I95320,I95303);
nor I_5459 (I95337,I95272,I95320);
nor I_5460 (I95354,I94978,I95337);
DFFARX1 I_5461 (I95354,I2507,I94944,I94930,);
nor I_5462 (I95385,I95038,I95320);
nor I_5463 (I94918,I95233,I95385);
nor I_5464 (I94927,I95168,I95303);
nor I_5465 (I94915,I95038,I95303);
not I_5466 (I95471,I2514);
DFFARX1 I_5467 (I272878,I2507,I95471,I95497,);
not I_5468 (I95505,I95497);
nand I_5469 (I95522,I272860,I272875);
and I_5470 (I95539,I95522,I272851);
DFFARX1 I_5471 (I95539,I2507,I95471,I95565,);
DFFARX1 I_5472 (I272854,I2507,I95471,I95582,);
and I_5473 (I95590,I95582,I272869);
nor I_5474 (I95607,I95565,I95590);
DFFARX1 I_5475 (I95607,I2507,I95471,I95439,);
nand I_5476 (I95638,I95582,I272869);
nand I_5477 (I95655,I95505,I95638);
not I_5478 (I95451,I95655);
DFFARX1 I_5479 (I272872,I2507,I95471,I95695,);
DFFARX1 I_5480 (I95695,I2507,I95471,I95460,);
nand I_5481 (I95717,I272851,I272863);
and I_5482 (I95734,I95717,I272857);
DFFARX1 I_5483 (I95734,I2507,I95471,I95760,);
DFFARX1 I_5484 (I95760,I2507,I95471,I95777,);
not I_5485 (I95463,I95777);
not I_5486 (I95799,I95760);
nand I_5487 (I95448,I95799,I95638);
nor I_5488 (I95830,I272866,I272863);
not I_5489 (I95847,I95830);
nor I_5490 (I95864,I95799,I95847);
nor I_5491 (I95881,I95505,I95864);
DFFARX1 I_5492 (I95881,I2507,I95471,I95457,);
nor I_5493 (I95912,I95565,I95847);
nor I_5494 (I95445,I95760,I95912);
nor I_5495 (I95454,I95695,I95830);
nor I_5496 (I95442,I95565,I95830);
not I_5497 (I95998,I2514);
DFFARX1 I_5498 (I370373,I2507,I95998,I96024,);
not I_5499 (I96032,I96024);
nand I_5500 (I96049,I370355,I370370);
and I_5501 (I96066,I96049,I370346);
DFFARX1 I_5502 (I96066,I2507,I95998,I96092,);
DFFARX1 I_5503 (I370349,I2507,I95998,I96109,);
and I_5504 (I96117,I96109,I370364);
nor I_5505 (I96134,I96092,I96117);
DFFARX1 I_5506 (I96134,I2507,I95998,I95966,);
nand I_5507 (I96165,I96109,I370364);
nand I_5508 (I96182,I96032,I96165);
not I_5509 (I95978,I96182);
DFFARX1 I_5510 (I370367,I2507,I95998,I96222,);
DFFARX1 I_5511 (I96222,I2507,I95998,I95987,);
nand I_5512 (I96244,I370346,I370358);
and I_5513 (I96261,I96244,I370352);
DFFARX1 I_5514 (I96261,I2507,I95998,I96287,);
DFFARX1 I_5515 (I96287,I2507,I95998,I96304,);
not I_5516 (I95990,I96304);
not I_5517 (I96326,I96287);
nand I_5518 (I95975,I96326,I96165);
nor I_5519 (I96357,I370361,I370358);
not I_5520 (I96374,I96357);
nor I_5521 (I96391,I96326,I96374);
nor I_5522 (I96408,I96032,I96391);
DFFARX1 I_5523 (I96408,I2507,I95998,I95984,);
nor I_5524 (I96439,I96092,I96374);
nor I_5525 (I95972,I96287,I96439);
nor I_5526 (I95981,I96222,I96357);
nor I_5527 (I95969,I96092,I96357);
not I_5528 (I96525,I2514);
DFFARX1 I_5529 (I1261133,I2507,I96525,I96551,);
not I_5530 (I96559,I96551);
nand I_5531 (I96576,I1261136,I1261130);
and I_5532 (I96593,I96576,I1261127);
DFFARX1 I_5533 (I96593,I2507,I96525,I96619,);
DFFARX1 I_5534 (I1261112,I2507,I96525,I96636,);
and I_5535 (I96644,I96636,I1261121);
nor I_5536 (I96661,I96619,I96644);
DFFARX1 I_5537 (I96661,I2507,I96525,I96493,);
nand I_5538 (I96692,I96636,I1261121);
nand I_5539 (I96709,I96559,I96692);
not I_5540 (I96505,I96709);
DFFARX1 I_5541 (I1261112,I2507,I96525,I96749,);
DFFARX1 I_5542 (I96749,I2507,I96525,I96514,);
nand I_5543 (I96771,I1261115,I1261118);
and I_5544 (I96788,I96771,I1261124);
DFFARX1 I_5545 (I96788,I2507,I96525,I96814,);
DFFARX1 I_5546 (I96814,I2507,I96525,I96831,);
not I_5547 (I96517,I96831);
not I_5548 (I96853,I96814);
nand I_5549 (I96502,I96853,I96692);
nor I_5550 (I96884,I1261115,I1261118);
not I_5551 (I96901,I96884);
nor I_5552 (I96918,I96853,I96901);
nor I_5553 (I96935,I96559,I96918);
DFFARX1 I_5554 (I96935,I2507,I96525,I96511,);
nor I_5555 (I96966,I96619,I96901);
nor I_5556 (I96499,I96814,I96966);
nor I_5557 (I96508,I96749,I96884);
nor I_5558 (I96496,I96619,I96884);
not I_5559 (I97052,I2514);
DFFARX1 I_5560 (I750376,I2507,I97052,I97078,);
not I_5561 (I97086,I97078);
nand I_5562 (I97103,I750367,I750385);
and I_5563 (I97120,I97103,I750364);
DFFARX1 I_5564 (I97120,I2507,I97052,I97146,);
DFFARX1 I_5565 (I750367,I2507,I97052,I97163,);
and I_5566 (I97171,I97163,I750370);
nor I_5567 (I97188,I97146,I97171);
DFFARX1 I_5568 (I97188,I2507,I97052,I97020,);
nand I_5569 (I97219,I97163,I750370);
nand I_5570 (I97236,I97086,I97219);
not I_5571 (I97032,I97236);
DFFARX1 I_5572 (I750364,I2507,I97052,I97276,);
DFFARX1 I_5573 (I97276,I2507,I97052,I97041,);
nand I_5574 (I97298,I750382,I750373);
and I_5575 (I97315,I97298,I750388);
DFFARX1 I_5576 (I97315,I2507,I97052,I97341,);
DFFARX1 I_5577 (I97341,I2507,I97052,I97358,);
not I_5578 (I97044,I97358);
not I_5579 (I97380,I97341);
nand I_5580 (I97029,I97380,I97219);
nor I_5581 (I97411,I750379,I750373);
not I_5582 (I97428,I97411);
nor I_5583 (I97445,I97380,I97428);
nor I_5584 (I97462,I97086,I97445);
DFFARX1 I_5585 (I97462,I2507,I97052,I97038,);
nor I_5586 (I97493,I97146,I97428);
nor I_5587 (I97026,I97341,I97493);
nor I_5588 (I97035,I97276,I97411);
nor I_5589 (I97023,I97146,I97411);
not I_5590 (I97579,I2514);
DFFARX1 I_5591 (I672346,I2507,I97579,I97605,);
not I_5592 (I97613,I97605);
nand I_5593 (I97630,I672337,I672355);
and I_5594 (I97647,I97630,I672334);
DFFARX1 I_5595 (I97647,I2507,I97579,I97673,);
DFFARX1 I_5596 (I672337,I2507,I97579,I97690,);
and I_5597 (I97698,I97690,I672340);
nor I_5598 (I97715,I97673,I97698);
DFFARX1 I_5599 (I97715,I2507,I97579,I97547,);
nand I_5600 (I97746,I97690,I672340);
nand I_5601 (I97763,I97613,I97746);
not I_5602 (I97559,I97763);
DFFARX1 I_5603 (I672334,I2507,I97579,I97803,);
DFFARX1 I_5604 (I97803,I2507,I97579,I97568,);
nand I_5605 (I97825,I672352,I672343);
and I_5606 (I97842,I97825,I672358);
DFFARX1 I_5607 (I97842,I2507,I97579,I97868,);
DFFARX1 I_5608 (I97868,I2507,I97579,I97885,);
not I_5609 (I97571,I97885);
not I_5610 (I97907,I97868);
nand I_5611 (I97556,I97907,I97746);
nor I_5612 (I97938,I672349,I672343);
not I_5613 (I97955,I97938);
nor I_5614 (I97972,I97907,I97955);
nor I_5615 (I97989,I97613,I97972);
DFFARX1 I_5616 (I97989,I2507,I97579,I97565,);
nor I_5617 (I98020,I97673,I97955);
nor I_5618 (I97553,I97868,I98020);
nor I_5619 (I97562,I97803,I97938);
nor I_5620 (I97550,I97673,I97938);
not I_5621 (I98106,I2514);
DFFARX1 I_5622 (I847052,I2507,I98106,I98132,);
not I_5623 (I98140,I98132);
nand I_5624 (I98157,I847049,I847064);
and I_5625 (I98174,I98157,I847046);
DFFARX1 I_5626 (I98174,I2507,I98106,I98200,);
DFFARX1 I_5627 (I847043,I2507,I98106,I98217,);
and I_5628 (I98225,I98217,I847043);
nor I_5629 (I98242,I98200,I98225);
DFFARX1 I_5630 (I98242,I2507,I98106,I98074,);
nand I_5631 (I98273,I98217,I847043);
nand I_5632 (I98290,I98140,I98273);
not I_5633 (I98086,I98290);
DFFARX1 I_5634 (I847046,I2507,I98106,I98330,);
DFFARX1 I_5635 (I98330,I2507,I98106,I98095,);
nand I_5636 (I98352,I847058,I847049);
and I_5637 (I98369,I98352,I847061);
DFFARX1 I_5638 (I98369,I2507,I98106,I98395,);
DFFARX1 I_5639 (I98395,I2507,I98106,I98412,);
not I_5640 (I98098,I98412);
not I_5641 (I98434,I98395);
nand I_5642 (I98083,I98434,I98273);
nor I_5643 (I98465,I847055,I847049);
not I_5644 (I98482,I98465);
nor I_5645 (I98499,I98434,I98482);
nor I_5646 (I98516,I98140,I98499);
DFFARX1 I_5647 (I98516,I2507,I98106,I98092,);
nor I_5648 (I98547,I98200,I98482);
nor I_5649 (I98080,I98395,I98547);
nor I_5650 (I98089,I98330,I98465);
nor I_5651 (I98077,I98200,I98465);
not I_5652 (I98633,I2514);
DFFARX1 I_5653 (I509562,I2507,I98633,I98659,);
not I_5654 (I98667,I98659);
nand I_5655 (I98684,I509583,I509577);
and I_5656 (I98701,I98684,I509559);
DFFARX1 I_5657 (I98701,I2507,I98633,I98727,);
DFFARX1 I_5658 (I509562,I2507,I98633,I98744,);
and I_5659 (I98752,I98744,I509571);
nor I_5660 (I98769,I98727,I98752);
DFFARX1 I_5661 (I98769,I2507,I98633,I98601,);
nand I_5662 (I98800,I98744,I509571);
nand I_5663 (I98817,I98667,I98800);
not I_5664 (I98613,I98817);
DFFARX1 I_5665 (I509568,I2507,I98633,I98857,);
DFFARX1 I_5666 (I98857,I2507,I98633,I98622,);
nand I_5667 (I98879,I509574,I509565);
and I_5668 (I98896,I98879,I509559);
DFFARX1 I_5669 (I98896,I2507,I98633,I98922,);
DFFARX1 I_5670 (I98922,I2507,I98633,I98939,);
not I_5671 (I98625,I98939);
not I_5672 (I98961,I98922);
nand I_5673 (I98610,I98961,I98800);
nor I_5674 (I98992,I509580,I509565);
not I_5675 (I99009,I98992);
nor I_5676 (I99026,I98961,I99009);
nor I_5677 (I99043,I98667,I99026);
DFFARX1 I_5678 (I99043,I2507,I98633,I98619,);
nor I_5679 (I99074,I98727,I99009);
nor I_5680 (I98607,I98922,I99074);
nor I_5681 (I98616,I98857,I98992);
nor I_5682 (I98604,I98727,I98992);
not I_5683 (I99160,I2514);
DFFARX1 I_5684 (I565413,I2507,I99160,I99186,);
not I_5685 (I99194,I99186);
nand I_5686 (I99211,I565425,I565410);
and I_5687 (I99228,I99211,I565404);
DFFARX1 I_5688 (I99228,I2507,I99160,I99254,);
DFFARX1 I_5689 (I565419,I2507,I99160,I99271,);
and I_5690 (I99279,I99271,I565407);
nor I_5691 (I99296,I99254,I99279);
DFFARX1 I_5692 (I99296,I2507,I99160,I99128,);
nand I_5693 (I99327,I99271,I565407);
nand I_5694 (I99344,I99194,I99327);
not I_5695 (I99140,I99344);
DFFARX1 I_5696 (I565416,I2507,I99160,I99384,);
DFFARX1 I_5697 (I99384,I2507,I99160,I99149,);
nand I_5698 (I99406,I565422,I565428);
and I_5699 (I99423,I99406,I565404);
DFFARX1 I_5700 (I99423,I2507,I99160,I99449,);
DFFARX1 I_5701 (I99449,I2507,I99160,I99466,);
not I_5702 (I99152,I99466);
not I_5703 (I99488,I99449);
nand I_5704 (I99137,I99488,I99327);
nor I_5705 (I99519,I565407,I565428);
not I_5706 (I99536,I99519);
nor I_5707 (I99553,I99488,I99536);
nor I_5708 (I99570,I99194,I99553);
DFFARX1 I_5709 (I99570,I2507,I99160,I99146,);
nor I_5710 (I99601,I99254,I99536);
nor I_5711 (I99134,I99449,I99601);
nor I_5712 (I99143,I99384,I99519);
nor I_5713 (I99131,I99254,I99519);
not I_5714 (I99687,I2514);
DFFARX1 I_5715 (I1636,I2507,I99687,I99713,);
not I_5716 (I99721,I99713);
nand I_5717 (I99738,I2124,I1700);
and I_5718 (I99755,I99738,I1476);
DFFARX1 I_5719 (I99755,I2507,I99687,I99781,);
DFFARX1 I_5720 (I2372,I2507,I99687,I99798,);
and I_5721 (I99806,I99798,I2348);
nor I_5722 (I99823,I99781,I99806);
DFFARX1 I_5723 (I99823,I2507,I99687,I99655,);
nand I_5724 (I99854,I99798,I2348);
nand I_5725 (I99871,I99721,I99854);
not I_5726 (I99667,I99871);
DFFARX1 I_5727 (I2452,I2507,I99687,I99911,);
DFFARX1 I_5728 (I99911,I2507,I99687,I99676,);
nand I_5729 (I99933,I2460,I2116);
and I_5730 (I99950,I99933,I2284);
DFFARX1 I_5731 (I99950,I2507,I99687,I99976,);
DFFARX1 I_5732 (I99976,I2507,I99687,I99993,);
not I_5733 (I99679,I99993);
not I_5734 (I100015,I99976);
nand I_5735 (I99664,I100015,I99854);
nor I_5736 (I100046,I1756,I2116);
not I_5737 (I100063,I100046);
nor I_5738 (I100080,I100015,I100063);
nor I_5739 (I100097,I99721,I100080);
DFFARX1 I_5740 (I100097,I2507,I99687,I99673,);
nor I_5741 (I100128,I99781,I100063);
nor I_5742 (I99661,I99976,I100128);
nor I_5743 (I99670,I99911,I100046);
nor I_5744 (I99658,I99781,I100046);
not I_5745 (I100214,I2514);
DFFARX1 I_5746 (I938614,I2507,I100214,I100240,);
not I_5747 (I100248,I100240);
nand I_5748 (I100265,I938632,I938626);
and I_5749 (I100282,I100265,I938605);
DFFARX1 I_5750 (I100282,I2507,I100214,I100308,);
DFFARX1 I_5751 (I938623,I2507,I100214,I100325,);
and I_5752 (I100333,I100325,I938608);
nor I_5753 (I100350,I100308,I100333);
DFFARX1 I_5754 (I100350,I2507,I100214,I100182,);
nand I_5755 (I100381,I100325,I938608);
nand I_5756 (I100398,I100248,I100381);
not I_5757 (I100194,I100398);
DFFARX1 I_5758 (I938620,I2507,I100214,I100438,);
DFFARX1 I_5759 (I100438,I2507,I100214,I100203,);
nand I_5760 (I100460,I938629,I938617);
and I_5761 (I100477,I100460,I938611);
DFFARX1 I_5762 (I100477,I2507,I100214,I100503,);
DFFARX1 I_5763 (I100503,I2507,I100214,I100520,);
not I_5764 (I100206,I100520);
not I_5765 (I100542,I100503);
nand I_5766 (I100191,I100542,I100381);
nor I_5767 (I100573,I938605,I938617);
not I_5768 (I100590,I100573);
nor I_5769 (I100607,I100542,I100590);
nor I_5770 (I100624,I100248,I100607);
DFFARX1 I_5771 (I100624,I2507,I100214,I100200,);
nor I_5772 (I100655,I100308,I100590);
nor I_5773 (I100188,I100503,I100655);
nor I_5774 (I100197,I100438,I100573);
nor I_5775 (I100185,I100308,I100573);
not I_5776 (I100741,I2514);
DFFARX1 I_5777 (I1167040,I2507,I100741,I100767,);
not I_5778 (I100775,I100767);
nand I_5779 (I100792,I1167055,I1167034);
and I_5780 (I100809,I100792,I1167037);
DFFARX1 I_5781 (I100809,I2507,I100741,I100835,);
DFFARX1 I_5782 (I1167058,I2507,I100741,I100852,);
and I_5783 (I100860,I100852,I1167037);
nor I_5784 (I100877,I100835,I100860);
DFFARX1 I_5785 (I100877,I2507,I100741,I100709,);
nand I_5786 (I100908,I100852,I1167037);
nand I_5787 (I100925,I100775,I100908);
not I_5788 (I100721,I100925);
DFFARX1 I_5789 (I1167034,I2507,I100741,I100965,);
DFFARX1 I_5790 (I100965,I2507,I100741,I100730,);
nand I_5791 (I100987,I1167046,I1167043);
and I_5792 (I101004,I100987,I1167049);
DFFARX1 I_5793 (I101004,I2507,I100741,I101030,);
DFFARX1 I_5794 (I101030,I2507,I100741,I101047,);
not I_5795 (I100733,I101047);
not I_5796 (I101069,I101030);
nand I_5797 (I100718,I101069,I100908);
nor I_5798 (I101100,I1167052,I1167043);
not I_5799 (I101117,I101100);
nor I_5800 (I101134,I101069,I101117);
nor I_5801 (I101151,I100775,I101134);
DFFARX1 I_5802 (I101151,I2507,I100741,I100727,);
nor I_5803 (I101182,I100835,I101117);
nor I_5804 (I100715,I101030,I101182);
nor I_5805 (I100724,I100965,I101100);
nor I_5806 (I100712,I100835,I101100);
not I_5807 (I101268,I2514);
DFFARX1 I_5808 (I1340429,I2507,I101268,I101294,);
not I_5809 (I101302,I101294);
nand I_5810 (I101319,I1340423,I1340444);
and I_5811 (I101336,I101319,I1340420);
DFFARX1 I_5812 (I101336,I2507,I101268,I101362,);
DFFARX1 I_5813 (I1340441,I2507,I101268,I101379,);
and I_5814 (I101387,I101379,I1340438);
nor I_5815 (I101404,I101362,I101387);
DFFARX1 I_5816 (I101404,I2507,I101268,I101236,);
nand I_5817 (I101435,I101379,I1340438);
nand I_5818 (I101452,I101302,I101435);
not I_5819 (I101248,I101452);
DFFARX1 I_5820 (I1340426,I2507,I101268,I101492,);
DFFARX1 I_5821 (I101492,I2507,I101268,I101257,);
nand I_5822 (I101514,I1340435,I1340432);
and I_5823 (I101531,I101514,I1340417);
DFFARX1 I_5824 (I101531,I2507,I101268,I101557,);
DFFARX1 I_5825 (I101557,I2507,I101268,I101574,);
not I_5826 (I101260,I101574);
not I_5827 (I101596,I101557);
nand I_5828 (I101245,I101596,I101435);
nor I_5829 (I101627,I1340417,I1340432);
not I_5830 (I101644,I101627);
nor I_5831 (I101661,I101596,I101644);
nor I_5832 (I101678,I101302,I101661);
DFFARX1 I_5833 (I101678,I2507,I101268,I101254,);
nor I_5834 (I101709,I101362,I101644);
nor I_5835 (I101242,I101557,I101709);
nor I_5836 (I101251,I101492,I101627);
nor I_5837 (I101239,I101362,I101627);
not I_5838 (I101795,I2514);
DFFARX1 I_5839 (I188322,I2507,I101795,I101821,);
not I_5840 (I101829,I101821);
nand I_5841 (I101846,I188316,I188310);
and I_5842 (I101863,I101846,I188331);
DFFARX1 I_5843 (I101863,I2507,I101795,I101889,);
DFFARX1 I_5844 (I188328,I2507,I101795,I101906,);
and I_5845 (I101914,I101906,I188325);
nor I_5846 (I101931,I101889,I101914);
DFFARX1 I_5847 (I101931,I2507,I101795,I101763,);
nand I_5848 (I101962,I101906,I188325);
nand I_5849 (I101979,I101829,I101962);
not I_5850 (I101775,I101979);
DFFARX1 I_5851 (I188310,I2507,I101795,I102019,);
DFFARX1 I_5852 (I102019,I2507,I101795,I101784,);
nand I_5853 (I102041,I188313,I188313);
and I_5854 (I102058,I102041,I188334);
DFFARX1 I_5855 (I102058,I2507,I101795,I102084,);
DFFARX1 I_5856 (I102084,I2507,I101795,I102101,);
not I_5857 (I101787,I102101);
not I_5858 (I102123,I102084);
nand I_5859 (I101772,I102123,I101962);
nor I_5860 (I102154,I188319,I188313);
not I_5861 (I102171,I102154);
nor I_5862 (I102188,I102123,I102171);
nor I_5863 (I102205,I101829,I102188);
DFFARX1 I_5864 (I102205,I2507,I101795,I101781,);
nor I_5865 (I102236,I101889,I102171);
nor I_5866 (I101769,I102084,I102236);
nor I_5867 (I101778,I102019,I102154);
nor I_5868 (I101766,I101889,I102154);
not I_5869 (I102322,I2514);
DFFARX1 I_5870 (I1336859,I2507,I102322,I102348,);
not I_5871 (I102356,I102348);
nand I_5872 (I102373,I1336853,I1336874);
and I_5873 (I102390,I102373,I1336850);
DFFARX1 I_5874 (I102390,I2507,I102322,I102416,);
DFFARX1 I_5875 (I1336871,I2507,I102322,I102433,);
and I_5876 (I102441,I102433,I1336868);
nor I_5877 (I102458,I102416,I102441);
DFFARX1 I_5878 (I102458,I2507,I102322,I102290,);
nand I_5879 (I102489,I102433,I1336868);
nand I_5880 (I102506,I102356,I102489);
not I_5881 (I102302,I102506);
DFFARX1 I_5882 (I1336856,I2507,I102322,I102546,);
DFFARX1 I_5883 (I102546,I2507,I102322,I102311,);
nand I_5884 (I102568,I1336865,I1336862);
and I_5885 (I102585,I102568,I1336847);
DFFARX1 I_5886 (I102585,I2507,I102322,I102611,);
DFFARX1 I_5887 (I102611,I2507,I102322,I102628,);
not I_5888 (I102314,I102628);
not I_5889 (I102650,I102611);
nand I_5890 (I102299,I102650,I102489);
nor I_5891 (I102681,I1336847,I1336862);
not I_5892 (I102698,I102681);
nor I_5893 (I102715,I102650,I102698);
nor I_5894 (I102732,I102356,I102715);
DFFARX1 I_5895 (I102732,I2507,I102322,I102308,);
nor I_5896 (I102763,I102416,I102698);
nor I_5897 (I102296,I102611,I102763);
nor I_5898 (I102305,I102546,I102681);
nor I_5899 (I102293,I102416,I102681);
not I_5900 (I102849,I2514);
DFFARX1 I_5901 (I235922,I2507,I102849,I102875,);
not I_5902 (I102883,I102875);
nand I_5903 (I102900,I235916,I235910);
and I_5904 (I102917,I102900,I235931);
DFFARX1 I_5905 (I102917,I2507,I102849,I102943,);
DFFARX1 I_5906 (I235928,I2507,I102849,I102960,);
and I_5907 (I102968,I102960,I235925);
nor I_5908 (I102985,I102943,I102968);
DFFARX1 I_5909 (I102985,I2507,I102849,I102817,);
nand I_5910 (I103016,I102960,I235925);
nand I_5911 (I103033,I102883,I103016);
not I_5912 (I102829,I103033);
DFFARX1 I_5913 (I235910,I2507,I102849,I103073,);
DFFARX1 I_5914 (I103073,I2507,I102849,I102838,);
nand I_5915 (I103095,I235913,I235913);
and I_5916 (I103112,I103095,I235934);
DFFARX1 I_5917 (I103112,I2507,I102849,I103138,);
DFFARX1 I_5918 (I103138,I2507,I102849,I103155,);
not I_5919 (I102841,I103155);
not I_5920 (I103177,I103138);
nand I_5921 (I102826,I103177,I103016);
nor I_5922 (I103208,I235919,I235913);
not I_5923 (I103225,I103208);
nor I_5924 (I103242,I103177,I103225);
nor I_5925 (I103259,I102883,I103242);
DFFARX1 I_5926 (I103259,I2507,I102849,I102835,);
nor I_5927 (I103290,I102943,I103225);
nor I_5928 (I102823,I103138,I103290);
nor I_5929 (I102832,I103073,I103208);
nor I_5930 (I102820,I102943,I103208);
not I_5931 (I103376,I2514);
DFFARX1 I_5932 (I923756,I2507,I103376,I103402,);
not I_5933 (I103410,I103402);
nand I_5934 (I103427,I923774,I923768);
and I_5935 (I103444,I103427,I923747);
DFFARX1 I_5936 (I103444,I2507,I103376,I103470,);
DFFARX1 I_5937 (I923765,I2507,I103376,I103487,);
and I_5938 (I103495,I103487,I923750);
nor I_5939 (I103512,I103470,I103495);
DFFARX1 I_5940 (I103512,I2507,I103376,I103344,);
nand I_5941 (I103543,I103487,I923750);
nand I_5942 (I103560,I103410,I103543);
not I_5943 (I103356,I103560);
DFFARX1 I_5944 (I923762,I2507,I103376,I103600,);
DFFARX1 I_5945 (I103600,I2507,I103376,I103365,);
nand I_5946 (I103622,I923771,I923759);
and I_5947 (I103639,I103622,I923753);
DFFARX1 I_5948 (I103639,I2507,I103376,I103665,);
DFFARX1 I_5949 (I103665,I2507,I103376,I103682,);
not I_5950 (I103368,I103682);
not I_5951 (I103704,I103665);
nand I_5952 (I103353,I103704,I103543);
nor I_5953 (I103735,I923747,I923759);
not I_5954 (I103752,I103735);
nor I_5955 (I103769,I103704,I103752);
nor I_5956 (I103786,I103410,I103769);
DFFARX1 I_5957 (I103786,I2507,I103376,I103362,);
nor I_5958 (I103817,I103470,I103752);
nor I_5959 (I103350,I103665,I103817);
nor I_5960 (I103359,I103600,I103735);
nor I_5961 (I103347,I103470,I103735);
not I_5962 (I103903,I2514);
DFFARX1 I_5963 (I1028096,I2507,I103903,I103929,);
not I_5964 (I103937,I103929);
nand I_5965 (I103954,I1028093,I1028099);
and I_5966 (I103971,I103954,I1028096);
DFFARX1 I_5967 (I103971,I2507,I103903,I103997,);
DFFARX1 I_5968 (I1028099,I2507,I103903,I104014,);
and I_5969 (I104022,I104014,I1028093);
nor I_5970 (I104039,I103997,I104022);
DFFARX1 I_5971 (I104039,I2507,I103903,I103871,);
nand I_5972 (I104070,I104014,I1028093);
nand I_5973 (I104087,I103937,I104070);
not I_5974 (I103883,I104087);
DFFARX1 I_5975 (I1028102,I2507,I103903,I104127,);
DFFARX1 I_5976 (I104127,I2507,I103903,I103892,);
nand I_5977 (I104149,I1028105,I1028114);
and I_5978 (I104166,I104149,I1028108);
DFFARX1 I_5979 (I104166,I2507,I103903,I104192,);
DFFARX1 I_5980 (I104192,I2507,I103903,I104209,);
not I_5981 (I103895,I104209);
not I_5982 (I104231,I104192);
nand I_5983 (I103880,I104231,I104070);
nor I_5984 (I104262,I1028111,I1028114);
not I_5985 (I104279,I104262);
nor I_5986 (I104296,I104231,I104279);
nor I_5987 (I104313,I103937,I104296);
DFFARX1 I_5988 (I104313,I2507,I103903,I103889,);
nor I_5989 (I104344,I103997,I104279);
nor I_5990 (I103877,I104192,I104344);
nor I_5991 (I103886,I104127,I104262);
nor I_5992 (I103874,I103997,I104262);
not I_5993 (I104430,I2514);
DFFARX1 I_5994 (I1356494,I2507,I104430,I104456,);
not I_5995 (I104464,I104456);
nand I_5996 (I104481,I1356488,I1356509);
and I_5997 (I104498,I104481,I1356485);
DFFARX1 I_5998 (I104498,I2507,I104430,I104524,);
DFFARX1 I_5999 (I1356506,I2507,I104430,I104541,);
and I_6000 (I104549,I104541,I1356503);
nor I_6001 (I104566,I104524,I104549);
DFFARX1 I_6002 (I104566,I2507,I104430,I104398,);
nand I_6003 (I104597,I104541,I1356503);
nand I_6004 (I104614,I104464,I104597);
not I_6005 (I104410,I104614);
DFFARX1 I_6006 (I1356491,I2507,I104430,I104654,);
DFFARX1 I_6007 (I104654,I2507,I104430,I104419,);
nand I_6008 (I104676,I1356500,I1356497);
and I_6009 (I104693,I104676,I1356482);
DFFARX1 I_6010 (I104693,I2507,I104430,I104719,);
DFFARX1 I_6011 (I104719,I2507,I104430,I104736,);
not I_6012 (I104422,I104736);
not I_6013 (I104758,I104719);
nand I_6014 (I104407,I104758,I104597);
nor I_6015 (I104789,I1356482,I1356497);
not I_6016 (I104806,I104789);
nor I_6017 (I104823,I104758,I104806);
nor I_6018 (I104840,I104464,I104823);
DFFARX1 I_6019 (I104840,I2507,I104430,I104416,);
nor I_6020 (I104871,I104524,I104806);
nor I_6021 (I104404,I104719,I104871);
nor I_6022 (I104413,I104654,I104789);
nor I_6023 (I104401,I104524,I104789);
not I_6024 (I104957,I2514);
DFFARX1 I_6025 (I911482,I2507,I104957,I104983,);
not I_6026 (I104991,I104983);
nand I_6027 (I105008,I911500,I911494);
and I_6028 (I105025,I105008,I911473);
DFFARX1 I_6029 (I105025,I2507,I104957,I105051,);
DFFARX1 I_6030 (I911491,I2507,I104957,I105068,);
and I_6031 (I105076,I105068,I911476);
nor I_6032 (I105093,I105051,I105076);
DFFARX1 I_6033 (I105093,I2507,I104957,I104925,);
nand I_6034 (I105124,I105068,I911476);
nand I_6035 (I105141,I104991,I105124);
not I_6036 (I104937,I105141);
DFFARX1 I_6037 (I911488,I2507,I104957,I105181,);
DFFARX1 I_6038 (I105181,I2507,I104957,I104946,);
nand I_6039 (I105203,I911497,I911485);
and I_6040 (I105220,I105203,I911479);
DFFARX1 I_6041 (I105220,I2507,I104957,I105246,);
DFFARX1 I_6042 (I105246,I2507,I104957,I105263,);
not I_6043 (I104949,I105263);
not I_6044 (I105285,I105246);
nand I_6045 (I104934,I105285,I105124);
nor I_6046 (I105316,I911473,I911485);
not I_6047 (I105333,I105316);
nor I_6048 (I105350,I105285,I105333);
nor I_6049 (I105367,I104991,I105350);
DFFARX1 I_6050 (I105367,I2507,I104957,I104943,);
nor I_6051 (I105398,I105051,I105333);
nor I_6052 (I104931,I105246,I105398);
nor I_6053 (I104940,I105181,I105316);
nor I_6054 (I104928,I105051,I105316);
not I_6055 (I105484,I2514);
DFFARX1 I_6056 (I1360659,I2507,I105484,I105510,);
not I_6057 (I105518,I105510);
nand I_6058 (I105535,I1360653,I1360674);
and I_6059 (I105552,I105535,I1360650);
DFFARX1 I_6060 (I105552,I2507,I105484,I105578,);
DFFARX1 I_6061 (I1360671,I2507,I105484,I105595,);
and I_6062 (I105603,I105595,I1360668);
nor I_6063 (I105620,I105578,I105603);
DFFARX1 I_6064 (I105620,I2507,I105484,I105452,);
nand I_6065 (I105651,I105595,I1360668);
nand I_6066 (I105668,I105518,I105651);
not I_6067 (I105464,I105668);
DFFARX1 I_6068 (I1360656,I2507,I105484,I105708,);
DFFARX1 I_6069 (I105708,I2507,I105484,I105473,);
nand I_6070 (I105730,I1360665,I1360662);
and I_6071 (I105747,I105730,I1360647);
DFFARX1 I_6072 (I105747,I2507,I105484,I105773,);
DFFARX1 I_6073 (I105773,I2507,I105484,I105790,);
not I_6074 (I105476,I105790);
not I_6075 (I105812,I105773);
nand I_6076 (I105461,I105812,I105651);
nor I_6077 (I105843,I1360647,I1360662);
not I_6078 (I105860,I105843);
nor I_6079 (I105877,I105812,I105860);
nor I_6080 (I105894,I105518,I105877);
DFFARX1 I_6081 (I105894,I2507,I105484,I105470,);
nor I_6082 (I105925,I105578,I105860);
nor I_6083 (I105458,I105773,I105925);
nor I_6084 (I105467,I105708,I105843);
nor I_6085 (I105455,I105578,I105843);
not I_6086 (I106011,I2514);
DFFARX1 I_6087 (I377249,I2507,I106011,I106037,);
not I_6088 (I106045,I106037);
nand I_6089 (I106062,I377243,I377234);
and I_6090 (I106079,I106062,I377255);
DFFARX1 I_6091 (I106079,I2507,I106011,I106105,);
DFFARX1 I_6092 (I377237,I2507,I106011,I106122,);
and I_6093 (I106130,I106122,I377231);
nor I_6094 (I106147,I106105,I106130);
DFFARX1 I_6095 (I106147,I2507,I106011,I105979,);
nand I_6096 (I106178,I106122,I377231);
nand I_6097 (I106195,I106045,I106178);
not I_6098 (I105991,I106195);
DFFARX1 I_6099 (I377231,I2507,I106011,I106235,);
DFFARX1 I_6100 (I106235,I2507,I106011,I106000,);
nand I_6101 (I106257,I377258,I377240);
and I_6102 (I106274,I106257,I377246);
DFFARX1 I_6103 (I106274,I2507,I106011,I106300,);
DFFARX1 I_6104 (I106300,I2507,I106011,I106317,);
not I_6105 (I106003,I106317);
not I_6106 (I106339,I106300);
nand I_6107 (I105988,I106339,I106178);
nor I_6108 (I106370,I377252,I377240);
not I_6109 (I106387,I106370);
nor I_6110 (I106404,I106339,I106387);
nor I_6111 (I106421,I106045,I106404);
DFFARX1 I_6112 (I106421,I2507,I106011,I105997,);
nor I_6113 (I106452,I106105,I106387);
nor I_6114 (I105985,I106300,I106452);
nor I_6115 (I105994,I106235,I106370);
nor I_6116 (I105982,I106105,I106370);
not I_6117 (I106538,I2514);
DFFARX1 I_6118 (I312930,I2507,I106538,I106564,);
not I_6119 (I106572,I106564);
nand I_6120 (I106589,I312912,I312927);
and I_6121 (I106606,I106589,I312903);
DFFARX1 I_6122 (I106606,I2507,I106538,I106632,);
DFFARX1 I_6123 (I312906,I2507,I106538,I106649,);
and I_6124 (I106657,I106649,I312921);
nor I_6125 (I106674,I106632,I106657);
DFFARX1 I_6126 (I106674,I2507,I106538,I106506,);
nand I_6127 (I106705,I106649,I312921);
nand I_6128 (I106722,I106572,I106705);
not I_6129 (I106518,I106722);
DFFARX1 I_6130 (I312924,I2507,I106538,I106762,);
DFFARX1 I_6131 (I106762,I2507,I106538,I106527,);
nand I_6132 (I106784,I312903,I312915);
and I_6133 (I106801,I106784,I312909);
DFFARX1 I_6134 (I106801,I2507,I106538,I106827,);
DFFARX1 I_6135 (I106827,I2507,I106538,I106844,);
not I_6136 (I106530,I106844);
not I_6137 (I106866,I106827);
nand I_6138 (I106515,I106866,I106705);
nor I_6139 (I106897,I312918,I312915);
not I_6140 (I106914,I106897);
nor I_6141 (I106931,I106866,I106914);
nor I_6142 (I106948,I106572,I106931);
DFFARX1 I_6143 (I106948,I2507,I106538,I106524,);
nor I_6144 (I106979,I106632,I106914);
nor I_6145 (I106512,I106827,I106979);
nor I_6146 (I106521,I106762,I106897);
nor I_6147 (I106509,I106632,I106897);
not I_6148 (I107065,I2514);
DFFARX1 I_6149 (I523247,I2507,I107065,I107091,);
not I_6150 (I107099,I107091);
nand I_6151 (I107116,I523268,I523262);
and I_6152 (I107133,I107116,I523244);
DFFARX1 I_6153 (I107133,I2507,I107065,I107159,);
DFFARX1 I_6154 (I523247,I2507,I107065,I107176,);
and I_6155 (I107184,I107176,I523256);
nor I_6156 (I107201,I107159,I107184);
DFFARX1 I_6157 (I107201,I2507,I107065,I107033,);
nand I_6158 (I107232,I107176,I523256);
nand I_6159 (I107249,I107099,I107232);
not I_6160 (I107045,I107249);
DFFARX1 I_6161 (I523253,I2507,I107065,I107289,);
DFFARX1 I_6162 (I107289,I2507,I107065,I107054,);
nand I_6163 (I107311,I523259,I523250);
and I_6164 (I107328,I107311,I523244);
DFFARX1 I_6165 (I107328,I2507,I107065,I107354,);
DFFARX1 I_6166 (I107354,I2507,I107065,I107371,);
not I_6167 (I107057,I107371);
not I_6168 (I107393,I107354);
nand I_6169 (I107042,I107393,I107232);
nor I_6170 (I107424,I523265,I523250);
not I_6171 (I107441,I107424);
nor I_6172 (I107458,I107393,I107441);
nor I_6173 (I107475,I107099,I107458);
DFFARX1 I_6174 (I107475,I2507,I107065,I107051,);
nor I_6175 (I107506,I107159,I107441);
nor I_6176 (I107039,I107354,I107506);
nor I_6177 (I107048,I107289,I107424);
nor I_6178 (I107036,I107159,I107424);
not I_6179 (I107592,I2514);
DFFARX1 I_6180 (I888872,I2507,I107592,I107618,);
not I_6181 (I107626,I107618);
nand I_6182 (I107643,I888890,I888884);
and I_6183 (I107660,I107643,I888863);
DFFARX1 I_6184 (I107660,I2507,I107592,I107686,);
DFFARX1 I_6185 (I888881,I2507,I107592,I107703,);
and I_6186 (I107711,I107703,I888866);
nor I_6187 (I107728,I107686,I107711);
DFFARX1 I_6188 (I107728,I2507,I107592,I107560,);
nand I_6189 (I107759,I107703,I888866);
nand I_6190 (I107776,I107626,I107759);
not I_6191 (I107572,I107776);
DFFARX1 I_6192 (I888878,I2507,I107592,I107816,);
DFFARX1 I_6193 (I107816,I2507,I107592,I107581,);
nand I_6194 (I107838,I888887,I888875);
and I_6195 (I107855,I107838,I888869);
DFFARX1 I_6196 (I107855,I2507,I107592,I107881,);
DFFARX1 I_6197 (I107881,I2507,I107592,I107898,);
not I_6198 (I107584,I107898);
not I_6199 (I107920,I107881);
nand I_6200 (I107569,I107920,I107759);
nor I_6201 (I107951,I888863,I888875);
not I_6202 (I107968,I107951);
nor I_6203 (I107985,I107920,I107968);
nor I_6204 (I108002,I107626,I107985);
DFFARX1 I_6205 (I108002,I2507,I107592,I107578,);
nor I_6206 (I108033,I107686,I107968);
nor I_6207 (I107566,I107881,I108033);
nor I_6208 (I107575,I107816,I107951);
nor I_6209 (I107563,I107686,I107951);
not I_6210 (I108119,I2514);
DFFARX1 I_6211 (I778542,I2507,I108119,I108145,);
not I_6212 (I108153,I108145);
nand I_6213 (I108170,I778539,I778554);
and I_6214 (I108187,I108170,I778536);
DFFARX1 I_6215 (I108187,I2507,I108119,I108213,);
DFFARX1 I_6216 (I778533,I2507,I108119,I108230,);
and I_6217 (I108238,I108230,I778533);
nor I_6218 (I108255,I108213,I108238);
DFFARX1 I_6219 (I108255,I2507,I108119,I108087,);
nand I_6220 (I108286,I108230,I778533);
nand I_6221 (I108303,I108153,I108286);
not I_6222 (I108099,I108303);
DFFARX1 I_6223 (I778536,I2507,I108119,I108343,);
DFFARX1 I_6224 (I108343,I2507,I108119,I108108,);
nand I_6225 (I108365,I778548,I778539);
and I_6226 (I108382,I108365,I778551);
DFFARX1 I_6227 (I108382,I2507,I108119,I108408,);
DFFARX1 I_6228 (I108408,I2507,I108119,I108425,);
not I_6229 (I108111,I108425);
not I_6230 (I108447,I108408);
nand I_6231 (I108096,I108447,I108286);
nor I_6232 (I108478,I778545,I778539);
not I_6233 (I108495,I108478);
nor I_6234 (I108512,I108447,I108495);
nor I_6235 (I108529,I108153,I108512);
DFFARX1 I_6236 (I108529,I2507,I108119,I108105,);
nor I_6237 (I108560,I108213,I108495);
nor I_6238 (I108093,I108408,I108560);
nor I_6239 (I108102,I108343,I108478);
nor I_6240 (I108090,I108213,I108478);
not I_6241 (I108646,I2514);
DFFARX1 I_6242 (I513132,I2507,I108646,I108672,);
not I_6243 (I108680,I108672);
nand I_6244 (I108697,I513153,I513147);
and I_6245 (I108714,I108697,I513129);
DFFARX1 I_6246 (I108714,I2507,I108646,I108740,);
DFFARX1 I_6247 (I513132,I2507,I108646,I108757,);
and I_6248 (I108765,I108757,I513141);
nor I_6249 (I108782,I108740,I108765);
DFFARX1 I_6250 (I108782,I2507,I108646,I108614,);
nand I_6251 (I108813,I108757,I513141);
nand I_6252 (I108830,I108680,I108813);
not I_6253 (I108626,I108830);
DFFARX1 I_6254 (I513138,I2507,I108646,I108870,);
DFFARX1 I_6255 (I108870,I2507,I108646,I108635,);
nand I_6256 (I108892,I513144,I513135);
and I_6257 (I108909,I108892,I513129);
DFFARX1 I_6258 (I108909,I2507,I108646,I108935,);
DFFARX1 I_6259 (I108935,I2507,I108646,I108952,);
not I_6260 (I108638,I108952);
not I_6261 (I108974,I108935);
nand I_6262 (I108623,I108974,I108813);
nor I_6263 (I109005,I513150,I513135);
not I_6264 (I109022,I109005);
nor I_6265 (I109039,I108974,I109022);
nor I_6266 (I109056,I108680,I109039);
DFFARX1 I_6267 (I109056,I2507,I108646,I108632,);
nor I_6268 (I109087,I108740,I109022);
nor I_6269 (I108620,I108935,I109087);
nor I_6270 (I108629,I108870,I109005);
nor I_6271 (I108617,I108740,I109005);
not I_6272 (I109173,I2514);
DFFARX1 I_6273 (I839674,I2507,I109173,I109199,);
not I_6274 (I109207,I109199);
nand I_6275 (I109224,I839671,I839686);
and I_6276 (I109241,I109224,I839668);
DFFARX1 I_6277 (I109241,I2507,I109173,I109267,);
DFFARX1 I_6278 (I839665,I2507,I109173,I109284,);
and I_6279 (I109292,I109284,I839665);
nor I_6280 (I109309,I109267,I109292);
DFFARX1 I_6281 (I109309,I2507,I109173,I109141,);
nand I_6282 (I109340,I109284,I839665);
nand I_6283 (I109357,I109207,I109340);
not I_6284 (I109153,I109357);
DFFARX1 I_6285 (I839668,I2507,I109173,I109397,);
DFFARX1 I_6286 (I109397,I2507,I109173,I109162,);
nand I_6287 (I109419,I839680,I839671);
and I_6288 (I109436,I109419,I839683);
DFFARX1 I_6289 (I109436,I2507,I109173,I109462,);
DFFARX1 I_6290 (I109462,I2507,I109173,I109479,);
not I_6291 (I109165,I109479);
not I_6292 (I109501,I109462);
nand I_6293 (I109150,I109501,I109340);
nor I_6294 (I109532,I839677,I839671);
not I_6295 (I109549,I109532);
nor I_6296 (I109566,I109501,I109549);
nor I_6297 (I109583,I109207,I109566);
DFFARX1 I_6298 (I109583,I2507,I109173,I109159,);
nor I_6299 (I109614,I109267,I109549);
nor I_6300 (I109147,I109462,I109614);
nor I_6301 (I109156,I109397,I109532);
nor I_6302 (I109144,I109267,I109532);
not I_6303 (I109700,I2514);
DFFARX1 I_6304 (I822283,I2507,I109700,I109726,);
not I_6305 (I109734,I109726);
nand I_6306 (I109751,I822280,I822295);
and I_6307 (I109768,I109751,I822277);
DFFARX1 I_6308 (I109768,I2507,I109700,I109794,);
DFFARX1 I_6309 (I822274,I2507,I109700,I109811,);
and I_6310 (I109819,I109811,I822274);
nor I_6311 (I109836,I109794,I109819);
DFFARX1 I_6312 (I109836,I2507,I109700,I109668,);
nand I_6313 (I109867,I109811,I822274);
nand I_6314 (I109884,I109734,I109867);
not I_6315 (I109680,I109884);
DFFARX1 I_6316 (I822277,I2507,I109700,I109924,);
DFFARX1 I_6317 (I109924,I2507,I109700,I109689,);
nand I_6318 (I109946,I822289,I822280);
and I_6319 (I109963,I109946,I822292);
DFFARX1 I_6320 (I109963,I2507,I109700,I109989,);
DFFARX1 I_6321 (I109989,I2507,I109700,I110006,);
not I_6322 (I109692,I110006);
not I_6323 (I110028,I109989);
nand I_6324 (I109677,I110028,I109867);
nor I_6325 (I110059,I822286,I822280);
not I_6326 (I110076,I110059);
nor I_6327 (I110093,I110028,I110076);
nor I_6328 (I110110,I109734,I110093);
DFFARX1 I_6329 (I110110,I2507,I109700,I109686,);
nor I_6330 (I110141,I109794,I110076);
nor I_6331 (I109674,I109989,I110141);
nor I_6332 (I109683,I109924,I110059);
nor I_6333 (I109671,I109794,I110059);
not I_6334 (I110227,I2514);
DFFARX1 I_6335 (I391393,I2507,I110227,I110253,);
not I_6336 (I110261,I110253);
nand I_6337 (I110278,I391387,I391378);
and I_6338 (I110295,I110278,I391399);
DFFARX1 I_6339 (I110295,I2507,I110227,I110321,);
DFFARX1 I_6340 (I391381,I2507,I110227,I110338,);
and I_6341 (I110346,I110338,I391375);
nor I_6342 (I110363,I110321,I110346);
DFFARX1 I_6343 (I110363,I2507,I110227,I110195,);
nand I_6344 (I110394,I110338,I391375);
nand I_6345 (I110411,I110261,I110394);
not I_6346 (I110207,I110411);
DFFARX1 I_6347 (I391375,I2507,I110227,I110451,);
DFFARX1 I_6348 (I110451,I2507,I110227,I110216,);
nand I_6349 (I110473,I391402,I391384);
and I_6350 (I110490,I110473,I391390);
DFFARX1 I_6351 (I110490,I2507,I110227,I110516,);
DFFARX1 I_6352 (I110516,I2507,I110227,I110533,);
not I_6353 (I110219,I110533);
not I_6354 (I110555,I110516);
nand I_6355 (I110204,I110555,I110394);
nor I_6356 (I110586,I391396,I391384);
not I_6357 (I110603,I110586);
nor I_6358 (I110620,I110555,I110603);
nor I_6359 (I110637,I110261,I110620);
DFFARX1 I_6360 (I110637,I2507,I110227,I110213,);
nor I_6361 (I110668,I110321,I110603);
nor I_6362 (I110201,I110516,I110668);
nor I_6363 (I110210,I110451,I110586);
nor I_6364 (I110198,I110321,I110586);
not I_6365 (I110754,I2514);
DFFARX1 I_6366 (I809108,I2507,I110754,I110780,);
not I_6367 (I110788,I110780);
nand I_6368 (I110805,I809105,I809120);
and I_6369 (I110822,I110805,I809102);
DFFARX1 I_6370 (I110822,I2507,I110754,I110848,);
DFFARX1 I_6371 (I809099,I2507,I110754,I110865,);
and I_6372 (I110873,I110865,I809099);
nor I_6373 (I110890,I110848,I110873);
DFFARX1 I_6374 (I110890,I2507,I110754,I110722,);
nand I_6375 (I110921,I110865,I809099);
nand I_6376 (I110938,I110788,I110921);
not I_6377 (I110734,I110938);
DFFARX1 I_6378 (I809102,I2507,I110754,I110978,);
DFFARX1 I_6379 (I110978,I2507,I110754,I110743,);
nand I_6380 (I111000,I809114,I809105);
and I_6381 (I111017,I111000,I809117);
DFFARX1 I_6382 (I111017,I2507,I110754,I111043,);
DFFARX1 I_6383 (I111043,I2507,I110754,I111060,);
not I_6384 (I110746,I111060);
not I_6385 (I111082,I111043);
nand I_6386 (I110731,I111082,I110921);
nor I_6387 (I111113,I809111,I809105);
not I_6388 (I111130,I111113);
nor I_6389 (I111147,I111082,I111130);
nor I_6390 (I111164,I110788,I111147);
DFFARX1 I_6391 (I111164,I2507,I110754,I110740,);
nor I_6392 (I111195,I110848,I111130);
nor I_6393 (I110728,I111043,I111195);
nor I_6394 (I110737,I110978,I111113);
nor I_6395 (I110725,I110848,I111113);
not I_6396 (I111281,I2514);
DFFARX1 I_6397 (I814905,I2507,I111281,I111307,);
not I_6398 (I111315,I111307);
nand I_6399 (I111332,I814902,I814917);
and I_6400 (I111349,I111332,I814899);
DFFARX1 I_6401 (I111349,I2507,I111281,I111375,);
DFFARX1 I_6402 (I814896,I2507,I111281,I111392,);
and I_6403 (I111400,I111392,I814896);
nor I_6404 (I111417,I111375,I111400);
DFFARX1 I_6405 (I111417,I2507,I111281,I111249,);
nand I_6406 (I111448,I111392,I814896);
nand I_6407 (I111465,I111315,I111448);
not I_6408 (I111261,I111465);
DFFARX1 I_6409 (I814899,I2507,I111281,I111505,);
DFFARX1 I_6410 (I111505,I2507,I111281,I111270,);
nand I_6411 (I111527,I814911,I814902);
and I_6412 (I111544,I111527,I814914);
DFFARX1 I_6413 (I111544,I2507,I111281,I111570,);
DFFARX1 I_6414 (I111570,I2507,I111281,I111587,);
not I_6415 (I111273,I111587);
not I_6416 (I111609,I111570);
nand I_6417 (I111258,I111609,I111448);
nor I_6418 (I111640,I814908,I814902);
not I_6419 (I111657,I111640);
nor I_6420 (I111674,I111609,I111657);
nor I_6421 (I111691,I111315,I111674);
DFFARX1 I_6422 (I111691,I2507,I111281,I111267,);
nor I_6423 (I111722,I111375,I111657);
nor I_6424 (I111255,I111570,I111722);
nor I_6425 (I111264,I111505,I111640);
nor I_6426 (I111252,I111375,I111640);
not I_6427 (I111808,I2514);
DFFARX1 I_6428 (I1386244,I2507,I111808,I111834,);
not I_6429 (I111842,I111834);
nand I_6430 (I111859,I1386238,I1386259);
and I_6431 (I111876,I111859,I1386235);
DFFARX1 I_6432 (I111876,I2507,I111808,I111902,);
DFFARX1 I_6433 (I1386256,I2507,I111808,I111919,);
and I_6434 (I111927,I111919,I1386253);
nor I_6435 (I111944,I111902,I111927);
DFFARX1 I_6436 (I111944,I2507,I111808,I111776,);
nand I_6437 (I111975,I111919,I1386253);
nand I_6438 (I111992,I111842,I111975);
not I_6439 (I111788,I111992);
DFFARX1 I_6440 (I1386241,I2507,I111808,I112032,);
DFFARX1 I_6441 (I112032,I2507,I111808,I111797,);
nand I_6442 (I112054,I1386250,I1386247);
and I_6443 (I112071,I112054,I1386232);
DFFARX1 I_6444 (I112071,I2507,I111808,I112097,);
DFFARX1 I_6445 (I112097,I2507,I111808,I112114,);
not I_6446 (I111800,I112114);
not I_6447 (I112136,I112097);
nand I_6448 (I111785,I112136,I111975);
nor I_6449 (I112167,I1386232,I1386247);
not I_6450 (I112184,I112167);
nor I_6451 (I112201,I112136,I112184);
nor I_6452 (I112218,I111842,I112201);
DFFARX1 I_6453 (I112218,I2507,I111808,I111794,);
nor I_6454 (I112249,I111902,I112184);
nor I_6455 (I111782,I112097,I112249);
nor I_6456 (I111791,I112032,I112167);
nor I_6457 (I111779,I111902,I112167);
not I_6458 (I112335,I2514);
DFFARX1 I_6459 (I410977,I2507,I112335,I112361,);
not I_6460 (I112369,I112361);
nand I_6461 (I112386,I410971,I410962);
and I_6462 (I112403,I112386,I410983);
DFFARX1 I_6463 (I112403,I2507,I112335,I112429,);
DFFARX1 I_6464 (I410965,I2507,I112335,I112446,);
and I_6465 (I112454,I112446,I410959);
nor I_6466 (I112471,I112429,I112454);
DFFARX1 I_6467 (I112471,I2507,I112335,I112303,);
nand I_6468 (I112502,I112446,I410959);
nand I_6469 (I112519,I112369,I112502);
not I_6470 (I112315,I112519);
DFFARX1 I_6471 (I410959,I2507,I112335,I112559,);
DFFARX1 I_6472 (I112559,I2507,I112335,I112324,);
nand I_6473 (I112581,I410986,I410968);
and I_6474 (I112598,I112581,I410974);
DFFARX1 I_6475 (I112598,I2507,I112335,I112624,);
DFFARX1 I_6476 (I112624,I2507,I112335,I112641,);
not I_6477 (I112327,I112641);
not I_6478 (I112663,I112624);
nand I_6479 (I112312,I112663,I112502);
nor I_6480 (I112694,I410980,I410968);
not I_6481 (I112711,I112694);
nor I_6482 (I112728,I112663,I112711);
nor I_6483 (I112745,I112369,I112728);
DFFARX1 I_6484 (I112745,I2507,I112335,I112321,);
nor I_6485 (I112776,I112429,I112711);
nor I_6486 (I112309,I112624,I112776);
nor I_6487 (I112318,I112559,I112694);
nor I_6488 (I112306,I112429,I112694);
not I_6489 (I112862,I2514);
DFFARX1 I_6490 (I1329719,I2507,I112862,I112888,);
not I_6491 (I112896,I112888);
nand I_6492 (I112913,I1329713,I1329734);
and I_6493 (I112930,I112913,I1329710);
DFFARX1 I_6494 (I112930,I2507,I112862,I112956,);
DFFARX1 I_6495 (I1329731,I2507,I112862,I112973,);
and I_6496 (I112981,I112973,I1329728);
nor I_6497 (I112998,I112956,I112981);
DFFARX1 I_6498 (I112998,I2507,I112862,I112830,);
nand I_6499 (I113029,I112973,I1329728);
nand I_6500 (I113046,I112896,I113029);
not I_6501 (I112842,I113046);
DFFARX1 I_6502 (I1329716,I2507,I112862,I113086,);
DFFARX1 I_6503 (I113086,I2507,I112862,I112851,);
nand I_6504 (I113108,I1329725,I1329722);
and I_6505 (I113125,I113108,I1329707);
DFFARX1 I_6506 (I113125,I2507,I112862,I113151,);
DFFARX1 I_6507 (I113151,I2507,I112862,I113168,);
not I_6508 (I112854,I113168);
not I_6509 (I113190,I113151);
nand I_6510 (I112839,I113190,I113029);
nor I_6511 (I113221,I1329707,I1329722);
not I_6512 (I113238,I113221);
nor I_6513 (I113255,I113190,I113238);
nor I_6514 (I113272,I112896,I113255);
DFFARX1 I_6515 (I113272,I2507,I112862,I112848,);
nor I_6516 (I113303,I112956,I113238);
nor I_6517 (I112836,I113151,I113303);
nor I_6518 (I112845,I113086,I113221);
nor I_6519 (I112833,I112956,I113221);
not I_6520 (I113389,I2514);
DFFARX1 I_6521 (I18521,I2507,I113389,I113415,);
not I_6522 (I113423,I113415);
nand I_6523 (I113440,I18509,I18515);
and I_6524 (I113457,I113440,I18518);
DFFARX1 I_6525 (I113457,I2507,I113389,I113483,);
DFFARX1 I_6526 (I18500,I2507,I113389,I113500,);
and I_6527 (I113508,I113500,I18506);
nor I_6528 (I113525,I113483,I113508);
DFFARX1 I_6529 (I113525,I2507,I113389,I113357,);
nand I_6530 (I113556,I113500,I18506);
nand I_6531 (I113573,I113423,I113556);
not I_6532 (I113369,I113573);
DFFARX1 I_6533 (I18500,I2507,I113389,I113613,);
DFFARX1 I_6534 (I113613,I2507,I113389,I113378,);
nand I_6535 (I113635,I18503,I18497);
and I_6536 (I113652,I113635,I18512);
DFFARX1 I_6537 (I113652,I2507,I113389,I113678,);
DFFARX1 I_6538 (I113678,I2507,I113389,I113695,);
not I_6539 (I113381,I113695);
not I_6540 (I113717,I113678);
nand I_6541 (I113366,I113717,I113556);
nor I_6542 (I113748,I18497,I18497);
not I_6543 (I113765,I113748);
nor I_6544 (I113782,I113717,I113765);
nor I_6545 (I113799,I113423,I113782);
DFFARX1 I_6546 (I113799,I2507,I113389,I113375,);
nor I_6547 (I113830,I113483,I113765);
nor I_6548 (I113363,I113678,I113830);
nor I_6549 (I113372,I113613,I113748);
nor I_6550 (I113360,I113483,I113748);
not I_6551 (I113916,I2514);
DFFARX1 I_6552 (I705292,I2507,I113916,I113942,);
not I_6553 (I113950,I113942);
nand I_6554 (I113967,I705283,I705301);
and I_6555 (I113984,I113967,I705280);
DFFARX1 I_6556 (I113984,I2507,I113916,I114010,);
DFFARX1 I_6557 (I705283,I2507,I113916,I114027,);
and I_6558 (I114035,I114027,I705286);
nor I_6559 (I114052,I114010,I114035);
DFFARX1 I_6560 (I114052,I2507,I113916,I113884,);
nand I_6561 (I114083,I114027,I705286);
nand I_6562 (I114100,I113950,I114083);
not I_6563 (I113896,I114100);
DFFARX1 I_6564 (I705280,I2507,I113916,I114140,);
DFFARX1 I_6565 (I114140,I2507,I113916,I113905,);
nand I_6566 (I114162,I705298,I705289);
and I_6567 (I114179,I114162,I705304);
DFFARX1 I_6568 (I114179,I2507,I113916,I114205,);
DFFARX1 I_6569 (I114205,I2507,I113916,I114222,);
not I_6570 (I113908,I114222);
not I_6571 (I114244,I114205);
nand I_6572 (I113893,I114244,I114083);
nor I_6573 (I114275,I705295,I705289);
not I_6574 (I114292,I114275);
nor I_6575 (I114309,I114244,I114292);
nor I_6576 (I114326,I113950,I114309);
DFFARX1 I_6577 (I114326,I2507,I113916,I113902,);
nor I_6578 (I114357,I114010,I114292);
nor I_6579 (I113890,I114205,I114357);
nor I_6580 (I113899,I114140,I114275);
nor I_6581 (I113887,I114010,I114275);
not I_6582 (I114443,I2514);
DFFARX1 I_6583 (I1241704,I2507,I114443,I114469,);
not I_6584 (I114477,I114469);
nand I_6585 (I114494,I1241698,I1241719);
and I_6586 (I114511,I114494,I1241710);
DFFARX1 I_6587 (I114511,I2507,I114443,I114537,);
DFFARX1 I_6588 (I1241701,I2507,I114443,I114554,);
and I_6589 (I114562,I114554,I1241713);
nor I_6590 (I114579,I114537,I114562);
DFFARX1 I_6591 (I114579,I2507,I114443,I114411,);
nand I_6592 (I114610,I114554,I1241713);
nand I_6593 (I114627,I114477,I114610);
not I_6594 (I114423,I114627);
DFFARX1 I_6595 (I1241701,I2507,I114443,I114667,);
DFFARX1 I_6596 (I114667,I2507,I114443,I114432,);
nand I_6597 (I114689,I1241722,I1241707);
and I_6598 (I114706,I114689,I1241698);
DFFARX1 I_6599 (I114706,I2507,I114443,I114732,);
DFFARX1 I_6600 (I114732,I2507,I114443,I114749,);
not I_6601 (I114435,I114749);
not I_6602 (I114771,I114732);
nand I_6603 (I114420,I114771,I114610);
nor I_6604 (I114802,I1241716,I1241707);
not I_6605 (I114819,I114802);
nor I_6606 (I114836,I114771,I114819);
nor I_6607 (I114853,I114477,I114836);
DFFARX1 I_6608 (I114853,I2507,I114443,I114429,);
nor I_6609 (I114884,I114537,I114819);
nor I_6610 (I114417,I114732,I114884);
nor I_6611 (I114426,I114667,I114802);
nor I_6612 (I114414,I114537,I114802);
not I_6613 (I114970,I2514);
DFFARX1 I_6614 (I326105,I2507,I114970,I114996,);
not I_6615 (I115004,I114996);
nand I_6616 (I115021,I326087,I326102);
and I_6617 (I115038,I115021,I326078);
DFFARX1 I_6618 (I115038,I2507,I114970,I115064,);
DFFARX1 I_6619 (I326081,I2507,I114970,I115081,);
and I_6620 (I115089,I115081,I326096);
nor I_6621 (I115106,I115064,I115089);
DFFARX1 I_6622 (I115106,I2507,I114970,I114938,);
nand I_6623 (I115137,I115081,I326096);
nand I_6624 (I115154,I115004,I115137);
not I_6625 (I114950,I115154);
DFFARX1 I_6626 (I326099,I2507,I114970,I115194,);
DFFARX1 I_6627 (I115194,I2507,I114970,I114959,);
nand I_6628 (I115216,I326078,I326090);
and I_6629 (I115233,I115216,I326084);
DFFARX1 I_6630 (I115233,I2507,I114970,I115259,);
DFFARX1 I_6631 (I115259,I2507,I114970,I115276,);
not I_6632 (I114962,I115276);
not I_6633 (I115298,I115259);
nand I_6634 (I114947,I115298,I115137);
nor I_6635 (I115329,I326093,I326090);
not I_6636 (I115346,I115329);
nor I_6637 (I115363,I115298,I115346);
nor I_6638 (I115380,I115004,I115363);
DFFARX1 I_6639 (I115380,I2507,I114970,I114956,);
nor I_6640 (I115411,I115064,I115346);
nor I_6641 (I114944,I115259,I115411);
nor I_6642 (I114953,I115194,I115329);
nor I_6643 (I114941,I115064,I115329);
not I_6644 (I115497,I2514);
DFFARX1 I_6645 (I376705,I2507,I115497,I115523,);
not I_6646 (I115531,I115523);
nand I_6647 (I115548,I376699,I376690);
and I_6648 (I115565,I115548,I376711);
DFFARX1 I_6649 (I115565,I2507,I115497,I115591,);
DFFARX1 I_6650 (I376693,I2507,I115497,I115608,);
and I_6651 (I115616,I115608,I376687);
nor I_6652 (I115633,I115591,I115616);
DFFARX1 I_6653 (I115633,I2507,I115497,I115465,);
nand I_6654 (I115664,I115608,I376687);
nand I_6655 (I115681,I115531,I115664);
not I_6656 (I115477,I115681);
DFFARX1 I_6657 (I376687,I2507,I115497,I115721,);
DFFARX1 I_6658 (I115721,I2507,I115497,I115486,);
nand I_6659 (I115743,I376714,I376696);
and I_6660 (I115760,I115743,I376702);
DFFARX1 I_6661 (I115760,I2507,I115497,I115786,);
DFFARX1 I_6662 (I115786,I2507,I115497,I115803,);
not I_6663 (I115489,I115803);
not I_6664 (I115825,I115786);
nand I_6665 (I115474,I115825,I115664);
nor I_6666 (I115856,I376708,I376696);
not I_6667 (I115873,I115856);
nor I_6668 (I115890,I115825,I115873);
nor I_6669 (I115907,I115531,I115890);
DFFARX1 I_6670 (I115907,I2507,I115497,I115483,);
nor I_6671 (I115938,I115591,I115873);
nor I_6672 (I115471,I115786,I115938);
nor I_6673 (I115480,I115721,I115856);
nor I_6674 (I115468,I115591,I115856);
not I_6675 (I116024,I2514);
DFFARX1 I_6676 (I157977,I2507,I116024,I116050,);
not I_6677 (I116058,I116050);
nand I_6678 (I116075,I157971,I157965);
and I_6679 (I116092,I116075,I157986);
DFFARX1 I_6680 (I116092,I2507,I116024,I116118,);
DFFARX1 I_6681 (I157983,I2507,I116024,I116135,);
and I_6682 (I116143,I116135,I157980);
nor I_6683 (I116160,I116118,I116143);
DFFARX1 I_6684 (I116160,I2507,I116024,I115992,);
nand I_6685 (I116191,I116135,I157980);
nand I_6686 (I116208,I116058,I116191);
not I_6687 (I116004,I116208);
DFFARX1 I_6688 (I157965,I2507,I116024,I116248,);
DFFARX1 I_6689 (I116248,I2507,I116024,I116013,);
nand I_6690 (I116270,I157968,I157968);
and I_6691 (I116287,I116270,I157989);
DFFARX1 I_6692 (I116287,I2507,I116024,I116313,);
DFFARX1 I_6693 (I116313,I2507,I116024,I116330,);
not I_6694 (I116016,I116330);
not I_6695 (I116352,I116313);
nand I_6696 (I116001,I116352,I116191);
nor I_6697 (I116383,I157974,I157968);
not I_6698 (I116400,I116383);
nor I_6699 (I116417,I116352,I116400);
nor I_6700 (I116434,I116058,I116417);
DFFARX1 I_6701 (I116434,I2507,I116024,I116010,);
nor I_6702 (I116465,I116118,I116400);
nor I_6703 (I115998,I116313,I116465);
nor I_6704 (I116007,I116248,I116383);
nor I_6705 (I115995,I116118,I116383);
not I_6706 (I116551,I2514);
DFFARX1 I_6707 (I798568,I2507,I116551,I116577,);
not I_6708 (I116585,I116577);
nand I_6709 (I116602,I798565,I798580);
and I_6710 (I116619,I116602,I798562);
DFFARX1 I_6711 (I116619,I2507,I116551,I116645,);
DFFARX1 I_6712 (I798559,I2507,I116551,I116662,);
and I_6713 (I116670,I116662,I798559);
nor I_6714 (I116687,I116645,I116670);
DFFARX1 I_6715 (I116687,I2507,I116551,I116519,);
nand I_6716 (I116718,I116662,I798559);
nand I_6717 (I116735,I116585,I116718);
not I_6718 (I116531,I116735);
DFFARX1 I_6719 (I798562,I2507,I116551,I116775,);
DFFARX1 I_6720 (I116775,I2507,I116551,I116540,);
nand I_6721 (I116797,I798574,I798565);
and I_6722 (I116814,I116797,I798577);
DFFARX1 I_6723 (I116814,I2507,I116551,I116840,);
DFFARX1 I_6724 (I116840,I2507,I116551,I116857,);
not I_6725 (I116543,I116857);
not I_6726 (I116879,I116840);
nand I_6727 (I116528,I116879,I116718);
nor I_6728 (I116910,I798571,I798565);
not I_6729 (I116927,I116910);
nor I_6730 (I116944,I116879,I116927);
nor I_6731 (I116961,I116585,I116944);
DFFARX1 I_6732 (I116961,I2507,I116551,I116537,);
nor I_6733 (I116992,I116645,I116927);
nor I_6734 (I116525,I116840,I116992);
nor I_6735 (I116534,I116775,I116910);
nor I_6736 (I116522,I116645,I116910);
not I_6737 (I117078,I2514);
DFFARX1 I_6738 (I494209,I2507,I117078,I117104,);
not I_6739 (I117112,I117104);
nand I_6740 (I117129,I494203,I494194);
and I_6741 (I117146,I117129,I494215);
DFFARX1 I_6742 (I117146,I2507,I117078,I117172,);
DFFARX1 I_6743 (I494197,I2507,I117078,I117189,);
and I_6744 (I117197,I117189,I494191);
nor I_6745 (I117214,I117172,I117197);
DFFARX1 I_6746 (I117214,I2507,I117078,I117046,);
nand I_6747 (I117245,I117189,I494191);
nand I_6748 (I117262,I117112,I117245);
not I_6749 (I117058,I117262);
DFFARX1 I_6750 (I494191,I2507,I117078,I117302,);
DFFARX1 I_6751 (I117302,I2507,I117078,I117067,);
nand I_6752 (I117324,I494218,I494200);
and I_6753 (I117341,I117324,I494206);
DFFARX1 I_6754 (I117341,I2507,I117078,I117367,);
DFFARX1 I_6755 (I117367,I2507,I117078,I117384,);
not I_6756 (I117070,I117384);
not I_6757 (I117406,I117367);
nand I_6758 (I117055,I117406,I117245);
nor I_6759 (I117437,I494212,I494200);
not I_6760 (I117454,I117437);
nor I_6761 (I117471,I117406,I117454);
nor I_6762 (I117488,I117112,I117471);
DFFARX1 I_6763 (I117488,I2507,I117078,I117064,);
nor I_6764 (I117519,I117172,I117454);
nor I_6765 (I117052,I117367,I117519);
nor I_6766 (I117061,I117302,I117437);
nor I_6767 (I117049,I117172,I117437);
not I_6768 (I117605,I2514);
DFFARX1 I_6769 (I894040,I2507,I117605,I117631,);
not I_6770 (I117639,I117631);
nand I_6771 (I117656,I894058,I894052);
and I_6772 (I117673,I117656,I894031);
DFFARX1 I_6773 (I117673,I2507,I117605,I117699,);
DFFARX1 I_6774 (I894049,I2507,I117605,I117716,);
and I_6775 (I117724,I117716,I894034);
nor I_6776 (I117741,I117699,I117724);
DFFARX1 I_6777 (I117741,I2507,I117605,I117573,);
nand I_6778 (I117772,I117716,I894034);
nand I_6779 (I117789,I117639,I117772);
not I_6780 (I117585,I117789);
DFFARX1 I_6781 (I894046,I2507,I117605,I117829,);
DFFARX1 I_6782 (I117829,I2507,I117605,I117594,);
nand I_6783 (I117851,I894055,I894043);
and I_6784 (I117868,I117851,I894037);
DFFARX1 I_6785 (I117868,I2507,I117605,I117894,);
DFFARX1 I_6786 (I117894,I2507,I117605,I117911,);
not I_6787 (I117597,I117911);
not I_6788 (I117933,I117894);
nand I_6789 (I117582,I117933,I117772);
nor I_6790 (I117964,I894031,I894043);
not I_6791 (I117981,I117964);
nor I_6792 (I117998,I117933,I117981);
nor I_6793 (I118015,I117639,I117998);
DFFARX1 I_6794 (I118015,I2507,I117605,I117591,);
nor I_6795 (I118046,I117699,I117981);
nor I_6796 (I117579,I117894,I118046);
nor I_6797 (I117588,I117829,I117964);
nor I_6798 (I117576,I117699,I117964);
not I_6799 (I118132,I2514);
DFFARX1 I_6800 (I843890,I2507,I118132,I118158,);
not I_6801 (I118166,I118158);
nand I_6802 (I118183,I843887,I843902);
and I_6803 (I118200,I118183,I843884);
DFFARX1 I_6804 (I118200,I2507,I118132,I118226,);
DFFARX1 I_6805 (I843881,I2507,I118132,I118243,);
and I_6806 (I118251,I118243,I843881);
nor I_6807 (I118268,I118226,I118251);
DFFARX1 I_6808 (I118268,I2507,I118132,I118100,);
nand I_6809 (I118299,I118243,I843881);
nand I_6810 (I118316,I118166,I118299);
not I_6811 (I118112,I118316);
DFFARX1 I_6812 (I843884,I2507,I118132,I118356,);
DFFARX1 I_6813 (I118356,I2507,I118132,I118121,);
nand I_6814 (I118378,I843896,I843887);
and I_6815 (I118395,I118378,I843899);
DFFARX1 I_6816 (I118395,I2507,I118132,I118421,);
DFFARX1 I_6817 (I118421,I2507,I118132,I118438,);
not I_6818 (I118124,I118438);
not I_6819 (I118460,I118421);
nand I_6820 (I118109,I118460,I118299);
nor I_6821 (I118491,I843893,I843887);
not I_6822 (I118508,I118491);
nor I_6823 (I118525,I118460,I118508);
nor I_6824 (I118542,I118166,I118525);
DFFARX1 I_6825 (I118542,I2507,I118132,I118118,);
nor I_6826 (I118573,I118226,I118508);
nor I_6827 (I118106,I118421,I118573);
nor I_6828 (I118115,I118356,I118491);
nor I_6829 (I118103,I118226,I118491);
not I_6830 (I118659,I2514);
DFFARX1 I_6831 (I380513,I2507,I118659,I118685,);
not I_6832 (I118693,I118685);
nand I_6833 (I118710,I380507,I380498);
and I_6834 (I118727,I118710,I380519);
DFFARX1 I_6835 (I118727,I2507,I118659,I118753,);
DFFARX1 I_6836 (I380501,I2507,I118659,I118770,);
and I_6837 (I118778,I118770,I380495);
nor I_6838 (I118795,I118753,I118778);
DFFARX1 I_6839 (I118795,I2507,I118659,I118627,);
nand I_6840 (I118826,I118770,I380495);
nand I_6841 (I118843,I118693,I118826);
not I_6842 (I118639,I118843);
DFFARX1 I_6843 (I380495,I2507,I118659,I118883,);
DFFARX1 I_6844 (I118883,I2507,I118659,I118648,);
nand I_6845 (I118905,I380522,I380504);
and I_6846 (I118922,I118905,I380510);
DFFARX1 I_6847 (I118922,I2507,I118659,I118948,);
DFFARX1 I_6848 (I118948,I2507,I118659,I118965,);
not I_6849 (I118651,I118965);
not I_6850 (I118987,I118948);
nand I_6851 (I118636,I118987,I118826);
nor I_6852 (I119018,I380516,I380504);
not I_6853 (I119035,I119018);
nor I_6854 (I119052,I118987,I119035);
nor I_6855 (I119069,I118693,I119052);
DFFARX1 I_6856 (I119069,I2507,I118659,I118645,);
nor I_6857 (I119100,I118753,I119035);
nor I_6858 (I118633,I118948,I119100);
nor I_6859 (I118642,I118883,I119018);
nor I_6860 (I118630,I118753,I119018);
not I_6861 (I119186,I2514);
DFFARX1 I_6862 (I1192472,I2507,I119186,I119212,);
not I_6863 (I119220,I119212);
nand I_6864 (I119237,I1192487,I1192466);
and I_6865 (I119254,I119237,I1192469);
DFFARX1 I_6866 (I119254,I2507,I119186,I119280,);
DFFARX1 I_6867 (I1192490,I2507,I119186,I119297,);
and I_6868 (I119305,I119297,I1192469);
nor I_6869 (I119322,I119280,I119305);
DFFARX1 I_6870 (I119322,I2507,I119186,I119154,);
nand I_6871 (I119353,I119297,I1192469);
nand I_6872 (I119370,I119220,I119353);
not I_6873 (I119166,I119370);
DFFARX1 I_6874 (I1192466,I2507,I119186,I119410,);
DFFARX1 I_6875 (I119410,I2507,I119186,I119175,);
nand I_6876 (I119432,I1192478,I1192475);
and I_6877 (I119449,I119432,I1192481);
DFFARX1 I_6878 (I119449,I2507,I119186,I119475,);
DFFARX1 I_6879 (I119475,I2507,I119186,I119492,);
not I_6880 (I119178,I119492);
not I_6881 (I119514,I119475);
nand I_6882 (I119163,I119514,I119353);
nor I_6883 (I119545,I1192484,I1192475);
not I_6884 (I119562,I119545);
nor I_6885 (I119579,I119514,I119562);
nor I_6886 (I119596,I119220,I119579);
DFFARX1 I_6887 (I119596,I2507,I119186,I119172,);
nor I_6888 (I119627,I119280,I119562);
nor I_6889 (I119160,I119475,I119627);
nor I_6890 (I119169,I119410,I119545);
nor I_6891 (I119157,I119280,I119545);
not I_6892 (I119713,I2514);
DFFARX1 I_6893 (I300809,I2507,I119713,I119739,);
not I_6894 (I119747,I119739);
nand I_6895 (I119764,I300791,I300806);
and I_6896 (I119781,I119764,I300782);
DFFARX1 I_6897 (I119781,I2507,I119713,I119807,);
DFFARX1 I_6898 (I300785,I2507,I119713,I119824,);
and I_6899 (I119832,I119824,I300800);
nor I_6900 (I119849,I119807,I119832);
DFFARX1 I_6901 (I119849,I2507,I119713,I119681,);
nand I_6902 (I119880,I119824,I300800);
nand I_6903 (I119897,I119747,I119880);
not I_6904 (I119693,I119897);
DFFARX1 I_6905 (I300803,I2507,I119713,I119937,);
DFFARX1 I_6906 (I119937,I2507,I119713,I119702,);
nand I_6907 (I119959,I300782,I300794);
and I_6908 (I119976,I119959,I300788);
DFFARX1 I_6909 (I119976,I2507,I119713,I120002,);
DFFARX1 I_6910 (I120002,I2507,I119713,I120019,);
not I_6911 (I119705,I120019);
not I_6912 (I120041,I120002);
nand I_6913 (I119690,I120041,I119880);
nor I_6914 (I120072,I300797,I300794);
not I_6915 (I120089,I120072);
nor I_6916 (I120106,I120041,I120089);
nor I_6917 (I120123,I119747,I120106);
DFFARX1 I_6918 (I120123,I2507,I119713,I119699,);
nor I_6919 (I120154,I119807,I120089);
nor I_6920 (I119687,I120002,I120154);
nor I_6921 (I119696,I119937,I120072);
nor I_6922 (I119684,I119807,I120072);
not I_6923 (I120240,I2514);
DFFARX1 I_6924 (I503612,I2507,I120240,I120266,);
not I_6925 (I120274,I120266);
nand I_6926 (I120291,I503633,I503627);
and I_6927 (I120308,I120291,I503609);
DFFARX1 I_6928 (I120308,I2507,I120240,I120334,);
DFFARX1 I_6929 (I503612,I2507,I120240,I120351,);
and I_6930 (I120359,I120351,I503621);
nor I_6931 (I120376,I120334,I120359);
DFFARX1 I_6932 (I120376,I2507,I120240,I120208,);
nand I_6933 (I120407,I120351,I503621);
nand I_6934 (I120424,I120274,I120407);
not I_6935 (I120220,I120424);
DFFARX1 I_6936 (I503618,I2507,I120240,I120464,);
DFFARX1 I_6937 (I120464,I2507,I120240,I120229,);
nand I_6938 (I120486,I503624,I503615);
and I_6939 (I120503,I120486,I503609);
DFFARX1 I_6940 (I120503,I2507,I120240,I120529,);
DFFARX1 I_6941 (I120529,I2507,I120240,I120546,);
not I_6942 (I120232,I120546);
not I_6943 (I120568,I120529);
nand I_6944 (I120217,I120568,I120407);
nor I_6945 (I120599,I503630,I503615);
not I_6946 (I120616,I120599);
nor I_6947 (I120633,I120568,I120616);
nor I_6948 (I120650,I120274,I120633);
DFFARX1 I_6949 (I120650,I2507,I120240,I120226,);
nor I_6950 (I120681,I120334,I120616);
nor I_6951 (I120214,I120529,I120681);
nor I_6952 (I120223,I120464,I120599);
nor I_6953 (I120211,I120334,I120599);
not I_6954 (I120767,I2514);
DFFARX1 I_6955 (I375116,I2507,I120767,I120793,);
not I_6956 (I120801,I120793);
nand I_6957 (I120818,I375098,I375113);
and I_6958 (I120835,I120818,I375089);
DFFARX1 I_6959 (I120835,I2507,I120767,I120861,);
DFFARX1 I_6960 (I375092,I2507,I120767,I120878,);
and I_6961 (I120886,I120878,I375107);
nor I_6962 (I120903,I120861,I120886);
DFFARX1 I_6963 (I120903,I2507,I120767,I120735,);
nand I_6964 (I120934,I120878,I375107);
nand I_6965 (I120951,I120801,I120934);
not I_6966 (I120747,I120951);
DFFARX1 I_6967 (I375110,I2507,I120767,I120991,);
DFFARX1 I_6968 (I120991,I2507,I120767,I120756,);
nand I_6969 (I121013,I375089,I375101);
and I_6970 (I121030,I121013,I375095);
DFFARX1 I_6971 (I121030,I2507,I120767,I121056,);
DFFARX1 I_6972 (I121056,I2507,I120767,I121073,);
not I_6973 (I120759,I121073);
not I_6974 (I121095,I121056);
nand I_6975 (I120744,I121095,I120934);
nor I_6976 (I121126,I375104,I375101);
not I_6977 (I121143,I121126);
nor I_6978 (I121160,I121095,I121143);
nor I_6979 (I121177,I120801,I121160);
DFFARX1 I_6980 (I121177,I2507,I120767,I120753,);
nor I_6981 (I121208,I120861,I121143);
nor I_6982 (I120741,I121056,I121208);
nor I_6983 (I120750,I120991,I121126);
nor I_6984 (I120738,I120861,I121126);
not I_6985 (I121294,I2514);
DFFARX1 I_6986 (I812270,I2507,I121294,I121320,);
not I_6987 (I121328,I121320);
nand I_6988 (I121345,I812267,I812282);
and I_6989 (I121362,I121345,I812264);
DFFARX1 I_6990 (I121362,I2507,I121294,I121388,);
DFFARX1 I_6991 (I812261,I2507,I121294,I121405,);
and I_6992 (I121413,I121405,I812261);
nor I_6993 (I121430,I121388,I121413);
DFFARX1 I_6994 (I121430,I2507,I121294,I121262,);
nand I_6995 (I121461,I121405,I812261);
nand I_6996 (I121478,I121328,I121461);
not I_6997 (I121274,I121478);
DFFARX1 I_6998 (I812264,I2507,I121294,I121518,);
DFFARX1 I_6999 (I121518,I2507,I121294,I121283,);
nand I_7000 (I121540,I812276,I812267);
and I_7001 (I121557,I121540,I812279);
DFFARX1 I_7002 (I121557,I2507,I121294,I121583,);
DFFARX1 I_7003 (I121583,I2507,I121294,I121600,);
not I_7004 (I121286,I121600);
not I_7005 (I121622,I121583);
nand I_7006 (I121271,I121622,I121461);
nor I_7007 (I121653,I812273,I812267);
not I_7008 (I121670,I121653);
nor I_7009 (I121687,I121622,I121670);
nor I_7010 (I121704,I121328,I121687);
DFFARX1 I_7011 (I121704,I2507,I121294,I121280,);
nor I_7012 (I121735,I121388,I121670);
nor I_7013 (I121268,I121583,I121735);
nor I_7014 (I121277,I121518,I121653);
nor I_7015 (I121265,I121388,I121653);
not I_7016 (I121821,I2514);
DFFARX1 I_7017 (I800676,I2507,I121821,I121847,);
not I_7018 (I121855,I121847);
nand I_7019 (I121872,I800673,I800688);
and I_7020 (I121889,I121872,I800670);
DFFARX1 I_7021 (I121889,I2507,I121821,I121915,);
DFFARX1 I_7022 (I800667,I2507,I121821,I121932,);
and I_7023 (I121940,I121932,I800667);
nor I_7024 (I121957,I121915,I121940);
DFFARX1 I_7025 (I121957,I2507,I121821,I121789,);
nand I_7026 (I121988,I121932,I800667);
nand I_7027 (I122005,I121855,I121988);
not I_7028 (I121801,I122005);
DFFARX1 I_7029 (I800670,I2507,I121821,I122045,);
DFFARX1 I_7030 (I122045,I2507,I121821,I121810,);
nand I_7031 (I122067,I800682,I800673);
and I_7032 (I122084,I122067,I800685);
DFFARX1 I_7033 (I122084,I2507,I121821,I122110,);
DFFARX1 I_7034 (I122110,I2507,I121821,I122127,);
not I_7035 (I121813,I122127);
not I_7036 (I122149,I122110);
nand I_7037 (I121798,I122149,I121988);
nor I_7038 (I122180,I800679,I800673);
not I_7039 (I122197,I122180);
nor I_7040 (I122214,I122149,I122197);
nor I_7041 (I122231,I121855,I122214);
DFFARX1 I_7042 (I122231,I2507,I121821,I121807,);
nor I_7043 (I122262,I121915,I122197);
nor I_7044 (I121795,I122110,I122262);
nor I_7045 (I121804,I122045,I122180);
nor I_7046 (I121792,I121915,I122180);
not I_7047 (I122348,I2514);
DFFARX1 I_7048 (I1223752,I2507,I122348,I122374,);
not I_7049 (I122382,I122374);
nand I_7050 (I122399,I1223746,I1223767);
and I_7051 (I122416,I122399,I1223758);
DFFARX1 I_7052 (I122416,I2507,I122348,I122442,);
DFFARX1 I_7053 (I1223749,I2507,I122348,I122459,);
and I_7054 (I122467,I122459,I1223761);
nor I_7055 (I122484,I122442,I122467);
DFFARX1 I_7056 (I122484,I2507,I122348,I122316,);
nand I_7057 (I122515,I122459,I1223761);
nand I_7058 (I122532,I122382,I122515);
not I_7059 (I122328,I122532);
DFFARX1 I_7060 (I1223749,I2507,I122348,I122572,);
DFFARX1 I_7061 (I122572,I2507,I122348,I122337,);
nand I_7062 (I122594,I1223770,I1223755);
and I_7063 (I122611,I122594,I1223746);
DFFARX1 I_7064 (I122611,I2507,I122348,I122637,);
DFFARX1 I_7065 (I122637,I2507,I122348,I122654,);
not I_7066 (I122340,I122654);
not I_7067 (I122676,I122637);
nand I_7068 (I122325,I122676,I122515);
nor I_7069 (I122707,I1223764,I1223755);
not I_7070 (I122724,I122707);
nor I_7071 (I122741,I122676,I122724);
nor I_7072 (I122758,I122382,I122741);
DFFARX1 I_7073 (I122758,I2507,I122348,I122334,);
nor I_7074 (I122789,I122442,I122724);
nor I_7075 (I122322,I122637,I122789);
nor I_7076 (I122331,I122572,I122707);
nor I_7077 (I122319,I122442,I122707);
not I_7078 (I122875,I2514);
DFFARX1 I_7079 (I948950,I2507,I122875,I122901,);
not I_7080 (I122909,I122901);
nand I_7081 (I122926,I948968,I948962);
and I_7082 (I122943,I122926,I948941);
DFFARX1 I_7083 (I122943,I2507,I122875,I122969,);
DFFARX1 I_7084 (I948959,I2507,I122875,I122986,);
and I_7085 (I122994,I122986,I948944);
nor I_7086 (I123011,I122969,I122994);
DFFARX1 I_7087 (I123011,I2507,I122875,I122843,);
nand I_7088 (I123042,I122986,I948944);
nand I_7089 (I123059,I122909,I123042);
not I_7090 (I122855,I123059);
DFFARX1 I_7091 (I948956,I2507,I122875,I123099,);
DFFARX1 I_7092 (I123099,I2507,I122875,I122864,);
nand I_7093 (I123121,I948965,I948953);
and I_7094 (I123138,I123121,I948947);
DFFARX1 I_7095 (I123138,I2507,I122875,I123164,);
DFFARX1 I_7096 (I123164,I2507,I122875,I123181,);
not I_7097 (I122867,I123181);
not I_7098 (I123203,I123164);
nand I_7099 (I122852,I123203,I123042);
nor I_7100 (I123234,I948941,I948953);
not I_7101 (I123251,I123234);
nor I_7102 (I123268,I123203,I123251);
nor I_7103 (I123285,I122909,I123268);
DFFARX1 I_7104 (I123285,I2507,I122875,I122861,);
nor I_7105 (I123316,I122969,I123251);
nor I_7106 (I122849,I123164,I123316);
nor I_7107 (I122858,I123099,I123234);
nor I_7108 (I122846,I122969,I123234);
not I_7109 (I123402,I2514);
DFFARX1 I_7110 (I580441,I2507,I123402,I123428,);
not I_7111 (I123436,I123428);
nand I_7112 (I123453,I580453,I580438);
and I_7113 (I123470,I123453,I580432);
DFFARX1 I_7114 (I123470,I2507,I123402,I123496,);
DFFARX1 I_7115 (I580447,I2507,I123402,I123513,);
and I_7116 (I123521,I123513,I580435);
nor I_7117 (I123538,I123496,I123521);
DFFARX1 I_7118 (I123538,I2507,I123402,I123370,);
nand I_7119 (I123569,I123513,I580435);
nand I_7120 (I123586,I123436,I123569);
not I_7121 (I123382,I123586);
DFFARX1 I_7122 (I580444,I2507,I123402,I123626,);
DFFARX1 I_7123 (I123626,I2507,I123402,I123391,);
nand I_7124 (I123648,I580450,I580456);
and I_7125 (I123665,I123648,I580432);
DFFARX1 I_7126 (I123665,I2507,I123402,I123691,);
DFFARX1 I_7127 (I123691,I2507,I123402,I123708,);
not I_7128 (I123394,I123708);
not I_7129 (I123730,I123691);
nand I_7130 (I123379,I123730,I123569);
nor I_7131 (I123761,I580435,I580456);
not I_7132 (I123778,I123761);
nor I_7133 (I123795,I123730,I123778);
nor I_7134 (I123812,I123436,I123795);
DFFARX1 I_7135 (I123812,I2507,I123402,I123388,);
nor I_7136 (I123843,I123496,I123778);
nor I_7137 (I123376,I123691,I123843);
nor I_7138 (I123385,I123626,I123761);
nor I_7139 (I123373,I123496,I123761);
not I_7140 (I123929,I2514);
DFFARX1 I_7141 (I217477,I2507,I123929,I123955,);
not I_7142 (I123963,I123955);
nand I_7143 (I123980,I217471,I217465);
and I_7144 (I123997,I123980,I217486);
DFFARX1 I_7145 (I123997,I2507,I123929,I124023,);
DFFARX1 I_7146 (I217483,I2507,I123929,I124040,);
and I_7147 (I124048,I124040,I217480);
nor I_7148 (I124065,I124023,I124048);
DFFARX1 I_7149 (I124065,I2507,I123929,I123897,);
nand I_7150 (I124096,I124040,I217480);
nand I_7151 (I124113,I123963,I124096);
not I_7152 (I123909,I124113);
DFFARX1 I_7153 (I217465,I2507,I123929,I124153,);
DFFARX1 I_7154 (I124153,I2507,I123929,I123918,);
nand I_7155 (I124175,I217468,I217468);
and I_7156 (I124192,I124175,I217489);
DFFARX1 I_7157 (I124192,I2507,I123929,I124218,);
DFFARX1 I_7158 (I124218,I2507,I123929,I124235,);
not I_7159 (I123921,I124235);
not I_7160 (I124257,I124218);
nand I_7161 (I123906,I124257,I124096);
nor I_7162 (I124288,I217474,I217468);
not I_7163 (I124305,I124288);
nor I_7164 (I124322,I124257,I124305);
nor I_7165 (I124339,I123963,I124322);
DFFARX1 I_7166 (I124339,I2507,I123929,I123915,);
nor I_7167 (I124370,I124023,I124305);
nor I_7168 (I123903,I124218,I124370);
nor I_7169 (I123912,I124153,I124288);
nor I_7170 (I123900,I124023,I124288);
not I_7171 (I124456,I2514);
DFFARX1 I_7172 (I1031462,I2507,I124456,I124482,);
not I_7173 (I124490,I124482);
nand I_7174 (I124507,I1031459,I1031465);
and I_7175 (I124524,I124507,I1031462);
DFFARX1 I_7176 (I124524,I2507,I124456,I124550,);
DFFARX1 I_7177 (I1031465,I2507,I124456,I124567,);
and I_7178 (I124575,I124567,I1031459);
nor I_7179 (I124592,I124550,I124575);
DFFARX1 I_7180 (I124592,I2507,I124456,I124424,);
nand I_7181 (I124623,I124567,I1031459);
nand I_7182 (I124640,I124490,I124623);
not I_7183 (I124436,I124640);
DFFARX1 I_7184 (I1031468,I2507,I124456,I124680,);
DFFARX1 I_7185 (I124680,I2507,I124456,I124445,);
nand I_7186 (I124702,I1031471,I1031480);
and I_7187 (I124719,I124702,I1031474);
DFFARX1 I_7188 (I124719,I2507,I124456,I124745,);
DFFARX1 I_7189 (I124745,I2507,I124456,I124762,);
not I_7190 (I124448,I124762);
not I_7191 (I124784,I124745);
nand I_7192 (I124433,I124784,I124623);
nor I_7193 (I124815,I1031477,I1031480);
not I_7194 (I124832,I124815);
nor I_7195 (I124849,I124784,I124832);
nor I_7196 (I124866,I124490,I124849);
DFFARX1 I_7197 (I124866,I2507,I124456,I124442,);
nor I_7198 (I124897,I124550,I124832);
nor I_7199 (I124430,I124745,I124897);
nor I_7200 (I124439,I124680,I124815);
nor I_7201 (I124427,I124550,I124815);
not I_7202 (I124983,I2514);
DFFARX1 I_7203 (I878145,I2507,I124983,I125009,);
not I_7204 (I125017,I125009);
nand I_7205 (I125034,I878142,I878157);
and I_7206 (I125051,I125034,I878139);
DFFARX1 I_7207 (I125051,I2507,I124983,I125077,);
DFFARX1 I_7208 (I878136,I2507,I124983,I125094,);
and I_7209 (I125102,I125094,I878136);
nor I_7210 (I125119,I125077,I125102);
DFFARX1 I_7211 (I125119,I2507,I124983,I124951,);
nand I_7212 (I125150,I125094,I878136);
nand I_7213 (I125167,I125017,I125150);
not I_7214 (I124963,I125167);
DFFARX1 I_7215 (I878139,I2507,I124983,I125207,);
DFFARX1 I_7216 (I125207,I2507,I124983,I124972,);
nand I_7217 (I125229,I878151,I878142);
and I_7218 (I125246,I125229,I878154);
DFFARX1 I_7219 (I125246,I2507,I124983,I125272,);
DFFARX1 I_7220 (I125272,I2507,I124983,I125289,);
not I_7221 (I124975,I125289);
not I_7222 (I125311,I125272);
nand I_7223 (I124960,I125311,I125150);
nor I_7224 (I125342,I878148,I878142);
not I_7225 (I125359,I125342);
nor I_7226 (I125376,I125311,I125359);
nor I_7227 (I125393,I125017,I125376);
DFFARX1 I_7228 (I125393,I2507,I124983,I124969,);
nor I_7229 (I125424,I125077,I125359);
nor I_7230 (I124957,I125272,I125424);
nor I_7231 (I124966,I125207,I125342);
nor I_7232 (I124954,I125077,I125342);
not I_7233 (I125510,I2514);
DFFARX1 I_7234 (I671768,I2507,I125510,I125536,);
not I_7235 (I125544,I125536);
nand I_7236 (I125561,I671759,I671777);
and I_7237 (I125578,I125561,I671756);
DFFARX1 I_7238 (I125578,I2507,I125510,I125604,);
DFFARX1 I_7239 (I671759,I2507,I125510,I125621,);
and I_7240 (I125629,I125621,I671762);
nor I_7241 (I125646,I125604,I125629);
DFFARX1 I_7242 (I125646,I2507,I125510,I125478,);
nand I_7243 (I125677,I125621,I671762);
nand I_7244 (I125694,I125544,I125677);
not I_7245 (I125490,I125694);
DFFARX1 I_7246 (I671756,I2507,I125510,I125734,);
DFFARX1 I_7247 (I125734,I2507,I125510,I125499,);
nand I_7248 (I125756,I671774,I671765);
and I_7249 (I125773,I125756,I671780);
DFFARX1 I_7250 (I125773,I2507,I125510,I125799,);
DFFARX1 I_7251 (I125799,I2507,I125510,I125816,);
not I_7252 (I125502,I125816);
not I_7253 (I125838,I125799);
nand I_7254 (I125487,I125838,I125677);
nor I_7255 (I125869,I671771,I671765);
not I_7256 (I125886,I125869);
nor I_7257 (I125903,I125838,I125886);
nor I_7258 (I125920,I125544,I125903);
DFFARX1 I_7259 (I125920,I2507,I125510,I125496,);
nor I_7260 (I125951,I125604,I125886);
nor I_7261 (I125484,I125799,I125951);
nor I_7262 (I125493,I125734,I125869);
nor I_7263 (I125481,I125604,I125869);
not I_7264 (I126037,I2514);
DFFARX1 I_7265 (I418049,I2507,I126037,I126063,);
not I_7266 (I126071,I126063);
nand I_7267 (I126088,I418043,I418034);
and I_7268 (I126105,I126088,I418055);
DFFARX1 I_7269 (I126105,I2507,I126037,I126131,);
DFFARX1 I_7270 (I418037,I2507,I126037,I126148,);
and I_7271 (I126156,I126148,I418031);
nor I_7272 (I126173,I126131,I126156);
DFFARX1 I_7273 (I126173,I2507,I126037,I126005,);
nand I_7274 (I126204,I126148,I418031);
nand I_7275 (I126221,I126071,I126204);
not I_7276 (I126017,I126221);
DFFARX1 I_7277 (I418031,I2507,I126037,I126261,);
DFFARX1 I_7278 (I126261,I2507,I126037,I126026,);
nand I_7279 (I126283,I418058,I418040);
and I_7280 (I126300,I126283,I418046);
DFFARX1 I_7281 (I126300,I2507,I126037,I126326,);
DFFARX1 I_7282 (I126326,I2507,I126037,I126343,);
not I_7283 (I126029,I126343);
not I_7284 (I126365,I126326);
nand I_7285 (I126014,I126365,I126204);
nor I_7286 (I126396,I418052,I418040);
not I_7287 (I126413,I126396);
nor I_7288 (I126430,I126365,I126413);
nor I_7289 (I126447,I126071,I126430);
DFFARX1 I_7290 (I126447,I2507,I126037,I126023,);
nor I_7291 (I126478,I126131,I126413);
nor I_7292 (I126011,I126326,I126478);
nor I_7293 (I126020,I126261,I126396);
nor I_7294 (I126008,I126131,I126396);
not I_7295 (I126564,I2514);
DFFARX1 I_7296 (I1079762,I2507,I126564,I126590,);
not I_7297 (I126598,I126590);
nand I_7298 (I126615,I1079777,I1079756);
and I_7299 (I126632,I126615,I1079759);
DFFARX1 I_7300 (I126632,I2507,I126564,I126658,);
DFFARX1 I_7301 (I1079780,I2507,I126564,I126675,);
and I_7302 (I126683,I126675,I1079759);
nor I_7303 (I126700,I126658,I126683);
DFFARX1 I_7304 (I126700,I2507,I126564,I126532,);
nand I_7305 (I126731,I126675,I1079759);
nand I_7306 (I126748,I126598,I126731);
not I_7307 (I126544,I126748);
DFFARX1 I_7308 (I1079756,I2507,I126564,I126788,);
DFFARX1 I_7309 (I126788,I2507,I126564,I126553,);
nand I_7310 (I126810,I1079768,I1079765);
and I_7311 (I126827,I126810,I1079771);
DFFARX1 I_7312 (I126827,I2507,I126564,I126853,);
DFFARX1 I_7313 (I126853,I2507,I126564,I126870,);
not I_7314 (I126556,I126870);
not I_7315 (I126892,I126853);
nand I_7316 (I126541,I126892,I126731);
nor I_7317 (I126923,I1079774,I1079765);
not I_7318 (I126940,I126923);
nor I_7319 (I126957,I126892,I126940);
nor I_7320 (I126974,I126598,I126957);
DFFARX1 I_7321 (I126974,I2507,I126564,I126550,);
nor I_7322 (I127005,I126658,I126940);
nor I_7323 (I126538,I126853,I127005);
nor I_7324 (I126547,I126788,I126923);
nor I_7325 (I126535,I126658,I126923);
not I_7326 (I127091,I2514);
DFFARX1 I_7327 (I1291767,I2507,I127091,I127117,);
not I_7328 (I127125,I127117);
nand I_7329 (I127142,I1291770,I1291764);
and I_7330 (I127159,I127142,I1291761);
DFFARX1 I_7331 (I127159,I2507,I127091,I127185,);
DFFARX1 I_7332 (I1291746,I2507,I127091,I127202,);
and I_7333 (I127210,I127202,I1291755);
nor I_7334 (I127227,I127185,I127210);
DFFARX1 I_7335 (I127227,I2507,I127091,I127059,);
nand I_7336 (I127258,I127202,I1291755);
nand I_7337 (I127275,I127125,I127258);
not I_7338 (I127071,I127275);
DFFARX1 I_7339 (I1291746,I2507,I127091,I127315,);
DFFARX1 I_7340 (I127315,I2507,I127091,I127080,);
nand I_7341 (I127337,I1291749,I1291752);
and I_7342 (I127354,I127337,I1291758);
DFFARX1 I_7343 (I127354,I2507,I127091,I127380,);
DFFARX1 I_7344 (I127380,I2507,I127091,I127397,);
not I_7345 (I127083,I127397);
not I_7346 (I127419,I127380);
nand I_7347 (I127068,I127419,I127258);
nor I_7348 (I127450,I1291749,I1291752);
not I_7349 (I127467,I127450);
nor I_7350 (I127484,I127419,I127467);
nor I_7351 (I127501,I127125,I127484);
DFFARX1 I_7352 (I127501,I2507,I127091,I127077,);
nor I_7353 (I127532,I127185,I127467);
nor I_7354 (I127065,I127380,I127532);
nor I_7355 (I127074,I127315,I127450);
nor I_7356 (I127062,I127185,I127450);
not I_7357 (I127618,I2514);
DFFARX1 I_7358 (I494753,I2507,I127618,I127644,);
not I_7359 (I127652,I127644);
nand I_7360 (I127669,I494747,I494738);
and I_7361 (I127686,I127669,I494759);
DFFARX1 I_7362 (I127686,I2507,I127618,I127712,);
DFFARX1 I_7363 (I494741,I2507,I127618,I127729,);
and I_7364 (I127737,I127729,I494735);
nor I_7365 (I127754,I127712,I127737);
DFFARX1 I_7366 (I127754,I2507,I127618,I127586,);
nand I_7367 (I127785,I127729,I494735);
nand I_7368 (I127802,I127652,I127785);
not I_7369 (I127598,I127802);
DFFARX1 I_7370 (I494735,I2507,I127618,I127842,);
DFFARX1 I_7371 (I127842,I2507,I127618,I127607,);
nand I_7372 (I127864,I494762,I494744);
and I_7373 (I127881,I127864,I494750);
DFFARX1 I_7374 (I127881,I2507,I127618,I127907,);
DFFARX1 I_7375 (I127907,I2507,I127618,I127924,);
not I_7376 (I127610,I127924);
not I_7377 (I127946,I127907);
nand I_7378 (I127595,I127946,I127785);
nor I_7379 (I127977,I494756,I494744);
not I_7380 (I127994,I127977);
nor I_7381 (I128011,I127946,I127994);
nor I_7382 (I128028,I127652,I128011);
DFFARX1 I_7383 (I128028,I2507,I127618,I127604,);
nor I_7384 (I128059,I127712,I127994);
nor I_7385 (I127592,I127907,I128059);
nor I_7386 (I127601,I127842,I127977);
nor I_7387 (I127589,I127712,I127977);
not I_7388 (I128145,I2514);
DFFARX1 I_7389 (I235327,I2507,I128145,I128171,);
not I_7390 (I128179,I128171);
nand I_7391 (I128196,I235321,I235315);
and I_7392 (I128213,I128196,I235336);
DFFARX1 I_7393 (I128213,I2507,I128145,I128239,);
DFFARX1 I_7394 (I235333,I2507,I128145,I128256,);
and I_7395 (I128264,I128256,I235330);
nor I_7396 (I128281,I128239,I128264);
DFFARX1 I_7397 (I128281,I2507,I128145,I128113,);
nand I_7398 (I128312,I128256,I235330);
nand I_7399 (I128329,I128179,I128312);
not I_7400 (I128125,I128329);
DFFARX1 I_7401 (I235315,I2507,I128145,I128369,);
DFFARX1 I_7402 (I128369,I2507,I128145,I128134,);
nand I_7403 (I128391,I235318,I235318);
and I_7404 (I128408,I128391,I235339);
DFFARX1 I_7405 (I128408,I2507,I128145,I128434,);
DFFARX1 I_7406 (I128434,I2507,I128145,I128451,);
not I_7407 (I128137,I128451);
not I_7408 (I128473,I128434);
nand I_7409 (I128122,I128473,I128312);
nor I_7410 (I128504,I235324,I235318);
not I_7411 (I128521,I128504);
nor I_7412 (I128538,I128473,I128521);
nor I_7413 (I128555,I128179,I128538);
DFFARX1 I_7414 (I128555,I2507,I128145,I128131,);
nor I_7415 (I128586,I128239,I128521);
nor I_7416 (I128119,I128434,I128586);
nor I_7417 (I128128,I128369,I128504);
nor I_7418 (I128116,I128239,I128504);
not I_7419 (I128672,I2514);
DFFARX1 I_7420 (I16413,I2507,I128672,I128698,);
not I_7421 (I128706,I128698);
nand I_7422 (I128723,I16401,I16407);
and I_7423 (I128740,I128723,I16410);
DFFARX1 I_7424 (I128740,I2507,I128672,I128766,);
DFFARX1 I_7425 (I16392,I2507,I128672,I128783,);
and I_7426 (I128791,I128783,I16398);
nor I_7427 (I128808,I128766,I128791);
DFFARX1 I_7428 (I128808,I2507,I128672,I128640,);
nand I_7429 (I128839,I128783,I16398);
nand I_7430 (I128856,I128706,I128839);
not I_7431 (I128652,I128856);
DFFARX1 I_7432 (I16392,I2507,I128672,I128896,);
DFFARX1 I_7433 (I128896,I2507,I128672,I128661,);
nand I_7434 (I128918,I16395,I16389);
and I_7435 (I128935,I128918,I16404);
DFFARX1 I_7436 (I128935,I2507,I128672,I128961,);
DFFARX1 I_7437 (I128961,I2507,I128672,I128978,);
not I_7438 (I128664,I128978);
not I_7439 (I129000,I128961);
nand I_7440 (I128649,I129000,I128839);
nor I_7441 (I129031,I16389,I16389);
not I_7442 (I129048,I129031);
nor I_7443 (I129065,I129000,I129048);
nor I_7444 (I129082,I128706,I129065);
DFFARX1 I_7445 (I129082,I2507,I128672,I128658,);
nor I_7446 (I129113,I128766,I129048);
nor I_7447 (I128646,I128961,I129113);
nor I_7448 (I128655,I128896,I129031);
nor I_7449 (I128643,I128766,I129031);
not I_7450 (I129199,I2514);
DFFARX1 I_7451 (I798041,I2507,I129199,I129225,);
not I_7452 (I129233,I129225);
nand I_7453 (I129250,I798038,I798053);
and I_7454 (I129267,I129250,I798035);
DFFARX1 I_7455 (I129267,I2507,I129199,I129293,);
DFFARX1 I_7456 (I798032,I2507,I129199,I129310,);
and I_7457 (I129318,I129310,I798032);
nor I_7458 (I129335,I129293,I129318);
DFFARX1 I_7459 (I129335,I2507,I129199,I129167,);
nand I_7460 (I129366,I129310,I798032);
nand I_7461 (I129383,I129233,I129366);
not I_7462 (I129179,I129383);
DFFARX1 I_7463 (I798035,I2507,I129199,I129423,);
DFFARX1 I_7464 (I129423,I2507,I129199,I129188,);
nand I_7465 (I129445,I798047,I798038);
and I_7466 (I129462,I129445,I798050);
DFFARX1 I_7467 (I129462,I2507,I129199,I129488,);
DFFARX1 I_7468 (I129488,I2507,I129199,I129505,);
not I_7469 (I129191,I129505);
not I_7470 (I129527,I129488);
nand I_7471 (I129176,I129527,I129366);
nor I_7472 (I129558,I798044,I798038);
not I_7473 (I129575,I129558);
nor I_7474 (I129592,I129527,I129575);
nor I_7475 (I129609,I129233,I129592);
DFFARX1 I_7476 (I129609,I2507,I129199,I129185,);
nor I_7477 (I129640,I129293,I129575);
nor I_7478 (I129173,I129488,I129640);
nor I_7479 (I129182,I129423,I129558);
nor I_7480 (I129170,I129293,I129558);
not I_7481 (I129726,I2514);
DFFARX1 I_7482 (I753266,I2507,I129726,I129752,);
not I_7483 (I129760,I129752);
nand I_7484 (I129777,I753257,I753275);
and I_7485 (I129794,I129777,I753254);
DFFARX1 I_7486 (I129794,I2507,I129726,I129820,);
DFFARX1 I_7487 (I753257,I2507,I129726,I129837,);
and I_7488 (I129845,I129837,I753260);
nor I_7489 (I129862,I129820,I129845);
DFFARX1 I_7490 (I129862,I2507,I129726,I129694,);
nand I_7491 (I129893,I129837,I753260);
nand I_7492 (I129910,I129760,I129893);
not I_7493 (I129706,I129910);
DFFARX1 I_7494 (I753254,I2507,I129726,I129950,);
DFFARX1 I_7495 (I129950,I2507,I129726,I129715,);
nand I_7496 (I129972,I753272,I753263);
and I_7497 (I129989,I129972,I753278);
DFFARX1 I_7498 (I129989,I2507,I129726,I130015,);
DFFARX1 I_7499 (I130015,I2507,I129726,I130032,);
not I_7500 (I129718,I130032);
not I_7501 (I130054,I130015);
nand I_7502 (I129703,I130054,I129893);
nor I_7503 (I130085,I753269,I753263);
not I_7504 (I130102,I130085);
nor I_7505 (I130119,I130054,I130102);
nor I_7506 (I130136,I129760,I130119);
DFFARX1 I_7507 (I130136,I2507,I129726,I129712,);
nor I_7508 (I130167,I129820,I130102);
nor I_7509 (I129700,I130015,I130167);
nor I_7510 (I129709,I129950,I130085);
nor I_7511 (I129697,I129820,I130085);
not I_7512 (I130253,I2514);
DFFARX1 I_7513 (I1064156,I2507,I130253,I130279,);
not I_7514 (I130287,I130279);
nand I_7515 (I130304,I1064171,I1064150);
and I_7516 (I130321,I130304,I1064153);
DFFARX1 I_7517 (I130321,I2507,I130253,I130347,);
DFFARX1 I_7518 (I1064174,I2507,I130253,I130364,);
and I_7519 (I130372,I130364,I1064153);
nor I_7520 (I130389,I130347,I130372);
DFFARX1 I_7521 (I130389,I2507,I130253,I130221,);
nand I_7522 (I130420,I130364,I1064153);
nand I_7523 (I130437,I130287,I130420);
not I_7524 (I130233,I130437);
DFFARX1 I_7525 (I1064150,I2507,I130253,I130477,);
DFFARX1 I_7526 (I130477,I2507,I130253,I130242,);
nand I_7527 (I130499,I1064162,I1064159);
and I_7528 (I130516,I130499,I1064165);
DFFARX1 I_7529 (I130516,I2507,I130253,I130542,);
DFFARX1 I_7530 (I130542,I2507,I130253,I130559,);
not I_7531 (I130245,I130559);
not I_7532 (I130581,I130542);
nand I_7533 (I130230,I130581,I130420);
nor I_7534 (I130612,I1064168,I1064159);
not I_7535 (I130629,I130612);
nor I_7536 (I130646,I130581,I130629);
nor I_7537 (I130663,I130287,I130646);
DFFARX1 I_7538 (I130663,I2507,I130253,I130239,);
nor I_7539 (I130694,I130347,I130629);
nor I_7540 (I130227,I130542,I130694);
nor I_7541 (I130236,I130477,I130612);
nor I_7542 (I130224,I130347,I130612);
not I_7543 (I130780,I2514);
DFFARX1 I_7544 (I1209064,I2507,I130780,I130806,);
not I_7545 (I130814,I130806);
nand I_7546 (I130831,I1209058,I1209079);
and I_7547 (I130848,I130831,I1209070);
DFFARX1 I_7548 (I130848,I2507,I130780,I130874,);
DFFARX1 I_7549 (I1209061,I2507,I130780,I130891,);
and I_7550 (I130899,I130891,I1209073);
nor I_7551 (I130916,I130874,I130899);
DFFARX1 I_7552 (I130916,I2507,I130780,I130748,);
nand I_7553 (I130947,I130891,I1209073);
nand I_7554 (I130964,I130814,I130947);
not I_7555 (I130760,I130964);
DFFARX1 I_7556 (I1209061,I2507,I130780,I131004,);
DFFARX1 I_7557 (I131004,I2507,I130780,I130769,);
nand I_7558 (I131026,I1209082,I1209067);
and I_7559 (I131043,I131026,I1209058);
DFFARX1 I_7560 (I131043,I2507,I130780,I131069,);
DFFARX1 I_7561 (I131069,I2507,I130780,I131086,);
not I_7562 (I130772,I131086);
not I_7563 (I131108,I131069);
nand I_7564 (I130757,I131108,I130947);
nor I_7565 (I131139,I1209076,I1209067);
not I_7566 (I131156,I131139);
nor I_7567 (I131173,I131108,I131156);
nor I_7568 (I131190,I130814,I131173);
DFFARX1 I_7569 (I131190,I2507,I130780,I130766,);
nor I_7570 (I131221,I130874,I131156);
nor I_7571 (I130754,I131069,I131221);
nor I_7572 (I130763,I131004,I131139);
nor I_7573 (I130751,I130874,I131139);
not I_7574 (I131307,I2514);
DFFARX1 I_7575 (I21156,I2507,I131307,I131333,);
not I_7576 (I131341,I131333);
nand I_7577 (I131358,I21144,I21150);
and I_7578 (I131375,I131358,I21153);
DFFARX1 I_7579 (I131375,I2507,I131307,I131401,);
DFFARX1 I_7580 (I21135,I2507,I131307,I131418,);
and I_7581 (I131426,I131418,I21141);
nor I_7582 (I131443,I131401,I131426);
DFFARX1 I_7583 (I131443,I2507,I131307,I131275,);
nand I_7584 (I131474,I131418,I21141);
nand I_7585 (I131491,I131341,I131474);
not I_7586 (I131287,I131491);
DFFARX1 I_7587 (I21135,I2507,I131307,I131531,);
DFFARX1 I_7588 (I131531,I2507,I131307,I131296,);
nand I_7589 (I131553,I21138,I21132);
and I_7590 (I131570,I131553,I21147);
DFFARX1 I_7591 (I131570,I2507,I131307,I131596,);
DFFARX1 I_7592 (I131596,I2507,I131307,I131613,);
not I_7593 (I131299,I131613);
not I_7594 (I131635,I131596);
nand I_7595 (I131284,I131635,I131474);
nor I_7596 (I131666,I21132,I21132);
not I_7597 (I131683,I131666);
nor I_7598 (I131700,I131635,I131683);
nor I_7599 (I131717,I131341,I131700);
DFFARX1 I_7600 (I131717,I2507,I131307,I131293,);
nor I_7601 (I131748,I131401,I131683);
nor I_7602 (I131281,I131596,I131748);
nor I_7603 (I131290,I131531,I131666);
nor I_7604 (I131278,I131401,I131666);
not I_7605 (I131834,I2514);
DFFARX1 I_7606 (I1353519,I2507,I131834,I131860,);
not I_7607 (I131868,I131860);
nand I_7608 (I131885,I1353513,I1353534);
and I_7609 (I131902,I131885,I1353510);
DFFARX1 I_7610 (I131902,I2507,I131834,I131928,);
DFFARX1 I_7611 (I1353531,I2507,I131834,I131945,);
and I_7612 (I131953,I131945,I1353528);
nor I_7613 (I131970,I131928,I131953);
DFFARX1 I_7614 (I131970,I2507,I131834,I131802,);
nand I_7615 (I132001,I131945,I1353528);
nand I_7616 (I132018,I131868,I132001);
not I_7617 (I131814,I132018);
DFFARX1 I_7618 (I1353516,I2507,I131834,I132058,);
DFFARX1 I_7619 (I132058,I2507,I131834,I131823,);
nand I_7620 (I132080,I1353525,I1353522);
and I_7621 (I132097,I132080,I1353507);
DFFARX1 I_7622 (I132097,I2507,I131834,I132123,);
DFFARX1 I_7623 (I132123,I2507,I131834,I132140,);
not I_7624 (I131826,I132140);
not I_7625 (I132162,I132123);
nand I_7626 (I131811,I132162,I132001);
nor I_7627 (I132193,I1353507,I1353522);
not I_7628 (I132210,I132193);
nor I_7629 (I132227,I132162,I132210);
nor I_7630 (I132244,I131868,I132227);
DFFARX1 I_7631 (I132244,I2507,I131834,I131820,);
nor I_7632 (I132275,I131928,I132210);
nor I_7633 (I131808,I132123,I132275);
nor I_7634 (I131817,I132058,I132193);
nor I_7635 (I131805,I131928,I132193);
not I_7636 (I132361,I2514);
DFFARX1 I_7637 (I596047,I2507,I132361,I132387,);
not I_7638 (I132395,I132387);
nand I_7639 (I132412,I596059,I596044);
and I_7640 (I132429,I132412,I596038);
DFFARX1 I_7641 (I132429,I2507,I132361,I132455,);
DFFARX1 I_7642 (I596053,I2507,I132361,I132472,);
and I_7643 (I132480,I132472,I596041);
nor I_7644 (I132497,I132455,I132480);
DFFARX1 I_7645 (I132497,I2507,I132361,I132329,);
nand I_7646 (I132528,I132472,I596041);
nand I_7647 (I132545,I132395,I132528);
not I_7648 (I132341,I132545);
DFFARX1 I_7649 (I596050,I2507,I132361,I132585,);
DFFARX1 I_7650 (I132585,I2507,I132361,I132350,);
nand I_7651 (I132607,I596056,I596062);
and I_7652 (I132624,I132607,I596038);
DFFARX1 I_7653 (I132624,I2507,I132361,I132650,);
DFFARX1 I_7654 (I132650,I2507,I132361,I132667,);
not I_7655 (I132353,I132667);
not I_7656 (I132689,I132650);
nand I_7657 (I132338,I132689,I132528);
nor I_7658 (I132720,I596041,I596062);
not I_7659 (I132737,I132720);
nor I_7660 (I132754,I132689,I132737);
nor I_7661 (I132771,I132395,I132754);
DFFARX1 I_7662 (I132771,I2507,I132361,I132347,);
nor I_7663 (I132802,I132455,I132737);
nor I_7664 (I132335,I132650,I132802);
nor I_7665 (I132344,I132585,I132720);
nor I_7666 (I132332,I132455,I132720);
not I_7667 (I132888,I2514);
DFFARX1 I_7668 (I1098836,I2507,I132888,I132914,);
not I_7669 (I132922,I132914);
nand I_7670 (I132939,I1098851,I1098830);
and I_7671 (I132956,I132939,I1098833);
DFFARX1 I_7672 (I132956,I2507,I132888,I132982,);
DFFARX1 I_7673 (I1098854,I2507,I132888,I132999,);
and I_7674 (I133007,I132999,I1098833);
nor I_7675 (I133024,I132982,I133007);
DFFARX1 I_7676 (I133024,I2507,I132888,I132856,);
nand I_7677 (I133055,I132999,I1098833);
nand I_7678 (I133072,I132922,I133055);
not I_7679 (I132868,I133072);
DFFARX1 I_7680 (I1098830,I2507,I132888,I133112,);
DFFARX1 I_7681 (I133112,I2507,I132888,I132877,);
nand I_7682 (I133134,I1098842,I1098839);
and I_7683 (I133151,I133134,I1098845);
DFFARX1 I_7684 (I133151,I2507,I132888,I133177,);
DFFARX1 I_7685 (I133177,I2507,I132888,I133194,);
not I_7686 (I132880,I133194);
not I_7687 (I133216,I133177);
nand I_7688 (I132865,I133216,I133055);
nor I_7689 (I133247,I1098848,I1098839);
not I_7690 (I133264,I133247);
nor I_7691 (I133281,I133216,I133264);
nor I_7692 (I133298,I132922,I133281);
DFFARX1 I_7693 (I133298,I2507,I132888,I132874,);
nor I_7694 (I133329,I132982,I133264);
nor I_7695 (I132862,I133177,I133329);
nor I_7696 (I132871,I133112,I133247);
nor I_7697 (I132859,I132982,I133247);
not I_7698 (I133415,I2514);
DFFARX1 I_7699 (I864443,I2507,I133415,I133441,);
not I_7700 (I133449,I133441);
nand I_7701 (I133466,I864440,I864455);
and I_7702 (I133483,I133466,I864437);
DFFARX1 I_7703 (I133483,I2507,I133415,I133509,);
DFFARX1 I_7704 (I864434,I2507,I133415,I133526,);
and I_7705 (I133534,I133526,I864434);
nor I_7706 (I133551,I133509,I133534);
DFFARX1 I_7707 (I133551,I2507,I133415,I133383,);
nand I_7708 (I133582,I133526,I864434);
nand I_7709 (I133599,I133449,I133582);
not I_7710 (I133395,I133599);
DFFARX1 I_7711 (I864437,I2507,I133415,I133639,);
DFFARX1 I_7712 (I133639,I2507,I133415,I133404,);
nand I_7713 (I133661,I864449,I864440);
and I_7714 (I133678,I133661,I864452);
DFFARX1 I_7715 (I133678,I2507,I133415,I133704,);
DFFARX1 I_7716 (I133704,I2507,I133415,I133721,);
not I_7717 (I133407,I133721);
not I_7718 (I133743,I133704);
nand I_7719 (I133392,I133743,I133582);
nor I_7720 (I133774,I864446,I864440);
not I_7721 (I133791,I133774);
nor I_7722 (I133808,I133743,I133791);
nor I_7723 (I133825,I133449,I133808);
DFFARX1 I_7724 (I133825,I2507,I133415,I133401,);
nor I_7725 (I133856,I133509,I133791);
nor I_7726 (I133389,I133704,I133856);
nor I_7727 (I133398,I133639,I133774);
nor I_7728 (I133386,I133509,I133774);
not I_7729 (I133942,I2514);
DFFARX1 I_7730 (I956056,I2507,I133942,I133968,);
not I_7731 (I133976,I133968);
nand I_7732 (I133993,I956074,I956068);
and I_7733 (I134010,I133993,I956047);
DFFARX1 I_7734 (I134010,I2507,I133942,I134036,);
DFFARX1 I_7735 (I956065,I2507,I133942,I134053,);
and I_7736 (I134061,I134053,I956050);
nor I_7737 (I134078,I134036,I134061);
DFFARX1 I_7738 (I134078,I2507,I133942,I133910,);
nand I_7739 (I134109,I134053,I956050);
nand I_7740 (I134126,I133976,I134109);
not I_7741 (I133922,I134126);
DFFARX1 I_7742 (I956062,I2507,I133942,I134166,);
DFFARX1 I_7743 (I134166,I2507,I133942,I133931,);
nand I_7744 (I134188,I956071,I956059);
and I_7745 (I134205,I134188,I956053);
DFFARX1 I_7746 (I134205,I2507,I133942,I134231,);
DFFARX1 I_7747 (I134231,I2507,I133942,I134248,);
not I_7748 (I133934,I134248);
not I_7749 (I134270,I134231);
nand I_7750 (I133919,I134270,I134109);
nor I_7751 (I134301,I956047,I956059);
not I_7752 (I134318,I134301);
nor I_7753 (I134335,I134270,I134318);
nor I_7754 (I134352,I133976,I134335);
DFFARX1 I_7755 (I134352,I2507,I133942,I133928,);
nor I_7756 (I134383,I134036,I134318);
nor I_7757 (I133916,I134231,I134383);
nor I_7758 (I133925,I134166,I134301);
nor I_7759 (I133913,I134036,I134301);
not I_7760 (I134469,I2514);
DFFARX1 I_7761 (I1112708,I2507,I134469,I134495,);
not I_7762 (I134503,I134495);
nand I_7763 (I134520,I1112723,I1112702);
and I_7764 (I134537,I134520,I1112705);
DFFARX1 I_7765 (I134537,I2507,I134469,I134563,);
DFFARX1 I_7766 (I1112726,I2507,I134469,I134580,);
and I_7767 (I134588,I134580,I1112705);
nor I_7768 (I134605,I134563,I134588);
DFFARX1 I_7769 (I134605,I2507,I134469,I134437,);
nand I_7770 (I134636,I134580,I1112705);
nand I_7771 (I134653,I134503,I134636);
not I_7772 (I134449,I134653);
DFFARX1 I_7773 (I1112702,I2507,I134469,I134693,);
DFFARX1 I_7774 (I134693,I2507,I134469,I134458,);
nand I_7775 (I134715,I1112714,I1112711);
and I_7776 (I134732,I134715,I1112717);
DFFARX1 I_7777 (I134732,I2507,I134469,I134758,);
DFFARX1 I_7778 (I134758,I2507,I134469,I134775,);
not I_7779 (I134461,I134775);
not I_7780 (I134797,I134758);
nand I_7781 (I134446,I134797,I134636);
nor I_7782 (I134828,I1112720,I1112711);
not I_7783 (I134845,I134828);
nor I_7784 (I134862,I134797,I134845);
nor I_7785 (I134879,I134503,I134862);
DFFARX1 I_7786 (I134879,I2507,I134469,I134455,);
nor I_7787 (I134910,I134563,I134845);
nor I_7788 (I134443,I134758,I134910);
nor I_7789 (I134452,I134693,I134828);
nor I_7790 (I134440,I134563,I134828);
not I_7791 (I134996,I2514);
DFFARX1 I_7792 (I549229,I2507,I134996,I135022,);
not I_7793 (I135030,I135022);
nand I_7794 (I135047,I549241,I549226);
and I_7795 (I135064,I135047,I549220);
DFFARX1 I_7796 (I135064,I2507,I134996,I135090,);
DFFARX1 I_7797 (I549235,I2507,I134996,I135107,);
and I_7798 (I135115,I135107,I549223);
nor I_7799 (I135132,I135090,I135115);
DFFARX1 I_7800 (I135132,I2507,I134996,I134964,);
nand I_7801 (I135163,I135107,I549223);
nand I_7802 (I135180,I135030,I135163);
not I_7803 (I134976,I135180);
DFFARX1 I_7804 (I549232,I2507,I134996,I135220,);
DFFARX1 I_7805 (I135220,I2507,I134996,I134985,);
nand I_7806 (I135242,I549238,I549244);
and I_7807 (I135259,I135242,I549220);
DFFARX1 I_7808 (I135259,I2507,I134996,I135285,);
DFFARX1 I_7809 (I135285,I2507,I134996,I135302,);
not I_7810 (I134988,I135302);
not I_7811 (I135324,I135285);
nand I_7812 (I134973,I135324,I135163);
nor I_7813 (I135355,I549223,I549244);
not I_7814 (I135372,I135355);
nor I_7815 (I135389,I135324,I135372);
nor I_7816 (I135406,I135030,I135389);
DFFARX1 I_7817 (I135406,I2507,I134996,I134982,);
nor I_7818 (I135437,I135090,I135372);
nor I_7819 (I134970,I135285,I135437);
nor I_7820 (I134979,I135220,I135355);
nor I_7821 (I134967,I135090,I135355);
not I_7822 (I135523,I2514);
DFFARX1 I_7823 (I365630,I2507,I135523,I135549,);
not I_7824 (I135557,I135549);
nand I_7825 (I135574,I365612,I365627);
and I_7826 (I135591,I135574,I365603);
DFFARX1 I_7827 (I135591,I2507,I135523,I135617,);
DFFARX1 I_7828 (I365606,I2507,I135523,I135634,);
and I_7829 (I135642,I135634,I365621);
nor I_7830 (I135659,I135617,I135642);
DFFARX1 I_7831 (I135659,I2507,I135523,I135491,);
nand I_7832 (I135690,I135634,I365621);
nand I_7833 (I135707,I135557,I135690);
not I_7834 (I135503,I135707);
DFFARX1 I_7835 (I365624,I2507,I135523,I135747,);
DFFARX1 I_7836 (I135747,I2507,I135523,I135512,);
nand I_7837 (I135769,I365603,I365615);
and I_7838 (I135786,I135769,I365609);
DFFARX1 I_7839 (I135786,I2507,I135523,I135812,);
DFFARX1 I_7840 (I135812,I2507,I135523,I135829,);
not I_7841 (I135515,I135829);
not I_7842 (I135851,I135812);
nand I_7843 (I135500,I135851,I135690);
nor I_7844 (I135882,I365618,I365615);
not I_7845 (I135899,I135882);
nor I_7846 (I135916,I135851,I135899);
nor I_7847 (I135933,I135557,I135916);
DFFARX1 I_7848 (I135933,I2507,I135523,I135509,);
nor I_7849 (I135964,I135617,I135899);
nor I_7850 (I135497,I135812,I135964);
nor I_7851 (I135506,I135747,I135882);
nor I_7852 (I135494,I135617,I135882);
not I_7853 (I136050,I2514);
DFFARX1 I_7854 (I605873,I2507,I136050,I136076,);
not I_7855 (I136084,I136076);
nand I_7856 (I136101,I605885,I605870);
and I_7857 (I136118,I136101,I605864);
DFFARX1 I_7858 (I136118,I2507,I136050,I136144,);
DFFARX1 I_7859 (I605879,I2507,I136050,I136161,);
and I_7860 (I136169,I136161,I605867);
nor I_7861 (I136186,I136144,I136169);
DFFARX1 I_7862 (I136186,I2507,I136050,I136018,);
nand I_7863 (I136217,I136161,I605867);
nand I_7864 (I136234,I136084,I136217);
not I_7865 (I136030,I136234);
DFFARX1 I_7866 (I605876,I2507,I136050,I136274,);
DFFARX1 I_7867 (I136274,I2507,I136050,I136039,);
nand I_7868 (I136296,I605882,I605888);
and I_7869 (I136313,I136296,I605864);
DFFARX1 I_7870 (I136313,I2507,I136050,I136339,);
DFFARX1 I_7871 (I136339,I2507,I136050,I136356,);
not I_7872 (I136042,I136356);
not I_7873 (I136378,I136339);
nand I_7874 (I136027,I136378,I136217);
nor I_7875 (I136409,I605867,I605888);
not I_7876 (I136426,I136409);
nor I_7877 (I136443,I136378,I136426);
nor I_7878 (I136460,I136084,I136443);
DFFARX1 I_7879 (I136460,I2507,I136050,I136036,);
nor I_7880 (I136491,I136144,I136426);
nor I_7881 (I136024,I136339,I136491);
nor I_7882 (I136033,I136274,I136409);
nor I_7883 (I136021,I136144,I136409);
not I_7884 (I136580,I2514);
DFFARX1 I_7885 (I460487,I2507,I136580,I136606,);
not I_7886 (I136614,I136606);
DFFARX1 I_7887 (I460481,I2507,I136580,I136640,);
not I_7888 (I136648,I460478);
or I_7889 (I136665,I460469,I460478);
nor I_7890 (I136682,I136640,I460469);
nand I_7891 (I136557,I136648,I136682);
nor I_7892 (I136713,I460472,I460469);
nand I_7893 (I136551,I136713,I136648);
not I_7894 (I136744,I460475);
nand I_7895 (I136761,I136648,I136744);
nor I_7896 (I136778,I460463,I460490);
not I_7897 (I136795,I136778);
nor I_7898 (I136812,I136795,I136761);
nor I_7899 (I136829,I136713,I136812);
DFFARX1 I_7900 (I136829,I2507,I136580,I136566,);
nor I_7901 (I136563,I136778,I136665);
DFFARX1 I_7902 (I136778,I2507,I136580,I136569,);
nor I_7903 (I136888,I136744,I460463);
nor I_7904 (I136905,I136888,I460478);
nor I_7905 (I136922,I460466,I460463);
DFFARX1 I_7906 (I136922,I2507,I136580,I136948,);
nor I_7907 (I136548,I136948,I136905);
DFFARX1 I_7908 (I136948,I2507,I136580,I136979,);
nand I_7909 (I136987,I136979,I460484);
nor I_7910 (I136572,I136614,I136987);
not I_7911 (I137018,I136948);
nand I_7912 (I137035,I137018,I460484);
nor I_7913 (I137052,I136614,I137035);
nor I_7914 (I136554,I136640,I137052);
nor I_7915 (I137083,I460466,I460472);
nor I_7916 (I137100,I136640,I137083);
DFFARX1 I_7917 (I137100,I2507,I136580,I136545,);
and I_7918 (I136560,I136713,I460466);
not I_7919 (I137175,I2514);
DFFARX1 I_7920 (I197259,I2507,I137175,I137201,);
not I_7921 (I137209,I137201);
DFFARX1 I_7922 (I197253,I2507,I137175,I137235,);
not I_7923 (I137243,I197238);
or I_7924 (I137260,I197247,I197238);
nor I_7925 (I137277,I137235,I197247);
nand I_7926 (I137152,I137243,I137277);
nor I_7927 (I137308,I197235,I197247);
nand I_7928 (I137146,I137308,I137243);
not I_7929 (I137339,I197241);
nand I_7930 (I137356,I137243,I137339);
nor I_7931 (I137373,I197244,I197256);
not I_7932 (I137390,I137373);
nor I_7933 (I137407,I137390,I137356);
nor I_7934 (I137424,I137308,I137407);
DFFARX1 I_7935 (I137424,I2507,I137175,I137161,);
nor I_7936 (I137158,I137373,I137260);
DFFARX1 I_7937 (I137373,I2507,I137175,I137164,);
nor I_7938 (I137483,I137339,I197244);
nor I_7939 (I137500,I137483,I197238);
nor I_7940 (I137517,I197250,I197238);
DFFARX1 I_7941 (I137517,I2507,I137175,I137543,);
nor I_7942 (I137143,I137543,I137500);
DFFARX1 I_7943 (I137543,I2507,I137175,I137574,);
nand I_7944 (I137582,I137574,I197235);
nor I_7945 (I137167,I137209,I137582);
not I_7946 (I137613,I137543);
nand I_7947 (I137630,I137613,I197235);
nor I_7948 (I137647,I137209,I137630);
nor I_7949 (I137149,I137235,I137647);
nor I_7950 (I137678,I197250,I197235);
nor I_7951 (I137695,I137235,I137678);
DFFARX1 I_7952 (I137695,I2507,I137175,I137140,);
and I_7953 (I137155,I137308,I197250);
not I_7954 (I137770,I2514);
DFFARX1 I_7955 (I526231,I2507,I137770,I137796,);
not I_7956 (I137804,I137796);
DFFARX1 I_7957 (I526237,I2507,I137770,I137830,);
not I_7958 (I137838,I526219);
or I_7959 (I137855,I526243,I526219);
nor I_7960 (I137872,I137830,I526243);
nand I_7961 (I137747,I137838,I137872);
nor I_7962 (I137903,I526234,I526243);
nand I_7963 (I137741,I137903,I137838);
not I_7964 (I137934,I526225);
nand I_7965 (I137951,I137838,I137934);
nor I_7966 (I137968,I526228,I526222);
not I_7967 (I137985,I137968);
nor I_7968 (I138002,I137985,I137951);
nor I_7969 (I138019,I137903,I138002);
DFFARX1 I_7970 (I138019,I2507,I137770,I137756,);
nor I_7971 (I137753,I137968,I137855);
DFFARX1 I_7972 (I137968,I2507,I137770,I137759,);
nor I_7973 (I138078,I137934,I526228);
nor I_7974 (I138095,I138078,I526219);
nor I_7975 (I138112,I526240,I526219);
DFFARX1 I_7976 (I138112,I2507,I137770,I138138,);
nor I_7977 (I137738,I138138,I138095);
DFFARX1 I_7978 (I138138,I2507,I137770,I138169,);
nand I_7979 (I138177,I138169,I526222);
nor I_7980 (I137762,I137804,I138177);
not I_7981 (I138208,I138138);
nand I_7982 (I138225,I138208,I526222);
nor I_7983 (I138242,I137804,I138225);
nor I_7984 (I137744,I137830,I138242);
nor I_7985 (I138273,I526240,I526234);
nor I_7986 (I138290,I137830,I138273);
DFFARX1 I_7987 (I138290,I2507,I137770,I137735,);
and I_7988 (I137750,I137903,I526240);
not I_7989 (I138365,I2514);
DFFARX1 I_7990 (I601255,I2507,I138365,I138391,);
not I_7991 (I138399,I138391);
DFFARX1 I_7992 (I601240,I2507,I138365,I138425,);
not I_7993 (I138433,I601264);
or I_7994 (I138450,I601243,I601264);
nor I_7995 (I138467,I138425,I601243);
nand I_7996 (I138342,I138433,I138467);
nor I_7997 (I138498,I601246,I601243);
nand I_7998 (I138336,I138498,I138433);
not I_7999 (I138529,I601249);
nand I_8000 (I138546,I138433,I138529);
nor I_8001 (I138563,I601252,I601258);
not I_8002 (I138580,I138563);
nor I_8003 (I138597,I138580,I138546);
nor I_8004 (I138614,I138498,I138597);
DFFARX1 I_8005 (I138614,I2507,I138365,I138351,);
nor I_8006 (I138348,I138563,I138450);
DFFARX1 I_8007 (I138563,I2507,I138365,I138354,);
nor I_8008 (I138673,I138529,I601252);
nor I_8009 (I138690,I138673,I601264);
nor I_8010 (I138707,I601261,I601243);
DFFARX1 I_8011 (I138707,I2507,I138365,I138733,);
nor I_8012 (I138333,I138733,I138690);
DFFARX1 I_8013 (I138733,I2507,I138365,I138764,);
nand I_8014 (I138772,I138764,I601240);
nor I_8015 (I138357,I138399,I138772);
not I_8016 (I138803,I138733);
nand I_8017 (I138820,I138803,I601240);
nor I_8018 (I138837,I138399,I138820);
nor I_8019 (I138339,I138425,I138837);
nor I_8020 (I138868,I601261,I601246);
nor I_8021 (I138885,I138425,I138868);
DFFARX1 I_8022 (I138885,I2507,I138365,I138330,);
and I_8023 (I138345,I138498,I601261);
not I_8024 (I138960,I2514);
DFFARX1 I_8025 (I279711,I2507,I138960,I138986,);
not I_8026 (I138994,I138986);
DFFARX1 I_8027 (I279708,I2507,I138960,I139020,);
not I_8028 (I139028,I279705);
or I_8029 (I139045,I279717,I279705);
nor I_8030 (I139062,I139020,I279717);
nand I_8031 (I138937,I139028,I139062);
nor I_8032 (I139093,I279726,I279717);
nand I_8033 (I138931,I139093,I139028);
not I_8034 (I139124,I279723);
nand I_8035 (I139141,I139028,I139124);
nor I_8036 (I139158,I279702,I279702);
not I_8037 (I139175,I139158);
nor I_8038 (I139192,I139175,I139141);
nor I_8039 (I139209,I139093,I139192);
DFFARX1 I_8040 (I139209,I2507,I138960,I138946,);
nor I_8041 (I138943,I139158,I139045);
DFFARX1 I_8042 (I139158,I2507,I138960,I138949,);
nor I_8043 (I139268,I139124,I279702);
nor I_8044 (I139285,I139268,I279705);
nor I_8045 (I139302,I279714,I279729);
DFFARX1 I_8046 (I139302,I2507,I138960,I139328,);
nor I_8047 (I138928,I139328,I139285);
DFFARX1 I_8048 (I139328,I2507,I138960,I139359,);
nand I_8049 (I139367,I139359,I279720);
nor I_8050 (I138952,I138994,I139367);
not I_8051 (I139398,I139328);
nand I_8052 (I139415,I139398,I279720);
nor I_8053 (I139432,I138994,I139415);
nor I_8054 (I138934,I139020,I139432);
nor I_8055 (I139463,I279714,I279726);
nor I_8056 (I139480,I139020,I139463);
DFFARX1 I_8057 (I139480,I2507,I138960,I138925,);
and I_8058 (I138940,I139093,I279714);
not I_8059 (I139555,I2514);
DFFARX1 I_8060 (I489863,I2507,I139555,I139581,);
not I_8061 (I139589,I139581);
DFFARX1 I_8062 (I489857,I2507,I139555,I139615,);
not I_8063 (I139623,I489854);
or I_8064 (I139640,I489845,I489854);
nor I_8065 (I139657,I139615,I489845);
nand I_8066 (I139532,I139623,I139657);
nor I_8067 (I139688,I489848,I489845);
nand I_8068 (I139526,I139688,I139623);
not I_8069 (I139719,I489851);
nand I_8070 (I139736,I139623,I139719);
nor I_8071 (I139753,I489839,I489866);
not I_8072 (I139770,I139753);
nor I_8073 (I139787,I139770,I139736);
nor I_8074 (I139804,I139688,I139787);
DFFARX1 I_8075 (I139804,I2507,I139555,I139541,);
nor I_8076 (I139538,I139753,I139640);
DFFARX1 I_8077 (I139753,I2507,I139555,I139544,);
nor I_8078 (I139863,I139719,I489839);
nor I_8079 (I139880,I139863,I489854);
nor I_8080 (I139897,I489842,I489839);
DFFARX1 I_8081 (I139897,I2507,I139555,I139923,);
nor I_8082 (I139523,I139923,I139880);
DFFARX1 I_8083 (I139923,I2507,I139555,I139954,);
nand I_8084 (I139962,I139954,I489860);
nor I_8085 (I139547,I139589,I139962);
not I_8086 (I139993,I139923);
nand I_8087 (I140010,I139993,I489860);
nor I_8088 (I140027,I139589,I140010);
nor I_8089 (I139529,I139615,I140027);
nor I_8090 (I140058,I489842,I489848);
nor I_8091 (I140075,I139615,I140058);
DFFARX1 I_8092 (I140075,I2507,I139555,I139520,);
and I_8093 (I139535,I139688,I489842);
not I_8094 (I140150,I2514);
DFFARX1 I_8095 (I2260,I2507,I140150,I140176,);
not I_8096 (I140184,I140176);
DFFARX1 I_8097 (I2236,I2507,I140150,I140210,);
not I_8098 (I140218,I1820);
or I_8099 (I140235,I1980,I1820);
nor I_8100 (I140252,I140210,I1980);
nand I_8101 (I140127,I140218,I140252);
nor I_8102 (I140283,I1580,I1980);
nand I_8103 (I140121,I140283,I140218);
not I_8104 (I140314,I2268);
nand I_8105 (I140331,I140218,I140314);
nor I_8106 (I140348,I1452,I1596);
not I_8107 (I140365,I140348);
nor I_8108 (I140382,I140365,I140331);
nor I_8109 (I140399,I140283,I140382);
DFFARX1 I_8110 (I140399,I2507,I140150,I140136,);
nor I_8111 (I140133,I140348,I140235);
DFFARX1 I_8112 (I140348,I2507,I140150,I140139,);
nor I_8113 (I140458,I140314,I1452);
nor I_8114 (I140475,I140458,I1820);
nor I_8115 (I140492,I2020,I1380);
DFFARX1 I_8116 (I140492,I2507,I140150,I140518,);
nor I_8117 (I140118,I140518,I140475);
DFFARX1 I_8118 (I140518,I2507,I140150,I140549,);
nand I_8119 (I140557,I140549,I1436);
nor I_8120 (I140142,I140184,I140557);
not I_8121 (I140588,I140518);
nand I_8122 (I140605,I140588,I1436);
nor I_8123 (I140622,I140184,I140605);
nor I_8124 (I140124,I140210,I140622);
nor I_8125 (I140653,I2020,I1580);
nor I_8126 (I140670,I140210,I140653);
DFFARX1 I_8127 (I140670,I2507,I140150,I140115,);
and I_8128 (I140130,I140283,I2020);
not I_8129 (I140745,I2514);
DFFARX1 I_8130 (I102838,I2507,I140745,I140771,);
not I_8131 (I140779,I140771);
DFFARX1 I_8132 (I102832,I2507,I140745,I140805,);
not I_8133 (I140813,I102841);
or I_8134 (I140830,I102826,I102841);
nor I_8135 (I140847,I140805,I102826);
nand I_8136 (I140722,I140813,I140847);
nor I_8137 (I140878,I102817,I102826);
nand I_8138 (I140716,I140878,I140813);
not I_8139 (I140909,I102817);
nand I_8140 (I140926,I140813,I140909);
nor I_8141 (I140943,I102820,I102835);
not I_8142 (I140960,I140943);
nor I_8143 (I140977,I140960,I140926);
nor I_8144 (I140994,I140878,I140977);
DFFARX1 I_8145 (I140994,I2507,I140745,I140731,);
nor I_8146 (I140728,I140943,I140830);
DFFARX1 I_8147 (I140943,I2507,I140745,I140734,);
nor I_8148 (I141053,I140909,I102820);
nor I_8149 (I141070,I141053,I102841);
nor I_8150 (I141087,I102820,I102829);
DFFARX1 I_8151 (I141087,I2507,I140745,I141113,);
nor I_8152 (I140713,I141113,I141070);
DFFARX1 I_8153 (I141113,I2507,I140745,I141144,);
nand I_8154 (I141152,I141144,I102823);
nor I_8155 (I140737,I140779,I141152);
not I_8156 (I141183,I141113);
nand I_8157 (I141200,I141183,I102823);
nor I_8158 (I141217,I140779,I141200);
nor I_8159 (I140719,I140805,I141217);
nor I_8160 (I141248,I102820,I102817);
nor I_8161 (I141265,I140805,I141248);
DFFARX1 I_8162 (I141265,I2507,I140745,I140710,);
and I_8163 (I140725,I140878,I102820);
not I_8164 (I141340,I2514);
DFFARX1 I_8165 (I449063,I2507,I141340,I141366,);
not I_8166 (I141374,I141366);
DFFARX1 I_8167 (I449057,I2507,I141340,I141400,);
not I_8168 (I141408,I449054);
or I_8169 (I141425,I449045,I449054);
nor I_8170 (I141442,I141400,I449045);
nand I_8171 (I141317,I141408,I141442);
nor I_8172 (I141473,I449048,I449045);
nand I_8173 (I141311,I141473,I141408);
not I_8174 (I141504,I449051);
nand I_8175 (I141521,I141408,I141504);
nor I_8176 (I141538,I449039,I449066);
not I_8177 (I141555,I141538);
nor I_8178 (I141572,I141555,I141521);
nor I_8179 (I141589,I141473,I141572);
DFFARX1 I_8180 (I141589,I2507,I141340,I141326,);
nor I_8181 (I141323,I141538,I141425);
DFFARX1 I_8182 (I141538,I2507,I141340,I141329,);
nor I_8183 (I141648,I141504,I449039);
nor I_8184 (I141665,I141648,I449054);
nor I_8185 (I141682,I449042,I449039);
DFFARX1 I_8186 (I141682,I2507,I141340,I141708,);
nor I_8187 (I141308,I141708,I141665);
DFFARX1 I_8188 (I141708,I2507,I141340,I141739,);
nand I_8189 (I141747,I141739,I449060);
nor I_8190 (I141332,I141374,I141747);
not I_8191 (I141778,I141708);
nand I_8192 (I141795,I141778,I449060);
nor I_8193 (I141812,I141374,I141795);
nor I_8194 (I141314,I141400,I141812);
nor I_8195 (I141843,I449042,I449048);
nor I_8196 (I141860,I141400,I141843);
DFFARX1 I_8197 (I141860,I2507,I141340,I141305,);
and I_8198 (I141320,I141473,I449042);
not I_8199 (I141935,I2514);
DFFARX1 I_8200 (I1084383,I2507,I141935,I141961,);
not I_8201 (I141969,I141961);
DFFARX1 I_8202 (I1084380,I2507,I141935,I141995,);
not I_8203 (I142003,I1084389);
or I_8204 (I142020,I1084380,I1084389);
nor I_8205 (I142037,I141995,I1084380);
nand I_8206 (I141912,I142003,I142037);
nor I_8207 (I142068,I1084392,I1084380);
nand I_8208 (I141906,I142068,I142003);
not I_8209 (I142099,I1084386);
nand I_8210 (I142116,I142003,I142099);
nor I_8211 (I142133,I1084383,I1084401);
not I_8212 (I142150,I142133);
nor I_8213 (I142167,I142150,I142116);
nor I_8214 (I142184,I142068,I142167);
DFFARX1 I_8215 (I142184,I2507,I141935,I141921,);
nor I_8216 (I141918,I142133,I142020);
DFFARX1 I_8217 (I142133,I2507,I141935,I141924,);
nor I_8218 (I142243,I142099,I1084383);
nor I_8219 (I142260,I142243,I1084389);
nor I_8220 (I142277,I1084404,I1084398);
DFFARX1 I_8221 (I142277,I2507,I141935,I142303,);
nor I_8222 (I141903,I142303,I142260);
DFFARX1 I_8223 (I142303,I2507,I141935,I142334,);
nand I_8224 (I142342,I142334,I1084395);
nor I_8225 (I141927,I141969,I142342);
not I_8226 (I142373,I142303);
nand I_8227 (I142390,I142373,I1084395);
nor I_8228 (I142407,I141969,I142390);
nor I_8229 (I141909,I141995,I142407);
nor I_8230 (I142438,I1084404,I1084392);
nor I_8231 (I142455,I141995,I142438);
DFFARX1 I_8232 (I142455,I2507,I141935,I141900,);
and I_8233 (I141915,I142068,I1084404);
not I_8234 (I142530,I2514);
DFFARX1 I_8235 (I712216,I2507,I142530,I142556,);
not I_8236 (I142564,I142556);
DFFARX1 I_8237 (I712237,I2507,I142530,I142590,);
not I_8238 (I142598,I712216);
or I_8239 (I142615,I712228,I712216);
nor I_8240 (I142632,I142590,I712228);
nand I_8241 (I142507,I142598,I142632);
nor I_8242 (I142663,I712225,I712228);
nand I_8243 (I142501,I142663,I142598);
not I_8244 (I142694,I712234);
nand I_8245 (I142711,I142598,I142694);
nor I_8246 (I142728,I712219,I712219);
not I_8247 (I142745,I142728);
nor I_8248 (I142762,I142745,I142711);
nor I_8249 (I142779,I142663,I142762);
DFFARX1 I_8250 (I142779,I2507,I142530,I142516,);
nor I_8251 (I142513,I142728,I142615);
DFFARX1 I_8252 (I142728,I2507,I142530,I142519,);
nor I_8253 (I142838,I142694,I712219);
nor I_8254 (I142855,I142838,I712216);
nor I_8255 (I142872,I712240,I712222);
DFFARX1 I_8256 (I142872,I2507,I142530,I142898,);
nor I_8257 (I142498,I142898,I142855);
DFFARX1 I_8258 (I142898,I2507,I142530,I142929,);
nand I_8259 (I142937,I142929,I712231);
nor I_8260 (I142522,I142564,I142937);
not I_8261 (I142968,I142898);
nand I_8262 (I142985,I142968,I712231);
nor I_8263 (I143002,I142564,I142985);
nor I_8264 (I142504,I142590,I143002);
nor I_8265 (I143033,I712240,I712225);
nor I_8266 (I143050,I142590,I143033);
DFFARX1 I_8267 (I143050,I2507,I142530,I142495,);
and I_8268 (I142510,I142663,I712240);
not I_8269 (I143125,I2514);
DFFARX1 I_8270 (I697188,I2507,I143125,I143151,);
not I_8271 (I143159,I143151);
DFFARX1 I_8272 (I697209,I2507,I143125,I143185,);
not I_8273 (I143193,I697188);
or I_8274 (I143210,I697200,I697188);
nor I_8275 (I143227,I143185,I697200);
nand I_8276 (I143102,I143193,I143227);
nor I_8277 (I143258,I697197,I697200);
nand I_8278 (I143096,I143258,I143193);
not I_8279 (I143289,I697206);
nand I_8280 (I143306,I143193,I143289);
nor I_8281 (I143323,I697191,I697191);
not I_8282 (I143340,I143323);
nor I_8283 (I143357,I143340,I143306);
nor I_8284 (I143374,I143258,I143357);
DFFARX1 I_8285 (I143374,I2507,I143125,I143111,);
nor I_8286 (I143108,I143323,I143210);
DFFARX1 I_8287 (I143323,I2507,I143125,I143114,);
nor I_8288 (I143433,I143289,I697191);
nor I_8289 (I143450,I143433,I697188);
nor I_8290 (I143467,I697212,I697194);
DFFARX1 I_8291 (I143467,I2507,I143125,I143493,);
nor I_8292 (I143093,I143493,I143450);
DFFARX1 I_8293 (I143493,I2507,I143125,I143524,);
nand I_8294 (I143532,I143524,I697203);
nor I_8295 (I143117,I143159,I143532);
not I_8296 (I143563,I143493);
nand I_8297 (I143580,I143563,I697203);
nor I_8298 (I143597,I143159,I143580);
nor I_8299 (I143099,I143185,I143597);
nor I_8300 (I143628,I697212,I697197);
nor I_8301 (I143645,I143185,I143628);
DFFARX1 I_8302 (I143645,I2507,I143125,I143090,);
and I_8303 (I143105,I143258,I697212);
not I_8304 (I143720,I2514);
DFFARX1 I_8305 (I652104,I2507,I143720,I143746,);
not I_8306 (I143754,I143746);
DFFARX1 I_8307 (I652125,I2507,I143720,I143780,);
not I_8308 (I143788,I652104);
or I_8309 (I143805,I652116,I652104);
nor I_8310 (I143822,I143780,I652116);
nand I_8311 (I143697,I143788,I143822);
nor I_8312 (I143853,I652113,I652116);
nand I_8313 (I143691,I143853,I143788);
not I_8314 (I143884,I652122);
nand I_8315 (I143901,I143788,I143884);
nor I_8316 (I143918,I652107,I652107);
not I_8317 (I143935,I143918);
nor I_8318 (I143952,I143935,I143901);
nor I_8319 (I143969,I143853,I143952);
DFFARX1 I_8320 (I143969,I2507,I143720,I143706,);
nor I_8321 (I143703,I143918,I143805);
DFFARX1 I_8322 (I143918,I2507,I143720,I143709,);
nor I_8323 (I144028,I143884,I652107);
nor I_8324 (I144045,I144028,I652104);
nor I_8325 (I144062,I652128,I652110);
DFFARX1 I_8326 (I144062,I2507,I143720,I144088,);
nor I_8327 (I143688,I144088,I144045);
DFFARX1 I_8328 (I144088,I2507,I143720,I144119,);
nand I_8329 (I144127,I144119,I652119);
nor I_8330 (I143712,I143754,I144127);
not I_8331 (I144158,I144088);
nand I_8332 (I144175,I144158,I652119);
nor I_8333 (I144192,I143754,I144175);
nor I_8334 (I143694,I143780,I144192);
nor I_8335 (I144223,I652128,I652113);
nor I_8336 (I144240,I143780,I144223);
DFFARX1 I_8337 (I144240,I2507,I143720,I143685,);
and I_8338 (I143700,I143853,I652128);
not I_8339 (I144315,I2514);
DFFARX1 I_8340 (I604723,I2507,I144315,I144341,);
not I_8341 (I144349,I144341);
DFFARX1 I_8342 (I604708,I2507,I144315,I144375,);
not I_8343 (I144383,I604732);
or I_8344 (I144400,I604711,I604732);
nor I_8345 (I144417,I144375,I604711);
nand I_8346 (I144292,I144383,I144417);
nor I_8347 (I144448,I604714,I604711);
nand I_8348 (I144286,I144448,I144383);
not I_8349 (I144479,I604717);
nand I_8350 (I144496,I144383,I144479);
nor I_8351 (I144513,I604720,I604726);
not I_8352 (I144530,I144513);
nor I_8353 (I144547,I144530,I144496);
nor I_8354 (I144564,I144448,I144547);
DFFARX1 I_8355 (I144564,I2507,I144315,I144301,);
nor I_8356 (I144298,I144513,I144400);
DFFARX1 I_8357 (I144513,I2507,I144315,I144304,);
nor I_8358 (I144623,I144479,I604720);
nor I_8359 (I144640,I144623,I604732);
nor I_8360 (I144657,I604729,I604711);
DFFARX1 I_8361 (I144657,I2507,I144315,I144683,);
nor I_8362 (I144283,I144683,I144640);
DFFARX1 I_8363 (I144683,I2507,I144315,I144714,);
nand I_8364 (I144722,I144714,I604708);
nor I_8365 (I144307,I144349,I144722);
not I_8366 (I144753,I144683);
nand I_8367 (I144770,I144753,I604708);
nor I_8368 (I144787,I144349,I144770);
nor I_8369 (I144289,I144375,I144787);
nor I_8370 (I144818,I604729,I604714);
nor I_8371 (I144835,I144375,I144818);
DFFARX1 I_8372 (I144835,I2507,I144315,I144280,);
and I_8373 (I144295,I144448,I604729);
not I_8374 (I144910,I2514);
DFFARX1 I_8375 (I567731,I2507,I144910,I144936,);
not I_8376 (I144944,I144936);
DFFARX1 I_8377 (I567716,I2507,I144910,I144970,);
not I_8378 (I144978,I567740);
or I_8379 (I144995,I567719,I567740);
nor I_8380 (I145012,I144970,I567719);
nand I_8381 (I144887,I144978,I145012);
nor I_8382 (I145043,I567722,I567719);
nand I_8383 (I144881,I145043,I144978);
not I_8384 (I145074,I567725);
nand I_8385 (I145091,I144978,I145074);
nor I_8386 (I145108,I567728,I567734);
not I_8387 (I145125,I145108);
nor I_8388 (I145142,I145125,I145091);
nor I_8389 (I145159,I145043,I145142);
DFFARX1 I_8390 (I145159,I2507,I144910,I144896,);
nor I_8391 (I144893,I145108,I144995);
DFFARX1 I_8392 (I145108,I2507,I144910,I144899,);
nor I_8393 (I145218,I145074,I567728);
nor I_8394 (I145235,I145218,I567740);
nor I_8395 (I145252,I567737,I567719);
DFFARX1 I_8396 (I145252,I2507,I144910,I145278,);
nor I_8397 (I144878,I145278,I145235);
DFFARX1 I_8398 (I145278,I2507,I144910,I145309,);
nand I_8399 (I145317,I145309,I567716);
nor I_8400 (I144902,I144944,I145317);
not I_8401 (I145348,I145278);
nand I_8402 (I145365,I145348,I567716);
nor I_8403 (I145382,I144944,I145365);
nor I_8404 (I144884,I144970,I145382);
nor I_8405 (I145413,I567737,I567722);
nor I_8406 (I145430,I144970,I145413);
DFFARX1 I_8407 (I145430,I2507,I144910,I144875,);
and I_8408 (I144890,I145043,I567737);
not I_8409 (I145505,I2514);
DFFARX1 I_8410 (I231769,I2507,I145505,I145531,);
not I_8411 (I145539,I145531);
DFFARX1 I_8412 (I231763,I2507,I145505,I145565,);
not I_8413 (I145573,I231748);
or I_8414 (I145590,I231757,I231748);
nor I_8415 (I145607,I145565,I231757);
nand I_8416 (I145482,I145573,I145607);
nor I_8417 (I145638,I231745,I231757);
nand I_8418 (I145476,I145638,I145573);
not I_8419 (I145669,I231751);
nand I_8420 (I145686,I145573,I145669);
nor I_8421 (I145703,I231754,I231766);
not I_8422 (I145720,I145703);
nor I_8423 (I145737,I145720,I145686);
nor I_8424 (I145754,I145638,I145737);
DFFARX1 I_8425 (I145754,I2507,I145505,I145491,);
nor I_8426 (I145488,I145703,I145590);
DFFARX1 I_8427 (I145703,I2507,I145505,I145494,);
nor I_8428 (I145813,I145669,I231754);
nor I_8429 (I145830,I145813,I231748);
nor I_8430 (I145847,I231760,I231748);
DFFARX1 I_8431 (I145847,I2507,I145505,I145873,);
nor I_8432 (I145473,I145873,I145830);
DFFARX1 I_8433 (I145873,I2507,I145505,I145904,);
nand I_8434 (I145912,I145904,I231745);
nor I_8435 (I145497,I145539,I145912);
not I_8436 (I145943,I145873);
nand I_8437 (I145960,I145943,I231745);
nor I_8438 (I145977,I145539,I145960);
nor I_8439 (I145479,I145565,I145977);
nor I_8440 (I146008,I231760,I231745);
nor I_8441 (I146025,I145565,I146008);
DFFARX1 I_8442 (I146025,I2507,I145505,I145470,);
and I_8443 (I145485,I145638,I231760);
not I_8444 (I146100,I2514);
DFFARX1 I_8445 (I498266,I2507,I146100,I146126,);
not I_8446 (I146134,I146126);
DFFARX1 I_8447 (I498272,I2507,I146100,I146160,);
not I_8448 (I146168,I498254);
or I_8449 (I146185,I498278,I498254);
nor I_8450 (I146202,I146160,I498278);
nand I_8451 (I146077,I146168,I146202);
nor I_8452 (I146233,I498269,I498278);
nand I_8453 (I146071,I146233,I146168);
not I_8454 (I146264,I498260);
nand I_8455 (I146281,I146168,I146264);
nor I_8456 (I146298,I498263,I498257);
not I_8457 (I146315,I146298);
nor I_8458 (I146332,I146315,I146281);
nor I_8459 (I146349,I146233,I146332);
DFFARX1 I_8460 (I146349,I2507,I146100,I146086,);
nor I_8461 (I146083,I146298,I146185);
DFFARX1 I_8462 (I146298,I2507,I146100,I146089,);
nor I_8463 (I146408,I146264,I498263);
nor I_8464 (I146425,I146408,I498254);
nor I_8465 (I146442,I498275,I498254);
DFFARX1 I_8466 (I146442,I2507,I146100,I146468,);
nor I_8467 (I146068,I146468,I146425);
DFFARX1 I_8468 (I146468,I2507,I146100,I146499,);
nand I_8469 (I146507,I146499,I498257);
nor I_8470 (I146092,I146134,I146507);
not I_8471 (I146538,I146468);
nand I_8472 (I146555,I146538,I498257);
nor I_8473 (I146572,I146134,I146555);
nor I_8474 (I146074,I146160,I146572);
nor I_8475 (I146603,I498275,I498269);
nor I_8476 (I146620,I146160,I146603);
DFFARX1 I_8477 (I146620,I2507,I146100,I146065,);
and I_8478 (I146080,I146233,I498275);
not I_8479 (I146695,I2514);
DFFARX1 I_8480 (I850738,I2507,I146695,I146721,);
not I_8481 (I146729,I146721);
DFFARX1 I_8482 (I850738,I2507,I146695,I146755,);
not I_8483 (I146763,I850735);
or I_8484 (I146780,I850747,I850735);
nor I_8485 (I146797,I146755,I850747);
nand I_8486 (I146672,I146763,I146797);
nor I_8487 (I146828,I850741,I850747);
nand I_8488 (I146666,I146828,I146763);
not I_8489 (I146859,I850753);
nand I_8490 (I146876,I146763,I146859);
nor I_8491 (I146893,I850744,I850732);
not I_8492 (I146910,I146893);
nor I_8493 (I146927,I146910,I146876);
nor I_8494 (I146944,I146828,I146927);
DFFARX1 I_8495 (I146944,I2507,I146695,I146681,);
nor I_8496 (I146678,I146893,I146780);
DFFARX1 I_8497 (I146893,I2507,I146695,I146684,);
nor I_8498 (I147003,I146859,I850744);
nor I_8499 (I147020,I147003,I850735);
nor I_8500 (I147037,I850735,I850732);
DFFARX1 I_8501 (I147037,I2507,I146695,I147063,);
nor I_8502 (I146663,I147063,I147020);
DFFARX1 I_8503 (I147063,I2507,I146695,I147094,);
nand I_8504 (I147102,I147094,I850750);
nor I_8505 (I146687,I146729,I147102);
not I_8506 (I147133,I147063);
nand I_8507 (I147150,I147133,I850750);
nor I_8508 (I147167,I146729,I147150);
nor I_8509 (I146669,I146755,I147167);
nor I_8510 (I147198,I850735,I850741);
nor I_8511 (I147215,I146755,I147198);
DFFARX1 I_8512 (I147215,I2507,I146695,I146660,);
and I_8513 (I146675,I146828,I850735);
not I_8514 (I147290,I2514);
DFFARX1 I_8515 (I225224,I2507,I147290,I147316,);
not I_8516 (I147324,I147316);
DFFARX1 I_8517 (I225218,I2507,I147290,I147350,);
not I_8518 (I147358,I225203);
or I_8519 (I147375,I225212,I225203);
nor I_8520 (I147392,I147350,I225212);
nand I_8521 (I147267,I147358,I147392);
nor I_8522 (I147423,I225200,I225212);
nand I_8523 (I147261,I147423,I147358);
not I_8524 (I147454,I225206);
nand I_8525 (I147471,I147358,I147454);
nor I_8526 (I147488,I225209,I225221);
not I_8527 (I147505,I147488);
nor I_8528 (I147522,I147505,I147471);
nor I_8529 (I147539,I147423,I147522);
DFFARX1 I_8530 (I147539,I2507,I147290,I147276,);
nor I_8531 (I147273,I147488,I147375);
DFFARX1 I_8532 (I147488,I2507,I147290,I147279,);
nor I_8533 (I147598,I147454,I225209);
nor I_8534 (I147615,I147598,I225203);
nor I_8535 (I147632,I225215,I225203);
DFFARX1 I_8536 (I147632,I2507,I147290,I147658,);
nor I_8537 (I147258,I147658,I147615);
DFFARX1 I_8538 (I147658,I2507,I147290,I147689,);
nand I_8539 (I147697,I147689,I225200);
nor I_8540 (I147282,I147324,I147697);
not I_8541 (I147728,I147658);
nand I_8542 (I147745,I147728,I225200);
nor I_8543 (I147762,I147324,I147745);
nor I_8544 (I147264,I147350,I147762);
nor I_8545 (I147793,I225215,I225200);
nor I_8546 (I147810,I147350,I147793);
DFFARX1 I_8547 (I147810,I2507,I147290,I147255,);
and I_8548 (I147270,I147423,I225215);
not I_8549 (I147885,I2514);
DFFARX1 I_8550 (I105473,I2507,I147885,I147911,);
not I_8551 (I147919,I147911);
DFFARX1 I_8552 (I105467,I2507,I147885,I147945,);
not I_8553 (I147953,I105476);
or I_8554 (I147970,I105461,I105476);
nor I_8555 (I147987,I147945,I105461);
nand I_8556 (I147862,I147953,I147987);
nor I_8557 (I148018,I105452,I105461);
nand I_8558 (I147856,I148018,I147953);
not I_8559 (I148049,I105452);
nand I_8560 (I148066,I147953,I148049);
nor I_8561 (I148083,I105455,I105470);
not I_8562 (I148100,I148083);
nor I_8563 (I148117,I148100,I148066);
nor I_8564 (I148134,I148018,I148117);
DFFARX1 I_8565 (I148134,I2507,I147885,I147871,);
nor I_8566 (I147868,I148083,I147970);
DFFARX1 I_8567 (I148083,I2507,I147885,I147874,);
nor I_8568 (I148193,I148049,I105455);
nor I_8569 (I148210,I148193,I105476);
nor I_8570 (I148227,I105455,I105464);
DFFARX1 I_8571 (I148227,I2507,I147885,I148253,);
nor I_8572 (I147853,I148253,I148210);
DFFARX1 I_8573 (I148253,I2507,I147885,I148284,);
nand I_8574 (I148292,I148284,I105458);
nor I_8575 (I147877,I147919,I148292);
not I_8576 (I148323,I148253);
nand I_8577 (I148340,I148323,I105458);
nor I_8578 (I148357,I147919,I148340);
nor I_8579 (I147859,I147945,I148357);
nor I_8580 (I148388,I105455,I105452);
nor I_8581 (I148405,I147945,I148388);
DFFARX1 I_8582 (I148405,I2507,I147885,I147850,);
and I_8583 (I147865,I148018,I105455);
not I_8584 (I148477,I2514);
DFFARX1 I_8585 (I621485,I2507,I148477,I148503,);
DFFARX1 I_8586 (I148503,I2507,I148477,I148520,);
not I_8587 (I148469,I148520);
not I_8588 (I148542,I148503);
DFFARX1 I_8589 (I621476,I2507,I148477,I148568,);
not I_8590 (I148576,I148568);
and I_8591 (I148593,I148542,I621494);
not I_8592 (I148610,I621491);
nand I_8593 (I148627,I148610,I621494);
not I_8594 (I148644,I621470);
nor I_8595 (I148661,I148644,I621473);
nand I_8596 (I148678,I148661,I621482);
nor I_8597 (I148695,I148678,I148627);
DFFARX1 I_8598 (I148695,I2507,I148477,I148445,);
not I_8599 (I148726,I148678);
not I_8600 (I148743,I621473);
nand I_8601 (I148760,I148743,I621494);
nor I_8602 (I148777,I621473,I621491);
nand I_8603 (I148457,I148593,I148777);
nand I_8604 (I148451,I148542,I621473);
nand I_8605 (I148822,I148644,I621488);
DFFARX1 I_8606 (I148822,I2507,I148477,I148466,);
DFFARX1 I_8607 (I148822,I2507,I148477,I148460,);
not I_8608 (I148867,I621488);
nor I_8609 (I148884,I148867,I621470);
and I_8610 (I148901,I148884,I621479);
or I_8611 (I148918,I148901,I621473);
DFFARX1 I_8612 (I148918,I2507,I148477,I148944,);
nand I_8613 (I148952,I148944,I148610);
nor I_8614 (I148454,I148952,I148760);
nor I_8615 (I148448,I148944,I148576);
DFFARX1 I_8616 (I148944,I2507,I148477,I149006,);
not I_8617 (I149014,I149006);
nor I_8618 (I148463,I149014,I148726);
not I_8619 (I149072,I2514);
DFFARX1 I_8620 (I490951,I2507,I149072,I149098,);
DFFARX1 I_8621 (I149098,I2507,I149072,I149115,);
not I_8622 (I149064,I149115);
not I_8623 (I149137,I149098);
DFFARX1 I_8624 (I490939,I2507,I149072,I149163,);
not I_8625 (I149171,I149163);
and I_8626 (I149188,I149137,I490948);
not I_8627 (I149205,I490945);
nand I_8628 (I149222,I149205,I490948);
not I_8629 (I149239,I490936);
nor I_8630 (I149256,I149239,I490942);
nand I_8631 (I149273,I149256,I490927);
nor I_8632 (I149290,I149273,I149222);
DFFARX1 I_8633 (I149290,I2507,I149072,I149040,);
not I_8634 (I149321,I149273);
not I_8635 (I149338,I490942);
nand I_8636 (I149355,I149338,I490948);
nor I_8637 (I149372,I490942,I490945);
nand I_8638 (I149052,I149188,I149372);
nand I_8639 (I149046,I149137,I490942);
nand I_8640 (I149417,I149239,I490927);
DFFARX1 I_8641 (I149417,I2507,I149072,I149061,);
DFFARX1 I_8642 (I149417,I2507,I149072,I149055,);
not I_8643 (I149462,I490927);
nor I_8644 (I149479,I149462,I490933);
and I_8645 (I149496,I149479,I490930);
or I_8646 (I149513,I149496,I490954);
DFFARX1 I_8647 (I149513,I2507,I149072,I149539,);
nand I_8648 (I149547,I149539,I149205);
nor I_8649 (I149049,I149547,I149355);
nor I_8650 (I149043,I149539,I149171);
DFFARX1 I_8651 (I149539,I2507,I149072,I149601,);
not I_8652 (I149609,I149601);
nor I_8653 (I149058,I149609,I149321);
not I_8654 (I149667,I2514);
DFFARX1 I_8655 (I1134666,I2507,I149667,I149693,);
DFFARX1 I_8656 (I149693,I2507,I149667,I149710,);
not I_8657 (I149659,I149710);
not I_8658 (I149732,I149693);
DFFARX1 I_8659 (I1134666,I2507,I149667,I149758,);
not I_8660 (I149766,I149758);
and I_8661 (I149783,I149732,I1134669);
not I_8662 (I149800,I1134681);
nand I_8663 (I149817,I149800,I1134669);
not I_8664 (I149834,I1134687);
nor I_8665 (I149851,I149834,I1134678);
nand I_8666 (I149868,I149851,I1134684);
nor I_8667 (I149885,I149868,I149817);
DFFARX1 I_8668 (I149885,I2507,I149667,I149635,);
not I_8669 (I149916,I149868);
not I_8670 (I149933,I1134678);
nand I_8671 (I149950,I149933,I1134669);
nor I_8672 (I149967,I1134678,I1134681);
nand I_8673 (I149647,I149783,I149967);
nand I_8674 (I149641,I149732,I1134678);
nand I_8675 (I150012,I149834,I1134675);
DFFARX1 I_8676 (I150012,I2507,I149667,I149656,);
DFFARX1 I_8677 (I150012,I2507,I149667,I149650,);
not I_8678 (I150057,I1134675);
nor I_8679 (I150074,I150057,I1134672);
and I_8680 (I150091,I150074,I1134690);
or I_8681 (I150108,I150091,I1134669);
DFFARX1 I_8682 (I150108,I2507,I149667,I150134,);
nand I_8683 (I150142,I150134,I149800);
nor I_8684 (I149644,I150142,I149950);
nor I_8685 (I149638,I150134,I149766);
DFFARX1 I_8686 (I150134,I2507,I149667,I150196,);
not I_8687 (I150204,I150196);
nor I_8688 (I149653,I150204,I149916);
not I_8689 (I150262,I2514);
DFFARX1 I_8690 (I510166,I2507,I150262,I150288,);
DFFARX1 I_8691 (I150288,I2507,I150262,I150305,);
not I_8692 (I150254,I150305);
not I_8693 (I150327,I150288);
DFFARX1 I_8694 (I510160,I2507,I150262,I150353,);
not I_8695 (I150361,I150353);
and I_8696 (I150378,I150327,I510175);
not I_8697 (I150395,I510172);
nand I_8698 (I150412,I150395,I510175);
not I_8699 (I150429,I510163);
nor I_8700 (I150446,I150429,I510154);
nand I_8701 (I150463,I150446,I510157);
nor I_8702 (I150480,I150463,I150412);
DFFARX1 I_8703 (I150480,I2507,I150262,I150230,);
not I_8704 (I150511,I150463);
not I_8705 (I150528,I510154);
nand I_8706 (I150545,I150528,I510175);
nor I_8707 (I150562,I510154,I510172);
nand I_8708 (I150242,I150378,I150562);
nand I_8709 (I150236,I150327,I510154);
nand I_8710 (I150607,I150429,I510178);
DFFARX1 I_8711 (I150607,I2507,I150262,I150251,);
DFFARX1 I_8712 (I150607,I2507,I150262,I150245,);
not I_8713 (I150652,I510178);
nor I_8714 (I150669,I150652,I510169);
and I_8715 (I150686,I150669,I510154);
or I_8716 (I150703,I150686,I510157);
DFFARX1 I_8717 (I150703,I2507,I150262,I150729,);
nand I_8718 (I150737,I150729,I150395);
nor I_8719 (I150239,I150737,I150545);
nor I_8720 (I150233,I150729,I150361);
DFFARX1 I_8721 (I150729,I2507,I150262,I150791,);
not I_8722 (I150799,I150791);
nor I_8723 (I150248,I150799,I150511);
not I_8724 (I150857,I2514);
DFFARX1 I_8725 (I335564,I2507,I150857,I150883,);
DFFARX1 I_8726 (I150883,I2507,I150857,I150900,);
not I_8727 (I150849,I150900);
not I_8728 (I150922,I150883);
DFFARX1 I_8729 (I335579,I2507,I150857,I150948,);
not I_8730 (I150956,I150948);
and I_8731 (I150973,I150922,I335576);
not I_8732 (I150990,I335564);
nand I_8733 (I151007,I150990,I335576);
not I_8734 (I151024,I335573);
nor I_8735 (I151041,I151024,I335588);
nand I_8736 (I151058,I151041,I335585);
nor I_8737 (I151075,I151058,I151007);
DFFARX1 I_8738 (I151075,I2507,I150857,I150825,);
not I_8739 (I151106,I151058);
not I_8740 (I151123,I335588);
nand I_8741 (I151140,I151123,I335576);
nor I_8742 (I151157,I335588,I335564);
nand I_8743 (I150837,I150973,I151157);
nand I_8744 (I150831,I150922,I335588);
nand I_8745 (I151202,I151024,I335582);
DFFARX1 I_8746 (I151202,I2507,I150857,I150846,);
DFFARX1 I_8747 (I151202,I2507,I150857,I150840,);
not I_8748 (I151247,I335582);
nor I_8749 (I151264,I151247,I335570);
and I_8750 (I151281,I151264,I335591);
or I_8751 (I151298,I151281,I335567);
DFFARX1 I_8752 (I151298,I2507,I150857,I151324,);
nand I_8753 (I151332,I151324,I150990);
nor I_8754 (I150834,I151332,I151140);
nor I_8755 (I150828,I151324,I150956);
DFFARX1 I_8756 (I151324,I2507,I150857,I151386,);
not I_8757 (I151394,I151386);
nor I_8758 (I150843,I151394,I151106);
not I_8759 (I151452,I2514);
DFFARX1 I_8760 (I786444,I2507,I151452,I151478,);
DFFARX1 I_8761 (I151478,I2507,I151452,I151495,);
not I_8762 (I151444,I151495);
not I_8763 (I151517,I151478);
DFFARX1 I_8764 (I786438,I2507,I151452,I151543,);
not I_8765 (I151551,I151543);
and I_8766 (I151568,I151517,I786456);
not I_8767 (I151585,I786444);
nand I_8768 (I151602,I151585,I786456);
not I_8769 (I151619,I786438);
nor I_8770 (I151636,I151619,I786450);
nand I_8771 (I151653,I151636,I786441);
nor I_8772 (I151670,I151653,I151602);
DFFARX1 I_8773 (I151670,I2507,I151452,I151420,);
not I_8774 (I151701,I151653);
not I_8775 (I151718,I786450);
nand I_8776 (I151735,I151718,I786456);
nor I_8777 (I151752,I786450,I786444);
nand I_8778 (I151432,I151568,I151752);
nand I_8779 (I151426,I151517,I786450);
nand I_8780 (I151797,I151619,I786453);
DFFARX1 I_8781 (I151797,I2507,I151452,I151441,);
DFFARX1 I_8782 (I151797,I2507,I151452,I151435,);
not I_8783 (I151842,I786453);
nor I_8784 (I151859,I151842,I786459);
and I_8785 (I151876,I151859,I786441);
or I_8786 (I151893,I151876,I786447);
DFFARX1 I_8787 (I151893,I2507,I151452,I151919,);
nand I_8788 (I151927,I151919,I151585);
nor I_8789 (I151429,I151927,I151735);
nor I_8790 (I151423,I151919,I151551);
DFFARX1 I_8791 (I151919,I2507,I151452,I151981,);
not I_8792 (I151989,I151981);
nor I_8793 (I151438,I151989,I151701);
not I_8794 (I152047,I2514);
DFFARX1 I_8795 (I890170,I2507,I152047,I152073,);
DFFARX1 I_8796 (I152073,I2507,I152047,I152090,);
not I_8797 (I152039,I152090);
not I_8798 (I152112,I152073);
DFFARX1 I_8799 (I890179,I2507,I152047,I152138,);
not I_8800 (I152146,I152138);
and I_8801 (I152163,I152112,I890167);
not I_8802 (I152180,I890158);
nand I_8803 (I152197,I152180,I890167);
not I_8804 (I152214,I890164);
nor I_8805 (I152231,I152214,I890182);
nand I_8806 (I152248,I152231,I890155);
nor I_8807 (I152265,I152248,I152197);
DFFARX1 I_8808 (I152265,I2507,I152047,I152015,);
not I_8809 (I152296,I152248);
not I_8810 (I152313,I890182);
nand I_8811 (I152330,I152313,I890167);
nor I_8812 (I152347,I890182,I890158);
nand I_8813 (I152027,I152163,I152347);
nand I_8814 (I152021,I152112,I890182);
nand I_8815 (I152392,I152214,I890161);
DFFARX1 I_8816 (I152392,I2507,I152047,I152036,);
DFFARX1 I_8817 (I152392,I2507,I152047,I152030,);
not I_8818 (I152437,I890161);
nor I_8819 (I152454,I152437,I890173);
and I_8820 (I152471,I152454,I890155);
or I_8821 (I152488,I152471,I890176);
DFFARX1 I_8822 (I152488,I2507,I152047,I152514,);
nand I_8823 (I152522,I152514,I152180);
nor I_8824 (I152024,I152522,I152330);
nor I_8825 (I152018,I152514,I152146);
DFFARX1 I_8826 (I152514,I2507,I152047,I152576,);
not I_8827 (I152584,I152576);
nor I_8828 (I152033,I152584,I152296);
not I_8829 (I152642,I2514);
DFFARX1 I_8830 (I1376733,I2507,I152642,I152668,);
DFFARX1 I_8831 (I152668,I2507,I152642,I152685,);
not I_8832 (I152634,I152685);
not I_8833 (I152707,I152668);
DFFARX1 I_8834 (I1376724,I2507,I152642,I152733,);
not I_8835 (I152741,I152733);
and I_8836 (I152758,I152707,I1376718);
not I_8837 (I152775,I1376712);
nand I_8838 (I152792,I152775,I1376718);
not I_8839 (I152809,I1376739);
nor I_8840 (I152826,I152809,I1376712);
nand I_8841 (I152843,I152826,I1376736);
nor I_8842 (I152860,I152843,I152792);
DFFARX1 I_8843 (I152860,I2507,I152642,I152610,);
not I_8844 (I152891,I152843);
not I_8845 (I152908,I1376712);
nand I_8846 (I152925,I152908,I1376718);
nor I_8847 (I152942,I1376712,I1376712);
nand I_8848 (I152622,I152758,I152942);
nand I_8849 (I152616,I152707,I1376712);
nand I_8850 (I152987,I152809,I1376721);
DFFARX1 I_8851 (I152987,I2507,I152642,I152631,);
DFFARX1 I_8852 (I152987,I2507,I152642,I152625,);
not I_8853 (I153032,I1376721);
nor I_8854 (I153049,I153032,I1376727);
and I_8855 (I153066,I153049,I1376730);
or I_8856 (I153083,I153066,I1376715);
DFFARX1 I_8857 (I153083,I2507,I152642,I153109,);
nand I_8858 (I153117,I153109,I152775);
nor I_8859 (I152619,I153117,I152925);
nor I_8860 (I152613,I153109,I152741);
DFFARX1 I_8861 (I153109,I2507,I152642,I153171,);
not I_8862 (I153179,I153171);
nor I_8863 (I152628,I153179,I152891);
not I_8864 (I153237,I2514);
DFFARX1 I_8865 (I323443,I2507,I153237,I153263,);
DFFARX1 I_8866 (I153263,I2507,I153237,I153280,);
not I_8867 (I153229,I153280);
not I_8868 (I153302,I153263);
DFFARX1 I_8869 (I323458,I2507,I153237,I153328,);
not I_8870 (I153336,I153328);
and I_8871 (I153353,I153302,I323455);
not I_8872 (I153370,I323443);
nand I_8873 (I153387,I153370,I323455);
not I_8874 (I153404,I323452);
nor I_8875 (I153421,I153404,I323467);
nand I_8876 (I153438,I153421,I323464);
nor I_8877 (I153455,I153438,I153387);
DFFARX1 I_8878 (I153455,I2507,I153237,I153205,);
not I_8879 (I153486,I153438);
not I_8880 (I153503,I323467);
nand I_8881 (I153520,I153503,I323455);
nor I_8882 (I153537,I323467,I323443);
nand I_8883 (I153217,I153353,I153537);
nand I_8884 (I153211,I153302,I323467);
nand I_8885 (I153582,I153404,I323461);
DFFARX1 I_8886 (I153582,I2507,I153237,I153226,);
DFFARX1 I_8887 (I153582,I2507,I153237,I153220,);
not I_8888 (I153627,I323461);
nor I_8889 (I153644,I153627,I323449);
and I_8890 (I153661,I153644,I323470);
or I_8891 (I153678,I153661,I323446);
DFFARX1 I_8892 (I153678,I2507,I153237,I153704,);
nand I_8893 (I153712,I153704,I153370);
nor I_8894 (I153214,I153712,I153520);
nor I_8895 (I153208,I153704,I153336);
DFFARX1 I_8896 (I153704,I2507,I153237,I153766,);
not I_8897 (I153774,I153766);
nor I_8898 (I153223,I153774,I153486);
not I_8899 (I153832,I2514);
DFFARX1 I_8900 (I935390,I2507,I153832,I153858,);
DFFARX1 I_8901 (I153858,I2507,I153832,I153875,);
not I_8902 (I153824,I153875);
not I_8903 (I153897,I153858);
DFFARX1 I_8904 (I935399,I2507,I153832,I153923,);
not I_8905 (I153931,I153923);
and I_8906 (I153948,I153897,I935387);
not I_8907 (I153965,I935378);
nand I_8908 (I153982,I153965,I935387);
not I_8909 (I153999,I935384);
nor I_8910 (I154016,I153999,I935402);
nand I_8911 (I154033,I154016,I935375);
nor I_8912 (I154050,I154033,I153982);
DFFARX1 I_8913 (I154050,I2507,I153832,I153800,);
not I_8914 (I154081,I154033);
not I_8915 (I154098,I935402);
nand I_8916 (I154115,I154098,I935387);
nor I_8917 (I154132,I935402,I935378);
nand I_8918 (I153812,I153948,I154132);
nand I_8919 (I153806,I153897,I935402);
nand I_8920 (I154177,I153999,I935381);
DFFARX1 I_8921 (I154177,I2507,I153832,I153821,);
DFFARX1 I_8922 (I154177,I2507,I153832,I153815,);
not I_8923 (I154222,I935381);
nor I_8924 (I154239,I154222,I935393);
and I_8925 (I154256,I154239,I935375);
or I_8926 (I154273,I154256,I935396);
DFFARX1 I_8927 (I154273,I2507,I153832,I154299,);
nand I_8928 (I154307,I154299,I153965);
nor I_8929 (I153809,I154307,I154115);
nor I_8930 (I153803,I154299,I153931);
DFFARX1 I_8931 (I154299,I2507,I153832,I154361,);
not I_8932 (I154369,I154361);
nor I_8933 (I153818,I154369,I154081);
not I_8934 (I154427,I2514);
DFFARX1 I_8935 (I1080334,I2507,I154427,I154453,);
DFFARX1 I_8936 (I154453,I2507,I154427,I154470,);
not I_8937 (I154419,I154470);
not I_8938 (I154492,I154453);
DFFARX1 I_8939 (I1080334,I2507,I154427,I154518,);
not I_8940 (I154526,I154518);
and I_8941 (I154543,I154492,I1080337);
not I_8942 (I154560,I1080349);
nand I_8943 (I154577,I154560,I1080337);
not I_8944 (I154594,I1080355);
nor I_8945 (I154611,I154594,I1080346);
nand I_8946 (I154628,I154611,I1080352);
nor I_8947 (I154645,I154628,I154577);
DFFARX1 I_8948 (I154645,I2507,I154427,I154395,);
not I_8949 (I154676,I154628);
not I_8950 (I154693,I1080346);
nand I_8951 (I154710,I154693,I1080337);
nor I_8952 (I154727,I1080346,I1080349);
nand I_8953 (I154407,I154543,I154727);
nand I_8954 (I154401,I154492,I1080346);
nand I_8955 (I154772,I154594,I1080343);
DFFARX1 I_8956 (I154772,I2507,I154427,I154416,);
DFFARX1 I_8957 (I154772,I2507,I154427,I154410,);
not I_8958 (I154817,I1080343);
nor I_8959 (I154834,I154817,I1080340);
and I_8960 (I154851,I154834,I1080358);
or I_8961 (I154868,I154851,I1080337);
DFFARX1 I_8962 (I154868,I2507,I154427,I154894,);
nand I_8963 (I154902,I154894,I154560);
nor I_8964 (I154404,I154902,I154710);
nor I_8965 (I154398,I154894,I154526);
DFFARX1 I_8966 (I154894,I2507,I154427,I154956,);
not I_8967 (I154964,I154956);
nor I_8968 (I154413,I154964,I154676);
not I_8969 (I155022,I2514);
DFFARX1 I_8970 (I1916,I2507,I155022,I155048,);
DFFARX1 I_8971 (I155048,I2507,I155022,I155065,);
not I_8972 (I155014,I155065);
not I_8973 (I155087,I155048);
DFFARX1 I_8974 (I1732,I2507,I155022,I155113,);
not I_8975 (I155121,I155113);
and I_8976 (I155138,I155087,I2252);
not I_8977 (I155155,I1892);
nand I_8978 (I155172,I155155,I2252);
not I_8979 (I155189,I1524);
nor I_8980 (I155206,I155189,I1668);
nand I_8981 (I155223,I155206,I1588);
nor I_8982 (I155240,I155223,I155172);
DFFARX1 I_8983 (I155240,I2507,I155022,I154990,);
not I_8984 (I155271,I155223);
not I_8985 (I155288,I1668);
nand I_8986 (I155305,I155288,I2252);
nor I_8987 (I155322,I1668,I1892);
nand I_8988 (I155002,I155138,I155322);
nand I_8989 (I154996,I155087,I1668);
nand I_8990 (I155367,I155189,I2204);
DFFARX1 I_8991 (I155367,I2507,I155022,I155011,);
DFFARX1 I_8992 (I155367,I2507,I155022,I155005,);
not I_8993 (I155412,I2204);
nor I_8994 (I155429,I155412,I1932);
and I_8995 (I155446,I155429,I2468);
or I_8996 (I155463,I155446,I1844);
DFFARX1 I_8997 (I155463,I2507,I155022,I155489,);
nand I_8998 (I155497,I155489,I155155);
nor I_8999 (I154999,I155497,I155305);
nor I_9000 (I154993,I155489,I155121);
DFFARX1 I_9001 (I155489,I2507,I155022,I155551,);
not I_9002 (I155559,I155551);
nor I_9003 (I155008,I155559,I155271);
not I_9004 (I155617,I2514);
DFFARX1 I_9005 (I1071086,I2507,I155617,I155643,);
DFFARX1 I_9006 (I155643,I2507,I155617,I155660,);
not I_9007 (I155609,I155660);
not I_9008 (I155682,I155643);
DFFARX1 I_9009 (I1071086,I2507,I155617,I155708,);
not I_9010 (I155716,I155708);
and I_9011 (I155733,I155682,I1071089);
not I_9012 (I155750,I1071101);
nand I_9013 (I155767,I155750,I1071089);
not I_9014 (I155784,I1071107);
nor I_9015 (I155801,I155784,I1071098);
nand I_9016 (I155818,I155801,I1071104);
nor I_9017 (I155835,I155818,I155767);
DFFARX1 I_9018 (I155835,I2507,I155617,I155585,);
not I_9019 (I155866,I155818);
not I_9020 (I155883,I1071098);
nand I_9021 (I155900,I155883,I1071089);
nor I_9022 (I155917,I1071098,I1071101);
nand I_9023 (I155597,I155733,I155917);
nand I_9024 (I155591,I155682,I1071098);
nand I_9025 (I155962,I155784,I1071095);
DFFARX1 I_9026 (I155962,I2507,I155617,I155606,);
DFFARX1 I_9027 (I155962,I2507,I155617,I155600,);
not I_9028 (I156007,I1071095);
nor I_9029 (I156024,I156007,I1071092);
and I_9030 (I156041,I156024,I1071110);
or I_9031 (I156058,I156041,I1071089);
DFFARX1 I_9032 (I156058,I2507,I155617,I156084,);
nand I_9033 (I156092,I156084,I155750);
nor I_9034 (I155594,I156092,I155900);
nor I_9035 (I155588,I156084,I155716);
DFFARX1 I_9036 (I156084,I2507,I155617,I156146,);
not I_9037 (I156154,I156146);
nor I_9038 (I155603,I156154,I155866);
not I_9039 (I156212,I2514);
DFFARX1 I_9040 (I1382088,I2507,I156212,I156238,);
DFFARX1 I_9041 (I156238,I2507,I156212,I156255,);
not I_9042 (I156204,I156255);
not I_9043 (I156277,I156238);
DFFARX1 I_9044 (I1382079,I2507,I156212,I156303,);
not I_9045 (I156311,I156303);
and I_9046 (I156328,I156277,I1382073);
not I_9047 (I156345,I1382067);
nand I_9048 (I156362,I156345,I1382073);
not I_9049 (I156379,I1382094);
nor I_9050 (I156396,I156379,I1382067);
nand I_9051 (I156413,I156396,I1382091);
nor I_9052 (I156430,I156413,I156362);
DFFARX1 I_9053 (I156430,I2507,I156212,I156180,);
not I_9054 (I156461,I156413);
not I_9055 (I156478,I1382067);
nand I_9056 (I156495,I156478,I1382073);
nor I_9057 (I156512,I1382067,I1382067);
nand I_9058 (I156192,I156328,I156512);
nand I_9059 (I156186,I156277,I1382067);
nand I_9060 (I156557,I156379,I1382076);
DFFARX1 I_9061 (I156557,I2507,I156212,I156201,);
DFFARX1 I_9062 (I156557,I2507,I156212,I156195,);
not I_9063 (I156602,I1382076);
nor I_9064 (I156619,I156602,I1382082);
and I_9065 (I156636,I156619,I1382085);
or I_9066 (I156653,I156636,I1382070);
DFFARX1 I_9067 (I156653,I2507,I156212,I156679,);
nand I_9068 (I156687,I156679,I156345);
nor I_9069 (I156189,I156687,I156495);
nor I_9070 (I156183,I156679,I156311);
DFFARX1 I_9071 (I156679,I2507,I156212,I156741,);
not I_9072 (I156749,I156741);
nor I_9073 (I156198,I156749,I156461);
not I_9074 (I156807,I2514);
DFFARX1 I_9075 (I392487,I2507,I156807,I156833,);
DFFARX1 I_9076 (I156833,I2507,I156807,I156850,);
not I_9077 (I156799,I156850);
not I_9078 (I156872,I156833);
DFFARX1 I_9079 (I392475,I2507,I156807,I156898,);
not I_9080 (I156906,I156898);
and I_9081 (I156923,I156872,I392484);
not I_9082 (I156940,I392481);
nand I_9083 (I156957,I156940,I392484);
not I_9084 (I156974,I392472);
nor I_9085 (I156991,I156974,I392478);
nand I_9086 (I157008,I156991,I392463);
nor I_9087 (I157025,I157008,I156957);
DFFARX1 I_9088 (I157025,I2507,I156807,I156775,);
not I_9089 (I157056,I157008);
not I_9090 (I157073,I392478);
nand I_9091 (I157090,I157073,I392484);
nor I_9092 (I157107,I392478,I392481);
nand I_9093 (I156787,I156923,I157107);
nand I_9094 (I156781,I156872,I392478);
nand I_9095 (I157152,I156974,I392463);
DFFARX1 I_9096 (I157152,I2507,I156807,I156796,);
DFFARX1 I_9097 (I157152,I2507,I156807,I156790,);
not I_9098 (I157197,I392463);
nor I_9099 (I157214,I157197,I392469);
and I_9100 (I157231,I157214,I392466);
or I_9101 (I157248,I157231,I392490);
DFFARX1 I_9102 (I157248,I2507,I156807,I157274,);
nand I_9103 (I157282,I157274,I156940);
nor I_9104 (I156784,I157282,I157090);
nor I_9105 (I156778,I157274,I156906);
DFFARX1 I_9106 (I157274,I2507,I156807,I157336,);
not I_9107 (I157344,I157336);
nor I_9108 (I156793,I157344,I157056);
not I_9109 (I157402,I2514);
DFFARX1 I_9110 (I1246612,I2507,I157402,I157428,);
DFFARX1 I_9111 (I157428,I2507,I157402,I157445,);
not I_9112 (I157394,I157445);
not I_9113 (I157467,I157428);
DFFARX1 I_9114 (I1246597,I2507,I157402,I157493,);
not I_9115 (I157501,I157493);
and I_9116 (I157518,I157467,I1246615);
not I_9117 (I157535,I1246597);
nand I_9118 (I157552,I157535,I1246615);
not I_9119 (I157569,I1246618);
nor I_9120 (I157586,I157569,I1246609);
nand I_9121 (I157603,I157586,I1246606);
nor I_9122 (I157620,I157603,I157552);
DFFARX1 I_9123 (I157620,I2507,I157402,I157370,);
not I_9124 (I157651,I157603);
not I_9125 (I157668,I1246609);
nand I_9126 (I157685,I157668,I1246615);
nor I_9127 (I157702,I1246609,I1246597);
nand I_9128 (I157382,I157518,I157702);
nand I_9129 (I157376,I157467,I1246609);
nand I_9130 (I157747,I157569,I1246603);
DFFARX1 I_9131 (I157747,I2507,I157402,I157391,);
DFFARX1 I_9132 (I157747,I2507,I157402,I157385,);
not I_9133 (I157792,I1246603);
nor I_9134 (I157809,I157792,I1246594);
and I_9135 (I157826,I157809,I1246600);
or I_9136 (I157843,I157826,I1246594);
DFFARX1 I_9137 (I157843,I2507,I157402,I157869,);
nand I_9138 (I157877,I157869,I157535);
nor I_9139 (I157379,I157877,I157685);
nor I_9140 (I157373,I157869,I157501);
DFFARX1 I_9141 (I157869,I2507,I157402,I157931,);
not I_9142 (I157939,I157931);
nor I_9143 (I157388,I157939,I157651);
not I_9144 (I157997,I2514);
DFFARX1 I_9145 (I638822,I2507,I157997,I158023,);
DFFARX1 I_9146 (I158023,I2507,I157997,I158040,);
not I_9147 (I157989,I158040);
not I_9148 (I158062,I158023);
DFFARX1 I_9149 (I638819,I2507,I157997,I158088,);
not I_9150 (I158096,I158088);
and I_9151 (I158113,I158062,I638825);
not I_9152 (I158130,I638810);
nand I_9153 (I158147,I158130,I638825);
not I_9154 (I158164,I638813);
nor I_9155 (I158181,I158164,I638834);
nand I_9156 (I158198,I158181,I638831);
nor I_9157 (I158215,I158198,I158147);
DFFARX1 I_9158 (I158215,I2507,I157997,I157965,);
not I_9159 (I158246,I158198);
not I_9160 (I158263,I638834);
nand I_9161 (I158280,I158263,I638825);
nor I_9162 (I158297,I638834,I638810);
nand I_9163 (I157977,I158113,I158297);
nand I_9164 (I157971,I158062,I638834);
nand I_9165 (I158342,I158164,I638810);
DFFARX1 I_9166 (I158342,I2507,I157997,I157986,);
DFFARX1 I_9167 (I158342,I2507,I157997,I157980,);
not I_9168 (I158387,I638810);
nor I_9169 (I158404,I158387,I638816);
and I_9170 (I158421,I158404,I638828);
or I_9171 (I158438,I158421,I638813);
DFFARX1 I_9172 (I158438,I2507,I157997,I158464,);
nand I_9173 (I158472,I158464,I158130);
nor I_9174 (I157974,I158472,I158280);
nor I_9175 (I157968,I158464,I158096);
DFFARX1 I_9176 (I158464,I2507,I157997,I158526,);
not I_9177 (I158534,I158526);
nor I_9178 (I157983,I158534,I158246);
not I_9179 (I158592,I2514);
DFFARX1 I_9180 (I1149116,I2507,I158592,I158618,);
DFFARX1 I_9181 (I158618,I2507,I158592,I158635,);
not I_9182 (I158584,I158635);
not I_9183 (I158657,I158618);
DFFARX1 I_9184 (I1149116,I2507,I158592,I158683,);
not I_9185 (I158691,I158683);
and I_9186 (I158708,I158657,I1149119);
not I_9187 (I158725,I1149131);
nand I_9188 (I158742,I158725,I1149119);
not I_9189 (I158759,I1149137);
nor I_9190 (I158776,I158759,I1149128);
nand I_9191 (I158793,I158776,I1149134);
nor I_9192 (I158810,I158793,I158742);
DFFARX1 I_9193 (I158810,I2507,I158592,I158560,);
not I_9194 (I158841,I158793);
not I_9195 (I158858,I1149128);
nand I_9196 (I158875,I158858,I1149119);
nor I_9197 (I158892,I1149128,I1149131);
nand I_9198 (I158572,I158708,I158892);
nand I_9199 (I158566,I158657,I1149128);
nand I_9200 (I158937,I158759,I1149125);
DFFARX1 I_9201 (I158937,I2507,I158592,I158581,);
DFFARX1 I_9202 (I158937,I2507,I158592,I158575,);
not I_9203 (I158982,I1149125);
nor I_9204 (I158999,I158982,I1149122);
and I_9205 (I159016,I158999,I1149140);
or I_9206 (I159033,I159016,I1149119);
DFFARX1 I_9207 (I159033,I2507,I158592,I159059,);
nand I_9208 (I159067,I159059,I158725);
nor I_9209 (I158569,I159067,I158875);
nor I_9210 (I158563,I159059,I158691);
DFFARX1 I_9211 (I159059,I2507,I158592,I159121,);
not I_9212 (I159129,I159121);
nor I_9213 (I158578,I159129,I158841);
not I_9214 (I159187,I2514);
DFFARX1 I_9215 (I1359478,I2507,I159187,I159213,);
DFFARX1 I_9216 (I159213,I2507,I159187,I159230,);
not I_9217 (I159179,I159230);
not I_9218 (I159252,I159213);
DFFARX1 I_9219 (I1359469,I2507,I159187,I159278,);
not I_9220 (I159286,I159278);
and I_9221 (I159303,I159252,I1359463);
not I_9222 (I159320,I1359457);
nand I_9223 (I159337,I159320,I1359463);
not I_9224 (I159354,I1359484);
nor I_9225 (I159371,I159354,I1359457);
nand I_9226 (I159388,I159371,I1359481);
nor I_9227 (I159405,I159388,I159337);
DFFARX1 I_9228 (I159405,I2507,I159187,I159155,);
not I_9229 (I159436,I159388);
not I_9230 (I159453,I1359457);
nand I_9231 (I159470,I159453,I1359463);
nor I_9232 (I159487,I1359457,I1359457);
nand I_9233 (I159167,I159303,I159487);
nand I_9234 (I159161,I159252,I1359457);
nand I_9235 (I159532,I159354,I1359466);
DFFARX1 I_9236 (I159532,I2507,I159187,I159176,);
DFFARX1 I_9237 (I159532,I2507,I159187,I159170,);
not I_9238 (I159577,I1359466);
nor I_9239 (I159594,I159577,I1359472);
and I_9240 (I159611,I159594,I1359475);
or I_9241 (I159628,I159611,I1359460);
DFFARX1 I_9242 (I159628,I2507,I159187,I159654,);
nand I_9243 (I159662,I159654,I159320);
nor I_9244 (I159164,I159662,I159470);
nor I_9245 (I159158,I159654,I159286);
DFFARX1 I_9246 (I159654,I2507,I159187,I159716,);
not I_9247 (I159724,I159716);
nor I_9248 (I159173,I159724,I159436);
not I_9249 (I159782,I2514);
DFFARX1 I_9250 (I1129464,I2507,I159782,I159808,);
DFFARX1 I_9251 (I159808,I2507,I159782,I159825,);
not I_9252 (I159774,I159825);
not I_9253 (I159847,I159808);
DFFARX1 I_9254 (I1129464,I2507,I159782,I159873,);
not I_9255 (I159881,I159873);
and I_9256 (I159898,I159847,I1129467);
not I_9257 (I159915,I1129479);
nand I_9258 (I159932,I159915,I1129467);
not I_9259 (I159949,I1129485);
nor I_9260 (I159966,I159949,I1129476);
nand I_9261 (I159983,I159966,I1129482);
nor I_9262 (I160000,I159983,I159932);
DFFARX1 I_9263 (I160000,I2507,I159782,I159750,);
not I_9264 (I160031,I159983);
not I_9265 (I160048,I1129476);
nand I_9266 (I160065,I160048,I1129467);
nor I_9267 (I160082,I1129476,I1129479);
nand I_9268 (I159762,I159898,I160082);
nand I_9269 (I159756,I159847,I1129476);
nand I_9270 (I160127,I159949,I1129473);
DFFARX1 I_9271 (I160127,I2507,I159782,I159771,);
DFFARX1 I_9272 (I160127,I2507,I159782,I159765,);
not I_9273 (I160172,I1129473);
nor I_9274 (I160189,I160172,I1129470);
and I_9275 (I160206,I160189,I1129488);
or I_9276 (I160223,I160206,I1129467);
DFFARX1 I_9277 (I160223,I2507,I159782,I160249,);
nand I_9278 (I160257,I160249,I159915);
nor I_9279 (I159759,I160257,I160065);
nor I_9280 (I159753,I160249,I159881);
DFFARX1 I_9281 (I160249,I2507,I159782,I160311,);
not I_9282 (I160319,I160311);
nor I_9283 (I159768,I160319,I160031);
not I_9284 (I160377,I2514);
DFFARX1 I_9285 (I1360073,I2507,I160377,I160403,);
DFFARX1 I_9286 (I160403,I2507,I160377,I160420,);
not I_9287 (I160369,I160420);
not I_9288 (I160442,I160403);
DFFARX1 I_9289 (I1360064,I2507,I160377,I160468,);
not I_9290 (I160476,I160468);
and I_9291 (I160493,I160442,I1360058);
not I_9292 (I160510,I1360052);
nand I_9293 (I160527,I160510,I1360058);
not I_9294 (I160544,I1360079);
nor I_9295 (I160561,I160544,I1360052);
nand I_9296 (I160578,I160561,I1360076);
nor I_9297 (I160595,I160578,I160527);
DFFARX1 I_9298 (I160595,I2507,I160377,I160345,);
not I_9299 (I160626,I160578);
not I_9300 (I160643,I1360052);
nand I_9301 (I160660,I160643,I1360058);
nor I_9302 (I160677,I1360052,I1360052);
nand I_9303 (I160357,I160493,I160677);
nand I_9304 (I160351,I160442,I1360052);
nand I_9305 (I160722,I160544,I1360061);
DFFARX1 I_9306 (I160722,I2507,I160377,I160366,);
DFFARX1 I_9307 (I160722,I2507,I160377,I160360,);
not I_9308 (I160767,I1360061);
nor I_9309 (I160784,I160767,I1360067);
and I_9310 (I160801,I160784,I1360070);
or I_9311 (I160818,I160801,I1360055);
DFFARX1 I_9312 (I160818,I2507,I160377,I160844,);
nand I_9313 (I160852,I160844,I160510);
nor I_9314 (I160354,I160852,I160660);
nor I_9315 (I160348,I160844,I160476);
DFFARX1 I_9316 (I160844,I2507,I160377,I160906,);
not I_9317 (I160914,I160906);
nor I_9318 (I160363,I160914,I160626);
not I_9319 (I160972,I2514);
DFFARX1 I_9320 (I94921,I2507,I160972,I160998,);
DFFARX1 I_9321 (I160998,I2507,I160972,I161015,);
not I_9322 (I160964,I161015);
not I_9323 (I161037,I160998);
DFFARX1 I_9324 (I94915,I2507,I160972,I161063,);
not I_9325 (I161071,I161063);
and I_9326 (I161088,I161037,I94912);
not I_9327 (I161105,I94933);
nand I_9328 (I161122,I161105,I94912);
not I_9329 (I161139,I94927);
nor I_9330 (I161156,I161139,I94918);
nand I_9331 (I161173,I161156,I94924);
nor I_9332 (I161190,I161173,I161122);
DFFARX1 I_9333 (I161190,I2507,I160972,I160940,);
not I_9334 (I161221,I161173);
not I_9335 (I161238,I94918);
nand I_9336 (I161255,I161238,I94912);
nor I_9337 (I161272,I94918,I94933);
nand I_9338 (I160952,I161088,I161272);
nand I_9339 (I160946,I161037,I94918);
nand I_9340 (I161317,I161139,I94912);
DFFARX1 I_9341 (I161317,I2507,I160972,I160961,);
DFFARX1 I_9342 (I161317,I2507,I160972,I160955,);
not I_9343 (I161362,I94912);
nor I_9344 (I161379,I161362,I94930);
and I_9345 (I161396,I161379,I94936);
or I_9346 (I161413,I161396,I94915);
DFFARX1 I_9347 (I161413,I2507,I160972,I161439,);
nand I_9348 (I161447,I161439,I161105);
nor I_9349 (I160949,I161447,I161255);
nor I_9350 (I160943,I161439,I161071);
DFFARX1 I_9351 (I161439,I2507,I160972,I161501,);
not I_9352 (I161509,I161501);
nor I_9353 (I160958,I161509,I161221);
not I_9354 (I161567,I2514);
DFFARX1 I_9355 (I127595,I2507,I161567,I161593,);
DFFARX1 I_9356 (I161593,I2507,I161567,I161610,);
not I_9357 (I161559,I161610);
not I_9358 (I161632,I161593);
DFFARX1 I_9359 (I127589,I2507,I161567,I161658,);
not I_9360 (I161666,I161658);
and I_9361 (I161683,I161632,I127586);
not I_9362 (I161700,I127607);
nand I_9363 (I161717,I161700,I127586);
not I_9364 (I161734,I127601);
nor I_9365 (I161751,I161734,I127592);
nand I_9366 (I161768,I161751,I127598);
nor I_9367 (I161785,I161768,I161717);
DFFARX1 I_9368 (I161785,I2507,I161567,I161535,);
not I_9369 (I161816,I161768);
not I_9370 (I161833,I127592);
nand I_9371 (I161850,I161833,I127586);
nor I_9372 (I161867,I127592,I127607);
nand I_9373 (I161547,I161683,I161867);
nand I_9374 (I161541,I161632,I127592);
nand I_9375 (I161912,I161734,I127586);
DFFARX1 I_9376 (I161912,I2507,I161567,I161556,);
DFFARX1 I_9377 (I161912,I2507,I161567,I161550,);
not I_9378 (I161957,I127586);
nor I_9379 (I161974,I161957,I127604);
and I_9380 (I161991,I161974,I127610);
or I_9381 (I162008,I161991,I127589);
DFFARX1 I_9382 (I162008,I2507,I161567,I162034,);
nand I_9383 (I162042,I162034,I161700);
nor I_9384 (I161544,I162042,I161850);
nor I_9385 (I161538,I162034,I161666);
DFFARX1 I_9386 (I162034,I2507,I161567,I162096,);
not I_9387 (I162104,I162096);
nor I_9388 (I161553,I162104,I161816);
not I_9389 (I162162,I2514);
DFFARX1 I_9390 (I642290,I2507,I162162,I162188,);
DFFARX1 I_9391 (I162188,I2507,I162162,I162205,);
not I_9392 (I162154,I162205);
not I_9393 (I162227,I162188);
DFFARX1 I_9394 (I642287,I2507,I162162,I162253,);
not I_9395 (I162261,I162253);
and I_9396 (I162278,I162227,I642293);
not I_9397 (I162295,I642278);
nand I_9398 (I162312,I162295,I642293);
not I_9399 (I162329,I642281);
nor I_9400 (I162346,I162329,I642302);
nand I_9401 (I162363,I162346,I642299);
nor I_9402 (I162380,I162363,I162312);
DFFARX1 I_9403 (I162380,I2507,I162162,I162130,);
not I_9404 (I162411,I162363);
not I_9405 (I162428,I642302);
nand I_9406 (I162445,I162428,I642293);
nor I_9407 (I162462,I642302,I642278);
nand I_9408 (I162142,I162278,I162462);
nand I_9409 (I162136,I162227,I642302);
nand I_9410 (I162507,I162329,I642278);
DFFARX1 I_9411 (I162507,I2507,I162162,I162151,);
DFFARX1 I_9412 (I162507,I2507,I162162,I162145,);
not I_9413 (I162552,I642278);
nor I_9414 (I162569,I162552,I642284);
and I_9415 (I162586,I162569,I642296);
or I_9416 (I162603,I162586,I642281);
DFFARX1 I_9417 (I162603,I2507,I162162,I162629,);
nand I_9418 (I162637,I162629,I162295);
nor I_9419 (I162139,I162637,I162445);
nor I_9420 (I162133,I162629,I162261);
DFFARX1 I_9421 (I162629,I2507,I162162,I162691,);
not I_9422 (I162699,I162691);
nor I_9423 (I162148,I162699,I162411);
not I_9424 (I162757,I2514);
DFFARX1 I_9425 (I1313663,I2507,I162757,I162783,);
DFFARX1 I_9426 (I162783,I2507,I162757,I162800,);
not I_9427 (I162749,I162800);
not I_9428 (I162822,I162783);
DFFARX1 I_9429 (I1313654,I2507,I162757,I162848,);
not I_9430 (I162856,I162848);
and I_9431 (I162873,I162822,I1313648);
not I_9432 (I162890,I1313642);
nand I_9433 (I162907,I162890,I1313648);
not I_9434 (I162924,I1313669);
nor I_9435 (I162941,I162924,I1313642);
nand I_9436 (I162958,I162941,I1313666);
nor I_9437 (I162975,I162958,I162907);
DFFARX1 I_9438 (I162975,I2507,I162757,I162725,);
not I_9439 (I163006,I162958);
not I_9440 (I163023,I1313642);
nand I_9441 (I163040,I163023,I1313648);
nor I_9442 (I163057,I1313642,I1313642);
nand I_9443 (I162737,I162873,I163057);
nand I_9444 (I162731,I162822,I1313642);
nand I_9445 (I163102,I162924,I1313651);
DFFARX1 I_9446 (I163102,I2507,I162757,I162746,);
DFFARX1 I_9447 (I163102,I2507,I162757,I162740,);
not I_9448 (I163147,I1313651);
nor I_9449 (I163164,I163147,I1313657);
and I_9450 (I163181,I163164,I1313660);
or I_9451 (I163198,I163181,I1313645);
DFFARX1 I_9452 (I163198,I2507,I162757,I163224,);
nand I_9453 (I163232,I163224,I162890);
nor I_9454 (I162734,I163232,I163040);
nor I_9455 (I162728,I163224,I162856);
DFFARX1 I_9456 (I163224,I2507,I162757,I163286,);
not I_9457 (I163294,I163286);
nor I_9458 (I162743,I163294,I163006);
not I_9459 (I163352,I2514);
DFFARX1 I_9460 (I686218,I2507,I163352,I163378,);
DFFARX1 I_9461 (I163378,I2507,I163352,I163395,);
not I_9462 (I163344,I163395);
not I_9463 (I163417,I163378);
DFFARX1 I_9464 (I686215,I2507,I163352,I163443,);
not I_9465 (I163451,I163443);
and I_9466 (I163468,I163417,I686221);
not I_9467 (I163485,I686206);
nand I_9468 (I163502,I163485,I686221);
not I_9469 (I163519,I686209);
nor I_9470 (I163536,I163519,I686230);
nand I_9471 (I163553,I163536,I686227);
nor I_9472 (I163570,I163553,I163502);
DFFARX1 I_9473 (I163570,I2507,I163352,I163320,);
not I_9474 (I163601,I163553);
not I_9475 (I163618,I686230);
nand I_9476 (I163635,I163618,I686221);
nor I_9477 (I163652,I686230,I686206);
nand I_9478 (I163332,I163468,I163652);
nand I_9479 (I163326,I163417,I686230);
nand I_9480 (I163697,I163519,I686206);
DFFARX1 I_9481 (I163697,I2507,I163352,I163341,);
DFFARX1 I_9482 (I163697,I2507,I163352,I163335,);
not I_9483 (I163742,I686206);
nor I_9484 (I163759,I163742,I686212);
and I_9485 (I163776,I163759,I686224);
or I_9486 (I163793,I163776,I686209);
DFFARX1 I_9487 (I163793,I2507,I163352,I163819,);
nand I_9488 (I163827,I163819,I163485);
nor I_9489 (I163329,I163827,I163635);
nor I_9490 (I163323,I163819,I163451);
DFFARX1 I_9491 (I163819,I2507,I163352,I163881,);
not I_9492 (I163889,I163881);
nor I_9493 (I163338,I163889,I163601);
not I_9494 (I163947,I2514);
DFFARX1 I_9495 (I1395178,I2507,I163947,I163973,);
DFFARX1 I_9496 (I163973,I2507,I163947,I163990,);
not I_9497 (I163939,I163990);
not I_9498 (I164012,I163973);
DFFARX1 I_9499 (I1395169,I2507,I163947,I164038,);
not I_9500 (I164046,I164038);
and I_9501 (I164063,I164012,I1395163);
not I_9502 (I164080,I1395157);
nand I_9503 (I164097,I164080,I1395163);
not I_9504 (I164114,I1395184);
nor I_9505 (I164131,I164114,I1395157);
nand I_9506 (I164148,I164131,I1395181);
nor I_9507 (I164165,I164148,I164097);
DFFARX1 I_9508 (I164165,I2507,I163947,I163915,);
not I_9509 (I164196,I164148);
not I_9510 (I164213,I1395157);
nand I_9511 (I164230,I164213,I1395163);
nor I_9512 (I164247,I1395157,I1395157);
nand I_9513 (I163927,I164063,I164247);
nand I_9514 (I163921,I164012,I1395157);
nand I_9515 (I164292,I164114,I1395166);
DFFARX1 I_9516 (I164292,I2507,I163947,I163936,);
DFFARX1 I_9517 (I164292,I2507,I163947,I163930,);
not I_9518 (I164337,I1395166);
nor I_9519 (I164354,I164337,I1395172);
and I_9520 (I164371,I164354,I1395175);
or I_9521 (I164388,I164371,I1395160);
DFFARX1 I_9522 (I164388,I2507,I163947,I164414,);
nand I_9523 (I164422,I164414,I164080);
nor I_9524 (I163924,I164422,I164230);
nor I_9525 (I163918,I164414,I164046);
DFFARX1 I_9526 (I164414,I2507,I163947,I164476,);
not I_9527 (I164484,I164476);
nor I_9528 (I163933,I164484,I164196);
not I_9529 (I164542,I2514);
DFFARX1 I_9530 (I620329,I2507,I164542,I164568,);
DFFARX1 I_9531 (I164568,I2507,I164542,I164585,);
not I_9532 (I164534,I164585);
not I_9533 (I164607,I164568);
DFFARX1 I_9534 (I620320,I2507,I164542,I164633,);
not I_9535 (I164641,I164633);
and I_9536 (I164658,I164607,I620338);
not I_9537 (I164675,I620335);
nand I_9538 (I164692,I164675,I620338);
not I_9539 (I164709,I620314);
nor I_9540 (I164726,I164709,I620317);
nand I_9541 (I164743,I164726,I620326);
nor I_9542 (I164760,I164743,I164692);
DFFARX1 I_9543 (I164760,I2507,I164542,I164510,);
not I_9544 (I164791,I164743);
not I_9545 (I164808,I620317);
nand I_9546 (I164825,I164808,I620338);
nor I_9547 (I164842,I620317,I620335);
nand I_9548 (I164522,I164658,I164842);
nand I_9549 (I164516,I164607,I620317);
nand I_9550 (I164887,I164709,I620332);
DFFARX1 I_9551 (I164887,I2507,I164542,I164531,);
DFFARX1 I_9552 (I164887,I2507,I164542,I164525,);
not I_9553 (I164932,I620332);
nor I_9554 (I164949,I164932,I620314);
and I_9555 (I164966,I164949,I620323);
or I_9556 (I164983,I164966,I620317);
DFFARX1 I_9557 (I164983,I2507,I164542,I165009,);
nand I_9558 (I165017,I165009,I164675);
nor I_9559 (I164519,I165017,I164825);
nor I_9560 (I164513,I165009,I164641);
DFFARX1 I_9561 (I165009,I2507,I164542,I165071,);
not I_9562 (I165079,I165071);
nor I_9563 (I164528,I165079,I164791);
not I_9564 (I165137,I2514);
DFFARX1 I_9565 (I346104,I2507,I165137,I165163,);
DFFARX1 I_9566 (I165163,I2507,I165137,I165180,);
not I_9567 (I165129,I165180);
not I_9568 (I165202,I165163);
DFFARX1 I_9569 (I346119,I2507,I165137,I165228,);
not I_9570 (I165236,I165228);
and I_9571 (I165253,I165202,I346116);
not I_9572 (I165270,I346104);
nand I_9573 (I165287,I165270,I346116);
not I_9574 (I165304,I346113);
nor I_9575 (I165321,I165304,I346128);
nand I_9576 (I165338,I165321,I346125);
nor I_9577 (I165355,I165338,I165287);
DFFARX1 I_9578 (I165355,I2507,I165137,I165105,);
not I_9579 (I165386,I165338);
not I_9580 (I165403,I346128);
nand I_9581 (I165420,I165403,I346116);
nor I_9582 (I165437,I346128,I346104);
nand I_9583 (I165117,I165253,I165437);
nand I_9584 (I165111,I165202,I346128);
nand I_9585 (I165482,I165304,I346122);
DFFARX1 I_9586 (I165482,I2507,I165137,I165126,);
DFFARX1 I_9587 (I165482,I2507,I165137,I165120,);
not I_9588 (I165527,I346122);
nor I_9589 (I165544,I165527,I346110);
and I_9590 (I165561,I165544,I346131);
or I_9591 (I165578,I165561,I346107);
DFFARX1 I_9592 (I165578,I2507,I165137,I165604,);
nand I_9593 (I165612,I165604,I165270);
nor I_9594 (I165114,I165612,I165420);
nor I_9595 (I165108,I165604,I165236);
DFFARX1 I_9596 (I165604,I2507,I165137,I165666,);
not I_9597 (I165674,I165666);
nor I_9598 (I165123,I165674,I165386);
not I_9599 (I165732,I2514);
DFFARX1 I_9600 (I1395773,I2507,I165732,I165758,);
DFFARX1 I_9601 (I165758,I2507,I165732,I165775,);
not I_9602 (I165724,I165775);
not I_9603 (I165797,I165758);
DFFARX1 I_9604 (I1395764,I2507,I165732,I165823,);
not I_9605 (I165831,I165823);
and I_9606 (I165848,I165797,I1395758);
not I_9607 (I165865,I1395752);
nand I_9608 (I165882,I165865,I1395758);
not I_9609 (I165899,I1395779);
nor I_9610 (I165916,I165899,I1395752);
nand I_9611 (I165933,I165916,I1395776);
nor I_9612 (I165950,I165933,I165882);
DFFARX1 I_9613 (I165950,I2507,I165732,I165700,);
not I_9614 (I165981,I165933);
not I_9615 (I165998,I1395752);
nand I_9616 (I166015,I165998,I1395758);
nor I_9617 (I166032,I1395752,I1395752);
nand I_9618 (I165712,I165848,I166032);
nand I_9619 (I165706,I165797,I1395752);
nand I_9620 (I166077,I165899,I1395761);
DFFARX1 I_9621 (I166077,I2507,I165732,I165721,);
DFFARX1 I_9622 (I166077,I2507,I165732,I165715,);
not I_9623 (I166122,I1395761);
nor I_9624 (I166139,I166122,I1395767);
and I_9625 (I166156,I166139,I1395770);
or I_9626 (I166173,I166156,I1395755);
DFFARX1 I_9627 (I166173,I2507,I165732,I166199,);
nand I_9628 (I166207,I166199,I165865);
nor I_9629 (I165709,I166207,I166015);
nor I_9630 (I165703,I166199,I165831);
DFFARX1 I_9631 (I166199,I2507,I165732,I166261,);
not I_9632 (I166269,I166261);
nor I_9633 (I165718,I166269,I165981);
not I_9634 (I166327,I2514);
DFFARX1 I_9635 (I82273,I2507,I166327,I166353,);
DFFARX1 I_9636 (I166353,I2507,I166327,I166370,);
not I_9637 (I166319,I166370);
not I_9638 (I166392,I166353);
DFFARX1 I_9639 (I82267,I2507,I166327,I166418,);
not I_9640 (I166426,I166418);
and I_9641 (I166443,I166392,I82264);
not I_9642 (I166460,I82285);
nand I_9643 (I166477,I166460,I82264);
not I_9644 (I166494,I82279);
nor I_9645 (I166511,I166494,I82270);
nand I_9646 (I166528,I166511,I82276);
nor I_9647 (I166545,I166528,I166477);
DFFARX1 I_9648 (I166545,I2507,I166327,I166295,);
not I_9649 (I166576,I166528);
not I_9650 (I166593,I82270);
nand I_9651 (I166610,I166593,I82264);
nor I_9652 (I166627,I82270,I82285);
nand I_9653 (I166307,I166443,I166627);
nand I_9654 (I166301,I166392,I82270);
nand I_9655 (I166672,I166494,I82264);
DFFARX1 I_9656 (I166672,I2507,I166327,I166316,);
DFFARX1 I_9657 (I166672,I2507,I166327,I166310,);
not I_9658 (I166717,I82264);
nor I_9659 (I166734,I166717,I82282);
and I_9660 (I166751,I166734,I82288);
or I_9661 (I166768,I166751,I82267);
DFFARX1 I_9662 (I166768,I2507,I166327,I166794,);
nand I_9663 (I166802,I166794,I166460);
nor I_9664 (I166304,I166802,I166610);
nor I_9665 (I166298,I166794,I166426);
DFFARX1 I_9666 (I166794,I2507,I166327,I166856,);
not I_9667 (I166864,I166856);
nor I_9668 (I166313,I166864,I166576);
not I_9669 (I166922,I2514);
DFFARX1 I_9670 (I643446,I2507,I166922,I166948,);
DFFARX1 I_9671 (I166948,I2507,I166922,I166965,);
not I_9672 (I166914,I166965);
not I_9673 (I166987,I166948);
DFFARX1 I_9674 (I643443,I2507,I166922,I167013,);
not I_9675 (I167021,I167013);
and I_9676 (I167038,I166987,I643449);
not I_9677 (I167055,I643434);
nand I_9678 (I167072,I167055,I643449);
not I_9679 (I167089,I643437);
nor I_9680 (I167106,I167089,I643458);
nand I_9681 (I167123,I167106,I643455);
nor I_9682 (I167140,I167123,I167072);
DFFARX1 I_9683 (I167140,I2507,I166922,I166890,);
not I_9684 (I167171,I167123);
not I_9685 (I167188,I643458);
nand I_9686 (I167205,I167188,I643449);
nor I_9687 (I167222,I643458,I643434);
nand I_9688 (I166902,I167038,I167222);
nand I_9689 (I166896,I166987,I643458);
nand I_9690 (I167267,I167089,I643434);
DFFARX1 I_9691 (I167267,I2507,I166922,I166911,);
DFFARX1 I_9692 (I167267,I2507,I166922,I166905,);
not I_9693 (I167312,I643434);
nor I_9694 (I167329,I167312,I643440);
and I_9695 (I167346,I167329,I643452);
or I_9696 (I167363,I167346,I643437);
DFFARX1 I_9697 (I167363,I2507,I166922,I167389,);
nand I_9698 (I167397,I167389,I167055);
nor I_9699 (I166899,I167397,I167205);
nor I_9700 (I166893,I167389,I167021);
DFFARX1 I_9701 (I167389,I2507,I166922,I167451,);
not I_9702 (I167459,I167451);
nor I_9703 (I166908,I167459,I167171);
not I_9704 (I167517,I2514);
DFFARX1 I_9705 (I388135,I2507,I167517,I167543,);
DFFARX1 I_9706 (I167543,I2507,I167517,I167560,);
not I_9707 (I167509,I167560);
not I_9708 (I167582,I167543);
DFFARX1 I_9709 (I388123,I2507,I167517,I167608,);
not I_9710 (I167616,I167608);
and I_9711 (I167633,I167582,I388132);
not I_9712 (I167650,I388129);
nand I_9713 (I167667,I167650,I388132);
not I_9714 (I167684,I388120);
nor I_9715 (I167701,I167684,I388126);
nand I_9716 (I167718,I167701,I388111);
nor I_9717 (I167735,I167718,I167667);
DFFARX1 I_9718 (I167735,I2507,I167517,I167485,);
not I_9719 (I167766,I167718);
not I_9720 (I167783,I388126);
nand I_9721 (I167800,I167783,I388132);
nor I_9722 (I167817,I388126,I388129);
nand I_9723 (I167497,I167633,I167817);
nand I_9724 (I167491,I167582,I388126);
nand I_9725 (I167862,I167684,I388111);
DFFARX1 I_9726 (I167862,I2507,I167517,I167506,);
DFFARX1 I_9727 (I167862,I2507,I167517,I167500,);
not I_9728 (I167907,I388111);
nor I_9729 (I167924,I167907,I388117);
and I_9730 (I167941,I167924,I388114);
or I_9731 (I167958,I167941,I388138);
DFFARX1 I_9732 (I167958,I2507,I167517,I167984,);
nand I_9733 (I167992,I167984,I167650);
nor I_9734 (I167494,I167992,I167800);
nor I_9735 (I167488,I167984,I167616);
DFFARX1 I_9736 (I167984,I2507,I167517,I168046,);
not I_9737 (I168054,I168046);
nor I_9738 (I167503,I168054,I167766);
not I_9739 (I168112,I2514);
DFFARX1 I_9740 (I1190732,I2507,I168112,I168138,);
DFFARX1 I_9741 (I168138,I2507,I168112,I168155,);
not I_9742 (I168104,I168155);
not I_9743 (I168177,I168138);
DFFARX1 I_9744 (I1190732,I2507,I168112,I168203,);
not I_9745 (I168211,I168203);
and I_9746 (I168228,I168177,I1190735);
not I_9747 (I168245,I1190747);
nand I_9748 (I168262,I168245,I1190735);
not I_9749 (I168279,I1190753);
nor I_9750 (I168296,I168279,I1190744);
nand I_9751 (I168313,I168296,I1190750);
nor I_9752 (I168330,I168313,I168262);
DFFARX1 I_9753 (I168330,I2507,I168112,I168080,);
not I_9754 (I168361,I168313);
not I_9755 (I168378,I1190744);
nand I_9756 (I168395,I168378,I1190735);
nor I_9757 (I168412,I1190744,I1190747);
nand I_9758 (I168092,I168228,I168412);
nand I_9759 (I168086,I168177,I1190744);
nand I_9760 (I168457,I168279,I1190741);
DFFARX1 I_9761 (I168457,I2507,I168112,I168101,);
DFFARX1 I_9762 (I168457,I2507,I168112,I168095,);
not I_9763 (I168502,I1190741);
nor I_9764 (I168519,I168502,I1190738);
and I_9765 (I168536,I168519,I1190756);
or I_9766 (I168553,I168536,I1190735);
DFFARX1 I_9767 (I168553,I2507,I168112,I168579,);
nand I_9768 (I168587,I168579,I168245);
nor I_9769 (I168089,I168587,I168395);
nor I_9770 (I168083,I168579,I168211);
DFFARX1 I_9771 (I168579,I2507,I168112,I168641,);
not I_9772 (I168649,I168641);
nor I_9773 (I168098,I168649,I168361);
not I_9774 (I168707,I2514);
DFFARX1 I_9775 (I257041,I2507,I168707,I168733,);
DFFARX1 I_9776 (I168733,I2507,I168707,I168750,);
not I_9777 (I168699,I168750);
not I_9778 (I168772,I168733);
DFFARX1 I_9779 (I257056,I2507,I168707,I168798,);
not I_9780 (I168806,I168798);
and I_9781 (I168823,I168772,I257053);
not I_9782 (I168840,I257041);
nand I_9783 (I168857,I168840,I257053);
not I_9784 (I168874,I257050);
nor I_9785 (I168891,I168874,I257065);
nand I_9786 (I168908,I168891,I257062);
nor I_9787 (I168925,I168908,I168857);
DFFARX1 I_9788 (I168925,I2507,I168707,I168675,);
not I_9789 (I168956,I168908);
not I_9790 (I168973,I257065);
nand I_9791 (I168990,I168973,I257053);
nor I_9792 (I169007,I257065,I257041);
nand I_9793 (I168687,I168823,I169007);
nand I_9794 (I168681,I168772,I257065);
nand I_9795 (I169052,I168874,I257059);
DFFARX1 I_9796 (I169052,I2507,I168707,I168696,);
DFFARX1 I_9797 (I169052,I2507,I168707,I168690,);
not I_9798 (I169097,I257059);
nor I_9799 (I169114,I169097,I257047);
and I_9800 (I169131,I169114,I257068);
or I_9801 (I169148,I169131,I257044);
DFFARX1 I_9802 (I169148,I2507,I168707,I169174,);
nand I_9803 (I169182,I169174,I168840);
nor I_9804 (I168684,I169182,I168990);
nor I_9805 (I168678,I169174,I168806);
DFFARX1 I_9806 (I169174,I2507,I168707,I169236,);
not I_9807 (I169244,I169236);
nor I_9808 (I168693,I169244,I168956);
not I_9809 (I169302,I2514);
DFFARX1 I_9810 (I430023,I2507,I169302,I169328,);
DFFARX1 I_9811 (I169328,I2507,I169302,I169345,);
not I_9812 (I169294,I169345);
not I_9813 (I169367,I169328);
DFFARX1 I_9814 (I430011,I2507,I169302,I169393,);
not I_9815 (I169401,I169393);
and I_9816 (I169418,I169367,I430020);
not I_9817 (I169435,I430017);
nand I_9818 (I169452,I169435,I430020);
not I_9819 (I169469,I430008);
nor I_9820 (I169486,I169469,I430014);
nand I_9821 (I169503,I169486,I429999);
nor I_9822 (I169520,I169503,I169452);
DFFARX1 I_9823 (I169520,I2507,I169302,I169270,);
not I_9824 (I169551,I169503);
not I_9825 (I169568,I430014);
nand I_9826 (I169585,I169568,I430020);
nor I_9827 (I169602,I430014,I430017);
nand I_9828 (I169282,I169418,I169602);
nand I_9829 (I169276,I169367,I430014);
nand I_9830 (I169647,I169469,I429999);
DFFARX1 I_9831 (I169647,I2507,I169302,I169291,);
DFFARX1 I_9832 (I169647,I2507,I169302,I169285,);
not I_9833 (I169692,I429999);
nor I_9834 (I169709,I169692,I430005);
and I_9835 (I169726,I169709,I430002);
or I_9836 (I169743,I169726,I430026);
DFFARX1 I_9837 (I169743,I2507,I169302,I169769,);
nand I_9838 (I169777,I169769,I169435);
nor I_9839 (I169279,I169777,I169585);
nor I_9840 (I169273,I169769,I169401);
DFFARX1 I_9841 (I169769,I2507,I169302,I169831,);
not I_9842 (I169839,I169831);
nor I_9843 (I169288,I169839,I169551);
not I_9844 (I169897,I2514);
DFFARX1 I_9845 (I847576,I2507,I169897,I169923,);
DFFARX1 I_9846 (I169923,I2507,I169897,I169940,);
not I_9847 (I169889,I169940);
not I_9848 (I169962,I169923);
DFFARX1 I_9849 (I847570,I2507,I169897,I169988,);
not I_9850 (I169996,I169988);
and I_9851 (I170013,I169962,I847588);
not I_9852 (I170030,I847576);
nand I_9853 (I170047,I170030,I847588);
not I_9854 (I170064,I847570);
nor I_9855 (I170081,I170064,I847582);
nand I_9856 (I170098,I170081,I847573);
nor I_9857 (I170115,I170098,I170047);
DFFARX1 I_9858 (I170115,I2507,I169897,I169865,);
not I_9859 (I170146,I170098);
not I_9860 (I170163,I847582);
nand I_9861 (I170180,I170163,I847588);
nor I_9862 (I170197,I847582,I847576);
nand I_9863 (I169877,I170013,I170197);
nand I_9864 (I169871,I169962,I847582);
nand I_9865 (I170242,I170064,I847585);
DFFARX1 I_9866 (I170242,I2507,I169897,I169886,);
DFFARX1 I_9867 (I170242,I2507,I169897,I169880,);
not I_9868 (I170287,I847585);
nor I_9869 (I170304,I170287,I847591);
and I_9870 (I170321,I170304,I847573);
or I_9871 (I170338,I170321,I847579);
DFFARX1 I_9872 (I170338,I2507,I169897,I170364,);
nand I_9873 (I170372,I170364,I170030);
nor I_9874 (I169874,I170372,I170180);
nor I_9875 (I169868,I170364,I169996);
DFFARX1 I_9876 (I170364,I2507,I169897,I170426,);
not I_9877 (I170434,I170426);
nor I_9878 (I169883,I170434,I170146);
not I_9879 (I170492,I2514);
DFFARX1 I_9880 (I36966,I2507,I170492,I170518,);
DFFARX1 I_9881 (I170518,I2507,I170492,I170535,);
not I_9882 (I170484,I170535);
not I_9883 (I170557,I170518);
DFFARX1 I_9884 (I36942,I2507,I170492,I170583,);
not I_9885 (I170591,I170583);
and I_9886 (I170608,I170557,I36957);
not I_9887 (I170625,I36945);
nand I_9888 (I170642,I170625,I36957);
not I_9889 (I170659,I36948);
nor I_9890 (I170676,I170659,I36960);
nand I_9891 (I170693,I170676,I36951);
nor I_9892 (I170710,I170693,I170642);
DFFARX1 I_9893 (I170710,I2507,I170492,I170460,);
not I_9894 (I170741,I170693);
not I_9895 (I170758,I36960);
nand I_9896 (I170775,I170758,I36957);
nor I_9897 (I170792,I36960,I36945);
nand I_9898 (I170472,I170608,I170792);
nand I_9899 (I170466,I170557,I36960);
nand I_9900 (I170837,I170659,I36954);
DFFARX1 I_9901 (I170837,I2507,I170492,I170481,);
DFFARX1 I_9902 (I170837,I2507,I170492,I170475,);
not I_9903 (I170882,I36954);
nor I_9904 (I170899,I170882,I36945);
and I_9905 (I170916,I170899,I36942);
or I_9906 (I170933,I170916,I36963);
DFFARX1 I_9907 (I170933,I2507,I170492,I170959,);
nand I_9908 (I170967,I170959,I170625);
nor I_9909 (I170469,I170967,I170775);
nor I_9910 (I170463,I170959,I170591);
DFFARX1 I_9911 (I170959,I2507,I170492,I171021,);
not I_9912 (I171029,I171021);
nor I_9913 (I170478,I171029,I170741);
not I_9914 (I171087,I2514);
DFFARX1 I_9915 (I117582,I2507,I171087,I171113,);
DFFARX1 I_9916 (I171113,I2507,I171087,I171130,);
not I_9917 (I171079,I171130);
not I_9918 (I171152,I171113);
DFFARX1 I_9919 (I117576,I2507,I171087,I171178,);
not I_9920 (I171186,I171178);
and I_9921 (I171203,I171152,I117573);
not I_9922 (I171220,I117594);
nand I_9923 (I171237,I171220,I117573);
not I_9924 (I171254,I117588);
nor I_9925 (I171271,I171254,I117579);
nand I_9926 (I171288,I171271,I117585);
nor I_9927 (I171305,I171288,I171237);
DFFARX1 I_9928 (I171305,I2507,I171087,I171055,);
not I_9929 (I171336,I171288);
not I_9930 (I171353,I117579);
nand I_9931 (I171370,I171353,I117573);
nor I_9932 (I171387,I117579,I117594);
nand I_9933 (I171067,I171203,I171387);
nand I_9934 (I171061,I171152,I117579);
nand I_9935 (I171432,I171254,I117573);
DFFARX1 I_9936 (I171432,I2507,I171087,I171076,);
DFFARX1 I_9937 (I171432,I2507,I171087,I171070,);
not I_9938 (I171477,I117573);
nor I_9939 (I171494,I171477,I117591);
and I_9940 (I171511,I171494,I117597);
or I_9941 (I171528,I171511,I117576);
DFFARX1 I_9942 (I171528,I2507,I171087,I171554,);
nand I_9943 (I171562,I171554,I171220);
nor I_9944 (I171064,I171562,I171370);
nor I_9945 (I171058,I171554,I171186);
DFFARX1 I_9946 (I171554,I2507,I171087,I171616,);
not I_9947 (I171624,I171616);
nor I_9948 (I171073,I171624,I171336);
not I_9949 (I171682,I2514);
DFFARX1 I_9950 (I660786,I2507,I171682,I171708,);
DFFARX1 I_9951 (I171708,I2507,I171682,I171725,);
not I_9952 (I171674,I171725);
not I_9953 (I171747,I171708);
DFFARX1 I_9954 (I660783,I2507,I171682,I171773,);
not I_9955 (I171781,I171773);
and I_9956 (I171798,I171747,I660789);
not I_9957 (I171815,I660774);
nand I_9958 (I171832,I171815,I660789);
not I_9959 (I171849,I660777);
nor I_9960 (I171866,I171849,I660798);
nand I_9961 (I171883,I171866,I660795);
nor I_9962 (I171900,I171883,I171832);
DFFARX1 I_9963 (I171900,I2507,I171682,I171650,);
not I_9964 (I171931,I171883);
not I_9965 (I171948,I660798);
nand I_9966 (I171965,I171948,I660789);
nor I_9967 (I171982,I660798,I660774);
nand I_9968 (I171662,I171798,I171982);
nand I_9969 (I171656,I171747,I660798);
nand I_9970 (I172027,I171849,I660774);
DFFARX1 I_9971 (I172027,I2507,I171682,I171671,);
DFFARX1 I_9972 (I172027,I2507,I171682,I171665,);
not I_9973 (I172072,I660774);
nor I_9974 (I172089,I172072,I660780);
and I_9975 (I172106,I172089,I660792);
or I_9976 (I172123,I172106,I660777);
DFFARX1 I_9977 (I172123,I2507,I171682,I172149,);
nand I_9978 (I172157,I172149,I171815);
nor I_9979 (I171659,I172157,I171965);
nor I_9980 (I171653,I172149,I171781);
DFFARX1 I_9981 (I172149,I2507,I171682,I172211,);
not I_9982 (I172219,I172211);
nor I_9983 (I171668,I172219,I171931);
not I_9984 (I172277,I2514);
DFFARX1 I_9985 (I1272097,I2507,I172277,I172303,);
DFFARX1 I_9986 (I172303,I2507,I172277,I172320,);
not I_9987 (I172269,I172320);
not I_9988 (I172342,I172303);
DFFARX1 I_9989 (I1272109,I2507,I172277,I172368,);
not I_9990 (I172376,I172368);
and I_9991 (I172393,I172342,I1272103);
not I_9992 (I172410,I1272115);
nand I_9993 (I172427,I172410,I1272103);
not I_9994 (I172444,I1272100);
nor I_9995 (I172461,I172444,I1272112);
nand I_9996 (I172478,I172461,I1272094);
nor I_9997 (I172495,I172478,I172427);
DFFARX1 I_9998 (I172495,I2507,I172277,I172245,);
not I_9999 (I172526,I172478);
not I_10000 (I172543,I1272112);
nand I_10001 (I172560,I172543,I1272103);
nor I_10002 (I172577,I1272112,I1272115);
nand I_10003 (I172257,I172393,I172577);
nand I_10004 (I172251,I172342,I1272112);
nand I_10005 (I172622,I172444,I1272106);
DFFARX1 I_10006 (I172622,I2507,I172277,I172266,);
DFFARX1 I_10007 (I172622,I2507,I172277,I172260,);
not I_10008 (I172667,I1272106);
nor I_10009 (I172684,I172667,I1272097);
and I_10010 (I172701,I172684,I1272094);
or I_10011 (I172718,I172701,I1272118);
DFFARX1 I_10012 (I172718,I2507,I172277,I172744,);
nand I_10013 (I172752,I172744,I172410);
nor I_10014 (I172254,I172752,I172560);
nor I_10015 (I172248,I172744,I172376);
DFFARX1 I_10016 (I172744,I2507,I172277,I172806,);
not I_10017 (I172814,I172806);
nor I_10018 (I172263,I172814,I172526);
not I_10019 (I172872,I2514);
DFFARX1 I_10020 (I1073398,I2507,I172872,I172898,);
DFFARX1 I_10021 (I172898,I2507,I172872,I172915,);
not I_10022 (I172864,I172915);
not I_10023 (I172937,I172898);
DFFARX1 I_10024 (I1073398,I2507,I172872,I172963,);
not I_10025 (I172971,I172963);
and I_10026 (I172988,I172937,I1073401);
not I_10027 (I173005,I1073413);
nand I_10028 (I173022,I173005,I1073401);
not I_10029 (I173039,I1073419);
nor I_10030 (I173056,I173039,I1073410);
nand I_10031 (I173073,I173056,I1073416);
nor I_10032 (I173090,I173073,I173022);
DFFARX1 I_10033 (I173090,I2507,I172872,I172840,);
not I_10034 (I173121,I173073);
not I_10035 (I173138,I1073410);
nand I_10036 (I173155,I173138,I1073401);
nor I_10037 (I173172,I1073410,I1073413);
nand I_10038 (I172852,I172988,I173172);
nand I_10039 (I172846,I172937,I1073410);
nand I_10040 (I173217,I173039,I1073407);
DFFARX1 I_10041 (I173217,I2507,I172872,I172861,);
DFFARX1 I_10042 (I173217,I2507,I172872,I172855,);
not I_10043 (I173262,I1073407);
nor I_10044 (I173279,I173262,I1073404);
and I_10045 (I173296,I173279,I1073422);
or I_10046 (I173313,I173296,I1073401);
DFFARX1 I_10047 (I173313,I2507,I172872,I173339,);
nand I_10048 (I173347,I173339,I173005);
nor I_10049 (I172849,I173347,I173155);
nor I_10050 (I172843,I173339,I172971);
DFFARX1 I_10051 (I173339,I2507,I172872,I173401,);
not I_10052 (I173409,I173401);
nor I_10053 (I172858,I173409,I173121);
not I_10054 (I173467,I2514);
DFFARX1 I_10055 (I444711,I2507,I173467,I173493,);
DFFARX1 I_10056 (I173493,I2507,I173467,I173510,);
not I_10057 (I173459,I173510);
not I_10058 (I173532,I173493);
DFFARX1 I_10059 (I444699,I2507,I173467,I173558,);
not I_10060 (I173566,I173558);
and I_10061 (I173583,I173532,I444708);
not I_10062 (I173600,I444705);
nand I_10063 (I173617,I173600,I444708);
not I_10064 (I173634,I444696);
nor I_10065 (I173651,I173634,I444702);
nand I_10066 (I173668,I173651,I444687);
nor I_10067 (I173685,I173668,I173617);
DFFARX1 I_10068 (I173685,I2507,I173467,I173435,);
not I_10069 (I173716,I173668);
not I_10070 (I173733,I444702);
nand I_10071 (I173750,I173733,I444708);
nor I_10072 (I173767,I444702,I444705);
nand I_10073 (I173447,I173583,I173767);
nand I_10074 (I173441,I173532,I444702);
nand I_10075 (I173812,I173634,I444687);
DFFARX1 I_10076 (I173812,I2507,I173467,I173456,);
DFFARX1 I_10077 (I173812,I2507,I173467,I173450,);
not I_10078 (I173857,I444687);
nor I_10079 (I173874,I173857,I444693);
and I_10080 (I173891,I173874,I444690);
or I_10081 (I173908,I173891,I444714);
DFFARX1 I_10082 (I173908,I2507,I173467,I173934,);
nand I_10083 (I173942,I173934,I173600);
nor I_10084 (I173444,I173942,I173750);
nor I_10085 (I173438,I173934,I173566);
DFFARX1 I_10086 (I173934,I2507,I173467,I173996,);
not I_10087 (I174004,I173996);
nor I_10088 (I173453,I174004,I173716);
not I_10089 (I174062,I2514);
DFFARX1 I_10090 (I1012949,I2507,I174062,I174088,);
DFFARX1 I_10091 (I174088,I2507,I174062,I174105,);
not I_10092 (I174054,I174105);
not I_10093 (I174127,I174088);
DFFARX1 I_10094 (I1012958,I2507,I174062,I174153,);
not I_10095 (I174161,I174153);
and I_10096 (I174178,I174127,I1012952);
not I_10097 (I174195,I1012946);
nand I_10098 (I174212,I174195,I1012952);
not I_10099 (I174229,I1012961);
nor I_10100 (I174246,I174229,I1012949);
nand I_10101 (I174263,I174246,I1012955);
nor I_10102 (I174280,I174263,I174212);
DFFARX1 I_10103 (I174280,I2507,I174062,I174030,);
not I_10104 (I174311,I174263);
not I_10105 (I174328,I1012949);
nand I_10106 (I174345,I174328,I1012952);
nor I_10107 (I174362,I1012949,I1012946);
nand I_10108 (I174042,I174178,I174362);
nand I_10109 (I174036,I174127,I1012949);
nand I_10110 (I174407,I174229,I1012952);
DFFARX1 I_10111 (I174407,I2507,I174062,I174051,);
DFFARX1 I_10112 (I174407,I2507,I174062,I174045,);
not I_10113 (I174452,I1012952);
nor I_10114 (I174469,I174452,I1012967);
and I_10115 (I174486,I174469,I1012964);
or I_10116 (I174503,I174486,I1012946);
DFFARX1 I_10117 (I174503,I2507,I174062,I174529,);
nand I_10118 (I174537,I174529,I174195);
nor I_10119 (I174039,I174537,I174345);
nor I_10120 (I174033,I174529,I174161);
DFFARX1 I_10121 (I174529,I2507,I174062,I174591,);
not I_10122 (I174599,I174591);
nor I_10123 (I174048,I174599,I174311);
not I_10124 (I174657,I2514);
DFFARX1 I_10125 (I575245,I2507,I174657,I174683,);
DFFARX1 I_10126 (I174683,I2507,I174657,I174700,);
not I_10127 (I174649,I174700);
not I_10128 (I174722,I174683);
DFFARX1 I_10129 (I575236,I2507,I174657,I174748,);
not I_10130 (I174756,I174748);
and I_10131 (I174773,I174722,I575254);
not I_10132 (I174790,I575251);
nand I_10133 (I174807,I174790,I575254);
not I_10134 (I174824,I575230);
nor I_10135 (I174841,I174824,I575233);
nand I_10136 (I174858,I174841,I575242);
nor I_10137 (I174875,I174858,I174807);
DFFARX1 I_10138 (I174875,I2507,I174657,I174625,);
not I_10139 (I174906,I174858);
not I_10140 (I174923,I575233);
nand I_10141 (I174940,I174923,I575254);
nor I_10142 (I174957,I575233,I575251);
nand I_10143 (I174637,I174773,I174957);
nand I_10144 (I174631,I174722,I575233);
nand I_10145 (I175002,I174824,I575248);
DFFARX1 I_10146 (I175002,I2507,I174657,I174646,);
DFFARX1 I_10147 (I175002,I2507,I174657,I174640,);
not I_10148 (I175047,I575248);
nor I_10149 (I175064,I175047,I575230);
and I_10150 (I175081,I175064,I575239);
or I_10151 (I175098,I175081,I575233);
DFFARX1 I_10152 (I175098,I2507,I174657,I175124,);
nand I_10153 (I175132,I175124,I174790);
nor I_10154 (I174634,I175132,I174940);
nor I_10155 (I174628,I175124,I174756);
DFFARX1 I_10156 (I175124,I2507,I174657,I175186,);
not I_10157 (I175194,I175186);
nor I_10158 (I174643,I175194,I174906);
not I_10159 (I175252,I2514);
DFFARX1 I_10160 (I521471,I2507,I175252,I175278,);
DFFARX1 I_10161 (I175278,I2507,I175252,I175295,);
not I_10162 (I175244,I175295);
not I_10163 (I175317,I175278);
DFFARX1 I_10164 (I521465,I2507,I175252,I175343,);
not I_10165 (I175351,I175343);
and I_10166 (I175368,I175317,I521480);
not I_10167 (I175385,I521477);
nand I_10168 (I175402,I175385,I521480);
not I_10169 (I175419,I521468);
nor I_10170 (I175436,I175419,I521459);
nand I_10171 (I175453,I175436,I521462);
nor I_10172 (I175470,I175453,I175402);
DFFARX1 I_10173 (I175470,I2507,I175252,I175220,);
not I_10174 (I175501,I175453);
not I_10175 (I175518,I521459);
nand I_10176 (I175535,I175518,I521480);
nor I_10177 (I175552,I521459,I521477);
nand I_10178 (I175232,I175368,I175552);
nand I_10179 (I175226,I175317,I521459);
nand I_10180 (I175597,I175419,I521483);
DFFARX1 I_10181 (I175597,I2507,I175252,I175241,);
DFFARX1 I_10182 (I175597,I2507,I175252,I175235,);
not I_10183 (I175642,I521483);
nor I_10184 (I175659,I175642,I521474);
and I_10185 (I175676,I175659,I521459);
or I_10186 (I175693,I175676,I521462);
DFFARX1 I_10187 (I175693,I2507,I175252,I175719,);
nand I_10188 (I175727,I175719,I175385);
nor I_10189 (I175229,I175727,I175535);
nor I_10190 (I175223,I175719,I175351);
DFFARX1 I_10191 (I175719,I2507,I175252,I175781,);
not I_10192 (I175789,I175781);
nor I_10193 (I175238,I175789,I175501);
not I_10194 (I175847,I2514);
DFFARX1 I_10195 (I607035,I2507,I175847,I175873,);
DFFARX1 I_10196 (I175873,I2507,I175847,I175890,);
not I_10197 (I175839,I175890);
not I_10198 (I175912,I175873);
DFFARX1 I_10199 (I607026,I2507,I175847,I175938,);
not I_10200 (I175946,I175938);
and I_10201 (I175963,I175912,I607044);
not I_10202 (I175980,I607041);
nand I_10203 (I175997,I175980,I607044);
not I_10204 (I176014,I607020);
nor I_10205 (I176031,I176014,I607023);
nand I_10206 (I176048,I176031,I607032);
nor I_10207 (I176065,I176048,I175997);
DFFARX1 I_10208 (I176065,I2507,I175847,I175815,);
not I_10209 (I176096,I176048);
not I_10210 (I176113,I607023);
nand I_10211 (I176130,I176113,I607044);
nor I_10212 (I176147,I607023,I607041);
nand I_10213 (I175827,I175963,I176147);
nand I_10214 (I175821,I175912,I607023);
nand I_10215 (I176192,I176014,I607038);
DFFARX1 I_10216 (I176192,I2507,I175847,I175836,);
DFFARX1 I_10217 (I176192,I2507,I175847,I175830,);
not I_10218 (I176237,I607038);
nor I_10219 (I176254,I176237,I607020);
and I_10220 (I176271,I176254,I607029);
or I_10221 (I176288,I176271,I607023);
DFFARX1 I_10222 (I176288,I2507,I175847,I176314,);
nand I_10223 (I176322,I176314,I175980);
nor I_10224 (I175824,I176322,I176130);
nor I_10225 (I175818,I176314,I175946);
DFFARX1 I_10226 (I176314,I2507,I175847,I176376,);
not I_10227 (I176384,I176376);
nor I_10228 (I175833,I176384,I176096);
not I_10229 (I176442,I2514);
DFFARX1 I_10230 (I1314853,I2507,I176442,I176468,);
DFFARX1 I_10231 (I176468,I2507,I176442,I176485,);
not I_10232 (I176434,I176485);
not I_10233 (I176507,I176468);
DFFARX1 I_10234 (I1314844,I2507,I176442,I176533,);
not I_10235 (I176541,I176533);
and I_10236 (I176558,I176507,I1314838);
not I_10237 (I176575,I1314832);
nand I_10238 (I176592,I176575,I1314838);
not I_10239 (I176609,I1314859);
nor I_10240 (I176626,I176609,I1314832);
nand I_10241 (I176643,I176626,I1314856);
nor I_10242 (I176660,I176643,I176592);
DFFARX1 I_10243 (I176660,I2507,I176442,I176410,);
not I_10244 (I176691,I176643);
not I_10245 (I176708,I1314832);
nand I_10246 (I176725,I176708,I1314838);
nor I_10247 (I176742,I1314832,I1314832);
nand I_10248 (I176422,I176558,I176742);
nand I_10249 (I176416,I176507,I1314832);
nand I_10250 (I176787,I176609,I1314841);
DFFARX1 I_10251 (I176787,I2507,I176442,I176431,);
DFFARX1 I_10252 (I176787,I2507,I176442,I176425,);
not I_10253 (I176832,I1314841);
nor I_10254 (I176849,I176832,I1314847);
and I_10255 (I176866,I176849,I1314850);
or I_10256 (I176883,I176866,I1314835);
DFFARX1 I_10257 (I176883,I2507,I176442,I176909,);
nand I_10258 (I176917,I176909,I176575);
nor I_10259 (I176419,I176917,I176725);
nor I_10260 (I176413,I176909,I176541);
DFFARX1 I_10261 (I176909,I2507,I176442,I176971,);
not I_10262 (I176979,I176971);
nor I_10263 (I176428,I176979,I176691);
not I_10264 (I177037,I2514);
DFFARX1 I_10265 (I519686,I2507,I177037,I177063,);
DFFARX1 I_10266 (I177063,I2507,I177037,I177080,);
not I_10267 (I177029,I177080);
not I_10268 (I177102,I177063);
DFFARX1 I_10269 (I519680,I2507,I177037,I177128,);
not I_10270 (I177136,I177128);
and I_10271 (I177153,I177102,I519695);
not I_10272 (I177170,I519692);
nand I_10273 (I177187,I177170,I519695);
not I_10274 (I177204,I519683);
nor I_10275 (I177221,I177204,I519674);
nand I_10276 (I177238,I177221,I519677);
nor I_10277 (I177255,I177238,I177187);
DFFARX1 I_10278 (I177255,I2507,I177037,I177005,);
not I_10279 (I177286,I177238);
not I_10280 (I177303,I519674);
nand I_10281 (I177320,I177303,I519695);
nor I_10282 (I177337,I519674,I519692);
nand I_10283 (I177017,I177153,I177337);
nand I_10284 (I177011,I177102,I519674);
nand I_10285 (I177382,I177204,I519698);
DFFARX1 I_10286 (I177382,I2507,I177037,I177026,);
DFFARX1 I_10287 (I177382,I2507,I177037,I177020,);
not I_10288 (I177427,I519698);
nor I_10289 (I177444,I177427,I519689);
and I_10290 (I177461,I177444,I519674);
or I_10291 (I177478,I177461,I519677);
DFFARX1 I_10292 (I177478,I2507,I177037,I177504,);
nand I_10293 (I177512,I177504,I177170);
nor I_10294 (I177014,I177512,I177320);
nor I_10295 (I177008,I177504,I177136);
DFFARX1 I_10296 (I177504,I2507,I177037,I177566,);
not I_10297 (I177574,I177566);
nor I_10298 (I177023,I177574,I177286);
not I_10299 (I177632,I2514);
DFFARX1 I_10300 (I687952,I2507,I177632,I177658,);
DFFARX1 I_10301 (I177658,I2507,I177632,I177675,);
not I_10302 (I177624,I177675);
not I_10303 (I177697,I177658);
DFFARX1 I_10304 (I687949,I2507,I177632,I177723,);
not I_10305 (I177731,I177723);
and I_10306 (I177748,I177697,I687955);
not I_10307 (I177765,I687940);
nand I_10308 (I177782,I177765,I687955);
not I_10309 (I177799,I687943);
nor I_10310 (I177816,I177799,I687964);
nand I_10311 (I177833,I177816,I687961);
nor I_10312 (I177850,I177833,I177782);
DFFARX1 I_10313 (I177850,I2507,I177632,I177600,);
not I_10314 (I177881,I177833);
not I_10315 (I177898,I687964);
nand I_10316 (I177915,I177898,I687955);
nor I_10317 (I177932,I687964,I687940);
nand I_10318 (I177612,I177748,I177932);
nand I_10319 (I177606,I177697,I687964);
nand I_10320 (I177977,I177799,I687940);
DFFARX1 I_10321 (I177977,I2507,I177632,I177621,);
DFFARX1 I_10322 (I177977,I2507,I177632,I177615,);
not I_10323 (I178022,I687940);
nor I_10324 (I178039,I178022,I687946);
and I_10325 (I178056,I178039,I687958);
or I_10326 (I178073,I178056,I687943);
DFFARX1 I_10327 (I178073,I2507,I177632,I178099,);
nand I_10328 (I178107,I178099,I177765);
nor I_10329 (I177609,I178107,I177915);
nor I_10330 (I177603,I178099,I177731);
DFFARX1 I_10331 (I178099,I2507,I177632,I178161,);
not I_10332 (I178169,I178161);
nor I_10333 (I177618,I178169,I177881);
not I_10334 (I178227,I2514);
DFFARX1 I_10335 (I1051658,I2507,I178227,I178253,);
DFFARX1 I_10336 (I178253,I2507,I178227,I178270,);
not I_10337 (I178219,I178270);
not I_10338 (I178292,I178253);
DFFARX1 I_10339 (I1051667,I2507,I178227,I178318,);
not I_10340 (I178326,I178318);
and I_10341 (I178343,I178292,I1051661);
not I_10342 (I178360,I1051655);
nand I_10343 (I178377,I178360,I1051661);
not I_10344 (I178394,I1051670);
nor I_10345 (I178411,I178394,I1051658);
nand I_10346 (I178428,I178411,I1051664);
nor I_10347 (I178445,I178428,I178377);
DFFARX1 I_10348 (I178445,I2507,I178227,I178195,);
not I_10349 (I178476,I178428);
not I_10350 (I178493,I1051658);
nand I_10351 (I178510,I178493,I1051661);
nor I_10352 (I178527,I1051658,I1051655);
nand I_10353 (I178207,I178343,I178527);
nand I_10354 (I178201,I178292,I1051658);
nand I_10355 (I178572,I178394,I1051661);
DFFARX1 I_10356 (I178572,I2507,I178227,I178216,);
DFFARX1 I_10357 (I178572,I2507,I178227,I178210,);
not I_10358 (I178617,I1051661);
nor I_10359 (I178634,I178617,I1051676);
and I_10360 (I178651,I178634,I1051673);
or I_10361 (I178668,I178651,I1051655);
DFFARX1 I_10362 (I178668,I2507,I178227,I178694,);
nand I_10363 (I178702,I178694,I178360);
nor I_10364 (I178204,I178702,I178510);
nor I_10365 (I178198,I178694,I178326);
DFFARX1 I_10366 (I178694,I2507,I178227,I178756,);
not I_10367 (I178764,I178756);
nor I_10368 (I178213,I178764,I178476);
not I_10369 (I178822,I2514);
DFFARX1 I_10370 (I976734,I2507,I178822,I178848,);
DFFARX1 I_10371 (I178848,I2507,I178822,I178865,);
not I_10372 (I178814,I178865);
not I_10373 (I178887,I178848);
DFFARX1 I_10374 (I976743,I2507,I178822,I178913,);
not I_10375 (I178921,I178913);
and I_10376 (I178938,I178887,I976731);
not I_10377 (I178955,I976722);
nand I_10378 (I178972,I178955,I976731);
not I_10379 (I178989,I976728);
nor I_10380 (I179006,I178989,I976746);
nand I_10381 (I179023,I179006,I976719);
nor I_10382 (I179040,I179023,I178972);
DFFARX1 I_10383 (I179040,I2507,I178822,I178790,);
not I_10384 (I179071,I179023);
not I_10385 (I179088,I976746);
nand I_10386 (I179105,I179088,I976731);
nor I_10387 (I179122,I976746,I976722);
nand I_10388 (I178802,I178938,I179122);
nand I_10389 (I178796,I178887,I976746);
nand I_10390 (I179167,I178989,I976725);
DFFARX1 I_10391 (I179167,I2507,I178822,I178811,);
DFFARX1 I_10392 (I179167,I2507,I178822,I178805,);
not I_10393 (I179212,I976725);
nor I_10394 (I179229,I179212,I976737);
and I_10395 (I179246,I179229,I976719);
or I_10396 (I179263,I179246,I976740);
DFFARX1 I_10397 (I179263,I2507,I178822,I179289,);
nand I_10398 (I179297,I179289,I178955);
nor I_10399 (I178799,I179297,I179105);
nor I_10400 (I178793,I179289,I178921);
DFFARX1 I_10401 (I179289,I2507,I178822,I179351,);
not I_10402 (I179359,I179351);
nor I_10403 (I178808,I179359,I179071);
not I_10404 (I179417,I2514);
DFFARX1 I_10405 (I842833,I2507,I179417,I179443,);
DFFARX1 I_10406 (I179443,I2507,I179417,I179460,);
not I_10407 (I179409,I179460);
not I_10408 (I179482,I179443);
DFFARX1 I_10409 (I842827,I2507,I179417,I179508,);
not I_10410 (I179516,I179508);
and I_10411 (I179533,I179482,I842845);
not I_10412 (I179550,I842833);
nand I_10413 (I179567,I179550,I842845);
not I_10414 (I179584,I842827);
nor I_10415 (I179601,I179584,I842839);
nand I_10416 (I179618,I179601,I842830);
nor I_10417 (I179635,I179618,I179567);
DFFARX1 I_10418 (I179635,I2507,I179417,I179385,);
not I_10419 (I179666,I179618);
not I_10420 (I179683,I842839);
nand I_10421 (I179700,I179683,I842845);
nor I_10422 (I179717,I842839,I842833);
nand I_10423 (I179397,I179533,I179717);
nand I_10424 (I179391,I179482,I842839);
nand I_10425 (I179762,I179584,I842842);
DFFARX1 I_10426 (I179762,I2507,I179417,I179406,);
DFFARX1 I_10427 (I179762,I2507,I179417,I179400,);
not I_10428 (I179807,I842842);
nor I_10429 (I179824,I179807,I842848);
and I_10430 (I179841,I179824,I842830);
or I_10431 (I179858,I179841,I842836);
DFFARX1 I_10432 (I179858,I2507,I179417,I179884,);
nand I_10433 (I179892,I179884,I179550);
nor I_10434 (I179394,I179892,I179700);
nor I_10435 (I179388,I179884,I179516);
DFFARX1 I_10436 (I179884,I2507,I179417,I179946,);
not I_10437 (I179954,I179946);
nor I_10438 (I179403,I179954,I179666);
not I_10439 (I180012,I2514);
DFFARX1 I_10440 (I61720,I2507,I180012,I180038,);
DFFARX1 I_10441 (I180038,I2507,I180012,I180055,);
not I_10442 (I180004,I180055);
not I_10443 (I180077,I180038);
DFFARX1 I_10444 (I61714,I2507,I180012,I180103,);
not I_10445 (I180111,I180103);
and I_10446 (I180128,I180077,I61711);
not I_10447 (I180145,I61732);
nand I_10448 (I180162,I180145,I61711);
not I_10449 (I180179,I61726);
nor I_10450 (I180196,I180179,I61717);
nand I_10451 (I180213,I180196,I61723);
nor I_10452 (I180230,I180213,I180162);
DFFARX1 I_10453 (I180230,I2507,I180012,I179980,);
not I_10454 (I180261,I180213);
not I_10455 (I180278,I61717);
nand I_10456 (I180295,I180278,I61711);
nor I_10457 (I180312,I61717,I61732);
nand I_10458 (I179992,I180128,I180312);
nand I_10459 (I179986,I180077,I61717);
nand I_10460 (I180357,I180179,I61711);
DFFARX1 I_10461 (I180357,I2507,I180012,I180001,);
DFFARX1 I_10462 (I180357,I2507,I180012,I179995,);
not I_10463 (I180402,I61711);
nor I_10464 (I180419,I180402,I61729);
and I_10465 (I180436,I180419,I61735);
or I_10466 (I180453,I180436,I61714);
DFFARX1 I_10467 (I180453,I2507,I180012,I180479,);
nand I_10468 (I180487,I180479,I180145);
nor I_10469 (I179989,I180487,I180295);
nor I_10470 (I179983,I180479,I180111);
DFFARX1 I_10471 (I180479,I2507,I180012,I180541,);
not I_10472 (I180549,I180541);
nor I_10473 (I179998,I180549,I180261);
not I_10474 (I180607,I2514);
DFFARX1 I_10475 (I686796,I2507,I180607,I180633,);
DFFARX1 I_10476 (I180633,I2507,I180607,I180650,);
not I_10477 (I180599,I180650);
not I_10478 (I180672,I180633);
DFFARX1 I_10479 (I686793,I2507,I180607,I180698,);
not I_10480 (I180706,I180698);
and I_10481 (I180723,I180672,I686799);
not I_10482 (I180740,I686784);
nand I_10483 (I180757,I180740,I686799);
not I_10484 (I180774,I686787);
nor I_10485 (I180791,I180774,I686808);
nand I_10486 (I180808,I180791,I686805);
nor I_10487 (I180825,I180808,I180757);
DFFARX1 I_10488 (I180825,I2507,I180607,I180575,);
not I_10489 (I180856,I180808);
not I_10490 (I180873,I686808);
nand I_10491 (I180890,I180873,I686799);
nor I_10492 (I180907,I686808,I686784);
nand I_10493 (I180587,I180723,I180907);
nand I_10494 (I180581,I180672,I686808);
nand I_10495 (I180952,I180774,I686784);
DFFARX1 I_10496 (I180952,I2507,I180607,I180596,);
DFFARX1 I_10497 (I180952,I2507,I180607,I180590,);
not I_10498 (I180997,I686784);
nor I_10499 (I181014,I180997,I686790);
and I_10500 (I181031,I181014,I686802);
or I_10501 (I181048,I181031,I686787);
DFFARX1 I_10502 (I181048,I2507,I180607,I181074,);
nand I_10503 (I181082,I181074,I180740);
nor I_10504 (I180584,I181082,I180890);
nor I_10505 (I180578,I181074,I180706);
DFFARX1 I_10506 (I181074,I2507,I180607,I181136,);
not I_10507 (I181144,I181136);
nor I_10508 (I180593,I181144,I180856);
not I_10509 (I181202,I2514);
DFFARX1 I_10510 (I414791,I2507,I181202,I181228,);
DFFARX1 I_10511 (I181228,I2507,I181202,I181245,);
not I_10512 (I181194,I181245);
not I_10513 (I181267,I181228);
DFFARX1 I_10514 (I414779,I2507,I181202,I181293,);
not I_10515 (I181301,I181293);
and I_10516 (I181318,I181267,I414788);
not I_10517 (I181335,I414785);
nand I_10518 (I181352,I181335,I414788);
not I_10519 (I181369,I414776);
nor I_10520 (I181386,I181369,I414782);
nand I_10521 (I181403,I181386,I414767);
nor I_10522 (I181420,I181403,I181352);
DFFARX1 I_10523 (I181420,I2507,I181202,I181170,);
not I_10524 (I181451,I181403);
not I_10525 (I181468,I414782);
nand I_10526 (I181485,I181468,I414788);
nor I_10527 (I181502,I414782,I414785);
nand I_10528 (I181182,I181318,I181502);
nand I_10529 (I181176,I181267,I414782);
nand I_10530 (I181547,I181369,I414767);
DFFARX1 I_10531 (I181547,I2507,I181202,I181191,);
DFFARX1 I_10532 (I181547,I2507,I181202,I181185,);
not I_10533 (I181592,I414767);
nor I_10534 (I181609,I181592,I414773);
and I_10535 (I181626,I181609,I414770);
or I_10536 (I181643,I181626,I414794);
DFFARX1 I_10537 (I181643,I2507,I181202,I181669,);
nand I_10538 (I181677,I181669,I181335);
nor I_10539 (I181179,I181677,I181485);
nor I_10540 (I181173,I181669,I181301);
DFFARX1 I_10541 (I181669,I2507,I181202,I181731,);
not I_10542 (I181739,I181731);
nor I_10543 (I181188,I181739,I181451);
not I_10544 (I181797,I2514);
DFFARX1 I_10545 (I310268,I2507,I181797,I181823,);
DFFARX1 I_10546 (I181823,I2507,I181797,I181840,);
not I_10547 (I181789,I181840);
not I_10548 (I181862,I181823);
DFFARX1 I_10549 (I310283,I2507,I181797,I181888,);
not I_10550 (I181896,I181888);
and I_10551 (I181913,I181862,I310280);
not I_10552 (I181930,I310268);
nand I_10553 (I181947,I181930,I310280);
not I_10554 (I181964,I310277);
nor I_10555 (I181981,I181964,I310292);
nand I_10556 (I181998,I181981,I310289);
nor I_10557 (I182015,I181998,I181947);
DFFARX1 I_10558 (I182015,I2507,I181797,I181765,);
not I_10559 (I182046,I181998);
not I_10560 (I182063,I310292);
nand I_10561 (I182080,I182063,I310280);
nor I_10562 (I182097,I310292,I310268);
nand I_10563 (I181777,I181913,I182097);
nand I_10564 (I181771,I181862,I310292);
nand I_10565 (I182142,I181964,I310286);
DFFARX1 I_10566 (I182142,I2507,I181797,I181786,);
DFFARX1 I_10567 (I182142,I2507,I181797,I181780,);
not I_10568 (I182187,I310286);
nor I_10569 (I182204,I182187,I310274);
and I_10570 (I182221,I182204,I310295);
or I_10571 (I182238,I182221,I310271);
DFFARX1 I_10572 (I182238,I2507,I181797,I182264,);
nand I_10573 (I182272,I182264,I181930);
nor I_10574 (I181774,I182272,I182080);
nor I_10575 (I181768,I182264,I181896);
DFFARX1 I_10576 (I182264,I2507,I181797,I182326,);
not I_10577 (I182334,I182326);
nor I_10578 (I181783,I182334,I182046);
not I_10579 (I182392,I2514);
DFFARX1 I_10580 (I1121950,I2507,I182392,I182418,);
DFFARX1 I_10581 (I182418,I2507,I182392,I182435,);
not I_10582 (I182384,I182435);
not I_10583 (I182457,I182418);
DFFARX1 I_10584 (I1121950,I2507,I182392,I182483,);
not I_10585 (I182491,I182483);
and I_10586 (I182508,I182457,I1121953);
not I_10587 (I182525,I1121965);
nand I_10588 (I182542,I182525,I1121953);
not I_10589 (I182559,I1121971);
nor I_10590 (I182576,I182559,I1121962);
nand I_10591 (I182593,I182576,I1121968);
nor I_10592 (I182610,I182593,I182542);
DFFARX1 I_10593 (I182610,I2507,I182392,I182360,);
not I_10594 (I182641,I182593);
not I_10595 (I182658,I1121962);
nand I_10596 (I182675,I182658,I1121953);
nor I_10597 (I182692,I1121962,I1121965);
nand I_10598 (I182372,I182508,I182692);
nand I_10599 (I182366,I182457,I1121962);
nand I_10600 (I182737,I182559,I1121959);
DFFARX1 I_10601 (I182737,I2507,I182392,I182381,);
DFFARX1 I_10602 (I182737,I2507,I182392,I182375,);
not I_10603 (I182782,I1121959);
nor I_10604 (I182799,I182782,I1121956);
and I_10605 (I182816,I182799,I1121974);
or I_10606 (I182833,I182816,I1121953);
DFFARX1 I_10607 (I182833,I2507,I182392,I182859,);
nand I_10608 (I182867,I182859,I182525);
nor I_10609 (I182369,I182867,I182675);
nor I_10610 (I182363,I182859,I182491);
DFFARX1 I_10611 (I182859,I2507,I182392,I182921,);
not I_10612 (I182929,I182921);
nor I_10613 (I182378,I182929,I182641);
not I_10614 (I182987,I2514);
DFFARX1 I_10615 (I668878,I2507,I182987,I183013,);
DFFARX1 I_10616 (I183013,I2507,I182987,I183030,);
not I_10617 (I182979,I183030);
not I_10618 (I183052,I183013);
DFFARX1 I_10619 (I668875,I2507,I182987,I183078,);
not I_10620 (I183086,I183078);
and I_10621 (I183103,I183052,I668881);
not I_10622 (I183120,I668866);
nand I_10623 (I183137,I183120,I668881);
not I_10624 (I183154,I668869);
nor I_10625 (I183171,I183154,I668890);
nand I_10626 (I183188,I183171,I668887);
nor I_10627 (I183205,I183188,I183137);
DFFARX1 I_10628 (I183205,I2507,I182987,I182955,);
not I_10629 (I183236,I183188);
not I_10630 (I183253,I668890);
nand I_10631 (I183270,I183253,I668881);
nor I_10632 (I183287,I668890,I668866);
nand I_10633 (I182967,I183103,I183287);
nand I_10634 (I182961,I183052,I668890);
nand I_10635 (I183332,I183154,I668866);
DFFARX1 I_10636 (I183332,I2507,I182987,I182976,);
DFFARX1 I_10637 (I183332,I2507,I182987,I182970,);
not I_10638 (I183377,I668866);
nor I_10639 (I183394,I183377,I668872);
and I_10640 (I183411,I183394,I668884);
or I_10641 (I183428,I183411,I668869);
DFFARX1 I_10642 (I183428,I2507,I182987,I183454,);
nand I_10643 (I183462,I183454,I183120);
nor I_10644 (I182964,I183462,I183270);
nor I_10645 (I182958,I183454,I183086);
DFFARX1 I_10646 (I183454,I2507,I182987,I183516,);
not I_10647 (I183524,I183516);
nor I_10648 (I182973,I183524,I183236);
not I_10649 (I183582,I2514);
DFFARX1 I_10650 (I1168768,I2507,I183582,I183608,);
DFFARX1 I_10651 (I183608,I2507,I183582,I183625,);
not I_10652 (I183574,I183625);
not I_10653 (I183647,I183608);
DFFARX1 I_10654 (I1168768,I2507,I183582,I183673,);
not I_10655 (I183681,I183673);
and I_10656 (I183698,I183647,I1168771);
not I_10657 (I183715,I1168783);
nand I_10658 (I183732,I183715,I1168771);
not I_10659 (I183749,I1168789);
nor I_10660 (I183766,I183749,I1168780);
nand I_10661 (I183783,I183766,I1168786);
nor I_10662 (I183800,I183783,I183732);
DFFARX1 I_10663 (I183800,I2507,I183582,I183550,);
not I_10664 (I183831,I183783);
not I_10665 (I183848,I1168780);
nand I_10666 (I183865,I183848,I1168771);
nor I_10667 (I183882,I1168780,I1168783);
nand I_10668 (I183562,I183698,I183882);
nand I_10669 (I183556,I183647,I1168780);
nand I_10670 (I183927,I183749,I1168777);
DFFARX1 I_10671 (I183927,I2507,I183582,I183571,);
DFFARX1 I_10672 (I183927,I2507,I183582,I183565,);
not I_10673 (I183972,I1168777);
nor I_10674 (I183989,I183972,I1168774);
and I_10675 (I184006,I183989,I1168792);
or I_10676 (I184023,I184006,I1168771);
DFFARX1 I_10677 (I184023,I2507,I183582,I184049,);
nand I_10678 (I184057,I184049,I183715);
nor I_10679 (I183559,I184057,I183865);
nor I_10680 (I183553,I184049,I183681);
DFFARX1 I_10681 (I184049,I2507,I183582,I184111,);
not I_10682 (I184119,I184111);
nor I_10683 (I183568,I184119,I183831);
not I_10684 (I184177,I2514);
DFFARX1 I_10685 (I91232,I2507,I184177,I184203,);
DFFARX1 I_10686 (I184203,I2507,I184177,I184220,);
not I_10687 (I184169,I184220);
not I_10688 (I184242,I184203);
DFFARX1 I_10689 (I91226,I2507,I184177,I184268,);
not I_10690 (I184276,I184268);
and I_10691 (I184293,I184242,I91223);
not I_10692 (I184310,I91244);
nand I_10693 (I184327,I184310,I91223);
not I_10694 (I184344,I91238);
nor I_10695 (I184361,I184344,I91229);
nand I_10696 (I184378,I184361,I91235);
nor I_10697 (I184395,I184378,I184327);
DFFARX1 I_10698 (I184395,I2507,I184177,I184145,);
not I_10699 (I184426,I184378);
not I_10700 (I184443,I91229);
nand I_10701 (I184460,I184443,I91223);
nor I_10702 (I184477,I91229,I91244);
nand I_10703 (I184157,I184293,I184477);
nand I_10704 (I184151,I184242,I91229);
nand I_10705 (I184522,I184344,I91223);
DFFARX1 I_10706 (I184522,I2507,I184177,I184166,);
DFFARX1 I_10707 (I184522,I2507,I184177,I184160,);
not I_10708 (I184567,I91223);
nor I_10709 (I184584,I184567,I91241);
and I_10710 (I184601,I184584,I91247);
or I_10711 (I184618,I184601,I91226);
DFFARX1 I_10712 (I184618,I2507,I184177,I184644,);
nand I_10713 (I184652,I184644,I184310);
nor I_10714 (I184154,I184652,I184460);
nor I_10715 (I184148,I184644,I184276);
DFFARX1 I_10716 (I184644,I2507,I184177,I184706,);
not I_10717 (I184714,I184706);
nor I_10718 (I184163,I184714,I184426);
not I_10719 (I184772,I2514);
DFFARX1 I_10720 (I280229,I2507,I184772,I184798,);
DFFARX1 I_10721 (I184798,I2507,I184772,I184815,);
not I_10722 (I184764,I184815);
not I_10723 (I184837,I184798);
DFFARX1 I_10724 (I280244,I2507,I184772,I184863,);
not I_10725 (I184871,I184863);
and I_10726 (I184888,I184837,I280241);
not I_10727 (I184905,I280229);
nand I_10728 (I184922,I184905,I280241);
not I_10729 (I184939,I280238);
nor I_10730 (I184956,I184939,I280253);
nand I_10731 (I184973,I184956,I280250);
nor I_10732 (I184990,I184973,I184922);
DFFARX1 I_10733 (I184990,I2507,I184772,I184740,);
not I_10734 (I185021,I184973);
not I_10735 (I185038,I280253);
nand I_10736 (I185055,I185038,I280241);
nor I_10737 (I185072,I280253,I280229);
nand I_10738 (I184752,I184888,I185072);
nand I_10739 (I184746,I184837,I280253);
nand I_10740 (I185117,I184939,I280247);
DFFARX1 I_10741 (I185117,I2507,I184772,I184761,);
DFFARX1 I_10742 (I185117,I2507,I184772,I184755,);
not I_10743 (I185162,I280247);
nor I_10744 (I185179,I185162,I280235);
and I_10745 (I185196,I185179,I280256);
or I_10746 (I185213,I185196,I280232);
DFFARX1 I_10747 (I185213,I2507,I184772,I185239,);
nand I_10748 (I185247,I185239,I184905);
nor I_10749 (I184749,I185247,I185055);
nor I_10750 (I184743,I185239,I184871);
DFFARX1 I_10751 (I185239,I2507,I184772,I185301,);
not I_10752 (I185309,I185301);
nor I_10753 (I184758,I185309,I185021);
not I_10754 (I185367,I2514);
DFFARX1 I_10755 (I46452,I2507,I185367,I185393,);
DFFARX1 I_10756 (I185393,I2507,I185367,I185410,);
not I_10757 (I185359,I185410);
not I_10758 (I185432,I185393);
DFFARX1 I_10759 (I46428,I2507,I185367,I185458,);
not I_10760 (I185466,I185458);
and I_10761 (I185483,I185432,I46443);
not I_10762 (I185500,I46431);
nand I_10763 (I185517,I185500,I46443);
not I_10764 (I185534,I46434);
nor I_10765 (I185551,I185534,I46446);
nand I_10766 (I185568,I185551,I46437);
nor I_10767 (I185585,I185568,I185517);
DFFARX1 I_10768 (I185585,I2507,I185367,I185335,);
not I_10769 (I185616,I185568);
not I_10770 (I185633,I46446);
nand I_10771 (I185650,I185633,I46443);
nor I_10772 (I185667,I46446,I46431);
nand I_10773 (I185347,I185483,I185667);
nand I_10774 (I185341,I185432,I46446);
nand I_10775 (I185712,I185534,I46440);
DFFARX1 I_10776 (I185712,I2507,I185367,I185356,);
DFFARX1 I_10777 (I185712,I2507,I185367,I185350,);
not I_10778 (I185757,I46440);
nor I_10779 (I185774,I185757,I46431);
and I_10780 (I185791,I185774,I46428);
or I_10781 (I185808,I185791,I46449);
DFFARX1 I_10782 (I185808,I2507,I185367,I185834,);
nand I_10783 (I185842,I185834,I185500);
nor I_10784 (I185344,I185842,I185650);
nor I_10785 (I185338,I185834,I185466);
DFFARX1 I_10786 (I185834,I2507,I185367,I185896,);
not I_10787 (I185904,I185896);
nor I_10788 (I185353,I185904,I185616);
not I_10789 (I185962,I2514);
DFFARX1 I_10790 (I316065,I2507,I185962,I185988,);
DFFARX1 I_10791 (I185988,I2507,I185962,I186005,);
not I_10792 (I185954,I186005);
not I_10793 (I186027,I185988);
DFFARX1 I_10794 (I316080,I2507,I185962,I186053,);
not I_10795 (I186061,I186053);
and I_10796 (I186078,I186027,I316077);
not I_10797 (I186095,I316065);
nand I_10798 (I186112,I186095,I316077);
not I_10799 (I186129,I316074);
nor I_10800 (I186146,I186129,I316089);
nand I_10801 (I186163,I186146,I316086);
nor I_10802 (I186180,I186163,I186112);
DFFARX1 I_10803 (I186180,I2507,I185962,I185930,);
not I_10804 (I186211,I186163);
not I_10805 (I186228,I316089);
nand I_10806 (I186245,I186228,I316077);
nor I_10807 (I186262,I316089,I316065);
nand I_10808 (I185942,I186078,I186262);
nand I_10809 (I185936,I186027,I316089);
nand I_10810 (I186307,I186129,I316083);
DFFARX1 I_10811 (I186307,I2507,I185962,I185951,);
DFFARX1 I_10812 (I186307,I2507,I185962,I185945,);
not I_10813 (I186352,I316083);
nor I_10814 (I186369,I186352,I316071);
and I_10815 (I186386,I186369,I316092);
or I_10816 (I186403,I186386,I316068);
DFFARX1 I_10817 (I186403,I2507,I185962,I186429,);
nand I_10818 (I186437,I186429,I186095);
nor I_10819 (I185939,I186437,I186245);
nor I_10820 (I185933,I186429,I186061);
DFFARX1 I_10821 (I186429,I2507,I185962,I186491,);
not I_10822 (I186499,I186491);
nor I_10823 (I185948,I186499,I186211);
not I_10824 (I186557,I2514);
DFFARX1 I_10825 (I1301446,I2507,I186557,I186583,);
DFFARX1 I_10826 (I186583,I2507,I186557,I186600,);
not I_10827 (I186549,I186600);
not I_10828 (I186622,I186583);
DFFARX1 I_10829 (I1301419,I2507,I186557,I186648,);
not I_10830 (I186656,I186648);
and I_10831 (I186673,I186622,I1301443);
not I_10832 (I186690,I1301440);
nand I_10833 (I186707,I186690,I1301443);
not I_10834 (I186724,I1301419);
nor I_10835 (I186741,I186724,I1301437);
nand I_10836 (I186758,I186741,I1301425);
nor I_10837 (I186775,I186758,I186707);
DFFARX1 I_10838 (I186775,I2507,I186557,I186525,);
not I_10839 (I186806,I186758);
not I_10840 (I186823,I1301437);
nand I_10841 (I186840,I186823,I1301443);
nor I_10842 (I186857,I1301437,I1301440);
nand I_10843 (I186537,I186673,I186857);
nand I_10844 (I186531,I186622,I1301437);
nand I_10845 (I186902,I186724,I1301431);
DFFARX1 I_10846 (I186902,I2507,I186557,I186546,);
DFFARX1 I_10847 (I186902,I2507,I186557,I186540,);
not I_10848 (I186947,I1301431);
nor I_10849 (I186964,I186947,I1301434);
and I_10850 (I186981,I186964,I1301422);
or I_10851 (I186998,I186981,I1301428);
DFFARX1 I_10852 (I186998,I2507,I186557,I187024,);
nand I_10853 (I187032,I187024,I186690);
nor I_10854 (I186534,I187032,I186840);
nor I_10855 (I186528,I187024,I186656);
DFFARX1 I_10856 (I187024,I2507,I186557,I187086,);
not I_10857 (I187094,I187086);
nor I_10858 (I186543,I187094,I186806);
not I_10859 (I187152,I2514);
DFFARX1 I_10860 (I1321398,I2507,I187152,I187178,);
DFFARX1 I_10861 (I187178,I2507,I187152,I187195,);
not I_10862 (I187144,I187195);
not I_10863 (I187217,I187178);
DFFARX1 I_10864 (I1321389,I2507,I187152,I187243,);
not I_10865 (I187251,I187243);
and I_10866 (I187268,I187217,I1321383);
not I_10867 (I187285,I1321377);
nand I_10868 (I187302,I187285,I1321383);
not I_10869 (I187319,I1321404);
nor I_10870 (I187336,I187319,I1321377);
nand I_10871 (I187353,I187336,I1321401);
nor I_10872 (I187370,I187353,I187302);
DFFARX1 I_10873 (I187370,I2507,I187152,I187120,);
not I_10874 (I187401,I187353);
not I_10875 (I187418,I1321377);
nand I_10876 (I187435,I187418,I1321383);
nor I_10877 (I187452,I1321377,I1321377);
nand I_10878 (I187132,I187268,I187452);
nand I_10879 (I187126,I187217,I1321377);
nand I_10880 (I187497,I187319,I1321386);
DFFARX1 I_10881 (I187497,I2507,I187152,I187141,);
DFFARX1 I_10882 (I187497,I2507,I187152,I187135,);
not I_10883 (I187542,I1321386);
nor I_10884 (I187559,I187542,I1321392);
and I_10885 (I187576,I187559,I1321395);
or I_10886 (I187593,I187576,I1321380);
DFFARX1 I_10887 (I187593,I2507,I187152,I187619,);
nand I_10888 (I187627,I187619,I187285);
nor I_10889 (I187129,I187627,I187435);
nor I_10890 (I187123,I187619,I187251);
DFFARX1 I_10891 (I187619,I2507,I187152,I187681,);
not I_10892 (I187689,I187681);
nor I_10893 (I187138,I187689,I187401);
not I_10894 (I187747,I2514);
DFFARX1 I_10895 (I1065306,I2507,I187747,I187773,);
DFFARX1 I_10896 (I187773,I2507,I187747,I187790,);
not I_10897 (I187739,I187790);
not I_10898 (I187812,I187773);
DFFARX1 I_10899 (I1065306,I2507,I187747,I187838,);
not I_10900 (I187846,I187838);
and I_10901 (I187863,I187812,I1065309);
not I_10902 (I187880,I1065321);
nand I_10903 (I187897,I187880,I1065309);
not I_10904 (I187914,I1065327);
nor I_10905 (I187931,I187914,I1065318);
nand I_10906 (I187948,I187931,I1065324);
nor I_10907 (I187965,I187948,I187897);
DFFARX1 I_10908 (I187965,I2507,I187747,I187715,);
not I_10909 (I187996,I187948);
not I_10910 (I188013,I1065318);
nand I_10911 (I188030,I188013,I1065309);
nor I_10912 (I188047,I1065318,I1065321);
nand I_10913 (I187727,I187863,I188047);
nand I_10914 (I187721,I187812,I1065318);
nand I_10915 (I188092,I187914,I1065315);
DFFARX1 I_10916 (I188092,I2507,I187747,I187736,);
DFFARX1 I_10917 (I188092,I2507,I187747,I187730,);
not I_10918 (I188137,I1065315);
nor I_10919 (I188154,I188137,I1065312);
and I_10920 (I188171,I188154,I1065330);
or I_10921 (I188188,I188171,I1065309);
DFFARX1 I_10922 (I188188,I2507,I187747,I188214,);
nand I_10923 (I188222,I188214,I187880);
nor I_10924 (I187724,I188222,I188030);
nor I_10925 (I187718,I188214,I187846);
DFFARX1 I_10926 (I188214,I2507,I187747,I188276,);
not I_10927 (I188284,I188276);
nor I_10928 (I187733,I188284,I187996);
not I_10929 (I188342,I2514);
DFFARX1 I_10930 (I77003,I2507,I188342,I188368,);
DFFARX1 I_10931 (I188368,I2507,I188342,I188385,);
not I_10932 (I188334,I188385);
not I_10933 (I188407,I188368);
DFFARX1 I_10934 (I76997,I2507,I188342,I188433,);
not I_10935 (I188441,I188433);
and I_10936 (I188458,I188407,I76994);
not I_10937 (I188475,I77015);
nand I_10938 (I188492,I188475,I76994);
not I_10939 (I188509,I77009);
nor I_10940 (I188526,I188509,I77000);
nand I_10941 (I188543,I188526,I77006);
nor I_10942 (I188560,I188543,I188492);
DFFARX1 I_10943 (I188560,I2507,I188342,I188310,);
not I_10944 (I188591,I188543);
not I_10945 (I188608,I77000);
nand I_10946 (I188625,I188608,I76994);
nor I_10947 (I188642,I77000,I77015);
nand I_10948 (I188322,I188458,I188642);
nand I_10949 (I188316,I188407,I77000);
nand I_10950 (I188687,I188509,I76994);
DFFARX1 I_10951 (I188687,I2507,I188342,I188331,);
DFFARX1 I_10952 (I188687,I2507,I188342,I188325,);
not I_10953 (I188732,I76994);
nor I_10954 (I188749,I188732,I77012);
and I_10955 (I188766,I188749,I77018);
or I_10956 (I188783,I188766,I76997);
DFFARX1 I_10957 (I188783,I2507,I188342,I188809,);
nand I_10958 (I188817,I188809,I188475);
nor I_10959 (I188319,I188817,I188625);
nor I_10960 (I188313,I188809,I188441);
DFFARX1 I_10961 (I188809,I2507,I188342,I188871,);
not I_10962 (I188879,I188871);
nor I_10963 (I188328,I188879,I188591);
not I_10964 (I188937,I2514);
DFFARX1 I_10965 (I1043804,I2507,I188937,I188963,);
DFFARX1 I_10966 (I188963,I2507,I188937,I188980,);
not I_10967 (I188929,I188980);
not I_10968 (I189002,I188963);
DFFARX1 I_10969 (I1043813,I2507,I188937,I189028,);
not I_10970 (I189036,I189028);
and I_10971 (I189053,I189002,I1043807);
not I_10972 (I189070,I1043801);
nand I_10973 (I189087,I189070,I1043807);
not I_10974 (I189104,I1043816);
nor I_10975 (I189121,I189104,I1043804);
nand I_10976 (I189138,I189121,I1043810);
nor I_10977 (I189155,I189138,I189087);
DFFARX1 I_10978 (I189155,I2507,I188937,I188905,);
not I_10979 (I189186,I189138);
not I_10980 (I189203,I1043804);
nand I_10981 (I189220,I189203,I1043807);
nor I_10982 (I189237,I1043804,I1043801);
nand I_10983 (I188917,I189053,I189237);
nand I_10984 (I188911,I189002,I1043804);
nand I_10985 (I189282,I189104,I1043807);
DFFARX1 I_10986 (I189282,I2507,I188937,I188926,);
DFFARX1 I_10987 (I189282,I2507,I188937,I188920,);
not I_10988 (I189327,I1043807);
nor I_10989 (I189344,I189327,I1043822);
and I_10990 (I189361,I189344,I1043819);
or I_10991 (I189378,I189361,I1043801);
DFFARX1 I_10992 (I189378,I2507,I188937,I189404,);
nand I_10993 (I189412,I189404,I189070);
nor I_10994 (I188914,I189412,I189220);
nor I_10995 (I188908,I189404,I189036);
DFFARX1 I_10996 (I189404,I2507,I188937,I189466,);
not I_10997 (I189474,I189466);
nor I_10998 (I188923,I189474,I189186);
not I_10999 (I189532,I2514);
DFFARX1 I_11000 (I590273,I2507,I189532,I189558,);
DFFARX1 I_11001 (I189558,I2507,I189532,I189575,);
not I_11002 (I189524,I189575);
not I_11003 (I189597,I189558);
DFFARX1 I_11004 (I590264,I2507,I189532,I189623,);
not I_11005 (I189631,I189623);
and I_11006 (I189648,I189597,I590282);
not I_11007 (I189665,I590279);
nand I_11008 (I189682,I189665,I590282);
not I_11009 (I189699,I590258);
nor I_11010 (I189716,I189699,I590261);
nand I_11011 (I189733,I189716,I590270);
nor I_11012 (I189750,I189733,I189682);
DFFARX1 I_11013 (I189750,I2507,I189532,I189500,);
not I_11014 (I189781,I189733);
not I_11015 (I189798,I590261);
nand I_11016 (I189815,I189798,I590282);
nor I_11017 (I189832,I590261,I590279);
nand I_11018 (I189512,I189648,I189832);
nand I_11019 (I189506,I189597,I590261);
nand I_11020 (I189877,I189699,I590276);
DFFARX1 I_11021 (I189877,I2507,I189532,I189521,);
DFFARX1 I_11022 (I189877,I2507,I189532,I189515,);
not I_11023 (I189922,I590276);
nor I_11024 (I189939,I189922,I590258);
and I_11025 (I189956,I189939,I590267);
or I_11026 (I189973,I189956,I590261);
DFFARX1 I_11027 (I189973,I2507,I189532,I189999,);
nand I_11028 (I190007,I189999,I189665);
nor I_11029 (I189509,I190007,I189815);
nor I_11030 (I189503,I189999,I189631);
DFFARX1 I_11031 (I189999,I2507,I189532,I190061,);
not I_11032 (I190069,I190061);
nor I_11033 (I189518,I190069,I189781);
not I_11034 (I190127,I2514);
DFFARX1 I_11035 (I796457,I2507,I190127,I190153,);
DFFARX1 I_11036 (I190153,I2507,I190127,I190170,);
not I_11037 (I190119,I190170);
not I_11038 (I190192,I190153);
DFFARX1 I_11039 (I796451,I2507,I190127,I190218,);
not I_11040 (I190226,I190218);
and I_11041 (I190243,I190192,I796469);
not I_11042 (I190260,I796457);
nand I_11043 (I190277,I190260,I796469);
not I_11044 (I190294,I796451);
nor I_11045 (I190311,I190294,I796463);
nand I_11046 (I190328,I190311,I796454);
nor I_11047 (I190345,I190328,I190277);
DFFARX1 I_11048 (I190345,I2507,I190127,I190095,);
not I_11049 (I190376,I190328);
not I_11050 (I190393,I796463);
nand I_11051 (I190410,I190393,I796469);
nor I_11052 (I190427,I796463,I796457);
nand I_11053 (I190107,I190243,I190427);
nand I_11054 (I190101,I190192,I796463);
nand I_11055 (I190472,I190294,I796466);
DFFARX1 I_11056 (I190472,I2507,I190127,I190116,);
DFFARX1 I_11057 (I190472,I2507,I190127,I190110,);
not I_11058 (I190517,I796466);
nor I_11059 (I190534,I190517,I796472);
and I_11060 (I190551,I190534,I796454);
or I_11061 (I190568,I190551,I796460);
DFFARX1 I_11062 (I190568,I2507,I190127,I190594,);
nand I_11063 (I190602,I190594,I190260);
nor I_11064 (I190104,I190602,I190410);
nor I_11065 (I190098,I190594,I190226);
DFFARX1 I_11066 (I190594,I2507,I190127,I190656,);
not I_11067 (I190664,I190656);
nor I_11068 (I190113,I190664,I190376);
not I_11069 (I190722,I2514);
DFFARX1 I_11070 (I1155474,I2507,I190722,I190748,);
DFFARX1 I_11071 (I190748,I2507,I190722,I190765,);
not I_11072 (I190714,I190765);
not I_11073 (I190787,I190748);
DFFARX1 I_11074 (I1155474,I2507,I190722,I190813,);
not I_11075 (I190821,I190813);
and I_11076 (I190838,I190787,I1155477);
not I_11077 (I190855,I1155489);
nand I_11078 (I190872,I190855,I1155477);
not I_11079 (I190889,I1155495);
nor I_11080 (I190906,I190889,I1155486);
nand I_11081 (I190923,I190906,I1155492);
nor I_11082 (I190940,I190923,I190872);
DFFARX1 I_11083 (I190940,I2507,I190722,I190690,);
not I_11084 (I190971,I190923);
not I_11085 (I190988,I1155486);
nand I_11086 (I191005,I190988,I1155477);
nor I_11087 (I191022,I1155486,I1155489);
nand I_11088 (I190702,I190838,I191022);
nand I_11089 (I190696,I190787,I1155486);
nand I_11090 (I191067,I190889,I1155483);
DFFARX1 I_11091 (I191067,I2507,I190722,I190711,);
DFFARX1 I_11092 (I191067,I2507,I190722,I190705,);
not I_11093 (I191112,I1155483);
nor I_11094 (I191129,I191112,I1155480);
and I_11095 (I191146,I191129,I1155498);
or I_11096 (I191163,I191146,I1155477);
DFFARX1 I_11097 (I191163,I2507,I190722,I191189,);
nand I_11098 (I191197,I191189,I190855);
nor I_11099 (I190699,I191197,I191005);
nor I_11100 (I190693,I191189,I190821);
DFFARX1 I_11101 (I191189,I2507,I190722,I191251,);
not I_11102 (I191259,I191251);
nor I_11103 (I190708,I191259,I190971);
not I_11104 (I191317,I2514);
DFFARX1 I_11105 (I366130,I2507,I191317,I191343,);
DFFARX1 I_11106 (I191343,I2507,I191317,I191360,);
not I_11107 (I191309,I191360);
not I_11108 (I191382,I191343);
DFFARX1 I_11109 (I366145,I2507,I191317,I191408,);
not I_11110 (I191416,I191408);
and I_11111 (I191433,I191382,I366142);
not I_11112 (I191450,I366130);
nand I_11113 (I191467,I191450,I366142);
not I_11114 (I191484,I366139);
nor I_11115 (I191501,I191484,I366154);
nand I_11116 (I191518,I191501,I366151);
nor I_11117 (I191535,I191518,I191467);
DFFARX1 I_11118 (I191535,I2507,I191317,I191285,);
not I_11119 (I191566,I191518);
not I_11120 (I191583,I366154);
nand I_11121 (I191600,I191583,I366142);
nor I_11122 (I191617,I366154,I366130);
nand I_11123 (I191297,I191433,I191617);
nand I_11124 (I191291,I191382,I366154);
nand I_11125 (I191662,I191484,I366148);
DFFARX1 I_11126 (I191662,I2507,I191317,I191306,);
DFFARX1 I_11127 (I191662,I2507,I191317,I191300,);
not I_11128 (I191707,I366148);
nor I_11129 (I191724,I191707,I366136);
and I_11130 (I191741,I191724,I366157);
or I_11131 (I191758,I191741,I366133);
DFFARX1 I_11132 (I191758,I2507,I191317,I191784,);
nand I_11133 (I191792,I191784,I191450);
nor I_11134 (I191294,I191792,I191600);
nor I_11135 (I191288,I191784,I191416);
DFFARX1 I_11136 (I191784,I2507,I191317,I191846,);
not I_11137 (I191854,I191846);
nor I_11138 (I191303,I191854,I191566);
not I_11139 (I191912,I2514);
DFFARX1 I_11140 (I258095,I2507,I191912,I191938,);
DFFARX1 I_11141 (I191938,I2507,I191912,I191955,);
not I_11142 (I191904,I191955);
not I_11143 (I191977,I191938);
DFFARX1 I_11144 (I258110,I2507,I191912,I192003,);
not I_11145 (I192011,I192003);
and I_11146 (I192028,I191977,I258107);
not I_11147 (I192045,I258095);
nand I_11148 (I192062,I192045,I258107);
not I_11149 (I192079,I258104);
nor I_11150 (I192096,I192079,I258119);
nand I_11151 (I192113,I192096,I258116);
nor I_11152 (I192130,I192113,I192062);
DFFARX1 I_11153 (I192130,I2507,I191912,I191880,);
not I_11154 (I192161,I192113);
not I_11155 (I192178,I258119);
nand I_11156 (I192195,I192178,I258107);
nor I_11157 (I192212,I258119,I258095);
nand I_11158 (I191892,I192028,I192212);
nand I_11159 (I191886,I191977,I258119);
nand I_11160 (I192257,I192079,I258113);
DFFARX1 I_11161 (I192257,I2507,I191912,I191901,);
DFFARX1 I_11162 (I192257,I2507,I191912,I191895,);
not I_11163 (I192302,I258113);
nor I_11164 (I192319,I192302,I258101);
and I_11165 (I192336,I192319,I258122);
or I_11166 (I192353,I192336,I258098);
DFFARX1 I_11167 (I192353,I2507,I191912,I192379,);
nand I_11168 (I192387,I192379,I192045);
nor I_11169 (I191889,I192387,I192195);
nor I_11170 (I191883,I192379,I192011);
DFFARX1 I_11171 (I192379,I2507,I191912,I192441,);
not I_11172 (I192449,I192441);
nor I_11173 (I191898,I192449,I192161);
not I_11174 (I192507,I2514);
DFFARX1 I_11175 (I524446,I2507,I192507,I192533,);
DFFARX1 I_11176 (I192533,I2507,I192507,I192550,);
not I_11177 (I192499,I192550);
not I_11178 (I192572,I192533);
DFFARX1 I_11179 (I524440,I2507,I192507,I192598,);
not I_11180 (I192606,I192598);
and I_11181 (I192623,I192572,I524455);
not I_11182 (I192640,I524452);
nand I_11183 (I192657,I192640,I524455);
not I_11184 (I192674,I524443);
nor I_11185 (I192691,I192674,I524434);
nand I_11186 (I192708,I192691,I524437);
nor I_11187 (I192725,I192708,I192657);
DFFARX1 I_11188 (I192725,I2507,I192507,I192475,);
not I_11189 (I192756,I192708);
not I_11190 (I192773,I524434);
nand I_11191 (I192790,I192773,I524455);
nor I_11192 (I192807,I524434,I524452);
nand I_11193 (I192487,I192623,I192807);
nand I_11194 (I192481,I192572,I524434);
nand I_11195 (I192852,I192674,I524458);
DFFARX1 I_11196 (I192852,I2507,I192507,I192496,);
DFFARX1 I_11197 (I192852,I2507,I192507,I192490,);
not I_11198 (I192897,I524458);
nor I_11199 (I192914,I192897,I524449);
and I_11200 (I192931,I192914,I524434);
or I_11201 (I192948,I192931,I524437);
DFFARX1 I_11202 (I192948,I2507,I192507,I192974,);
nand I_11203 (I192982,I192974,I192640);
nor I_11204 (I192484,I192982,I192790);
nor I_11205 (I192478,I192974,I192606);
DFFARX1 I_11206 (I192974,I2507,I192507,I193036,);
not I_11207 (I193044,I193036);
nor I_11208 (I192493,I193044,I192756);
not I_11209 (I193102,I2514);
DFFARX1 I_11210 (I844941,I2507,I193102,I193128,);
DFFARX1 I_11211 (I193128,I2507,I193102,I193145,);
not I_11212 (I193094,I193145);
not I_11213 (I193167,I193128);
DFFARX1 I_11214 (I844935,I2507,I193102,I193193,);
not I_11215 (I193201,I193193);
and I_11216 (I193218,I193167,I844953);
not I_11217 (I193235,I844941);
nand I_11218 (I193252,I193235,I844953);
not I_11219 (I193269,I844935);
nor I_11220 (I193286,I193269,I844947);
nand I_11221 (I193303,I193286,I844938);
nor I_11222 (I193320,I193303,I193252);
DFFARX1 I_11223 (I193320,I2507,I193102,I193070,);
not I_11224 (I193351,I193303);
not I_11225 (I193368,I844947);
nand I_11226 (I193385,I193368,I844953);
nor I_11227 (I193402,I844947,I844941);
nand I_11228 (I193082,I193218,I193402);
nand I_11229 (I193076,I193167,I844947);
nand I_11230 (I193447,I193269,I844950);
DFFARX1 I_11231 (I193447,I2507,I193102,I193091,);
DFFARX1 I_11232 (I193447,I2507,I193102,I193085,);
not I_11233 (I193492,I844950);
nor I_11234 (I193509,I193492,I844956);
and I_11235 (I193526,I193509,I844938);
or I_11236 (I193543,I193526,I844944);
DFFARX1 I_11237 (I193543,I2507,I193102,I193569,);
nand I_11238 (I193577,I193569,I193235);
nor I_11239 (I193079,I193577,I193385);
nor I_11240 (I193073,I193569,I193201);
DFFARX1 I_11241 (I193569,I2507,I193102,I193631,);
not I_11242 (I193639,I193631);
nor I_11243 (I193088,I193639,I193351);
not I_11244 (I193697,I2514);
DFFARX1 I_11245 (I670612,I2507,I193697,I193723,);
DFFARX1 I_11246 (I193723,I2507,I193697,I193740,);
not I_11247 (I193689,I193740);
not I_11248 (I193762,I193723);
DFFARX1 I_11249 (I670609,I2507,I193697,I193788,);
not I_11250 (I193796,I193788);
and I_11251 (I193813,I193762,I670615);
not I_11252 (I193830,I670600);
nand I_11253 (I193847,I193830,I670615);
not I_11254 (I193864,I670603);
nor I_11255 (I193881,I193864,I670624);
nand I_11256 (I193898,I193881,I670621);
nor I_11257 (I193915,I193898,I193847);
DFFARX1 I_11258 (I193915,I2507,I193697,I193665,);
not I_11259 (I193946,I193898);
not I_11260 (I193963,I670624);
nand I_11261 (I193980,I193963,I670615);
nor I_11262 (I193997,I670624,I670600);
nand I_11263 (I193677,I193813,I193997);
nand I_11264 (I193671,I193762,I670624);
nand I_11265 (I194042,I193864,I670600);
DFFARX1 I_11266 (I194042,I2507,I193697,I193686,);
DFFARX1 I_11267 (I194042,I2507,I193697,I193680,);
not I_11268 (I194087,I670600);
nor I_11269 (I194104,I194087,I670606);
and I_11270 (I194121,I194104,I670618);
or I_11271 (I194138,I194121,I670603);
DFFARX1 I_11272 (I194138,I2507,I193697,I194164,);
nand I_11273 (I194172,I194164,I193830);
nor I_11274 (I193674,I194172,I193980);
nor I_11275 (I193668,I194164,I193796);
DFFARX1 I_11276 (I194164,I2507,I193697,I194226,);
not I_11277 (I194234,I194226);
nor I_11278 (I193683,I194234,I193946);
not I_11279 (I194292,I2514);
DFFARX1 I_11280 (I1342818,I2507,I194292,I194318,);
DFFARX1 I_11281 (I194318,I2507,I194292,I194335,);
not I_11282 (I194284,I194335);
not I_11283 (I194357,I194318);
DFFARX1 I_11284 (I1342809,I2507,I194292,I194383,);
not I_11285 (I194391,I194383);
and I_11286 (I194408,I194357,I1342803);
not I_11287 (I194425,I1342797);
nand I_11288 (I194442,I194425,I1342803);
not I_11289 (I194459,I1342824);
nor I_11290 (I194476,I194459,I1342797);
nand I_11291 (I194493,I194476,I1342821);
nor I_11292 (I194510,I194493,I194442);
DFFARX1 I_11293 (I194510,I2507,I194292,I194260,);
not I_11294 (I194541,I194493);
not I_11295 (I194558,I1342797);
nand I_11296 (I194575,I194558,I1342803);
nor I_11297 (I194592,I1342797,I1342797);
nand I_11298 (I194272,I194408,I194592);
nand I_11299 (I194266,I194357,I1342797);
nand I_11300 (I194637,I194459,I1342806);
DFFARX1 I_11301 (I194637,I2507,I194292,I194281,);
DFFARX1 I_11302 (I194637,I2507,I194292,I194275,);
not I_11303 (I194682,I1342806);
nor I_11304 (I194699,I194682,I1342812);
and I_11305 (I194716,I194699,I1342815);
or I_11306 (I194733,I194716,I1342800);
DFFARX1 I_11307 (I194733,I2507,I194292,I194759,);
nand I_11308 (I194767,I194759,I194425);
nor I_11309 (I194269,I194767,I194575);
nor I_11310 (I194263,I194759,I194391);
DFFARX1 I_11311 (I194759,I2507,I194292,I194821,);
not I_11312 (I194829,I194821);
nor I_11313 (I194278,I194829,I194541);
not I_11314 (I194887,I2514);
DFFARX1 I_11315 (I1184374,I2507,I194887,I194913,);
DFFARX1 I_11316 (I194913,I2507,I194887,I194930,);
not I_11317 (I194879,I194930);
not I_11318 (I194952,I194913);
DFFARX1 I_11319 (I1184374,I2507,I194887,I194978,);
not I_11320 (I194986,I194978);
and I_11321 (I195003,I194952,I1184377);
not I_11322 (I195020,I1184389);
nand I_11323 (I195037,I195020,I1184377);
not I_11324 (I195054,I1184395);
nor I_11325 (I195071,I195054,I1184386);
nand I_11326 (I195088,I195071,I1184392);
nor I_11327 (I195105,I195088,I195037);
DFFARX1 I_11328 (I195105,I2507,I194887,I194855,);
not I_11329 (I195136,I195088);
not I_11330 (I195153,I1184386);
nand I_11331 (I195170,I195153,I1184377);
nor I_11332 (I195187,I1184386,I1184389);
nand I_11333 (I194867,I195003,I195187);
nand I_11334 (I194861,I194952,I1184386);
nand I_11335 (I195232,I195054,I1184383);
DFFARX1 I_11336 (I195232,I2507,I194887,I194876,);
DFFARX1 I_11337 (I195232,I2507,I194887,I194870,);
not I_11338 (I195277,I1184383);
nor I_11339 (I195294,I195277,I1184380);
and I_11340 (I195311,I195294,I1184398);
or I_11341 (I195328,I195311,I1184377);
DFFARX1 I_11342 (I195328,I2507,I194887,I195354,);
nand I_11343 (I195362,I195354,I195020);
nor I_11344 (I194864,I195362,I195170);
nor I_11345 (I194858,I195354,I194986);
DFFARX1 I_11346 (I195354,I2507,I194887,I195416,);
not I_11347 (I195424,I195416);
nor I_11348 (I194873,I195424,I195136);
not I_11349 (I195482,I2514);
DFFARX1 I_11350 (I574667,I2507,I195482,I195508,);
DFFARX1 I_11351 (I195508,I2507,I195482,I195525,);
not I_11352 (I195474,I195525);
not I_11353 (I195547,I195508);
DFFARX1 I_11354 (I574658,I2507,I195482,I195573,);
not I_11355 (I195581,I195573);
and I_11356 (I195598,I195547,I574676);
not I_11357 (I195615,I574673);
nand I_11358 (I195632,I195615,I574676);
not I_11359 (I195649,I574652);
nor I_11360 (I195666,I195649,I574655);
nand I_11361 (I195683,I195666,I574664);
nor I_11362 (I195700,I195683,I195632);
DFFARX1 I_11363 (I195700,I2507,I195482,I195450,);
not I_11364 (I195731,I195683);
not I_11365 (I195748,I574655);
nand I_11366 (I195765,I195748,I574676);
nor I_11367 (I195782,I574655,I574673);
nand I_11368 (I195462,I195598,I195782);
nand I_11369 (I195456,I195547,I574655);
nand I_11370 (I195827,I195649,I574670);
DFFARX1 I_11371 (I195827,I2507,I195482,I195471,);
DFFARX1 I_11372 (I195827,I2507,I195482,I195465,);
not I_11373 (I195872,I574670);
nor I_11374 (I195889,I195872,I574652);
and I_11375 (I195906,I195889,I574661);
or I_11376 (I195923,I195906,I574655);
DFFARX1 I_11377 (I195923,I2507,I195482,I195949,);
nand I_11378 (I195957,I195949,I195615);
nor I_11379 (I195459,I195957,I195765);
nor I_11380 (I195453,I195949,I195581);
DFFARX1 I_11381 (I195949,I2507,I195482,I196011,);
not I_11382 (I196019,I196011);
nor I_11383 (I195468,I196019,I195731);
not I_11384 (I196077,I2514);
DFFARX1 I_11385 (I874980,I2507,I196077,I196103,);
DFFARX1 I_11386 (I196103,I2507,I196077,I196120,);
not I_11387 (I196069,I196120);
not I_11388 (I196142,I196103);
DFFARX1 I_11389 (I874974,I2507,I196077,I196168,);
not I_11390 (I196176,I196168);
and I_11391 (I196193,I196142,I874992);
not I_11392 (I196210,I874980);
nand I_11393 (I196227,I196210,I874992);
not I_11394 (I196244,I874974);
nor I_11395 (I196261,I196244,I874986);
nand I_11396 (I196278,I196261,I874977);
nor I_11397 (I196295,I196278,I196227);
DFFARX1 I_11398 (I196295,I2507,I196077,I196045,);
not I_11399 (I196326,I196278);
not I_11400 (I196343,I874986);
nand I_11401 (I196360,I196343,I874992);
nor I_11402 (I196377,I874986,I874980);
nand I_11403 (I196057,I196193,I196377);
nand I_11404 (I196051,I196142,I874986);
nand I_11405 (I196422,I196244,I874989);
DFFARX1 I_11406 (I196422,I2507,I196077,I196066,);
DFFARX1 I_11407 (I196422,I2507,I196077,I196060,);
not I_11408 (I196467,I874989);
nor I_11409 (I196484,I196467,I874995);
and I_11410 (I196501,I196484,I874977);
or I_11411 (I196518,I196501,I874983);
DFFARX1 I_11412 (I196518,I2507,I196077,I196544,);
nand I_11413 (I196552,I196544,I196210);
nor I_11414 (I196054,I196552,I196360);
nor I_11415 (I196048,I196544,I196176);
DFFARX1 I_11416 (I196544,I2507,I196077,I196606,);
not I_11417 (I196614,I196606);
nor I_11418 (I196063,I196614,I196326);
not I_11419 (I196672,I2514);
DFFARX1 I_11420 (I545189,I2507,I196672,I196698,);
DFFARX1 I_11421 (I196698,I2507,I196672,I196715,);
not I_11422 (I196664,I196715);
not I_11423 (I196737,I196698);
DFFARX1 I_11424 (I545180,I2507,I196672,I196763,);
not I_11425 (I196771,I196763);
and I_11426 (I196788,I196737,I545198);
not I_11427 (I196805,I545195);
nand I_11428 (I196822,I196805,I545198);
not I_11429 (I196839,I545174);
nor I_11430 (I196856,I196839,I545177);
nand I_11431 (I196873,I196856,I545186);
nor I_11432 (I196890,I196873,I196822);
DFFARX1 I_11433 (I196890,I2507,I196672,I196640,);
not I_11434 (I196921,I196873);
not I_11435 (I196938,I545177);
nand I_11436 (I196955,I196938,I545198);
nor I_11437 (I196972,I545177,I545195);
nand I_11438 (I196652,I196788,I196972);
nand I_11439 (I196646,I196737,I545177);
nand I_11440 (I197017,I196839,I545192);
DFFARX1 I_11441 (I197017,I2507,I196672,I196661,);
DFFARX1 I_11442 (I197017,I2507,I196672,I196655,);
not I_11443 (I197062,I545192);
nor I_11444 (I197079,I197062,I545174);
and I_11445 (I197096,I197079,I545183);
or I_11446 (I197113,I197096,I545177);
DFFARX1 I_11447 (I197113,I2507,I196672,I197139,);
nand I_11448 (I197147,I197139,I196805);
nor I_11449 (I196649,I197147,I196955);
nor I_11450 (I196643,I197139,I196771);
DFFARX1 I_11451 (I197139,I2507,I196672,I197201,);
not I_11452 (I197209,I197201);
nor I_11453 (I196658,I197209,I196921);
not I_11454 (I197267,I2514);
DFFARX1 I_11455 (I308160,I2507,I197267,I197293,);
DFFARX1 I_11456 (I197293,I2507,I197267,I197310,);
not I_11457 (I197259,I197310);
not I_11458 (I197332,I197293);
DFFARX1 I_11459 (I308175,I2507,I197267,I197358,);
not I_11460 (I197366,I197358);
and I_11461 (I197383,I197332,I308172);
not I_11462 (I197400,I308160);
nand I_11463 (I197417,I197400,I308172);
not I_11464 (I197434,I308169);
nor I_11465 (I197451,I197434,I308184);
nand I_11466 (I197468,I197451,I308181);
nor I_11467 (I197485,I197468,I197417);
DFFARX1 I_11468 (I197485,I2507,I197267,I197235,);
not I_11469 (I197516,I197468);
not I_11470 (I197533,I308184);
nand I_11471 (I197550,I197533,I308172);
nor I_11472 (I197567,I308184,I308160);
nand I_11473 (I197247,I197383,I197567);
nand I_11474 (I197241,I197332,I308184);
nand I_11475 (I197612,I197434,I308178);
DFFARX1 I_11476 (I197612,I2507,I197267,I197256,);
DFFARX1 I_11477 (I197612,I2507,I197267,I197250,);
not I_11478 (I197657,I308178);
nor I_11479 (I197674,I197657,I308166);
and I_11480 (I197691,I197674,I308187);
or I_11481 (I197708,I197691,I308163);
DFFARX1 I_11482 (I197708,I2507,I197267,I197734,);
nand I_11483 (I197742,I197734,I197400);
nor I_11484 (I197244,I197742,I197550);
nor I_11485 (I197238,I197734,I197366);
DFFARX1 I_11486 (I197734,I2507,I197267,I197796,);
not I_11487 (I197804,I197796);
nor I_11488 (I197253,I197804,I197516);
not I_11489 (I197862,I2514);
DFFARX1 I_11490 (I992238,I2507,I197862,I197888,);
DFFARX1 I_11491 (I197888,I2507,I197862,I197905,);
not I_11492 (I197854,I197905);
not I_11493 (I197927,I197888);
DFFARX1 I_11494 (I992247,I2507,I197862,I197953,);
not I_11495 (I197961,I197953);
and I_11496 (I197978,I197927,I992235);
not I_11497 (I197995,I992226);
nand I_11498 (I198012,I197995,I992235);
not I_11499 (I198029,I992232);
nor I_11500 (I198046,I198029,I992250);
nand I_11501 (I198063,I198046,I992223);
nor I_11502 (I198080,I198063,I198012);
DFFARX1 I_11503 (I198080,I2507,I197862,I197830,);
not I_11504 (I198111,I198063);
not I_11505 (I198128,I992250);
nand I_11506 (I198145,I198128,I992235);
nor I_11507 (I198162,I992250,I992226);
nand I_11508 (I197842,I197978,I198162);
nand I_11509 (I197836,I197927,I992250);
nand I_11510 (I198207,I198029,I992229);
DFFARX1 I_11511 (I198207,I2507,I197862,I197851,);
DFFARX1 I_11512 (I198207,I2507,I197862,I197845,);
not I_11513 (I198252,I992229);
nor I_11514 (I198269,I198252,I992241);
and I_11515 (I198286,I198269,I992223);
or I_11516 (I198303,I198286,I992244);
DFFARX1 I_11517 (I198303,I2507,I197862,I198329,);
nand I_11518 (I198337,I198329,I197995);
nor I_11519 (I197839,I198337,I198145);
nor I_11520 (I197833,I198329,I197961);
DFFARX1 I_11521 (I198329,I2507,I197862,I198391,);
not I_11522 (I198399,I198391);
nor I_11523 (I197848,I198399,I198111);
not I_11524 (I198457,I2514);
DFFARX1 I_11525 (I634776,I2507,I198457,I198483,);
DFFARX1 I_11526 (I198483,I2507,I198457,I198500,);
not I_11527 (I198449,I198500);
not I_11528 (I198522,I198483);
DFFARX1 I_11529 (I634773,I2507,I198457,I198548,);
not I_11530 (I198556,I198548);
and I_11531 (I198573,I198522,I634779);
not I_11532 (I198590,I634764);
nand I_11533 (I198607,I198590,I634779);
not I_11534 (I198624,I634767);
nor I_11535 (I198641,I198624,I634788);
nand I_11536 (I198658,I198641,I634785);
nor I_11537 (I198675,I198658,I198607);
DFFARX1 I_11538 (I198675,I2507,I198457,I198425,);
not I_11539 (I198706,I198658);
not I_11540 (I198723,I634788);
nand I_11541 (I198740,I198723,I634779);
nor I_11542 (I198757,I634788,I634764);
nand I_11543 (I198437,I198573,I198757);
nand I_11544 (I198431,I198522,I634788);
nand I_11545 (I198802,I198624,I634764);
DFFARX1 I_11546 (I198802,I2507,I198457,I198446,);
DFFARX1 I_11547 (I198802,I2507,I198457,I198440,);
not I_11548 (I198847,I634764);
nor I_11549 (I198864,I198847,I634770);
and I_11550 (I198881,I198864,I634782);
or I_11551 (I198898,I198881,I634767);
DFFARX1 I_11552 (I198898,I2507,I198457,I198924,);
nand I_11553 (I198932,I198924,I198590);
nor I_11554 (I198434,I198932,I198740);
nor I_11555 (I198428,I198924,I198556);
DFFARX1 I_11556 (I198924,I2507,I198457,I198986,);
not I_11557 (I198994,I198986);
nor I_11558 (I198443,I198994,I198706);
not I_11559 (I199052,I2514);
DFFARX1 I_11560 (I1273831,I2507,I199052,I199078,);
DFFARX1 I_11561 (I199078,I2507,I199052,I199095,);
not I_11562 (I199044,I199095);
not I_11563 (I199117,I199078);
DFFARX1 I_11564 (I1273843,I2507,I199052,I199143,);
not I_11565 (I199151,I199143);
and I_11566 (I199168,I199117,I1273837);
not I_11567 (I199185,I1273849);
nand I_11568 (I199202,I199185,I1273837);
not I_11569 (I199219,I1273834);
nor I_11570 (I199236,I199219,I1273846);
nand I_11571 (I199253,I199236,I1273828);
nor I_11572 (I199270,I199253,I199202);
DFFARX1 I_11573 (I199270,I2507,I199052,I199020,);
not I_11574 (I199301,I199253);
not I_11575 (I199318,I1273846);
nand I_11576 (I199335,I199318,I1273837);
nor I_11577 (I199352,I1273846,I1273849);
nand I_11578 (I199032,I199168,I199352);
nand I_11579 (I199026,I199117,I1273846);
nand I_11580 (I199397,I199219,I1273840);
DFFARX1 I_11581 (I199397,I2507,I199052,I199041,);
DFFARX1 I_11582 (I199397,I2507,I199052,I199035,);
not I_11583 (I199442,I1273840);
nor I_11584 (I199459,I199442,I1273831);
and I_11585 (I199476,I199459,I1273828);
or I_11586 (I199493,I199476,I1273852);
DFFARX1 I_11587 (I199493,I2507,I199052,I199519,);
nand I_11588 (I199527,I199519,I199185);
nor I_11589 (I199029,I199527,I199335);
nor I_11590 (I199023,I199519,I199151);
DFFARX1 I_11591 (I199519,I2507,I199052,I199581,);
not I_11592 (I199589,I199581);
nor I_11593 (I199038,I199589,I199301);
not I_11594 (I199647,I2514);
DFFARX1 I_11595 (I1258803,I2507,I199647,I199673,);
DFFARX1 I_11596 (I199673,I2507,I199647,I199690,);
not I_11597 (I199639,I199690);
not I_11598 (I199712,I199673);
DFFARX1 I_11599 (I1258815,I2507,I199647,I199738,);
not I_11600 (I199746,I199738);
and I_11601 (I199763,I199712,I1258809);
not I_11602 (I199780,I1258821);
nand I_11603 (I199797,I199780,I1258809);
not I_11604 (I199814,I1258806);
nor I_11605 (I199831,I199814,I1258818);
nand I_11606 (I199848,I199831,I1258800);
nor I_11607 (I199865,I199848,I199797);
DFFARX1 I_11608 (I199865,I2507,I199647,I199615,);
not I_11609 (I199896,I199848);
not I_11610 (I199913,I1258818);
nand I_11611 (I199930,I199913,I1258809);
nor I_11612 (I199947,I1258818,I1258821);
nand I_11613 (I199627,I199763,I199947);
nand I_11614 (I199621,I199712,I1258818);
nand I_11615 (I199992,I199814,I1258812);
DFFARX1 I_11616 (I199992,I2507,I199647,I199636,);
DFFARX1 I_11617 (I199992,I2507,I199647,I199630,);
not I_11618 (I200037,I1258812);
nor I_11619 (I200054,I200037,I1258803);
and I_11620 (I200071,I200054,I1258800);
or I_11621 (I200088,I200071,I1258824);
DFFARX1 I_11622 (I200088,I2507,I199647,I200114,);
nand I_11623 (I200122,I200114,I199780);
nor I_11624 (I199624,I200122,I199930);
nor I_11625 (I199618,I200114,I199746);
DFFARX1 I_11626 (I200114,I2507,I199647,I200176,);
not I_11627 (I200184,I200176);
nor I_11628 (I199633,I200184,I199896);
not I_11629 (I200242,I2514);
DFFARX1 I_11630 (I1312473,I2507,I200242,I200268,);
DFFARX1 I_11631 (I200268,I2507,I200242,I200285,);
not I_11632 (I200234,I200285);
not I_11633 (I200307,I200268);
DFFARX1 I_11634 (I1312464,I2507,I200242,I200333,);
not I_11635 (I200341,I200333);
and I_11636 (I200358,I200307,I1312458);
not I_11637 (I200375,I1312452);
nand I_11638 (I200392,I200375,I1312458);
not I_11639 (I200409,I1312479);
nor I_11640 (I200426,I200409,I1312452);
nand I_11641 (I200443,I200426,I1312476);
nor I_11642 (I200460,I200443,I200392);
DFFARX1 I_11643 (I200460,I2507,I200242,I200210,);
not I_11644 (I200491,I200443);
not I_11645 (I200508,I1312452);
nand I_11646 (I200525,I200508,I1312458);
nor I_11647 (I200542,I1312452,I1312452);
nand I_11648 (I200222,I200358,I200542);
nand I_11649 (I200216,I200307,I1312452);
nand I_11650 (I200587,I200409,I1312461);
DFFARX1 I_11651 (I200587,I2507,I200242,I200231,);
DFFARX1 I_11652 (I200587,I2507,I200242,I200225,);
not I_11653 (I200632,I1312461);
nor I_11654 (I200649,I200632,I1312467);
and I_11655 (I200666,I200649,I1312470);
or I_11656 (I200683,I200666,I1312455);
DFFARX1 I_11657 (I200683,I2507,I200242,I200709,);
nand I_11658 (I200717,I200709,I200375);
nor I_11659 (I200219,I200717,I200525);
nor I_11660 (I200213,I200709,I200341);
DFFARX1 I_11661 (I200709,I2507,I200242,I200771,);
not I_11662 (I200779,I200771);
nor I_11663 (I200228,I200779,I200491);
not I_11664 (I200837,I2514);
DFFARX1 I_11665 (I372981,I2507,I200837,I200863,);
DFFARX1 I_11666 (I200863,I2507,I200837,I200880,);
not I_11667 (I200829,I200880);
not I_11668 (I200902,I200863);
DFFARX1 I_11669 (I372996,I2507,I200837,I200928,);
not I_11670 (I200936,I200928);
and I_11671 (I200953,I200902,I372993);
not I_11672 (I200970,I372981);
nand I_11673 (I200987,I200970,I372993);
not I_11674 (I201004,I372990);
nor I_11675 (I201021,I201004,I373005);
nand I_11676 (I201038,I201021,I373002);
nor I_11677 (I201055,I201038,I200987);
DFFARX1 I_11678 (I201055,I2507,I200837,I200805,);
not I_11679 (I201086,I201038);
not I_11680 (I201103,I373005);
nand I_11681 (I201120,I201103,I372993);
nor I_11682 (I201137,I373005,I372981);
nand I_11683 (I200817,I200953,I201137);
nand I_11684 (I200811,I200902,I373005);
nand I_11685 (I201182,I201004,I372999);
DFFARX1 I_11686 (I201182,I2507,I200837,I200826,);
DFFARX1 I_11687 (I201182,I2507,I200837,I200820,);
not I_11688 (I201227,I372999);
nor I_11689 (I201244,I201227,I372987);
and I_11690 (I201261,I201244,I373008);
or I_11691 (I201278,I201261,I372984);
DFFARX1 I_11692 (I201278,I2507,I200837,I201304,);
nand I_11693 (I201312,I201304,I200970);
nor I_11694 (I200814,I201312,I201120);
nor I_11695 (I200808,I201304,I200936);
DFFARX1 I_11696 (I201304,I2507,I200837,I201366,);
not I_11697 (I201374,I201366);
nor I_11698 (I200823,I201374,I201086);
not I_11699 (I201432,I2514);
DFFARX1 I_11700 (I525041,I2507,I201432,I201458,);
DFFARX1 I_11701 (I201458,I2507,I201432,I201475,);
not I_11702 (I201424,I201475);
not I_11703 (I201497,I201458);
DFFARX1 I_11704 (I525035,I2507,I201432,I201523,);
not I_11705 (I201531,I201523);
and I_11706 (I201548,I201497,I525050);
not I_11707 (I201565,I525047);
nand I_11708 (I201582,I201565,I525050);
not I_11709 (I201599,I525038);
nor I_11710 (I201616,I201599,I525029);
nand I_11711 (I201633,I201616,I525032);
nor I_11712 (I201650,I201633,I201582);
DFFARX1 I_11713 (I201650,I2507,I201432,I201400,);
not I_11714 (I201681,I201633);
not I_11715 (I201698,I525029);
nand I_11716 (I201715,I201698,I525050);
nor I_11717 (I201732,I525029,I525047);
nand I_11718 (I201412,I201548,I201732);
nand I_11719 (I201406,I201497,I525029);
nand I_11720 (I201777,I201599,I525053);
DFFARX1 I_11721 (I201777,I2507,I201432,I201421,);
DFFARX1 I_11722 (I201777,I2507,I201432,I201415,);
not I_11723 (I201822,I525053);
nor I_11724 (I201839,I201822,I525044);
and I_11725 (I201856,I201839,I525029);
or I_11726 (I201873,I201856,I525032);
DFFARX1 I_11727 (I201873,I2507,I201432,I201899,);
nand I_11728 (I201907,I201899,I201565);
nor I_11729 (I201409,I201907,I201715);
nor I_11730 (I201403,I201899,I201531);
DFFARX1 I_11731 (I201899,I2507,I201432,I201961,);
not I_11732 (I201969,I201961);
nor I_11733 (I201418,I201969,I201681);
not I_11734 (I202027,I2514);
DFFARX1 I_11735 (I1161832,I2507,I202027,I202053,);
DFFARX1 I_11736 (I202053,I2507,I202027,I202070,);
not I_11737 (I202019,I202070);
not I_11738 (I202092,I202053);
DFFARX1 I_11739 (I1161832,I2507,I202027,I202118,);
not I_11740 (I202126,I202118);
and I_11741 (I202143,I202092,I1161835);
not I_11742 (I202160,I1161847);
nand I_11743 (I202177,I202160,I1161835);
not I_11744 (I202194,I1161853);
nor I_11745 (I202211,I202194,I1161844);
nand I_11746 (I202228,I202211,I1161850);
nor I_11747 (I202245,I202228,I202177);
DFFARX1 I_11748 (I202245,I2507,I202027,I201995,);
not I_11749 (I202276,I202228);
not I_11750 (I202293,I1161844);
nand I_11751 (I202310,I202293,I1161835);
nor I_11752 (I202327,I1161844,I1161847);
nand I_11753 (I202007,I202143,I202327);
nand I_11754 (I202001,I202092,I1161844);
nand I_11755 (I202372,I202194,I1161841);
DFFARX1 I_11756 (I202372,I2507,I202027,I202016,);
DFFARX1 I_11757 (I202372,I2507,I202027,I202010,);
not I_11758 (I202417,I1161841);
nor I_11759 (I202434,I202417,I1161838);
and I_11760 (I202451,I202434,I1161856);
or I_11761 (I202468,I202451,I1161835);
DFFARX1 I_11762 (I202468,I2507,I202027,I202494,);
nand I_11763 (I202502,I202494,I202160);
nor I_11764 (I202004,I202502,I202310);
nor I_11765 (I201998,I202494,I202126);
DFFARX1 I_11766 (I202494,I2507,I202027,I202556,);
not I_11767 (I202564,I202556);
nor I_11768 (I202013,I202564,I202276);
not I_11769 (I202622,I2514);
DFFARX1 I_11770 (I829131,I2507,I202622,I202648,);
DFFARX1 I_11771 (I202648,I2507,I202622,I202665,);
not I_11772 (I202614,I202665);
not I_11773 (I202687,I202648);
DFFARX1 I_11774 (I829125,I2507,I202622,I202713,);
not I_11775 (I202721,I202713);
and I_11776 (I202738,I202687,I829143);
not I_11777 (I202755,I829131);
nand I_11778 (I202772,I202755,I829143);
not I_11779 (I202789,I829125);
nor I_11780 (I202806,I202789,I829137);
nand I_11781 (I202823,I202806,I829128);
nor I_11782 (I202840,I202823,I202772);
DFFARX1 I_11783 (I202840,I2507,I202622,I202590,);
not I_11784 (I202871,I202823);
not I_11785 (I202888,I829137);
nand I_11786 (I202905,I202888,I829143);
nor I_11787 (I202922,I829137,I829131);
nand I_11788 (I202602,I202738,I202922);
nand I_11789 (I202596,I202687,I829137);
nand I_11790 (I202967,I202789,I829140);
DFFARX1 I_11791 (I202967,I2507,I202622,I202611,);
DFFARX1 I_11792 (I202967,I2507,I202622,I202605,);
not I_11793 (I203012,I829140);
nor I_11794 (I203029,I203012,I829146);
and I_11795 (I203046,I203029,I829128);
or I_11796 (I203063,I203046,I829134);
DFFARX1 I_11797 (I203063,I2507,I202622,I203089,);
nand I_11798 (I203097,I203089,I202755);
nor I_11799 (I202599,I203097,I202905);
nor I_11800 (I202593,I203089,I202721);
DFFARX1 I_11801 (I203089,I2507,I202622,I203151,);
not I_11802 (I203159,I203151);
nor I_11803 (I202608,I203159,I202871);
not I_11804 (I203217,I2514);
DFFARX1 I_11805 (I1375543,I2507,I203217,I203243,);
DFFARX1 I_11806 (I203243,I2507,I203217,I203260,);
not I_11807 (I203209,I203260);
not I_11808 (I203282,I203243);
DFFARX1 I_11809 (I1375534,I2507,I203217,I203308,);
not I_11810 (I203316,I203308);
and I_11811 (I203333,I203282,I1375528);
not I_11812 (I203350,I1375522);
nand I_11813 (I203367,I203350,I1375528);
not I_11814 (I203384,I1375549);
nor I_11815 (I203401,I203384,I1375522);
nand I_11816 (I203418,I203401,I1375546);
nor I_11817 (I203435,I203418,I203367);
DFFARX1 I_11818 (I203435,I2507,I203217,I203185,);
not I_11819 (I203466,I203418);
not I_11820 (I203483,I1375522);
nand I_11821 (I203500,I203483,I1375528);
nor I_11822 (I203517,I1375522,I1375522);
nand I_11823 (I203197,I203333,I203517);
nand I_11824 (I203191,I203282,I1375522);
nand I_11825 (I203562,I203384,I1375531);
DFFARX1 I_11826 (I203562,I2507,I203217,I203206,);
DFFARX1 I_11827 (I203562,I2507,I203217,I203200,);
not I_11828 (I203607,I1375531);
nor I_11829 (I203624,I203607,I1375537);
and I_11830 (I203641,I203624,I1375540);
or I_11831 (I203658,I203641,I1375525);
DFFARX1 I_11832 (I203658,I2507,I203217,I203684,);
nand I_11833 (I203692,I203684,I203350);
nor I_11834 (I203194,I203692,I203500);
nor I_11835 (I203188,I203684,I203316);
DFFARX1 I_11836 (I203684,I2507,I203217,I203746,);
not I_11837 (I203754,I203746);
nor I_11838 (I203203,I203754,I203466);
not I_11839 (I203812,I2514);
DFFARX1 I_11840 (I483335,I2507,I203812,I203838,);
DFFARX1 I_11841 (I203838,I2507,I203812,I203855,);
not I_11842 (I203804,I203855);
not I_11843 (I203877,I203838);
DFFARX1 I_11844 (I483323,I2507,I203812,I203903,);
not I_11845 (I203911,I203903);
and I_11846 (I203928,I203877,I483332);
not I_11847 (I203945,I483329);
nand I_11848 (I203962,I203945,I483332);
not I_11849 (I203979,I483320);
nor I_11850 (I203996,I203979,I483326);
nand I_11851 (I204013,I203996,I483311);
nor I_11852 (I204030,I204013,I203962);
DFFARX1 I_11853 (I204030,I2507,I203812,I203780,);
not I_11854 (I204061,I204013);
not I_11855 (I204078,I483326);
nand I_11856 (I204095,I204078,I483332);
nor I_11857 (I204112,I483326,I483329);
nand I_11858 (I203792,I203928,I204112);
nand I_11859 (I203786,I203877,I483326);
nand I_11860 (I204157,I203979,I483311);
DFFARX1 I_11861 (I204157,I2507,I203812,I203801,);
DFFARX1 I_11862 (I204157,I2507,I203812,I203795,);
not I_11863 (I204202,I483311);
nor I_11864 (I204219,I204202,I483317);
and I_11865 (I204236,I204219,I483314);
or I_11866 (I204253,I204236,I483338);
DFFARX1 I_11867 (I204253,I2507,I203812,I204279,);
nand I_11868 (I204287,I204279,I203945);
nor I_11869 (I203789,I204287,I204095);
nor I_11870 (I203783,I204279,I203911);
DFFARX1 I_11871 (I204279,I2507,I203812,I204341,);
not I_11872 (I204349,I204341);
nor I_11873 (I203798,I204349,I204061);
not I_11874 (I204407,I2514);
DFFARX1 I_11875 (I838090,I2507,I204407,I204433,);
DFFARX1 I_11876 (I204433,I2507,I204407,I204450,);
not I_11877 (I204399,I204450);
not I_11878 (I204472,I204433);
DFFARX1 I_11879 (I838084,I2507,I204407,I204498,);
not I_11880 (I204506,I204498);
and I_11881 (I204523,I204472,I838102);
not I_11882 (I204540,I838090);
nand I_11883 (I204557,I204540,I838102);
not I_11884 (I204574,I838084);
nor I_11885 (I204591,I204574,I838096);
nand I_11886 (I204608,I204591,I838087);
nor I_11887 (I204625,I204608,I204557);
DFFARX1 I_11888 (I204625,I2507,I204407,I204375,);
not I_11889 (I204656,I204608);
not I_11890 (I204673,I838096);
nand I_11891 (I204690,I204673,I838102);
nor I_11892 (I204707,I838096,I838090);
nand I_11893 (I204387,I204523,I204707);
nand I_11894 (I204381,I204472,I838096);
nand I_11895 (I204752,I204574,I838099);
DFFARX1 I_11896 (I204752,I2507,I204407,I204396,);
DFFARX1 I_11897 (I204752,I2507,I204407,I204390,);
not I_11898 (I204797,I838099);
nor I_11899 (I204814,I204797,I838105);
and I_11900 (I204831,I204814,I838087);
or I_11901 (I204848,I204831,I838093);
DFFARX1 I_11902 (I204848,I2507,I204407,I204874,);
nand I_11903 (I204882,I204874,I204540);
nor I_11904 (I204384,I204882,I204690);
nor I_11905 (I204378,I204874,I204506);
DFFARX1 I_11906 (I204874,I2507,I204407,I204936,);
not I_11907 (I204944,I204936);
nor I_11908 (I204393,I204944,I204656);
not I_11909 (I205002,I2514);
DFFARX1 I_11910 (I608769,I2507,I205002,I205028,);
DFFARX1 I_11911 (I205028,I2507,I205002,I205045,);
not I_11912 (I204994,I205045);
not I_11913 (I205067,I205028);
DFFARX1 I_11914 (I608760,I2507,I205002,I205093,);
not I_11915 (I205101,I205093);
and I_11916 (I205118,I205067,I608778);
not I_11917 (I205135,I608775);
nand I_11918 (I205152,I205135,I608778);
not I_11919 (I205169,I608754);
nor I_11920 (I205186,I205169,I608757);
nand I_11921 (I205203,I205186,I608766);
nor I_11922 (I205220,I205203,I205152);
DFFARX1 I_11923 (I205220,I2507,I205002,I204970,);
not I_11924 (I205251,I205203);
not I_11925 (I205268,I608757);
nand I_11926 (I205285,I205268,I608778);
nor I_11927 (I205302,I608757,I608775);
nand I_11928 (I204982,I205118,I205302);
nand I_11929 (I204976,I205067,I608757);
nand I_11930 (I205347,I205169,I608772);
DFFARX1 I_11931 (I205347,I2507,I205002,I204991,);
DFFARX1 I_11932 (I205347,I2507,I205002,I204985,);
not I_11933 (I205392,I608772);
nor I_11934 (I205409,I205392,I608754);
and I_11935 (I205426,I205409,I608763);
or I_11936 (I205443,I205426,I608757);
DFFARX1 I_11937 (I205443,I2507,I205002,I205469,);
nand I_11938 (I205477,I205469,I205135);
nor I_11939 (I204979,I205477,I205285);
nor I_11940 (I204973,I205469,I205101);
DFFARX1 I_11941 (I205469,I2507,I205002,I205531,);
not I_11942 (I205539,I205531);
nor I_11943 (I204988,I205539,I205251);
not I_11944 (I205597,I2514);
DFFARX1 I_11945 (I1300324,I2507,I205597,I205623,);
DFFARX1 I_11946 (I205623,I2507,I205597,I205640,);
not I_11947 (I205589,I205640);
not I_11948 (I205662,I205623);
DFFARX1 I_11949 (I1300297,I2507,I205597,I205688,);
not I_11950 (I205696,I205688);
and I_11951 (I205713,I205662,I1300321);
not I_11952 (I205730,I1300318);
nand I_11953 (I205747,I205730,I1300321);
not I_11954 (I205764,I1300297);
nor I_11955 (I205781,I205764,I1300315);
nand I_11956 (I205798,I205781,I1300303);
nor I_11957 (I205815,I205798,I205747);
DFFARX1 I_11958 (I205815,I2507,I205597,I205565,);
not I_11959 (I205846,I205798);
not I_11960 (I205863,I1300315);
nand I_11961 (I205880,I205863,I1300321);
nor I_11962 (I205897,I1300315,I1300318);
nand I_11963 (I205577,I205713,I205897);
nand I_11964 (I205571,I205662,I1300315);
nand I_11965 (I205942,I205764,I1300309);
DFFARX1 I_11966 (I205942,I2507,I205597,I205586,);
DFFARX1 I_11967 (I205942,I2507,I205597,I205580,);
not I_11968 (I205987,I1300309);
nor I_11969 (I206004,I205987,I1300312);
and I_11970 (I206021,I206004,I1300300);
or I_11971 (I206038,I206021,I1300306);
DFFARX1 I_11972 (I206038,I2507,I205597,I206064,);
nand I_11973 (I206072,I206064,I205730);
nor I_11974 (I205574,I206072,I205880);
nor I_11975 (I205568,I206064,I205696);
DFFARX1 I_11976 (I206064,I2507,I205597,I206126,);
not I_11977 (I206134,I206126);
nor I_11978 (I205583,I206134,I205846);
not I_11979 (I206192,I2514);
DFFARX1 I_11980 (I866548,I2507,I206192,I206218,);
DFFARX1 I_11981 (I206218,I2507,I206192,I206235,);
not I_11982 (I206184,I206235);
not I_11983 (I206257,I206218);
DFFARX1 I_11984 (I866542,I2507,I206192,I206283,);
not I_11985 (I206291,I206283);
and I_11986 (I206308,I206257,I866560);
not I_11987 (I206325,I866548);
nand I_11988 (I206342,I206325,I866560);
not I_11989 (I206359,I866542);
nor I_11990 (I206376,I206359,I866554);
nand I_11991 (I206393,I206376,I866545);
nor I_11992 (I206410,I206393,I206342);
DFFARX1 I_11993 (I206410,I2507,I206192,I206160,);
not I_11994 (I206441,I206393);
not I_11995 (I206458,I866554);
nand I_11996 (I206475,I206458,I866560);
nor I_11997 (I206492,I866554,I866548);
nand I_11998 (I206172,I206308,I206492);
nand I_11999 (I206166,I206257,I866554);
nand I_12000 (I206537,I206359,I866557);
DFFARX1 I_12001 (I206537,I2507,I206192,I206181,);
DFFARX1 I_12002 (I206537,I2507,I206192,I206175,);
not I_12003 (I206582,I866557);
nor I_12004 (I206599,I206582,I866563);
and I_12005 (I206616,I206599,I866545);
or I_12006 (I206633,I206616,I866551);
DFFARX1 I_12007 (I206633,I2507,I206192,I206659,);
nand I_12008 (I206667,I206659,I206325);
nor I_12009 (I206169,I206667,I206475);
nor I_12010 (I206163,I206659,I206291);
DFFARX1 I_12011 (I206659,I2507,I206192,I206721,);
not I_12012 (I206729,I206721);
nor I_12013 (I206178,I206729,I206441);
not I_12014 (I206787,I2514);
DFFARX1 I_12015 (I562529,I2507,I206787,I206813,);
DFFARX1 I_12016 (I206813,I2507,I206787,I206830,);
not I_12017 (I206779,I206830);
not I_12018 (I206852,I206813);
DFFARX1 I_12019 (I562520,I2507,I206787,I206878,);
not I_12020 (I206886,I206878);
and I_12021 (I206903,I206852,I562538);
not I_12022 (I206920,I562535);
nand I_12023 (I206937,I206920,I562538);
not I_12024 (I206954,I562514);
nor I_12025 (I206971,I206954,I562517);
nand I_12026 (I206988,I206971,I562526);
nor I_12027 (I207005,I206988,I206937);
DFFARX1 I_12028 (I207005,I2507,I206787,I206755,);
not I_12029 (I207036,I206988);
not I_12030 (I207053,I562517);
nand I_12031 (I207070,I207053,I562538);
nor I_12032 (I207087,I562517,I562535);
nand I_12033 (I206767,I206903,I207087);
nand I_12034 (I206761,I206852,I562517);
nand I_12035 (I207132,I206954,I562532);
DFFARX1 I_12036 (I207132,I2507,I206787,I206776,);
DFFARX1 I_12037 (I207132,I2507,I206787,I206770,);
not I_12038 (I207177,I562532);
nor I_12039 (I207194,I207177,I562514);
and I_12040 (I207211,I207194,I562523);
or I_12041 (I207228,I207211,I562517);
DFFARX1 I_12042 (I207228,I2507,I206787,I207254,);
nand I_12043 (I207262,I207254,I206920);
nor I_12044 (I206764,I207262,I207070);
nor I_12045 (I206758,I207254,I206886);
DFFARX1 I_12046 (I207254,I2507,I206787,I207316,);
not I_12047 (I207324,I207316);
nor I_12048 (I206773,I207324,I207036);
not I_12049 (I207382,I2514);
DFFARX1 I_12050 (I1352933,I2507,I207382,I207408,);
DFFARX1 I_12051 (I207408,I2507,I207382,I207425,);
not I_12052 (I207374,I207425);
not I_12053 (I207447,I207408);
DFFARX1 I_12054 (I1352924,I2507,I207382,I207473,);
not I_12055 (I207481,I207473);
and I_12056 (I207498,I207447,I1352918);
not I_12057 (I207515,I1352912);
nand I_12058 (I207532,I207515,I1352918);
not I_12059 (I207549,I1352939);
nor I_12060 (I207566,I207549,I1352912);
nand I_12061 (I207583,I207566,I1352936);
nor I_12062 (I207600,I207583,I207532);
DFFARX1 I_12063 (I207600,I2507,I207382,I207350,);
not I_12064 (I207631,I207583);
not I_12065 (I207648,I1352912);
nand I_12066 (I207665,I207648,I1352918);
nor I_12067 (I207682,I1352912,I1352912);
nand I_12068 (I207362,I207498,I207682);
nand I_12069 (I207356,I207447,I1352912);
nand I_12070 (I207727,I207549,I1352921);
DFFARX1 I_12071 (I207727,I2507,I207382,I207371,);
DFFARX1 I_12072 (I207727,I2507,I207382,I207365,);
not I_12073 (I207772,I1352921);
nor I_12074 (I207789,I207772,I1352927);
and I_12075 (I207806,I207789,I1352930);
or I_12076 (I207823,I207806,I1352915);
DFFARX1 I_12077 (I207823,I2507,I207382,I207849,);
nand I_12078 (I207857,I207849,I207515);
nor I_12079 (I207359,I207857,I207665);
nor I_12080 (I207353,I207849,I207481);
DFFARX1 I_12081 (I207849,I2507,I207382,I207911,);
not I_12082 (I207919,I207911);
nor I_12083 (I207368,I207919,I207631);
not I_12084 (I207977,I2514);
DFFARX1 I_12085 (I1267473,I2507,I207977,I208003,);
DFFARX1 I_12086 (I208003,I2507,I207977,I208020,);
not I_12087 (I207969,I208020);
not I_12088 (I208042,I208003);
DFFARX1 I_12089 (I1267485,I2507,I207977,I208068,);
not I_12090 (I208076,I208068);
and I_12091 (I208093,I208042,I1267479);
not I_12092 (I208110,I1267491);
nand I_12093 (I208127,I208110,I1267479);
not I_12094 (I208144,I1267476);
nor I_12095 (I208161,I208144,I1267488);
nand I_12096 (I208178,I208161,I1267470);
nor I_12097 (I208195,I208178,I208127);
DFFARX1 I_12098 (I208195,I2507,I207977,I207945,);
not I_12099 (I208226,I208178);
not I_12100 (I208243,I1267488);
nand I_12101 (I208260,I208243,I1267479);
nor I_12102 (I208277,I1267488,I1267491);
nand I_12103 (I207957,I208093,I208277);
nand I_12104 (I207951,I208042,I1267488);
nand I_12105 (I208322,I208144,I1267482);
DFFARX1 I_12106 (I208322,I2507,I207977,I207966,);
DFFARX1 I_12107 (I208322,I2507,I207977,I207960,);
not I_12108 (I208367,I1267482);
nor I_12109 (I208384,I208367,I1267473);
and I_12110 (I208401,I208384,I1267470);
or I_12111 (I208418,I208401,I1267494);
DFFARX1 I_12112 (I208418,I2507,I207977,I208444,);
nand I_12113 (I208452,I208444,I208110);
nor I_12114 (I207954,I208452,I208260);
nor I_12115 (I207948,I208444,I208076);
DFFARX1 I_12116 (I208444,I2507,I207977,I208506,);
not I_12117 (I208514,I208506);
nor I_12118 (I207963,I208514,I208226);
not I_12119 (I208572,I2514);
DFFARX1 I_12120 (I1269785,I2507,I208572,I208598,);
DFFARX1 I_12121 (I208598,I2507,I208572,I208615,);
not I_12122 (I208564,I208615);
not I_12123 (I208637,I208598);
DFFARX1 I_12124 (I1269797,I2507,I208572,I208663,);
not I_12125 (I208671,I208663);
and I_12126 (I208688,I208637,I1269791);
not I_12127 (I208705,I1269803);
nand I_12128 (I208722,I208705,I1269791);
not I_12129 (I208739,I1269788);
nor I_12130 (I208756,I208739,I1269800);
nand I_12131 (I208773,I208756,I1269782);
nor I_12132 (I208790,I208773,I208722);
DFFARX1 I_12133 (I208790,I2507,I208572,I208540,);
not I_12134 (I208821,I208773);
not I_12135 (I208838,I1269800);
nand I_12136 (I208855,I208838,I1269791);
nor I_12137 (I208872,I1269800,I1269803);
nand I_12138 (I208552,I208688,I208872);
nand I_12139 (I208546,I208637,I1269800);
nand I_12140 (I208917,I208739,I1269794);
DFFARX1 I_12141 (I208917,I2507,I208572,I208561,);
DFFARX1 I_12142 (I208917,I2507,I208572,I208555,);
not I_12143 (I208962,I1269794);
nor I_12144 (I208979,I208962,I1269785);
and I_12145 (I208996,I208979,I1269782);
or I_12146 (I209013,I208996,I1269806);
DFFARX1 I_12147 (I209013,I2507,I208572,I209039,);
nand I_12148 (I209047,I209039,I208705);
nor I_12149 (I208549,I209047,I208855);
nor I_12150 (I208543,I209039,I208671);
DFFARX1 I_12151 (I209039,I2507,I208572,I209101,);
not I_12152 (I209109,I209101);
nor I_12153 (I208558,I209109,I208821);
not I_12154 (I209167,I2514);
DFFARX1 I_12155 (I874453,I2507,I209167,I209193,);
DFFARX1 I_12156 (I209193,I2507,I209167,I209210,);
not I_12157 (I209159,I209210);
not I_12158 (I209232,I209193);
DFFARX1 I_12159 (I874447,I2507,I209167,I209258,);
not I_12160 (I209266,I209258);
and I_12161 (I209283,I209232,I874465);
not I_12162 (I209300,I874453);
nand I_12163 (I209317,I209300,I874465);
not I_12164 (I209334,I874447);
nor I_12165 (I209351,I209334,I874459);
nand I_12166 (I209368,I209351,I874450);
nor I_12167 (I209385,I209368,I209317);
DFFARX1 I_12168 (I209385,I2507,I209167,I209135,);
not I_12169 (I209416,I209368);
not I_12170 (I209433,I874459);
nand I_12171 (I209450,I209433,I874465);
nor I_12172 (I209467,I874459,I874453);
nand I_12173 (I209147,I209283,I209467);
nand I_12174 (I209141,I209232,I874459);
nand I_12175 (I209512,I209334,I874462);
DFFARX1 I_12176 (I209512,I2507,I209167,I209156,);
DFFARX1 I_12177 (I209512,I2507,I209167,I209150,);
not I_12178 (I209557,I874462);
nor I_12179 (I209574,I209557,I874468);
and I_12180 (I209591,I209574,I874450);
or I_12181 (I209608,I209591,I874456);
DFFARX1 I_12182 (I209608,I2507,I209167,I209634,);
nand I_12183 (I209642,I209634,I209300);
nor I_12184 (I209144,I209642,I209450);
nor I_12185 (I209138,I209634,I209266);
DFFARX1 I_12186 (I209634,I2507,I209167,I209696,);
not I_12187 (I209704,I209696);
nor I_12188 (I209153,I209704,I209416);
not I_12189 (I209762,I2514);
DFFARX1 I_12190 (I548657,I2507,I209762,I209788,);
DFFARX1 I_12191 (I209788,I2507,I209762,I209805,);
not I_12192 (I209754,I209805);
not I_12193 (I209827,I209788);
DFFARX1 I_12194 (I548648,I2507,I209762,I209853,);
not I_12195 (I209861,I209853);
and I_12196 (I209878,I209827,I548666);
not I_12197 (I209895,I548663);
nand I_12198 (I209912,I209895,I548666);
not I_12199 (I209929,I548642);
nor I_12200 (I209946,I209929,I548645);
nand I_12201 (I209963,I209946,I548654);
nor I_12202 (I209980,I209963,I209912);
DFFARX1 I_12203 (I209980,I2507,I209762,I209730,);
not I_12204 (I210011,I209963);
not I_12205 (I210028,I548645);
nand I_12206 (I210045,I210028,I548666);
nor I_12207 (I210062,I548645,I548663);
nand I_12208 (I209742,I209878,I210062);
nand I_12209 (I209736,I209827,I548645);
nand I_12210 (I210107,I209929,I548660);
DFFARX1 I_12211 (I210107,I2507,I209762,I209751,);
DFFARX1 I_12212 (I210107,I2507,I209762,I209745,);
not I_12213 (I210152,I548660);
nor I_12214 (I210169,I210152,I548642);
and I_12215 (I210186,I210169,I548651);
or I_12216 (I210203,I210186,I548645);
DFFARX1 I_12217 (I210203,I2507,I209762,I210229,);
nand I_12218 (I210237,I210229,I209895);
nor I_12219 (I209739,I210237,I210045);
nor I_12220 (I209733,I210229,I209861);
DFFARX1 I_12221 (I210229,I2507,I209762,I210291,);
not I_12222 (I210299,I210291);
nor I_12223 (I209748,I210299,I210011);
not I_12224 (I210357,I2514);
DFFARX1 I_12225 (I1114436,I2507,I210357,I210383,);
DFFARX1 I_12226 (I210383,I2507,I210357,I210400,);
not I_12227 (I210349,I210400);
not I_12228 (I210422,I210383);
DFFARX1 I_12229 (I1114436,I2507,I210357,I210448,);
not I_12230 (I210456,I210448);
and I_12231 (I210473,I210422,I1114439);
not I_12232 (I210490,I1114451);
nand I_12233 (I210507,I210490,I1114439);
not I_12234 (I210524,I1114457);
nor I_12235 (I210541,I210524,I1114448);
nand I_12236 (I210558,I210541,I1114454);
nor I_12237 (I210575,I210558,I210507);
DFFARX1 I_12238 (I210575,I2507,I210357,I210325,);
not I_12239 (I210606,I210558);
not I_12240 (I210623,I1114448);
nand I_12241 (I210640,I210623,I1114439);
nor I_12242 (I210657,I1114448,I1114451);
nand I_12243 (I210337,I210473,I210657);
nand I_12244 (I210331,I210422,I1114448);
nand I_12245 (I210702,I210524,I1114445);
DFFARX1 I_12246 (I210702,I2507,I210357,I210346,);
DFFARX1 I_12247 (I210702,I2507,I210357,I210340,);
not I_12248 (I210747,I1114445);
nor I_12249 (I210764,I210747,I1114442);
and I_12250 (I210781,I210764,I1114460);
or I_12251 (I210798,I210781,I1114439);
DFFARX1 I_12252 (I210798,I2507,I210357,I210824,);
nand I_12253 (I210832,I210824,I210490);
nor I_12254 (I210334,I210832,I210640);
nor I_12255 (I210328,I210824,I210456);
DFFARX1 I_12256 (I210824,I2507,I210357,I210886,);
not I_12257 (I210894,I210886);
nor I_12258 (I210343,I210894,I210606);
not I_12259 (I210952,I2514);
DFFARX1 I_12260 (I1086692,I2507,I210952,I210978,);
DFFARX1 I_12261 (I210978,I2507,I210952,I210995,);
not I_12262 (I210944,I210995);
not I_12263 (I211017,I210978);
DFFARX1 I_12264 (I1086692,I2507,I210952,I211043,);
not I_12265 (I211051,I211043);
and I_12266 (I211068,I211017,I1086695);
not I_12267 (I211085,I1086707);
nand I_12268 (I211102,I211085,I1086695);
not I_12269 (I211119,I1086713);
nor I_12270 (I211136,I211119,I1086704);
nand I_12271 (I211153,I211136,I1086710);
nor I_12272 (I211170,I211153,I211102);
DFFARX1 I_12273 (I211170,I2507,I210952,I210920,);
not I_12274 (I211201,I211153);
not I_12275 (I211218,I1086704);
nand I_12276 (I211235,I211218,I1086695);
nor I_12277 (I211252,I1086704,I1086707);
nand I_12278 (I210932,I211068,I211252);
nand I_12279 (I210926,I211017,I1086704);
nand I_12280 (I211297,I211119,I1086701);
DFFARX1 I_12281 (I211297,I2507,I210952,I210941,);
DFFARX1 I_12282 (I211297,I2507,I210952,I210935,);
not I_12283 (I211342,I1086701);
nor I_12284 (I211359,I211342,I1086698);
and I_12285 (I211376,I211359,I1086716);
or I_12286 (I211393,I211376,I1086695);
DFFARX1 I_12287 (I211393,I2507,I210952,I211419,);
nand I_12288 (I211427,I211419,I211085);
nor I_12289 (I210929,I211427,I211235);
nor I_12290 (I210923,I211419,I211051);
DFFARX1 I_12291 (I211419,I2507,I210952,I211481,);
not I_12292 (I211489,I211481);
nor I_12293 (I210938,I211489,I211201);
not I_12294 (I211547,I2514);
DFFARX1 I_12295 (I648648,I2507,I211547,I211573,);
DFFARX1 I_12296 (I211573,I2507,I211547,I211590,);
not I_12297 (I211539,I211590);
not I_12298 (I211612,I211573);
DFFARX1 I_12299 (I648645,I2507,I211547,I211638,);
not I_12300 (I211646,I211638);
and I_12301 (I211663,I211612,I648651);
not I_12302 (I211680,I648636);
nand I_12303 (I211697,I211680,I648651);
not I_12304 (I211714,I648639);
nor I_12305 (I211731,I211714,I648660);
nand I_12306 (I211748,I211731,I648657);
nor I_12307 (I211765,I211748,I211697);
DFFARX1 I_12308 (I211765,I2507,I211547,I211515,);
not I_12309 (I211796,I211748);
not I_12310 (I211813,I648660);
nand I_12311 (I211830,I211813,I648651);
nor I_12312 (I211847,I648660,I648636);
nand I_12313 (I211527,I211663,I211847);
nand I_12314 (I211521,I211612,I648660);
nand I_12315 (I211892,I211714,I648636);
DFFARX1 I_12316 (I211892,I2507,I211547,I211536,);
DFFARX1 I_12317 (I211892,I2507,I211547,I211530,);
not I_12318 (I211937,I648636);
nor I_12319 (I211954,I211937,I648642);
and I_12320 (I211971,I211954,I648654);
or I_12321 (I211988,I211971,I648639);
DFFARX1 I_12322 (I211988,I2507,I211547,I212014,);
nand I_12323 (I212022,I212014,I211680);
nor I_12324 (I211524,I212022,I211830);
nor I_12325 (I211518,I212014,I211646);
DFFARX1 I_12326 (I212014,I2507,I211547,I212076,);
not I_12327 (I212084,I212076);
nor I_12328 (I211533,I212084,I211796);
not I_12329 (I212142,I2514);
DFFARX1 I_12330 (I447431,I2507,I212142,I212168,);
DFFARX1 I_12331 (I212168,I2507,I212142,I212185,);
not I_12332 (I212134,I212185);
not I_12333 (I212207,I212168);
DFFARX1 I_12334 (I447419,I2507,I212142,I212233,);
not I_12335 (I212241,I212233);
and I_12336 (I212258,I212207,I447428);
not I_12337 (I212275,I447425);
nand I_12338 (I212292,I212275,I447428);
not I_12339 (I212309,I447416);
nor I_12340 (I212326,I212309,I447422);
nand I_12341 (I212343,I212326,I447407);
nor I_12342 (I212360,I212343,I212292);
DFFARX1 I_12343 (I212360,I2507,I212142,I212110,);
not I_12344 (I212391,I212343);
not I_12345 (I212408,I447422);
nand I_12346 (I212425,I212408,I447428);
nor I_12347 (I212442,I447422,I447425);
nand I_12348 (I212122,I212258,I212442);
nand I_12349 (I212116,I212207,I447422);
nand I_12350 (I212487,I212309,I447407);
DFFARX1 I_12351 (I212487,I2507,I212142,I212131,);
DFFARX1 I_12352 (I212487,I2507,I212142,I212125,);
not I_12353 (I212532,I447407);
nor I_12354 (I212549,I212532,I447413);
and I_12355 (I212566,I212549,I447410);
or I_12356 (I212583,I212566,I447434);
DFFARX1 I_12357 (I212583,I2507,I212142,I212609,);
nand I_12358 (I212617,I212609,I212275);
nor I_12359 (I212119,I212617,I212425);
nor I_12360 (I212113,I212609,I212241);
DFFARX1 I_12361 (I212609,I2507,I212142,I212671,);
not I_12362 (I212679,I212671);
nor I_12363 (I212128,I212679,I212391);
not I_12364 (I212737,I2514);
DFFARX1 I_12365 (I886294,I2507,I212737,I212763,);
DFFARX1 I_12366 (I212763,I2507,I212737,I212780,);
not I_12367 (I212729,I212780);
not I_12368 (I212802,I212763);
DFFARX1 I_12369 (I886303,I2507,I212737,I212828,);
not I_12370 (I212836,I212828);
and I_12371 (I212853,I212802,I886291);
not I_12372 (I212870,I886282);
nand I_12373 (I212887,I212870,I886291);
not I_12374 (I212904,I886288);
nor I_12375 (I212921,I212904,I886306);
nand I_12376 (I212938,I212921,I886279);
nor I_12377 (I212955,I212938,I212887);
DFFARX1 I_12378 (I212955,I2507,I212737,I212705,);
not I_12379 (I212986,I212938);
not I_12380 (I213003,I886306);
nand I_12381 (I213020,I213003,I886291);
nor I_12382 (I213037,I886306,I886282);
nand I_12383 (I212717,I212853,I213037);
nand I_12384 (I212711,I212802,I886306);
nand I_12385 (I213082,I212904,I886285);
DFFARX1 I_12386 (I213082,I2507,I212737,I212726,);
DFFARX1 I_12387 (I213082,I2507,I212737,I212720,);
not I_12388 (I213127,I886285);
nor I_12389 (I213144,I213127,I886297);
and I_12390 (I213161,I213144,I886279);
or I_12391 (I213178,I213161,I886300);
DFFARX1 I_12392 (I213178,I2507,I212737,I213204,);
nand I_12393 (I213212,I213204,I212870);
nor I_12394 (I212714,I213212,I213020);
nor I_12395 (I212708,I213204,I212836);
DFFARX1 I_12396 (I213204,I2507,I212737,I213266,);
not I_12397 (I213274,I213266);
nor I_12398 (I212723,I213274,I212986);
not I_12399 (I213332,I2514);
DFFARX1 I_12400 (I88597,I2507,I213332,I213358,);
DFFARX1 I_12401 (I213358,I2507,I213332,I213375,);
not I_12402 (I213324,I213375);
not I_12403 (I213397,I213358);
DFFARX1 I_12404 (I88591,I2507,I213332,I213423,);
not I_12405 (I213431,I213423);
and I_12406 (I213448,I213397,I88588);
not I_12407 (I213465,I88609);
nand I_12408 (I213482,I213465,I88588);
not I_12409 (I213499,I88603);
nor I_12410 (I213516,I213499,I88594);
nand I_12411 (I213533,I213516,I88600);
nor I_12412 (I213550,I213533,I213482);
DFFARX1 I_12413 (I213550,I2507,I213332,I213300,);
not I_12414 (I213581,I213533);
not I_12415 (I213598,I88594);
nand I_12416 (I213615,I213598,I88588);
nor I_12417 (I213632,I88594,I88609);
nand I_12418 (I213312,I213448,I213632);
nand I_12419 (I213306,I213397,I88594);
nand I_12420 (I213677,I213499,I88588);
DFFARX1 I_12421 (I213677,I2507,I213332,I213321,);
DFFARX1 I_12422 (I213677,I2507,I213332,I213315,);
not I_12423 (I213722,I88588);
nor I_12424 (I213739,I213722,I88606);
and I_12425 (I213756,I213739,I88612);
or I_12426 (I213773,I213756,I88591);
DFFARX1 I_12427 (I213773,I2507,I213332,I213799,);
nand I_12428 (I213807,I213799,I213465);
nor I_12429 (I213309,I213807,I213615);
nor I_12430 (I213303,I213799,I213431);
DFFARX1 I_12431 (I213799,I2507,I213332,I213861,);
not I_12432 (I213869,I213861);
nor I_12433 (I213318,I213869,I213581);
not I_12434 (I213927,I2514);
DFFARX1 I_12435 (I1334488,I2507,I213927,I213953,);
DFFARX1 I_12436 (I213953,I2507,I213927,I213970,);
not I_12437 (I213919,I213970);
not I_12438 (I213992,I213953);
DFFARX1 I_12439 (I1334479,I2507,I213927,I214018,);
not I_12440 (I214026,I214018);
and I_12441 (I214043,I213992,I1334473);
not I_12442 (I214060,I1334467);
nand I_12443 (I214077,I214060,I1334473);
not I_12444 (I214094,I1334494);
nor I_12445 (I214111,I214094,I1334467);
nand I_12446 (I214128,I214111,I1334491);
nor I_12447 (I214145,I214128,I214077);
DFFARX1 I_12448 (I214145,I2507,I213927,I213895,);
not I_12449 (I214176,I214128);
not I_12450 (I214193,I1334467);
nand I_12451 (I214210,I214193,I1334473);
nor I_12452 (I214227,I1334467,I1334467);
nand I_12453 (I213907,I214043,I214227);
nand I_12454 (I213901,I213992,I1334467);
nand I_12455 (I214272,I214094,I1334476);
DFFARX1 I_12456 (I214272,I2507,I213927,I213916,);
DFFARX1 I_12457 (I214272,I2507,I213927,I213910,);
not I_12458 (I214317,I1334476);
nor I_12459 (I214334,I214317,I1334482);
and I_12460 (I214351,I214334,I1334485);
or I_12461 (I214368,I214351,I1334470);
DFFARX1 I_12462 (I214368,I2507,I213927,I214394,);
nand I_12463 (I214402,I214394,I214060);
nor I_12464 (I213904,I214402,I214210);
nor I_12465 (I213898,I214394,I214026);
DFFARX1 I_12466 (I214394,I2507,I213927,I214456,);
not I_12467 (I214464,I214456);
nor I_12468 (I213913,I214464,I214176);
not I_12469 (I214522,I2514);
DFFARX1 I_12470 (I522066,I2507,I214522,I214548,);
DFFARX1 I_12471 (I214548,I2507,I214522,I214565,);
not I_12472 (I214514,I214565);
not I_12473 (I214587,I214548);
DFFARX1 I_12474 (I522060,I2507,I214522,I214613,);
not I_12475 (I214621,I214613);
and I_12476 (I214638,I214587,I522075);
not I_12477 (I214655,I522072);
nand I_12478 (I214672,I214655,I522075);
not I_12479 (I214689,I522063);
nor I_12480 (I214706,I214689,I522054);
nand I_12481 (I214723,I214706,I522057);
nor I_12482 (I214740,I214723,I214672);
DFFARX1 I_12483 (I214740,I2507,I214522,I214490,);
not I_12484 (I214771,I214723);
not I_12485 (I214788,I522054);
nand I_12486 (I214805,I214788,I522075);
nor I_12487 (I214822,I522054,I522072);
nand I_12488 (I214502,I214638,I214822);
nand I_12489 (I214496,I214587,I522054);
nand I_12490 (I214867,I214689,I522078);
DFFARX1 I_12491 (I214867,I2507,I214522,I214511,);
DFFARX1 I_12492 (I214867,I2507,I214522,I214505,);
not I_12493 (I214912,I522078);
nor I_12494 (I214929,I214912,I522069);
and I_12495 (I214946,I214929,I522054);
or I_12496 (I214963,I214946,I522057);
DFFARX1 I_12497 (I214963,I2507,I214522,I214989,);
nand I_12498 (I214997,I214989,I214655);
nor I_12499 (I214499,I214997,I214805);
nor I_12500 (I214493,I214989,I214621);
DFFARX1 I_12501 (I214989,I2507,I214522,I215051,);
not I_12502 (I215059,I215051);
nor I_12503 (I214508,I215059,I214771);
not I_12504 (I215117,I2514);
DFFARX1 I_12505 (I120744,I2507,I215117,I215143,);
DFFARX1 I_12506 (I215143,I2507,I215117,I215160,);
not I_12507 (I215109,I215160);
not I_12508 (I215182,I215143);
DFFARX1 I_12509 (I120738,I2507,I215117,I215208,);
not I_12510 (I215216,I215208);
and I_12511 (I215233,I215182,I120735);
not I_12512 (I215250,I120756);
nand I_12513 (I215267,I215250,I120735);
not I_12514 (I215284,I120750);
nor I_12515 (I215301,I215284,I120741);
nand I_12516 (I215318,I215301,I120747);
nor I_12517 (I215335,I215318,I215267);
DFFARX1 I_12518 (I215335,I2507,I215117,I215085,);
not I_12519 (I215366,I215318);
not I_12520 (I215383,I120741);
nand I_12521 (I215400,I215383,I120735);
nor I_12522 (I215417,I120741,I120756);
nand I_12523 (I215097,I215233,I215417);
nand I_12524 (I215091,I215182,I120741);
nand I_12525 (I215462,I215284,I120735);
DFFARX1 I_12526 (I215462,I2507,I215117,I215106,);
DFFARX1 I_12527 (I215462,I2507,I215117,I215100,);
not I_12528 (I215507,I120735);
nor I_12529 (I215524,I215507,I120753);
and I_12530 (I215541,I215524,I120759);
or I_12531 (I215558,I215541,I120738);
DFFARX1 I_12532 (I215558,I2507,I215117,I215584,);
nand I_12533 (I215592,I215584,I215250);
nor I_12534 (I215094,I215592,I215400);
nor I_12535 (I215088,I215584,I215216);
DFFARX1 I_12536 (I215584,I2507,I215117,I215646,);
not I_12537 (I215654,I215646);
nor I_12538 (I215103,I215654,I215366);
not I_12539 (I215712,I2514);
DFFARX1 I_12540 (I1044926,I2507,I215712,I215738,);
DFFARX1 I_12541 (I215738,I2507,I215712,I215755,);
not I_12542 (I215704,I215755);
not I_12543 (I215777,I215738);
DFFARX1 I_12544 (I1044935,I2507,I215712,I215803,);
not I_12545 (I215811,I215803);
and I_12546 (I215828,I215777,I1044929);
not I_12547 (I215845,I1044923);
nand I_12548 (I215862,I215845,I1044929);
not I_12549 (I215879,I1044938);
nor I_12550 (I215896,I215879,I1044926);
nand I_12551 (I215913,I215896,I1044932);
nor I_12552 (I215930,I215913,I215862);
DFFARX1 I_12553 (I215930,I2507,I215712,I215680,);
not I_12554 (I215961,I215913);
not I_12555 (I215978,I1044926);
nand I_12556 (I215995,I215978,I1044929);
nor I_12557 (I216012,I1044926,I1044923);
nand I_12558 (I215692,I215828,I216012);
nand I_12559 (I215686,I215777,I1044926);
nand I_12560 (I216057,I215879,I1044929);
DFFARX1 I_12561 (I216057,I2507,I215712,I215701,);
DFFARX1 I_12562 (I216057,I2507,I215712,I215695,);
not I_12563 (I216102,I1044929);
nor I_12564 (I216119,I216102,I1044944);
and I_12565 (I216136,I216119,I1044941);
or I_12566 (I216153,I216136,I1044923);
DFFARX1 I_12567 (I216153,I2507,I215712,I216179,);
nand I_12568 (I216187,I216179,I215845);
nor I_12569 (I215689,I216187,I215995);
nor I_12570 (I215683,I216179,I215811);
DFFARX1 I_12571 (I216179,I2507,I215712,I216241,);
not I_12572 (I216249,I216241);
nor I_12573 (I215698,I216249,I215961);
not I_12574 (I216307,I2514);
DFFARX1 I_12575 (I696044,I2507,I216307,I216333,);
DFFARX1 I_12576 (I216333,I2507,I216307,I216350,);
not I_12577 (I216299,I216350);
not I_12578 (I216372,I216333);
DFFARX1 I_12579 (I696041,I2507,I216307,I216398,);
not I_12580 (I216406,I216398);
and I_12581 (I216423,I216372,I696047);
not I_12582 (I216440,I696032);
nand I_12583 (I216457,I216440,I696047);
not I_12584 (I216474,I696035);
nor I_12585 (I216491,I216474,I696056);
nand I_12586 (I216508,I216491,I696053);
nor I_12587 (I216525,I216508,I216457);
DFFARX1 I_12588 (I216525,I2507,I216307,I216275,);
not I_12589 (I216556,I216508);
not I_12590 (I216573,I696056);
nand I_12591 (I216590,I216573,I696047);
nor I_12592 (I216607,I696056,I696032);
nand I_12593 (I216287,I216423,I216607);
nand I_12594 (I216281,I216372,I696056);
nand I_12595 (I216652,I216474,I696032);
DFFARX1 I_12596 (I216652,I2507,I216307,I216296,);
DFFARX1 I_12597 (I216652,I2507,I216307,I216290,);
not I_12598 (I216697,I696032);
nor I_12599 (I216714,I216697,I696038);
and I_12600 (I216731,I216714,I696050);
or I_12601 (I216748,I216731,I696035);
DFFARX1 I_12602 (I216748,I2507,I216307,I216774,);
nand I_12603 (I216782,I216774,I216440);
nor I_12604 (I216284,I216782,I216590);
nor I_12605 (I216278,I216774,I216406);
DFFARX1 I_12606 (I216774,I2507,I216307,I216836,);
not I_12607 (I216844,I216836);
nor I_12608 (I216293,I216844,I216556);
not I_12609 (I216902,I2514);
DFFARX1 I_12610 (I1198824,I2507,I216902,I216928,);
DFFARX1 I_12611 (I216928,I2507,I216902,I216945,);
not I_12612 (I216894,I216945);
not I_12613 (I216967,I216928);
DFFARX1 I_12614 (I1198824,I2507,I216902,I216993,);
not I_12615 (I217001,I216993);
and I_12616 (I217018,I216967,I1198827);
not I_12617 (I217035,I1198839);
nand I_12618 (I217052,I217035,I1198827);
not I_12619 (I217069,I1198845);
nor I_12620 (I217086,I217069,I1198836);
nand I_12621 (I217103,I217086,I1198842);
nor I_12622 (I217120,I217103,I217052);
DFFARX1 I_12623 (I217120,I2507,I216902,I216870,);
not I_12624 (I217151,I217103);
not I_12625 (I217168,I1198836);
nand I_12626 (I217185,I217168,I1198827);
nor I_12627 (I217202,I1198836,I1198839);
nand I_12628 (I216882,I217018,I217202);
nand I_12629 (I216876,I216967,I1198836);
nand I_12630 (I217247,I217069,I1198833);
DFFARX1 I_12631 (I217247,I2507,I216902,I216891,);
DFFARX1 I_12632 (I217247,I2507,I216902,I216885,);
not I_12633 (I217292,I1198833);
nor I_12634 (I217309,I217292,I1198830);
and I_12635 (I217326,I217309,I1198848);
or I_12636 (I217343,I217326,I1198827);
DFFARX1 I_12637 (I217343,I2507,I216902,I217369,);
nand I_12638 (I217377,I217369,I217035);
nor I_12639 (I216879,I217377,I217185);
nor I_12640 (I216873,I217369,I217001);
DFFARX1 I_12641 (I217369,I2507,I216902,I217431,);
not I_12642 (I217439,I217431);
nor I_12643 (I216888,I217439,I217151);
not I_12644 (I217497,I2514);
DFFARX1 I_12645 (I54342,I2507,I217497,I217523,);
DFFARX1 I_12646 (I217523,I2507,I217497,I217540,);
not I_12647 (I217489,I217540);
not I_12648 (I217562,I217523);
DFFARX1 I_12649 (I54336,I2507,I217497,I217588,);
not I_12650 (I217596,I217588);
and I_12651 (I217613,I217562,I54333);
not I_12652 (I217630,I54354);
nand I_12653 (I217647,I217630,I54333);
not I_12654 (I217664,I54348);
nor I_12655 (I217681,I217664,I54339);
nand I_12656 (I217698,I217681,I54345);
nor I_12657 (I217715,I217698,I217647);
DFFARX1 I_12658 (I217715,I2507,I217497,I217465,);
not I_12659 (I217746,I217698);
not I_12660 (I217763,I54339);
nand I_12661 (I217780,I217763,I54333);
nor I_12662 (I217797,I54339,I54354);
nand I_12663 (I217477,I217613,I217797);
nand I_12664 (I217471,I217562,I54339);
nand I_12665 (I217842,I217664,I54333);
DFFARX1 I_12666 (I217842,I2507,I217497,I217486,);
DFFARX1 I_12667 (I217842,I2507,I217497,I217480,);
not I_12668 (I217887,I54333);
nor I_12669 (I217904,I217887,I54351);
and I_12670 (I217921,I217904,I54357);
or I_12671 (I217938,I217921,I54336);
DFFARX1 I_12672 (I217938,I2507,I217497,I217964,);
nand I_12673 (I217972,I217964,I217630);
nor I_12674 (I217474,I217972,I217780);
nor I_12675 (I217468,I217964,I217596);
DFFARX1 I_12676 (I217964,I2507,I217497,I218026,);
not I_12677 (I218034,I218026);
nor I_12678 (I217483,I218034,I217746);
not I_12679 (I218092,I2514);
DFFARX1 I_12680 (I852319,I2507,I218092,I218118,);
DFFARX1 I_12681 (I218118,I2507,I218092,I218135,);
not I_12682 (I218084,I218135);
not I_12683 (I218157,I218118);
DFFARX1 I_12684 (I852313,I2507,I218092,I218183,);
not I_12685 (I218191,I218183);
and I_12686 (I218208,I218157,I852331);
not I_12687 (I218225,I852319);
nand I_12688 (I218242,I218225,I852331);
not I_12689 (I218259,I852313);
nor I_12690 (I218276,I218259,I852325);
nand I_12691 (I218293,I218276,I852316);
nor I_12692 (I218310,I218293,I218242);
DFFARX1 I_12693 (I218310,I2507,I218092,I218060,);
not I_12694 (I218341,I218293);
not I_12695 (I218358,I852325);
nand I_12696 (I218375,I218358,I852331);
nor I_12697 (I218392,I852325,I852319);
nand I_12698 (I218072,I218208,I218392);
nand I_12699 (I218066,I218157,I852325);
nand I_12700 (I218437,I218259,I852328);
DFFARX1 I_12701 (I218437,I2507,I218092,I218081,);
DFFARX1 I_12702 (I218437,I2507,I218092,I218075,);
not I_12703 (I218482,I852328);
nor I_12704 (I218499,I218482,I852334);
and I_12705 (I218516,I218499,I852316);
or I_12706 (I218533,I218516,I852322);
DFFARX1 I_12707 (I218533,I2507,I218092,I218559,);
nand I_12708 (I218567,I218559,I218225);
nor I_12709 (I218069,I218567,I218375);
nor I_12710 (I218063,I218559,I218191);
DFFARX1 I_12711 (I218559,I2507,I218092,I218621,);
not I_12712 (I218629,I218621);
nor I_12713 (I218078,I218629,I218341);
not I_12714 (I218687,I2514);
DFFARX1 I_12715 (I1209620,I2507,I218687,I218713,);
DFFARX1 I_12716 (I218713,I2507,I218687,I218730,);
not I_12717 (I218679,I218730);
not I_12718 (I218752,I218713);
DFFARX1 I_12719 (I1209605,I2507,I218687,I218778,);
not I_12720 (I218786,I218778);
and I_12721 (I218803,I218752,I1209623);
not I_12722 (I218820,I1209605);
nand I_12723 (I218837,I218820,I1209623);
not I_12724 (I218854,I1209626);
nor I_12725 (I218871,I218854,I1209617);
nand I_12726 (I218888,I218871,I1209614);
nor I_12727 (I218905,I218888,I218837);
DFFARX1 I_12728 (I218905,I2507,I218687,I218655,);
not I_12729 (I218936,I218888);
not I_12730 (I218953,I1209617);
nand I_12731 (I218970,I218953,I1209623);
nor I_12732 (I218987,I1209617,I1209605);
nand I_12733 (I218667,I218803,I218987);
nand I_12734 (I218661,I218752,I1209617);
nand I_12735 (I219032,I218854,I1209611);
DFFARX1 I_12736 (I219032,I2507,I218687,I218676,);
DFFARX1 I_12737 (I219032,I2507,I218687,I218670,);
not I_12738 (I219077,I1209611);
nor I_12739 (I219094,I219077,I1209602);
and I_12740 (I219111,I219094,I1209608);
or I_12741 (I219128,I219111,I1209602);
DFFARX1 I_12742 (I219128,I2507,I218687,I219154,);
nand I_12743 (I219162,I219154,I218820);
nor I_12744 (I218664,I219162,I218970);
nor I_12745 (I218658,I219154,I218786);
DFFARX1 I_12746 (I219154,I2507,I218687,I219216,);
not I_12747 (I219224,I219216);
nor I_12748 (I218673,I219224,I218936);
not I_12749 (I219282,I2514);
DFFARX1 I_12750 (I760780,I2507,I219282,I219308,);
DFFARX1 I_12751 (I219308,I2507,I219282,I219325,);
not I_12752 (I219274,I219325);
not I_12753 (I219347,I219308);
DFFARX1 I_12754 (I760777,I2507,I219282,I219373,);
not I_12755 (I219381,I219373);
and I_12756 (I219398,I219347,I760783);
not I_12757 (I219415,I760768);
nand I_12758 (I219432,I219415,I760783);
not I_12759 (I219449,I760771);
nor I_12760 (I219466,I219449,I760792);
nand I_12761 (I219483,I219466,I760789);
nor I_12762 (I219500,I219483,I219432);
DFFARX1 I_12763 (I219500,I2507,I219282,I219250,);
not I_12764 (I219531,I219483);
not I_12765 (I219548,I760792);
nand I_12766 (I219565,I219548,I760783);
nor I_12767 (I219582,I760792,I760768);
nand I_12768 (I219262,I219398,I219582);
nand I_12769 (I219256,I219347,I760792);
nand I_12770 (I219627,I219449,I760768);
DFFARX1 I_12771 (I219627,I2507,I219282,I219271,);
DFFARX1 I_12772 (I219627,I2507,I219282,I219265,);
not I_12773 (I219672,I760768);
nor I_12774 (I219689,I219672,I760774);
and I_12775 (I219706,I219689,I760786);
or I_12776 (I219723,I219706,I760771);
DFFARX1 I_12777 (I219723,I2507,I219282,I219749,);
nand I_12778 (I219757,I219749,I219415);
nor I_12779 (I219259,I219757,I219565);
nor I_12780 (I219253,I219749,I219381);
DFFARX1 I_12781 (I219749,I2507,I219282,I219811,);
not I_12782 (I219819,I219811);
nor I_12783 (I219268,I219819,I219531);
not I_12784 (I219877,I2514);
DFFARX1 I_12785 (I488231,I2507,I219877,I219903,);
DFFARX1 I_12786 (I219903,I2507,I219877,I219920,);
not I_12787 (I219869,I219920);
not I_12788 (I219942,I219903);
DFFARX1 I_12789 (I488219,I2507,I219877,I219968,);
not I_12790 (I219976,I219968);
and I_12791 (I219993,I219942,I488228);
not I_12792 (I220010,I488225);
nand I_12793 (I220027,I220010,I488228);
not I_12794 (I220044,I488216);
nor I_12795 (I220061,I220044,I488222);
nand I_12796 (I220078,I220061,I488207);
nor I_12797 (I220095,I220078,I220027);
DFFARX1 I_12798 (I220095,I2507,I219877,I219845,);
not I_12799 (I220126,I220078);
not I_12800 (I220143,I488222);
nand I_12801 (I220160,I220143,I488228);
nor I_12802 (I220177,I488222,I488225);
nand I_12803 (I219857,I219993,I220177);
nand I_12804 (I219851,I219942,I488222);
nand I_12805 (I220222,I220044,I488207);
DFFARX1 I_12806 (I220222,I2507,I219877,I219866,);
DFFARX1 I_12807 (I220222,I2507,I219877,I219860,);
not I_12808 (I220267,I488207);
nor I_12809 (I220284,I220267,I488213);
and I_12810 (I220301,I220284,I488210);
or I_12811 (I220318,I220301,I488234);
DFFARX1 I_12812 (I220318,I2507,I219877,I220344,);
nand I_12813 (I220352,I220344,I220010);
nor I_12814 (I219854,I220352,I220160);
nor I_12815 (I219848,I220344,I219976);
DFFARX1 I_12816 (I220344,I2507,I219877,I220406,);
not I_12817 (I220414,I220406);
nor I_12818 (I219863,I220414,I220126);
not I_12819 (I220472,I2514);
DFFARX1 I_12820 (I1262849,I2507,I220472,I220498,);
DFFARX1 I_12821 (I220498,I2507,I220472,I220515,);
not I_12822 (I220464,I220515);
not I_12823 (I220537,I220498);
DFFARX1 I_12824 (I1262861,I2507,I220472,I220563,);
not I_12825 (I220571,I220563);
and I_12826 (I220588,I220537,I1262855);
not I_12827 (I220605,I1262867);
nand I_12828 (I220622,I220605,I1262855);
not I_12829 (I220639,I1262852);
nor I_12830 (I220656,I220639,I1262864);
nand I_12831 (I220673,I220656,I1262846);
nor I_12832 (I220690,I220673,I220622);
DFFARX1 I_12833 (I220690,I2507,I220472,I220440,);
not I_12834 (I220721,I220673);
not I_12835 (I220738,I1262864);
nand I_12836 (I220755,I220738,I1262855);
nor I_12837 (I220772,I1262864,I1262867);
nand I_12838 (I220452,I220588,I220772);
nand I_12839 (I220446,I220537,I1262864);
nand I_12840 (I220817,I220639,I1262858);
DFFARX1 I_12841 (I220817,I2507,I220472,I220461,);
DFFARX1 I_12842 (I220817,I2507,I220472,I220455,);
not I_12843 (I220862,I1262858);
nor I_12844 (I220879,I220862,I1262849);
and I_12845 (I220896,I220879,I1262846);
or I_12846 (I220913,I220896,I1262870);
DFFARX1 I_12847 (I220913,I2507,I220472,I220939,);
nand I_12848 (I220947,I220939,I220605);
nor I_12849 (I220449,I220947,I220755);
nor I_12850 (I220443,I220939,I220571);
DFFARX1 I_12851 (I220939,I2507,I220472,I221001,);
not I_12852 (I221009,I221001);
nor I_12853 (I220458,I221009,I220721);
not I_12854 (I221067,I2514);
DFFARX1 I_12855 (I1160676,I2507,I221067,I221093,);
DFFARX1 I_12856 (I221093,I2507,I221067,I221110,);
not I_12857 (I221059,I221110);
not I_12858 (I221132,I221093);
DFFARX1 I_12859 (I1160676,I2507,I221067,I221158,);
not I_12860 (I221166,I221158);
and I_12861 (I221183,I221132,I1160679);
not I_12862 (I221200,I1160691);
nand I_12863 (I221217,I221200,I1160679);
not I_12864 (I221234,I1160697);
nor I_12865 (I221251,I221234,I1160688);
nand I_12866 (I221268,I221251,I1160694);
nor I_12867 (I221285,I221268,I221217);
DFFARX1 I_12868 (I221285,I2507,I221067,I221035,);
not I_12869 (I221316,I221268);
not I_12870 (I221333,I1160688);
nand I_12871 (I221350,I221333,I1160679);
nor I_12872 (I221367,I1160688,I1160691);
nand I_12873 (I221047,I221183,I221367);
nand I_12874 (I221041,I221132,I1160688);
nand I_12875 (I221412,I221234,I1160685);
DFFARX1 I_12876 (I221412,I2507,I221067,I221056,);
DFFARX1 I_12877 (I221412,I2507,I221067,I221050,);
not I_12878 (I221457,I1160685);
nor I_12879 (I221474,I221457,I1160682);
and I_12880 (I221491,I221474,I1160700);
or I_12881 (I221508,I221491,I1160679);
DFFARX1 I_12882 (I221508,I2507,I221067,I221534,);
nand I_12883 (I221542,I221534,I221200);
nor I_12884 (I221044,I221542,I221350);
nor I_12885 (I221038,I221534,I221166);
DFFARX1 I_12886 (I221534,I2507,I221067,I221596,);
not I_12887 (I221604,I221596);
nor I_12888 (I221053,I221604,I221316);
not I_12889 (I221662,I2514);
DFFARX1 I_12890 (I723788,I2507,I221662,I221688,);
DFFARX1 I_12891 (I221688,I2507,I221662,I221705,);
not I_12892 (I221654,I221705);
not I_12893 (I221727,I221688);
DFFARX1 I_12894 (I723785,I2507,I221662,I221753,);
not I_12895 (I221761,I221753);
and I_12896 (I221778,I221727,I723791);
not I_12897 (I221795,I723776);
nand I_12898 (I221812,I221795,I723791);
not I_12899 (I221829,I723779);
nor I_12900 (I221846,I221829,I723800);
nand I_12901 (I221863,I221846,I723797);
nor I_12902 (I221880,I221863,I221812);
DFFARX1 I_12903 (I221880,I2507,I221662,I221630,);
not I_12904 (I221911,I221863);
not I_12905 (I221928,I723800);
nand I_12906 (I221945,I221928,I723791);
nor I_12907 (I221962,I723800,I723776);
nand I_12908 (I221642,I221778,I221962);
nand I_12909 (I221636,I221727,I723800);
nand I_12910 (I222007,I221829,I723776);
DFFARX1 I_12911 (I222007,I2507,I221662,I221651,);
DFFARX1 I_12912 (I222007,I2507,I221662,I221645,);
not I_12913 (I222052,I723776);
nor I_12914 (I222069,I222052,I723782);
and I_12915 (I222086,I222069,I723794);
or I_12916 (I222103,I222086,I723779);
DFFARX1 I_12917 (I222103,I2507,I221662,I222129,);
nand I_12918 (I222137,I222129,I221795);
nor I_12919 (I221639,I222137,I221945);
nor I_12920 (I221633,I222129,I221761);
DFFARX1 I_12921 (I222129,I2507,I221662,I222191,);
not I_12922 (I222199,I222191);
nor I_12923 (I221648,I222199,I221911);
not I_12924 (I222257,I2514);
DFFARX1 I_12925 (I871818,I2507,I222257,I222283,);
DFFARX1 I_12926 (I222283,I2507,I222257,I222300,);
not I_12927 (I222249,I222300);
not I_12928 (I222322,I222283);
DFFARX1 I_12929 (I871812,I2507,I222257,I222348,);
not I_12930 (I222356,I222348);
and I_12931 (I222373,I222322,I871830);
not I_12932 (I222390,I871818);
nand I_12933 (I222407,I222390,I871830);
not I_12934 (I222424,I871812);
nor I_12935 (I222441,I222424,I871824);
nand I_12936 (I222458,I222441,I871815);
nor I_12937 (I222475,I222458,I222407);
DFFARX1 I_12938 (I222475,I2507,I222257,I222225,);
not I_12939 (I222506,I222458);
not I_12940 (I222523,I871824);
nand I_12941 (I222540,I222523,I871830);
nor I_12942 (I222557,I871824,I871818);
nand I_12943 (I222237,I222373,I222557);
nand I_12944 (I222231,I222322,I871824);
nand I_12945 (I222602,I222424,I871827);
DFFARX1 I_12946 (I222602,I2507,I222257,I222246,);
DFFARX1 I_12947 (I222602,I2507,I222257,I222240,);
not I_12948 (I222647,I871827);
nor I_12949 (I222664,I222647,I871833);
and I_12950 (I222681,I222664,I871815);
or I_12951 (I222698,I222681,I871821);
DFFARX1 I_12952 (I222698,I2507,I222257,I222724,);
nand I_12953 (I222732,I222724,I222390);
nor I_12954 (I222234,I222732,I222540);
nor I_12955 (I222228,I222724,I222356);
DFFARX1 I_12956 (I222724,I2507,I222257,I222786,);
not I_12957 (I222794,I222786);
nor I_12958 (I222243,I222794,I222506);
not I_12959 (I222852,I2514);
DFFARX1 I_12960 (I470823,I2507,I222852,I222878,);
DFFARX1 I_12961 (I222878,I2507,I222852,I222895,);
not I_12962 (I222844,I222895);
not I_12963 (I222917,I222878);
DFFARX1 I_12964 (I470811,I2507,I222852,I222943,);
not I_12965 (I222951,I222943);
and I_12966 (I222968,I222917,I470820);
not I_12967 (I222985,I470817);
nand I_12968 (I223002,I222985,I470820);
not I_12969 (I223019,I470808);
nor I_12970 (I223036,I223019,I470814);
nand I_12971 (I223053,I223036,I470799);
nor I_12972 (I223070,I223053,I223002);
DFFARX1 I_12973 (I223070,I2507,I222852,I222820,);
not I_12974 (I223101,I223053);
not I_12975 (I223118,I470814);
nand I_12976 (I223135,I223118,I470820);
nor I_12977 (I223152,I470814,I470817);
nand I_12978 (I222832,I222968,I223152);
nand I_12979 (I222826,I222917,I470814);
nand I_12980 (I223197,I223019,I470799);
DFFARX1 I_12981 (I223197,I2507,I222852,I222841,);
DFFARX1 I_12982 (I223197,I2507,I222852,I222835,);
not I_12983 (I223242,I470799);
nor I_12984 (I223259,I223242,I470805);
and I_12985 (I223276,I223259,I470802);
or I_12986 (I223293,I223276,I470826);
DFFARX1 I_12987 (I223293,I2507,I222852,I223319,);
nand I_12988 (I223327,I223319,I222985);
nor I_12989 (I222829,I223327,I223135);
nor I_12990 (I222823,I223319,I222951);
DFFARX1 I_12991 (I223319,I2507,I222852,I223381,);
not I_12992 (I223389,I223381);
nor I_12993 (I222838,I223389,I223101);
not I_12994 (I223447,I2514);
DFFARX1 I_12995 (I1088426,I2507,I223447,I223473,);
DFFARX1 I_12996 (I223473,I2507,I223447,I223490,);
not I_12997 (I223439,I223490);
not I_12998 (I223512,I223473);
DFFARX1 I_12999 (I1088426,I2507,I223447,I223538,);
not I_13000 (I223546,I223538);
and I_13001 (I223563,I223512,I1088429);
not I_13002 (I223580,I1088441);
nand I_13003 (I223597,I223580,I1088429);
not I_13004 (I223614,I1088447);
nor I_13005 (I223631,I223614,I1088438);
nand I_13006 (I223648,I223631,I1088444);
nor I_13007 (I223665,I223648,I223597);
DFFARX1 I_13008 (I223665,I2507,I223447,I223415,);
not I_13009 (I223696,I223648);
not I_13010 (I223713,I1088438);
nand I_13011 (I223730,I223713,I1088429);
nor I_13012 (I223747,I1088438,I1088441);
nand I_13013 (I223427,I223563,I223747);
nand I_13014 (I223421,I223512,I1088438);
nand I_13015 (I223792,I223614,I1088435);
DFFARX1 I_13016 (I223792,I2507,I223447,I223436,);
DFFARX1 I_13017 (I223792,I2507,I223447,I223430,);
not I_13018 (I223837,I1088435);
nor I_13019 (I223854,I223837,I1088432);
and I_13020 (I223871,I223854,I1088450);
or I_13021 (I223888,I223871,I1088429);
DFFARX1 I_13022 (I223888,I2507,I223447,I223914,);
nand I_13023 (I223922,I223914,I223580);
nor I_13024 (I223424,I223922,I223730);
nor I_13025 (I223418,I223914,I223546);
DFFARX1 I_13026 (I223914,I2507,I223447,I223976,);
not I_13027 (I223984,I223976);
nor I_13028 (I223433,I223984,I223696);
not I_13029 (I224042,I2514);
DFFARX1 I_13030 (I850211,I2507,I224042,I224068,);
DFFARX1 I_13031 (I224068,I2507,I224042,I224085,);
not I_13032 (I224034,I224085);
not I_13033 (I224107,I224068);
DFFARX1 I_13034 (I850205,I2507,I224042,I224133,);
not I_13035 (I224141,I224133);
and I_13036 (I224158,I224107,I850223);
not I_13037 (I224175,I850211);
nand I_13038 (I224192,I224175,I850223);
not I_13039 (I224209,I850205);
nor I_13040 (I224226,I224209,I850217);
nand I_13041 (I224243,I224226,I850208);
nor I_13042 (I224260,I224243,I224192);
DFFARX1 I_13043 (I224260,I2507,I224042,I224010,);
not I_13044 (I224291,I224243);
not I_13045 (I224308,I850217);
nand I_13046 (I224325,I224308,I850223);
nor I_13047 (I224342,I850217,I850211);
nand I_13048 (I224022,I224158,I224342);
nand I_13049 (I224016,I224107,I850217);
nand I_13050 (I224387,I224209,I850220);
DFFARX1 I_13051 (I224387,I2507,I224042,I224031,);
DFFARX1 I_13052 (I224387,I2507,I224042,I224025,);
not I_13053 (I224432,I850220);
nor I_13054 (I224449,I224432,I850226);
and I_13055 (I224466,I224449,I850208);
or I_13056 (I224483,I224466,I850214);
DFFARX1 I_13057 (I224483,I2507,I224042,I224509,);
nand I_13058 (I224517,I224509,I224175);
nor I_13059 (I224019,I224517,I224325);
nor I_13060 (I224013,I224509,I224141);
DFFARX1 I_13061 (I224509,I2507,I224042,I224571,);
not I_13062 (I224579,I224571);
nor I_13063 (I224028,I224579,I224291);
not I_13064 (I224637,I2514);
DFFARX1 I_13065 (I785390,I2507,I224637,I224663,);
DFFARX1 I_13066 (I224663,I2507,I224637,I224680,);
not I_13067 (I224629,I224680);
not I_13068 (I224702,I224663);
DFFARX1 I_13069 (I785384,I2507,I224637,I224728,);
not I_13070 (I224736,I224728);
and I_13071 (I224753,I224702,I785402);
not I_13072 (I224770,I785390);
nand I_13073 (I224787,I224770,I785402);
not I_13074 (I224804,I785384);
nor I_13075 (I224821,I224804,I785396);
nand I_13076 (I224838,I224821,I785387);
nor I_13077 (I224855,I224838,I224787);
DFFARX1 I_13078 (I224855,I2507,I224637,I224605,);
not I_13079 (I224886,I224838);
not I_13080 (I224903,I785396);
nand I_13081 (I224920,I224903,I785402);
nor I_13082 (I224937,I785396,I785390);
nand I_13083 (I224617,I224753,I224937);
nand I_13084 (I224611,I224702,I785396);
nand I_13085 (I224982,I224804,I785399);
DFFARX1 I_13086 (I224982,I2507,I224637,I224626,);
DFFARX1 I_13087 (I224982,I2507,I224637,I224620,);
not I_13088 (I225027,I785399);
nor I_13089 (I225044,I225027,I785405);
and I_13090 (I225061,I225044,I785387);
or I_13091 (I225078,I225061,I785393);
DFFARX1 I_13092 (I225078,I2507,I224637,I225104,);
nand I_13093 (I225112,I225104,I224770);
nor I_13094 (I224614,I225112,I224920);
nor I_13095 (I224608,I225104,I224736);
DFFARX1 I_13096 (I225104,I2507,I224637,I225166,);
not I_13097 (I225174,I225166);
nor I_13098 (I224623,I225174,I224886);
not I_13099 (I225232,I2514);
DFFARX1 I_13100 (I361914,I2507,I225232,I225258,);
DFFARX1 I_13101 (I225258,I2507,I225232,I225275,);
not I_13102 (I225224,I225275);
not I_13103 (I225297,I225258);
DFFARX1 I_13104 (I361929,I2507,I225232,I225323,);
not I_13105 (I225331,I225323);
and I_13106 (I225348,I225297,I361926);
not I_13107 (I225365,I361914);
nand I_13108 (I225382,I225365,I361926);
not I_13109 (I225399,I361923);
nor I_13110 (I225416,I225399,I361938);
nand I_13111 (I225433,I225416,I361935);
nor I_13112 (I225450,I225433,I225382);
DFFARX1 I_13113 (I225450,I2507,I225232,I225200,);
not I_13114 (I225481,I225433);
not I_13115 (I225498,I361938);
nand I_13116 (I225515,I225498,I361926);
nor I_13117 (I225532,I361938,I361914);
nand I_13118 (I225212,I225348,I225532);
nand I_13119 (I225206,I225297,I361938);
nand I_13120 (I225577,I225399,I361932);
DFFARX1 I_13121 (I225577,I2507,I225232,I225221,);
DFFARX1 I_13122 (I225577,I2507,I225232,I225215,);
not I_13123 (I225622,I361932);
nor I_13124 (I225639,I225622,I361920);
and I_13125 (I225656,I225639,I361941);
or I_13126 (I225673,I225656,I361917);
DFFARX1 I_13127 (I225673,I2507,I225232,I225699,);
nand I_13128 (I225707,I225699,I225365);
nor I_13129 (I225209,I225707,I225515);
nor I_13130 (I225203,I225699,I225331);
DFFARX1 I_13131 (I225699,I2507,I225232,I225761,);
not I_13132 (I225769,I225761);
nor I_13133 (I225218,I225769,I225481);
not I_13134 (I225827,I2514);
DFFARX1 I_13135 (I1058948,I2507,I225827,I225853,);
DFFARX1 I_13136 (I225853,I2507,I225827,I225870,);
not I_13137 (I225819,I225870);
not I_13138 (I225892,I225853);
DFFARX1 I_13139 (I1058948,I2507,I225827,I225918,);
not I_13140 (I225926,I225918);
and I_13141 (I225943,I225892,I1058951);
not I_13142 (I225960,I1058963);
nand I_13143 (I225977,I225960,I1058951);
not I_13144 (I225994,I1058969);
nor I_13145 (I226011,I225994,I1058960);
nand I_13146 (I226028,I226011,I1058966);
nor I_13147 (I226045,I226028,I225977);
DFFARX1 I_13148 (I226045,I2507,I225827,I225795,);
not I_13149 (I226076,I226028);
not I_13150 (I226093,I1058960);
nand I_13151 (I226110,I226093,I1058951);
nor I_13152 (I226127,I1058960,I1058963);
nand I_13153 (I225807,I225943,I226127);
nand I_13154 (I225801,I225892,I1058960);
nand I_13155 (I226172,I225994,I1058957);
DFFARX1 I_13156 (I226172,I2507,I225827,I225816,);
DFFARX1 I_13157 (I226172,I2507,I225827,I225810,);
not I_13158 (I226217,I1058957);
nor I_13159 (I226234,I226217,I1058954);
and I_13160 (I226251,I226234,I1058972);
or I_13161 (I226268,I226251,I1058951);
DFFARX1 I_13162 (I226268,I2507,I225827,I226294,);
nand I_13163 (I226302,I226294,I225960);
nor I_13164 (I225804,I226302,I226110);
nor I_13165 (I225798,I226294,I225926);
DFFARX1 I_13166 (I226294,I2507,I225827,I226356,);
not I_13167 (I226364,I226356);
nor I_13168 (I225813,I226364,I226076);
not I_13169 (I226422,I2514);
DFFARX1 I_13170 (I381607,I2507,I226422,I226448,);
DFFARX1 I_13171 (I226448,I2507,I226422,I226465,);
not I_13172 (I226414,I226465);
not I_13173 (I226487,I226448);
DFFARX1 I_13174 (I381595,I2507,I226422,I226513,);
not I_13175 (I226521,I226513);
and I_13176 (I226538,I226487,I381604);
not I_13177 (I226555,I381601);
nand I_13178 (I226572,I226555,I381604);
not I_13179 (I226589,I381592);
nor I_13180 (I226606,I226589,I381598);
nand I_13181 (I226623,I226606,I381583);
nor I_13182 (I226640,I226623,I226572);
DFFARX1 I_13183 (I226640,I2507,I226422,I226390,);
not I_13184 (I226671,I226623);
not I_13185 (I226688,I381598);
nand I_13186 (I226705,I226688,I381604);
nor I_13187 (I226722,I381598,I381601);
nand I_13188 (I226402,I226538,I226722);
nand I_13189 (I226396,I226487,I381598);
nand I_13190 (I226767,I226589,I381583);
DFFARX1 I_13191 (I226767,I2507,I226422,I226411,);
DFFARX1 I_13192 (I226767,I2507,I226422,I226405,);
not I_13193 (I226812,I381583);
nor I_13194 (I226829,I226812,I381589);
and I_13195 (I226846,I226829,I381586);
or I_13196 (I226863,I226846,I381610);
DFFARX1 I_13197 (I226863,I2507,I226422,I226889,);
nand I_13198 (I226897,I226889,I226555);
nor I_13199 (I226399,I226897,I226705);
nor I_13200 (I226393,I226889,I226521);
DFFARX1 I_13201 (I226889,I2507,I226422,I226951,);
not I_13202 (I226959,I226951);
nor I_13203 (I226408,I226959,I226671);
not I_13204 (I227017,I2514);
DFFARX1 I_13205 (I628418,I2507,I227017,I227043,);
DFFARX1 I_13206 (I227043,I2507,I227017,I227060,);
not I_13207 (I227009,I227060);
not I_13208 (I227082,I227043);
DFFARX1 I_13209 (I628415,I2507,I227017,I227108,);
not I_13210 (I227116,I227108);
and I_13211 (I227133,I227082,I628421);
not I_13212 (I227150,I628406);
nand I_13213 (I227167,I227150,I628421);
not I_13214 (I227184,I628409);
nor I_13215 (I227201,I227184,I628430);
nand I_13216 (I227218,I227201,I628427);
nor I_13217 (I227235,I227218,I227167);
DFFARX1 I_13218 (I227235,I2507,I227017,I226985,);
not I_13219 (I227266,I227218);
not I_13220 (I227283,I628430);
nand I_13221 (I227300,I227283,I628421);
nor I_13222 (I227317,I628430,I628406);
nand I_13223 (I226997,I227133,I227317);
nand I_13224 (I226991,I227082,I628430);
nand I_13225 (I227362,I227184,I628406);
DFFARX1 I_13226 (I227362,I2507,I227017,I227006,);
DFFARX1 I_13227 (I227362,I2507,I227017,I227000,);
not I_13228 (I227407,I628406);
nor I_13229 (I227424,I227407,I628412);
and I_13230 (I227441,I227424,I628424);
or I_13231 (I227458,I227441,I628409);
DFFARX1 I_13232 (I227458,I2507,I227017,I227484,);
nand I_13233 (I227492,I227484,I227150);
nor I_13234 (I226994,I227492,I227300);
nor I_13235 (I226988,I227484,I227116);
DFFARX1 I_13236 (I227484,I2507,I227017,I227546,);
not I_13237 (I227554,I227546);
nor I_13238 (I227003,I227554,I227266);
not I_13239 (I227612,I2514);
DFFARX1 I_13240 (I1319613,I2507,I227612,I227638,);
DFFARX1 I_13241 (I227638,I2507,I227612,I227655,);
not I_13242 (I227604,I227655);
not I_13243 (I227677,I227638);
DFFARX1 I_13244 (I1319604,I2507,I227612,I227703,);
not I_13245 (I227711,I227703);
and I_13246 (I227728,I227677,I1319598);
not I_13247 (I227745,I1319592);
nand I_13248 (I227762,I227745,I1319598);
not I_13249 (I227779,I1319619);
nor I_13250 (I227796,I227779,I1319592);
nand I_13251 (I227813,I227796,I1319616);
nor I_13252 (I227830,I227813,I227762);
DFFARX1 I_13253 (I227830,I2507,I227612,I227580,);
not I_13254 (I227861,I227813);
not I_13255 (I227878,I1319592);
nand I_13256 (I227895,I227878,I1319598);
nor I_13257 (I227912,I1319592,I1319592);
nand I_13258 (I227592,I227728,I227912);
nand I_13259 (I227586,I227677,I1319592);
nand I_13260 (I227957,I227779,I1319601);
DFFARX1 I_13261 (I227957,I2507,I227612,I227601,);
DFFARX1 I_13262 (I227957,I2507,I227612,I227595,);
not I_13263 (I228002,I1319601);
nor I_13264 (I228019,I228002,I1319607);
and I_13265 (I228036,I228019,I1319610);
or I_13266 (I228053,I228036,I1319595);
DFFARX1 I_13267 (I228053,I2507,I227612,I228079,);
nand I_13268 (I228087,I228079,I227745);
nor I_13269 (I227589,I228087,I227895);
nor I_13270 (I227583,I228079,I227711);
DFFARX1 I_13271 (I228079,I2507,I227612,I228141,);
not I_13272 (I228149,I228141);
nor I_13273 (I227598,I228149,I227861);
not I_13274 (I228207,I2514);
DFFARX1 I_13275 (I541106,I2507,I228207,I228233,);
DFFARX1 I_13276 (I228233,I2507,I228207,I228250,);
not I_13277 (I228199,I228250);
not I_13278 (I228272,I228233);
DFFARX1 I_13279 (I541100,I2507,I228207,I228298,);
not I_13280 (I228306,I228298);
and I_13281 (I228323,I228272,I541115);
not I_13282 (I228340,I541112);
nand I_13283 (I228357,I228340,I541115);
not I_13284 (I228374,I541103);
nor I_13285 (I228391,I228374,I541094);
nand I_13286 (I228408,I228391,I541097);
nor I_13287 (I228425,I228408,I228357);
DFFARX1 I_13288 (I228425,I2507,I228207,I228175,);
not I_13289 (I228456,I228408);
not I_13290 (I228473,I541094);
nand I_13291 (I228490,I228473,I541115);
nor I_13292 (I228507,I541094,I541112);
nand I_13293 (I228187,I228323,I228507);
nand I_13294 (I228181,I228272,I541094);
nand I_13295 (I228552,I228374,I541118);
DFFARX1 I_13296 (I228552,I2507,I228207,I228196,);
DFFARX1 I_13297 (I228552,I2507,I228207,I228190,);
not I_13298 (I228597,I541118);
nor I_13299 (I228614,I228597,I541109);
and I_13300 (I228631,I228614,I541094);
or I_13301 (I228648,I228631,I541097);
DFFARX1 I_13302 (I228648,I2507,I228207,I228674,);
nand I_13303 (I228682,I228674,I228340);
nor I_13304 (I228184,I228682,I228490);
nor I_13305 (I228178,I228674,I228306);
DFFARX1 I_13306 (I228674,I2507,I228207,I228736,);
not I_13307 (I228744,I228736);
nor I_13308 (I228193,I228744,I228456);
not I_13309 (I228802,I2514);
DFFARX1 I_13310 (I715696,I2507,I228802,I228828,);
DFFARX1 I_13311 (I228828,I2507,I228802,I228845,);
not I_13312 (I228794,I228845);
not I_13313 (I228867,I228828);
DFFARX1 I_13314 (I715693,I2507,I228802,I228893,);
not I_13315 (I228901,I228893);
and I_13316 (I228918,I228867,I715699);
not I_13317 (I228935,I715684);
nand I_13318 (I228952,I228935,I715699);
not I_13319 (I228969,I715687);
nor I_13320 (I228986,I228969,I715708);
nand I_13321 (I229003,I228986,I715705);
nor I_13322 (I229020,I229003,I228952);
DFFARX1 I_13323 (I229020,I2507,I228802,I228770,);
not I_13324 (I229051,I229003);
not I_13325 (I229068,I715708);
nand I_13326 (I229085,I229068,I715699);
nor I_13327 (I229102,I715708,I715684);
nand I_13328 (I228782,I228918,I229102);
nand I_13329 (I228776,I228867,I715708);
nand I_13330 (I229147,I228969,I715684);
DFFARX1 I_13331 (I229147,I2507,I228802,I228791,);
DFFARX1 I_13332 (I229147,I2507,I228802,I228785,);
not I_13333 (I229192,I715684);
nor I_13334 (I229209,I229192,I715690);
and I_13335 (I229226,I229209,I715702);
or I_13336 (I229243,I229226,I715687);
DFFARX1 I_13337 (I229243,I2507,I228802,I229269,);
nand I_13338 (I229277,I229269,I228935);
nor I_13339 (I228779,I229277,I229085);
nor I_13340 (I228773,I229269,I228901);
DFFARX1 I_13341 (I229269,I2507,I228802,I229331,);
not I_13342 (I229339,I229331);
nor I_13343 (I228788,I229339,I229051);
not I_13344 (I229397,I2514);
DFFARX1 I_13345 (I917302,I2507,I229397,I229423,);
DFFARX1 I_13346 (I229423,I2507,I229397,I229440,);
not I_13347 (I229389,I229440);
not I_13348 (I229462,I229423);
DFFARX1 I_13349 (I917311,I2507,I229397,I229488,);
not I_13350 (I229496,I229488);
and I_13351 (I229513,I229462,I917299);
not I_13352 (I229530,I917290);
nand I_13353 (I229547,I229530,I917299);
not I_13354 (I229564,I917296);
nor I_13355 (I229581,I229564,I917314);
nand I_13356 (I229598,I229581,I917287);
nor I_13357 (I229615,I229598,I229547);
DFFARX1 I_13358 (I229615,I2507,I229397,I229365,);
not I_13359 (I229646,I229598);
not I_13360 (I229663,I917314);
nand I_13361 (I229680,I229663,I917299);
nor I_13362 (I229697,I917314,I917290);
nand I_13363 (I229377,I229513,I229697);
nand I_13364 (I229371,I229462,I917314);
nand I_13365 (I229742,I229564,I917293);
DFFARX1 I_13366 (I229742,I2507,I229397,I229386,);
DFFARX1 I_13367 (I229742,I2507,I229397,I229380,);
not I_13368 (I229787,I917293);
nor I_13369 (I229804,I229787,I917305);
and I_13370 (I229821,I229804,I917287);
or I_13371 (I229838,I229821,I917308);
DFFARX1 I_13372 (I229838,I2507,I229397,I229864,);
nand I_13373 (I229872,I229864,I229530);
nor I_13374 (I229374,I229872,I229680);
nor I_13375 (I229368,I229864,I229496);
DFFARX1 I_13376 (I229864,I2507,I229397,I229926,);
not I_13377 (I229934,I229926);
nor I_13378 (I229383,I229934,I229646);
not I_13379 (I229992,I2514);
DFFARX1 I_13380 (I919240,I2507,I229992,I230018,);
DFFARX1 I_13381 (I230018,I2507,I229992,I230035,);
not I_13382 (I229984,I230035);
not I_13383 (I230057,I230018);
DFFARX1 I_13384 (I919249,I2507,I229992,I230083,);
not I_13385 (I230091,I230083);
and I_13386 (I230108,I230057,I919237);
not I_13387 (I230125,I919228);
nand I_13388 (I230142,I230125,I919237);
not I_13389 (I230159,I919234);
nor I_13390 (I230176,I230159,I919252);
nand I_13391 (I230193,I230176,I919225);
nor I_13392 (I230210,I230193,I230142);
DFFARX1 I_13393 (I230210,I2507,I229992,I229960,);
not I_13394 (I230241,I230193);
not I_13395 (I230258,I919252);
nand I_13396 (I230275,I230258,I919237);
nor I_13397 (I230292,I919252,I919228);
nand I_13398 (I229972,I230108,I230292);
nand I_13399 (I229966,I230057,I919252);
nand I_13400 (I230337,I230159,I919231);
DFFARX1 I_13401 (I230337,I2507,I229992,I229981,);
DFFARX1 I_13402 (I230337,I2507,I229992,I229975,);
not I_13403 (I230382,I919231);
nor I_13404 (I230399,I230382,I919243);
and I_13405 (I230416,I230399,I919225);
or I_13406 (I230433,I230416,I919246);
DFFARX1 I_13407 (I230433,I2507,I229992,I230459,);
nand I_13408 (I230467,I230459,I230125);
nor I_13409 (I229969,I230467,I230275);
nor I_13410 (I229963,I230459,I230091);
DFFARX1 I_13411 (I230459,I2507,I229992,I230521,);
not I_13412 (I230529,I230521);
nor I_13413 (I229978,I230529,I230241);
not I_13414 (I230587,I2514);
DFFARX1 I_13415 (I1222676,I2507,I230587,I230613,);
DFFARX1 I_13416 (I230613,I2507,I230587,I230630,);
not I_13417 (I230579,I230630);
not I_13418 (I230652,I230613);
DFFARX1 I_13419 (I1222661,I2507,I230587,I230678,);
not I_13420 (I230686,I230678);
and I_13421 (I230703,I230652,I1222679);
not I_13422 (I230720,I1222661);
nand I_13423 (I230737,I230720,I1222679);
not I_13424 (I230754,I1222682);
nor I_13425 (I230771,I230754,I1222673);
nand I_13426 (I230788,I230771,I1222670);
nor I_13427 (I230805,I230788,I230737);
DFFARX1 I_13428 (I230805,I2507,I230587,I230555,);
not I_13429 (I230836,I230788);
not I_13430 (I230853,I1222673);
nand I_13431 (I230870,I230853,I1222679);
nor I_13432 (I230887,I1222673,I1222661);
nand I_13433 (I230567,I230703,I230887);
nand I_13434 (I230561,I230652,I1222673);
nand I_13435 (I230932,I230754,I1222667);
DFFARX1 I_13436 (I230932,I2507,I230587,I230576,);
DFFARX1 I_13437 (I230932,I2507,I230587,I230570,);
not I_13438 (I230977,I1222667);
nor I_13439 (I230994,I230977,I1222658);
and I_13440 (I231011,I230994,I1222664);
or I_13441 (I231028,I231011,I1222658);
DFFARX1 I_13442 (I231028,I2507,I230587,I231054,);
nand I_13443 (I231062,I231054,I230720);
nor I_13444 (I230564,I231062,I230870);
nor I_13445 (I230558,I231054,I230686);
DFFARX1 I_13446 (I231054,I2507,I230587,I231116,);
not I_13447 (I231124,I231116);
nor I_13448 (I230573,I231124,I230836);
not I_13449 (I231182,I2514);
DFFARX1 I_13450 (I903736,I2507,I231182,I231208,);
DFFARX1 I_13451 (I231208,I2507,I231182,I231225,);
not I_13452 (I231174,I231225);
not I_13453 (I231247,I231208);
DFFARX1 I_13454 (I903745,I2507,I231182,I231273,);
not I_13455 (I231281,I231273);
and I_13456 (I231298,I231247,I903733);
not I_13457 (I231315,I903724);
nand I_13458 (I231332,I231315,I903733);
not I_13459 (I231349,I903730);
nor I_13460 (I231366,I231349,I903748);
nand I_13461 (I231383,I231366,I903721);
nor I_13462 (I231400,I231383,I231332);
DFFARX1 I_13463 (I231400,I2507,I231182,I231150,);
not I_13464 (I231431,I231383);
not I_13465 (I231448,I903748);
nand I_13466 (I231465,I231448,I903733);
nor I_13467 (I231482,I903748,I903724);
nand I_13468 (I231162,I231298,I231482);
nand I_13469 (I231156,I231247,I903748);
nand I_13470 (I231527,I231349,I903727);
DFFARX1 I_13471 (I231527,I2507,I231182,I231171,);
DFFARX1 I_13472 (I231527,I2507,I231182,I231165,);
not I_13473 (I231572,I903727);
nor I_13474 (I231589,I231572,I903739);
and I_13475 (I231606,I231589,I903721);
or I_13476 (I231623,I231606,I903742);
DFFARX1 I_13477 (I231623,I2507,I231182,I231649,);
nand I_13478 (I231657,I231649,I231315);
nor I_13479 (I231159,I231657,I231465);
nor I_13480 (I231153,I231649,I231281);
DFFARX1 I_13481 (I231649,I2507,I231182,I231711,);
not I_13482 (I231719,I231711);
nor I_13483 (I231168,I231719,I231431);
not I_13484 (I231777,I2514);
DFFARX1 I_13485 (I596631,I2507,I231777,I231803,);
DFFARX1 I_13486 (I231803,I2507,I231777,I231820,);
not I_13487 (I231769,I231820);
not I_13488 (I231842,I231803);
DFFARX1 I_13489 (I596622,I2507,I231777,I231868,);
not I_13490 (I231876,I231868);
and I_13491 (I231893,I231842,I596640);
not I_13492 (I231910,I596637);
nand I_13493 (I231927,I231910,I596640);
not I_13494 (I231944,I596616);
nor I_13495 (I231961,I231944,I596619);
nand I_13496 (I231978,I231961,I596628);
nor I_13497 (I231995,I231978,I231927);
DFFARX1 I_13498 (I231995,I2507,I231777,I231745,);
not I_13499 (I232026,I231978);
not I_13500 (I232043,I596619);
nand I_13501 (I232060,I232043,I596640);
nor I_13502 (I232077,I596619,I596637);
nand I_13503 (I231757,I231893,I232077);
nand I_13504 (I231751,I231842,I596619);
nand I_13505 (I232122,I231944,I596634);
DFFARX1 I_13506 (I232122,I2507,I231777,I231766,);
DFFARX1 I_13507 (I232122,I2507,I231777,I231760,);
not I_13508 (I232167,I596634);
nor I_13509 (I232184,I232167,I596616);
and I_13510 (I232201,I232184,I596625);
or I_13511 (I232218,I232201,I596619);
DFFARX1 I_13512 (I232218,I2507,I231777,I232244,);
nand I_13513 (I232252,I232244,I231910);
nor I_13514 (I231754,I232252,I232060);
nor I_13515 (I231748,I232244,I231876);
DFFARX1 I_13516 (I232244,I2507,I231777,I232306,);
not I_13517 (I232314,I232306);
nor I_13518 (I231763,I232314,I232026);
not I_13519 (I232372,I2514);
DFFARX1 I_13520 (I1266895,I2507,I232372,I232398,);
DFFARX1 I_13521 (I232398,I2507,I232372,I232415,);
not I_13522 (I232364,I232415);
not I_13523 (I232437,I232398);
DFFARX1 I_13524 (I1266907,I2507,I232372,I232463,);
not I_13525 (I232471,I232463);
and I_13526 (I232488,I232437,I1266901);
not I_13527 (I232505,I1266913);
nand I_13528 (I232522,I232505,I1266901);
not I_13529 (I232539,I1266898);
nor I_13530 (I232556,I232539,I1266910);
nand I_13531 (I232573,I232556,I1266892);
nor I_13532 (I232590,I232573,I232522);
DFFARX1 I_13533 (I232590,I2507,I232372,I232340,);
not I_13534 (I232621,I232573);
not I_13535 (I232638,I1266910);
nand I_13536 (I232655,I232638,I1266901);
nor I_13537 (I232672,I1266910,I1266913);
nand I_13538 (I232352,I232488,I232672);
nand I_13539 (I232346,I232437,I1266910);
nand I_13540 (I232717,I232539,I1266904);
DFFARX1 I_13541 (I232717,I2507,I232372,I232361,);
DFFARX1 I_13542 (I232717,I2507,I232372,I232355,);
not I_13543 (I232762,I1266904);
nor I_13544 (I232779,I232762,I1266895);
and I_13545 (I232796,I232779,I1266892);
or I_13546 (I232813,I232796,I1266916);
DFFARX1 I_13547 (I232813,I2507,I232372,I232839,);
nand I_13548 (I232847,I232839,I232505);
nor I_13549 (I232349,I232847,I232655);
nor I_13550 (I232343,I232839,I232471);
DFFARX1 I_13551 (I232839,I2507,I232372,I232901,);
not I_13552 (I232909,I232901);
nor I_13553 (I232358,I232909,I232621);
not I_13554 (I232967,I2514);
DFFARX1 I_13555 (I1383278,I2507,I232967,I232993,);
DFFARX1 I_13556 (I232993,I2507,I232967,I233010,);
not I_13557 (I232959,I233010);
not I_13558 (I233032,I232993);
DFFARX1 I_13559 (I1383269,I2507,I232967,I233058,);
not I_13560 (I233066,I233058);
and I_13561 (I233083,I233032,I1383263);
not I_13562 (I233100,I1383257);
nand I_13563 (I233117,I233100,I1383263);
not I_13564 (I233134,I1383284);
nor I_13565 (I233151,I233134,I1383257);
nand I_13566 (I233168,I233151,I1383281);
nor I_13567 (I233185,I233168,I233117);
DFFARX1 I_13568 (I233185,I2507,I232967,I232935,);
not I_13569 (I233216,I233168);
not I_13570 (I233233,I1383257);
nand I_13571 (I233250,I233233,I1383263);
nor I_13572 (I233267,I1383257,I1383257);
nand I_13573 (I232947,I233083,I233267);
nand I_13574 (I232941,I233032,I1383257);
nand I_13575 (I233312,I233134,I1383266);
DFFARX1 I_13576 (I233312,I2507,I232967,I232956,);
DFFARX1 I_13577 (I233312,I2507,I232967,I232950,);
not I_13578 (I233357,I1383266);
nor I_13579 (I233374,I233357,I1383272);
and I_13580 (I233391,I233374,I1383275);
or I_13581 (I233408,I233391,I1383260);
DFFARX1 I_13582 (I233408,I2507,I232967,I233434,);
nand I_13583 (I233442,I233434,I233100);
nor I_13584 (I232944,I233442,I233250);
nor I_13585 (I232938,I233434,I233066);
DFFARX1 I_13586 (I233434,I2507,I232967,I233496,);
not I_13587 (I233504,I233496);
nor I_13588 (I232953,I233504,I233216);
not I_13589 (I233562,I2514);
DFFARX1 I_13590 (I358752,I2507,I233562,I233588,);
DFFARX1 I_13591 (I233588,I2507,I233562,I233605,);
not I_13592 (I233554,I233605);
not I_13593 (I233627,I233588);
DFFARX1 I_13594 (I358767,I2507,I233562,I233653,);
not I_13595 (I233661,I233653);
and I_13596 (I233678,I233627,I358764);
not I_13597 (I233695,I358752);
nand I_13598 (I233712,I233695,I358764);
not I_13599 (I233729,I358761);
nor I_13600 (I233746,I233729,I358776);
nand I_13601 (I233763,I233746,I358773);
nor I_13602 (I233780,I233763,I233712);
DFFARX1 I_13603 (I233780,I2507,I233562,I233530,);
not I_13604 (I233811,I233763);
not I_13605 (I233828,I358776);
nand I_13606 (I233845,I233828,I358764);
nor I_13607 (I233862,I358776,I358752);
nand I_13608 (I233542,I233678,I233862);
nand I_13609 (I233536,I233627,I358776);
nand I_13610 (I233907,I233729,I358770);
DFFARX1 I_13611 (I233907,I2507,I233562,I233551,);
DFFARX1 I_13612 (I233907,I2507,I233562,I233545,);
not I_13613 (I233952,I358770);
nor I_13614 (I233969,I233952,I358758);
and I_13615 (I233986,I233969,I358779);
or I_13616 (I234003,I233986,I358755);
DFFARX1 I_13617 (I234003,I2507,I233562,I234029,);
nand I_13618 (I234037,I234029,I233695);
nor I_13619 (I233539,I234037,I233845);
nor I_13620 (I233533,I234029,I233661);
DFFARX1 I_13621 (I234029,I2507,I233562,I234091,);
not I_13622 (I234099,I234091);
nor I_13623 (I233548,I234099,I233811);
not I_13624 (I234157,I2514);
DFFARX1 I_13625 (I624953,I2507,I234157,I234183,);
DFFARX1 I_13626 (I234183,I2507,I234157,I234200,);
not I_13627 (I234149,I234200);
not I_13628 (I234222,I234183);
DFFARX1 I_13629 (I624944,I2507,I234157,I234248,);
not I_13630 (I234256,I234248);
and I_13631 (I234273,I234222,I624962);
not I_13632 (I234290,I624959);
nand I_13633 (I234307,I234290,I624962);
not I_13634 (I234324,I624938);
nor I_13635 (I234341,I234324,I624941);
nand I_13636 (I234358,I234341,I624950);
nor I_13637 (I234375,I234358,I234307);
DFFARX1 I_13638 (I234375,I2507,I234157,I234125,);
not I_13639 (I234406,I234358);
not I_13640 (I234423,I624941);
nand I_13641 (I234440,I234423,I624962);
nor I_13642 (I234457,I624941,I624959);
nand I_13643 (I234137,I234273,I234457);
nand I_13644 (I234131,I234222,I624941);
nand I_13645 (I234502,I234324,I624956);
DFFARX1 I_13646 (I234502,I2507,I234157,I234146,);
DFFARX1 I_13647 (I234502,I2507,I234157,I234140,);
not I_13648 (I234547,I624956);
nor I_13649 (I234564,I234547,I624938);
and I_13650 (I234581,I234564,I624947);
or I_13651 (I234598,I234581,I624941);
DFFARX1 I_13652 (I234598,I2507,I234157,I234624,);
nand I_13653 (I234632,I234624,I234290);
nor I_13654 (I234134,I234632,I234440);
nor I_13655 (I234128,I234624,I234256);
DFFARX1 I_13656 (I234624,I2507,I234157,I234686,);
not I_13657 (I234694,I234686);
nor I_13658 (I234143,I234694,I234406);
not I_13659 (I234752,I2514);
DFFARX1 I_13660 (I461575,I2507,I234752,I234778,);
DFFARX1 I_13661 (I234778,I2507,I234752,I234795,);
not I_13662 (I234744,I234795);
not I_13663 (I234817,I234778);
DFFARX1 I_13664 (I461563,I2507,I234752,I234843,);
not I_13665 (I234851,I234843);
and I_13666 (I234868,I234817,I461572);
not I_13667 (I234885,I461569);
nand I_13668 (I234902,I234885,I461572);
not I_13669 (I234919,I461560);
nor I_13670 (I234936,I234919,I461566);
nand I_13671 (I234953,I234936,I461551);
nor I_13672 (I234970,I234953,I234902);
DFFARX1 I_13673 (I234970,I2507,I234752,I234720,);
not I_13674 (I235001,I234953);
not I_13675 (I235018,I461566);
nand I_13676 (I235035,I235018,I461572);
nor I_13677 (I235052,I461566,I461569);
nand I_13678 (I234732,I234868,I235052);
nand I_13679 (I234726,I234817,I461566);
nand I_13680 (I235097,I234919,I461551);
DFFARX1 I_13681 (I235097,I2507,I234752,I234741,);
DFFARX1 I_13682 (I235097,I2507,I234752,I234735,);
not I_13683 (I235142,I461551);
nor I_13684 (I235159,I235142,I461557);
and I_13685 (I235176,I235159,I461554);
or I_13686 (I235193,I235176,I461578);
DFFARX1 I_13687 (I235193,I2507,I234752,I235219,);
nand I_13688 (I235227,I235219,I234885);
nor I_13689 (I234729,I235227,I235035);
nor I_13690 (I234723,I235219,I234851);
DFFARX1 I_13691 (I235219,I2507,I234752,I235281,);
not I_13692 (I235289,I235281);
nor I_13693 (I234738,I235289,I235001);
not I_13694 (I235347,I2514);
DFFARX1 I_13695 (I487687,I2507,I235347,I235373,);
DFFARX1 I_13696 (I235373,I2507,I235347,I235390,);
not I_13697 (I235339,I235390);
not I_13698 (I235412,I235373);
DFFARX1 I_13699 (I487675,I2507,I235347,I235438,);
not I_13700 (I235446,I235438);
and I_13701 (I235463,I235412,I487684);
not I_13702 (I235480,I487681);
nand I_13703 (I235497,I235480,I487684);
not I_13704 (I235514,I487672);
nor I_13705 (I235531,I235514,I487678);
nand I_13706 (I235548,I235531,I487663);
nor I_13707 (I235565,I235548,I235497);
DFFARX1 I_13708 (I235565,I2507,I235347,I235315,);
not I_13709 (I235596,I235548);
not I_13710 (I235613,I487678);
nand I_13711 (I235630,I235613,I487684);
nor I_13712 (I235647,I487678,I487681);
nand I_13713 (I235327,I235463,I235647);
nand I_13714 (I235321,I235412,I487678);
nand I_13715 (I235692,I235514,I487663);
DFFARX1 I_13716 (I235692,I2507,I235347,I235336,);
DFFARX1 I_13717 (I235692,I2507,I235347,I235330,);
not I_13718 (I235737,I487663);
nor I_13719 (I235754,I235737,I487669);
and I_13720 (I235771,I235754,I487666);
or I_13721 (I235788,I235771,I487690);
DFFARX1 I_13722 (I235788,I2507,I235347,I235814,);
nand I_13723 (I235822,I235814,I235480);
nor I_13724 (I235324,I235822,I235630);
nor I_13725 (I235318,I235814,I235446);
DFFARX1 I_13726 (I235814,I2507,I235347,I235876,);
not I_13727 (I235884,I235876);
nor I_13728 (I235333,I235884,I235596);
not I_13729 (I235942,I2514);
DFFARX1 I_13730 (I378343,I2507,I235942,I235968,);
DFFARX1 I_13731 (I235968,I2507,I235942,I235985,);
not I_13732 (I235934,I235985);
not I_13733 (I236007,I235968);
DFFARX1 I_13734 (I378331,I2507,I235942,I236033,);
not I_13735 (I236041,I236033);
and I_13736 (I236058,I236007,I378340);
not I_13737 (I236075,I378337);
nand I_13738 (I236092,I236075,I378340);
not I_13739 (I236109,I378328);
nor I_13740 (I236126,I236109,I378334);
nand I_13741 (I236143,I236126,I378319);
nor I_13742 (I236160,I236143,I236092);
DFFARX1 I_13743 (I236160,I2507,I235942,I235910,);
not I_13744 (I236191,I236143);
not I_13745 (I236208,I378334);
nand I_13746 (I236225,I236208,I378340);
nor I_13747 (I236242,I378334,I378337);
nand I_13748 (I235922,I236058,I236242);
nand I_13749 (I235916,I236007,I378334);
nand I_13750 (I236287,I236109,I378319);
DFFARX1 I_13751 (I236287,I2507,I235942,I235931,);
DFFARX1 I_13752 (I236287,I2507,I235942,I235925,);
not I_13753 (I236332,I378319);
nor I_13754 (I236349,I236332,I378325);
and I_13755 (I236366,I236349,I378322);
or I_13756 (I236383,I236366,I378346);
DFFARX1 I_13757 (I236383,I2507,I235942,I236409,);
nand I_13758 (I236417,I236409,I236075);
nor I_13759 (I235919,I236417,I236225);
nor I_13760 (I235913,I236409,I236041);
DFFARX1 I_13761 (I236409,I2507,I235942,I236471,);
not I_13762 (I236479,I236471);
nor I_13763 (I235928,I236479,I236191);
not I_13764 (I236537,I2514);
DFFARX1 I_13765 (I974150,I2507,I236537,I236563,);
DFFARX1 I_13766 (I236563,I2507,I236537,I236580,);
not I_13767 (I236529,I236580);
not I_13768 (I236602,I236563);
DFFARX1 I_13769 (I974159,I2507,I236537,I236628,);
not I_13770 (I236636,I236628);
and I_13771 (I236653,I236602,I974147);
not I_13772 (I236670,I974138);
nand I_13773 (I236687,I236670,I974147);
not I_13774 (I236704,I974144);
nor I_13775 (I236721,I236704,I974162);
nand I_13776 (I236738,I236721,I974135);
nor I_13777 (I236755,I236738,I236687);
DFFARX1 I_13778 (I236755,I2507,I236537,I236505,);
not I_13779 (I236786,I236738);
not I_13780 (I236803,I974162);
nand I_13781 (I236820,I236803,I974147);
nor I_13782 (I236837,I974162,I974138);
nand I_13783 (I236517,I236653,I236837);
nand I_13784 (I236511,I236602,I974162);
nand I_13785 (I236882,I236704,I974141);
DFFARX1 I_13786 (I236882,I2507,I236537,I236526,);
DFFARX1 I_13787 (I236882,I2507,I236537,I236520,);
not I_13788 (I236927,I974141);
nor I_13789 (I236944,I236927,I974153);
and I_13790 (I236961,I236944,I974135);
or I_13791 (I236978,I236961,I974156);
DFFARX1 I_13792 (I236978,I2507,I236537,I237004,);
nand I_13793 (I237012,I237004,I236670);
nor I_13794 (I236514,I237012,I236820);
nor I_13795 (I236508,I237004,I236636);
DFFARX1 I_13796 (I237004,I2507,I236537,I237066,);
not I_13797 (I237074,I237066);
nor I_13798 (I236523,I237074,I236786);
not I_13799 (I237132,I2514);
DFFARX1 I_13800 (I1074554,I2507,I237132,I237158,);
DFFARX1 I_13801 (I237158,I2507,I237132,I237175,);
not I_13802 (I237124,I237175);
not I_13803 (I237197,I237158);
DFFARX1 I_13804 (I1074554,I2507,I237132,I237223,);
not I_13805 (I237231,I237223);
and I_13806 (I237248,I237197,I1074557);
not I_13807 (I237265,I1074569);
nand I_13808 (I237282,I237265,I1074557);
not I_13809 (I237299,I1074575);
nor I_13810 (I237316,I237299,I1074566);
nand I_13811 (I237333,I237316,I1074572);
nor I_13812 (I237350,I237333,I237282);
DFFARX1 I_13813 (I237350,I2507,I237132,I237100,);
not I_13814 (I237381,I237333);
not I_13815 (I237398,I1074566);
nand I_13816 (I237415,I237398,I1074557);
nor I_13817 (I237432,I1074566,I1074569);
nand I_13818 (I237112,I237248,I237432);
nand I_13819 (I237106,I237197,I1074566);
nand I_13820 (I237477,I237299,I1074563);
DFFARX1 I_13821 (I237477,I2507,I237132,I237121,);
DFFARX1 I_13822 (I237477,I2507,I237132,I237115,);
not I_13823 (I237522,I1074563);
nor I_13824 (I237539,I237522,I1074560);
and I_13825 (I237556,I237539,I1074578);
or I_13826 (I237573,I237556,I1074557);
DFFARX1 I_13827 (I237573,I2507,I237132,I237599,);
nand I_13828 (I237607,I237599,I237265);
nor I_13829 (I237109,I237607,I237415);
nor I_13830 (I237103,I237599,I237231);
DFFARX1 I_13831 (I237599,I2507,I237132,I237661,);
not I_13832 (I237669,I237661);
nor I_13833 (I237118,I237669,I237381);
not I_13834 (I237727,I2514);
DFFARX1 I_13835 (I937974,I2507,I237727,I237753,);
DFFARX1 I_13836 (I237753,I2507,I237727,I237770,);
not I_13837 (I237719,I237770);
not I_13838 (I237792,I237753);
DFFARX1 I_13839 (I937983,I2507,I237727,I237818,);
not I_13840 (I237826,I237818);
and I_13841 (I237843,I237792,I937971);
not I_13842 (I237860,I937962);
nand I_13843 (I237877,I237860,I937971);
not I_13844 (I237894,I937968);
nor I_13845 (I237911,I237894,I937986);
nand I_13846 (I237928,I237911,I937959);
nor I_13847 (I237945,I237928,I237877);
DFFARX1 I_13848 (I237945,I2507,I237727,I237695,);
not I_13849 (I237976,I237928);
not I_13850 (I237993,I937986);
nand I_13851 (I238010,I237993,I937971);
nor I_13852 (I238027,I937986,I937962);
nand I_13853 (I237707,I237843,I238027);
nand I_13854 (I237701,I237792,I937986);
nand I_13855 (I238072,I237894,I937965);
DFFARX1 I_13856 (I238072,I2507,I237727,I237716,);
DFFARX1 I_13857 (I238072,I2507,I237727,I237710,);
not I_13858 (I238117,I937965);
nor I_13859 (I238134,I238117,I937977);
and I_13860 (I238151,I238134,I937959);
or I_13861 (I238168,I238151,I937980);
DFFARX1 I_13862 (I238168,I2507,I237727,I238194,);
nand I_13863 (I238202,I238194,I237860);
nor I_13864 (I237704,I238202,I238010);
nor I_13865 (I237698,I238194,I237826);
DFFARX1 I_13866 (I238194,I2507,I237727,I238256,);
not I_13867 (I238264,I238256);
nor I_13868 (I237713,I238264,I237976);
not I_13869 (I238322,I2514);
DFFARX1 I_13870 (I266527,I2507,I238322,I238348,);
DFFARX1 I_13871 (I238348,I2507,I238322,I238365,);
not I_13872 (I238314,I238365);
not I_13873 (I238387,I238348);
DFFARX1 I_13874 (I266542,I2507,I238322,I238413,);
not I_13875 (I238421,I238413);
and I_13876 (I238438,I238387,I266539);
not I_13877 (I238455,I266527);
nand I_13878 (I238472,I238455,I266539);
not I_13879 (I238489,I266536);
nor I_13880 (I238506,I238489,I266551);
nand I_13881 (I238523,I238506,I266548);
nor I_13882 (I238540,I238523,I238472);
DFFARX1 I_13883 (I238540,I2507,I238322,I238290,);
not I_13884 (I238571,I238523);
not I_13885 (I238588,I266551);
nand I_13886 (I238605,I238588,I266539);
nor I_13887 (I238622,I266551,I266527);
nand I_13888 (I238302,I238438,I238622);
nand I_13889 (I238296,I238387,I266551);
nand I_13890 (I238667,I238489,I266545);
DFFARX1 I_13891 (I238667,I2507,I238322,I238311,);
DFFARX1 I_13892 (I238667,I2507,I238322,I238305,);
not I_13893 (I238712,I266545);
nor I_13894 (I238729,I238712,I266533);
and I_13895 (I238746,I238729,I266554);
or I_13896 (I238763,I238746,I266530);
DFFARX1 I_13897 (I238763,I2507,I238322,I238789,);
nand I_13898 (I238797,I238789,I238455);
nor I_13899 (I238299,I238797,I238605);
nor I_13900 (I238293,I238789,I238421);
DFFARX1 I_13901 (I238789,I2507,I238322,I238851,);
not I_13902 (I238859,I238851);
nor I_13903 (I238308,I238859,I238571);
not I_13904 (I238917,I2514);
DFFARX1 I_13905 (I493671,I2507,I238917,I238943,);
DFFARX1 I_13906 (I238943,I2507,I238917,I238960,);
not I_13907 (I238909,I238960);
not I_13908 (I238982,I238943);
DFFARX1 I_13909 (I493659,I2507,I238917,I239008,);
not I_13910 (I239016,I239008);
and I_13911 (I239033,I238982,I493668);
not I_13912 (I239050,I493665);
nand I_13913 (I239067,I239050,I493668);
not I_13914 (I239084,I493656);
nor I_13915 (I239101,I239084,I493662);
nand I_13916 (I239118,I239101,I493647);
nor I_13917 (I239135,I239118,I239067);
DFFARX1 I_13918 (I239135,I2507,I238917,I238885,);
not I_13919 (I239166,I239118);
not I_13920 (I239183,I493662);
nand I_13921 (I239200,I239183,I493668);
nor I_13922 (I239217,I493662,I493665);
nand I_13923 (I238897,I239033,I239217);
nand I_13924 (I238891,I238982,I493662);
nand I_13925 (I239262,I239084,I493647);
DFFARX1 I_13926 (I239262,I2507,I238917,I238906,);
DFFARX1 I_13927 (I239262,I2507,I238917,I238900,);
not I_13928 (I239307,I493647);
nor I_13929 (I239324,I239307,I493653);
and I_13930 (I239341,I239324,I493650);
or I_13931 (I239358,I239341,I493674);
DFFARX1 I_13932 (I239358,I2507,I238917,I239384,);
nand I_13933 (I239392,I239384,I239050);
nor I_13934 (I238894,I239392,I239200);
nor I_13935 (I238888,I239384,I239016);
DFFARX1 I_13936 (I239384,I2507,I238917,I239446,);
not I_13937 (I239454,I239446);
nor I_13938 (I238903,I239454,I239166);
not I_13939 (I239512,I2514);
DFFARX1 I_13940 (I65936,I2507,I239512,I239538,);
DFFARX1 I_13941 (I239538,I2507,I239512,I239555,);
not I_13942 (I239504,I239555);
not I_13943 (I239577,I239538);
DFFARX1 I_13944 (I65930,I2507,I239512,I239603,);
not I_13945 (I239611,I239603);
and I_13946 (I239628,I239577,I65927);
not I_13947 (I239645,I65948);
nand I_13948 (I239662,I239645,I65927);
not I_13949 (I239679,I65942);
nor I_13950 (I239696,I239679,I65933);
nand I_13951 (I239713,I239696,I65939);
nor I_13952 (I239730,I239713,I239662);
DFFARX1 I_13953 (I239730,I2507,I239512,I239480,);
not I_13954 (I239761,I239713);
not I_13955 (I239778,I65933);
nand I_13956 (I239795,I239778,I65927);
nor I_13957 (I239812,I65933,I65948);
nand I_13958 (I239492,I239628,I239812);
nand I_13959 (I239486,I239577,I65933);
nand I_13960 (I239857,I239679,I65927);
DFFARX1 I_13961 (I239857,I2507,I239512,I239501,);
DFFARX1 I_13962 (I239857,I2507,I239512,I239495,);
not I_13963 (I239902,I65927);
nor I_13964 (I239919,I239902,I65945);
and I_13965 (I239936,I239919,I65951);
or I_13966 (I239953,I239936,I65930);
DFFARX1 I_13967 (I239953,I2507,I239512,I239979,);
nand I_13968 (I239987,I239979,I239645);
nor I_13969 (I239489,I239987,I239795);
nor I_13970 (I239483,I239979,I239611);
DFFARX1 I_13971 (I239979,I2507,I239512,I240041,);
not I_13972 (I240049,I240041);
nor I_13973 (I239498,I240049,I239761);
not I_13974 (I240107,I2514);
DFFARX1 I_13975 (I1290593,I2507,I240107,I240133,);
DFFARX1 I_13976 (I240133,I2507,I240107,I240150,);
not I_13977 (I240099,I240150);
not I_13978 (I240172,I240133);
DFFARX1 I_13979 (I1290605,I2507,I240107,I240198,);
not I_13980 (I240206,I240198);
and I_13981 (I240223,I240172,I1290599);
not I_13982 (I240240,I1290611);
nand I_13983 (I240257,I240240,I1290599);
not I_13984 (I240274,I1290596);
nor I_13985 (I240291,I240274,I1290608);
nand I_13986 (I240308,I240291,I1290590);
nor I_13987 (I240325,I240308,I240257);
DFFARX1 I_13988 (I240325,I2507,I240107,I240075,);
not I_13989 (I240356,I240308);
not I_13990 (I240373,I1290608);
nand I_13991 (I240390,I240373,I1290599);
nor I_13992 (I240407,I1290608,I1290611);
nand I_13993 (I240087,I240223,I240407);
nand I_13994 (I240081,I240172,I1290608);
nand I_13995 (I240452,I240274,I1290602);
DFFARX1 I_13996 (I240452,I2507,I240107,I240096,);
DFFARX1 I_13997 (I240452,I2507,I240107,I240090,);
not I_13998 (I240497,I1290602);
nor I_13999 (I240514,I240497,I1290593);
and I_14000 (I240531,I240514,I1290590);
or I_14001 (I240548,I240531,I1290614);
DFFARX1 I_14002 (I240548,I2507,I240107,I240574,);
nand I_14003 (I240582,I240574,I240240);
nor I_14004 (I240084,I240582,I240390);
nor I_14005 (I240078,I240574,I240206);
DFFARX1 I_14006 (I240574,I2507,I240107,I240636,);
not I_14007 (I240644,I240636);
nor I_14008 (I240093,I240644,I240356);
not I_14009 (I240702,I2514);
DFFARX1 I_14010 (I894692,I2507,I240702,I240728,);
DFFARX1 I_14011 (I240728,I2507,I240702,I240745,);
not I_14012 (I240694,I240745);
not I_14013 (I240767,I240728);
DFFARX1 I_14014 (I894701,I2507,I240702,I240793,);
not I_14015 (I240801,I240793);
and I_14016 (I240818,I240767,I894689);
not I_14017 (I240835,I894680);
nand I_14018 (I240852,I240835,I894689);
not I_14019 (I240869,I894686);
nor I_14020 (I240886,I240869,I894704);
nand I_14021 (I240903,I240886,I894677);
nor I_14022 (I240920,I240903,I240852);
DFFARX1 I_14023 (I240920,I2507,I240702,I240670,);
not I_14024 (I240951,I240903);
not I_14025 (I240968,I894704);
nand I_14026 (I240985,I240968,I894689);
nor I_14027 (I241002,I894704,I894680);
nand I_14028 (I240682,I240818,I241002);
nand I_14029 (I240676,I240767,I894704);
nand I_14030 (I241047,I240869,I894683);
DFFARX1 I_14031 (I241047,I2507,I240702,I240691,);
DFFARX1 I_14032 (I241047,I2507,I240702,I240685,);
not I_14033 (I241092,I894683);
nor I_14034 (I241109,I241092,I894695);
and I_14035 (I241126,I241109,I894677);
or I_14036 (I241143,I241126,I894698);
DFFARX1 I_14037 (I241143,I2507,I240702,I241169,);
nand I_14038 (I241177,I241169,I240835);
nor I_14039 (I240679,I241177,I240985);
nor I_14040 (I240673,I241169,I240801);
DFFARX1 I_14041 (I241169,I2507,I240702,I241231,);
not I_14042 (I241239,I241231);
nor I_14043 (I240688,I241239,I240951);
not I_14044 (I241297,I2514);
DFFARX1 I_14045 (I22210,I2507,I241297,I241323,);
DFFARX1 I_14046 (I241323,I2507,I241297,I241340,);
not I_14047 (I241289,I241340);
not I_14048 (I241362,I241323);
DFFARX1 I_14049 (I22186,I2507,I241297,I241388,);
not I_14050 (I241396,I241388);
and I_14051 (I241413,I241362,I22201);
not I_14052 (I241430,I22189);
nand I_14053 (I241447,I241430,I22201);
not I_14054 (I241464,I22192);
nor I_14055 (I241481,I241464,I22204);
nand I_14056 (I241498,I241481,I22195);
nor I_14057 (I241515,I241498,I241447);
DFFARX1 I_14058 (I241515,I2507,I241297,I241265,);
not I_14059 (I241546,I241498);
not I_14060 (I241563,I22204);
nand I_14061 (I241580,I241563,I22201);
nor I_14062 (I241597,I22204,I22189);
nand I_14063 (I241277,I241413,I241597);
nand I_14064 (I241271,I241362,I22204);
nand I_14065 (I241642,I241464,I22198);
DFFARX1 I_14066 (I241642,I2507,I241297,I241286,);
DFFARX1 I_14067 (I241642,I2507,I241297,I241280,);
not I_14068 (I241687,I22198);
nor I_14069 (I241704,I241687,I22189);
and I_14070 (I241721,I241704,I22186);
or I_14071 (I241738,I241721,I22207);
DFFARX1 I_14072 (I241738,I2507,I241297,I241764,);
nand I_14073 (I241772,I241764,I241430);
nor I_14074 (I241274,I241772,I241580);
nor I_14075 (I241268,I241764,I241396);
DFFARX1 I_14076 (I241764,I2507,I241297,I241826,);
not I_14077 (I241834,I241826);
nor I_14078 (I241283,I241834,I241546);
not I_14079 (I241892,I2514);
DFFARX1 I_14080 (I129703,I2507,I241892,I241918,);
DFFARX1 I_14081 (I241918,I2507,I241892,I241935,);
not I_14082 (I241884,I241935);
not I_14083 (I241957,I241918);
DFFARX1 I_14084 (I129697,I2507,I241892,I241983,);
not I_14085 (I241991,I241983);
and I_14086 (I242008,I241957,I129694);
not I_14087 (I242025,I129715);
nand I_14088 (I242042,I242025,I129694);
not I_14089 (I242059,I129709);
nor I_14090 (I242076,I242059,I129700);
nand I_14091 (I242093,I242076,I129706);
nor I_14092 (I242110,I242093,I242042);
DFFARX1 I_14093 (I242110,I2507,I241892,I241860,);
not I_14094 (I242141,I242093);
not I_14095 (I242158,I129700);
nand I_14096 (I242175,I242158,I129694);
nor I_14097 (I242192,I129700,I129715);
nand I_14098 (I241872,I242008,I242192);
nand I_14099 (I241866,I241957,I129700);
nand I_14100 (I242237,I242059,I129694);
DFFARX1 I_14101 (I242237,I2507,I241892,I241881,);
DFFARX1 I_14102 (I242237,I2507,I241892,I241875,);
not I_14103 (I242282,I129694);
nor I_14104 (I242299,I242282,I129712);
and I_14105 (I242316,I242299,I129718);
or I_14106 (I242333,I242316,I129697);
DFFARX1 I_14107 (I242333,I2507,I241892,I242359,);
nand I_14108 (I242367,I242359,I242025);
nor I_14109 (I241869,I242367,I242175);
nor I_14110 (I241863,I242359,I241991);
DFFARX1 I_14111 (I242359,I2507,I241892,I242421,);
not I_14112 (I242429,I242421);
nor I_14113 (I241878,I242429,I242141);
not I_14114 (I242487,I2514);
DFFARX1 I_14115 (I331875,I2507,I242487,I242513,);
DFFARX1 I_14116 (I242513,I2507,I242487,I242530,);
not I_14117 (I242479,I242530);
not I_14118 (I242552,I242513);
DFFARX1 I_14119 (I331890,I2507,I242487,I242578,);
not I_14120 (I242586,I242578);
and I_14121 (I242603,I242552,I331887);
not I_14122 (I242620,I331875);
nand I_14123 (I242637,I242620,I331887);
not I_14124 (I242654,I331884);
nor I_14125 (I242671,I242654,I331899);
nand I_14126 (I242688,I242671,I331896);
nor I_14127 (I242705,I242688,I242637);
DFFARX1 I_14128 (I242705,I2507,I242487,I242455,);
not I_14129 (I242736,I242688);
not I_14130 (I242753,I331899);
nand I_14131 (I242770,I242753,I331887);
nor I_14132 (I242787,I331899,I331875);
nand I_14133 (I242467,I242603,I242787);
nand I_14134 (I242461,I242552,I331899);
nand I_14135 (I242832,I242654,I331893);
DFFARX1 I_14136 (I242832,I2507,I242487,I242476,);
DFFARX1 I_14137 (I242832,I2507,I242487,I242470,);
not I_14138 (I242877,I331893);
nor I_14139 (I242894,I242877,I331881);
and I_14140 (I242911,I242894,I331902);
or I_14141 (I242928,I242911,I331878);
DFFARX1 I_14142 (I242928,I2507,I242487,I242954,);
nand I_14143 (I242962,I242954,I242620);
nor I_14144 (I242464,I242962,I242770);
nor I_14145 (I242458,I242954,I242586);
DFFARX1 I_14146 (I242954,I2507,I242487,I243016,);
not I_14147 (I243024,I243016);
nor I_14148 (I242473,I243024,I242736);
not I_14149 (I243082,I2514);
DFFARX1 I_14150 (I75949,I2507,I243082,I243108,);
DFFARX1 I_14151 (I243108,I2507,I243082,I243125,);
not I_14152 (I243074,I243125);
not I_14153 (I243147,I243108);
DFFARX1 I_14154 (I75943,I2507,I243082,I243173,);
not I_14155 (I243181,I243173);
and I_14156 (I243198,I243147,I75940);
not I_14157 (I243215,I75961);
nand I_14158 (I243232,I243215,I75940);
not I_14159 (I243249,I75955);
nor I_14160 (I243266,I243249,I75946);
nand I_14161 (I243283,I243266,I75952);
nor I_14162 (I243300,I243283,I243232);
DFFARX1 I_14163 (I243300,I2507,I243082,I243050,);
not I_14164 (I243331,I243283);
not I_14165 (I243348,I75946);
nand I_14166 (I243365,I243348,I75940);
nor I_14167 (I243382,I75946,I75961);
nand I_14168 (I243062,I243198,I243382);
nand I_14169 (I243056,I243147,I75946);
nand I_14170 (I243427,I243249,I75940);
DFFARX1 I_14171 (I243427,I2507,I243082,I243071,);
DFFARX1 I_14172 (I243427,I2507,I243082,I243065,);
not I_14173 (I243472,I75940);
nor I_14174 (I243489,I243472,I75958);
and I_14175 (I243506,I243489,I75964);
or I_14176 (I243523,I243506,I75943);
DFFARX1 I_14177 (I243523,I2507,I243082,I243549,);
nand I_14178 (I243557,I243549,I243215);
nor I_14179 (I243059,I243557,I243365);
nor I_14180 (I243053,I243549,I243181);
DFFARX1 I_14181 (I243549,I2507,I243082,I243611,);
not I_14182 (I243619,I243611);
nor I_14183 (I243068,I243619,I243331);
not I_14184 (I243677,I2514);
DFFARX1 I_14185 (I901152,I2507,I243677,I243703,);
DFFARX1 I_14186 (I243703,I2507,I243677,I243720,);
not I_14187 (I243669,I243720);
not I_14188 (I243742,I243703);
DFFARX1 I_14189 (I901161,I2507,I243677,I243768,);
not I_14190 (I243776,I243768);
and I_14191 (I243793,I243742,I901149);
not I_14192 (I243810,I901140);
nand I_14193 (I243827,I243810,I901149);
not I_14194 (I243844,I901146);
nor I_14195 (I243861,I243844,I901164);
nand I_14196 (I243878,I243861,I901137);
nor I_14197 (I243895,I243878,I243827);
DFFARX1 I_14198 (I243895,I2507,I243677,I243645,);
not I_14199 (I243926,I243878);
not I_14200 (I243943,I901164);
nand I_14201 (I243960,I243943,I901149);
nor I_14202 (I243977,I901164,I901140);
nand I_14203 (I243657,I243793,I243977);
nand I_14204 (I243651,I243742,I901164);
nand I_14205 (I244022,I243844,I901143);
DFFARX1 I_14206 (I244022,I2507,I243677,I243666,);
DFFARX1 I_14207 (I244022,I2507,I243677,I243660,);
not I_14208 (I244067,I901143);
nor I_14209 (I244084,I244067,I901155);
and I_14210 (I244101,I244084,I901137);
or I_14211 (I244118,I244101,I901158);
DFFARX1 I_14212 (I244118,I2507,I243677,I244144,);
nand I_14213 (I244152,I244144,I243810);
nor I_14214 (I243654,I244152,I243960);
nor I_14215 (I243648,I244144,I243776);
DFFARX1 I_14216 (I244144,I2507,I243677,I244206,);
not I_14217 (I244214,I244206);
nor I_14218 (I243663,I244214,I243926);
not I_14219 (I244272,I2514);
DFFARX1 I_14220 (I1351148,I2507,I244272,I244298,);
DFFARX1 I_14221 (I244298,I2507,I244272,I244315,);
not I_14222 (I244264,I244315);
not I_14223 (I244337,I244298);
DFFARX1 I_14224 (I1351139,I2507,I244272,I244363,);
not I_14225 (I244371,I244363);
and I_14226 (I244388,I244337,I1351133);
not I_14227 (I244405,I1351127);
nand I_14228 (I244422,I244405,I1351133);
not I_14229 (I244439,I1351154);
nor I_14230 (I244456,I244439,I1351127);
nand I_14231 (I244473,I244456,I1351151);
nor I_14232 (I244490,I244473,I244422);
DFFARX1 I_14233 (I244490,I2507,I244272,I244240,);
not I_14234 (I244521,I244473);
not I_14235 (I244538,I1351127);
nand I_14236 (I244555,I244538,I1351133);
nor I_14237 (I244572,I1351127,I1351127);
nand I_14238 (I244252,I244388,I244572);
nand I_14239 (I244246,I244337,I1351127);
nand I_14240 (I244617,I244439,I1351136);
DFFARX1 I_14241 (I244617,I2507,I244272,I244261,);
DFFARX1 I_14242 (I244617,I2507,I244272,I244255,);
not I_14243 (I244662,I1351136);
nor I_14244 (I244679,I244662,I1351142);
and I_14245 (I244696,I244679,I1351145);
or I_14246 (I244713,I244696,I1351130);
DFFARX1 I_14247 (I244713,I2507,I244272,I244739,);
nand I_14248 (I244747,I244739,I244405);
nor I_14249 (I244249,I244747,I244555);
nor I_14250 (I244243,I244739,I244371);
DFFARX1 I_14251 (I244739,I2507,I244272,I244801,);
not I_14252 (I244809,I244801);
nor I_14253 (I244258,I244809,I244521);
not I_14254 (I244867,I2514);
DFFARX1 I_14255 (I482247,I2507,I244867,I244893,);
DFFARX1 I_14256 (I244893,I2507,I244867,I244910,);
not I_14257 (I244859,I244910);
not I_14258 (I244932,I244893);
DFFARX1 I_14259 (I482235,I2507,I244867,I244958,);
not I_14260 (I244966,I244958);
and I_14261 (I244983,I244932,I482244);
not I_14262 (I245000,I482241);
nand I_14263 (I245017,I245000,I482244);
not I_14264 (I245034,I482232);
nor I_14265 (I245051,I245034,I482238);
nand I_14266 (I245068,I245051,I482223);
nor I_14267 (I245085,I245068,I245017);
DFFARX1 I_14268 (I245085,I2507,I244867,I244835,);
not I_14269 (I245116,I245068);
not I_14270 (I245133,I482238);
nand I_14271 (I245150,I245133,I482244);
nor I_14272 (I245167,I482238,I482241);
nand I_14273 (I244847,I244983,I245167);
nand I_14274 (I244841,I244932,I482238);
nand I_14275 (I245212,I245034,I482223);
DFFARX1 I_14276 (I245212,I2507,I244867,I244856,);
DFFARX1 I_14277 (I245212,I2507,I244867,I244850,);
not I_14278 (I245257,I482223);
nor I_14279 (I245274,I245257,I482229);
and I_14280 (I245291,I245274,I482226);
or I_14281 (I245308,I245291,I482250);
DFFARX1 I_14282 (I245308,I2507,I244867,I245334,);
nand I_14283 (I245342,I245334,I245000);
nor I_14284 (I244844,I245342,I245150);
nor I_14285 (I244838,I245334,I244966);
DFFARX1 I_14286 (I245334,I2507,I244867,I245396,);
not I_14287 (I245404,I245396);
nor I_14288 (I244853,I245404,I245116);
not I_14289 (I245462,I2514);
DFFARX1 I_14290 (I419143,I2507,I245462,I245488,);
DFFARX1 I_14291 (I245488,I2507,I245462,I245505,);
not I_14292 (I245454,I245505);
not I_14293 (I245527,I245488);
DFFARX1 I_14294 (I419131,I2507,I245462,I245553,);
not I_14295 (I245561,I245553);
and I_14296 (I245578,I245527,I419140);
not I_14297 (I245595,I419137);
nand I_14298 (I245612,I245595,I419140);
not I_14299 (I245629,I419128);
nor I_14300 (I245646,I245629,I419134);
nand I_14301 (I245663,I245646,I419119);
nor I_14302 (I245680,I245663,I245612);
DFFARX1 I_14303 (I245680,I2507,I245462,I245430,);
not I_14304 (I245711,I245663);
not I_14305 (I245728,I419134);
nand I_14306 (I245745,I245728,I419140);
nor I_14307 (I245762,I419134,I419137);
nand I_14308 (I245442,I245578,I245762);
nand I_14309 (I245436,I245527,I419134);
nand I_14310 (I245807,I245629,I419119);
DFFARX1 I_14311 (I245807,I2507,I245462,I245451,);
DFFARX1 I_14312 (I245807,I2507,I245462,I245445,);
not I_14313 (I245852,I419119);
nor I_14314 (I245869,I245852,I419125);
and I_14315 (I245886,I245869,I419122);
or I_14316 (I245903,I245886,I419146);
DFFARX1 I_14317 (I245903,I2507,I245462,I245929,);
nand I_14318 (I245937,I245929,I245595);
nor I_14319 (I245439,I245937,I245745);
nor I_14320 (I245433,I245929,I245561);
DFFARX1 I_14321 (I245929,I2507,I245462,I245991,);
not I_14322 (I245999,I245991);
nor I_14323 (I245448,I245999,I245711);
not I_14324 (I246057,I2514);
DFFARX1 I_14325 (I35912,I2507,I246057,I246083,);
DFFARX1 I_14326 (I246083,I2507,I246057,I246100,);
not I_14327 (I246049,I246100);
not I_14328 (I246122,I246083);
DFFARX1 I_14329 (I35888,I2507,I246057,I246148,);
not I_14330 (I246156,I246148);
and I_14331 (I246173,I246122,I35903);
not I_14332 (I246190,I35891);
nand I_14333 (I246207,I246190,I35903);
not I_14334 (I246224,I35894);
nor I_14335 (I246241,I246224,I35906);
nand I_14336 (I246258,I246241,I35897);
nor I_14337 (I246275,I246258,I246207);
DFFARX1 I_14338 (I246275,I2507,I246057,I246025,);
not I_14339 (I246306,I246258);
not I_14340 (I246323,I35906);
nand I_14341 (I246340,I246323,I35903);
nor I_14342 (I246357,I35906,I35891);
nand I_14343 (I246037,I246173,I246357);
nand I_14344 (I246031,I246122,I35906);
nand I_14345 (I246402,I246224,I35900);
DFFARX1 I_14346 (I246402,I2507,I246057,I246046,);
DFFARX1 I_14347 (I246402,I2507,I246057,I246040,);
not I_14348 (I246447,I35900);
nor I_14349 (I246464,I246447,I35891);
and I_14350 (I246481,I246464,I35888);
or I_14351 (I246498,I246481,I35909);
DFFARX1 I_14352 (I246498,I2507,I246057,I246524,);
nand I_14353 (I246532,I246524,I246190);
nor I_14354 (I246034,I246532,I246340);
nor I_14355 (I246028,I246524,I246156);
DFFARX1 I_14356 (I246524,I2507,I246057,I246586,);
not I_14357 (I246594,I246586);
nor I_14358 (I246043,I246594,I246306);
not I_14359 (I246652,I2514);
DFFARX1 I_14360 (I303944,I2507,I246652,I246678,);
DFFARX1 I_14361 (I246678,I2507,I246652,I246695,);
not I_14362 (I246644,I246695);
not I_14363 (I246717,I246678);
DFFARX1 I_14364 (I303959,I2507,I246652,I246743,);
not I_14365 (I246751,I246743);
and I_14366 (I246768,I246717,I303956);
not I_14367 (I246785,I303944);
nand I_14368 (I246802,I246785,I303956);
not I_14369 (I246819,I303953);
nor I_14370 (I246836,I246819,I303968);
nand I_14371 (I246853,I246836,I303965);
nor I_14372 (I246870,I246853,I246802);
DFFARX1 I_14373 (I246870,I2507,I246652,I246620,);
not I_14374 (I246901,I246853);
not I_14375 (I246918,I303968);
nand I_14376 (I246935,I246918,I303956);
nor I_14377 (I246952,I303968,I303944);
nand I_14378 (I246632,I246768,I246952);
nand I_14379 (I246626,I246717,I303968);
nand I_14380 (I246997,I246819,I303962);
DFFARX1 I_14381 (I246997,I2507,I246652,I246641,);
DFFARX1 I_14382 (I246997,I2507,I246652,I246635,);
not I_14383 (I247042,I303962);
nor I_14384 (I247059,I247042,I303950);
and I_14385 (I247076,I247059,I303971);
or I_14386 (I247093,I247076,I303947);
DFFARX1 I_14387 (I247093,I2507,I246652,I247119,);
nand I_14388 (I247127,I247119,I246785);
nor I_14389 (I246629,I247127,I246935);
nor I_14390 (I246623,I247119,I246751);
DFFARX1 I_14391 (I247119,I2507,I246652,I247181,);
not I_14392 (I247189,I247181);
nor I_14393 (I246638,I247189,I246901);
not I_14394 (I247247,I2514);
DFFARX1 I_14395 (I132865,I2507,I247247,I247273,);
DFFARX1 I_14396 (I247273,I2507,I247247,I247290,);
not I_14397 (I247239,I247290);
not I_14398 (I247312,I247273);
DFFARX1 I_14399 (I132859,I2507,I247247,I247338,);
not I_14400 (I247346,I247338);
and I_14401 (I247363,I247312,I132856);
not I_14402 (I247380,I132877);
nand I_14403 (I247397,I247380,I132856);
not I_14404 (I247414,I132871);
nor I_14405 (I247431,I247414,I132862);
nand I_14406 (I247448,I247431,I132868);
nor I_14407 (I247465,I247448,I247397);
DFFARX1 I_14408 (I247465,I2507,I247247,I247215,);
not I_14409 (I247496,I247448);
not I_14410 (I247513,I132862);
nand I_14411 (I247530,I247513,I132856);
nor I_14412 (I247547,I132862,I132877);
nand I_14413 (I247227,I247363,I247547);
nand I_14414 (I247221,I247312,I132862);
nand I_14415 (I247592,I247414,I132856);
DFFARX1 I_14416 (I247592,I2507,I247247,I247236,);
DFFARX1 I_14417 (I247592,I2507,I247247,I247230,);
not I_14418 (I247637,I132856);
nor I_14419 (I247654,I247637,I132874);
and I_14420 (I247671,I247654,I132880);
or I_14421 (I247688,I247671,I132859);
DFFARX1 I_14422 (I247688,I2507,I247247,I247714,);
nand I_14423 (I247722,I247714,I247380);
nor I_14424 (I247224,I247722,I247530);
nor I_14425 (I247218,I247714,I247346);
DFFARX1 I_14426 (I247714,I2507,I247247,I247776,);
not I_14427 (I247784,I247776);
nor I_14428 (I247233,I247784,I247496);
not I_14429 (I247842,I2514);
DFFARX1 I_14430 (I264946,I2507,I247842,I247868,);
DFFARX1 I_14431 (I247868,I2507,I247842,I247885,);
not I_14432 (I247834,I247885);
not I_14433 (I247907,I247868);
DFFARX1 I_14434 (I264961,I2507,I247842,I247933,);
not I_14435 (I247941,I247933);
and I_14436 (I247958,I247907,I264958);
not I_14437 (I247975,I264946);
nand I_14438 (I247992,I247975,I264958);
not I_14439 (I248009,I264955);
nor I_14440 (I248026,I248009,I264970);
nand I_14441 (I248043,I248026,I264967);
nor I_14442 (I248060,I248043,I247992);
DFFARX1 I_14443 (I248060,I2507,I247842,I247810,);
not I_14444 (I248091,I248043);
not I_14445 (I248108,I264970);
nand I_14446 (I248125,I248108,I264958);
nor I_14447 (I248142,I264970,I264946);
nand I_14448 (I247822,I247958,I248142);
nand I_14449 (I247816,I247907,I264970);
nand I_14450 (I248187,I248009,I264964);
DFFARX1 I_14451 (I248187,I2507,I247842,I247831,);
DFFARX1 I_14452 (I248187,I2507,I247842,I247825,);
not I_14453 (I248232,I264964);
nor I_14454 (I248249,I248232,I264952);
and I_14455 (I248266,I248249,I264973);
or I_14456 (I248283,I248266,I264949);
DFFARX1 I_14457 (I248283,I2507,I247842,I248309,);
nand I_14458 (I248317,I248309,I247975);
nor I_14459 (I247819,I248317,I248125);
nor I_14460 (I247813,I248309,I247941);
DFFARX1 I_14461 (I248309,I2507,I247842,I248371,);
not I_14462 (I248379,I248371);
nor I_14463 (I247828,I248379,I248091);
not I_14464 (I248437,I2514);
DFFARX1 I_14465 (I1349958,I2507,I248437,I248463,);
DFFARX1 I_14466 (I248463,I2507,I248437,I248480,);
not I_14467 (I248429,I248480);
not I_14468 (I248502,I248463);
DFFARX1 I_14469 (I1349949,I2507,I248437,I248528,);
not I_14470 (I248536,I248528);
and I_14471 (I248553,I248502,I1349943);
not I_14472 (I248570,I1349937);
nand I_14473 (I248587,I248570,I1349943);
not I_14474 (I248604,I1349964);
nor I_14475 (I248621,I248604,I1349937);
nand I_14476 (I248638,I248621,I1349961);
nor I_14477 (I248655,I248638,I248587);
DFFARX1 I_14478 (I248655,I2507,I248437,I248405,);
not I_14479 (I248686,I248638);
not I_14480 (I248703,I1349937);
nand I_14481 (I248720,I248703,I1349943);
nor I_14482 (I248737,I1349937,I1349937);
nand I_14483 (I248417,I248553,I248737);
nand I_14484 (I248411,I248502,I1349937);
nand I_14485 (I248782,I248604,I1349946);
DFFARX1 I_14486 (I248782,I2507,I248437,I248426,);
DFFARX1 I_14487 (I248782,I2507,I248437,I248420,);
not I_14488 (I248827,I1349946);
nor I_14489 (I248844,I248827,I1349952);
and I_14490 (I248861,I248844,I1349955);
or I_14491 (I248878,I248861,I1349940);
DFFARX1 I_14492 (I248878,I2507,I248437,I248904,);
nand I_14493 (I248912,I248904,I248570);
nor I_14494 (I248414,I248912,I248720);
nor I_14495 (I248408,I248904,I248536);
DFFARX1 I_14496 (I248904,I2507,I248437,I248966,);
not I_14497 (I248974,I248966);
nor I_14498 (I248423,I248974,I248686);
not I_14499 (I249032,I2514);
DFFARX1 I_14500 (I464295,I2507,I249032,I249058,);
DFFARX1 I_14501 (I249058,I2507,I249032,I249075,);
not I_14502 (I249024,I249075);
not I_14503 (I249097,I249058);
DFFARX1 I_14504 (I464283,I2507,I249032,I249123,);
not I_14505 (I249131,I249123);
and I_14506 (I249148,I249097,I464292);
not I_14507 (I249165,I464289);
nand I_14508 (I249182,I249165,I464292);
not I_14509 (I249199,I464280);
nor I_14510 (I249216,I249199,I464286);
nand I_14511 (I249233,I249216,I464271);
nor I_14512 (I249250,I249233,I249182);
DFFARX1 I_14513 (I249250,I2507,I249032,I249000,);
not I_14514 (I249281,I249233);
not I_14515 (I249298,I464286);
nand I_14516 (I249315,I249298,I464292);
nor I_14517 (I249332,I464286,I464289);
nand I_14518 (I249012,I249148,I249332);
nand I_14519 (I249006,I249097,I464286);
nand I_14520 (I249377,I249199,I464271);
DFFARX1 I_14521 (I249377,I2507,I249032,I249021,);
DFFARX1 I_14522 (I249377,I2507,I249032,I249015,);
not I_14523 (I249422,I464271);
nor I_14524 (I249439,I249422,I464277);
and I_14525 (I249456,I249439,I464274);
or I_14526 (I249473,I249456,I464298);
DFFARX1 I_14527 (I249473,I2507,I249032,I249499,);
nand I_14528 (I249507,I249499,I249165);
nor I_14529 (I249009,I249507,I249315);
nor I_14530 (I249003,I249499,I249131);
DFFARX1 I_14531 (I249499,I2507,I249032,I249561,);
not I_14532 (I249569,I249561);
nor I_14533 (I249018,I249569,I249281);
not I_14534 (I249627,I2514);
DFFARX1 I_14535 (I1186686,I2507,I249627,I249653,);
DFFARX1 I_14536 (I249653,I2507,I249627,I249670,);
not I_14537 (I249619,I249670);
not I_14538 (I249692,I249653);
DFFARX1 I_14539 (I1186686,I2507,I249627,I249718,);
not I_14540 (I249726,I249718);
and I_14541 (I249743,I249692,I1186689);
not I_14542 (I249760,I1186701);
nand I_14543 (I249777,I249760,I1186689);
not I_14544 (I249794,I1186707);
nor I_14545 (I249811,I249794,I1186698);
nand I_14546 (I249828,I249811,I1186704);
nor I_14547 (I249845,I249828,I249777);
DFFARX1 I_14548 (I249845,I2507,I249627,I249595,);
not I_14549 (I249876,I249828);
not I_14550 (I249893,I1186698);
nand I_14551 (I249910,I249893,I1186689);
nor I_14552 (I249927,I1186698,I1186701);
nand I_14553 (I249607,I249743,I249927);
nand I_14554 (I249601,I249692,I1186698);
nand I_14555 (I249972,I249794,I1186695);
DFFARX1 I_14556 (I249972,I2507,I249627,I249616,);
DFFARX1 I_14557 (I249972,I2507,I249627,I249610,);
not I_14558 (I250017,I1186695);
nor I_14559 (I250034,I250017,I1186692);
and I_14560 (I250051,I250034,I1186710);
or I_14561 (I250068,I250051,I1186689);
DFFARX1 I_14562 (I250068,I2507,I249627,I250094,);
nand I_14563 (I250102,I250094,I249760);
nor I_14564 (I249604,I250102,I249910);
nor I_14565 (I249598,I250094,I249726);
DFFARX1 I_14566 (I250094,I2507,I249627,I250156,);
not I_14567 (I250164,I250156);
nor I_14568 (I249613,I250164,I249876);
not I_14569 (I250225,I2514);
DFFARX1 I_14570 (I1320208,I2507,I250225,I250251,);
nand I_14571 (I250259,I1320187,I1320187);
and I_14572 (I250276,I250259,I1320214);
DFFARX1 I_14573 (I250276,I2507,I250225,I250302,);
nor I_14574 (I250193,I250302,I250251);
not I_14575 (I250324,I250302);
DFFARX1 I_14576 (I1320202,I2507,I250225,I250350,);
nand I_14577 (I250358,I250350,I1320205);
not I_14578 (I250375,I250358);
DFFARX1 I_14579 (I250375,I2507,I250225,I250401,);
not I_14580 (I250217,I250401);
nor I_14581 (I250423,I250251,I250358);
nor I_14582 (I250199,I250302,I250423);
DFFARX1 I_14583 (I1320196,I2507,I250225,I250463,);
DFFARX1 I_14584 (I250463,I2507,I250225,I250480,);
not I_14585 (I250488,I250480);
not I_14586 (I250505,I250463);
nand I_14587 (I250202,I250505,I250324);
nand I_14588 (I250536,I1320193,I1320190);
and I_14589 (I250553,I250536,I1320211);
DFFARX1 I_14590 (I250553,I2507,I250225,I250579,);
nor I_14591 (I250587,I250579,I250251);
DFFARX1 I_14592 (I250587,I2507,I250225,I250190,);
DFFARX1 I_14593 (I250579,I2507,I250225,I250208,);
nor I_14594 (I250632,I1320199,I1320190);
not I_14595 (I250649,I250632);
nor I_14596 (I250211,I250488,I250649);
nand I_14597 (I250196,I250505,I250649);
nor I_14598 (I250205,I250251,I250632);
DFFARX1 I_14599 (I250632,I2507,I250225,I250214,);
not I_14600 (I250752,I2514);
DFFARX1 I_14601 (I1244980,I2507,I250752,I250778,);
nand I_14602 (I250786,I1244962,I1244986);
and I_14603 (I250803,I250786,I1244977);
DFFARX1 I_14604 (I250803,I2507,I250752,I250829,);
nor I_14605 (I250720,I250829,I250778);
not I_14606 (I250851,I250829);
DFFARX1 I_14607 (I1244983,I2507,I250752,I250877,);
nand I_14608 (I250885,I250877,I1244971);
not I_14609 (I250902,I250885);
DFFARX1 I_14610 (I250902,I2507,I250752,I250928,);
not I_14611 (I250744,I250928);
nor I_14612 (I250950,I250778,I250885);
nor I_14613 (I250726,I250829,I250950);
DFFARX1 I_14614 (I1244962,I2507,I250752,I250990,);
DFFARX1 I_14615 (I250990,I2507,I250752,I251007,);
not I_14616 (I251015,I251007);
not I_14617 (I251032,I250990);
nand I_14618 (I250729,I251032,I250851);
nand I_14619 (I251063,I1244968,I1244965);
and I_14620 (I251080,I251063,I1244974);
DFFARX1 I_14621 (I251080,I2507,I250752,I251106,);
nor I_14622 (I251114,I251106,I250778);
DFFARX1 I_14623 (I251114,I2507,I250752,I250717,);
DFFARX1 I_14624 (I251106,I2507,I250752,I250735,);
nor I_14625 (I251159,I1244965,I1244965);
not I_14626 (I251176,I251159);
nor I_14627 (I250738,I251015,I251176);
nand I_14628 (I250723,I251032,I251176);
nor I_14629 (I250732,I250778,I251159);
DFFARX1 I_14630 (I251159,I2507,I250752,I250741,);
not I_14631 (I251279,I2514);
DFFARX1 I_14632 (I805413,I2507,I251279,I251305,);
nand I_14633 (I251313,I805416,I805410);
and I_14634 (I251330,I251313,I805422);
DFFARX1 I_14635 (I251330,I2507,I251279,I251356,);
nor I_14636 (I251247,I251356,I251305);
not I_14637 (I251378,I251356);
DFFARX1 I_14638 (I805425,I2507,I251279,I251404,);
nand I_14639 (I251412,I251404,I805416);
not I_14640 (I251429,I251412);
DFFARX1 I_14641 (I251429,I2507,I251279,I251455,);
not I_14642 (I251271,I251455);
nor I_14643 (I251477,I251305,I251412);
nor I_14644 (I251253,I251356,I251477);
DFFARX1 I_14645 (I805428,I2507,I251279,I251517,);
DFFARX1 I_14646 (I251517,I2507,I251279,I251534,);
not I_14647 (I251542,I251534);
not I_14648 (I251559,I251517);
nand I_14649 (I251256,I251559,I251378);
nand I_14650 (I251590,I805410,I805419);
and I_14651 (I251607,I251590,I805413);
DFFARX1 I_14652 (I251607,I2507,I251279,I251633,);
nor I_14653 (I251641,I251633,I251305);
DFFARX1 I_14654 (I251641,I2507,I251279,I251244,);
DFFARX1 I_14655 (I251633,I2507,I251279,I251262,);
nor I_14656 (I251686,I805431,I805419);
not I_14657 (I251703,I251686);
nor I_14658 (I251265,I251542,I251703);
nand I_14659 (I251250,I251559,I251703);
nor I_14660 (I251259,I251305,I251686);
DFFARX1 I_14661 (I251686,I2507,I251279,I251268,);
not I_14662 (I251806,I2514);
DFFARX1 I_14663 (I171650,I2507,I251806,I251832,);
nand I_14664 (I251840,I171650,I171656);
and I_14665 (I251857,I251840,I171674);
DFFARX1 I_14666 (I251857,I2507,I251806,I251883,);
nor I_14667 (I251774,I251883,I251832);
not I_14668 (I251905,I251883);
DFFARX1 I_14669 (I171662,I2507,I251806,I251931,);
nand I_14670 (I251939,I251931,I171659);
not I_14671 (I251956,I251939);
DFFARX1 I_14672 (I251956,I2507,I251806,I251982,);
not I_14673 (I251798,I251982);
nor I_14674 (I252004,I251832,I251939);
nor I_14675 (I251780,I251883,I252004);
DFFARX1 I_14676 (I171668,I2507,I251806,I252044,);
DFFARX1 I_14677 (I252044,I2507,I251806,I252061,);
not I_14678 (I252069,I252061);
not I_14679 (I252086,I252044);
nand I_14680 (I251783,I252086,I251905);
nand I_14681 (I252117,I171653,I171653);
and I_14682 (I252134,I252117,I171665);
DFFARX1 I_14683 (I252134,I2507,I251806,I252160,);
nor I_14684 (I252168,I252160,I251832);
DFFARX1 I_14685 (I252168,I2507,I251806,I251771,);
DFFARX1 I_14686 (I252160,I2507,I251806,I251789,);
nor I_14687 (I252213,I171671,I171653);
not I_14688 (I252230,I252213);
nor I_14689 (I251792,I252069,I252230);
nand I_14690 (I251777,I252086,I252230);
nor I_14691 (I251786,I251832,I252213);
DFFARX1 I_14692 (I252213,I2507,I251806,I251795,);
not I_14693 (I252333,I2514);
DFFARX1 I_14694 (I851789,I2507,I252333,I252359,);
nand I_14695 (I252367,I851792,I851786);
and I_14696 (I252384,I252367,I851798);
DFFARX1 I_14697 (I252384,I2507,I252333,I252410,);
nor I_14698 (I252301,I252410,I252359);
not I_14699 (I252432,I252410);
DFFARX1 I_14700 (I851801,I2507,I252333,I252458,);
nand I_14701 (I252466,I252458,I851792);
not I_14702 (I252483,I252466);
DFFARX1 I_14703 (I252483,I2507,I252333,I252509,);
not I_14704 (I252325,I252509);
nor I_14705 (I252531,I252359,I252466);
nor I_14706 (I252307,I252410,I252531);
DFFARX1 I_14707 (I851804,I2507,I252333,I252571,);
DFFARX1 I_14708 (I252571,I2507,I252333,I252588,);
not I_14709 (I252596,I252588);
not I_14710 (I252613,I252571);
nand I_14711 (I252310,I252613,I252432);
nand I_14712 (I252644,I851786,I851795);
and I_14713 (I252661,I252644,I851789);
DFFARX1 I_14714 (I252661,I2507,I252333,I252687,);
nor I_14715 (I252695,I252687,I252359);
DFFARX1 I_14716 (I252695,I2507,I252333,I252298,);
DFFARX1 I_14717 (I252687,I2507,I252333,I252316,);
nor I_14718 (I252740,I851807,I851795);
not I_14719 (I252757,I252740);
nor I_14720 (I252319,I252596,I252757);
nand I_14721 (I252304,I252613,I252757);
nor I_14722 (I252313,I252359,I252740);
DFFARX1 I_14723 (I252740,I2507,I252333,I252322,);
not I_14724 (I252860,I2514);
DFFARX1 I_14725 (I112306,I2507,I252860,I252886,);
nand I_14726 (I252894,I112318,I112327);
and I_14727 (I252911,I252894,I112306);
DFFARX1 I_14728 (I252911,I2507,I252860,I252937,);
nor I_14729 (I252828,I252937,I252886);
not I_14730 (I252959,I252937);
DFFARX1 I_14731 (I112321,I2507,I252860,I252985,);
nand I_14732 (I252993,I252985,I112309);
not I_14733 (I253010,I252993);
DFFARX1 I_14734 (I253010,I2507,I252860,I253036,);
not I_14735 (I252852,I253036);
nor I_14736 (I253058,I252886,I252993);
nor I_14737 (I252834,I252937,I253058);
DFFARX1 I_14738 (I112312,I2507,I252860,I253098,);
DFFARX1 I_14739 (I253098,I2507,I252860,I253115,);
not I_14740 (I253123,I253115);
not I_14741 (I253140,I253098);
nand I_14742 (I252837,I253140,I252959);
nand I_14743 (I253171,I112303,I112303);
and I_14744 (I253188,I253171,I112315);
DFFARX1 I_14745 (I253188,I2507,I252860,I253214,);
nor I_14746 (I253222,I253214,I252886);
DFFARX1 I_14747 (I253222,I2507,I252860,I252825,);
DFFARX1 I_14748 (I253214,I2507,I252860,I252843,);
nor I_14749 (I253267,I112324,I112303);
not I_14750 (I253284,I253267);
nor I_14751 (I252846,I253123,I253284);
nand I_14752 (I252831,I253140,I253284);
nor I_14753 (I252840,I252886,I253267);
DFFARX1 I_14754 (I253267,I2507,I252860,I252849,);
not I_14755 (I253387,I2514);
DFFARX1 I_14756 (I584493,I2507,I253387,I253413,);
nand I_14757 (I253421,I584478,I584481);
and I_14758 (I253438,I253421,I584496);
DFFARX1 I_14759 (I253438,I2507,I253387,I253464,);
nor I_14760 (I253355,I253464,I253413);
not I_14761 (I253486,I253464);
DFFARX1 I_14762 (I584490,I2507,I253387,I253512,);
nand I_14763 (I253520,I253512,I584481);
not I_14764 (I253537,I253520);
DFFARX1 I_14765 (I253537,I2507,I253387,I253563,);
not I_14766 (I253379,I253563);
nor I_14767 (I253585,I253413,I253520);
nor I_14768 (I253361,I253464,I253585);
DFFARX1 I_14769 (I584487,I2507,I253387,I253625,);
DFFARX1 I_14770 (I253625,I2507,I253387,I253642,);
not I_14771 (I253650,I253642);
not I_14772 (I253667,I253625);
nand I_14773 (I253364,I253667,I253486);
nand I_14774 (I253698,I584502,I584478);
and I_14775 (I253715,I253698,I584499);
DFFARX1 I_14776 (I253715,I2507,I253387,I253741,);
nor I_14777 (I253749,I253741,I253413);
DFFARX1 I_14778 (I253749,I2507,I253387,I253352,);
DFFARX1 I_14779 (I253741,I2507,I253387,I253370,);
nor I_14780 (I253794,I584484,I584478);
not I_14781 (I253811,I253794);
nor I_14782 (I253373,I253650,I253811);
nand I_14783 (I253358,I253667,I253811);
nor I_14784 (I253367,I253413,I253794);
DFFARX1 I_14785 (I253794,I2507,I253387,I253376,);
not I_14786 (I253914,I2514);
DFFARX1 I_14787 (I1060682,I2507,I253914,I253940,);
nand I_14788 (I253948,I1060697,I1060682);
and I_14789 (I253965,I253948,I1060700);
DFFARX1 I_14790 (I253965,I2507,I253914,I253991,);
nor I_14791 (I253882,I253991,I253940);
not I_14792 (I254013,I253991);
DFFARX1 I_14793 (I1060706,I2507,I253914,I254039,);
nand I_14794 (I254047,I254039,I1060688);
not I_14795 (I254064,I254047);
DFFARX1 I_14796 (I254064,I2507,I253914,I254090,);
not I_14797 (I253906,I254090);
nor I_14798 (I254112,I253940,I254047);
nor I_14799 (I253888,I253991,I254112);
DFFARX1 I_14800 (I1060685,I2507,I253914,I254152,);
DFFARX1 I_14801 (I254152,I2507,I253914,I254169,);
not I_14802 (I254177,I254169);
not I_14803 (I254194,I254152);
nand I_14804 (I253891,I254194,I254013);
nand I_14805 (I254225,I1060685,I1060691);
and I_14806 (I254242,I254225,I1060703);
DFFARX1 I_14807 (I254242,I2507,I253914,I254268,);
nor I_14808 (I254276,I254268,I253940);
DFFARX1 I_14809 (I254276,I2507,I253914,I253879,);
DFFARX1 I_14810 (I254268,I2507,I253914,I253897,);
nor I_14811 (I254321,I1060694,I1060691);
not I_14812 (I254338,I254321);
nor I_14813 (I253900,I254177,I254338);
nand I_14814 (I253885,I254194,I254338);
nor I_14815 (I253894,I253940,I254321);
DFFARX1 I_14816 (I254321,I2507,I253914,I253903,);
not I_14817 (I254441,I2514);
DFFARX1 I_14818 (I1341033,I2507,I254441,I254467,);
nand I_14819 (I254475,I1341012,I1341012);
and I_14820 (I254492,I254475,I1341039);
DFFARX1 I_14821 (I254492,I2507,I254441,I254518,);
nor I_14822 (I254409,I254518,I254467);
not I_14823 (I254540,I254518);
DFFARX1 I_14824 (I1341027,I2507,I254441,I254566,);
nand I_14825 (I254574,I254566,I1341030);
not I_14826 (I254591,I254574);
DFFARX1 I_14827 (I254591,I2507,I254441,I254617,);
not I_14828 (I254433,I254617);
nor I_14829 (I254639,I254467,I254574);
nor I_14830 (I254415,I254518,I254639);
DFFARX1 I_14831 (I1341021,I2507,I254441,I254679,);
DFFARX1 I_14832 (I254679,I2507,I254441,I254696,);
not I_14833 (I254704,I254696);
not I_14834 (I254721,I254679);
nand I_14835 (I254418,I254721,I254540);
nand I_14836 (I254752,I1341018,I1341015);
and I_14837 (I254769,I254752,I1341036);
DFFARX1 I_14838 (I254769,I2507,I254441,I254795,);
nor I_14839 (I254803,I254795,I254467);
DFFARX1 I_14840 (I254803,I2507,I254441,I254406,);
DFFARX1 I_14841 (I254795,I2507,I254441,I254424,);
nor I_14842 (I254848,I1341024,I1341015);
not I_14843 (I254865,I254848);
nor I_14844 (I254427,I254704,I254865);
nand I_14845 (I254412,I254721,I254865);
nor I_14846 (I254421,I254467,I254848);
DFFARX1 I_14847 (I254848,I2507,I254441,I254430,);
not I_14848 (I254968,I2514);
DFFARX1 I_14849 (I925042,I2507,I254968,I254994,);
nand I_14850 (I255002,I925039,I925057);
and I_14851 (I255019,I255002,I925048);
DFFARX1 I_14852 (I255019,I2507,I254968,I255045,);
nor I_14853 (I254936,I255045,I254994);
not I_14854 (I255067,I255045);
DFFARX1 I_14855 (I925063,I2507,I254968,I255093,);
nand I_14856 (I255101,I255093,I925045);
not I_14857 (I255118,I255101);
DFFARX1 I_14858 (I255118,I2507,I254968,I255144,);
not I_14859 (I254960,I255144);
nor I_14860 (I255166,I254994,I255101);
nor I_14861 (I254942,I255045,I255166);
DFFARX1 I_14862 (I925051,I2507,I254968,I255206,);
DFFARX1 I_14863 (I255206,I2507,I254968,I255223,);
not I_14864 (I255231,I255223);
not I_14865 (I255248,I255206);
nand I_14866 (I254945,I255248,I255067);
nand I_14867 (I255279,I925039,I925066);
and I_14868 (I255296,I255279,I925054);
DFFARX1 I_14869 (I255296,I2507,I254968,I255322,);
nor I_14870 (I255330,I255322,I254994);
DFFARX1 I_14871 (I255330,I2507,I254968,I254933,);
DFFARX1 I_14872 (I255322,I2507,I254968,I254951,);
nor I_14873 (I255375,I925060,I925066);
not I_14874 (I255392,I255375);
nor I_14875 (I254954,I255231,I255392);
nand I_14876 (I254939,I255248,I255392);
nor I_14877 (I254948,I254994,I255375);
DFFARX1 I_14878 (I255375,I2507,I254968,I254957,);
not I_14879 (I255495,I2514);
DFFARX1 I_14880 (I1082646,I2507,I255495,I255521,);
nand I_14881 (I255529,I1082661,I1082646);
and I_14882 (I255546,I255529,I1082664);
DFFARX1 I_14883 (I255546,I2507,I255495,I255572,);
nor I_14884 (I255463,I255572,I255521);
not I_14885 (I255594,I255572);
DFFARX1 I_14886 (I1082670,I2507,I255495,I255620,);
nand I_14887 (I255628,I255620,I1082652);
not I_14888 (I255645,I255628);
DFFARX1 I_14889 (I255645,I2507,I255495,I255671,);
not I_14890 (I255487,I255671);
nor I_14891 (I255693,I255521,I255628);
nor I_14892 (I255469,I255572,I255693);
DFFARX1 I_14893 (I1082649,I2507,I255495,I255733,);
DFFARX1 I_14894 (I255733,I2507,I255495,I255750,);
not I_14895 (I255758,I255750);
not I_14896 (I255775,I255733);
nand I_14897 (I255472,I255775,I255594);
nand I_14898 (I255806,I1082649,I1082655);
and I_14899 (I255823,I255806,I1082667);
DFFARX1 I_14900 (I255823,I2507,I255495,I255849,);
nor I_14901 (I255857,I255849,I255521);
DFFARX1 I_14902 (I255857,I2507,I255495,I255460,);
DFFARX1 I_14903 (I255849,I2507,I255495,I255478,);
nor I_14904 (I255902,I1082658,I1082655);
not I_14905 (I255919,I255902);
nor I_14906 (I255481,I255758,I255919);
nand I_14907 (I255466,I255775,I255919);
nor I_14908 (I255475,I255521,I255902);
DFFARX1 I_14909 (I255902,I2507,I255495,I255484,);
not I_14910 (I256022,I2514);
DFFARX1 I_14911 (I1231380,I2507,I256022,I256048,);
nand I_14912 (I256056,I1231362,I1231386);
and I_14913 (I256073,I256056,I1231377);
DFFARX1 I_14914 (I256073,I2507,I256022,I256099,);
nor I_14915 (I255990,I256099,I256048);
not I_14916 (I256121,I256099);
DFFARX1 I_14917 (I1231383,I2507,I256022,I256147,);
nand I_14918 (I256155,I256147,I1231371);
not I_14919 (I256172,I256155);
DFFARX1 I_14920 (I256172,I2507,I256022,I256198,);
not I_14921 (I256014,I256198);
nor I_14922 (I256220,I256048,I256155);
nor I_14923 (I255996,I256099,I256220);
DFFARX1 I_14924 (I1231362,I2507,I256022,I256260,);
DFFARX1 I_14925 (I256260,I2507,I256022,I256277,);
not I_14926 (I256285,I256277);
not I_14927 (I256302,I256260);
nand I_14928 (I255999,I256302,I256121);
nand I_14929 (I256333,I1231368,I1231365);
and I_14930 (I256350,I256333,I1231374);
DFFARX1 I_14931 (I256350,I2507,I256022,I256376,);
nor I_14932 (I256384,I256376,I256048);
DFFARX1 I_14933 (I256384,I2507,I256022,I255987,);
DFFARX1 I_14934 (I256376,I2507,I256022,I256005,);
nor I_14935 (I256429,I1231365,I1231365);
not I_14936 (I256446,I256429);
nor I_14937 (I256008,I256285,I256446);
nand I_14938 (I255993,I256302,I256446);
nor I_14939 (I256002,I256048,I256429);
DFFARX1 I_14940 (I256429,I2507,I256022,I256011,);
not I_14941 (I256549,I2514);
DFFARX1 I_14942 (I136021,I2507,I256549,I256575,);
nand I_14943 (I256583,I136033,I136042);
and I_14944 (I256600,I256583,I136021);
DFFARX1 I_14945 (I256600,I2507,I256549,I256626,);
nor I_14946 (I256517,I256626,I256575);
not I_14947 (I256648,I256626);
DFFARX1 I_14948 (I136036,I2507,I256549,I256674,);
nand I_14949 (I256682,I256674,I136024);
not I_14950 (I256699,I256682);
DFFARX1 I_14951 (I256699,I2507,I256549,I256725,);
not I_14952 (I256541,I256725);
nor I_14953 (I256747,I256575,I256682);
nor I_14954 (I256523,I256626,I256747);
DFFARX1 I_14955 (I136027,I2507,I256549,I256787,);
DFFARX1 I_14956 (I256787,I2507,I256549,I256804,);
not I_14957 (I256812,I256804);
not I_14958 (I256829,I256787);
nand I_14959 (I256526,I256829,I256648);
nand I_14960 (I256860,I136018,I136018);
and I_14961 (I256877,I256860,I136030);
DFFARX1 I_14962 (I256877,I2507,I256549,I256903,);
nor I_14963 (I256911,I256903,I256575);
DFFARX1 I_14964 (I256911,I2507,I256549,I256514,);
DFFARX1 I_14965 (I256903,I2507,I256549,I256532,);
nor I_14966 (I256956,I136039,I136018);
not I_14967 (I256973,I256956);
nor I_14968 (I256535,I256812,I256973);
nand I_14969 (I256520,I256829,I256973);
nor I_14970 (I256529,I256575,I256956);
DFFARX1 I_14971 (I256956,I2507,I256549,I256538,);
not I_14972 (I257076,I2514);
DFFARX1 I_14973 (I549813,I2507,I257076,I257102,);
nand I_14974 (I257110,I549798,I549801);
and I_14975 (I257127,I257110,I549816);
DFFARX1 I_14976 (I257127,I2507,I257076,I257153,);
nor I_14977 (I257044,I257153,I257102);
not I_14978 (I257175,I257153);
DFFARX1 I_14979 (I549810,I2507,I257076,I257201,);
nand I_14980 (I257209,I257201,I549801);
not I_14981 (I257226,I257209);
DFFARX1 I_14982 (I257226,I2507,I257076,I257252,);
not I_14983 (I257068,I257252);
nor I_14984 (I257274,I257102,I257209);
nor I_14985 (I257050,I257153,I257274);
DFFARX1 I_14986 (I549807,I2507,I257076,I257314,);
DFFARX1 I_14987 (I257314,I2507,I257076,I257331,);
not I_14988 (I257339,I257331);
not I_14989 (I257356,I257314);
nand I_14990 (I257053,I257356,I257175);
nand I_14991 (I257387,I549822,I549798);
and I_14992 (I257404,I257387,I549819);
DFFARX1 I_14993 (I257404,I2507,I257076,I257430,);
nor I_14994 (I257438,I257430,I257102);
DFFARX1 I_14995 (I257438,I2507,I257076,I257041,);
DFFARX1 I_14996 (I257430,I2507,I257076,I257059,);
nor I_14997 (I257483,I549804,I549798);
not I_14998 (I257500,I257483);
nor I_14999 (I257062,I257339,I257500);
nand I_15000 (I257047,I257356,I257500);
nor I_15001 (I257056,I257102,I257483);
DFFARX1 I_15002 (I257483,I2507,I257076,I257065,);
not I_15003 (I257603,I2514);
DFFARX1 I_15004 (I1321993,I2507,I257603,I257629,);
nand I_15005 (I257637,I1321972,I1321972);
and I_15006 (I257654,I257637,I1321999);
DFFARX1 I_15007 (I257654,I2507,I257603,I257680,);
nor I_15008 (I257571,I257680,I257629);
not I_15009 (I257702,I257680);
DFFARX1 I_15010 (I1321987,I2507,I257603,I257728,);
nand I_15011 (I257736,I257728,I1321990);
not I_15012 (I257753,I257736);
DFFARX1 I_15013 (I257753,I2507,I257603,I257779,);
not I_15014 (I257595,I257779);
nor I_15015 (I257801,I257629,I257736);
nor I_15016 (I257577,I257680,I257801);
DFFARX1 I_15017 (I1321981,I2507,I257603,I257841,);
DFFARX1 I_15018 (I257841,I2507,I257603,I257858,);
not I_15019 (I257866,I257858);
not I_15020 (I257883,I257841);
nand I_15021 (I257580,I257883,I257702);
nand I_15022 (I257914,I1321978,I1321975);
and I_15023 (I257931,I257914,I1321996);
DFFARX1 I_15024 (I257931,I2507,I257603,I257957,);
nor I_15025 (I257965,I257957,I257629);
DFFARX1 I_15026 (I257965,I2507,I257603,I257568,);
DFFARX1 I_15027 (I257957,I2507,I257603,I257586,);
nor I_15028 (I258010,I1321984,I1321975);
not I_15029 (I258027,I258010);
nor I_15030 (I257589,I257866,I258027);
nand I_15031 (I257574,I257883,I258027);
nor I_15032 (I257583,I257629,I258010);
DFFARX1 I_15033 (I258010,I2507,I257603,I257592,);
not I_15034 (I258130,I2514);
DFFARX1 I_15035 (I633042,I2507,I258130,I258156,);
nand I_15036 (I258164,I633033,I633048);
and I_15037 (I258181,I258164,I633054);
DFFARX1 I_15038 (I258181,I2507,I258130,I258207,);
nor I_15039 (I258098,I258207,I258156);
not I_15040 (I258229,I258207);
DFFARX1 I_15041 (I633039,I2507,I258130,I258255,);
nand I_15042 (I258263,I258255,I633033);
not I_15043 (I258280,I258263);
DFFARX1 I_15044 (I258280,I2507,I258130,I258306,);
not I_15045 (I258122,I258306);
nor I_15046 (I258328,I258156,I258263);
nor I_15047 (I258104,I258207,I258328);
DFFARX1 I_15048 (I633036,I2507,I258130,I258368,);
DFFARX1 I_15049 (I258368,I2507,I258130,I258385,);
not I_15050 (I258393,I258385);
not I_15051 (I258410,I258368);
nand I_15052 (I258107,I258410,I258229);
nand I_15053 (I258441,I633030,I633045);
and I_15054 (I258458,I258441,I633030);
DFFARX1 I_15055 (I258458,I2507,I258130,I258484,);
nor I_15056 (I258492,I258484,I258156);
DFFARX1 I_15057 (I258492,I2507,I258130,I258095,);
DFFARX1 I_15058 (I258484,I2507,I258130,I258113,);
nor I_15059 (I258537,I633051,I633045);
not I_15060 (I258554,I258537);
nor I_15061 (I258116,I258393,I258554);
nand I_15062 (I258101,I258410,I258554);
nor I_15063 (I258110,I258156,I258537);
DFFARX1 I_15064 (I258537,I2507,I258130,I258119,);
not I_15065 (I258657,I2514);
DFFARX1 I_15066 (I14808,I2507,I258657,I258683,);
nand I_15067 (I258691,I14832,I14811);
and I_15068 (I258708,I258691,I14808);
DFFARX1 I_15069 (I258708,I2507,I258657,I258734,);
nor I_15070 (I258625,I258734,I258683);
not I_15071 (I258756,I258734);
DFFARX1 I_15072 (I14814,I2507,I258657,I258782,);
nand I_15073 (I258790,I258782,I14823);
not I_15074 (I258807,I258790);
DFFARX1 I_15075 (I258807,I2507,I258657,I258833,);
not I_15076 (I258649,I258833);
nor I_15077 (I258855,I258683,I258790);
nor I_15078 (I258631,I258734,I258855);
DFFARX1 I_15079 (I14817,I2507,I258657,I258895,);
DFFARX1 I_15080 (I258895,I2507,I258657,I258912,);
not I_15081 (I258920,I258912);
not I_15082 (I258937,I258895);
nand I_15083 (I258634,I258937,I258756);
nand I_15084 (I258968,I14829,I14811);
and I_15085 (I258985,I258968,I14820);
DFFARX1 I_15086 (I258985,I2507,I258657,I259011,);
nor I_15087 (I259019,I259011,I258683);
DFFARX1 I_15088 (I259019,I2507,I258657,I258622,);
DFFARX1 I_15089 (I259011,I2507,I258657,I258640,);
nor I_15090 (I259064,I14826,I14811);
not I_15091 (I259081,I259064);
nor I_15092 (I258643,I258920,I259081);
nand I_15093 (I258628,I258937,I259081);
nor I_15094 (I258637,I258683,I259064);
DFFARX1 I_15095 (I259064,I2507,I258657,I258646,);
not I_15096 (I259184,I2514);
DFFARX1 I_15097 (I204970,I2507,I259184,I259210,);
nand I_15098 (I259218,I204970,I204976);
and I_15099 (I259235,I259218,I204994);
DFFARX1 I_15100 (I259235,I2507,I259184,I259261,);
nor I_15101 (I259152,I259261,I259210);
not I_15102 (I259283,I259261);
DFFARX1 I_15103 (I204982,I2507,I259184,I259309,);
nand I_15104 (I259317,I259309,I204979);
not I_15105 (I259334,I259317);
DFFARX1 I_15106 (I259334,I2507,I259184,I259360,);
not I_15107 (I259176,I259360);
nor I_15108 (I259382,I259210,I259317);
nor I_15109 (I259158,I259261,I259382);
DFFARX1 I_15110 (I204988,I2507,I259184,I259422,);
DFFARX1 I_15111 (I259422,I2507,I259184,I259439,);
not I_15112 (I259447,I259439);
not I_15113 (I259464,I259422);
nand I_15114 (I259161,I259464,I259283);
nand I_15115 (I259495,I204973,I204973);
and I_15116 (I259512,I259495,I204985);
DFFARX1 I_15117 (I259512,I2507,I259184,I259538,);
nor I_15118 (I259546,I259538,I259210);
DFFARX1 I_15119 (I259546,I2507,I259184,I259149,);
DFFARX1 I_15120 (I259538,I2507,I259184,I259167,);
nor I_15121 (I259591,I204991,I204973);
not I_15122 (I259608,I259591);
nor I_15123 (I259170,I259447,I259608);
nand I_15124 (I259155,I259464,I259608);
nor I_15125 (I259164,I259210,I259591);
DFFARX1 I_15126 (I259591,I2507,I259184,I259173,);
not I_15127 (I259711,I2514);
DFFARX1 I_15128 (I184145,I2507,I259711,I259737,);
nand I_15129 (I259745,I184145,I184151);
and I_15130 (I259762,I259745,I184169);
DFFARX1 I_15131 (I259762,I2507,I259711,I259788,);
nor I_15132 (I259679,I259788,I259737);
not I_15133 (I259810,I259788);
DFFARX1 I_15134 (I184157,I2507,I259711,I259836,);
nand I_15135 (I259844,I259836,I184154);
not I_15136 (I259861,I259844);
DFFARX1 I_15137 (I259861,I2507,I259711,I259887,);
not I_15138 (I259703,I259887);
nor I_15139 (I259909,I259737,I259844);
nor I_15140 (I259685,I259788,I259909);
DFFARX1 I_15141 (I184163,I2507,I259711,I259949,);
DFFARX1 I_15142 (I259949,I2507,I259711,I259966,);
not I_15143 (I259974,I259966);
not I_15144 (I259991,I259949);
nand I_15145 (I259688,I259991,I259810);
nand I_15146 (I260022,I184148,I184148);
and I_15147 (I260039,I260022,I184160);
DFFARX1 I_15148 (I260039,I2507,I259711,I260065,);
nor I_15149 (I260073,I260065,I259737);
DFFARX1 I_15150 (I260073,I2507,I259711,I259676,);
DFFARX1 I_15151 (I260065,I2507,I259711,I259694,);
nor I_15152 (I260118,I184166,I184148);
not I_15153 (I260135,I260118);
nor I_15154 (I259697,I259974,I260135);
nand I_15155 (I259682,I259991,I260135);
nor I_15156 (I259691,I259737,I260118);
DFFARX1 I_15157 (I260118,I2507,I259711,I259700,);
not I_15158 (I260238,I2514);
DFFARX1 I_15159 (I1295229,I2507,I260238,I260264,);
nand I_15160 (I260272,I1295226,I1295217);
and I_15161 (I260289,I260272,I1295214);
DFFARX1 I_15162 (I260289,I2507,I260238,I260315,);
nor I_15163 (I260206,I260315,I260264);
not I_15164 (I260337,I260315);
DFFARX1 I_15165 (I1295223,I2507,I260238,I260363,);
nand I_15166 (I260371,I260363,I1295232);
not I_15167 (I260388,I260371);
DFFARX1 I_15168 (I260388,I2507,I260238,I260414,);
not I_15169 (I260230,I260414);
nor I_15170 (I260436,I260264,I260371);
nor I_15171 (I260212,I260315,I260436);
DFFARX1 I_15172 (I1295235,I2507,I260238,I260476,);
DFFARX1 I_15173 (I260476,I2507,I260238,I260493,);
not I_15174 (I260501,I260493);
not I_15175 (I260518,I260476);
nand I_15176 (I260215,I260518,I260337);
nand I_15177 (I260549,I1295214,I1295220);
and I_15178 (I260566,I260549,I1295238);
DFFARX1 I_15179 (I260566,I2507,I260238,I260592,);
nor I_15180 (I260600,I260592,I260264);
DFFARX1 I_15181 (I260600,I2507,I260238,I260203,);
DFFARX1 I_15182 (I260592,I2507,I260238,I260221,);
nor I_15183 (I260645,I1295217,I1295220);
not I_15184 (I260662,I260645);
nor I_15185 (I260224,I260501,I260662);
nand I_15186 (I260209,I260518,I260662);
nor I_15187 (I260218,I260264,I260645);
DFFARX1 I_15188 (I260645,I2507,I260238,I260227,);
not I_15189 (I260765,I2514);
DFFARX1 I_15190 (I43266,I2507,I260765,I260791,);
nand I_15191 (I260799,I43290,I43269);
and I_15192 (I260816,I260799,I43266);
DFFARX1 I_15193 (I260816,I2507,I260765,I260842,);
nor I_15194 (I260733,I260842,I260791);
not I_15195 (I260864,I260842);
DFFARX1 I_15196 (I43272,I2507,I260765,I260890,);
nand I_15197 (I260898,I260890,I43281);
not I_15198 (I260915,I260898);
DFFARX1 I_15199 (I260915,I2507,I260765,I260941,);
not I_15200 (I260757,I260941);
nor I_15201 (I260963,I260791,I260898);
nor I_15202 (I260739,I260842,I260963);
DFFARX1 I_15203 (I43275,I2507,I260765,I261003,);
DFFARX1 I_15204 (I261003,I2507,I260765,I261020,);
not I_15205 (I261028,I261020);
not I_15206 (I261045,I261003);
nand I_15207 (I260742,I261045,I260864);
nand I_15208 (I261076,I43287,I43269);
and I_15209 (I261093,I261076,I43278);
DFFARX1 I_15210 (I261093,I2507,I260765,I261119,);
nor I_15211 (I261127,I261119,I260791);
DFFARX1 I_15212 (I261127,I2507,I260765,I260730,);
DFFARX1 I_15213 (I261119,I2507,I260765,I260748,);
nor I_15214 (I261172,I43284,I43269);
not I_15215 (I261189,I261172);
nor I_15216 (I260751,I261028,I261189);
nand I_15217 (I260736,I261045,I261189);
nor I_15218 (I260745,I260791,I261172);
DFFARX1 I_15219 (I261172,I2507,I260765,I260754,);
not I_15220 (I261292,I2514);
DFFARX1 I_15221 (I705870,I2507,I261292,I261318,);
nand I_15222 (I261326,I705861,I705876);
and I_15223 (I261343,I261326,I705882);
DFFARX1 I_15224 (I261343,I2507,I261292,I261369,);
nor I_15225 (I261260,I261369,I261318);
not I_15226 (I261391,I261369);
DFFARX1 I_15227 (I705867,I2507,I261292,I261417,);
nand I_15228 (I261425,I261417,I705861);
not I_15229 (I261442,I261425);
DFFARX1 I_15230 (I261442,I2507,I261292,I261468,);
not I_15231 (I261284,I261468);
nor I_15232 (I261490,I261318,I261425);
nor I_15233 (I261266,I261369,I261490);
DFFARX1 I_15234 (I705864,I2507,I261292,I261530,);
DFFARX1 I_15235 (I261530,I2507,I261292,I261547,);
not I_15236 (I261555,I261547);
not I_15237 (I261572,I261530);
nand I_15238 (I261269,I261572,I261391);
nand I_15239 (I261603,I705858,I705873);
and I_15240 (I261620,I261603,I705858);
DFFARX1 I_15241 (I261620,I2507,I261292,I261646,);
nor I_15242 (I261654,I261646,I261318);
DFFARX1 I_15243 (I261654,I2507,I261292,I261257,);
DFFARX1 I_15244 (I261646,I2507,I261292,I261275,);
nor I_15245 (I261699,I705879,I705873);
not I_15246 (I261716,I261699);
nor I_15247 (I261278,I261555,I261716);
nand I_15248 (I261263,I261572,I261716);
nor I_15249 (I261272,I261318,I261699);
DFFARX1 I_15250 (I261699,I2507,I261292,I261281,);
not I_15251 (I261819,I2514);
DFFARX1 I_15252 (I972200,I2507,I261819,I261845,);
nand I_15253 (I261853,I972197,I972215);
and I_15254 (I261870,I261853,I972206);
DFFARX1 I_15255 (I261870,I2507,I261819,I261896,);
nor I_15256 (I261787,I261896,I261845);
not I_15257 (I261918,I261896);
DFFARX1 I_15258 (I972221,I2507,I261819,I261944,);
nand I_15259 (I261952,I261944,I972203);
not I_15260 (I261969,I261952);
DFFARX1 I_15261 (I261969,I2507,I261819,I261995,);
not I_15262 (I261811,I261995);
nor I_15263 (I262017,I261845,I261952);
nor I_15264 (I261793,I261896,I262017);
DFFARX1 I_15265 (I972209,I2507,I261819,I262057,);
DFFARX1 I_15266 (I262057,I2507,I261819,I262074,);
not I_15267 (I262082,I262074);
not I_15268 (I262099,I262057);
nand I_15269 (I261796,I262099,I261918);
nand I_15270 (I262130,I972197,I972224);
and I_15271 (I262147,I262130,I972212);
DFFARX1 I_15272 (I262147,I2507,I261819,I262173,);
nor I_15273 (I262181,I262173,I261845);
DFFARX1 I_15274 (I262181,I2507,I261819,I261784,);
DFFARX1 I_15275 (I262173,I2507,I261819,I261802,);
nor I_15276 (I262226,I972218,I972224);
not I_15277 (I262243,I262226);
nor I_15278 (I261805,I262082,I262243);
nand I_15279 (I261790,I262099,I262243);
nor I_15280 (I261799,I261845,I262226);
DFFARX1 I_15281 (I262226,I2507,I261819,I261808,);
not I_15282 (I262346,I2514);
DFFARX1 I_15283 (I512537,I2507,I262346,I262372,);
nand I_15284 (I262380,I512537,I512549);
and I_15285 (I262397,I262380,I512534);
DFFARX1 I_15286 (I262397,I2507,I262346,I262423,);
nor I_15287 (I262314,I262423,I262372);
not I_15288 (I262445,I262423);
DFFARX1 I_15289 (I512558,I2507,I262346,I262471,);
nand I_15290 (I262479,I262471,I512555);
not I_15291 (I262496,I262479);
DFFARX1 I_15292 (I262496,I2507,I262346,I262522,);
not I_15293 (I262338,I262522);
nor I_15294 (I262544,I262372,I262479);
nor I_15295 (I262320,I262423,I262544);
DFFARX1 I_15296 (I512546,I2507,I262346,I262584,);
DFFARX1 I_15297 (I262584,I2507,I262346,I262601,);
not I_15298 (I262609,I262601);
not I_15299 (I262626,I262584);
nand I_15300 (I262323,I262626,I262445);
nand I_15301 (I262657,I512534,I512543);
and I_15302 (I262674,I262657,I512552);
DFFARX1 I_15303 (I262674,I2507,I262346,I262700,);
nor I_15304 (I262708,I262700,I262372);
DFFARX1 I_15305 (I262708,I2507,I262346,I262311,);
DFFARX1 I_15306 (I262700,I2507,I262346,I262329,);
nor I_15307 (I262753,I512540,I512543);
not I_15308 (I262770,I262753);
nor I_15309 (I262332,I262609,I262770);
nand I_15310 (I262317,I262626,I262770);
nor I_15311 (I262326,I262372,I262753);
DFFARX1 I_15312 (I262753,I2507,I262346,I262335,);
not I_15313 (I262873,I2514);
DFFARX1 I_15314 (I674658,I2507,I262873,I262899,);
nand I_15315 (I262907,I674649,I674664);
and I_15316 (I262924,I262907,I674670);
DFFARX1 I_15317 (I262924,I2507,I262873,I262950,);
nor I_15318 (I262841,I262950,I262899);
not I_15319 (I262972,I262950);
DFFARX1 I_15320 (I674655,I2507,I262873,I262998,);
nand I_15321 (I263006,I262998,I674649);
not I_15322 (I263023,I263006);
DFFARX1 I_15323 (I263023,I2507,I262873,I263049,);
not I_15324 (I262865,I263049);
nor I_15325 (I263071,I262899,I263006);
nor I_15326 (I262847,I262950,I263071);
DFFARX1 I_15327 (I674652,I2507,I262873,I263111,);
DFFARX1 I_15328 (I263111,I2507,I262873,I263128,);
not I_15329 (I263136,I263128);
not I_15330 (I263153,I263111);
nand I_15331 (I262850,I263153,I262972);
nand I_15332 (I263184,I674646,I674661);
and I_15333 (I263201,I263184,I674646);
DFFARX1 I_15334 (I263201,I2507,I262873,I263227,);
nor I_15335 (I263235,I263227,I262899);
DFFARX1 I_15336 (I263235,I2507,I262873,I262838,);
DFFARX1 I_15337 (I263227,I2507,I262873,I262856,);
nor I_15338 (I263280,I674667,I674661);
not I_15339 (I263297,I263280);
nor I_15340 (I262859,I263136,I263297);
nand I_15341 (I262844,I263153,I263297);
nor I_15342 (I262853,I262899,I263280);
DFFARX1 I_15343 (I263280,I2507,I262873,I262862,);
not I_15344 (I263400,I2514);
DFFARX1 I_15345 (I965740,I2507,I263400,I263426,);
nand I_15346 (I263434,I965737,I965755);
and I_15347 (I263451,I263434,I965746);
DFFARX1 I_15348 (I263451,I2507,I263400,I263477,);
nor I_15349 (I263368,I263477,I263426);
not I_15350 (I263499,I263477);
DFFARX1 I_15351 (I965761,I2507,I263400,I263525,);
nand I_15352 (I263533,I263525,I965743);
not I_15353 (I263550,I263533);
DFFARX1 I_15354 (I263550,I2507,I263400,I263576,);
not I_15355 (I263392,I263576);
nor I_15356 (I263598,I263426,I263533);
nor I_15357 (I263374,I263477,I263598);
DFFARX1 I_15358 (I965749,I2507,I263400,I263638,);
DFFARX1 I_15359 (I263638,I2507,I263400,I263655,);
not I_15360 (I263663,I263655);
not I_15361 (I263680,I263638);
nand I_15362 (I263377,I263680,I263499);
nand I_15363 (I263711,I965737,I965764);
and I_15364 (I263728,I263711,I965752);
DFFARX1 I_15365 (I263728,I2507,I263400,I263754,);
nor I_15366 (I263762,I263754,I263426);
DFFARX1 I_15367 (I263762,I2507,I263400,I263365,);
DFFARX1 I_15368 (I263754,I2507,I263400,I263383,);
nor I_15369 (I263807,I965758,I965764);
not I_15370 (I263824,I263807);
nor I_15371 (I263386,I263663,I263824);
nand I_15372 (I263371,I263680,I263824);
nor I_15373 (I263380,I263426,I263807);
DFFARX1 I_15374 (I263807,I2507,I263400,I263389,);
not I_15375 (I263927,I2514);
DFFARX1 I_15376 (I704714,I2507,I263927,I263953,);
nand I_15377 (I263961,I704705,I704720);
and I_15378 (I263978,I263961,I704726);
DFFARX1 I_15379 (I263978,I2507,I263927,I264004,);
nor I_15380 (I263895,I264004,I263953);
not I_15381 (I264026,I264004);
DFFARX1 I_15382 (I704711,I2507,I263927,I264052,);
nand I_15383 (I264060,I264052,I704705);
not I_15384 (I264077,I264060);
DFFARX1 I_15385 (I264077,I2507,I263927,I264103,);
not I_15386 (I263919,I264103);
nor I_15387 (I264125,I263953,I264060);
nor I_15388 (I263901,I264004,I264125);
DFFARX1 I_15389 (I704708,I2507,I263927,I264165,);
DFFARX1 I_15390 (I264165,I2507,I263927,I264182,);
not I_15391 (I264190,I264182);
not I_15392 (I264207,I264165);
nand I_15393 (I263904,I264207,I264026);
nand I_15394 (I264238,I704702,I704717);
and I_15395 (I264255,I264238,I704702);
DFFARX1 I_15396 (I264255,I2507,I263927,I264281,);
nor I_15397 (I264289,I264281,I263953);
DFFARX1 I_15398 (I264289,I2507,I263927,I263892,);
DFFARX1 I_15399 (I264281,I2507,I263927,I263910,);
nor I_15400 (I264334,I704723,I704717);
not I_15401 (I264351,I264334);
nor I_15402 (I263913,I264190,I264351);
nand I_15403 (I263898,I264207,I264351);
nor I_15404 (I263907,I263953,I264334);
DFFARX1 I_15405 (I264334,I2507,I263927,I263916,);
not I_15406 (I264454,I2514);
DFFARX1 I_15407 (I912122,I2507,I264454,I264480,);
nand I_15408 (I264488,I912119,I912137);
and I_15409 (I264505,I264488,I912128);
DFFARX1 I_15410 (I264505,I2507,I264454,I264531,);
nor I_15411 (I264422,I264531,I264480);
not I_15412 (I264553,I264531);
DFFARX1 I_15413 (I912143,I2507,I264454,I264579,);
nand I_15414 (I264587,I264579,I912125);
not I_15415 (I264604,I264587);
DFFARX1 I_15416 (I264604,I2507,I264454,I264630,);
not I_15417 (I264446,I264630);
nor I_15418 (I264652,I264480,I264587);
nor I_15419 (I264428,I264531,I264652);
DFFARX1 I_15420 (I912131,I2507,I264454,I264692,);
DFFARX1 I_15421 (I264692,I2507,I264454,I264709,);
not I_15422 (I264717,I264709);
not I_15423 (I264734,I264692);
nand I_15424 (I264431,I264734,I264553);
nand I_15425 (I264765,I912119,I912146);
and I_15426 (I264782,I264765,I912134);
DFFARX1 I_15427 (I264782,I2507,I264454,I264808,);
nor I_15428 (I264816,I264808,I264480);
DFFARX1 I_15429 (I264816,I2507,I264454,I264419,);
DFFARX1 I_15430 (I264808,I2507,I264454,I264437,);
nor I_15431 (I264861,I912140,I912146);
not I_15432 (I264878,I264861);
nor I_15433 (I264440,I264717,I264878);
nand I_15434 (I264425,I264734,I264878);
nor I_15435 (I264434,I264480,I264861);
DFFARX1 I_15436 (I264861,I2507,I264454,I264443,);
not I_15437 (I264981,I2514);
DFFARX1 I_15438 (I597787,I2507,I264981,I265007,);
nand I_15439 (I265015,I597772,I597775);
and I_15440 (I265032,I265015,I597790);
DFFARX1 I_15441 (I265032,I2507,I264981,I265058,);
nor I_15442 (I264949,I265058,I265007);
not I_15443 (I265080,I265058);
DFFARX1 I_15444 (I597784,I2507,I264981,I265106,);
nand I_15445 (I265114,I265106,I597775);
not I_15446 (I265131,I265114);
DFFARX1 I_15447 (I265131,I2507,I264981,I265157,);
not I_15448 (I264973,I265157);
nor I_15449 (I265179,I265007,I265114);
nor I_15450 (I264955,I265058,I265179);
DFFARX1 I_15451 (I597781,I2507,I264981,I265219,);
DFFARX1 I_15452 (I265219,I2507,I264981,I265236,);
not I_15453 (I265244,I265236);
not I_15454 (I265261,I265219);
nand I_15455 (I264958,I265261,I265080);
nand I_15456 (I265292,I597796,I597772);
and I_15457 (I265309,I265292,I597793);
DFFARX1 I_15458 (I265309,I2507,I264981,I265335,);
nor I_15459 (I265343,I265335,I265007);
DFFARX1 I_15460 (I265343,I2507,I264981,I264946,);
DFFARX1 I_15461 (I265335,I2507,I264981,I264964,);
nor I_15462 (I265388,I597778,I597772);
not I_15463 (I265405,I265388);
nor I_15464 (I264967,I265244,I265405);
nand I_15465 (I264952,I265261,I265405);
nor I_15466 (I264961,I265007,I265388);
DFFARX1 I_15467 (I265388,I2507,I264981,I264970,);
not I_15468 (I265508,I2514);
DFFARX1 I_15469 (I925688,I2507,I265508,I265534,);
nand I_15470 (I265542,I925685,I925703);
and I_15471 (I265559,I265542,I925694);
DFFARX1 I_15472 (I265559,I2507,I265508,I265585,);
nor I_15473 (I265476,I265585,I265534);
not I_15474 (I265607,I265585);
DFFARX1 I_15475 (I925709,I2507,I265508,I265633,);
nand I_15476 (I265641,I265633,I925691);
not I_15477 (I265658,I265641);
DFFARX1 I_15478 (I265658,I2507,I265508,I265684,);
not I_15479 (I265500,I265684);
nor I_15480 (I265706,I265534,I265641);
nor I_15481 (I265482,I265585,I265706);
DFFARX1 I_15482 (I925697,I2507,I265508,I265746,);
DFFARX1 I_15483 (I265746,I2507,I265508,I265763,);
not I_15484 (I265771,I265763);
not I_15485 (I265788,I265746);
nand I_15486 (I265485,I265788,I265607);
nand I_15487 (I265819,I925685,I925712);
and I_15488 (I265836,I265819,I925700);
DFFARX1 I_15489 (I265836,I2507,I265508,I265862,);
nor I_15490 (I265870,I265862,I265534);
DFFARX1 I_15491 (I265870,I2507,I265508,I265473,);
DFFARX1 I_15492 (I265862,I2507,I265508,I265491,);
nor I_15493 (I265915,I925706,I925712);
not I_15494 (I265932,I265915);
nor I_15495 (I265494,I265771,I265932);
nand I_15496 (I265479,I265788,I265932);
nor I_15497 (I265488,I265534,I265915);
DFFARX1 I_15498 (I265915,I2507,I265508,I265497,);
not I_15499 (I266035,I2514);
DFFARX1 I_15500 (I1063572,I2507,I266035,I266061,);
nand I_15501 (I266069,I1063587,I1063572);
and I_15502 (I266086,I266069,I1063590);
DFFARX1 I_15503 (I266086,I2507,I266035,I266112,);
nor I_15504 (I266003,I266112,I266061);
not I_15505 (I266134,I266112);
DFFARX1 I_15506 (I1063596,I2507,I266035,I266160,);
nand I_15507 (I266168,I266160,I1063578);
not I_15508 (I266185,I266168);
DFFARX1 I_15509 (I266185,I2507,I266035,I266211,);
not I_15510 (I266027,I266211);
nor I_15511 (I266233,I266061,I266168);
nor I_15512 (I266009,I266112,I266233);
DFFARX1 I_15513 (I1063575,I2507,I266035,I266273,);
DFFARX1 I_15514 (I266273,I2507,I266035,I266290,);
not I_15515 (I266298,I266290);
not I_15516 (I266315,I266273);
nand I_15517 (I266012,I266315,I266134);
nand I_15518 (I266346,I1063575,I1063581);
and I_15519 (I266363,I266346,I1063593);
DFFARX1 I_15520 (I266363,I2507,I266035,I266389,);
nor I_15521 (I266397,I266389,I266061);
DFFARX1 I_15522 (I266397,I2507,I266035,I266000,);
DFFARX1 I_15523 (I266389,I2507,I266035,I266018,);
nor I_15524 (I266442,I1063584,I1063581);
not I_15525 (I266459,I266442);
nor I_15526 (I266021,I266298,I266459);
nand I_15527 (I266006,I266315,I266459);
nor I_15528 (I266015,I266061,I266442);
DFFARX1 I_15529 (I266442,I2507,I266035,I266024,);
not I_15530 (I266562,I2514);
DFFARX1 I_15531 (I441435,I2507,I266562,I266588,);
nand I_15532 (I266596,I441447,I441426);
and I_15533 (I266613,I266596,I441450);
DFFARX1 I_15534 (I266613,I2507,I266562,I266639,);
nor I_15535 (I266530,I266639,I266588);
not I_15536 (I266661,I266639);
DFFARX1 I_15537 (I441441,I2507,I266562,I266687,);
nand I_15538 (I266695,I266687,I441423);
not I_15539 (I266712,I266695);
DFFARX1 I_15540 (I266712,I2507,I266562,I266738,);
not I_15541 (I266554,I266738);
nor I_15542 (I266760,I266588,I266695);
nor I_15543 (I266536,I266639,I266760);
DFFARX1 I_15544 (I441438,I2507,I266562,I266800,);
DFFARX1 I_15545 (I266800,I2507,I266562,I266817,);
not I_15546 (I266825,I266817);
not I_15547 (I266842,I266800);
nand I_15548 (I266539,I266842,I266661);
nand I_15549 (I266873,I441423,I441429);
and I_15550 (I266890,I266873,I441432);
DFFARX1 I_15551 (I266890,I2507,I266562,I266916,);
nor I_15552 (I266924,I266916,I266588);
DFFARX1 I_15553 (I266924,I2507,I266562,I266527,);
DFFARX1 I_15554 (I266916,I2507,I266562,I266545,);
nor I_15555 (I266969,I441444,I441429);
not I_15556 (I266986,I266969);
nor I_15557 (I266548,I266825,I266986);
nand I_15558 (I266533,I266842,I266986);
nor I_15559 (I266542,I266588,I266969);
DFFARX1 I_15560 (I266969,I2507,I266562,I266551,);
not I_15561 (I267089,I2514);
DFFARX1 I_15562 (I227580,I2507,I267089,I267115,);
nand I_15563 (I267123,I227580,I227586);
and I_15564 (I267140,I267123,I227604);
DFFARX1 I_15565 (I267140,I2507,I267089,I267166,);
nor I_15566 (I267057,I267166,I267115);
not I_15567 (I267188,I267166);
DFFARX1 I_15568 (I227592,I2507,I267089,I267214,);
nand I_15569 (I267222,I267214,I227589);
not I_15570 (I267239,I267222);
DFFARX1 I_15571 (I267239,I2507,I267089,I267265,);
not I_15572 (I267081,I267265);
nor I_15573 (I267287,I267115,I267222);
nor I_15574 (I267063,I267166,I267287);
DFFARX1 I_15575 (I227598,I2507,I267089,I267327,);
DFFARX1 I_15576 (I267327,I2507,I267089,I267344,);
not I_15577 (I267352,I267344);
not I_15578 (I267369,I267327);
nand I_15579 (I267066,I267369,I267188);
nand I_15580 (I267400,I227583,I227583);
and I_15581 (I267417,I267400,I227595);
DFFARX1 I_15582 (I267417,I2507,I267089,I267443,);
nor I_15583 (I267451,I267443,I267115);
DFFARX1 I_15584 (I267451,I2507,I267089,I267054,);
DFFARX1 I_15585 (I267443,I2507,I267089,I267072,);
nor I_15586 (I267496,I227601,I227583);
not I_15587 (I267513,I267496);
nor I_15588 (I267075,I267352,I267513);
nand I_15589 (I267060,I267369,I267513);
nor I_15590 (I267069,I267115,I267496);
DFFARX1 I_15591 (I267496,I2507,I267089,I267078,);
not I_15592 (I267616,I2514);
DFFARX1 I_15593 (I1011827,I2507,I267616,I267642,);
nand I_15594 (I267650,I1011824,I1011827);
and I_15595 (I267667,I267650,I1011836);
DFFARX1 I_15596 (I267667,I2507,I267616,I267693,);
nor I_15597 (I267584,I267693,I267642);
not I_15598 (I267715,I267693);
DFFARX1 I_15599 (I1011824,I2507,I267616,I267741,);
nand I_15600 (I267749,I267741,I1011842);
not I_15601 (I267766,I267749);
DFFARX1 I_15602 (I267766,I2507,I267616,I267792,);
not I_15603 (I267608,I267792);
nor I_15604 (I267814,I267642,I267749);
nor I_15605 (I267590,I267693,I267814);
DFFARX1 I_15606 (I1011830,I2507,I267616,I267854,);
DFFARX1 I_15607 (I267854,I2507,I267616,I267871,);
not I_15608 (I267879,I267871);
not I_15609 (I267896,I267854);
nand I_15610 (I267593,I267896,I267715);
nand I_15611 (I267927,I1011839,I1011845);
and I_15612 (I267944,I267927,I1011830);
DFFARX1 I_15613 (I267944,I2507,I267616,I267970,);
nor I_15614 (I267978,I267970,I267642);
DFFARX1 I_15615 (I267978,I2507,I267616,I267581,);
DFFARX1 I_15616 (I267970,I2507,I267616,I267599,);
nor I_15617 (I268023,I1011833,I1011845);
not I_15618 (I268040,I268023);
nor I_15619 (I267602,I267879,I268040);
nand I_15620 (I267587,I267896,I268040);
nor I_15621 (I267596,I267642,I268023);
DFFARX1 I_15622 (I268023,I2507,I267616,I267605,);
not I_15623 (I268143,I2514);
DFFARX1 I_15624 (I1119060,I2507,I268143,I268169,);
nand I_15625 (I268177,I1119075,I1119060);
and I_15626 (I268194,I268177,I1119078);
DFFARX1 I_15627 (I268194,I2507,I268143,I268220,);
nor I_15628 (I268111,I268220,I268169);
not I_15629 (I268242,I268220);
DFFARX1 I_15630 (I1119084,I2507,I268143,I268268,);
nand I_15631 (I268276,I268268,I1119066);
not I_15632 (I268293,I268276);
DFFARX1 I_15633 (I268293,I2507,I268143,I268319,);
not I_15634 (I268135,I268319);
nor I_15635 (I268341,I268169,I268276);
nor I_15636 (I268117,I268220,I268341);
DFFARX1 I_15637 (I1119063,I2507,I268143,I268381,);
DFFARX1 I_15638 (I268381,I2507,I268143,I268398,);
not I_15639 (I268406,I268398);
not I_15640 (I268423,I268381);
nand I_15641 (I268120,I268423,I268242);
nand I_15642 (I268454,I1119063,I1119069);
and I_15643 (I268471,I268454,I1119081);
DFFARX1 I_15644 (I268471,I2507,I268143,I268497,);
nor I_15645 (I268505,I268497,I268169);
DFFARX1 I_15646 (I268505,I2507,I268143,I268108,);
DFFARX1 I_15647 (I268497,I2507,I268143,I268126,);
nor I_15648 (I268550,I1119072,I1119069);
not I_15649 (I268567,I268550);
nor I_15650 (I268129,I268406,I268567);
nand I_15651 (I268114,I268423,I268567);
nor I_15652 (I268123,I268169,I268550);
DFFARX1 I_15653 (I268550,I2507,I268143,I268132,);
not I_15654 (I268670,I2514);
DFFARX1 I_15655 (I378875,I2507,I268670,I268696,);
nand I_15656 (I268704,I378887,I378866);
and I_15657 (I268721,I268704,I378890);
DFFARX1 I_15658 (I268721,I2507,I268670,I268747,);
nor I_15659 (I268638,I268747,I268696);
not I_15660 (I268769,I268747);
DFFARX1 I_15661 (I378881,I2507,I268670,I268795,);
nand I_15662 (I268803,I268795,I378863);
not I_15663 (I268820,I268803);
DFFARX1 I_15664 (I268820,I2507,I268670,I268846,);
not I_15665 (I268662,I268846);
nor I_15666 (I268868,I268696,I268803);
nor I_15667 (I268644,I268747,I268868);
DFFARX1 I_15668 (I378878,I2507,I268670,I268908,);
DFFARX1 I_15669 (I268908,I2507,I268670,I268925,);
not I_15670 (I268933,I268925);
not I_15671 (I268950,I268908);
nand I_15672 (I268647,I268950,I268769);
nand I_15673 (I268981,I378863,I378869);
and I_15674 (I268998,I268981,I378872);
DFFARX1 I_15675 (I268998,I2507,I268670,I269024,);
nor I_15676 (I269032,I269024,I268696);
DFFARX1 I_15677 (I269032,I2507,I268670,I268635,);
DFFARX1 I_15678 (I269024,I2507,I268670,I268653,);
nor I_15679 (I269077,I378884,I378869);
not I_15680 (I269094,I269077);
nor I_15681 (I268656,I268933,I269094);
nand I_15682 (I268641,I268950,I269094);
nor I_15683 (I268650,I268696,I269077);
DFFARX1 I_15684 (I269077,I2507,I268670,I268659,);
not I_15685 (I269197,I2514);
DFFARX1 I_15686 (I499447,I2507,I269197,I269223,);
nand I_15687 (I269231,I499447,I499459);
and I_15688 (I269248,I269231,I499444);
DFFARX1 I_15689 (I269248,I2507,I269197,I269274,);
nor I_15690 (I269165,I269274,I269223);
not I_15691 (I269296,I269274);
DFFARX1 I_15692 (I499468,I2507,I269197,I269322,);
nand I_15693 (I269330,I269322,I499465);
not I_15694 (I269347,I269330);
DFFARX1 I_15695 (I269347,I2507,I269197,I269373,);
not I_15696 (I269189,I269373);
nor I_15697 (I269395,I269223,I269330);
nor I_15698 (I269171,I269274,I269395);
DFFARX1 I_15699 (I499456,I2507,I269197,I269435,);
DFFARX1 I_15700 (I269435,I2507,I269197,I269452,);
not I_15701 (I269460,I269452);
not I_15702 (I269477,I269435);
nand I_15703 (I269174,I269477,I269296);
nand I_15704 (I269508,I499444,I499453);
and I_15705 (I269525,I269508,I499462);
DFFARX1 I_15706 (I269525,I2507,I269197,I269551,);
nor I_15707 (I269559,I269551,I269223);
DFFARX1 I_15708 (I269559,I2507,I269197,I269162,);
DFFARX1 I_15709 (I269551,I2507,I269197,I269180,);
nor I_15710 (I269604,I499450,I499453);
not I_15711 (I269621,I269604);
nor I_15712 (I269183,I269460,I269621);
nand I_15713 (I269168,I269477,I269621);
nor I_15714 (I269177,I269223,I269604);
DFFARX1 I_15715 (I269604,I2507,I269197,I269186,);
not I_15716 (I269724,I2514);
DFFARX1 I_15717 (I603567,I2507,I269724,I269750,);
nand I_15718 (I269758,I603552,I603555);
and I_15719 (I269775,I269758,I603570);
DFFARX1 I_15720 (I269775,I2507,I269724,I269801,);
nor I_15721 (I269692,I269801,I269750);
not I_15722 (I269823,I269801);
DFFARX1 I_15723 (I603564,I2507,I269724,I269849,);
nand I_15724 (I269857,I269849,I603555);
not I_15725 (I269874,I269857);
DFFARX1 I_15726 (I269874,I2507,I269724,I269900,);
not I_15727 (I269716,I269900);
nor I_15728 (I269922,I269750,I269857);
nor I_15729 (I269698,I269801,I269922);
DFFARX1 I_15730 (I603561,I2507,I269724,I269962,);
DFFARX1 I_15731 (I269962,I2507,I269724,I269979,);
not I_15732 (I269987,I269979);
not I_15733 (I270004,I269962);
nand I_15734 (I269701,I270004,I269823);
nand I_15735 (I270035,I603576,I603552);
and I_15736 (I270052,I270035,I603573);
DFFARX1 I_15737 (I270052,I2507,I269724,I270078,);
nor I_15738 (I270086,I270078,I269750);
DFFARX1 I_15739 (I270086,I2507,I269724,I269689,);
DFFARX1 I_15740 (I270078,I2507,I269724,I269707,);
nor I_15741 (I270131,I603558,I603552);
not I_15742 (I270148,I270131);
nor I_15743 (I269710,I269987,I270148);
nand I_15744 (I269695,I270004,I270148);
nor I_15745 (I269704,I269750,I270131);
DFFARX1 I_15746 (I270131,I2507,I269724,I269713,);
not I_15747 (I270251,I2514);
DFFARX1 I_15748 (I761358,I2507,I270251,I270277,);
nand I_15749 (I270285,I761349,I761364);
and I_15750 (I270302,I270285,I761370);
DFFARX1 I_15751 (I270302,I2507,I270251,I270328,);
nor I_15752 (I270219,I270328,I270277);
not I_15753 (I270350,I270328);
DFFARX1 I_15754 (I761355,I2507,I270251,I270376,);
nand I_15755 (I270384,I270376,I761349);
not I_15756 (I270401,I270384);
DFFARX1 I_15757 (I270401,I2507,I270251,I270427,);
not I_15758 (I270243,I270427);
nor I_15759 (I270449,I270277,I270384);
nor I_15760 (I270225,I270328,I270449);
DFFARX1 I_15761 (I761352,I2507,I270251,I270489,);
DFFARX1 I_15762 (I270489,I2507,I270251,I270506,);
not I_15763 (I270514,I270506);
not I_15764 (I270531,I270489);
nand I_15765 (I270228,I270531,I270350);
nand I_15766 (I270562,I761346,I761361);
and I_15767 (I270579,I270562,I761346);
DFFARX1 I_15768 (I270579,I2507,I270251,I270605,);
nor I_15769 (I270613,I270605,I270277);
DFFARX1 I_15770 (I270613,I2507,I270251,I270216,);
DFFARX1 I_15771 (I270605,I2507,I270251,I270234,);
nor I_15772 (I270658,I761367,I761361);
not I_15773 (I270675,I270658);
nor I_15774 (I270237,I270514,I270675);
nand I_15775 (I270222,I270531,I270675);
nor I_15776 (I270231,I270277,I270658);
DFFARX1 I_15777 (I270658,I2507,I270251,I270240,);
not I_15778 (I270778,I2514);
DFFARX1 I_15779 (I106509,I2507,I270778,I270804,);
nand I_15780 (I270812,I106521,I106530);
and I_15781 (I270829,I270812,I106509);
DFFARX1 I_15782 (I270829,I2507,I270778,I270855,);
nor I_15783 (I270746,I270855,I270804);
not I_15784 (I270877,I270855);
DFFARX1 I_15785 (I106524,I2507,I270778,I270903,);
nand I_15786 (I270911,I270903,I106512);
not I_15787 (I270928,I270911);
DFFARX1 I_15788 (I270928,I2507,I270778,I270954,);
not I_15789 (I270770,I270954);
nor I_15790 (I270976,I270804,I270911);
nor I_15791 (I270752,I270855,I270976);
DFFARX1 I_15792 (I106515,I2507,I270778,I271016,);
DFFARX1 I_15793 (I271016,I2507,I270778,I271033,);
not I_15794 (I271041,I271033);
not I_15795 (I271058,I271016);
nand I_15796 (I270755,I271058,I270877);
nand I_15797 (I271089,I106506,I106506);
and I_15798 (I271106,I271089,I106518);
DFFARX1 I_15799 (I271106,I2507,I270778,I271132,);
nor I_15800 (I271140,I271132,I270804);
DFFARX1 I_15801 (I271140,I2507,I270778,I270743,);
DFFARX1 I_15802 (I271132,I2507,I270778,I270761,);
nor I_15803 (I271185,I106527,I106506);
not I_15804 (I271202,I271185);
nor I_15805 (I270764,I271041,I271202);
nand I_15806 (I270749,I271058,I271202);
nor I_15807 (I270758,I270804,I271185);
DFFARX1 I_15808 (I271185,I2507,I270778,I270767,);
not I_15809 (I271305,I2514);
DFFARX1 I_15810 (I915998,I2507,I271305,I271331,);
nand I_15811 (I271339,I915995,I916013);
and I_15812 (I271356,I271339,I916004);
DFFARX1 I_15813 (I271356,I2507,I271305,I271382,);
nor I_15814 (I271273,I271382,I271331);
not I_15815 (I271404,I271382);
DFFARX1 I_15816 (I916019,I2507,I271305,I271430,);
nand I_15817 (I271438,I271430,I916001);
not I_15818 (I271455,I271438);
DFFARX1 I_15819 (I271455,I2507,I271305,I271481,);
not I_15820 (I271297,I271481);
nor I_15821 (I271503,I271331,I271438);
nor I_15822 (I271279,I271382,I271503);
DFFARX1 I_15823 (I916007,I2507,I271305,I271543,);
DFFARX1 I_15824 (I271543,I2507,I271305,I271560,);
not I_15825 (I271568,I271560);
not I_15826 (I271585,I271543);
nand I_15827 (I271282,I271585,I271404);
nand I_15828 (I271616,I915995,I916022);
and I_15829 (I271633,I271616,I916010);
DFFARX1 I_15830 (I271633,I2507,I271305,I271659,);
nor I_15831 (I271667,I271659,I271331);
DFFARX1 I_15832 (I271667,I2507,I271305,I271270,);
DFFARX1 I_15833 (I271659,I2507,I271305,I271288,);
nor I_15834 (I271712,I916016,I916022);
not I_15835 (I271729,I271712);
nor I_15836 (I271291,I271568,I271729);
nand I_15837 (I271276,I271585,I271729);
nor I_15838 (I271285,I271331,I271712);
DFFARX1 I_15839 (I271712,I2507,I271305,I271294,);
not I_15840 (I271832,I2514);
DFFARX1 I_15841 (I568887,I2507,I271832,I271858,);
nand I_15842 (I271866,I568872,I568875);
and I_15843 (I271883,I271866,I568890);
DFFARX1 I_15844 (I271883,I2507,I271832,I271909,);
nor I_15845 (I271800,I271909,I271858);
not I_15846 (I271931,I271909);
DFFARX1 I_15847 (I568884,I2507,I271832,I271957,);
nand I_15848 (I271965,I271957,I568875);
not I_15849 (I271982,I271965);
DFFARX1 I_15850 (I271982,I2507,I271832,I272008,);
not I_15851 (I271824,I272008);
nor I_15852 (I272030,I271858,I271965);
nor I_15853 (I271806,I271909,I272030);
DFFARX1 I_15854 (I568881,I2507,I271832,I272070,);
DFFARX1 I_15855 (I272070,I2507,I271832,I272087,);
not I_15856 (I272095,I272087);
not I_15857 (I272112,I272070);
nand I_15858 (I271809,I272112,I271931);
nand I_15859 (I272143,I568896,I568872);
and I_15860 (I272160,I272143,I568893);
DFFARX1 I_15861 (I272160,I2507,I271832,I272186,);
nor I_15862 (I272194,I272186,I271858);
DFFARX1 I_15863 (I272194,I2507,I271832,I271797,);
DFFARX1 I_15864 (I272186,I2507,I271832,I271815,);
nor I_15865 (I272239,I568878,I568872);
not I_15866 (I272256,I272239);
nor I_15867 (I271818,I272095,I272256);
nand I_15868 (I271803,I272112,I272256);
nor I_15869 (I271812,I271858,I272239);
DFFARX1 I_15870 (I272239,I2507,I271832,I271821,);
not I_15871 (I272359,I2514);
DFFARX1 I_15872 (I906954,I2507,I272359,I272385,);
nand I_15873 (I272393,I906951,I906969);
and I_15874 (I272410,I272393,I906960);
DFFARX1 I_15875 (I272410,I2507,I272359,I272436,);
nor I_15876 (I272327,I272436,I272385);
not I_15877 (I272458,I272436);
DFFARX1 I_15878 (I906975,I2507,I272359,I272484,);
nand I_15879 (I272492,I272484,I906957);
not I_15880 (I272509,I272492);
DFFARX1 I_15881 (I272509,I2507,I272359,I272535,);
not I_15882 (I272351,I272535);
nor I_15883 (I272557,I272385,I272492);
nor I_15884 (I272333,I272436,I272557);
DFFARX1 I_15885 (I906963,I2507,I272359,I272597,);
DFFARX1 I_15886 (I272597,I2507,I272359,I272614,);
not I_15887 (I272622,I272614);
not I_15888 (I272639,I272597);
nand I_15889 (I272336,I272639,I272458);
nand I_15890 (I272670,I906951,I906978);
and I_15891 (I272687,I272670,I906966);
DFFARX1 I_15892 (I272687,I2507,I272359,I272713,);
nor I_15893 (I272721,I272713,I272385);
DFFARX1 I_15894 (I272721,I2507,I272359,I272324,);
DFFARX1 I_15895 (I272713,I2507,I272359,I272342,);
nor I_15896 (I272766,I906972,I906978);
not I_15897 (I272783,I272766);
nor I_15898 (I272345,I272622,I272783);
nand I_15899 (I272330,I272639,I272783);
nor I_15900 (I272339,I272385,I272766);
DFFARX1 I_15901 (I272766,I2507,I272359,I272348,);
not I_15902 (I272886,I2514);
DFFARX1 I_15903 (I1093050,I2507,I272886,I272912,);
nand I_15904 (I272920,I1093065,I1093050);
and I_15905 (I272937,I272920,I1093068);
DFFARX1 I_15906 (I272937,I2507,I272886,I272963,);
nor I_15907 (I272854,I272963,I272912);
not I_15908 (I272985,I272963);
DFFARX1 I_15909 (I1093074,I2507,I272886,I273011,);
nand I_15910 (I273019,I273011,I1093056);
not I_15911 (I273036,I273019);
DFFARX1 I_15912 (I273036,I2507,I272886,I273062,);
not I_15913 (I272878,I273062);
nor I_15914 (I273084,I272912,I273019);
nor I_15915 (I272860,I272963,I273084);
DFFARX1 I_15916 (I1093053,I2507,I272886,I273124,);
DFFARX1 I_15917 (I273124,I2507,I272886,I273141,);
not I_15918 (I273149,I273141);
not I_15919 (I273166,I273124);
nand I_15920 (I272863,I273166,I272985);
nand I_15921 (I273197,I1093053,I1093059);
and I_15922 (I273214,I273197,I1093071);
DFFARX1 I_15923 (I273214,I2507,I272886,I273240,);
nor I_15924 (I273248,I273240,I272912);
DFFARX1 I_15925 (I273248,I2507,I272886,I272851,);
DFFARX1 I_15926 (I273240,I2507,I272886,I272869,);
nor I_15927 (I273293,I1093062,I1093059);
not I_15928 (I273310,I273293);
nor I_15929 (I272872,I273149,I273310);
nand I_15930 (I272857,I273166,I273310);
nor I_15931 (I272866,I272912,I273293);
DFFARX1 I_15932 (I273293,I2507,I272886,I272875,);
not I_15933 (I273413,I2514);
DFFARX1 I_15934 (I33253,I2507,I273413,I273439,);
nand I_15935 (I273447,I33277,I33256);
and I_15936 (I273464,I273447,I33253);
DFFARX1 I_15937 (I273464,I2507,I273413,I273490,);
nor I_15938 (I273381,I273490,I273439);
not I_15939 (I273512,I273490);
DFFARX1 I_15940 (I33259,I2507,I273413,I273538,);
nand I_15941 (I273546,I273538,I33268);
not I_15942 (I273563,I273546);
DFFARX1 I_15943 (I273563,I2507,I273413,I273589,);
not I_15944 (I273405,I273589);
nor I_15945 (I273611,I273439,I273546);
nor I_15946 (I273387,I273490,I273611);
DFFARX1 I_15947 (I33262,I2507,I273413,I273651,);
DFFARX1 I_15948 (I273651,I2507,I273413,I273668,);
not I_15949 (I273676,I273668);
not I_15950 (I273693,I273651);
nand I_15951 (I273390,I273693,I273512);
nand I_15952 (I273724,I33274,I33256);
and I_15953 (I273741,I273724,I33265);
DFFARX1 I_15954 (I273741,I2507,I273413,I273767,);
nor I_15955 (I273775,I273767,I273439);
DFFARX1 I_15956 (I273775,I2507,I273413,I273378,);
DFFARX1 I_15957 (I273767,I2507,I273413,I273396,);
nor I_15958 (I273820,I33271,I33256);
not I_15959 (I273837,I273820);
nor I_15960 (I273399,I273676,I273837);
nand I_15961 (I273384,I273693,I273837);
nor I_15962 (I273393,I273439,I273820);
DFFARX1 I_15963 (I273820,I2507,I273413,I273402,);
not I_15964 (I273940,I2514);
DFFARX1 I_15965 (I172840,I2507,I273940,I273966,);
nand I_15966 (I273974,I172840,I172846);
and I_15967 (I273991,I273974,I172864);
DFFARX1 I_15968 (I273991,I2507,I273940,I274017,);
nor I_15969 (I273908,I274017,I273966);
not I_15970 (I274039,I274017);
DFFARX1 I_15971 (I172852,I2507,I273940,I274065,);
nand I_15972 (I274073,I274065,I172849);
not I_15973 (I274090,I274073);
DFFARX1 I_15974 (I274090,I2507,I273940,I274116,);
not I_15975 (I273932,I274116);
nor I_15976 (I274138,I273966,I274073);
nor I_15977 (I273914,I274017,I274138);
DFFARX1 I_15978 (I172858,I2507,I273940,I274178,);
DFFARX1 I_15979 (I274178,I2507,I273940,I274195,);
not I_15980 (I274203,I274195);
not I_15981 (I274220,I274178);
nand I_15982 (I273917,I274220,I274039);
nand I_15983 (I274251,I172843,I172843);
and I_15984 (I274268,I274251,I172855);
DFFARX1 I_15985 (I274268,I2507,I273940,I274294,);
nor I_15986 (I274302,I274294,I273966);
DFFARX1 I_15987 (I274302,I2507,I273940,I273905,);
DFFARX1 I_15988 (I274294,I2507,I273940,I273923,);
nor I_15989 (I274347,I172861,I172843);
not I_15990 (I274364,I274347);
nor I_15991 (I273926,I274203,I274364);
nand I_15992 (I273911,I274220,I274364);
nor I_15993 (I273920,I273966,I274347);
DFFARX1 I_15994 (I274347,I2507,I273940,I273929,);
not I_15995 (I274467,I2514);
DFFARX1 I_15996 (I542877,I2507,I274467,I274493,);
nand I_15997 (I274501,I542862,I542865);
and I_15998 (I274518,I274501,I542880);
DFFARX1 I_15999 (I274518,I2507,I274467,I274544,);
nor I_16000 (I274435,I274544,I274493);
not I_16001 (I274566,I274544);
DFFARX1 I_16002 (I542874,I2507,I274467,I274592,);
nand I_16003 (I274600,I274592,I542865);
not I_16004 (I274617,I274600);
DFFARX1 I_16005 (I274617,I2507,I274467,I274643,);
not I_16006 (I274459,I274643);
nor I_16007 (I274665,I274493,I274600);
nor I_16008 (I274441,I274544,I274665);
DFFARX1 I_16009 (I542871,I2507,I274467,I274705,);
DFFARX1 I_16010 (I274705,I2507,I274467,I274722,);
not I_16011 (I274730,I274722);
not I_16012 (I274747,I274705);
nand I_16013 (I274444,I274747,I274566);
nand I_16014 (I274778,I542886,I542862);
and I_16015 (I274795,I274778,I542883);
DFFARX1 I_16016 (I274795,I2507,I274467,I274821,);
nor I_16017 (I274829,I274821,I274493);
DFFARX1 I_16018 (I274829,I2507,I274467,I274432,);
DFFARX1 I_16019 (I274821,I2507,I274467,I274450,);
nor I_16020 (I274874,I542868,I542862);
not I_16021 (I274891,I274874);
nor I_16022 (I274453,I274730,I274891);
nand I_16023 (I274438,I274747,I274891);
nor I_16024 (I274447,I274493,I274874);
DFFARX1 I_16025 (I274874,I2507,I274467,I274456,);
not I_16026 (I274994,I2514);
DFFARX1 I_16027 (I823858,I2507,I274994,I275020,);
nand I_16028 (I275028,I823861,I823855);
and I_16029 (I275045,I275028,I823867);
DFFARX1 I_16030 (I275045,I2507,I274994,I275071,);
nor I_16031 (I274962,I275071,I275020);
not I_16032 (I275093,I275071);
DFFARX1 I_16033 (I823870,I2507,I274994,I275119,);
nand I_16034 (I275127,I275119,I823861);
not I_16035 (I275144,I275127);
DFFARX1 I_16036 (I275144,I2507,I274994,I275170,);
not I_16037 (I274986,I275170);
nor I_16038 (I275192,I275020,I275127);
nor I_16039 (I274968,I275071,I275192);
DFFARX1 I_16040 (I823873,I2507,I274994,I275232,);
DFFARX1 I_16041 (I275232,I2507,I274994,I275249,);
not I_16042 (I275257,I275249);
not I_16043 (I275274,I275232);
nand I_16044 (I274971,I275274,I275093);
nand I_16045 (I275305,I823855,I823864);
and I_16046 (I275322,I275305,I823858);
DFFARX1 I_16047 (I275322,I2507,I274994,I275348,);
nor I_16048 (I275356,I275348,I275020);
DFFARX1 I_16049 (I275356,I2507,I274994,I274959,);
DFFARX1 I_16050 (I275348,I2507,I274994,I274977,);
nor I_16051 (I275401,I823876,I823864);
not I_16052 (I275418,I275401);
nor I_16053 (I274980,I275257,I275418);
nand I_16054 (I274965,I275274,I275418);
nor I_16055 (I274974,I275020,I275401);
DFFARX1 I_16056 (I275401,I2507,I274994,I274983,);
not I_16057 (I275521,I2514);
DFFARX1 I_16058 (I594319,I2507,I275521,I275547,);
nand I_16059 (I275555,I594304,I594307);
and I_16060 (I275572,I275555,I594322);
DFFARX1 I_16061 (I275572,I2507,I275521,I275598,);
nor I_16062 (I275489,I275598,I275547);
not I_16063 (I275620,I275598);
DFFARX1 I_16064 (I594316,I2507,I275521,I275646,);
nand I_16065 (I275654,I275646,I594307);
not I_16066 (I275671,I275654);
DFFARX1 I_16067 (I275671,I2507,I275521,I275697,);
not I_16068 (I275513,I275697);
nor I_16069 (I275719,I275547,I275654);
nor I_16070 (I275495,I275598,I275719);
DFFARX1 I_16071 (I594313,I2507,I275521,I275759,);
DFFARX1 I_16072 (I275759,I2507,I275521,I275776,);
not I_16073 (I275784,I275776);
not I_16074 (I275801,I275759);
nand I_16075 (I275498,I275801,I275620);
nand I_16076 (I275832,I594328,I594304);
and I_16077 (I275849,I275832,I594325);
DFFARX1 I_16078 (I275849,I2507,I275521,I275875,);
nor I_16079 (I275883,I275875,I275547);
DFFARX1 I_16080 (I275883,I2507,I275521,I275486,);
DFFARX1 I_16081 (I275875,I2507,I275521,I275504,);
nor I_16082 (I275928,I594310,I594304);
not I_16083 (I275945,I275928);
nor I_16084 (I275507,I275784,I275945);
nand I_16085 (I275492,I275801,I275945);
nor I_16086 (I275501,I275547,I275928);
DFFARX1 I_16087 (I275928,I2507,I275521,I275510,);
not I_16088 (I276048,I2514);
DFFARX1 I_16089 (I1130042,I2507,I276048,I276074,);
nand I_16090 (I276082,I1130057,I1130042);
and I_16091 (I276099,I276082,I1130060);
DFFARX1 I_16092 (I276099,I2507,I276048,I276125,);
nor I_16093 (I276016,I276125,I276074);
not I_16094 (I276147,I276125);
DFFARX1 I_16095 (I1130066,I2507,I276048,I276173,);
nand I_16096 (I276181,I276173,I1130048);
not I_16097 (I276198,I276181);
DFFARX1 I_16098 (I276198,I2507,I276048,I276224,);
not I_16099 (I276040,I276224);
nor I_16100 (I276246,I276074,I276181);
nor I_16101 (I276022,I276125,I276246);
DFFARX1 I_16102 (I1130045,I2507,I276048,I276286,);
DFFARX1 I_16103 (I276286,I2507,I276048,I276303,);
not I_16104 (I276311,I276303);
not I_16105 (I276328,I276286);
nand I_16106 (I276025,I276328,I276147);
nand I_16107 (I276359,I1130045,I1130051);
and I_16108 (I276376,I276359,I1130063);
DFFARX1 I_16109 (I276376,I2507,I276048,I276402,);
nor I_16110 (I276410,I276402,I276074);
DFFARX1 I_16111 (I276410,I2507,I276048,I276013,);
DFFARX1 I_16112 (I276402,I2507,I276048,I276031,);
nor I_16113 (I276455,I1130054,I1130051);
not I_16114 (I276472,I276455);
nor I_16115 (I276034,I276311,I276472);
nand I_16116 (I276019,I276328,I276472);
nor I_16117 (I276028,I276074,I276455);
DFFARX1 I_16118 (I276455,I2507,I276048,I276037,);
not I_16119 (I276575,I2514);
DFFARX1 I_16120 (I1036511,I2507,I276575,I276601,);
nand I_16121 (I276609,I1036508,I1036511);
and I_16122 (I276626,I276609,I1036520);
DFFARX1 I_16123 (I276626,I2507,I276575,I276652,);
nor I_16124 (I276543,I276652,I276601);
not I_16125 (I276674,I276652);
DFFARX1 I_16126 (I1036508,I2507,I276575,I276700,);
nand I_16127 (I276708,I276700,I1036526);
not I_16128 (I276725,I276708);
DFFARX1 I_16129 (I276725,I2507,I276575,I276751,);
not I_16130 (I276567,I276751);
nor I_16131 (I276773,I276601,I276708);
nor I_16132 (I276549,I276652,I276773);
DFFARX1 I_16133 (I1036514,I2507,I276575,I276813,);
DFFARX1 I_16134 (I276813,I2507,I276575,I276830,);
not I_16135 (I276838,I276830);
not I_16136 (I276855,I276813);
nand I_16137 (I276552,I276855,I276674);
nand I_16138 (I276886,I1036523,I1036529);
and I_16139 (I276903,I276886,I1036514);
DFFARX1 I_16140 (I276903,I2507,I276575,I276929,);
nor I_16141 (I276937,I276929,I276601);
DFFARX1 I_16142 (I276937,I2507,I276575,I276540,);
DFFARX1 I_16143 (I276929,I2507,I276575,I276558,);
nor I_16144 (I276982,I1036517,I1036529);
not I_16145 (I276999,I276982);
nor I_16146 (I276561,I276838,I276999);
nand I_16147 (I276546,I276855,I276999);
nor I_16148 (I276555,I276601,I276982);
DFFARX1 I_16149 (I276982,I2507,I276575,I276564,);
not I_16150 (I277102,I2514);
DFFARX1 I_16151 (I78051,I2507,I277102,I277128,);
nand I_16152 (I277136,I78063,I78072);
and I_16153 (I277153,I277136,I78051);
DFFARX1 I_16154 (I277153,I2507,I277102,I277179,);
nor I_16155 (I277070,I277179,I277128);
not I_16156 (I277201,I277179);
DFFARX1 I_16157 (I78066,I2507,I277102,I277227,);
nand I_16158 (I277235,I277227,I78054);
not I_16159 (I277252,I277235);
DFFARX1 I_16160 (I277252,I2507,I277102,I277278,);
not I_16161 (I277094,I277278);
nor I_16162 (I277300,I277128,I277235);
nor I_16163 (I277076,I277179,I277300);
DFFARX1 I_16164 (I78057,I2507,I277102,I277340,);
DFFARX1 I_16165 (I277340,I2507,I277102,I277357,);
not I_16166 (I277365,I277357);
not I_16167 (I277382,I277340);
nand I_16168 (I277079,I277382,I277201);
nand I_16169 (I277413,I78048,I78048);
and I_16170 (I277430,I277413,I78060);
DFFARX1 I_16171 (I277430,I2507,I277102,I277456,);
nor I_16172 (I277464,I277456,I277128);
DFFARX1 I_16173 (I277464,I2507,I277102,I277067,);
DFFARX1 I_16174 (I277456,I2507,I277102,I277085,);
nor I_16175 (I277509,I78069,I78048);
not I_16176 (I277526,I277509);
nor I_16177 (I277088,I277365,I277526);
nand I_16178 (I277073,I277382,I277526);
nor I_16179 (I277082,I277128,I277509);
DFFARX1 I_16180 (I277509,I2507,I277102,I277091,);
not I_16181 (I277629,I2514);
DFFARX1 I_16182 (I186525,I2507,I277629,I277655,);
nand I_16183 (I277663,I186525,I186531);
and I_16184 (I277680,I277663,I186549);
DFFARX1 I_16185 (I277680,I2507,I277629,I277706,);
nor I_16186 (I277597,I277706,I277655);
not I_16187 (I277728,I277706);
DFFARX1 I_16188 (I186537,I2507,I277629,I277754,);
nand I_16189 (I277762,I277754,I186534);
not I_16190 (I277779,I277762);
DFFARX1 I_16191 (I277779,I2507,I277629,I277805,);
not I_16192 (I277621,I277805);
nor I_16193 (I277827,I277655,I277762);
nor I_16194 (I277603,I277706,I277827);
DFFARX1 I_16195 (I186543,I2507,I277629,I277867,);
DFFARX1 I_16196 (I277867,I2507,I277629,I277884,);
not I_16197 (I277892,I277884);
not I_16198 (I277909,I277867);
nand I_16199 (I277606,I277909,I277728);
nand I_16200 (I277940,I186528,I186528);
and I_16201 (I277957,I277940,I186540);
DFFARX1 I_16202 (I277957,I2507,I277629,I277983,);
nor I_16203 (I277991,I277983,I277655);
DFFARX1 I_16204 (I277991,I2507,I277629,I277594,);
DFFARX1 I_16205 (I277983,I2507,I277629,I277612,);
nor I_16206 (I278036,I186546,I186528);
not I_16207 (I278053,I278036);
nor I_16208 (I277615,I277892,I278053);
nand I_16209 (I277600,I277909,I278053);
nor I_16210 (I277609,I277655,I278036);
DFFARX1 I_16211 (I278036,I2507,I277629,I277618,);
not I_16212 (I278156,I2514);
DFFARX1 I_16213 (I453403,I2507,I278156,I278182,);
nand I_16214 (I278190,I453415,I453394);
and I_16215 (I278207,I278190,I453418);
DFFARX1 I_16216 (I278207,I2507,I278156,I278233,);
nor I_16217 (I278124,I278233,I278182);
not I_16218 (I278255,I278233);
DFFARX1 I_16219 (I453409,I2507,I278156,I278281,);
nand I_16220 (I278289,I278281,I453391);
not I_16221 (I278306,I278289);
DFFARX1 I_16222 (I278306,I2507,I278156,I278332,);
not I_16223 (I278148,I278332);
nor I_16224 (I278354,I278182,I278289);
nor I_16225 (I278130,I278233,I278354);
DFFARX1 I_16226 (I453406,I2507,I278156,I278394,);
DFFARX1 I_16227 (I278394,I2507,I278156,I278411,);
not I_16228 (I278419,I278411);
not I_16229 (I278436,I278394);
nand I_16230 (I278133,I278436,I278255);
nand I_16231 (I278467,I453391,I453397);
and I_16232 (I278484,I278467,I453400);
DFFARX1 I_16233 (I278484,I2507,I278156,I278510,);
nor I_16234 (I278518,I278510,I278182);
DFFARX1 I_16235 (I278518,I2507,I278156,I278121,);
DFFARX1 I_16236 (I278510,I2507,I278156,I278139,);
nor I_16237 (I278563,I453412,I453397);
not I_16238 (I278580,I278563);
nor I_16239 (I278142,I278419,I278580);
nand I_16240 (I278127,I278436,I278580);
nor I_16241 (I278136,I278182,I278563);
DFFARX1 I_16242 (I278563,I2507,I278156,I278145,);
not I_16243 (I278683,I2514);
DFFARX1 I_16244 (I1188998,I2507,I278683,I278709,);
nand I_16245 (I278717,I1189013,I1188998);
and I_16246 (I278734,I278717,I1189016);
DFFARX1 I_16247 (I278734,I2507,I278683,I278760,);
nor I_16248 (I278651,I278760,I278709);
not I_16249 (I278782,I278760);
DFFARX1 I_16250 (I1189022,I2507,I278683,I278808,);
nand I_16251 (I278816,I278808,I1189004);
not I_16252 (I278833,I278816);
DFFARX1 I_16253 (I278833,I2507,I278683,I278859,);
not I_16254 (I278675,I278859);
nor I_16255 (I278881,I278709,I278816);
nor I_16256 (I278657,I278760,I278881);
DFFARX1 I_16257 (I1189001,I2507,I278683,I278921,);
DFFARX1 I_16258 (I278921,I2507,I278683,I278938,);
not I_16259 (I278946,I278938);
not I_16260 (I278963,I278921);
nand I_16261 (I278660,I278963,I278782);
nand I_16262 (I278994,I1189001,I1189007);
and I_16263 (I279011,I278994,I1189019);
DFFARX1 I_16264 (I279011,I2507,I278683,I279037,);
nor I_16265 (I279045,I279037,I278709);
DFFARX1 I_16266 (I279045,I2507,I278683,I278648,);
DFFARX1 I_16267 (I279037,I2507,I278683,I278666,);
nor I_16268 (I279090,I1189010,I1189007);
not I_16269 (I279107,I279090);
nor I_16270 (I278669,I278946,I279107);
nand I_16271 (I278654,I278963,I279107);
nor I_16272 (I278663,I278709,I279090);
DFFARX1 I_16273 (I279090,I2507,I278683,I278672,);
not I_16274 (I279210,I2514);
DFFARX1 I_16275 (I1148538,I2507,I279210,I279236,);
nand I_16276 (I279244,I1148553,I1148538);
and I_16277 (I279261,I279244,I1148556);
DFFARX1 I_16278 (I279261,I2507,I279210,I279287,);
nor I_16279 (I279178,I279287,I279236);
not I_16280 (I279309,I279287);
DFFARX1 I_16281 (I1148562,I2507,I279210,I279335,);
nand I_16282 (I279343,I279335,I1148544);
not I_16283 (I279360,I279343);
DFFARX1 I_16284 (I279360,I2507,I279210,I279386,);
not I_16285 (I279202,I279386);
nor I_16286 (I279408,I279236,I279343);
nor I_16287 (I279184,I279287,I279408);
DFFARX1 I_16288 (I1148541,I2507,I279210,I279448,);
DFFARX1 I_16289 (I279448,I2507,I279210,I279465,);
not I_16290 (I279473,I279465);
not I_16291 (I279490,I279448);
nand I_16292 (I279187,I279490,I279309);
nand I_16293 (I279521,I1148541,I1148547);
and I_16294 (I279538,I279521,I1148559);
DFFARX1 I_16295 (I279538,I2507,I279210,I279564,);
nor I_16296 (I279572,I279564,I279236);
DFFARX1 I_16297 (I279572,I2507,I279210,I279175,);
DFFARX1 I_16298 (I279564,I2507,I279210,I279193,);
nor I_16299 (I279617,I1148550,I1148547);
not I_16300 (I279634,I279617);
nor I_16301 (I279196,I279473,I279634);
nand I_16302 (I279181,I279490,I279634);
nor I_16303 (I279190,I279236,I279617);
DFFARX1 I_16304 (I279617,I2507,I279210,I279199,);
not I_16305 (I279737,I2514);
DFFARX1 I_16306 (I1364238,I2507,I279737,I279763,);
nand I_16307 (I279771,I1364217,I1364217);
and I_16308 (I279788,I279771,I1364244);
DFFARX1 I_16309 (I279788,I2507,I279737,I279814,);
nor I_16310 (I279705,I279814,I279763);
not I_16311 (I279836,I279814);
DFFARX1 I_16312 (I1364232,I2507,I279737,I279862,);
nand I_16313 (I279870,I279862,I1364235);
not I_16314 (I279887,I279870);
DFFARX1 I_16315 (I279887,I2507,I279737,I279913,);
not I_16316 (I279729,I279913);
nor I_16317 (I279935,I279763,I279870);
nor I_16318 (I279711,I279814,I279935);
DFFARX1 I_16319 (I1364226,I2507,I279737,I279975,);
DFFARX1 I_16320 (I279975,I2507,I279737,I279992,);
not I_16321 (I280000,I279992);
not I_16322 (I280017,I279975);
nand I_16323 (I279714,I280017,I279836);
nand I_16324 (I280048,I1364223,I1364220);
and I_16325 (I280065,I280048,I1364241);
DFFARX1 I_16326 (I280065,I2507,I279737,I280091,);
nor I_16327 (I280099,I280091,I279763);
DFFARX1 I_16328 (I280099,I2507,I279737,I279702,);
DFFARX1 I_16329 (I280091,I2507,I279737,I279720,);
nor I_16330 (I280144,I1364229,I1364220);
not I_16331 (I280161,I280144);
nor I_16332 (I279723,I280000,I280161);
nand I_16333 (I279708,I280017,I280161);
nor I_16334 (I279717,I279763,I280144);
DFFARX1 I_16335 (I280144,I2507,I279737,I279726,);
not I_16336 (I280264,I2514);
DFFARX1 I_16337 (I832817,I2507,I280264,I280290,);
nand I_16338 (I280298,I832820,I832814);
and I_16339 (I280315,I280298,I832826);
DFFARX1 I_16340 (I280315,I2507,I280264,I280341,);
nor I_16341 (I280232,I280341,I280290);
not I_16342 (I280363,I280341);
DFFARX1 I_16343 (I832829,I2507,I280264,I280389,);
nand I_16344 (I280397,I280389,I832820);
not I_16345 (I280414,I280397);
DFFARX1 I_16346 (I280414,I2507,I280264,I280440,);
not I_16347 (I280256,I280440);
nor I_16348 (I280462,I280290,I280397);
nor I_16349 (I280238,I280341,I280462);
DFFARX1 I_16350 (I832832,I2507,I280264,I280502,);
DFFARX1 I_16351 (I280502,I2507,I280264,I280519,);
not I_16352 (I280527,I280519);
not I_16353 (I280544,I280502);
nand I_16354 (I280241,I280544,I280363);
nand I_16355 (I280575,I832814,I832823);
and I_16356 (I280592,I280575,I832817);
DFFARX1 I_16357 (I280592,I2507,I280264,I280618,);
nor I_16358 (I280626,I280618,I280290);
DFFARX1 I_16359 (I280626,I2507,I280264,I280229,);
DFFARX1 I_16360 (I280618,I2507,I280264,I280247,);
nor I_16361 (I280671,I832835,I832823);
not I_16362 (I280688,I280671);
nor I_16363 (I280250,I280527,I280688);
nand I_16364 (I280235,I280544,I280688);
nor I_16365 (I280244,I280290,I280671);
DFFARX1 I_16366 (I280671,I2507,I280264,I280253,);
not I_16367 (I280791,I2514);
DFFARX1 I_16368 (I131278,I2507,I280791,I280817,);
nand I_16369 (I280825,I131290,I131299);
and I_16370 (I280842,I280825,I131278);
DFFARX1 I_16371 (I280842,I2507,I280791,I280868,);
nor I_16372 (I280759,I280868,I280817);
not I_16373 (I280890,I280868);
DFFARX1 I_16374 (I131293,I2507,I280791,I280916,);
nand I_16375 (I280924,I280916,I131281);
not I_16376 (I280941,I280924);
DFFARX1 I_16377 (I280941,I2507,I280791,I280967,);
not I_16378 (I280783,I280967);
nor I_16379 (I280989,I280817,I280924);
nor I_16380 (I280765,I280868,I280989);
DFFARX1 I_16381 (I131284,I2507,I280791,I281029,);
DFFARX1 I_16382 (I281029,I2507,I280791,I281046,);
not I_16383 (I281054,I281046);
not I_16384 (I281071,I281029);
nand I_16385 (I280768,I281071,I280890);
nand I_16386 (I281102,I131275,I131275);
and I_16387 (I281119,I281102,I131287);
DFFARX1 I_16388 (I281119,I2507,I280791,I281145,);
nor I_16389 (I281153,I281145,I280817);
DFFARX1 I_16390 (I281153,I2507,I280791,I280756,);
DFFARX1 I_16391 (I281145,I2507,I280791,I280774,);
nor I_16392 (I281198,I131296,I131275);
not I_16393 (I281215,I281198);
nor I_16394 (I280777,I281054,I281215);
nand I_16395 (I280762,I281071,I281215);
nor I_16396 (I280771,I280817,I281198);
DFFARX1 I_16397 (I281198,I2507,I280791,I280780,);
not I_16398 (I281318,I2514);
DFFARX1 I_16399 (I683328,I2507,I281318,I281344,);
nand I_16400 (I281352,I683319,I683334);
and I_16401 (I281369,I281352,I683340);
DFFARX1 I_16402 (I281369,I2507,I281318,I281395,);
nor I_16403 (I281286,I281395,I281344);
not I_16404 (I281417,I281395);
DFFARX1 I_16405 (I683325,I2507,I281318,I281443,);
nand I_16406 (I281451,I281443,I683319);
not I_16407 (I281468,I281451);
DFFARX1 I_16408 (I281468,I2507,I281318,I281494,);
not I_16409 (I281310,I281494);
nor I_16410 (I281516,I281344,I281451);
nor I_16411 (I281292,I281395,I281516);
DFFARX1 I_16412 (I683322,I2507,I281318,I281556,);
DFFARX1 I_16413 (I281556,I2507,I281318,I281573,);
not I_16414 (I281581,I281573);
not I_16415 (I281598,I281556);
nand I_16416 (I281295,I281598,I281417);
nand I_16417 (I281629,I683316,I683331);
and I_16418 (I281646,I281629,I683316);
DFFARX1 I_16419 (I281646,I2507,I281318,I281672,);
nor I_16420 (I281680,I281672,I281344);
DFFARX1 I_16421 (I281680,I2507,I281318,I281283,);
DFFARX1 I_16422 (I281672,I2507,I281318,I281301,);
nor I_16423 (I281725,I683337,I683331);
not I_16424 (I281742,I281725);
nor I_16425 (I281304,I281581,I281742);
nand I_16426 (I281289,I281598,I281742);
nor I_16427 (I281298,I281344,I281725);
DFFARX1 I_16428 (I281725,I2507,I281318,I281307,);
not I_16429 (I281845,I2514);
DFFARX1 I_16430 (I791184,I2507,I281845,I281871,);
nand I_16431 (I281879,I791187,I791181);
and I_16432 (I281896,I281879,I791193);
DFFARX1 I_16433 (I281896,I2507,I281845,I281922,);
nor I_16434 (I281813,I281922,I281871);
not I_16435 (I281944,I281922);
DFFARX1 I_16436 (I791196,I2507,I281845,I281970,);
nand I_16437 (I281978,I281970,I791187);
not I_16438 (I281995,I281978);
DFFARX1 I_16439 (I281995,I2507,I281845,I282021,);
not I_16440 (I281837,I282021);
nor I_16441 (I282043,I281871,I281978);
nor I_16442 (I281819,I281922,I282043);
DFFARX1 I_16443 (I791199,I2507,I281845,I282083,);
DFFARX1 I_16444 (I282083,I2507,I281845,I282100,);
not I_16445 (I282108,I282100);
not I_16446 (I282125,I282083);
nand I_16447 (I281822,I282125,I281944);
nand I_16448 (I282156,I791181,I791190);
and I_16449 (I282173,I282156,I791184);
DFFARX1 I_16450 (I282173,I2507,I281845,I282199,);
nor I_16451 (I282207,I282199,I281871);
DFFARX1 I_16452 (I282207,I2507,I281845,I281810,);
DFFARX1 I_16453 (I282199,I2507,I281845,I281828,);
nor I_16454 (I282252,I791202,I791190);
not I_16455 (I282269,I282252);
nor I_16456 (I281831,I282108,I282269);
nand I_16457 (I281816,I282125,I282269);
nor I_16458 (I281825,I281871,I282252);
DFFARX1 I_16459 (I282252,I2507,I281845,I281834,);
not I_16460 (I282372,I2514);
DFFARX1 I_16461 (I637088,I2507,I282372,I282398,);
nand I_16462 (I282406,I637079,I637094);
and I_16463 (I282423,I282406,I637100);
DFFARX1 I_16464 (I282423,I2507,I282372,I282449,);
nor I_16465 (I282340,I282449,I282398);
not I_16466 (I282471,I282449);
DFFARX1 I_16467 (I637085,I2507,I282372,I282497,);
nand I_16468 (I282505,I282497,I637079);
not I_16469 (I282522,I282505);
DFFARX1 I_16470 (I282522,I2507,I282372,I282548,);
not I_16471 (I282364,I282548);
nor I_16472 (I282570,I282398,I282505);
nor I_16473 (I282346,I282449,I282570);
DFFARX1 I_16474 (I637082,I2507,I282372,I282610,);
DFFARX1 I_16475 (I282610,I2507,I282372,I282627,);
not I_16476 (I282635,I282627);
not I_16477 (I282652,I282610);
nand I_16478 (I282349,I282652,I282471);
nand I_16479 (I282683,I637076,I637091);
and I_16480 (I282700,I282683,I637076);
DFFARX1 I_16481 (I282700,I2507,I282372,I282726,);
nor I_16482 (I282734,I282726,I282398);
DFFARX1 I_16483 (I282734,I2507,I282372,I282337,);
DFFARX1 I_16484 (I282726,I2507,I282372,I282355,);
nor I_16485 (I282779,I637097,I637091);
not I_16486 (I282796,I282779);
nor I_16487 (I282358,I282635,I282796);
nand I_16488 (I282343,I282652,I282796);
nor I_16489 (I282352,I282398,I282779);
DFFARX1 I_16490 (I282779,I2507,I282372,I282361,);
not I_16491 (I282899,I2514);
DFFARX1 I_16492 (I738816,I2507,I282899,I282925,);
nand I_16493 (I282933,I738807,I738822);
and I_16494 (I282950,I282933,I738828);
DFFARX1 I_16495 (I282950,I2507,I282899,I282976,);
nor I_16496 (I282867,I282976,I282925);
not I_16497 (I282998,I282976);
DFFARX1 I_16498 (I738813,I2507,I282899,I283024,);
nand I_16499 (I283032,I283024,I738807);
not I_16500 (I283049,I283032);
DFFARX1 I_16501 (I283049,I2507,I282899,I283075,);
not I_16502 (I282891,I283075);
nor I_16503 (I283097,I282925,I283032);
nor I_16504 (I282873,I282976,I283097);
DFFARX1 I_16505 (I738810,I2507,I282899,I283137,);
DFFARX1 I_16506 (I283137,I2507,I282899,I283154,);
not I_16507 (I283162,I283154);
not I_16508 (I283179,I283137);
nand I_16509 (I282876,I283179,I282998);
nand I_16510 (I283210,I738804,I738819);
and I_16511 (I283227,I283210,I738804);
DFFARX1 I_16512 (I283227,I2507,I282899,I283253,);
nor I_16513 (I283261,I283253,I282925);
DFFARX1 I_16514 (I283261,I2507,I282899,I282864,);
DFFARX1 I_16515 (I283253,I2507,I282899,I282882,);
nor I_16516 (I283306,I738825,I738819);
not I_16517 (I283323,I283306);
nor I_16518 (I282885,I283162,I283323);
nand I_16519 (I282870,I283179,I283323);
nor I_16520 (I282879,I282925,I283306);
DFFARX1 I_16521 (I283306,I2507,I282899,I282888,);
not I_16522 (I283426,I2514);
DFFARX1 I_16523 (I45374,I2507,I283426,I283452,);
nand I_16524 (I283460,I45398,I45377);
and I_16525 (I283477,I283460,I45374);
DFFARX1 I_16526 (I283477,I2507,I283426,I283503,);
nor I_16527 (I283394,I283503,I283452);
not I_16528 (I283525,I283503);
DFFARX1 I_16529 (I45380,I2507,I283426,I283551,);
nand I_16530 (I283559,I283551,I45389);
not I_16531 (I283576,I283559);
DFFARX1 I_16532 (I283576,I2507,I283426,I283602,);
not I_16533 (I283418,I283602);
nor I_16534 (I283624,I283452,I283559);
nor I_16535 (I283400,I283503,I283624);
DFFARX1 I_16536 (I45383,I2507,I283426,I283664,);
DFFARX1 I_16537 (I283664,I2507,I283426,I283681,);
not I_16538 (I283689,I283681);
not I_16539 (I283706,I283664);
nand I_16540 (I283403,I283706,I283525);
nand I_16541 (I283737,I45395,I45377);
and I_16542 (I283754,I283737,I45386);
DFFARX1 I_16543 (I283754,I2507,I283426,I283780,);
nor I_16544 (I283788,I283780,I283452);
DFFARX1 I_16545 (I283788,I2507,I283426,I283391,);
DFFARX1 I_16546 (I283780,I2507,I283426,I283409,);
nor I_16547 (I283833,I45392,I45377);
not I_16548 (I283850,I283833);
nor I_16549 (I283412,I283689,I283850);
nand I_16550 (I283397,I283706,I283850);
nor I_16551 (I283406,I283452,I283833);
DFFARX1 I_16552 (I283833,I2507,I283426,I283415,);
not I_16553 (I283953,I2514);
DFFARX1 I_16554 (I1179172,I2507,I283953,I283979,);
nand I_16555 (I283987,I1179187,I1179172);
and I_16556 (I284004,I283987,I1179190);
DFFARX1 I_16557 (I284004,I2507,I283953,I284030,);
nor I_16558 (I283921,I284030,I283979);
not I_16559 (I284052,I284030);
DFFARX1 I_16560 (I1179196,I2507,I283953,I284078,);
nand I_16561 (I284086,I284078,I1179178);
not I_16562 (I284103,I284086);
DFFARX1 I_16563 (I284103,I2507,I283953,I284129,);
not I_16564 (I283945,I284129);
nor I_16565 (I284151,I283979,I284086);
nor I_16566 (I283927,I284030,I284151);
DFFARX1 I_16567 (I1179175,I2507,I283953,I284191,);
DFFARX1 I_16568 (I284191,I2507,I283953,I284208,);
not I_16569 (I284216,I284208);
not I_16570 (I284233,I284191);
nand I_16571 (I283930,I284233,I284052);
nand I_16572 (I284264,I1179175,I1179181);
and I_16573 (I284281,I284264,I1179193);
DFFARX1 I_16574 (I284281,I2507,I283953,I284307,);
nor I_16575 (I284315,I284307,I283979);
DFFARX1 I_16576 (I284315,I2507,I283953,I283918,);
DFFARX1 I_16577 (I284307,I2507,I283953,I283936,);
nor I_16578 (I284360,I1179184,I1179181);
not I_16579 (I284377,I284360);
nor I_16580 (I283939,I284216,I284377);
nand I_16581 (I283924,I284233,I284377);
nor I_16582 (I283933,I283979,I284360);
DFFARX1 I_16583 (I284360,I2507,I283953,I283942,);
not I_16584 (I284480,I2514);
DFFARX1 I_16585 (I1097096,I2507,I284480,I284506,);
nand I_16586 (I284514,I1097111,I1097096);
and I_16587 (I284531,I284514,I1097114);
DFFARX1 I_16588 (I284531,I2507,I284480,I284557,);
nor I_16589 (I284448,I284557,I284506);
not I_16590 (I284579,I284557);
DFFARX1 I_16591 (I1097120,I2507,I284480,I284605,);
nand I_16592 (I284613,I284605,I1097102);
not I_16593 (I284630,I284613);
DFFARX1 I_16594 (I284630,I2507,I284480,I284656,);
not I_16595 (I284472,I284656);
nor I_16596 (I284678,I284506,I284613);
nor I_16597 (I284454,I284557,I284678);
DFFARX1 I_16598 (I1097099,I2507,I284480,I284718,);
DFFARX1 I_16599 (I284718,I2507,I284480,I284735,);
not I_16600 (I284743,I284735);
not I_16601 (I284760,I284718);
nand I_16602 (I284457,I284760,I284579);
nand I_16603 (I284791,I1097099,I1097105);
and I_16604 (I284808,I284791,I1097117);
DFFARX1 I_16605 (I284808,I2507,I284480,I284834,);
nor I_16606 (I284842,I284834,I284506);
DFFARX1 I_16607 (I284842,I2507,I284480,I284445,);
DFFARX1 I_16608 (I284834,I2507,I284480,I284463,);
nor I_16609 (I284887,I1097108,I1097105);
not I_16610 (I284904,I284887);
nor I_16611 (I284466,I284743,I284904);
nand I_16612 (I284451,I284760,I284904);
nor I_16613 (I284460,I284506,I284887);
DFFARX1 I_16614 (I284887,I2507,I284480,I284469,);
not I_16615 (I285007,I2514);
DFFARX1 I_16616 (I237100,I2507,I285007,I285033,);
nand I_16617 (I285041,I237100,I237106);
and I_16618 (I285058,I285041,I237124);
DFFARX1 I_16619 (I285058,I2507,I285007,I285084,);
nor I_16620 (I284975,I285084,I285033);
not I_16621 (I285106,I285084);
DFFARX1 I_16622 (I237112,I2507,I285007,I285132,);
nand I_16623 (I285140,I285132,I237109);
not I_16624 (I285157,I285140);
DFFARX1 I_16625 (I285157,I2507,I285007,I285183,);
not I_16626 (I284999,I285183);
nor I_16627 (I285205,I285033,I285140);
nor I_16628 (I284981,I285084,I285205);
DFFARX1 I_16629 (I237118,I2507,I285007,I285245,);
DFFARX1 I_16630 (I285245,I2507,I285007,I285262,);
not I_16631 (I285270,I285262);
not I_16632 (I285287,I285245);
nand I_16633 (I284984,I285287,I285106);
nand I_16634 (I285318,I237103,I237103);
and I_16635 (I285335,I285318,I237115);
DFFARX1 I_16636 (I285335,I2507,I285007,I285361,);
nor I_16637 (I285369,I285361,I285033);
DFFARX1 I_16638 (I285369,I2507,I285007,I284972,);
DFFARX1 I_16639 (I285361,I2507,I285007,I284990,);
nor I_16640 (I285414,I237121,I237103);
not I_16641 (I285431,I285414);
nor I_16642 (I284993,I285270,I285431);
nand I_16643 (I284978,I285287,I285431);
nor I_16644 (I284987,I285033,I285414);
DFFARX1 I_16645 (I285414,I2507,I285007,I284996,);
not I_16646 (I285534,I2514);
DFFARX1 I_16647 (I1199980,I2507,I285534,I285560,);
nand I_16648 (I285568,I1199995,I1199980);
and I_16649 (I285585,I285568,I1199998);
DFFARX1 I_16650 (I285585,I2507,I285534,I285611,);
nor I_16651 (I285502,I285611,I285560);
not I_16652 (I285633,I285611);
DFFARX1 I_16653 (I1200004,I2507,I285534,I285659,);
nand I_16654 (I285667,I285659,I1199986);
not I_16655 (I285684,I285667);
DFFARX1 I_16656 (I285684,I2507,I285534,I285710,);
not I_16657 (I285526,I285710);
nor I_16658 (I285732,I285560,I285667);
nor I_16659 (I285508,I285611,I285732);
DFFARX1 I_16660 (I1199983,I2507,I285534,I285772,);
DFFARX1 I_16661 (I285772,I2507,I285534,I285789,);
not I_16662 (I285797,I285789);
not I_16663 (I285814,I285772);
nand I_16664 (I285511,I285814,I285633);
nand I_16665 (I285845,I1199983,I1199989);
and I_16666 (I285862,I285845,I1200001);
DFFARX1 I_16667 (I285862,I2507,I285534,I285888,);
nor I_16668 (I285896,I285888,I285560);
DFFARX1 I_16669 (I285896,I2507,I285534,I285499,);
DFFARX1 I_16670 (I285888,I2507,I285534,I285517,);
nor I_16671 (I285941,I1199992,I1199989);
not I_16672 (I285958,I285941);
nor I_16673 (I285520,I285797,I285958);
nand I_16674 (I285505,I285814,I285958);
nor I_16675 (I285514,I285560,I285941);
DFFARX1 I_16676 (I285941,I2507,I285534,I285523,);
not I_16677 (I286061,I2514);
DFFARX1 I_16678 (I480603,I2507,I286061,I286087,);
nand I_16679 (I286095,I480615,I480594);
and I_16680 (I286112,I286095,I480618);
DFFARX1 I_16681 (I286112,I2507,I286061,I286138,);
nor I_16682 (I286029,I286138,I286087);
not I_16683 (I286160,I286138);
DFFARX1 I_16684 (I480609,I2507,I286061,I286186,);
nand I_16685 (I286194,I286186,I480591);
not I_16686 (I286211,I286194);
DFFARX1 I_16687 (I286211,I2507,I286061,I286237,);
not I_16688 (I286053,I286237);
nor I_16689 (I286259,I286087,I286194);
nor I_16690 (I286035,I286138,I286259);
DFFARX1 I_16691 (I480606,I2507,I286061,I286299,);
DFFARX1 I_16692 (I286299,I2507,I286061,I286316,);
not I_16693 (I286324,I286316);
not I_16694 (I286341,I286299);
nand I_16695 (I286038,I286341,I286160);
nand I_16696 (I286372,I480591,I480597);
and I_16697 (I286389,I286372,I480600);
DFFARX1 I_16698 (I286389,I2507,I286061,I286415,);
nor I_16699 (I286423,I286415,I286087);
DFFARX1 I_16700 (I286423,I2507,I286061,I286026,);
DFFARX1 I_16701 (I286415,I2507,I286061,I286044,);
nor I_16702 (I286468,I480612,I480597);
not I_16703 (I286485,I286468);
nor I_16704 (I286047,I286324,I286485);
nand I_16705 (I286032,I286341,I286485);
nor I_16706 (I286041,I286087,I286468);
DFFARX1 I_16707 (I286468,I2507,I286061,I286050,);
not I_16708 (I286588,I2514);
DFFARX1 I_16709 (I1288293,I2507,I286588,I286614,);
nand I_16710 (I286622,I1288290,I1288281);
and I_16711 (I286639,I286622,I1288278);
DFFARX1 I_16712 (I286639,I2507,I286588,I286665,);
nor I_16713 (I286556,I286665,I286614);
not I_16714 (I286687,I286665);
DFFARX1 I_16715 (I1288287,I2507,I286588,I286713,);
nand I_16716 (I286721,I286713,I1288296);
not I_16717 (I286738,I286721);
DFFARX1 I_16718 (I286738,I2507,I286588,I286764,);
not I_16719 (I286580,I286764);
nor I_16720 (I286786,I286614,I286721);
nor I_16721 (I286562,I286665,I286786);
DFFARX1 I_16722 (I1288299,I2507,I286588,I286826,);
DFFARX1 I_16723 (I286826,I2507,I286588,I286843,);
not I_16724 (I286851,I286843);
not I_16725 (I286868,I286826);
nand I_16726 (I286565,I286868,I286687);
nand I_16727 (I286899,I1288278,I1288284);
and I_16728 (I286916,I286899,I1288302);
DFFARX1 I_16729 (I286916,I2507,I286588,I286942,);
nor I_16730 (I286950,I286942,I286614);
DFFARX1 I_16731 (I286950,I2507,I286588,I286553,);
DFFARX1 I_16732 (I286942,I2507,I286588,I286571,);
nor I_16733 (I286995,I1288281,I1288284);
not I_16734 (I287012,I286995);
nor I_16735 (I286574,I286851,I287012);
nand I_16736 (I286559,I286868,I287012);
nor I_16737 (I286568,I286614,I286995);
DFFARX1 I_16738 (I286995,I2507,I286588,I286577,);
not I_16739 (I287115,I2514);
DFFARX1 I_16740 (I1030340,I2507,I287115,I287141,);
nand I_16741 (I287149,I1030337,I1030340);
and I_16742 (I287166,I287149,I1030349);
DFFARX1 I_16743 (I287166,I2507,I287115,I287192,);
nor I_16744 (I287083,I287192,I287141);
not I_16745 (I287214,I287192);
DFFARX1 I_16746 (I1030337,I2507,I287115,I287240,);
nand I_16747 (I287248,I287240,I1030355);
not I_16748 (I287265,I287248);
DFFARX1 I_16749 (I287265,I2507,I287115,I287291,);
not I_16750 (I287107,I287291);
nor I_16751 (I287313,I287141,I287248);
nor I_16752 (I287089,I287192,I287313);
DFFARX1 I_16753 (I1030343,I2507,I287115,I287353,);
DFFARX1 I_16754 (I287353,I2507,I287115,I287370,);
not I_16755 (I287378,I287370);
not I_16756 (I287395,I287353);
nand I_16757 (I287092,I287395,I287214);
nand I_16758 (I287426,I1030352,I1030358);
and I_16759 (I287443,I287426,I1030343);
DFFARX1 I_16760 (I287443,I2507,I287115,I287469,);
nor I_16761 (I287477,I287469,I287141);
DFFARX1 I_16762 (I287477,I2507,I287115,I287080,);
DFFARX1 I_16763 (I287469,I2507,I287115,I287098,);
nor I_16764 (I287522,I1030346,I1030358);
not I_16765 (I287539,I287522);
nor I_16766 (I287101,I287378,I287539);
nand I_16767 (I287086,I287395,I287539);
nor I_16768 (I287095,I287141,I287522);
DFFARX1 I_16769 (I287522,I2507,I287115,I287104,);
not I_16770 (I287642,I2514);
DFFARX1 I_16771 (I456123,I2507,I287642,I287668,);
nand I_16772 (I287676,I456135,I456114);
and I_16773 (I287693,I287676,I456138);
DFFARX1 I_16774 (I287693,I2507,I287642,I287719,);
nor I_16775 (I287610,I287719,I287668);
not I_16776 (I287741,I287719);
DFFARX1 I_16777 (I456129,I2507,I287642,I287767,);
nand I_16778 (I287775,I287767,I456111);
not I_16779 (I287792,I287775);
DFFARX1 I_16780 (I287792,I2507,I287642,I287818,);
not I_16781 (I287634,I287818);
nor I_16782 (I287840,I287668,I287775);
nor I_16783 (I287616,I287719,I287840);
DFFARX1 I_16784 (I456126,I2507,I287642,I287880,);
DFFARX1 I_16785 (I287880,I2507,I287642,I287897,);
not I_16786 (I287905,I287897);
not I_16787 (I287922,I287880);
nand I_16788 (I287619,I287922,I287741);
nand I_16789 (I287953,I456111,I456117);
and I_16790 (I287970,I287953,I456120);
DFFARX1 I_16791 (I287970,I2507,I287642,I287996,);
nor I_16792 (I288004,I287996,I287668);
DFFARX1 I_16793 (I288004,I2507,I287642,I287607,);
DFFARX1 I_16794 (I287996,I2507,I287642,I287625,);
nor I_16795 (I288049,I456132,I456117);
not I_16796 (I288066,I288049);
nor I_16797 (I287628,I287905,I288066);
nand I_16798 (I287613,I287922,I288066);
nor I_16799 (I287622,I287668,I288049);
DFFARX1 I_16800 (I288049,I2507,I287642,I287631,);
not I_16801 (I288169,I2514);
DFFARX1 I_16802 (I1123684,I2507,I288169,I288195,);
nand I_16803 (I288203,I1123699,I1123684);
and I_16804 (I288220,I288203,I1123702);
DFFARX1 I_16805 (I288220,I2507,I288169,I288246,);
nor I_16806 (I288137,I288246,I288195);
not I_16807 (I288268,I288246);
DFFARX1 I_16808 (I1123708,I2507,I288169,I288294,);
nand I_16809 (I288302,I288294,I1123690);
not I_16810 (I288319,I288302);
DFFARX1 I_16811 (I288319,I2507,I288169,I288345,);
not I_16812 (I288161,I288345);
nor I_16813 (I288367,I288195,I288302);
nor I_16814 (I288143,I288246,I288367);
DFFARX1 I_16815 (I1123687,I2507,I288169,I288407,);
DFFARX1 I_16816 (I288407,I2507,I288169,I288424,);
not I_16817 (I288432,I288424);
not I_16818 (I288449,I288407);
nand I_16819 (I288146,I288449,I288268);
nand I_16820 (I288480,I1123687,I1123693);
and I_16821 (I288497,I288480,I1123705);
DFFARX1 I_16822 (I288497,I2507,I288169,I288523,);
nor I_16823 (I288531,I288523,I288195);
DFFARX1 I_16824 (I288531,I2507,I288169,I288134,);
DFFARX1 I_16825 (I288523,I2507,I288169,I288152,);
nor I_16826 (I288576,I1123696,I1123693);
not I_16827 (I288593,I288576);
nor I_16828 (I288155,I288432,I288593);
nand I_16829 (I288140,I288449,I288593);
nor I_16830 (I288149,I288195,I288576);
DFFARX1 I_16831 (I288576,I2507,I288169,I288158,);
not I_16832 (I288696,I2514);
DFFARX1 I_16833 (I792238,I2507,I288696,I288722,);
nand I_16834 (I288730,I792241,I792235);
and I_16835 (I288747,I288730,I792247);
DFFARX1 I_16836 (I288747,I2507,I288696,I288773,);
nor I_16837 (I288664,I288773,I288722);
not I_16838 (I288795,I288773);
DFFARX1 I_16839 (I792250,I2507,I288696,I288821,);
nand I_16840 (I288829,I288821,I792241);
not I_16841 (I288846,I288829);
DFFARX1 I_16842 (I288846,I2507,I288696,I288872,);
not I_16843 (I288688,I288872);
nor I_16844 (I288894,I288722,I288829);
nor I_16845 (I288670,I288773,I288894);
DFFARX1 I_16846 (I792253,I2507,I288696,I288934,);
DFFARX1 I_16847 (I288934,I2507,I288696,I288951,);
not I_16848 (I288959,I288951);
not I_16849 (I288976,I288934);
nand I_16850 (I288673,I288976,I288795);
nand I_16851 (I289007,I792235,I792244);
and I_16852 (I289024,I289007,I792238);
DFFARX1 I_16853 (I289024,I2507,I288696,I289050,);
nor I_16854 (I289058,I289050,I288722);
DFFARX1 I_16855 (I289058,I2507,I288696,I288661,);
DFFARX1 I_16856 (I289050,I2507,I288696,I288679,);
nor I_16857 (I289103,I792256,I792244);
not I_16858 (I289120,I289103);
nor I_16859 (I288682,I288959,I289120);
nand I_16860 (I288667,I288976,I289120);
nor I_16861 (I288676,I288722,I289103);
DFFARX1 I_16862 (I289103,I2507,I288696,I288685,);
not I_16863 (I289223,I2514);
DFFARX1 I_16864 (I2220,I2507,I289223,I289249,);
nand I_16865 (I289257,I2380,I1652);
and I_16866 (I289274,I289257,I1956);
DFFARX1 I_16867 (I289274,I2507,I289223,I289300,);
nor I_16868 (I289191,I289300,I289249);
not I_16869 (I289322,I289300);
DFFARX1 I_16870 (I2132,I2507,I289223,I289348,);
nand I_16871 (I289356,I289348,I2428);
not I_16872 (I289373,I289356);
DFFARX1 I_16873 (I289373,I2507,I289223,I289399,);
not I_16874 (I289215,I289399);
nor I_16875 (I289421,I289249,I289356);
nor I_16876 (I289197,I289300,I289421);
DFFARX1 I_16877 (I1572,I2507,I289223,I289461,);
DFFARX1 I_16878 (I289461,I2507,I289223,I289478,);
not I_16879 (I289486,I289478);
not I_16880 (I289503,I289461);
nand I_16881 (I289200,I289503,I289322);
nand I_16882 (I289534,I2492,I2420);
and I_16883 (I289551,I289534,I1628);
DFFARX1 I_16884 (I289551,I2507,I289223,I289577,);
nor I_16885 (I289585,I289577,I289249);
DFFARX1 I_16886 (I289585,I2507,I289223,I289188,);
DFFARX1 I_16887 (I289577,I2507,I289223,I289206,);
nor I_16888 (I289630,I1620,I2420);
not I_16889 (I289647,I289630);
nor I_16890 (I289209,I289486,I289647);
nand I_16891 (I289194,I289503,I289647);
nor I_16892 (I289203,I289249,I289630);
DFFARX1 I_16893 (I289630,I2507,I289223,I289212,);
not I_16894 (I289750,I2514);
DFFARX1 I_16895 (I400635,I2507,I289750,I289776,);
nand I_16896 (I289784,I400647,I400626);
and I_16897 (I289801,I289784,I400650);
DFFARX1 I_16898 (I289801,I2507,I289750,I289827,);
nor I_16899 (I289718,I289827,I289776);
not I_16900 (I289849,I289827);
DFFARX1 I_16901 (I400641,I2507,I289750,I289875,);
nand I_16902 (I289883,I289875,I400623);
not I_16903 (I289900,I289883);
DFFARX1 I_16904 (I289900,I2507,I289750,I289926,);
not I_16905 (I289742,I289926);
nor I_16906 (I289948,I289776,I289883);
nor I_16907 (I289724,I289827,I289948);
DFFARX1 I_16908 (I400638,I2507,I289750,I289988,);
DFFARX1 I_16909 (I289988,I2507,I289750,I290005,);
not I_16910 (I290013,I290005);
not I_16911 (I290030,I289988);
nand I_16912 (I289727,I290030,I289849);
nand I_16913 (I290061,I400623,I400629);
and I_16914 (I290078,I290061,I400632);
DFFARX1 I_16915 (I290078,I2507,I289750,I290104,);
nor I_16916 (I290112,I290104,I289776);
DFFARX1 I_16917 (I290112,I2507,I289750,I289715,);
DFFARX1 I_16918 (I290104,I2507,I289750,I289733,);
nor I_16919 (I290157,I400644,I400629);
not I_16920 (I290174,I290157);
nor I_16921 (I289736,I290013,I290174);
nand I_16922 (I289721,I290030,I290174);
nor I_16923 (I289730,I289776,I290157);
DFFARX1 I_16924 (I290157,I2507,I289750,I289739,);
not I_16925 (I290277,I2514);
DFFARX1 I_16926 (I891450,I2507,I290277,I290303,);
nand I_16927 (I290311,I891447,I891465);
and I_16928 (I290328,I290311,I891456);
DFFARX1 I_16929 (I290328,I2507,I290277,I290354,);
nor I_16930 (I290245,I290354,I290303);
not I_16931 (I290376,I290354);
DFFARX1 I_16932 (I891471,I2507,I290277,I290402,);
nand I_16933 (I290410,I290402,I891453);
not I_16934 (I290427,I290410);
DFFARX1 I_16935 (I290427,I2507,I290277,I290453,);
not I_16936 (I290269,I290453);
nor I_16937 (I290475,I290303,I290410);
nor I_16938 (I290251,I290354,I290475);
DFFARX1 I_16939 (I891459,I2507,I290277,I290515,);
DFFARX1 I_16940 (I290515,I2507,I290277,I290532,);
not I_16941 (I290540,I290532);
not I_16942 (I290557,I290515);
nand I_16943 (I290254,I290557,I290376);
nand I_16944 (I290588,I891447,I891474);
and I_16945 (I290605,I290588,I891462);
DFFARX1 I_16946 (I290605,I2507,I290277,I290631,);
nor I_16947 (I290639,I290631,I290303);
DFFARX1 I_16948 (I290639,I2507,I290277,I290242,);
DFFARX1 I_16949 (I290631,I2507,I290277,I290260,);
nor I_16950 (I290684,I891468,I891474);
not I_16951 (I290701,I290684);
nor I_16952 (I290263,I290540,I290701);
nand I_16953 (I290248,I290557,I290701);
nor I_16954 (I290257,I290303,I290684);
DFFARX1 I_16955 (I290684,I2507,I290277,I290266,);
not I_16956 (I290804,I2514);
DFFARX1 I_16957 (I462107,I2507,I290804,I290830,);
nand I_16958 (I290838,I462119,I462098);
and I_16959 (I290855,I290838,I462122);
DFFARX1 I_16960 (I290855,I2507,I290804,I290881,);
nor I_16961 (I290772,I290881,I290830);
not I_16962 (I290903,I290881);
DFFARX1 I_16963 (I462113,I2507,I290804,I290929,);
nand I_16964 (I290937,I290929,I462095);
not I_16965 (I290954,I290937);
DFFARX1 I_16966 (I290954,I2507,I290804,I290980,);
not I_16967 (I290796,I290980);
nor I_16968 (I291002,I290830,I290937);
nor I_16969 (I290778,I290881,I291002);
DFFARX1 I_16970 (I462110,I2507,I290804,I291042,);
DFFARX1 I_16971 (I291042,I2507,I290804,I291059,);
not I_16972 (I291067,I291059);
not I_16973 (I291084,I291042);
nand I_16974 (I290781,I291084,I290903);
nand I_16975 (I291115,I462095,I462101);
and I_16976 (I291132,I291115,I462104);
DFFARX1 I_16977 (I291132,I2507,I290804,I291158,);
nor I_16978 (I291166,I291158,I290830);
DFFARX1 I_16979 (I291166,I2507,I290804,I290769,);
DFFARX1 I_16980 (I291158,I2507,I290804,I290787,);
nor I_16981 (I291211,I462116,I462101);
not I_16982 (I291228,I291211);
nor I_16983 (I290790,I291067,I291228);
nand I_16984 (I290775,I291084,I291228);
nor I_16985 (I290784,I290830,I291211);
DFFARX1 I_16986 (I291211,I2507,I290804,I290793,);
not I_16987 (I291331,I2514);
DFFARX1 I_16988 (I843357,I2507,I291331,I291357,);
nand I_16989 (I291365,I843360,I843354);
and I_16990 (I291382,I291365,I843366);
DFFARX1 I_16991 (I291382,I2507,I291331,I291408,);
nor I_16992 (I291299,I291408,I291357);
not I_16993 (I291430,I291408);
DFFARX1 I_16994 (I843369,I2507,I291331,I291456,);
nand I_16995 (I291464,I291456,I843360);
not I_16996 (I291481,I291464);
DFFARX1 I_16997 (I291481,I2507,I291331,I291507,);
not I_16998 (I291323,I291507);
nor I_16999 (I291529,I291357,I291464);
nor I_17000 (I291305,I291408,I291529);
DFFARX1 I_17001 (I843372,I2507,I291331,I291569,);
DFFARX1 I_17002 (I291569,I2507,I291331,I291586,);
not I_17003 (I291594,I291586);
not I_17004 (I291611,I291569);
nand I_17005 (I291308,I291611,I291430);
nand I_17006 (I291642,I843354,I843363);
and I_17007 (I291659,I291642,I843357);
DFFARX1 I_17008 (I291659,I2507,I291331,I291685,);
nor I_17009 (I291693,I291685,I291357);
DFFARX1 I_17010 (I291693,I2507,I291331,I291296,);
DFFARX1 I_17011 (I291685,I2507,I291331,I291314,);
nor I_17012 (I291738,I843375,I843363);
not I_17013 (I291755,I291738);
nor I_17014 (I291317,I291594,I291755);
nand I_17015 (I291302,I291611,I291755);
nor I_17016 (I291311,I291357,I291738);
DFFARX1 I_17017 (I291738,I2507,I291331,I291320,);
not I_17018 (I291858,I2514);
DFFARX1 I_17019 (I192475,I2507,I291858,I291884,);
nand I_17020 (I291892,I192475,I192481);
and I_17021 (I291909,I291892,I192499);
DFFARX1 I_17022 (I291909,I2507,I291858,I291935,);
nor I_17023 (I291826,I291935,I291884);
not I_17024 (I291957,I291935);
DFFARX1 I_17025 (I192487,I2507,I291858,I291983,);
nand I_17026 (I291991,I291983,I192484);
not I_17027 (I292008,I291991);
DFFARX1 I_17028 (I292008,I2507,I291858,I292034,);
not I_17029 (I291850,I292034);
nor I_17030 (I292056,I291884,I291991);
nor I_17031 (I291832,I291935,I292056);
DFFARX1 I_17032 (I192493,I2507,I291858,I292096,);
DFFARX1 I_17033 (I292096,I2507,I291858,I292113,);
not I_17034 (I292121,I292113);
not I_17035 (I292138,I292096);
nand I_17036 (I291835,I292138,I291957);
nand I_17037 (I292169,I192478,I192478);
and I_17038 (I292186,I292169,I192490);
DFFARX1 I_17039 (I292186,I2507,I291858,I292212,);
nor I_17040 (I292220,I292212,I291884);
DFFARX1 I_17041 (I292220,I2507,I291858,I291823,);
DFFARX1 I_17042 (I292212,I2507,I291858,I291841,);
nor I_17043 (I292265,I192496,I192478);
not I_17044 (I292282,I292265);
nor I_17045 (I291844,I292121,I292282);
nand I_17046 (I291829,I292138,I292282);
nor I_17047 (I291838,I291884,I292265);
DFFARX1 I_17048 (I292265,I2507,I291858,I291847,);
not I_17049 (I292385,I2514);
DFFARX1 I_17050 (I1116170,I2507,I292385,I292411,);
nand I_17051 (I292419,I1116185,I1116170);
and I_17052 (I292436,I292419,I1116188);
DFFARX1 I_17053 (I292436,I2507,I292385,I292462,);
nor I_17054 (I292353,I292462,I292411);
not I_17055 (I292484,I292462);
DFFARX1 I_17056 (I1116194,I2507,I292385,I292510,);
nand I_17057 (I292518,I292510,I1116176);
not I_17058 (I292535,I292518);
DFFARX1 I_17059 (I292535,I2507,I292385,I292561,);
not I_17060 (I292377,I292561);
nor I_17061 (I292583,I292411,I292518);
nor I_17062 (I292359,I292462,I292583);
DFFARX1 I_17063 (I1116173,I2507,I292385,I292623,);
DFFARX1 I_17064 (I292623,I2507,I292385,I292640,);
not I_17065 (I292648,I292640);
not I_17066 (I292665,I292623);
nand I_17067 (I292362,I292665,I292484);
nand I_17068 (I292696,I1116173,I1116179);
and I_17069 (I292713,I292696,I1116191);
DFFARX1 I_17070 (I292713,I2507,I292385,I292739,);
nor I_17071 (I292747,I292739,I292411);
DFFARX1 I_17072 (I292747,I2507,I292385,I292350,);
DFFARX1 I_17073 (I292739,I2507,I292385,I292368,);
nor I_17074 (I292792,I1116182,I1116179);
not I_17075 (I292809,I292792);
nor I_17076 (I292371,I292648,I292809);
nand I_17077 (I292356,I292665,I292809);
nor I_17078 (I292365,I292411,I292792);
DFFARX1 I_17079 (I292792,I2507,I292385,I292374,);
not I_17080 (I292912,I2514);
DFFARX1 I_17081 (I480059,I2507,I292912,I292938,);
nand I_17082 (I292946,I480071,I480050);
and I_17083 (I292963,I292946,I480074);
DFFARX1 I_17084 (I292963,I2507,I292912,I292989,);
nor I_17085 (I292880,I292989,I292938);
not I_17086 (I293011,I292989);
DFFARX1 I_17087 (I480065,I2507,I292912,I293037,);
nand I_17088 (I293045,I293037,I480047);
not I_17089 (I293062,I293045);
DFFARX1 I_17090 (I293062,I2507,I292912,I293088,);
not I_17091 (I292904,I293088);
nor I_17092 (I293110,I292938,I293045);
nor I_17093 (I292886,I292989,I293110);
DFFARX1 I_17094 (I480062,I2507,I292912,I293150,);
DFFARX1 I_17095 (I293150,I2507,I292912,I293167,);
not I_17096 (I293175,I293167);
not I_17097 (I293192,I293150);
nand I_17098 (I292889,I293192,I293011);
nand I_17099 (I293223,I480047,I480053);
and I_17100 (I293240,I293223,I480056);
DFFARX1 I_17101 (I293240,I2507,I292912,I293266,);
nor I_17102 (I293274,I293266,I292938);
DFFARX1 I_17103 (I293274,I2507,I292912,I292877,);
DFFARX1 I_17104 (I293266,I2507,I292912,I292895,);
nor I_17105 (I293319,I480068,I480053);
not I_17106 (I293336,I293319);
nor I_17107 (I292898,I293175,I293336);
nand I_17108 (I292883,I293192,I293336);
nor I_17109 (I292892,I292938,I293319);
DFFARX1 I_17110 (I293319,I2507,I292912,I292901,);
not I_17111 (I293439,I2514);
DFFARX1 I_17112 (I589117,I2507,I293439,I293465,);
nand I_17113 (I293473,I589102,I589105);
and I_17114 (I293490,I293473,I589120);
DFFARX1 I_17115 (I293490,I2507,I293439,I293516,);
nor I_17116 (I293407,I293516,I293465);
not I_17117 (I293538,I293516);
DFFARX1 I_17118 (I589114,I2507,I293439,I293564,);
nand I_17119 (I293572,I293564,I589105);
not I_17120 (I293589,I293572);
DFFARX1 I_17121 (I293589,I2507,I293439,I293615,);
not I_17122 (I293431,I293615);
nor I_17123 (I293637,I293465,I293572);
nor I_17124 (I293413,I293516,I293637);
DFFARX1 I_17125 (I589111,I2507,I293439,I293677,);
DFFARX1 I_17126 (I293677,I2507,I293439,I293694,);
not I_17127 (I293702,I293694);
not I_17128 (I293719,I293677);
nand I_17129 (I293416,I293719,I293538);
nand I_17130 (I293750,I589126,I589102);
and I_17131 (I293767,I293750,I589123);
DFFARX1 I_17132 (I293767,I2507,I293439,I293793,);
nor I_17133 (I293801,I293793,I293465);
DFFARX1 I_17134 (I293801,I2507,I293439,I293404,);
DFFARX1 I_17135 (I293793,I2507,I293439,I293422,);
nor I_17136 (I293846,I589108,I589102);
not I_17137 (I293863,I293846);
nor I_17138 (I293425,I293702,I293863);
nand I_17139 (I293410,I293719,I293863);
nor I_17140 (I293419,I293465,I293846);
DFFARX1 I_17141 (I293846,I2507,I293439,I293428,);
not I_17142 (I293966,I2514);
DFFARX1 I_17143 (I910184,I2507,I293966,I293992,);
nand I_17144 (I294000,I910181,I910199);
and I_17145 (I294017,I294000,I910190);
DFFARX1 I_17146 (I294017,I2507,I293966,I294043,);
nor I_17147 (I293934,I294043,I293992);
not I_17148 (I294065,I294043);
DFFARX1 I_17149 (I910205,I2507,I293966,I294091,);
nand I_17150 (I294099,I294091,I910187);
not I_17151 (I294116,I294099);
DFFARX1 I_17152 (I294116,I2507,I293966,I294142,);
not I_17153 (I293958,I294142);
nor I_17154 (I294164,I293992,I294099);
nor I_17155 (I293940,I294043,I294164);
DFFARX1 I_17156 (I910193,I2507,I293966,I294204,);
DFFARX1 I_17157 (I294204,I2507,I293966,I294221,);
not I_17158 (I294229,I294221);
not I_17159 (I294246,I294204);
nand I_17160 (I293943,I294246,I294065);
nand I_17161 (I294277,I910181,I910208);
and I_17162 (I294294,I294277,I910196);
DFFARX1 I_17163 (I294294,I2507,I293966,I294320,);
nor I_17164 (I294328,I294320,I293992);
DFFARX1 I_17165 (I294328,I2507,I293966,I293931,);
DFFARX1 I_17166 (I294320,I2507,I293966,I293949,);
nor I_17167 (I294373,I910202,I910208);
not I_17168 (I294390,I294373);
nor I_17169 (I293952,I294229,I294390);
nand I_17170 (I293937,I294246,I294390);
nor I_17171 (I293946,I293992,I294373);
DFFARX1 I_17172 (I294373,I2507,I293966,I293955,);
not I_17173 (I294493,I2514);
DFFARX1 I_17174 (I1217236,I2507,I294493,I294519,);
nand I_17175 (I294527,I1217218,I1217242);
and I_17176 (I294544,I294527,I1217233);
DFFARX1 I_17177 (I294544,I2507,I294493,I294570,);
nor I_17178 (I294461,I294570,I294519);
not I_17179 (I294592,I294570);
DFFARX1 I_17180 (I1217239,I2507,I294493,I294618,);
nand I_17181 (I294626,I294618,I1217227);
not I_17182 (I294643,I294626);
DFFARX1 I_17183 (I294643,I2507,I294493,I294669,);
not I_17184 (I294485,I294669);
nor I_17185 (I294691,I294519,I294626);
nor I_17186 (I294467,I294570,I294691);
DFFARX1 I_17187 (I1217218,I2507,I294493,I294731,);
DFFARX1 I_17188 (I294731,I2507,I294493,I294748,);
not I_17189 (I294756,I294748);
not I_17190 (I294773,I294731);
nand I_17191 (I294470,I294773,I294592);
nand I_17192 (I294804,I1217224,I1217221);
and I_17193 (I294821,I294804,I1217230);
DFFARX1 I_17194 (I294821,I2507,I294493,I294847,);
nor I_17195 (I294855,I294847,I294519);
DFFARX1 I_17196 (I294855,I2507,I294493,I294458,);
DFFARX1 I_17197 (I294847,I2507,I294493,I294476,);
nor I_17198 (I294900,I1217221,I1217221);
not I_17199 (I294917,I294900);
nor I_17200 (I294479,I294756,I294917);
nand I_17201 (I294464,I294773,I294917);
nor I_17202 (I294473,I294519,I294900);
DFFARX1 I_17203 (I294900,I2507,I294493,I294482,);
not I_17204 (I295020,I2514);
DFFARX1 I_17205 (I194260,I2507,I295020,I295046,);
nand I_17206 (I295054,I194260,I194266);
and I_17207 (I295071,I295054,I194284);
DFFARX1 I_17208 (I295071,I2507,I295020,I295097,);
nor I_17209 (I294988,I295097,I295046);
not I_17210 (I295119,I295097);
DFFARX1 I_17211 (I194272,I2507,I295020,I295145,);
nand I_17212 (I295153,I295145,I194269);
not I_17213 (I295170,I295153);
DFFARX1 I_17214 (I295170,I2507,I295020,I295196,);
not I_17215 (I295012,I295196);
nor I_17216 (I295218,I295046,I295153);
nor I_17217 (I294994,I295097,I295218);
DFFARX1 I_17218 (I194278,I2507,I295020,I295258,);
DFFARX1 I_17219 (I295258,I2507,I295020,I295275,);
not I_17220 (I295283,I295275);
not I_17221 (I295300,I295258);
nand I_17222 (I294997,I295300,I295119);
nand I_17223 (I295331,I194263,I194263);
and I_17224 (I295348,I295331,I194275);
DFFARX1 I_17225 (I295348,I2507,I295020,I295374,);
nor I_17226 (I295382,I295374,I295046);
DFFARX1 I_17227 (I295382,I2507,I295020,I294985,);
DFFARX1 I_17228 (I295374,I2507,I295020,I295003,);
nor I_17229 (I295427,I194281,I194263);
not I_17230 (I295444,I295427);
nor I_17231 (I295006,I295283,I295444);
nand I_17232 (I294991,I295300,I295444);
nor I_17233 (I295000,I295046,I295427);
DFFARX1 I_17234 (I295427,I2507,I295020,I295009,);
not I_17235 (I295547,I2514);
DFFARX1 I_17236 (I226390,I2507,I295547,I295573,);
nand I_17237 (I295581,I226390,I226396);
and I_17238 (I295598,I295581,I226414);
DFFARX1 I_17239 (I295598,I2507,I295547,I295624,);
nor I_17240 (I295515,I295624,I295573);
not I_17241 (I295646,I295624);
DFFARX1 I_17242 (I226402,I2507,I295547,I295672,);
nand I_17243 (I295680,I295672,I226399);
not I_17244 (I295697,I295680);
DFFARX1 I_17245 (I295697,I2507,I295547,I295723,);
not I_17246 (I295539,I295723);
nor I_17247 (I295745,I295573,I295680);
nor I_17248 (I295521,I295624,I295745);
DFFARX1 I_17249 (I226408,I2507,I295547,I295785,);
DFFARX1 I_17250 (I295785,I2507,I295547,I295802,);
not I_17251 (I295810,I295802);
not I_17252 (I295827,I295785);
nand I_17253 (I295524,I295827,I295646);
nand I_17254 (I295858,I226393,I226393);
and I_17255 (I295875,I295858,I226405);
DFFARX1 I_17256 (I295875,I2507,I295547,I295901,);
nor I_17257 (I295909,I295901,I295573);
DFFARX1 I_17258 (I295909,I2507,I295547,I295512,);
DFFARX1 I_17259 (I295901,I2507,I295547,I295530,);
nor I_17260 (I295954,I226411,I226393);
not I_17261 (I295971,I295954);
nor I_17262 (I295533,I295810,I295971);
nand I_17263 (I295518,I295827,I295971);
nor I_17264 (I295527,I295573,I295954);
DFFARX1 I_17265 (I295954,I2507,I295547,I295536,);
not I_17266 (I296074,I2514);
DFFARX1 I_17267 (I713962,I2507,I296074,I296100,);
nand I_17268 (I296108,I713953,I713968);
and I_17269 (I296125,I296108,I713974);
DFFARX1 I_17270 (I296125,I2507,I296074,I296151,);
nor I_17271 (I296042,I296151,I296100);
not I_17272 (I296173,I296151);
DFFARX1 I_17273 (I713959,I2507,I296074,I296199,);
nand I_17274 (I296207,I296199,I713953);
not I_17275 (I296224,I296207);
DFFARX1 I_17276 (I296224,I2507,I296074,I296250,);
not I_17277 (I296066,I296250);
nor I_17278 (I296272,I296100,I296207);
nor I_17279 (I296048,I296151,I296272);
DFFARX1 I_17280 (I713956,I2507,I296074,I296312,);
DFFARX1 I_17281 (I296312,I2507,I296074,I296329,);
not I_17282 (I296337,I296329);
not I_17283 (I296354,I296312);
nand I_17284 (I296051,I296354,I296173);
nand I_17285 (I296385,I713950,I713965);
and I_17286 (I296402,I296385,I713950);
DFFARX1 I_17287 (I296402,I2507,I296074,I296428,);
nor I_17288 (I296436,I296428,I296100);
DFFARX1 I_17289 (I296436,I2507,I296074,I296039,);
DFFARX1 I_17290 (I296428,I2507,I296074,I296057,);
nor I_17291 (I296481,I713971,I713965);
not I_17292 (I296498,I296481);
nor I_17293 (I296060,I296337,I296498);
nand I_17294 (I296045,I296354,I296498);
nor I_17295 (I296054,I296100,I296481);
DFFARX1 I_17296 (I296481,I2507,I296074,I296063,);
not I_17297 (I296601,I2514);
DFFARX1 I_17298 (I1392798,I2507,I296601,I296627,);
nand I_17299 (I296635,I1392777,I1392777);
and I_17300 (I296652,I296635,I1392804);
DFFARX1 I_17301 (I296652,I2507,I296601,I296678,);
nor I_17302 (I296569,I296678,I296627);
not I_17303 (I296700,I296678);
DFFARX1 I_17304 (I1392792,I2507,I296601,I296726,);
nand I_17305 (I296734,I296726,I1392795);
not I_17306 (I296751,I296734);
DFFARX1 I_17307 (I296751,I2507,I296601,I296777,);
not I_17308 (I296593,I296777);
nor I_17309 (I296799,I296627,I296734);
nor I_17310 (I296575,I296678,I296799);
DFFARX1 I_17311 (I1392786,I2507,I296601,I296839,);
DFFARX1 I_17312 (I296839,I2507,I296601,I296856,);
not I_17313 (I296864,I296856);
not I_17314 (I296881,I296839);
nand I_17315 (I296578,I296881,I296700);
nand I_17316 (I296912,I1392783,I1392780);
and I_17317 (I296929,I296912,I1392801);
DFFARX1 I_17318 (I296929,I2507,I296601,I296955,);
nor I_17319 (I296963,I296955,I296627);
DFFARX1 I_17320 (I296963,I2507,I296601,I296566,);
DFFARX1 I_17321 (I296955,I2507,I296601,I296584,);
nor I_17322 (I297008,I1392789,I1392780);
not I_17323 (I297025,I297008);
nor I_17324 (I296587,I296864,I297025);
nand I_17325 (I296572,I296881,I297025);
nor I_17326 (I296581,I296627,I297008);
DFFARX1 I_17327 (I297008,I2507,I296601,I296590,);
not I_17328 (I297128,I2514);
DFFARX1 I_17329 (I905016,I2507,I297128,I297154,);
nand I_17330 (I297162,I905013,I905031);
and I_17331 (I297179,I297162,I905022);
DFFARX1 I_17332 (I297179,I2507,I297128,I297205,);
nor I_17333 (I297096,I297205,I297154);
not I_17334 (I297227,I297205);
DFFARX1 I_17335 (I905037,I2507,I297128,I297253,);
nand I_17336 (I297261,I297253,I905019);
not I_17337 (I297278,I297261);
DFFARX1 I_17338 (I297278,I2507,I297128,I297304,);
not I_17339 (I297120,I297304);
nor I_17340 (I297326,I297154,I297261);
nor I_17341 (I297102,I297205,I297326);
DFFARX1 I_17342 (I905025,I2507,I297128,I297366,);
DFFARX1 I_17343 (I297366,I2507,I297128,I297383,);
not I_17344 (I297391,I297383);
not I_17345 (I297408,I297366);
nand I_17346 (I297105,I297408,I297227);
nand I_17347 (I297439,I905013,I905040);
and I_17348 (I297456,I297439,I905028);
DFFARX1 I_17349 (I297456,I2507,I297128,I297482,);
nor I_17350 (I297490,I297482,I297154);
DFFARX1 I_17351 (I297490,I2507,I297128,I297093,);
DFFARX1 I_17352 (I297482,I2507,I297128,I297111,);
nor I_17353 (I297535,I905034,I905040);
not I_17354 (I297552,I297535);
nor I_17355 (I297114,I297391,I297552);
nand I_17356 (I297099,I297408,I297552);
nor I_17357 (I297108,I297154,I297535);
DFFARX1 I_17358 (I297535,I2507,I297128,I297117,);
not I_17359 (I297655,I2514);
DFFARX1 I_17360 (I388667,I2507,I297655,I297681,);
nand I_17361 (I297689,I388679,I388658);
and I_17362 (I297706,I297689,I388682);
DFFARX1 I_17363 (I297706,I2507,I297655,I297732,);
nor I_17364 (I297623,I297732,I297681);
not I_17365 (I297754,I297732);
DFFARX1 I_17366 (I388673,I2507,I297655,I297780,);
nand I_17367 (I297788,I297780,I388655);
not I_17368 (I297805,I297788);
DFFARX1 I_17369 (I297805,I2507,I297655,I297831,);
not I_17370 (I297647,I297831);
nor I_17371 (I297853,I297681,I297788);
nor I_17372 (I297629,I297732,I297853);
DFFARX1 I_17373 (I388670,I2507,I297655,I297893,);
DFFARX1 I_17374 (I297893,I2507,I297655,I297910,);
not I_17375 (I297918,I297910);
not I_17376 (I297935,I297893);
nand I_17377 (I297632,I297935,I297754);
nand I_17378 (I297966,I388655,I388661);
and I_17379 (I297983,I297966,I388664);
DFFARX1 I_17380 (I297983,I2507,I297655,I298009,);
nor I_17381 (I298017,I298009,I297681);
DFFARX1 I_17382 (I298017,I2507,I297655,I297620,);
DFFARX1 I_17383 (I298009,I2507,I297655,I297638,);
nor I_17384 (I298062,I388676,I388661);
not I_17385 (I298079,I298062);
nor I_17386 (I297641,I297918,I298079);
nand I_17387 (I297626,I297935,I298079);
nor I_17388 (I297635,I297681,I298062);
DFFARX1 I_17389 (I298062,I2507,I297655,I297644,);
not I_17390 (I298182,I2514);
DFFARX1 I_17391 (I611081,I2507,I298182,I298208,);
nand I_17392 (I298216,I611066,I611069);
and I_17393 (I298233,I298216,I611084);
DFFARX1 I_17394 (I298233,I2507,I298182,I298259,);
nor I_17395 (I298150,I298259,I298208);
not I_17396 (I298281,I298259);
DFFARX1 I_17397 (I611078,I2507,I298182,I298307,);
nand I_17398 (I298315,I298307,I611069);
not I_17399 (I298332,I298315);
DFFARX1 I_17400 (I298332,I2507,I298182,I298358,);
not I_17401 (I298174,I298358);
nor I_17402 (I298380,I298208,I298315);
nor I_17403 (I298156,I298259,I298380);
DFFARX1 I_17404 (I611075,I2507,I298182,I298420,);
DFFARX1 I_17405 (I298420,I2507,I298182,I298437,);
not I_17406 (I298445,I298437);
not I_17407 (I298462,I298420);
nand I_17408 (I298159,I298462,I298281);
nand I_17409 (I298493,I611090,I611066);
and I_17410 (I298510,I298493,I611087);
DFFARX1 I_17411 (I298510,I2507,I298182,I298536,);
nor I_17412 (I298544,I298536,I298208);
DFFARX1 I_17413 (I298544,I2507,I298182,I298147,);
DFFARX1 I_17414 (I298536,I2507,I298182,I298165,);
nor I_17415 (I298589,I611072,I611066);
not I_17416 (I298606,I298589);
nor I_17417 (I298168,I298445,I298606);
nand I_17418 (I298153,I298462,I298606);
nor I_17419 (I298162,I298208,I298589);
DFFARX1 I_17420 (I298589,I2507,I298182,I298171,);
not I_17421 (I298709,I2514);
DFFARX1 I_17422 (I576401,I2507,I298709,I298735,);
nand I_17423 (I298743,I576386,I576389);
and I_17424 (I298760,I298743,I576404);
DFFARX1 I_17425 (I298760,I2507,I298709,I298786,);
nor I_17426 (I298677,I298786,I298735);
not I_17427 (I298808,I298786);
DFFARX1 I_17428 (I576398,I2507,I298709,I298834,);
nand I_17429 (I298842,I298834,I576389);
not I_17430 (I298859,I298842);
DFFARX1 I_17431 (I298859,I2507,I298709,I298885,);
not I_17432 (I298701,I298885);
nor I_17433 (I298907,I298735,I298842);
nor I_17434 (I298683,I298786,I298907);
DFFARX1 I_17435 (I576395,I2507,I298709,I298947,);
DFFARX1 I_17436 (I298947,I2507,I298709,I298964,);
not I_17437 (I298972,I298964);
not I_17438 (I298989,I298947);
nand I_17439 (I298686,I298989,I298808);
nand I_17440 (I299020,I576410,I576386);
and I_17441 (I299037,I299020,I576407);
DFFARX1 I_17442 (I299037,I2507,I298709,I299063,);
nor I_17443 (I299071,I299063,I298735);
DFFARX1 I_17444 (I299071,I2507,I298709,I298674,);
DFFARX1 I_17445 (I299063,I2507,I298709,I298692,);
nor I_17446 (I299116,I576392,I576386);
not I_17447 (I299133,I299116);
nor I_17448 (I298695,I298972,I299133);
nand I_17449 (I298680,I298989,I299133);
nor I_17450 (I298689,I298735,I299116);
DFFARX1 I_17451 (I299116,I2507,I298709,I298698,);
not I_17452 (I299236,I2514);
DFFARX1 I_17453 (I474619,I2507,I299236,I299262,);
nand I_17454 (I299270,I474631,I474610);
and I_17455 (I299287,I299270,I474634);
DFFARX1 I_17456 (I299287,I2507,I299236,I299313,);
nor I_17457 (I299204,I299313,I299262);
not I_17458 (I299335,I299313);
DFFARX1 I_17459 (I474625,I2507,I299236,I299361,);
nand I_17460 (I299369,I299361,I474607);
not I_17461 (I299386,I299369);
DFFARX1 I_17462 (I299386,I2507,I299236,I299412,);
not I_17463 (I299228,I299412);
nor I_17464 (I299434,I299262,I299369);
nor I_17465 (I299210,I299313,I299434);
DFFARX1 I_17466 (I474622,I2507,I299236,I299474,);
DFFARX1 I_17467 (I299474,I2507,I299236,I299491,);
not I_17468 (I299499,I299491);
not I_17469 (I299516,I299474);
nand I_17470 (I299213,I299516,I299335);
nand I_17471 (I299547,I474607,I474613);
and I_17472 (I299564,I299547,I474616);
DFFARX1 I_17473 (I299564,I2507,I299236,I299590,);
nor I_17474 (I299598,I299590,I299262);
DFFARX1 I_17475 (I299598,I2507,I299236,I299201,);
DFFARX1 I_17476 (I299590,I2507,I299236,I299219,);
nor I_17477 (I299643,I474628,I474613);
not I_17478 (I299660,I299643);
nor I_17479 (I299222,I299499,I299660);
nand I_17480 (I299207,I299516,I299660);
nor I_17481 (I299216,I299262,I299643);
DFFARX1 I_17482 (I299643,I2507,I299236,I299225,);
not I_17483 (I299763,I2514);
DFFARX1 I_17484 (I731880,I2507,I299763,I299789,);
nand I_17485 (I299797,I731871,I731886);
and I_17486 (I299814,I299797,I731892);
DFFARX1 I_17487 (I299814,I2507,I299763,I299840,);
nor I_17488 (I299731,I299840,I299789);
not I_17489 (I299862,I299840);
DFFARX1 I_17490 (I731877,I2507,I299763,I299888,);
nand I_17491 (I299896,I299888,I731871);
not I_17492 (I299913,I299896);
DFFARX1 I_17493 (I299913,I2507,I299763,I299939,);
not I_17494 (I299755,I299939);
nor I_17495 (I299961,I299789,I299896);
nor I_17496 (I299737,I299840,I299961);
DFFARX1 I_17497 (I731874,I2507,I299763,I300001,);
DFFARX1 I_17498 (I300001,I2507,I299763,I300018,);
not I_17499 (I300026,I300018);
not I_17500 (I300043,I300001);
nand I_17501 (I299740,I300043,I299862);
nand I_17502 (I300074,I731868,I731883);
and I_17503 (I300091,I300074,I731868);
DFFARX1 I_17504 (I300091,I2507,I299763,I300117,);
nor I_17505 (I300125,I300117,I299789);
DFFARX1 I_17506 (I300125,I2507,I299763,I299728,);
DFFARX1 I_17507 (I300117,I2507,I299763,I299746,);
nor I_17508 (I300170,I731889,I731883);
not I_17509 (I300187,I300170);
nor I_17510 (I299749,I300026,I300187);
nand I_17511 (I299734,I300043,I300187);
nor I_17512 (I299743,I299789,I300170);
DFFARX1 I_17513 (I300170,I2507,I299763,I299752,);
not I_17514 (I300290,I2514);
DFFARX1 I_17515 (I990934,I2507,I300290,I300316,);
nand I_17516 (I300324,I990931,I990949);
and I_17517 (I300341,I300324,I990940);
DFFARX1 I_17518 (I300341,I2507,I300290,I300367,);
nor I_17519 (I300258,I300367,I300316);
not I_17520 (I300389,I300367);
DFFARX1 I_17521 (I990955,I2507,I300290,I300415,);
nand I_17522 (I300423,I300415,I990937);
not I_17523 (I300440,I300423);
DFFARX1 I_17524 (I300440,I2507,I300290,I300466,);
not I_17525 (I300282,I300466);
nor I_17526 (I300488,I300316,I300423);
nor I_17527 (I300264,I300367,I300488);
DFFARX1 I_17528 (I990943,I2507,I300290,I300528,);
DFFARX1 I_17529 (I300528,I2507,I300290,I300545,);
not I_17530 (I300553,I300545);
not I_17531 (I300570,I300528);
nand I_17532 (I300267,I300570,I300389);
nand I_17533 (I300601,I990931,I990958);
and I_17534 (I300618,I300601,I990946);
DFFARX1 I_17535 (I300618,I2507,I300290,I300644,);
nor I_17536 (I300652,I300644,I300316);
DFFARX1 I_17537 (I300652,I2507,I300290,I300255,);
DFFARX1 I_17538 (I300644,I2507,I300290,I300273,);
nor I_17539 (I300697,I990952,I990958);
not I_17540 (I300714,I300697);
nor I_17541 (I300276,I300553,I300714);
nand I_17542 (I300261,I300570,I300714);
nor I_17543 (I300270,I300316,I300697);
DFFARX1 I_17544 (I300697,I2507,I300290,I300279,);
not I_17545 (I300817,I2514);
DFFARX1 I_17546 (I394651,I2507,I300817,I300843,);
nand I_17547 (I300851,I394663,I394642);
and I_17548 (I300868,I300851,I394666);
DFFARX1 I_17549 (I300868,I2507,I300817,I300894,);
nor I_17550 (I300785,I300894,I300843);
not I_17551 (I300916,I300894);
DFFARX1 I_17552 (I394657,I2507,I300817,I300942,);
nand I_17553 (I300950,I300942,I394639);
not I_17554 (I300967,I300950);
DFFARX1 I_17555 (I300967,I2507,I300817,I300993,);
not I_17556 (I300809,I300993);
nor I_17557 (I301015,I300843,I300950);
nor I_17558 (I300791,I300894,I301015);
DFFARX1 I_17559 (I394654,I2507,I300817,I301055,);
DFFARX1 I_17560 (I301055,I2507,I300817,I301072,);
not I_17561 (I301080,I301072);
not I_17562 (I301097,I301055);
nand I_17563 (I300794,I301097,I300916);
nand I_17564 (I301128,I394639,I394645);
and I_17565 (I301145,I301128,I394648);
DFFARX1 I_17566 (I301145,I2507,I300817,I301171,);
nor I_17567 (I301179,I301171,I300843);
DFFARX1 I_17568 (I301179,I2507,I300817,I300782,);
DFFARX1 I_17569 (I301171,I2507,I300817,I300800,);
nor I_17570 (I301224,I394660,I394645);
not I_17571 (I301241,I301224);
nor I_17572 (I300803,I301080,I301241);
nand I_17573 (I300788,I301097,I301241);
nor I_17574 (I300797,I300843,I301224);
DFFARX1 I_17575 (I301224,I2507,I300817,I300806,);
not I_17576 (I301344,I2514);
DFFARX1 I_17577 (I638244,I2507,I301344,I301370,);
nand I_17578 (I301378,I638235,I638250);
and I_17579 (I301395,I301378,I638256);
DFFARX1 I_17580 (I301395,I2507,I301344,I301421,);
nor I_17581 (I301312,I301421,I301370);
not I_17582 (I301443,I301421);
DFFARX1 I_17583 (I638241,I2507,I301344,I301469,);
nand I_17584 (I301477,I301469,I638235);
not I_17585 (I301494,I301477);
DFFARX1 I_17586 (I301494,I2507,I301344,I301520,);
not I_17587 (I301336,I301520);
nor I_17588 (I301542,I301370,I301477);
nor I_17589 (I301318,I301421,I301542);
DFFARX1 I_17590 (I638238,I2507,I301344,I301582,);
DFFARX1 I_17591 (I301582,I2507,I301344,I301599,);
not I_17592 (I301607,I301599);
not I_17593 (I301624,I301582);
nand I_17594 (I301321,I301624,I301443);
nand I_17595 (I301655,I638232,I638247);
and I_17596 (I301672,I301655,I638232);
DFFARX1 I_17597 (I301672,I2507,I301344,I301698,);
nor I_17598 (I301706,I301698,I301370);
DFFARX1 I_17599 (I301706,I2507,I301344,I301309,);
DFFARX1 I_17600 (I301698,I2507,I301344,I301327,);
nor I_17601 (I301751,I638253,I638247);
not I_17602 (I301768,I301751);
nor I_17603 (I301330,I301607,I301768);
nand I_17604 (I301315,I301624,I301768);
nor I_17605 (I301324,I301370,I301751);
DFFARX1 I_17606 (I301751,I2507,I301344,I301333,);
not I_17607 (I301871,I2514);
DFFARX1 I_17608 (I814372,I2507,I301871,I301897,);
nand I_17609 (I301905,I814375,I814369);
and I_17610 (I301922,I301905,I814381);
DFFARX1 I_17611 (I301922,I2507,I301871,I301948,);
nor I_17612 (I301839,I301948,I301897);
not I_17613 (I301970,I301948);
DFFARX1 I_17614 (I814384,I2507,I301871,I301996,);
nand I_17615 (I302004,I301996,I814375);
not I_17616 (I302021,I302004);
DFFARX1 I_17617 (I302021,I2507,I301871,I302047,);
not I_17618 (I301863,I302047);
nor I_17619 (I302069,I301897,I302004);
nor I_17620 (I301845,I301948,I302069);
DFFARX1 I_17621 (I814387,I2507,I301871,I302109,);
DFFARX1 I_17622 (I302109,I2507,I301871,I302126,);
not I_17623 (I302134,I302126);
not I_17624 (I302151,I302109);
nand I_17625 (I301848,I302151,I301970);
nand I_17626 (I302182,I814369,I814378);
and I_17627 (I302199,I302182,I814372);
DFFARX1 I_17628 (I302199,I2507,I301871,I302225,);
nor I_17629 (I302233,I302225,I301897);
DFFARX1 I_17630 (I302233,I2507,I301871,I301836,);
DFFARX1 I_17631 (I302225,I2507,I301871,I301854,);
nor I_17632 (I302278,I814390,I814378);
not I_17633 (I302295,I302278);
nor I_17634 (I301857,I302134,I302295);
nand I_17635 (I301842,I302151,I302295);
nor I_17636 (I301851,I301897,I302278);
DFFARX1 I_17637 (I302278,I2507,I301871,I301860,);
not I_17638 (I302398,I2514);
DFFARX1 I_17639 (I978660,I2507,I302398,I302424,);
nand I_17640 (I302432,I978657,I978675);
and I_17641 (I302449,I302432,I978666);
DFFARX1 I_17642 (I302449,I2507,I302398,I302475,);
nor I_17643 (I302366,I302475,I302424);
not I_17644 (I302497,I302475);
DFFARX1 I_17645 (I978681,I2507,I302398,I302523,);
nand I_17646 (I302531,I302523,I978663);
not I_17647 (I302548,I302531);
DFFARX1 I_17648 (I302548,I2507,I302398,I302574,);
not I_17649 (I302390,I302574);
nor I_17650 (I302596,I302424,I302531);
nor I_17651 (I302372,I302475,I302596);
DFFARX1 I_17652 (I978669,I2507,I302398,I302636,);
DFFARX1 I_17653 (I302636,I2507,I302398,I302653,);
not I_17654 (I302661,I302653);
not I_17655 (I302678,I302636);
nand I_17656 (I302375,I302678,I302497);
nand I_17657 (I302709,I978657,I978684);
and I_17658 (I302726,I302709,I978672);
DFFARX1 I_17659 (I302726,I2507,I302398,I302752,);
nor I_17660 (I302760,I302752,I302424);
DFFARX1 I_17661 (I302760,I2507,I302398,I302363,);
DFFARX1 I_17662 (I302752,I2507,I302398,I302381,);
nor I_17663 (I302805,I978678,I978684);
not I_17664 (I302822,I302805);
nor I_17665 (I302384,I302661,I302822);
nand I_17666 (I302369,I302678,I302822);
nor I_17667 (I302378,I302424,I302805);
DFFARX1 I_17668 (I302805,I2507,I302398,I302387,);
not I_17669 (I302925,I2514);
DFFARX1 I_17670 (I98077,I2507,I302925,I302951,);
nand I_17671 (I302959,I98089,I98098);
and I_17672 (I302976,I302959,I98077);
DFFARX1 I_17673 (I302976,I2507,I302925,I303002,);
nor I_17674 (I302893,I303002,I302951);
not I_17675 (I303024,I303002);
DFFARX1 I_17676 (I98092,I2507,I302925,I303050,);
nand I_17677 (I303058,I303050,I98080);
not I_17678 (I303075,I303058);
DFFARX1 I_17679 (I303075,I2507,I302925,I303101,);
not I_17680 (I302917,I303101);
nor I_17681 (I303123,I302951,I303058);
nor I_17682 (I302899,I303002,I303123);
DFFARX1 I_17683 (I98083,I2507,I302925,I303163,);
DFFARX1 I_17684 (I303163,I2507,I302925,I303180,);
not I_17685 (I303188,I303180);
not I_17686 (I303205,I303163);
nand I_17687 (I302902,I303205,I303024);
nand I_17688 (I303236,I98074,I98074);
and I_17689 (I303253,I303236,I98086);
DFFARX1 I_17690 (I303253,I2507,I302925,I303279,);
nor I_17691 (I303287,I303279,I302951);
DFFARX1 I_17692 (I303287,I2507,I302925,I302890,);
DFFARX1 I_17693 (I303279,I2507,I302925,I302908,);
nor I_17694 (I303332,I98095,I98074);
not I_17695 (I303349,I303332);
nor I_17696 (I302911,I303188,I303349);
nand I_17697 (I302896,I303205,I303349);
nor I_17698 (I302905,I302951,I303332);
DFFARX1 I_17699 (I303332,I2507,I302925,I302914,);
not I_17700 (I303452,I2514);
DFFARX1 I_17701 (I411515,I2507,I303452,I303478,);
nand I_17702 (I303486,I411527,I411506);
and I_17703 (I303503,I303486,I411530);
DFFARX1 I_17704 (I303503,I2507,I303452,I303529,);
nor I_17705 (I303420,I303529,I303478);
not I_17706 (I303551,I303529);
DFFARX1 I_17707 (I411521,I2507,I303452,I303577,);
nand I_17708 (I303585,I303577,I411503);
not I_17709 (I303602,I303585);
DFFARX1 I_17710 (I303602,I2507,I303452,I303628,);
not I_17711 (I303444,I303628);
nor I_17712 (I303650,I303478,I303585);
nor I_17713 (I303426,I303529,I303650);
DFFARX1 I_17714 (I411518,I2507,I303452,I303690,);
DFFARX1 I_17715 (I303690,I2507,I303452,I303707,);
not I_17716 (I303715,I303707);
not I_17717 (I303732,I303690);
nand I_17718 (I303429,I303732,I303551);
nand I_17719 (I303763,I411503,I411509);
and I_17720 (I303780,I303763,I411512);
DFFARX1 I_17721 (I303780,I2507,I303452,I303806,);
nor I_17722 (I303814,I303806,I303478);
DFFARX1 I_17723 (I303814,I2507,I303452,I303417,);
DFFARX1 I_17724 (I303806,I2507,I303452,I303435,);
nor I_17725 (I303859,I411524,I411509);
not I_17726 (I303876,I303859);
nor I_17727 (I303438,I303715,I303876);
nand I_17728 (I303423,I303732,I303876);
nor I_17729 (I303432,I303478,I303859);
DFFARX1 I_17730 (I303859,I2507,I303452,I303441,);
not I_17731 (I303979,I2514);
DFFARX1 I_17732 (I863910,I2507,I303979,I304005,);
nand I_17733 (I304013,I863913,I863907);
and I_17734 (I304030,I304013,I863919);
DFFARX1 I_17735 (I304030,I2507,I303979,I304056,);
nor I_17736 (I303947,I304056,I304005);
not I_17737 (I304078,I304056);
DFFARX1 I_17738 (I863922,I2507,I303979,I304104,);
nand I_17739 (I304112,I304104,I863913);
not I_17740 (I304129,I304112);
DFFARX1 I_17741 (I304129,I2507,I303979,I304155,);
not I_17742 (I303971,I304155);
nor I_17743 (I304177,I304005,I304112);
nor I_17744 (I303953,I304056,I304177);
DFFARX1 I_17745 (I863925,I2507,I303979,I304217,);
DFFARX1 I_17746 (I304217,I2507,I303979,I304234,);
not I_17747 (I304242,I304234);
not I_17748 (I304259,I304217);
nand I_17749 (I303956,I304259,I304078);
nand I_17750 (I304290,I863907,I863916);
and I_17751 (I304307,I304290,I863910);
DFFARX1 I_17752 (I304307,I2507,I303979,I304333,);
nor I_17753 (I304341,I304333,I304005);
DFFARX1 I_17754 (I304341,I2507,I303979,I303944,);
DFFARX1 I_17755 (I304333,I2507,I303979,I303962,);
nor I_17756 (I304386,I863928,I863916);
not I_17757 (I304403,I304386);
nor I_17758 (I303965,I304242,I304403);
nand I_17759 (I303950,I304259,I304403);
nor I_17760 (I303959,I304005,I304386);
DFFARX1 I_17761 (I304386,I2507,I303979,I303968,);
not I_17762 (I304506,I2514);
DFFARX1 I_17763 (I178790,I2507,I304506,I304532,);
nand I_17764 (I304540,I178790,I178796);
and I_17765 (I304557,I304540,I178814);
DFFARX1 I_17766 (I304557,I2507,I304506,I304583,);
nor I_17767 (I304474,I304583,I304532);
not I_17768 (I304605,I304583);
DFFARX1 I_17769 (I178802,I2507,I304506,I304631,);
nand I_17770 (I304639,I304631,I178799);
not I_17771 (I304656,I304639);
DFFARX1 I_17772 (I304656,I2507,I304506,I304682,);
not I_17773 (I304498,I304682);
nor I_17774 (I304704,I304532,I304639);
nor I_17775 (I304480,I304583,I304704);
DFFARX1 I_17776 (I178808,I2507,I304506,I304744,);
DFFARX1 I_17777 (I304744,I2507,I304506,I304761,);
not I_17778 (I304769,I304761);
not I_17779 (I304786,I304744);
nand I_17780 (I304483,I304786,I304605);
nand I_17781 (I304817,I178793,I178793);
and I_17782 (I304834,I304817,I178805);
DFFARX1 I_17783 (I304834,I2507,I304506,I304860,);
nor I_17784 (I304868,I304860,I304532);
DFFARX1 I_17785 (I304868,I2507,I304506,I304471,);
DFFARX1 I_17786 (I304860,I2507,I304506,I304489,);
nor I_17787 (I304913,I178811,I178793);
not I_17788 (I304930,I304913);
nor I_17789 (I304492,I304769,I304930);
nand I_17790 (I304477,I304786,I304930);
nor I_17791 (I304486,I304532,I304913);
DFFARX1 I_17792 (I304913,I2507,I304506,I304495,);
not I_17793 (I305033,I2514);
DFFARX1 I_17794 (I495877,I2507,I305033,I305059,);
nand I_17795 (I305067,I495877,I495889);
and I_17796 (I305084,I305067,I495874);
DFFARX1 I_17797 (I305084,I2507,I305033,I305110,);
nor I_17798 (I305001,I305110,I305059);
not I_17799 (I305132,I305110);
DFFARX1 I_17800 (I495898,I2507,I305033,I305158,);
nand I_17801 (I305166,I305158,I495895);
not I_17802 (I305183,I305166);
DFFARX1 I_17803 (I305183,I2507,I305033,I305209,);
not I_17804 (I305025,I305209);
nor I_17805 (I305231,I305059,I305166);
nor I_17806 (I305007,I305110,I305231);
DFFARX1 I_17807 (I495886,I2507,I305033,I305271,);
DFFARX1 I_17808 (I305271,I2507,I305033,I305288,);
not I_17809 (I305296,I305288);
not I_17810 (I305313,I305271);
nand I_17811 (I305010,I305313,I305132);
nand I_17812 (I305344,I495874,I495883);
and I_17813 (I305361,I305344,I495892);
DFFARX1 I_17814 (I305361,I2507,I305033,I305387,);
nor I_17815 (I305395,I305387,I305059);
DFFARX1 I_17816 (I305395,I2507,I305033,I304998,);
DFFARX1 I_17817 (I305387,I2507,I305033,I305016,);
nor I_17818 (I305440,I495880,I495883);
not I_17819 (I305457,I305440);
nor I_17820 (I305019,I305296,I305457);
nand I_17821 (I305004,I305313,I305457);
nor I_17822 (I305013,I305059,I305440);
DFFARX1 I_17823 (I305440,I2507,I305033,I305022,);
not I_17824 (I305560,I2514);
DFFARX1 I_17825 (I127062,I2507,I305560,I305586,);
nand I_17826 (I305594,I127074,I127083);
and I_17827 (I305611,I305594,I127062);
DFFARX1 I_17828 (I305611,I2507,I305560,I305637,);
nor I_17829 (I305528,I305637,I305586);
not I_17830 (I305659,I305637);
DFFARX1 I_17831 (I127077,I2507,I305560,I305685,);
nand I_17832 (I305693,I305685,I127065);
not I_17833 (I305710,I305693);
DFFARX1 I_17834 (I305710,I2507,I305560,I305736,);
not I_17835 (I305552,I305736);
nor I_17836 (I305758,I305586,I305693);
nor I_17837 (I305534,I305637,I305758);
DFFARX1 I_17838 (I127068,I2507,I305560,I305798,);
DFFARX1 I_17839 (I305798,I2507,I305560,I305815,);
not I_17840 (I305823,I305815);
not I_17841 (I305840,I305798);
nand I_17842 (I305537,I305840,I305659);
nand I_17843 (I305871,I127059,I127059);
and I_17844 (I305888,I305871,I127071);
DFFARX1 I_17845 (I305888,I2507,I305560,I305914,);
nor I_17846 (I305922,I305914,I305586);
DFFARX1 I_17847 (I305922,I2507,I305560,I305525,);
DFFARX1 I_17848 (I305914,I2507,I305560,I305543,);
nor I_17849 (I305967,I127080,I127059);
not I_17850 (I305984,I305967);
nor I_17851 (I305546,I305823,I305984);
nand I_17852 (I305531,I305840,I305984);
nor I_17853 (I305540,I305586,I305967);
DFFARX1 I_17854 (I305967,I2507,I305560,I305549,);
not I_17855 (I306087,I2514);
DFFARX1 I_17856 (I664254,I2507,I306087,I306113,);
nand I_17857 (I306121,I664245,I664260);
and I_17858 (I306138,I306121,I664266);
DFFARX1 I_17859 (I306138,I2507,I306087,I306164,);
nor I_17860 (I306055,I306164,I306113);
not I_17861 (I306186,I306164);
DFFARX1 I_17862 (I664251,I2507,I306087,I306212,);
nand I_17863 (I306220,I306212,I664245);
not I_17864 (I306237,I306220);
DFFARX1 I_17865 (I306237,I2507,I306087,I306263,);
not I_17866 (I306079,I306263);
nor I_17867 (I306285,I306113,I306220);
nor I_17868 (I306061,I306164,I306285);
DFFARX1 I_17869 (I664248,I2507,I306087,I306325,);
DFFARX1 I_17870 (I306325,I2507,I306087,I306342,);
not I_17871 (I306350,I306342);
not I_17872 (I306367,I306325);
nand I_17873 (I306064,I306367,I306186);
nand I_17874 (I306398,I664242,I664257);
and I_17875 (I306415,I306398,I664242);
DFFARX1 I_17876 (I306415,I2507,I306087,I306441,);
nor I_17877 (I306449,I306441,I306113);
DFFARX1 I_17878 (I306449,I2507,I306087,I306052,);
DFFARX1 I_17879 (I306441,I2507,I306087,I306070,);
nor I_17880 (I306494,I664263,I664257);
not I_17881 (I306511,I306494);
nor I_17882 (I306073,I306350,I306511);
nand I_17883 (I306058,I306367,I306511);
nor I_17884 (I306067,I306113,I306494);
DFFARX1 I_17885 (I306494,I2507,I306087,I306076,);
not I_17886 (I306614,I2514);
DFFARX1 I_17887 (I873923,I2507,I306614,I306640,);
nand I_17888 (I306648,I873926,I873920);
and I_17889 (I306665,I306648,I873932);
DFFARX1 I_17890 (I306665,I2507,I306614,I306691,);
nor I_17891 (I306582,I306691,I306640);
not I_17892 (I306713,I306691);
DFFARX1 I_17893 (I873935,I2507,I306614,I306739,);
nand I_17894 (I306747,I306739,I873926);
not I_17895 (I306764,I306747);
DFFARX1 I_17896 (I306764,I2507,I306614,I306790,);
not I_17897 (I306606,I306790);
nor I_17898 (I306812,I306640,I306747);
nor I_17899 (I306588,I306691,I306812);
DFFARX1 I_17900 (I873938,I2507,I306614,I306852,);
DFFARX1 I_17901 (I306852,I2507,I306614,I306869,);
not I_17902 (I306877,I306869);
not I_17903 (I306894,I306852);
nand I_17904 (I306591,I306894,I306713);
nand I_17905 (I306925,I873920,I873929);
and I_17906 (I306942,I306925,I873923);
DFFARX1 I_17907 (I306942,I2507,I306614,I306968,);
nor I_17908 (I306976,I306968,I306640);
DFFARX1 I_17909 (I306976,I2507,I306614,I306579,);
DFFARX1 I_17910 (I306968,I2507,I306614,I306597,);
nor I_17911 (I307021,I873941,I873929);
not I_17912 (I307038,I307021);
nor I_17913 (I306600,I306877,I307038);
nand I_17914 (I306585,I306894,I307038);
nor I_17915 (I306594,I306640,I307021);
DFFARX1 I_17916 (I307021,I2507,I306614,I306603,);
not I_17917 (I307141,I2514);
DFFARX1 I_17918 (I778009,I2507,I307141,I307167,);
nand I_17919 (I307175,I778012,I778006);
and I_17920 (I307192,I307175,I778018);
DFFARX1 I_17921 (I307192,I2507,I307141,I307218,);
nor I_17922 (I307109,I307218,I307167);
not I_17923 (I307240,I307218);
DFFARX1 I_17924 (I778021,I2507,I307141,I307266,);
nand I_17925 (I307274,I307266,I778012);
not I_17926 (I307291,I307274);
DFFARX1 I_17927 (I307291,I2507,I307141,I307317,);
not I_17928 (I307133,I307317);
nor I_17929 (I307339,I307167,I307274);
nor I_17930 (I307115,I307218,I307339);
DFFARX1 I_17931 (I778024,I2507,I307141,I307379,);
DFFARX1 I_17932 (I307379,I2507,I307141,I307396,);
not I_17933 (I307404,I307396);
not I_17934 (I307421,I307379);
nand I_17935 (I307118,I307421,I307240);
nand I_17936 (I307452,I778006,I778015);
and I_17937 (I307469,I307452,I778009);
DFFARX1 I_17938 (I307469,I2507,I307141,I307495,);
nor I_17939 (I307503,I307495,I307167);
DFFARX1 I_17940 (I307503,I2507,I307141,I307106,);
DFFARX1 I_17941 (I307495,I2507,I307141,I307124,);
nor I_17942 (I307548,I778027,I778015);
not I_17943 (I307565,I307548);
nor I_17944 (I307127,I307404,I307565);
nand I_17945 (I307112,I307421,I307565);
nor I_17946 (I307121,I307167,I307548);
DFFARX1 I_17947 (I307548,I2507,I307141,I307130,);
not I_17948 (I307668,I2514);
DFFARX1 I_17949 (I876031,I2507,I307668,I307694,);
nand I_17950 (I307702,I876034,I876028);
and I_17951 (I307719,I307702,I876040);
DFFARX1 I_17952 (I307719,I2507,I307668,I307745,);
nor I_17953 (I307636,I307745,I307694);
not I_17954 (I307767,I307745);
DFFARX1 I_17955 (I876043,I2507,I307668,I307793,);
nand I_17956 (I307801,I307793,I876034);
not I_17957 (I307818,I307801);
DFFARX1 I_17958 (I307818,I2507,I307668,I307844,);
not I_17959 (I307660,I307844);
nor I_17960 (I307866,I307694,I307801);
nor I_17961 (I307642,I307745,I307866);
DFFARX1 I_17962 (I876046,I2507,I307668,I307906,);
DFFARX1 I_17963 (I307906,I2507,I307668,I307923,);
not I_17964 (I307931,I307923);
not I_17965 (I307948,I307906);
nand I_17966 (I307645,I307948,I307767);
nand I_17967 (I307979,I876028,I876037);
and I_17968 (I307996,I307979,I876031);
DFFARX1 I_17969 (I307996,I2507,I307668,I308022,);
nor I_17970 (I308030,I308022,I307694);
DFFARX1 I_17971 (I308030,I2507,I307668,I307633,);
DFFARX1 I_17972 (I308022,I2507,I307668,I307651,);
nor I_17973 (I308075,I876049,I876037);
not I_17974 (I308092,I308075);
nor I_17975 (I307654,I307931,I308092);
nand I_17976 (I307639,I307948,I308092);
nor I_17977 (I307648,I307694,I308075);
DFFARX1 I_17978 (I308075,I2507,I307668,I307657,);
not I_17979 (I308195,I2514);
DFFARX1 I_17980 (I551547,I2507,I308195,I308221,);
nand I_17981 (I308229,I551532,I551535);
and I_17982 (I308246,I308229,I551550);
DFFARX1 I_17983 (I308246,I2507,I308195,I308272,);
nor I_17984 (I308163,I308272,I308221);
not I_17985 (I308294,I308272);
DFFARX1 I_17986 (I551544,I2507,I308195,I308320,);
nand I_17987 (I308328,I308320,I551535);
not I_17988 (I308345,I308328);
DFFARX1 I_17989 (I308345,I2507,I308195,I308371,);
not I_17990 (I308187,I308371);
nor I_17991 (I308393,I308221,I308328);
nor I_17992 (I308169,I308272,I308393);
DFFARX1 I_17993 (I551541,I2507,I308195,I308433,);
DFFARX1 I_17994 (I308433,I2507,I308195,I308450,);
not I_17995 (I308458,I308450);
not I_17996 (I308475,I308433);
nand I_17997 (I308172,I308475,I308294);
nand I_17998 (I308506,I551556,I551532);
and I_17999 (I308523,I308506,I551553);
DFFARX1 I_18000 (I308523,I2507,I308195,I308549,);
nor I_18001 (I308557,I308549,I308221);
DFFARX1 I_18002 (I308557,I2507,I308195,I308160,);
DFFARX1 I_18003 (I308549,I2507,I308195,I308178,);
nor I_18004 (I308602,I551538,I551532);
not I_18005 (I308619,I308602);
nor I_18006 (I308181,I308458,I308619);
nand I_18007 (I308166,I308475,I308619);
nor I_18008 (I308175,I308221,I308602);
DFFARX1 I_18009 (I308602,I2507,I308195,I308184,);
not I_18010 (I308722,I2514);
DFFARX1 I_18011 (I968324,I2507,I308722,I308748,);
nand I_18012 (I308756,I968321,I968339);
and I_18013 (I308773,I308756,I968330);
DFFARX1 I_18014 (I308773,I2507,I308722,I308799,);
nor I_18015 (I308690,I308799,I308748);
not I_18016 (I308821,I308799);
DFFARX1 I_18017 (I968345,I2507,I308722,I308847,);
nand I_18018 (I308855,I308847,I968327);
not I_18019 (I308872,I308855);
DFFARX1 I_18020 (I308872,I2507,I308722,I308898,);
not I_18021 (I308714,I308898);
nor I_18022 (I308920,I308748,I308855);
nor I_18023 (I308696,I308799,I308920);
DFFARX1 I_18024 (I968333,I2507,I308722,I308960,);
DFFARX1 I_18025 (I308960,I2507,I308722,I308977,);
not I_18026 (I308985,I308977);
not I_18027 (I309002,I308960);
nand I_18028 (I308699,I309002,I308821);
nand I_18029 (I309033,I968321,I968348);
and I_18030 (I309050,I309033,I968336);
DFFARX1 I_18031 (I309050,I2507,I308722,I309076,);
nor I_18032 (I309084,I309076,I308748);
DFFARX1 I_18033 (I309084,I2507,I308722,I308687,);
DFFARX1 I_18034 (I309076,I2507,I308722,I308705,);
nor I_18035 (I309129,I968342,I968348);
not I_18036 (I309146,I309129);
nor I_18037 (I308708,I308985,I309146);
nand I_18038 (I308693,I309002,I309146);
nor I_18039 (I308702,I308748,I309129);
DFFARX1 I_18040 (I309129,I2507,I308722,I308711,);
not I_18041 (I309249,I2514);
DFFARX1 I_18042 (I711072,I2507,I309249,I309275,);
nand I_18043 (I309283,I711063,I711078);
and I_18044 (I309300,I309283,I711084);
DFFARX1 I_18045 (I309300,I2507,I309249,I309326,);
nor I_18046 (I309217,I309326,I309275);
not I_18047 (I309348,I309326);
DFFARX1 I_18048 (I711069,I2507,I309249,I309374,);
nand I_18049 (I309382,I309374,I711063);
not I_18050 (I309399,I309382);
DFFARX1 I_18051 (I309399,I2507,I309249,I309425,);
not I_18052 (I309241,I309425);
nor I_18053 (I309447,I309275,I309382);
nor I_18054 (I309223,I309326,I309447);
DFFARX1 I_18055 (I711066,I2507,I309249,I309487,);
DFFARX1 I_18056 (I309487,I2507,I309249,I309504,);
not I_18057 (I309512,I309504);
not I_18058 (I309529,I309487);
nand I_18059 (I309226,I309529,I309348);
nand I_18060 (I309560,I711060,I711075);
and I_18061 (I309577,I309560,I711060);
DFFARX1 I_18062 (I309577,I2507,I309249,I309603,);
nor I_18063 (I309611,I309603,I309275);
DFFARX1 I_18064 (I309611,I2507,I309249,I309214,);
DFFARX1 I_18065 (I309603,I2507,I309249,I309232,);
nor I_18066 (I309656,I711081,I711075);
not I_18067 (I309673,I309656);
nor I_18068 (I309235,I309512,I309673);
nand I_18069 (I309220,I309529,I309673);
nor I_18070 (I309229,I309275,I309656);
DFFARX1 I_18071 (I309656,I2507,I309249,I309238,);
not I_18072 (I309776,I2514);
DFFARX1 I_18073 (I966386,I2507,I309776,I309802,);
nand I_18074 (I309810,I966383,I966401);
and I_18075 (I309827,I309810,I966392);
DFFARX1 I_18076 (I309827,I2507,I309776,I309853,);
nor I_18077 (I309744,I309853,I309802);
not I_18078 (I309875,I309853);
DFFARX1 I_18079 (I966407,I2507,I309776,I309901,);
nand I_18080 (I309909,I309901,I966389);
not I_18081 (I309926,I309909);
DFFARX1 I_18082 (I309926,I2507,I309776,I309952,);
not I_18083 (I309768,I309952);
nor I_18084 (I309974,I309802,I309909);
nor I_18085 (I309750,I309853,I309974);
DFFARX1 I_18086 (I966395,I2507,I309776,I310014,);
DFFARX1 I_18087 (I310014,I2507,I309776,I310031,);
not I_18088 (I310039,I310031);
not I_18089 (I310056,I310014);
nand I_18090 (I309753,I310056,I309875);
nand I_18091 (I310087,I966383,I966410);
and I_18092 (I310104,I310087,I966398);
DFFARX1 I_18093 (I310104,I2507,I309776,I310130,);
nor I_18094 (I310138,I310130,I309802);
DFFARX1 I_18095 (I310138,I2507,I309776,I309741,);
DFFARX1 I_18096 (I310130,I2507,I309776,I309759,);
nor I_18097 (I310183,I966404,I966410);
not I_18098 (I310200,I310183);
nor I_18099 (I309762,I310039,I310200);
nand I_18100 (I309747,I310056,I310200);
nor I_18101 (I309756,I309802,I310183);
DFFARX1 I_18102 (I310183,I2507,I309776,I309765,);
not I_18103 (I310303,I2514);
DFFARX1 I_18104 (I436539,I2507,I310303,I310329,);
nand I_18105 (I310337,I436551,I436530);
and I_18106 (I310354,I310337,I436554);
DFFARX1 I_18107 (I310354,I2507,I310303,I310380,);
nor I_18108 (I310271,I310380,I310329);
not I_18109 (I310402,I310380);
DFFARX1 I_18110 (I436545,I2507,I310303,I310428,);
nand I_18111 (I310436,I310428,I436527);
not I_18112 (I310453,I310436);
DFFARX1 I_18113 (I310453,I2507,I310303,I310479,);
not I_18114 (I310295,I310479);
nor I_18115 (I310501,I310329,I310436);
nor I_18116 (I310277,I310380,I310501);
DFFARX1 I_18117 (I436542,I2507,I310303,I310541,);
DFFARX1 I_18118 (I310541,I2507,I310303,I310558,);
not I_18119 (I310566,I310558);
not I_18120 (I310583,I310541);
nand I_18121 (I310280,I310583,I310402);
nand I_18122 (I310614,I436527,I436533);
and I_18123 (I310631,I310614,I436536);
DFFARX1 I_18124 (I310631,I2507,I310303,I310657,);
nor I_18125 (I310665,I310657,I310329);
DFFARX1 I_18126 (I310665,I2507,I310303,I310268,);
DFFARX1 I_18127 (I310657,I2507,I310303,I310286,);
nor I_18128 (I310710,I436548,I436533);
not I_18129 (I310727,I310710);
nor I_18130 (I310289,I310566,I310727);
nand I_18131 (I310274,I310583,I310727);
nor I_18132 (I310283,I310329,I310710);
DFFARX1 I_18133 (I310710,I2507,I310303,I310292,);
not I_18134 (I310830,I2514);
DFFARX1 I_18135 (I1099408,I2507,I310830,I310856,);
nand I_18136 (I310864,I1099423,I1099408);
and I_18137 (I310881,I310864,I1099426);
DFFARX1 I_18138 (I310881,I2507,I310830,I310907,);
nor I_18139 (I310798,I310907,I310856);
not I_18140 (I310929,I310907);
DFFARX1 I_18141 (I1099432,I2507,I310830,I310955,);
nand I_18142 (I310963,I310955,I1099414);
not I_18143 (I310980,I310963);
DFFARX1 I_18144 (I310980,I2507,I310830,I311006,);
not I_18145 (I310822,I311006);
nor I_18146 (I311028,I310856,I310963);
nor I_18147 (I310804,I310907,I311028);
DFFARX1 I_18148 (I1099411,I2507,I310830,I311068,);
DFFARX1 I_18149 (I311068,I2507,I310830,I311085,);
not I_18150 (I311093,I311085);
not I_18151 (I311110,I311068);
nand I_18152 (I310807,I311110,I310929);
nand I_18153 (I311141,I1099411,I1099417);
and I_18154 (I311158,I311141,I1099429);
DFFARX1 I_18155 (I311158,I2507,I310830,I311184,);
nor I_18156 (I311192,I311184,I310856);
DFFARX1 I_18157 (I311192,I2507,I310830,I310795,);
DFFARX1 I_18158 (I311184,I2507,I310830,I310813,);
nor I_18159 (I311237,I1099420,I1099417);
not I_18160 (I311254,I311237);
nor I_18161 (I310816,I311093,I311254);
nand I_18162 (I310801,I311110,I311254);
nor I_18163 (I310810,I310856,I311237);
DFFARX1 I_18164 (I311237,I2507,I310830,I310819,);
not I_18165 (I311357,I2514);
DFFARX1 I_18166 (I130224,I2507,I311357,I311383,);
nand I_18167 (I311391,I130236,I130245);
and I_18168 (I311408,I311391,I130224);
DFFARX1 I_18169 (I311408,I2507,I311357,I311434,);
nor I_18170 (I311325,I311434,I311383);
not I_18171 (I311456,I311434);
DFFARX1 I_18172 (I130239,I2507,I311357,I311482,);
nand I_18173 (I311490,I311482,I130227);
not I_18174 (I311507,I311490);
DFFARX1 I_18175 (I311507,I2507,I311357,I311533,);
not I_18176 (I311349,I311533);
nor I_18177 (I311555,I311383,I311490);
nor I_18178 (I311331,I311434,I311555);
DFFARX1 I_18179 (I130230,I2507,I311357,I311595,);
DFFARX1 I_18180 (I311595,I2507,I311357,I311612,);
not I_18181 (I311620,I311612);
not I_18182 (I311637,I311595);
nand I_18183 (I311334,I311637,I311456);
nand I_18184 (I311668,I130221,I130221);
and I_18185 (I311685,I311668,I130233);
DFFARX1 I_18186 (I311685,I2507,I311357,I311711,);
nor I_18187 (I311719,I311711,I311383);
DFFARX1 I_18188 (I311719,I2507,I311357,I311322,);
DFFARX1 I_18189 (I311711,I2507,I311357,I311340,);
nor I_18190 (I311764,I130242,I130221);
not I_18191 (I311781,I311764);
nor I_18192 (I311343,I311620,I311781);
nand I_18193 (I311328,I311637,I311781);
nor I_18194 (I311337,I311383,I311764);
DFFARX1 I_18195 (I311764,I2507,I311357,I311346,);
not I_18196 (I311884,I2514);
DFFARX1 I_18197 (I1250964,I2507,I311884,I311910,);
nand I_18198 (I311918,I1250946,I1250970);
and I_18199 (I311935,I311918,I1250961);
DFFARX1 I_18200 (I311935,I2507,I311884,I311961,);
nor I_18201 (I311852,I311961,I311910);
not I_18202 (I311983,I311961);
DFFARX1 I_18203 (I1250967,I2507,I311884,I312009,);
nand I_18204 (I312017,I312009,I1250955);
not I_18205 (I312034,I312017);
DFFARX1 I_18206 (I312034,I2507,I311884,I312060,);
not I_18207 (I311876,I312060);
nor I_18208 (I312082,I311910,I312017);
nor I_18209 (I311858,I311961,I312082);
DFFARX1 I_18210 (I1250946,I2507,I311884,I312122,);
DFFARX1 I_18211 (I312122,I2507,I311884,I312139,);
not I_18212 (I312147,I312139);
not I_18213 (I312164,I312122);
nand I_18214 (I311861,I312164,I311983);
nand I_18215 (I312195,I1250952,I1250949);
and I_18216 (I312212,I312195,I1250958);
DFFARX1 I_18217 (I312212,I2507,I311884,I312238,);
nor I_18218 (I312246,I312238,I311910);
DFFARX1 I_18219 (I312246,I2507,I311884,I311849,);
DFFARX1 I_18220 (I312238,I2507,I311884,I311867,);
nor I_18221 (I312291,I1250949,I1250949);
not I_18222 (I312308,I312291);
nor I_18223 (I311870,I312147,I312308);
nand I_18224 (I311855,I312164,I312308);
nor I_18225 (I311864,I311910,I312291);
DFFARX1 I_18226 (I312291,I2507,I311884,I311873,);
not I_18227 (I312411,I2514);
DFFARX1 I_18228 (I1061838,I2507,I312411,I312437,);
nand I_18229 (I312445,I1061853,I1061838);
and I_18230 (I312462,I312445,I1061856);
DFFARX1 I_18231 (I312462,I2507,I312411,I312488,);
nor I_18232 (I312379,I312488,I312437);
not I_18233 (I312510,I312488);
DFFARX1 I_18234 (I1061862,I2507,I312411,I312536,);
nand I_18235 (I312544,I312536,I1061844);
not I_18236 (I312561,I312544);
DFFARX1 I_18237 (I312561,I2507,I312411,I312587,);
not I_18238 (I312403,I312587);
nor I_18239 (I312609,I312437,I312544);
nor I_18240 (I312385,I312488,I312609);
DFFARX1 I_18241 (I1061841,I2507,I312411,I312649,);
DFFARX1 I_18242 (I312649,I2507,I312411,I312666,);
not I_18243 (I312674,I312666);
not I_18244 (I312691,I312649);
nand I_18245 (I312388,I312691,I312510);
nand I_18246 (I312722,I1061841,I1061847);
and I_18247 (I312739,I312722,I1061859);
DFFARX1 I_18248 (I312739,I2507,I312411,I312765,);
nor I_18249 (I312773,I312765,I312437);
DFFARX1 I_18250 (I312773,I2507,I312411,I312376,);
DFFARX1 I_18251 (I312765,I2507,I312411,I312394,);
nor I_18252 (I312818,I1061850,I1061847);
not I_18253 (I312835,I312818);
nor I_18254 (I312397,I312674,I312835);
nand I_18255 (I312382,I312691,I312835);
nor I_18256 (I312391,I312437,I312818);
DFFARX1 I_18257 (I312818,I2507,I312411,I312400,);
not I_18258 (I312938,I2514);
DFFARX1 I_18259 (I952174,I2507,I312938,I312964,);
nand I_18260 (I312972,I952171,I952189);
and I_18261 (I312989,I312972,I952180);
DFFARX1 I_18262 (I312989,I2507,I312938,I313015,);
nor I_18263 (I312906,I313015,I312964);
not I_18264 (I313037,I313015);
DFFARX1 I_18265 (I952195,I2507,I312938,I313063,);
nand I_18266 (I313071,I313063,I952177);
not I_18267 (I313088,I313071);
DFFARX1 I_18268 (I313088,I2507,I312938,I313114,);
not I_18269 (I312930,I313114);
nor I_18270 (I313136,I312964,I313071);
nor I_18271 (I312912,I313015,I313136);
DFFARX1 I_18272 (I952183,I2507,I312938,I313176,);
DFFARX1 I_18273 (I313176,I2507,I312938,I313193,);
not I_18274 (I313201,I313193);
not I_18275 (I313218,I313176);
nand I_18276 (I312915,I313218,I313037);
nand I_18277 (I313249,I952171,I952198);
and I_18278 (I313266,I313249,I952186);
DFFARX1 I_18279 (I313266,I2507,I312938,I313292,);
nor I_18280 (I313300,I313292,I312964);
DFFARX1 I_18281 (I313300,I2507,I312938,I312903,);
DFFARX1 I_18282 (I313292,I2507,I312938,I312921,);
nor I_18283 (I313345,I952192,I952198);
not I_18284 (I313362,I313345);
nor I_18285 (I312924,I313201,I313362);
nand I_18286 (I312909,I313218,I313362);
nor I_18287 (I312918,I312964,I313345);
DFFARX1 I_18288 (I313345,I2507,I312938,I312927,);
not I_18289 (I313465,I2514);
DFFARX1 I_18290 (I572933,I2507,I313465,I313491,);
nand I_18291 (I313499,I572918,I572921);
and I_18292 (I313516,I313499,I572936);
DFFARX1 I_18293 (I313516,I2507,I313465,I313542,);
nor I_18294 (I313433,I313542,I313491);
not I_18295 (I313564,I313542);
DFFARX1 I_18296 (I572930,I2507,I313465,I313590,);
nand I_18297 (I313598,I313590,I572921);
not I_18298 (I313615,I313598);
DFFARX1 I_18299 (I313615,I2507,I313465,I313641,);
not I_18300 (I313457,I313641);
nor I_18301 (I313663,I313491,I313598);
nor I_18302 (I313439,I313542,I313663);
DFFARX1 I_18303 (I572927,I2507,I313465,I313703,);
DFFARX1 I_18304 (I313703,I2507,I313465,I313720,);
not I_18305 (I313728,I313720);
not I_18306 (I313745,I313703);
nand I_18307 (I313442,I313745,I313564);
nand I_18308 (I313776,I572942,I572918);
and I_18309 (I313793,I313776,I572939);
DFFARX1 I_18310 (I313793,I2507,I313465,I313819,);
nor I_18311 (I313827,I313819,I313491);
DFFARX1 I_18312 (I313827,I2507,I313465,I313430,);
DFFARX1 I_18313 (I313819,I2507,I313465,I313448,);
nor I_18314 (I313872,I572924,I572918);
not I_18315 (I313889,I313872);
nor I_18316 (I313451,I313728,I313889);
nand I_18317 (I313436,I313745,I313889);
nor I_18318 (I313445,I313491,I313872);
DFFARX1 I_18319 (I313872,I2507,I313465,I313454,);
not I_18320 (I313992,I2514);
DFFARX1 I_18321 (I12052,I2507,I313992,I314018,);
nand I_18322 (I314026,I12043,I12046);
and I_18323 (I314043,I314026,I12037);
DFFARX1 I_18324 (I314043,I2507,I313992,I314069,);
nor I_18325 (I313960,I314069,I314018);
not I_18326 (I314091,I314069);
DFFARX1 I_18327 (I12043,I2507,I313992,I314117,);
nand I_18328 (I314125,I314117,I12049);
not I_18329 (I314142,I314125);
DFFARX1 I_18330 (I314142,I2507,I313992,I314168,);
not I_18331 (I313984,I314168);
nor I_18332 (I314190,I314018,I314125);
nor I_18333 (I313966,I314069,I314190);
DFFARX1 I_18334 (I12040,I2507,I313992,I314230,);
DFFARX1 I_18335 (I314230,I2507,I313992,I314247,);
not I_18336 (I314255,I314247);
not I_18337 (I314272,I314230);
nand I_18338 (I313969,I314272,I314091);
nand I_18339 (I314303,I12040,I12055);
and I_18340 (I314320,I314303,I12037);
DFFARX1 I_18341 (I314320,I2507,I313992,I314346,);
nor I_18342 (I314354,I314346,I314018);
DFFARX1 I_18343 (I314354,I2507,I313992,I313957,);
DFFARX1 I_18344 (I314346,I2507,I313992,I313975,);
nor I_18345 (I314399,I12058,I12055);
not I_18346 (I314416,I314399);
nor I_18347 (I313978,I314255,I314416);
nand I_18348 (I313963,I314272,I314416);
nor I_18349 (I313972,I314018,I314399);
DFFARX1 I_18350 (I314399,I2507,I313992,I313981,);
not I_18351 (I314519,I2514);
DFFARX1 I_18352 (I953466,I2507,I314519,I314545,);
nand I_18353 (I314553,I953463,I953481);
and I_18354 (I314570,I314553,I953472);
DFFARX1 I_18355 (I314570,I2507,I314519,I314596,);
nor I_18356 (I314487,I314596,I314545);
not I_18357 (I314618,I314596);
DFFARX1 I_18358 (I953487,I2507,I314519,I314644,);
nand I_18359 (I314652,I314644,I953469);
not I_18360 (I314669,I314652);
DFFARX1 I_18361 (I314669,I2507,I314519,I314695,);
not I_18362 (I314511,I314695);
nor I_18363 (I314717,I314545,I314652);
nor I_18364 (I314493,I314596,I314717);
DFFARX1 I_18365 (I953475,I2507,I314519,I314757,);
DFFARX1 I_18366 (I314757,I2507,I314519,I314774,);
not I_18367 (I314782,I314774);
not I_18368 (I314799,I314757);
nand I_18369 (I314496,I314799,I314618);
nand I_18370 (I314830,I953463,I953490);
and I_18371 (I314847,I314830,I953478);
DFFARX1 I_18372 (I314847,I2507,I314519,I314873,);
nor I_18373 (I314881,I314873,I314545);
DFFARX1 I_18374 (I314881,I2507,I314519,I314484,);
DFFARX1 I_18375 (I314873,I2507,I314519,I314502,);
nor I_18376 (I314926,I953484,I953490);
not I_18377 (I314943,I314926);
nor I_18378 (I314505,I314782,I314943);
nand I_18379 (I314490,I314799,I314943);
nor I_18380 (I314499,I314545,I314926);
DFFARX1 I_18381 (I314926,I2507,I314519,I314508,);
not I_18382 (I315046,I2514);
DFFARX1 I_18383 (I53809,I2507,I315046,I315072,);
nand I_18384 (I315080,I53821,I53830);
and I_18385 (I315097,I315080,I53809);
DFFARX1 I_18386 (I315097,I2507,I315046,I315123,);
nor I_18387 (I315014,I315123,I315072);
not I_18388 (I315145,I315123);
DFFARX1 I_18389 (I53824,I2507,I315046,I315171,);
nand I_18390 (I315179,I315171,I53812);
not I_18391 (I315196,I315179);
DFFARX1 I_18392 (I315196,I2507,I315046,I315222,);
not I_18393 (I315038,I315222);
nor I_18394 (I315244,I315072,I315179);
nor I_18395 (I315020,I315123,I315244);
DFFARX1 I_18396 (I53815,I2507,I315046,I315284,);
DFFARX1 I_18397 (I315284,I2507,I315046,I315301,);
not I_18398 (I315309,I315301);
not I_18399 (I315326,I315284);
nand I_18400 (I315023,I315326,I315145);
nand I_18401 (I315357,I53806,I53806);
and I_18402 (I315374,I315357,I53818);
DFFARX1 I_18403 (I315374,I2507,I315046,I315400,);
nor I_18404 (I315408,I315400,I315072);
DFFARX1 I_18405 (I315408,I2507,I315046,I315011,);
DFFARX1 I_18406 (I315400,I2507,I315046,I315029,);
nor I_18407 (I315453,I53827,I53806);
not I_18408 (I315470,I315453);
nor I_18409 (I315032,I315309,I315470);
nand I_18410 (I315017,I315326,I315470);
nor I_18411 (I315026,I315072,I315453);
DFFARX1 I_18412 (I315453,I2507,I315046,I315035,);
not I_18413 (I315573,I2514);
DFFARX1 I_18414 (I804359,I2507,I315573,I315599,);
nand I_18415 (I315607,I804362,I804356);
and I_18416 (I315624,I315607,I804368);
DFFARX1 I_18417 (I315624,I2507,I315573,I315650,);
nor I_18418 (I315541,I315650,I315599);
not I_18419 (I315672,I315650);
DFFARX1 I_18420 (I804371,I2507,I315573,I315698,);
nand I_18421 (I315706,I315698,I804362);
not I_18422 (I315723,I315706);
DFFARX1 I_18423 (I315723,I2507,I315573,I315749,);
not I_18424 (I315565,I315749);
nor I_18425 (I315771,I315599,I315706);
nor I_18426 (I315547,I315650,I315771);
DFFARX1 I_18427 (I804374,I2507,I315573,I315811,);
DFFARX1 I_18428 (I315811,I2507,I315573,I315828,);
not I_18429 (I315836,I315828);
not I_18430 (I315853,I315811);
nand I_18431 (I315550,I315853,I315672);
nand I_18432 (I315884,I804356,I804365);
and I_18433 (I315901,I315884,I804359);
DFFARX1 I_18434 (I315901,I2507,I315573,I315927,);
nor I_18435 (I315935,I315927,I315599);
DFFARX1 I_18436 (I315935,I2507,I315573,I315538,);
DFFARX1 I_18437 (I315927,I2507,I315573,I315556,);
nor I_18438 (I315980,I804377,I804365);
not I_18439 (I315997,I315980);
nor I_18440 (I315559,I315836,I315997);
nand I_18441 (I315544,I315853,I315997);
nor I_18442 (I315553,I315599,I315980);
DFFARX1 I_18443 (I315980,I2507,I315573,I315562,);
not I_18444 (I316100,I2514);
DFFARX1 I_18445 (I1311878,I2507,I316100,I316126,);
nand I_18446 (I316134,I1311857,I1311857);
and I_18447 (I316151,I316134,I1311884);
DFFARX1 I_18448 (I316151,I2507,I316100,I316177,);
nor I_18449 (I316068,I316177,I316126);
not I_18450 (I316199,I316177);
DFFARX1 I_18451 (I1311872,I2507,I316100,I316225,);
nand I_18452 (I316233,I316225,I1311875);
not I_18453 (I316250,I316233);
DFFARX1 I_18454 (I316250,I2507,I316100,I316276,);
not I_18455 (I316092,I316276);
nor I_18456 (I316298,I316126,I316233);
nor I_18457 (I316074,I316177,I316298);
DFFARX1 I_18458 (I1311866,I2507,I316100,I316338,);
DFFARX1 I_18459 (I316338,I2507,I316100,I316355,);
not I_18460 (I316363,I316355);
not I_18461 (I316380,I316338);
nand I_18462 (I316077,I316380,I316199);
nand I_18463 (I316411,I1311863,I1311860);
and I_18464 (I316428,I316411,I1311881);
DFFARX1 I_18465 (I316428,I2507,I316100,I316454,);
nor I_18466 (I316462,I316454,I316126);
DFFARX1 I_18467 (I316462,I2507,I316100,I316065,);
DFFARX1 I_18468 (I316454,I2507,I316100,I316083,);
nor I_18469 (I316507,I1311869,I1311860);
not I_18470 (I316524,I316507);
nor I_18471 (I316086,I316363,I316524);
nand I_18472 (I316071,I316380,I316524);
nor I_18473 (I316080,I316126,I316507);
DFFARX1 I_18474 (I316507,I2507,I316100,I316089,);
not I_18475 (I316627,I2514);
DFFARX1 I_18476 (I1384468,I2507,I316627,I316653,);
nand I_18477 (I316661,I1384447,I1384447);
and I_18478 (I316678,I316661,I1384474);
DFFARX1 I_18479 (I316678,I2507,I316627,I316704,);
nor I_18480 (I316595,I316704,I316653);
not I_18481 (I316726,I316704);
DFFARX1 I_18482 (I1384462,I2507,I316627,I316752,);
nand I_18483 (I316760,I316752,I1384465);
not I_18484 (I316777,I316760);
DFFARX1 I_18485 (I316777,I2507,I316627,I316803,);
not I_18486 (I316619,I316803);
nor I_18487 (I316825,I316653,I316760);
nor I_18488 (I316601,I316704,I316825);
DFFARX1 I_18489 (I1384456,I2507,I316627,I316865,);
DFFARX1 I_18490 (I316865,I2507,I316627,I316882,);
not I_18491 (I316890,I316882);
not I_18492 (I316907,I316865);
nand I_18493 (I316604,I316907,I316726);
nand I_18494 (I316938,I1384453,I1384450);
and I_18495 (I316955,I316938,I1384471);
DFFARX1 I_18496 (I316955,I2507,I316627,I316981,);
nor I_18497 (I316989,I316981,I316653);
DFFARX1 I_18498 (I316989,I2507,I316627,I316592,);
DFFARX1 I_18499 (I316981,I2507,I316627,I316610,);
nor I_18500 (I317034,I1384459,I1384450);
not I_18501 (I317051,I317034);
nor I_18502 (I316613,I316890,I317051);
nand I_18503 (I316598,I316907,I317051);
nor I_18504 (I316607,I316653,I317034);
DFFARX1 I_18505 (I317034,I2507,I316627,I316616,);
not I_18506 (I317154,I2514);
DFFARX1 I_18507 (I1052219,I2507,I317154,I317180,);
nand I_18508 (I317188,I1052216,I1052219);
and I_18509 (I317205,I317188,I1052228);
DFFARX1 I_18510 (I317205,I2507,I317154,I317231,);
nor I_18511 (I317122,I317231,I317180);
not I_18512 (I317253,I317231);
DFFARX1 I_18513 (I1052216,I2507,I317154,I317279,);
nand I_18514 (I317287,I317279,I1052234);
not I_18515 (I317304,I317287);
DFFARX1 I_18516 (I317304,I2507,I317154,I317330,);
not I_18517 (I317146,I317330);
nor I_18518 (I317352,I317180,I317287);
nor I_18519 (I317128,I317231,I317352);
DFFARX1 I_18520 (I1052222,I2507,I317154,I317392,);
DFFARX1 I_18521 (I317392,I2507,I317154,I317409,);
not I_18522 (I317417,I317409);
not I_18523 (I317434,I317392);
nand I_18524 (I317131,I317434,I317253);
nand I_18525 (I317465,I1052231,I1052237);
and I_18526 (I317482,I317465,I1052222);
DFFARX1 I_18527 (I317482,I2507,I317154,I317508,);
nor I_18528 (I317516,I317508,I317180);
DFFARX1 I_18529 (I317516,I2507,I317154,I317119,);
DFFARX1 I_18530 (I317508,I2507,I317154,I317137,);
nor I_18531 (I317561,I1052225,I1052237);
not I_18532 (I317578,I317561);
nor I_18533 (I317140,I317417,I317578);
nand I_18534 (I317125,I317434,I317578);
nor I_18535 (I317134,I317180,I317561);
DFFARX1 I_18536 (I317561,I2507,I317154,I317143,);
not I_18537 (I317681,I2514);
DFFARX1 I_18538 (I83321,I2507,I317681,I317707,);
nand I_18539 (I317715,I83333,I83342);
and I_18540 (I317732,I317715,I83321);
DFFARX1 I_18541 (I317732,I2507,I317681,I317758,);
nor I_18542 (I317649,I317758,I317707);
not I_18543 (I317780,I317758);
DFFARX1 I_18544 (I83336,I2507,I317681,I317806,);
nand I_18545 (I317814,I317806,I83324);
not I_18546 (I317831,I317814);
DFFARX1 I_18547 (I317831,I2507,I317681,I317857,);
not I_18548 (I317673,I317857);
nor I_18549 (I317879,I317707,I317814);
nor I_18550 (I317655,I317758,I317879);
DFFARX1 I_18551 (I83327,I2507,I317681,I317919,);
DFFARX1 I_18552 (I317919,I2507,I317681,I317936,);
not I_18553 (I317944,I317936);
not I_18554 (I317961,I317919);
nand I_18555 (I317658,I317961,I317780);
nand I_18556 (I317992,I83318,I83318);
and I_18557 (I318009,I317992,I83330);
DFFARX1 I_18558 (I318009,I2507,I317681,I318035,);
nor I_18559 (I318043,I318035,I317707);
DFFARX1 I_18560 (I318043,I2507,I317681,I317646,);
DFFARX1 I_18561 (I318035,I2507,I317681,I317664,);
nor I_18562 (I318088,I83339,I83318);
not I_18563 (I318105,I318088);
nor I_18564 (I317667,I317944,I318105);
nand I_18565 (I317652,I317961,I318105);
nor I_18566 (I317661,I317707,I318088);
DFFARX1 I_18567 (I318088,I2507,I317681,I317670,);
not I_18568 (I318208,I2514);
DFFARX1 I_18569 (I1179750,I2507,I318208,I318234,);
nand I_18570 (I318242,I1179765,I1179750);
and I_18571 (I318259,I318242,I1179768);
DFFARX1 I_18572 (I318259,I2507,I318208,I318285,);
nor I_18573 (I318176,I318285,I318234);
not I_18574 (I318307,I318285);
DFFARX1 I_18575 (I1179774,I2507,I318208,I318333,);
nand I_18576 (I318341,I318333,I1179756);
not I_18577 (I318358,I318341);
DFFARX1 I_18578 (I318358,I2507,I318208,I318384,);
not I_18579 (I318200,I318384);
nor I_18580 (I318406,I318234,I318341);
nor I_18581 (I318182,I318285,I318406);
DFFARX1 I_18582 (I1179753,I2507,I318208,I318446,);
DFFARX1 I_18583 (I318446,I2507,I318208,I318463,);
not I_18584 (I318471,I318463);
not I_18585 (I318488,I318446);
nand I_18586 (I318185,I318488,I318307);
nand I_18587 (I318519,I1179753,I1179759);
and I_18588 (I318536,I318519,I1179771);
DFFARX1 I_18589 (I318536,I2507,I318208,I318562,);
nor I_18590 (I318570,I318562,I318234);
DFFARX1 I_18591 (I318570,I2507,I318208,I318173,);
DFFARX1 I_18592 (I318562,I2507,I318208,I318191,);
nor I_18593 (I318615,I1179762,I1179759);
not I_18594 (I318632,I318615);
nor I_18595 (I318194,I318471,I318632);
nand I_18596 (I318179,I318488,I318632);
nor I_18597 (I318188,I318234,I318615);
DFFARX1 I_18598 (I318615,I2507,I318208,I318197,);
not I_18599 (I318735,I2514);
DFFARX1 I_18600 (I1003854,I2507,I318735,I318761,);
nand I_18601 (I318769,I1003851,I1003869);
and I_18602 (I318786,I318769,I1003860);
DFFARX1 I_18603 (I318786,I2507,I318735,I318812,);
nor I_18604 (I318703,I318812,I318761);
not I_18605 (I318834,I318812);
DFFARX1 I_18606 (I1003875,I2507,I318735,I318860,);
nand I_18607 (I318868,I318860,I1003857);
not I_18608 (I318885,I318868);
DFFARX1 I_18609 (I318885,I2507,I318735,I318911,);
not I_18610 (I318727,I318911);
nor I_18611 (I318933,I318761,I318868);
nor I_18612 (I318709,I318812,I318933);
DFFARX1 I_18613 (I1003863,I2507,I318735,I318973,);
DFFARX1 I_18614 (I318973,I2507,I318735,I318990,);
not I_18615 (I318998,I318990);
not I_18616 (I319015,I318973);
nand I_18617 (I318712,I319015,I318834);
nand I_18618 (I319046,I1003851,I1003878);
and I_18619 (I319063,I319046,I1003866);
DFFARX1 I_18620 (I319063,I2507,I318735,I319089,);
nor I_18621 (I319097,I319089,I318761);
DFFARX1 I_18622 (I319097,I2507,I318735,I318700,);
DFFARX1 I_18623 (I319089,I2507,I318735,I318718,);
nor I_18624 (I319142,I1003872,I1003878);
not I_18625 (I319159,I319142);
nor I_18626 (I318721,I318998,I319159);
nand I_18627 (I318706,I319015,I319159);
nor I_18628 (I318715,I318761,I319142);
DFFARX1 I_18629 (I319142,I2507,I318735,I318724,);
not I_18630 (I319262,I2514);
DFFARX1 I_18631 (I1152006,I2507,I319262,I319288,);
nand I_18632 (I319296,I1152021,I1152006);
and I_18633 (I319313,I319296,I1152024);
DFFARX1 I_18634 (I319313,I2507,I319262,I319339,);
nor I_18635 (I319230,I319339,I319288);
not I_18636 (I319361,I319339);
DFFARX1 I_18637 (I1152030,I2507,I319262,I319387,);
nand I_18638 (I319395,I319387,I1152012);
not I_18639 (I319412,I319395);
DFFARX1 I_18640 (I319412,I2507,I319262,I319438,);
not I_18641 (I319254,I319438);
nor I_18642 (I319460,I319288,I319395);
nor I_18643 (I319236,I319339,I319460);
DFFARX1 I_18644 (I1152009,I2507,I319262,I319500,);
DFFARX1 I_18645 (I319500,I2507,I319262,I319517,);
not I_18646 (I319525,I319517);
not I_18647 (I319542,I319500);
nand I_18648 (I319239,I319542,I319361);
nand I_18649 (I319573,I1152009,I1152015);
and I_18650 (I319590,I319573,I1152027);
DFFARX1 I_18651 (I319590,I2507,I319262,I319616,);
nor I_18652 (I319624,I319616,I319288);
DFFARX1 I_18653 (I319624,I2507,I319262,I319227,);
DFFARX1 I_18654 (I319616,I2507,I319262,I319245,);
nor I_18655 (I319669,I1152018,I1152015);
not I_18656 (I319686,I319669);
nor I_18657 (I319248,I319525,I319686);
nand I_18658 (I319233,I319542,I319686);
nor I_18659 (I319242,I319288,I319669);
DFFARX1 I_18660 (I319669,I2507,I319262,I319251,);
not I_18661 (I319789,I2514);
DFFARX1 I_18662 (I412059,I2507,I319789,I319815,);
nand I_18663 (I319823,I412071,I412050);
and I_18664 (I319840,I319823,I412074);
DFFARX1 I_18665 (I319840,I2507,I319789,I319866,);
nor I_18666 (I319757,I319866,I319815);
not I_18667 (I319888,I319866);
DFFARX1 I_18668 (I412065,I2507,I319789,I319914,);
nand I_18669 (I319922,I319914,I412047);
not I_18670 (I319939,I319922);
DFFARX1 I_18671 (I319939,I2507,I319789,I319965,);
not I_18672 (I319781,I319965);
nor I_18673 (I319987,I319815,I319922);
nor I_18674 (I319763,I319866,I319987);
DFFARX1 I_18675 (I412062,I2507,I319789,I320027,);
DFFARX1 I_18676 (I320027,I2507,I319789,I320044,);
not I_18677 (I320052,I320044);
not I_18678 (I320069,I320027);
nand I_18679 (I319766,I320069,I319888);
nand I_18680 (I320100,I412047,I412053);
and I_18681 (I320117,I320100,I412056);
DFFARX1 I_18682 (I320117,I2507,I319789,I320143,);
nor I_18683 (I320151,I320143,I319815);
DFFARX1 I_18684 (I320151,I2507,I319789,I319754,);
DFFARX1 I_18685 (I320143,I2507,I319789,I319772,);
nor I_18686 (I320196,I412068,I412053);
not I_18687 (I320213,I320196);
nor I_18688 (I319775,I320052,I320213);
nand I_18689 (I319760,I320069,I320213);
nor I_18690 (I319769,I319815,I320196);
DFFARX1 I_18691 (I320196,I2507,I319789,I319778,);
not I_18692 (I320316,I2514);
DFFARX1 I_18693 (I535742,I2507,I320316,I320342,);
nand I_18694 (I320350,I535742,I535754);
and I_18695 (I320367,I320350,I535739);
DFFARX1 I_18696 (I320367,I2507,I320316,I320393,);
nor I_18697 (I320284,I320393,I320342);
not I_18698 (I320415,I320393);
DFFARX1 I_18699 (I535763,I2507,I320316,I320441,);
nand I_18700 (I320449,I320441,I535760);
not I_18701 (I320466,I320449);
DFFARX1 I_18702 (I320466,I2507,I320316,I320492,);
not I_18703 (I320308,I320492);
nor I_18704 (I320514,I320342,I320449);
nor I_18705 (I320290,I320393,I320514);
DFFARX1 I_18706 (I535751,I2507,I320316,I320554,);
DFFARX1 I_18707 (I320554,I2507,I320316,I320571,);
not I_18708 (I320579,I320571);
not I_18709 (I320596,I320554);
nand I_18710 (I320293,I320596,I320415);
nand I_18711 (I320627,I535739,I535748);
and I_18712 (I320644,I320627,I535757);
DFFARX1 I_18713 (I320644,I2507,I320316,I320670,);
nor I_18714 (I320678,I320670,I320342);
DFFARX1 I_18715 (I320678,I2507,I320316,I320281,);
DFFARX1 I_18716 (I320670,I2507,I320316,I320299,);
nor I_18717 (I320723,I535745,I535748);
not I_18718 (I320740,I320723);
nor I_18719 (I320302,I320579,I320740);
nand I_18720 (I320287,I320596,I320740);
nor I_18721 (I320296,I320342,I320723);
DFFARX1 I_18722 (I320723,I2507,I320316,I320305,);
not I_18723 (I320843,I2514);
DFFARX1 I_18724 (I1145648,I2507,I320843,I320869,);
nand I_18725 (I320877,I1145663,I1145648);
and I_18726 (I320894,I320877,I1145666);
DFFARX1 I_18727 (I320894,I2507,I320843,I320920,);
nor I_18728 (I320811,I320920,I320869);
not I_18729 (I320942,I320920);
DFFARX1 I_18730 (I1145672,I2507,I320843,I320968,);
nand I_18731 (I320976,I320968,I1145654);
not I_18732 (I320993,I320976);
DFFARX1 I_18733 (I320993,I2507,I320843,I321019,);
not I_18734 (I320835,I321019);
nor I_18735 (I321041,I320869,I320976);
nor I_18736 (I320817,I320920,I321041);
DFFARX1 I_18737 (I1145651,I2507,I320843,I321081,);
DFFARX1 I_18738 (I321081,I2507,I320843,I321098,);
not I_18739 (I321106,I321098);
not I_18740 (I321123,I321081);
nand I_18741 (I320820,I321123,I320942);
nand I_18742 (I321154,I1145651,I1145657);
and I_18743 (I321171,I321154,I1145669);
DFFARX1 I_18744 (I321171,I2507,I320843,I321197,);
nor I_18745 (I321205,I321197,I320869);
DFFARX1 I_18746 (I321205,I2507,I320843,I320808,);
DFFARX1 I_18747 (I321197,I2507,I320843,I320826,);
nor I_18748 (I321250,I1145660,I1145657);
not I_18749 (I321267,I321250);
nor I_18750 (I320829,I321106,I321267);
nand I_18751 (I320814,I321123,I321267);
nor I_18752 (I320823,I320869,I321250);
DFFARX1 I_18753 (I321250,I2507,I320843,I320832,);
not I_18754 (I321370,I2514);
DFFARX1 I_18755 (I849154,I2507,I321370,I321396,);
nand I_18756 (I321404,I849157,I849151);
and I_18757 (I321421,I321404,I849163);
DFFARX1 I_18758 (I321421,I2507,I321370,I321447,);
nor I_18759 (I321338,I321447,I321396);
not I_18760 (I321469,I321447);
DFFARX1 I_18761 (I849166,I2507,I321370,I321495,);
nand I_18762 (I321503,I321495,I849157);
not I_18763 (I321520,I321503);
DFFARX1 I_18764 (I321520,I2507,I321370,I321546,);
not I_18765 (I321362,I321546);
nor I_18766 (I321568,I321396,I321503);
nor I_18767 (I321344,I321447,I321568);
DFFARX1 I_18768 (I849169,I2507,I321370,I321608,);
DFFARX1 I_18769 (I321608,I2507,I321370,I321625,);
not I_18770 (I321633,I321625);
not I_18771 (I321650,I321608);
nand I_18772 (I321347,I321650,I321469);
nand I_18773 (I321681,I849151,I849160);
and I_18774 (I321698,I321681,I849154);
DFFARX1 I_18775 (I321698,I2507,I321370,I321724,);
nor I_18776 (I321732,I321724,I321396);
DFFARX1 I_18777 (I321732,I2507,I321370,I321335,);
DFFARX1 I_18778 (I321724,I2507,I321370,I321353,);
nor I_18779 (I321777,I849172,I849160);
not I_18780 (I321794,I321777);
nor I_18781 (I321356,I321633,I321794);
nand I_18782 (I321341,I321650,I321794);
nor I_18783 (I321350,I321396,I321777);
DFFARX1 I_18784 (I321777,I2507,I321370,I321359,);
not I_18785 (I321897,I2514);
DFFARX1 I_18786 (I382139,I2507,I321897,I321923,);
nand I_18787 (I321931,I382151,I382130);
and I_18788 (I321948,I321931,I382154);
DFFARX1 I_18789 (I321948,I2507,I321897,I321974,);
nor I_18790 (I321865,I321974,I321923);
not I_18791 (I321996,I321974);
DFFARX1 I_18792 (I382145,I2507,I321897,I322022,);
nand I_18793 (I322030,I322022,I382127);
not I_18794 (I322047,I322030);
DFFARX1 I_18795 (I322047,I2507,I321897,I322073,);
not I_18796 (I321889,I322073);
nor I_18797 (I322095,I321923,I322030);
nor I_18798 (I321871,I321974,I322095);
DFFARX1 I_18799 (I382142,I2507,I321897,I322135,);
DFFARX1 I_18800 (I322135,I2507,I321897,I322152,);
not I_18801 (I322160,I322152);
not I_18802 (I322177,I322135);
nand I_18803 (I321874,I322177,I321996);
nand I_18804 (I322208,I382127,I382133);
and I_18805 (I322225,I322208,I382136);
DFFARX1 I_18806 (I322225,I2507,I321897,I322251,);
nor I_18807 (I322259,I322251,I321923);
DFFARX1 I_18808 (I322259,I2507,I321897,I321862,);
DFFARX1 I_18809 (I322251,I2507,I321897,I321880,);
nor I_18810 (I322304,I382148,I382133);
not I_18811 (I322321,I322304);
nor I_18812 (I321883,I322160,I322321);
nand I_18813 (I321868,I322177,I322321);
nor I_18814 (I321877,I321923,I322304);
DFFARX1 I_18815 (I322304,I2507,I321897,I321886,);
not I_18816 (I322424,I2514);
DFFARX1 I_18817 (I175815,I2507,I322424,I322450,);
nand I_18818 (I322458,I175815,I175821);
and I_18819 (I322475,I322458,I175839);
DFFARX1 I_18820 (I322475,I2507,I322424,I322501,);
nor I_18821 (I322392,I322501,I322450);
not I_18822 (I322523,I322501);
DFFARX1 I_18823 (I175827,I2507,I322424,I322549,);
nand I_18824 (I322557,I322549,I175824);
not I_18825 (I322574,I322557);
DFFARX1 I_18826 (I322574,I2507,I322424,I322600,);
not I_18827 (I322416,I322600);
nor I_18828 (I322622,I322450,I322557);
nor I_18829 (I322398,I322501,I322622);
DFFARX1 I_18830 (I175833,I2507,I322424,I322662,);
DFFARX1 I_18831 (I322662,I2507,I322424,I322679,);
not I_18832 (I322687,I322679);
not I_18833 (I322704,I322662);
nand I_18834 (I322401,I322704,I322523);
nand I_18835 (I322735,I175818,I175818);
and I_18836 (I322752,I322735,I175830);
DFFARX1 I_18837 (I322752,I2507,I322424,I322778,);
nor I_18838 (I322786,I322778,I322450);
DFFARX1 I_18839 (I322786,I2507,I322424,I322389,);
DFFARX1 I_18840 (I322778,I2507,I322424,I322407,);
nor I_18841 (I322831,I175836,I175818);
not I_18842 (I322848,I322831);
nor I_18843 (I322410,I322687,I322848);
nand I_18844 (I322395,I322704,I322848);
nor I_18845 (I322404,I322450,I322831);
DFFARX1 I_18846 (I322831,I2507,I322424,I322413,);
not I_18847 (I322951,I2514);
DFFARX1 I_18848 (I1988,I2507,I322951,I322977,);
nand I_18849 (I322985,I2404,I1412);
and I_18850 (I323002,I322985,I1860);
DFFARX1 I_18851 (I323002,I2507,I322951,I323028,);
nor I_18852 (I322919,I323028,I322977);
not I_18853 (I323050,I323028);
DFFARX1 I_18854 (I1740,I2507,I322951,I323076,);
nand I_18855 (I323084,I323076,I1492);
not I_18856 (I323101,I323084);
DFFARX1 I_18857 (I323101,I2507,I322951,I323127,);
not I_18858 (I322943,I323127);
nor I_18859 (I323149,I322977,I323084);
nor I_18860 (I322925,I323028,I323149);
DFFARX1 I_18861 (I2332,I2507,I322951,I323189,);
DFFARX1 I_18862 (I323189,I2507,I322951,I323206,);
not I_18863 (I323214,I323206);
not I_18864 (I323231,I323189);
nand I_18865 (I322928,I323231,I323050);
nand I_18866 (I323262,I2228,I1500);
and I_18867 (I323279,I323262,I1396);
DFFARX1 I_18868 (I323279,I2507,I322951,I323305,);
nor I_18869 (I323313,I323305,I322977);
DFFARX1 I_18870 (I323313,I2507,I322951,I322916,);
DFFARX1 I_18871 (I323305,I2507,I322951,I322934,);
nor I_18872 (I323358,I1684,I1500);
not I_18873 (I323375,I323358);
nor I_18874 (I322937,I323214,I323375);
nand I_18875 (I322922,I323231,I323375);
nor I_18876 (I322931,I322977,I323358);
DFFARX1 I_18877 (I323358,I2507,I322951,I322940,);
not I_18878 (I323478,I2514);
DFFARX1 I_18879 (I1367213,I2507,I323478,I323504,);
nand I_18880 (I323512,I1367192,I1367192);
and I_18881 (I323529,I323512,I1367219);
DFFARX1 I_18882 (I323529,I2507,I323478,I323555,);
nor I_18883 (I323446,I323555,I323504);
not I_18884 (I323577,I323555);
DFFARX1 I_18885 (I1367207,I2507,I323478,I323603,);
nand I_18886 (I323611,I323603,I1367210);
not I_18887 (I323628,I323611);
DFFARX1 I_18888 (I323628,I2507,I323478,I323654,);
not I_18889 (I323470,I323654);
nor I_18890 (I323676,I323504,I323611);
nor I_18891 (I323452,I323555,I323676);
DFFARX1 I_18892 (I1367201,I2507,I323478,I323716,);
DFFARX1 I_18893 (I323716,I2507,I323478,I323733,);
not I_18894 (I323741,I323733);
not I_18895 (I323758,I323716);
nand I_18896 (I323455,I323758,I323577);
nand I_18897 (I323789,I1367198,I1367195);
and I_18898 (I323806,I323789,I1367216);
DFFARX1 I_18899 (I323806,I2507,I323478,I323832,);
nor I_18900 (I323840,I323832,I323504);
DFFARX1 I_18901 (I323840,I2507,I323478,I323443,);
DFFARX1 I_18902 (I323832,I2507,I323478,I323461,);
nor I_18903 (I323885,I1367204,I1367195);
not I_18904 (I323902,I323885);
nor I_18905 (I323464,I323741,I323902);
nand I_18906 (I323449,I323758,I323902);
nor I_18907 (I323458,I323504,I323885);
DFFARX1 I_18908 (I323885,I2507,I323478,I323467,);
not I_18909 (I324005,I2514);
DFFARX1 I_18910 (I451227,I2507,I324005,I324031,);
nand I_18911 (I324039,I451239,I451218);
and I_18912 (I324056,I324039,I451242);
DFFARX1 I_18913 (I324056,I2507,I324005,I324082,);
nor I_18914 (I323973,I324082,I324031);
not I_18915 (I324104,I324082);
DFFARX1 I_18916 (I451233,I2507,I324005,I324130,);
nand I_18917 (I324138,I324130,I451215);
not I_18918 (I324155,I324138);
DFFARX1 I_18919 (I324155,I2507,I324005,I324181,);
not I_18920 (I323997,I324181);
nor I_18921 (I324203,I324031,I324138);
nor I_18922 (I323979,I324082,I324203);
DFFARX1 I_18923 (I451230,I2507,I324005,I324243,);
DFFARX1 I_18924 (I324243,I2507,I324005,I324260,);
not I_18925 (I324268,I324260);
not I_18926 (I324285,I324243);
nand I_18927 (I323982,I324285,I324104);
nand I_18928 (I324316,I451215,I451221);
and I_18929 (I324333,I324316,I451224);
DFFARX1 I_18930 (I324333,I2507,I324005,I324359,);
nor I_18931 (I324367,I324359,I324031);
DFFARX1 I_18932 (I324367,I2507,I324005,I323970,);
DFFARX1 I_18933 (I324359,I2507,I324005,I323988,);
nor I_18934 (I324412,I451236,I451221);
not I_18935 (I324429,I324412);
nor I_18936 (I323991,I324268,I324429);
nand I_18937 (I323976,I324285,I324429);
nor I_18938 (I323985,I324031,I324412);
DFFARX1 I_18939 (I324412,I2507,I324005,I323994,);
not I_18940 (I324532,I2514);
DFFARX1 I_18941 (I774652,I2507,I324532,I324558,);
nand I_18942 (I324566,I774643,I774658);
and I_18943 (I324583,I324566,I774664);
DFFARX1 I_18944 (I324583,I2507,I324532,I324609,);
nor I_18945 (I324500,I324609,I324558);
not I_18946 (I324631,I324609);
DFFARX1 I_18947 (I774649,I2507,I324532,I324657,);
nand I_18948 (I324665,I324657,I774643);
not I_18949 (I324682,I324665);
DFFARX1 I_18950 (I324682,I2507,I324532,I324708,);
not I_18951 (I324524,I324708);
nor I_18952 (I324730,I324558,I324665);
nor I_18953 (I324506,I324609,I324730);
DFFARX1 I_18954 (I774646,I2507,I324532,I324770,);
DFFARX1 I_18955 (I324770,I2507,I324532,I324787,);
not I_18956 (I324795,I324787);
not I_18957 (I324812,I324770);
nand I_18958 (I324509,I324812,I324631);
nand I_18959 (I324843,I774640,I774655);
and I_18960 (I324860,I324843,I774640);
DFFARX1 I_18961 (I324860,I2507,I324532,I324886,);
nor I_18962 (I324894,I324886,I324558);
DFFARX1 I_18963 (I324894,I2507,I324532,I324497,);
DFFARX1 I_18964 (I324886,I2507,I324532,I324515,);
nor I_18965 (I324939,I774661,I774655);
not I_18966 (I324956,I324939);
nor I_18967 (I324518,I324795,I324956);
nand I_18968 (I324503,I324812,I324956);
nor I_18969 (I324512,I324558,I324939);
DFFARX1 I_18970 (I324939,I2507,I324532,I324521,);
not I_18971 (I325059,I2514);
DFFARX1 I_18972 (I90699,I2507,I325059,I325085,);
nand I_18973 (I325093,I90711,I90720);
and I_18974 (I325110,I325093,I90699);
DFFARX1 I_18975 (I325110,I2507,I325059,I325136,);
nor I_18976 (I325027,I325136,I325085);
not I_18977 (I325158,I325136);
DFFARX1 I_18978 (I90714,I2507,I325059,I325184,);
nand I_18979 (I325192,I325184,I90702);
not I_18980 (I325209,I325192);
DFFARX1 I_18981 (I325209,I2507,I325059,I325235,);
not I_18982 (I325051,I325235);
nor I_18983 (I325257,I325085,I325192);
nor I_18984 (I325033,I325136,I325257);
DFFARX1 I_18985 (I90705,I2507,I325059,I325297,);
DFFARX1 I_18986 (I325297,I2507,I325059,I325314,);
not I_18987 (I325322,I325314);
not I_18988 (I325339,I325297);
nand I_18989 (I325036,I325339,I325158);
nand I_18990 (I325370,I90696,I90696);
and I_18991 (I325387,I325370,I90708);
DFFARX1 I_18992 (I325387,I2507,I325059,I325413,);
nor I_18993 (I325421,I325413,I325085);
DFFARX1 I_18994 (I325421,I2507,I325059,I325024,);
DFFARX1 I_18995 (I325413,I2507,I325059,I325042,);
nor I_18996 (I325466,I90717,I90696);
not I_18997 (I325483,I325466);
nor I_18998 (I325045,I325322,I325483);
nand I_18999 (I325030,I325339,I325483);
nor I_19000 (I325039,I325085,I325466);
DFFARX1 I_19001 (I325466,I2507,I325059,I325048,);
not I_19002 (I325586,I2514);
DFFARX1 I_19003 (I387035,I2507,I325586,I325612,);
nand I_19004 (I325620,I387047,I387026);
and I_19005 (I325637,I325620,I387050);
DFFARX1 I_19006 (I325637,I2507,I325586,I325663,);
nor I_19007 (I325554,I325663,I325612);
not I_19008 (I325685,I325663);
DFFARX1 I_19009 (I387041,I2507,I325586,I325711,);
nand I_19010 (I325719,I325711,I387023);
not I_19011 (I325736,I325719);
DFFARX1 I_19012 (I325736,I2507,I325586,I325762,);
not I_19013 (I325578,I325762);
nor I_19014 (I325784,I325612,I325719);
nor I_19015 (I325560,I325663,I325784);
DFFARX1 I_19016 (I387038,I2507,I325586,I325824,);
DFFARX1 I_19017 (I325824,I2507,I325586,I325841,);
not I_19018 (I325849,I325841);
not I_19019 (I325866,I325824);
nand I_19020 (I325563,I325866,I325685);
nand I_19021 (I325897,I387023,I387029);
and I_19022 (I325914,I325897,I387032);
DFFARX1 I_19023 (I325914,I2507,I325586,I325940,);
nor I_19024 (I325948,I325940,I325612);
DFFARX1 I_19025 (I325948,I2507,I325586,I325551,);
DFFARX1 I_19026 (I325940,I2507,I325586,I325569,);
nor I_19027 (I325993,I387044,I387029);
not I_19028 (I326010,I325993);
nor I_19029 (I325572,I325849,I326010);
nand I_19030 (I325557,I325866,I326010);
nor I_19031 (I325566,I325612,I325993);
DFFARX1 I_19032 (I325993,I2507,I325586,I325575,);
not I_19033 (I326113,I2514);
DFFARX1 I_19034 (I1165300,I2507,I326113,I326139,);
nand I_19035 (I326147,I1165315,I1165300);
and I_19036 (I326164,I326147,I1165318);
DFFARX1 I_19037 (I326164,I2507,I326113,I326190,);
nor I_19038 (I326081,I326190,I326139);
not I_19039 (I326212,I326190);
DFFARX1 I_19040 (I1165324,I2507,I326113,I326238,);
nand I_19041 (I326246,I326238,I1165306);
not I_19042 (I326263,I326246);
DFFARX1 I_19043 (I326263,I2507,I326113,I326289,);
not I_19044 (I326105,I326289);
nor I_19045 (I326311,I326139,I326246);
nor I_19046 (I326087,I326190,I326311);
DFFARX1 I_19047 (I1165303,I2507,I326113,I326351,);
DFFARX1 I_19048 (I326351,I2507,I326113,I326368,);
not I_19049 (I326376,I326368);
not I_19050 (I326393,I326351);
nand I_19051 (I326090,I326393,I326212);
nand I_19052 (I326424,I1165303,I1165309);
and I_19053 (I326441,I326424,I1165321);
DFFARX1 I_19054 (I326441,I2507,I326113,I326467,);
nor I_19055 (I326475,I326467,I326139);
DFFARX1 I_19056 (I326475,I2507,I326113,I326078,);
DFFARX1 I_19057 (I326467,I2507,I326113,I326096,);
nor I_19058 (I326520,I1165312,I1165309);
not I_19059 (I326537,I326520);
nor I_19060 (I326099,I326376,I326537);
nand I_19061 (I326084,I326393,I326537);
nor I_19062 (I326093,I326139,I326520);
DFFARX1 I_19063 (I326520,I2507,I326113,I326102,);
not I_19064 (I326640,I2514);
DFFARX1 I_19065 (I627262,I2507,I326640,I326666,);
nand I_19066 (I326674,I627253,I627268);
and I_19067 (I326691,I326674,I627274);
DFFARX1 I_19068 (I326691,I2507,I326640,I326717,);
nor I_19069 (I326608,I326717,I326666);
not I_19070 (I326739,I326717);
DFFARX1 I_19071 (I627259,I2507,I326640,I326765,);
nand I_19072 (I326773,I326765,I627253);
not I_19073 (I326790,I326773);
DFFARX1 I_19074 (I326790,I2507,I326640,I326816,);
not I_19075 (I326632,I326816);
nor I_19076 (I326838,I326666,I326773);
nor I_19077 (I326614,I326717,I326838);
DFFARX1 I_19078 (I627256,I2507,I326640,I326878,);
DFFARX1 I_19079 (I326878,I2507,I326640,I326895,);
not I_19080 (I326903,I326895);
not I_19081 (I326920,I326878);
nand I_19082 (I326617,I326920,I326739);
nand I_19083 (I326951,I627250,I627265);
and I_19084 (I326968,I326951,I627250);
DFFARX1 I_19085 (I326968,I2507,I326640,I326994,);
nor I_19086 (I327002,I326994,I326666);
DFFARX1 I_19087 (I327002,I2507,I326640,I326605,);
DFFARX1 I_19088 (I326994,I2507,I326640,I326623,);
nor I_19089 (I327047,I627271,I627265);
not I_19090 (I327064,I327047);
nor I_19091 (I326626,I326903,I327064);
nand I_19092 (I326611,I326920,I327064);
nor I_19093 (I326620,I326666,I327047);
DFFARX1 I_19094 (I327047,I2507,I326640,I326629,);
not I_19095 (I327167,I2514);
DFFARX1 I_19096 (I222225,I2507,I327167,I327193,);
nand I_19097 (I327201,I222225,I222231);
and I_19098 (I327218,I327201,I222249);
DFFARX1 I_19099 (I327218,I2507,I327167,I327244,);
nor I_19100 (I327135,I327244,I327193);
not I_19101 (I327266,I327244);
DFFARX1 I_19102 (I222237,I2507,I327167,I327292,);
nand I_19103 (I327300,I327292,I222234);
not I_19104 (I327317,I327300);
DFFARX1 I_19105 (I327317,I2507,I327167,I327343,);
not I_19106 (I327159,I327343);
nor I_19107 (I327365,I327193,I327300);
nor I_19108 (I327141,I327244,I327365);
DFFARX1 I_19109 (I222243,I2507,I327167,I327405,);
DFFARX1 I_19110 (I327405,I2507,I327167,I327422,);
not I_19111 (I327430,I327422);
not I_19112 (I327447,I327405);
nand I_19113 (I327144,I327447,I327266);
nand I_19114 (I327478,I222228,I222228);
and I_19115 (I327495,I327478,I222240);
DFFARX1 I_19116 (I327495,I2507,I327167,I327521,);
nor I_19117 (I327529,I327521,I327193);
DFFARX1 I_19118 (I327529,I2507,I327167,I327132,);
DFFARX1 I_19119 (I327521,I2507,I327167,I327150,);
nor I_19120 (I327574,I222246,I222228);
not I_19121 (I327591,I327574);
nor I_19122 (I327153,I327430,I327591);
nand I_19123 (I327138,I327447,I327591);
nor I_19124 (I327147,I327193,I327574);
DFFARX1 I_19125 (I327574,I2507,I327167,I327156,);
not I_19126 (I327694,I2514);
DFFARX1 I_19127 (I1313068,I2507,I327694,I327720,);
nand I_19128 (I327728,I1313047,I1313047);
and I_19129 (I327745,I327728,I1313074);
DFFARX1 I_19130 (I327745,I2507,I327694,I327771,);
nor I_19131 (I327662,I327771,I327720);
not I_19132 (I327793,I327771);
DFFARX1 I_19133 (I1313062,I2507,I327694,I327819,);
nand I_19134 (I327827,I327819,I1313065);
not I_19135 (I327844,I327827);
DFFARX1 I_19136 (I327844,I2507,I327694,I327870,);
not I_19137 (I327686,I327870);
nor I_19138 (I327892,I327720,I327827);
nor I_19139 (I327668,I327771,I327892);
DFFARX1 I_19140 (I1313056,I2507,I327694,I327932,);
DFFARX1 I_19141 (I327932,I2507,I327694,I327949,);
not I_19142 (I327957,I327949);
not I_19143 (I327974,I327932);
nand I_19144 (I327671,I327974,I327793);
nand I_19145 (I328005,I1313053,I1313050);
and I_19146 (I328022,I328005,I1313071);
DFFARX1 I_19147 (I328022,I2507,I327694,I328048,);
nor I_19148 (I328056,I328048,I327720);
DFFARX1 I_19149 (I328056,I2507,I327694,I327659,);
DFFARX1 I_19150 (I328048,I2507,I327694,I327677,);
nor I_19151 (I328101,I1313059,I1313050);
not I_19152 (I328118,I328101);
nor I_19153 (I327680,I327957,I328118);
nand I_19154 (I327665,I327974,I328118);
nor I_19155 (I327674,I327720,I328101);
DFFARX1 I_19156 (I328101,I2507,I327694,I327683,);
not I_19157 (I328221,I2514);
DFFARX1 I_19158 (I657318,I2507,I328221,I328247,);
nand I_19159 (I328255,I657309,I657324);
and I_19160 (I328272,I328255,I657330);
DFFARX1 I_19161 (I328272,I2507,I328221,I328298,);
nor I_19162 (I328189,I328298,I328247);
not I_19163 (I328320,I328298);
DFFARX1 I_19164 (I657315,I2507,I328221,I328346,);
nand I_19165 (I328354,I328346,I657309);
not I_19166 (I328371,I328354);
DFFARX1 I_19167 (I328371,I2507,I328221,I328397,);
not I_19168 (I328213,I328397);
nor I_19169 (I328419,I328247,I328354);
nor I_19170 (I328195,I328298,I328419);
DFFARX1 I_19171 (I657312,I2507,I328221,I328459,);
DFFARX1 I_19172 (I328459,I2507,I328221,I328476,);
not I_19173 (I328484,I328476);
not I_19174 (I328501,I328459);
nand I_19175 (I328198,I328501,I328320);
nand I_19176 (I328532,I657306,I657321);
and I_19177 (I328549,I328532,I657306);
DFFARX1 I_19178 (I328549,I2507,I328221,I328575,);
nor I_19179 (I328583,I328575,I328247);
DFFARX1 I_19180 (I328583,I2507,I328221,I328186,);
DFFARX1 I_19181 (I328575,I2507,I328221,I328204,);
nor I_19182 (I328628,I657327,I657321);
not I_19183 (I328645,I328628);
nor I_19184 (I328207,I328484,I328645);
nand I_19185 (I328192,I328501,I328645);
nor I_19186 (I328201,I328247,I328628);
DFFARX1 I_19187 (I328628,I2507,I328221,I328210,);
not I_19188 (I328748,I2514);
DFFARX1 I_19189 (I102293,I2507,I328748,I328774,);
nand I_19190 (I328782,I102305,I102314);
and I_19191 (I328799,I328782,I102293);
DFFARX1 I_19192 (I328799,I2507,I328748,I328825,);
nor I_19193 (I328716,I328825,I328774);
not I_19194 (I328847,I328825);
DFFARX1 I_19195 (I102308,I2507,I328748,I328873,);
nand I_19196 (I328881,I328873,I102296);
not I_19197 (I328898,I328881);
DFFARX1 I_19198 (I328898,I2507,I328748,I328924,);
not I_19199 (I328740,I328924);
nor I_19200 (I328946,I328774,I328881);
nor I_19201 (I328722,I328825,I328946);
DFFARX1 I_19202 (I102299,I2507,I328748,I328986,);
DFFARX1 I_19203 (I328986,I2507,I328748,I329003,);
not I_19204 (I329011,I329003);
not I_19205 (I329028,I328986);
nand I_19206 (I328725,I329028,I328847);
nand I_19207 (I329059,I102290,I102290);
and I_19208 (I329076,I329059,I102302);
DFFARX1 I_19209 (I329076,I2507,I328748,I329102,);
nor I_19210 (I329110,I329102,I328774);
DFFARX1 I_19211 (I329110,I2507,I328748,I328713,);
DFFARX1 I_19212 (I329102,I2507,I328748,I328731,);
nor I_19213 (I329155,I102311,I102290);
not I_19214 (I329172,I329155);
nor I_19215 (I328734,I329011,I329172);
nand I_19216 (I328719,I329028,I329172);
nor I_19217 (I328728,I328774,I329155);
DFFARX1 I_19218 (I329155,I2507,I328748,I328737,);
not I_19219 (I329275,I2514);
DFFARX1 I_19220 (I52228,I2507,I329275,I329301,);
nand I_19221 (I329309,I52240,I52249);
and I_19222 (I329326,I329309,I52228);
DFFARX1 I_19223 (I329326,I2507,I329275,I329352,);
nor I_19224 (I329243,I329352,I329301);
not I_19225 (I329374,I329352);
DFFARX1 I_19226 (I52243,I2507,I329275,I329400,);
nand I_19227 (I329408,I329400,I52231);
not I_19228 (I329425,I329408);
DFFARX1 I_19229 (I329425,I2507,I329275,I329451,);
not I_19230 (I329267,I329451);
nor I_19231 (I329473,I329301,I329408);
nor I_19232 (I329249,I329352,I329473);
DFFARX1 I_19233 (I52234,I2507,I329275,I329513,);
DFFARX1 I_19234 (I329513,I2507,I329275,I329530,);
not I_19235 (I329538,I329530);
not I_19236 (I329555,I329513);
nand I_19237 (I329252,I329555,I329374);
nand I_19238 (I329586,I52225,I52225);
and I_19239 (I329603,I329586,I52237);
DFFARX1 I_19240 (I329603,I2507,I329275,I329629,);
nor I_19241 (I329637,I329629,I329301);
DFFARX1 I_19242 (I329637,I2507,I329275,I329240,);
DFFARX1 I_19243 (I329629,I2507,I329275,I329258,);
nor I_19244 (I329682,I52246,I52225);
not I_19245 (I329699,I329682);
nor I_19246 (I329261,I329538,I329699);
nand I_19247 (I329246,I329555,I329699);
nor I_19248 (I329255,I329301,I329682);
DFFARX1 I_19249 (I329682,I2507,I329275,I329264,);
not I_19250 (I329802,I2514);
DFFARX1 I_19251 (I1007730,I2507,I329802,I329828,);
nand I_19252 (I329836,I1007727,I1007745);
and I_19253 (I329853,I329836,I1007736);
DFFARX1 I_19254 (I329853,I2507,I329802,I329879,);
nor I_19255 (I329770,I329879,I329828);
not I_19256 (I329901,I329879);
DFFARX1 I_19257 (I1007751,I2507,I329802,I329927,);
nand I_19258 (I329935,I329927,I1007733);
not I_19259 (I329952,I329935);
DFFARX1 I_19260 (I329952,I2507,I329802,I329978,);
not I_19261 (I329794,I329978);
nor I_19262 (I330000,I329828,I329935);
nor I_19263 (I329776,I329879,I330000);
DFFARX1 I_19264 (I1007739,I2507,I329802,I330040,);
DFFARX1 I_19265 (I330040,I2507,I329802,I330057,);
not I_19266 (I330065,I330057);
not I_19267 (I330082,I330040);
nand I_19268 (I329779,I330082,I329901);
nand I_19269 (I330113,I1007727,I1007754);
and I_19270 (I330130,I330113,I1007742);
DFFARX1 I_19271 (I330130,I2507,I329802,I330156,);
nor I_19272 (I330164,I330156,I329828);
DFFARX1 I_19273 (I330164,I2507,I329802,I329767,);
DFFARX1 I_19274 (I330156,I2507,I329802,I329785,);
nor I_19275 (I330209,I1007748,I1007754);
not I_19276 (I330226,I330209);
nor I_19277 (I329788,I330065,I330226);
nand I_19278 (I329773,I330082,I330226);
nor I_19279 (I329782,I329828,I330209);
DFFARX1 I_19280 (I330209,I2507,I329802,I329791,);
not I_19281 (I330329,I2514);
DFFARX1 I_19282 (I1206356,I2507,I330329,I330355,);
nand I_19283 (I330363,I1206338,I1206362);
and I_19284 (I330380,I330363,I1206353);
DFFARX1 I_19285 (I330380,I2507,I330329,I330406,);
nor I_19286 (I330297,I330406,I330355);
not I_19287 (I330428,I330406);
DFFARX1 I_19288 (I1206359,I2507,I330329,I330454,);
nand I_19289 (I330462,I330454,I1206347);
not I_19290 (I330479,I330462);
DFFARX1 I_19291 (I330479,I2507,I330329,I330505,);
not I_19292 (I330321,I330505);
nor I_19293 (I330527,I330355,I330462);
nor I_19294 (I330303,I330406,I330527);
DFFARX1 I_19295 (I1206338,I2507,I330329,I330567,);
DFFARX1 I_19296 (I330567,I2507,I330329,I330584,);
not I_19297 (I330592,I330584);
not I_19298 (I330609,I330567);
nand I_19299 (I330306,I330609,I330428);
nand I_19300 (I330640,I1206344,I1206341);
and I_19301 (I330657,I330640,I1206350);
DFFARX1 I_19302 (I330657,I2507,I330329,I330683,);
nor I_19303 (I330691,I330683,I330355);
DFFARX1 I_19304 (I330691,I2507,I330329,I330294,);
DFFARX1 I_19305 (I330683,I2507,I330329,I330312,);
nor I_19306 (I330736,I1206341,I1206341);
not I_19307 (I330753,I330736);
nor I_19308 (I330315,I330592,I330753);
nand I_19309 (I330300,I330609,I330753);
nor I_19310 (I330309,I330355,I330736);
DFFARX1 I_19311 (I330736,I2507,I330329,I330318,);
not I_19312 (I330856,I2514);
DFFARX1 I_19313 (I394107,I2507,I330856,I330882,);
nand I_19314 (I330890,I394119,I394098);
and I_19315 (I330907,I330890,I394122);
DFFARX1 I_19316 (I330907,I2507,I330856,I330933,);
nor I_19317 (I330824,I330933,I330882);
not I_19318 (I330955,I330933);
DFFARX1 I_19319 (I394113,I2507,I330856,I330981,);
nand I_19320 (I330989,I330981,I394095);
not I_19321 (I331006,I330989);
DFFARX1 I_19322 (I331006,I2507,I330856,I331032,);
not I_19323 (I330848,I331032);
nor I_19324 (I331054,I330882,I330989);
nor I_19325 (I330830,I330933,I331054);
DFFARX1 I_19326 (I394110,I2507,I330856,I331094,);
DFFARX1 I_19327 (I331094,I2507,I330856,I331111,);
not I_19328 (I331119,I331111);
not I_19329 (I331136,I331094);
nand I_19330 (I330833,I331136,I330955);
nand I_19331 (I331167,I394095,I394101);
and I_19332 (I331184,I331167,I394104);
DFFARX1 I_19333 (I331184,I2507,I330856,I331210,);
nor I_19334 (I331218,I331210,I330882);
DFFARX1 I_19335 (I331218,I2507,I330856,I330821,);
DFFARX1 I_19336 (I331210,I2507,I330856,I330839,);
nor I_19337 (I331263,I394116,I394101);
not I_19338 (I331280,I331263);
nor I_19339 (I330842,I331119,I331280);
nand I_19340 (I330827,I331136,I331280);
nor I_19341 (I330836,I330882,I331263);
DFFARX1 I_19342 (I331263,I2507,I330856,I330845,);
not I_19343 (I331383,I2514);
DFFARX1 I_19344 (I1072820,I2507,I331383,I331409,);
nand I_19345 (I331417,I1072835,I1072820);
and I_19346 (I331434,I331417,I1072838);
DFFARX1 I_19347 (I331434,I2507,I331383,I331460,);
nor I_19348 (I331351,I331460,I331409);
not I_19349 (I331482,I331460);
DFFARX1 I_19350 (I1072844,I2507,I331383,I331508,);
nand I_19351 (I331516,I331508,I1072826);
not I_19352 (I331533,I331516);
DFFARX1 I_19353 (I331533,I2507,I331383,I331559,);
not I_19354 (I331375,I331559);
nor I_19355 (I331581,I331409,I331516);
nor I_19356 (I331357,I331460,I331581);
DFFARX1 I_19357 (I1072823,I2507,I331383,I331621,);
DFFARX1 I_19358 (I331621,I2507,I331383,I331638,);
not I_19359 (I331646,I331638);
not I_19360 (I331663,I331621);
nand I_19361 (I331360,I331663,I331482);
nand I_19362 (I331694,I1072823,I1072829);
and I_19363 (I331711,I331694,I1072841);
DFFARX1 I_19364 (I331711,I2507,I331383,I331737,);
nor I_19365 (I331745,I331737,I331409);
DFFARX1 I_19366 (I331745,I2507,I331383,I331348,);
DFFARX1 I_19367 (I331737,I2507,I331383,I331366,);
nor I_19368 (I331790,I1072832,I1072829);
not I_19369 (I331807,I331790);
nor I_19370 (I331369,I331646,I331807);
nand I_19371 (I331354,I331663,I331807);
nor I_19372 (I331363,I331409,I331790);
DFFARX1 I_19373 (I331790,I2507,I331383,I331372,);
not I_19374 (I331910,I2514);
DFFARX1 I_19375 (I735926,I2507,I331910,I331936,);
nand I_19376 (I331944,I735917,I735932);
and I_19377 (I331961,I331944,I735938);
DFFARX1 I_19378 (I331961,I2507,I331910,I331987,);
nor I_19379 (I331878,I331987,I331936);
not I_19380 (I332009,I331987);
DFFARX1 I_19381 (I735923,I2507,I331910,I332035,);
nand I_19382 (I332043,I332035,I735917);
not I_19383 (I332060,I332043);
DFFARX1 I_19384 (I332060,I2507,I331910,I332086,);
not I_19385 (I331902,I332086);
nor I_19386 (I332108,I331936,I332043);
nor I_19387 (I331884,I331987,I332108);
DFFARX1 I_19388 (I735920,I2507,I331910,I332148,);
DFFARX1 I_19389 (I332148,I2507,I331910,I332165,);
not I_19390 (I332173,I332165);
not I_19391 (I332190,I332148);
nand I_19392 (I331887,I332190,I332009);
nand I_19393 (I332221,I735914,I735929);
and I_19394 (I332238,I332221,I735914);
DFFARX1 I_19395 (I332238,I2507,I331910,I332264,);
nor I_19396 (I332272,I332264,I331936);
DFFARX1 I_19397 (I332272,I2507,I331910,I331875,);
DFFARX1 I_19398 (I332264,I2507,I331910,I331893,);
nor I_19399 (I332317,I735935,I735929);
not I_19400 (I332334,I332317);
nor I_19401 (I331896,I332173,I332334);
nand I_19402 (I331881,I332190,I332334);
nor I_19403 (I331890,I331936,I332317);
DFFARX1 I_19404 (I332317,I2507,I331910,I331899,);
not I_19405 (I332437,I2514);
DFFARX1 I_19406 (I212705,I2507,I332437,I332463,);
nand I_19407 (I332471,I212705,I212711);
and I_19408 (I332488,I332471,I212729);
DFFARX1 I_19409 (I332488,I2507,I332437,I332514,);
nor I_19410 (I332405,I332514,I332463);
not I_19411 (I332536,I332514);
DFFARX1 I_19412 (I212717,I2507,I332437,I332562,);
nand I_19413 (I332570,I332562,I212714);
not I_19414 (I332587,I332570);
DFFARX1 I_19415 (I332587,I2507,I332437,I332613,);
not I_19416 (I332429,I332613);
nor I_19417 (I332635,I332463,I332570);
nor I_19418 (I332411,I332514,I332635);
DFFARX1 I_19419 (I212723,I2507,I332437,I332675,);
DFFARX1 I_19420 (I332675,I2507,I332437,I332692,);
not I_19421 (I332700,I332692);
not I_19422 (I332717,I332675);
nand I_19423 (I332414,I332717,I332536);
nand I_19424 (I332748,I212708,I212708);
and I_19425 (I332765,I332748,I212720);
DFFARX1 I_19426 (I332765,I2507,I332437,I332791,);
nor I_19427 (I332799,I332791,I332463);
DFFARX1 I_19428 (I332799,I2507,I332437,I332402,);
DFFARX1 I_19429 (I332791,I2507,I332437,I332420,);
nor I_19430 (I332844,I212726,I212708);
not I_19431 (I332861,I332844);
nor I_19432 (I332423,I332700,I332861);
nand I_19433 (I332408,I332717,I332861);
nor I_19434 (I332417,I332463,I332844);
DFFARX1 I_19435 (I332844,I2507,I332437,I332426,);
not I_19436 (I332964,I2514);
DFFARX1 I_19437 (I38523,I2507,I332964,I332990,);
nand I_19438 (I332998,I38547,I38526);
and I_19439 (I333015,I332998,I38523);
DFFARX1 I_19440 (I333015,I2507,I332964,I333041,);
nor I_19441 (I332932,I333041,I332990);
not I_19442 (I333063,I333041);
DFFARX1 I_19443 (I38529,I2507,I332964,I333089,);
nand I_19444 (I333097,I333089,I38538);
not I_19445 (I333114,I333097);
DFFARX1 I_19446 (I333114,I2507,I332964,I333140,);
not I_19447 (I332956,I333140);
nor I_19448 (I333162,I332990,I333097);
nor I_19449 (I332938,I333041,I333162);
DFFARX1 I_19450 (I38532,I2507,I332964,I333202,);
DFFARX1 I_19451 (I333202,I2507,I332964,I333219,);
not I_19452 (I333227,I333219);
not I_19453 (I333244,I333202);
nand I_19454 (I332941,I333244,I333063);
nand I_19455 (I333275,I38544,I38526);
and I_19456 (I333292,I333275,I38535);
DFFARX1 I_19457 (I333292,I2507,I332964,I333318,);
nor I_19458 (I333326,I333318,I332990);
DFFARX1 I_19459 (I333326,I2507,I332964,I332929,);
DFFARX1 I_19460 (I333318,I2507,I332964,I332947,);
nor I_19461 (I333371,I38541,I38526);
not I_19462 (I333388,I333371);
nor I_19463 (I332950,I333227,I333388);
nand I_19464 (I332935,I333244,I333388);
nor I_19465 (I332944,I332990,I333371);
DFFARX1 I_19466 (I333371,I2507,I332964,I332953,);
not I_19467 (I333491,I2514);
DFFARX1 I_19468 (I196045,I2507,I333491,I333517,);
nand I_19469 (I333525,I196045,I196051);
and I_19470 (I333542,I333525,I196069);
DFFARX1 I_19471 (I333542,I2507,I333491,I333568,);
nor I_19472 (I333459,I333568,I333517);
not I_19473 (I333590,I333568);
DFFARX1 I_19474 (I196057,I2507,I333491,I333616,);
nand I_19475 (I333624,I333616,I196054);
not I_19476 (I333641,I333624);
DFFARX1 I_19477 (I333641,I2507,I333491,I333667,);
not I_19478 (I333483,I333667);
nor I_19479 (I333689,I333517,I333624);
nor I_19480 (I333465,I333568,I333689);
DFFARX1 I_19481 (I196063,I2507,I333491,I333729,);
DFFARX1 I_19482 (I333729,I2507,I333491,I333746,);
not I_19483 (I333754,I333746);
not I_19484 (I333771,I333729);
nand I_19485 (I333468,I333771,I333590);
nand I_19486 (I333802,I196048,I196048);
and I_19487 (I333819,I333802,I196060);
DFFARX1 I_19488 (I333819,I2507,I333491,I333845,);
nor I_19489 (I333853,I333845,I333517);
DFFARX1 I_19490 (I333853,I2507,I333491,I333456,);
DFFARX1 I_19491 (I333845,I2507,I333491,I333474,);
nor I_19492 (I333898,I196066,I196048);
not I_19493 (I333915,I333898);
nor I_19494 (I333477,I333754,I333915);
nand I_19495 (I333462,I333771,I333915);
nor I_19496 (I333471,I333517,I333898);
DFFARX1 I_19497 (I333898,I2507,I333491,I333480,);
not I_19498 (I334018,I2514);
DFFARX1 I_19499 (I861802,I2507,I334018,I334044,);
nand I_19500 (I334052,I861805,I861799);
and I_19501 (I334069,I334052,I861811);
DFFARX1 I_19502 (I334069,I2507,I334018,I334095,);
nor I_19503 (I333986,I334095,I334044);
not I_19504 (I334117,I334095);
DFFARX1 I_19505 (I861814,I2507,I334018,I334143,);
nand I_19506 (I334151,I334143,I861805);
not I_19507 (I334168,I334151);
DFFARX1 I_19508 (I334168,I2507,I334018,I334194,);
not I_19509 (I334010,I334194);
nor I_19510 (I334216,I334044,I334151);
nor I_19511 (I333992,I334095,I334216);
DFFARX1 I_19512 (I861817,I2507,I334018,I334256,);
DFFARX1 I_19513 (I334256,I2507,I334018,I334273,);
not I_19514 (I334281,I334273);
not I_19515 (I334298,I334256);
nand I_19516 (I333995,I334298,I334117);
nand I_19517 (I334329,I861799,I861808);
and I_19518 (I334346,I334329,I861802);
DFFARX1 I_19519 (I334346,I2507,I334018,I334372,);
nor I_19520 (I334380,I334372,I334044);
DFFARX1 I_19521 (I334380,I2507,I334018,I333983,);
DFFARX1 I_19522 (I334372,I2507,I334018,I334001,);
nor I_19523 (I334425,I861820,I861808);
not I_19524 (I334442,I334425);
nor I_19525 (I334004,I334281,I334442);
nand I_19526 (I333989,I334298,I334442);
nor I_19527 (I333998,I334044,I334425);
DFFARX1 I_19528 (I334425,I2507,I334018,I334007,);
not I_19529 (I334545,I2514);
DFFARX1 I_19530 (I452315,I2507,I334545,I334571,);
nand I_19531 (I334579,I452327,I452306);
and I_19532 (I334596,I334579,I452330);
DFFARX1 I_19533 (I334596,I2507,I334545,I334622,);
nor I_19534 (I334513,I334622,I334571);
not I_19535 (I334644,I334622);
DFFARX1 I_19536 (I452321,I2507,I334545,I334670,);
nand I_19537 (I334678,I334670,I452303);
not I_19538 (I334695,I334678);
DFFARX1 I_19539 (I334695,I2507,I334545,I334721,);
not I_19540 (I334537,I334721);
nor I_19541 (I334743,I334571,I334678);
nor I_19542 (I334519,I334622,I334743);
DFFARX1 I_19543 (I452318,I2507,I334545,I334783,);
DFFARX1 I_19544 (I334783,I2507,I334545,I334800,);
not I_19545 (I334808,I334800);
not I_19546 (I334825,I334783);
nand I_19547 (I334522,I334825,I334644);
nand I_19548 (I334856,I452303,I452309);
and I_19549 (I334873,I334856,I452312);
DFFARX1 I_19550 (I334873,I2507,I334545,I334899,);
nor I_19551 (I334907,I334899,I334571);
DFFARX1 I_19552 (I334907,I2507,I334545,I334510,);
DFFARX1 I_19553 (I334899,I2507,I334545,I334528,);
nor I_19554 (I334952,I452324,I452309);
not I_19555 (I334969,I334952);
nor I_19556 (I334531,I334808,I334969);
nand I_19557 (I334516,I334825,I334969);
nor I_19558 (I334525,I334571,I334952);
DFFARX1 I_19559 (I334952,I2507,I334545,I334534,);
not I_19560 (I335072,I2514);
DFFARX1 I_19561 (I915352,I2507,I335072,I335098,);
nand I_19562 (I335106,I915349,I915367);
and I_19563 (I335123,I335106,I915358);
DFFARX1 I_19564 (I335123,I2507,I335072,I335149,);
nor I_19565 (I335040,I335149,I335098);
not I_19566 (I335171,I335149);
DFFARX1 I_19567 (I915373,I2507,I335072,I335197,);
nand I_19568 (I335205,I335197,I915355);
not I_19569 (I335222,I335205);
DFFARX1 I_19570 (I335222,I2507,I335072,I335248,);
not I_19571 (I335064,I335248);
nor I_19572 (I335270,I335098,I335205);
nor I_19573 (I335046,I335149,I335270);
DFFARX1 I_19574 (I915361,I2507,I335072,I335310,);
DFFARX1 I_19575 (I335310,I2507,I335072,I335327,);
not I_19576 (I335335,I335327);
not I_19577 (I335352,I335310);
nand I_19578 (I335049,I335352,I335171);
nand I_19579 (I335383,I915349,I915376);
and I_19580 (I335400,I335383,I915364);
DFFARX1 I_19581 (I335400,I2507,I335072,I335426,);
nor I_19582 (I335434,I335426,I335098);
DFFARX1 I_19583 (I335434,I2507,I335072,I335037,);
DFFARX1 I_19584 (I335426,I2507,I335072,I335055,);
nor I_19585 (I335479,I915370,I915376);
not I_19586 (I335496,I335479);
nor I_19587 (I335058,I335335,I335496);
nand I_19588 (I335043,I335352,I335496);
nor I_19589 (I335052,I335098,I335479);
DFFARX1 I_19590 (I335479,I2507,I335072,I335061,);
not I_19591 (I335599,I2514);
DFFARX1 I_19592 (I1056146,I2507,I335599,I335625,);
nand I_19593 (I335633,I1056143,I1056146);
and I_19594 (I335650,I335633,I1056155);
DFFARX1 I_19595 (I335650,I2507,I335599,I335676,);
nor I_19596 (I335567,I335676,I335625);
not I_19597 (I335698,I335676);
DFFARX1 I_19598 (I1056143,I2507,I335599,I335724,);
nand I_19599 (I335732,I335724,I1056161);
not I_19600 (I335749,I335732);
DFFARX1 I_19601 (I335749,I2507,I335599,I335775,);
not I_19602 (I335591,I335775);
nor I_19603 (I335797,I335625,I335732);
nor I_19604 (I335573,I335676,I335797);
DFFARX1 I_19605 (I1056149,I2507,I335599,I335837,);
DFFARX1 I_19606 (I335837,I2507,I335599,I335854,);
not I_19607 (I335862,I335854);
not I_19608 (I335879,I335837);
nand I_19609 (I335576,I335879,I335698);
nand I_19610 (I335910,I1056158,I1056164);
and I_19611 (I335927,I335910,I1056149);
DFFARX1 I_19612 (I335927,I2507,I335599,I335953,);
nor I_19613 (I335961,I335953,I335625);
DFFARX1 I_19614 (I335961,I2507,I335599,I335564,);
DFFARX1 I_19615 (I335953,I2507,I335599,I335582,);
nor I_19616 (I336006,I1056152,I1056164);
not I_19617 (I336023,I336006);
nor I_19618 (I335585,I335862,I336023);
nand I_19619 (I335570,I335879,I336023);
nor I_19620 (I335579,I335625,I336006);
DFFARX1 I_19621 (I336006,I2507,I335599,I335588,);
not I_19622 (I336126,I2514);
DFFARX1 I_19623 (I909538,I2507,I336126,I336152,);
nand I_19624 (I336160,I909535,I909553);
and I_19625 (I336177,I336160,I909544);
DFFARX1 I_19626 (I336177,I2507,I336126,I336203,);
nor I_19627 (I336094,I336203,I336152);
not I_19628 (I336225,I336203);
DFFARX1 I_19629 (I909559,I2507,I336126,I336251,);
nand I_19630 (I336259,I336251,I909541);
not I_19631 (I336276,I336259);
DFFARX1 I_19632 (I336276,I2507,I336126,I336302,);
not I_19633 (I336118,I336302);
nor I_19634 (I336324,I336152,I336259);
nor I_19635 (I336100,I336203,I336324);
DFFARX1 I_19636 (I909547,I2507,I336126,I336364,);
DFFARX1 I_19637 (I336364,I2507,I336126,I336381,);
not I_19638 (I336389,I336381);
not I_19639 (I336406,I336364);
nand I_19640 (I336103,I336406,I336225);
nand I_19641 (I336437,I909535,I909562);
and I_19642 (I336454,I336437,I909550);
DFFARX1 I_19643 (I336454,I2507,I336126,I336480,);
nor I_19644 (I336488,I336480,I336152);
DFFARX1 I_19645 (I336488,I2507,I336126,I336091,);
DFFARX1 I_19646 (I336480,I2507,I336126,I336109,);
nor I_19647 (I336533,I909556,I909562);
not I_19648 (I336550,I336533);
nor I_19649 (I336112,I336389,I336550);
nand I_19650 (I336097,I336406,I336550);
nor I_19651 (I336106,I336152,I336533);
DFFARX1 I_19652 (I336533,I2507,I336126,I336115,);
not I_19653 (I336653,I2514);
DFFARX1 I_19654 (I1149694,I2507,I336653,I336679,);
nand I_19655 (I336687,I1149709,I1149694);
and I_19656 (I336704,I336687,I1149712);
DFFARX1 I_19657 (I336704,I2507,I336653,I336730,);
nor I_19658 (I336621,I336730,I336679);
not I_19659 (I336752,I336730);
DFFARX1 I_19660 (I1149718,I2507,I336653,I336778,);
nand I_19661 (I336786,I336778,I1149700);
not I_19662 (I336803,I336786);
DFFARX1 I_19663 (I336803,I2507,I336653,I336829,);
not I_19664 (I336645,I336829);
nor I_19665 (I336851,I336679,I336786);
nor I_19666 (I336627,I336730,I336851);
DFFARX1 I_19667 (I1149697,I2507,I336653,I336891,);
DFFARX1 I_19668 (I336891,I2507,I336653,I336908,);
not I_19669 (I336916,I336908);
not I_19670 (I336933,I336891);
nand I_19671 (I336630,I336933,I336752);
nand I_19672 (I336964,I1149697,I1149703);
and I_19673 (I336981,I336964,I1149715);
DFFARX1 I_19674 (I336981,I2507,I336653,I337007,);
nor I_19675 (I337015,I337007,I336679);
DFFARX1 I_19676 (I337015,I2507,I336653,I336618,);
DFFARX1 I_19677 (I337007,I2507,I336653,I336636,);
nor I_19678 (I337060,I1149706,I1149703);
not I_19679 (I337077,I337060);
nor I_19680 (I336639,I336916,I337077);
nand I_19681 (I336624,I336933,I337077);
nor I_19682 (I336633,I336679,I337060);
DFFARX1 I_19683 (I337060,I2507,I336653,I336642,);
not I_19684 (I337180,I2514);
DFFARX1 I_19685 (I1190154,I2507,I337180,I337206,);
nand I_19686 (I337214,I1190169,I1190154);
and I_19687 (I337231,I337214,I1190172);
DFFARX1 I_19688 (I337231,I2507,I337180,I337257,);
nor I_19689 (I337148,I337257,I337206);
not I_19690 (I337279,I337257);
DFFARX1 I_19691 (I1190178,I2507,I337180,I337305,);
nand I_19692 (I337313,I337305,I1190160);
not I_19693 (I337330,I337313);
DFFARX1 I_19694 (I337330,I2507,I337180,I337356,);
not I_19695 (I337172,I337356);
nor I_19696 (I337378,I337206,I337313);
nor I_19697 (I337154,I337257,I337378);
DFFARX1 I_19698 (I1190157,I2507,I337180,I337418,);
DFFARX1 I_19699 (I337418,I2507,I337180,I337435,);
not I_19700 (I337443,I337435);
not I_19701 (I337460,I337418);
nand I_19702 (I337157,I337460,I337279);
nand I_19703 (I337491,I1190157,I1190163);
and I_19704 (I337508,I337491,I1190175);
DFFARX1 I_19705 (I337508,I2507,I337180,I337534,);
nor I_19706 (I337542,I337534,I337206);
DFFARX1 I_19707 (I337542,I2507,I337180,I337145,);
DFFARX1 I_19708 (I337534,I2507,I337180,I337163,);
nor I_19709 (I337587,I1190166,I1190163);
not I_19710 (I337604,I337587);
nor I_19711 (I337166,I337443,I337604);
nand I_19712 (I337151,I337460,I337604);
nor I_19713 (I337160,I337206,I337587);
DFFARX1 I_19714 (I337587,I2507,I337180,I337169,);
not I_19715 (I337707,I2514);
DFFARX1 I_19716 (I508372,I2507,I337707,I337733,);
nand I_19717 (I337741,I508372,I508384);
and I_19718 (I337758,I337741,I508369);
DFFARX1 I_19719 (I337758,I2507,I337707,I337784,);
nor I_19720 (I337675,I337784,I337733);
not I_19721 (I337806,I337784);
DFFARX1 I_19722 (I508393,I2507,I337707,I337832,);
nand I_19723 (I337840,I337832,I508390);
not I_19724 (I337857,I337840);
DFFARX1 I_19725 (I337857,I2507,I337707,I337883,);
not I_19726 (I337699,I337883);
nor I_19727 (I337905,I337733,I337840);
nor I_19728 (I337681,I337784,I337905);
DFFARX1 I_19729 (I508381,I2507,I337707,I337945,);
DFFARX1 I_19730 (I337945,I2507,I337707,I337962,);
not I_19731 (I337970,I337962);
not I_19732 (I337987,I337945);
nand I_19733 (I337684,I337987,I337806);
nand I_19734 (I338018,I508369,I508378);
and I_19735 (I338035,I338018,I508387);
DFFARX1 I_19736 (I338035,I2507,I337707,I338061,);
nor I_19737 (I338069,I338061,I337733);
DFFARX1 I_19738 (I338069,I2507,I337707,I337672,);
DFFARX1 I_19739 (I338061,I2507,I337707,I337690,);
nor I_19740 (I338114,I508375,I508378);
not I_19741 (I338131,I338114);
nor I_19742 (I337693,I337970,I338131);
nand I_19743 (I337678,I337987,I338131);
nor I_19744 (I337687,I337733,I338114);
DFFARX1 I_19745 (I338114,I2507,I337707,I337696,);
not I_19746 (I338234,I2514);
DFFARX1 I_19747 (I1175126,I2507,I338234,I338260,);
nand I_19748 (I338268,I1175141,I1175126);
and I_19749 (I338285,I338268,I1175144);
DFFARX1 I_19750 (I338285,I2507,I338234,I338311,);
nor I_19751 (I338202,I338311,I338260);
not I_19752 (I338333,I338311);
DFFARX1 I_19753 (I1175150,I2507,I338234,I338359,);
nand I_19754 (I338367,I338359,I1175132);
not I_19755 (I338384,I338367);
DFFARX1 I_19756 (I338384,I2507,I338234,I338410,);
not I_19757 (I338226,I338410);
nor I_19758 (I338432,I338260,I338367);
nor I_19759 (I338208,I338311,I338432);
DFFARX1 I_19760 (I1175129,I2507,I338234,I338472,);
DFFARX1 I_19761 (I338472,I2507,I338234,I338489,);
not I_19762 (I338497,I338489);
not I_19763 (I338514,I338472);
nand I_19764 (I338211,I338514,I338333);
nand I_19765 (I338545,I1175129,I1175135);
and I_19766 (I338562,I338545,I1175147);
DFFARX1 I_19767 (I338562,I2507,I338234,I338588,);
nor I_19768 (I338596,I338588,I338260);
DFFARX1 I_19769 (I338596,I2507,I338234,I338199,);
DFFARX1 I_19770 (I338588,I2507,I338234,I338217,);
nor I_19771 (I338641,I1175138,I1175135);
not I_19772 (I338658,I338641);
nor I_19773 (I338220,I338497,I338658);
nand I_19774 (I338205,I338514,I338658);
nor I_19775 (I338214,I338260,I338641);
DFFARX1 I_19776 (I338641,I2507,I338234,I338223,);
not I_19777 (I338761,I2514);
DFFARX1 I_19778 (I573511,I2507,I338761,I338787,);
nand I_19779 (I338795,I573496,I573499);
and I_19780 (I338812,I338795,I573514);
DFFARX1 I_19781 (I338812,I2507,I338761,I338838,);
nor I_19782 (I338729,I338838,I338787);
not I_19783 (I338860,I338838);
DFFARX1 I_19784 (I573508,I2507,I338761,I338886,);
nand I_19785 (I338894,I338886,I573499);
not I_19786 (I338911,I338894);
DFFARX1 I_19787 (I338911,I2507,I338761,I338937,);
not I_19788 (I338753,I338937);
nor I_19789 (I338959,I338787,I338894);
nor I_19790 (I338735,I338838,I338959);
DFFARX1 I_19791 (I573505,I2507,I338761,I338999,);
DFFARX1 I_19792 (I338999,I2507,I338761,I339016,);
not I_19793 (I339024,I339016);
not I_19794 (I339041,I338999);
nand I_19795 (I338738,I339041,I338860);
nand I_19796 (I339072,I573520,I573496);
and I_19797 (I339089,I339072,I573517);
DFFARX1 I_19798 (I339089,I2507,I338761,I339115,);
nor I_19799 (I339123,I339115,I338787);
DFFARX1 I_19800 (I339123,I2507,I338761,I338726,);
DFFARX1 I_19801 (I339115,I2507,I338761,I338744,);
nor I_19802 (I339168,I573502,I573496);
not I_19803 (I339185,I339168);
nor I_19804 (I338747,I339024,I339185);
nand I_19805 (I338732,I339041,I339185);
nor I_19806 (I338741,I338787,I339168);
DFFARX1 I_19807 (I339168,I2507,I338761,I338750,);
not I_19808 (I339288,I2514);
DFFARX1 I_19809 (I1164144,I2507,I339288,I339314,);
nand I_19810 (I339322,I1164159,I1164144);
and I_19811 (I339339,I339322,I1164162);
DFFARX1 I_19812 (I339339,I2507,I339288,I339365,);
nor I_19813 (I339256,I339365,I339314);
not I_19814 (I339387,I339365);
DFFARX1 I_19815 (I1164168,I2507,I339288,I339413,);
nand I_19816 (I339421,I339413,I1164150);
not I_19817 (I339438,I339421);
DFFARX1 I_19818 (I339438,I2507,I339288,I339464,);
not I_19819 (I339280,I339464);
nor I_19820 (I339486,I339314,I339421);
nor I_19821 (I339262,I339365,I339486);
DFFARX1 I_19822 (I1164147,I2507,I339288,I339526,);
DFFARX1 I_19823 (I339526,I2507,I339288,I339543,);
not I_19824 (I339551,I339543);
not I_19825 (I339568,I339526);
nand I_19826 (I339265,I339568,I339387);
nand I_19827 (I339599,I1164147,I1164153);
and I_19828 (I339616,I339599,I1164165);
DFFARX1 I_19829 (I339616,I2507,I339288,I339642,);
nor I_19830 (I339650,I339642,I339314);
DFFARX1 I_19831 (I339650,I2507,I339288,I339253,);
DFFARX1 I_19832 (I339642,I2507,I339288,I339271,);
nor I_19833 (I339695,I1164156,I1164153);
not I_19834 (I339712,I339695);
nor I_19835 (I339274,I339551,I339712);
nand I_19836 (I339259,I339568,I339712);
nor I_19837 (I339268,I339314,I339695);
DFFARX1 I_19838 (I339695,I2507,I339288,I339277,);
not I_19839 (I339815,I2514);
DFFARX1 I_19840 (I1165878,I2507,I339815,I339841,);
nand I_19841 (I339849,I1165893,I1165878);
and I_19842 (I339866,I339849,I1165896);
DFFARX1 I_19843 (I339866,I2507,I339815,I339892,);
nor I_19844 (I339783,I339892,I339841);
not I_19845 (I339914,I339892);
DFFARX1 I_19846 (I1165902,I2507,I339815,I339940,);
nand I_19847 (I339948,I339940,I1165884);
not I_19848 (I339965,I339948);
DFFARX1 I_19849 (I339965,I2507,I339815,I339991,);
not I_19850 (I339807,I339991);
nor I_19851 (I340013,I339841,I339948);
nor I_19852 (I339789,I339892,I340013);
DFFARX1 I_19853 (I1165881,I2507,I339815,I340053,);
DFFARX1 I_19854 (I340053,I2507,I339815,I340070,);
not I_19855 (I340078,I340070);
not I_19856 (I340095,I340053);
nand I_19857 (I339792,I340095,I339914);
nand I_19858 (I340126,I1165881,I1165887);
and I_19859 (I340143,I340126,I1165899);
DFFARX1 I_19860 (I340143,I2507,I339815,I340169,);
nor I_19861 (I340177,I340169,I339841);
DFFARX1 I_19862 (I340177,I2507,I339815,I339780,);
DFFARX1 I_19863 (I340169,I2507,I339815,I339798,);
nor I_19864 (I340222,I1165890,I1165887);
not I_19865 (I340239,I340222);
nor I_19866 (I339801,I340078,I340239);
nand I_19867 (I339786,I340095,I340239);
nor I_19868 (I339795,I339841,I340222);
DFFARX1 I_19869 (I340222,I2507,I339815,I339804,);
not I_19870 (I340342,I2514);
DFFARX1 I_19871 (I739394,I2507,I340342,I340368,);
nand I_19872 (I340376,I739385,I739400);
and I_19873 (I340393,I340376,I739406);
DFFARX1 I_19874 (I340393,I2507,I340342,I340419,);
nor I_19875 (I340310,I340419,I340368);
not I_19876 (I340441,I340419);
DFFARX1 I_19877 (I739391,I2507,I340342,I340467,);
nand I_19878 (I340475,I340467,I739385);
not I_19879 (I340492,I340475);
DFFARX1 I_19880 (I340492,I2507,I340342,I340518,);
not I_19881 (I340334,I340518);
nor I_19882 (I340540,I340368,I340475);
nor I_19883 (I340316,I340419,I340540);
DFFARX1 I_19884 (I739388,I2507,I340342,I340580,);
DFFARX1 I_19885 (I340580,I2507,I340342,I340597,);
not I_19886 (I340605,I340597);
not I_19887 (I340622,I340580);
nand I_19888 (I340319,I340622,I340441);
nand I_19889 (I340653,I739382,I739397);
and I_19890 (I340670,I340653,I739382);
DFFARX1 I_19891 (I340670,I2507,I340342,I340696,);
nor I_19892 (I340704,I340696,I340368);
DFFARX1 I_19893 (I340704,I2507,I340342,I340307,);
DFFARX1 I_19894 (I340696,I2507,I340342,I340325,);
nor I_19895 (I340749,I739403,I739397);
not I_19896 (I340766,I340749);
nor I_19897 (I340328,I340605,I340766);
nand I_19898 (I340313,I340622,I340766);
nor I_19899 (I340322,I340368,I340749);
DFFARX1 I_19900 (I340749,I2507,I340342,I340331,);
not I_19901 (I340869,I2514);
DFFARX1 I_19902 (I1296370,I2507,I340869,I340895,);
nand I_19903 (I340903,I1296397,I1296373);
and I_19904 (I340920,I340903,I1296382);
DFFARX1 I_19905 (I340920,I2507,I340869,I340946,);
nor I_19906 (I340837,I340946,I340895);
not I_19907 (I340968,I340946);
DFFARX1 I_19908 (I1296370,I2507,I340869,I340994,);
nand I_19909 (I341002,I340994,I1296394);
not I_19910 (I341019,I341002);
DFFARX1 I_19911 (I341019,I2507,I340869,I341045,);
not I_19912 (I340861,I341045);
nor I_19913 (I341067,I340895,I341002);
nor I_19914 (I340843,I340946,I341067);
DFFARX1 I_19915 (I1296376,I2507,I340869,I341107,);
DFFARX1 I_19916 (I341107,I2507,I340869,I341124,);
not I_19917 (I341132,I341124);
not I_19918 (I341149,I341107);
nand I_19919 (I340846,I341149,I340968);
nand I_19920 (I341180,I1296391,I1296379);
and I_19921 (I341197,I341180,I1296385);
DFFARX1 I_19922 (I341197,I2507,I340869,I341223,);
nor I_19923 (I341231,I341223,I340895);
DFFARX1 I_19924 (I341231,I2507,I340869,I340834,);
DFFARX1 I_19925 (I341223,I2507,I340869,I340852,);
nor I_19926 (I341276,I1296388,I1296379);
not I_19927 (I341293,I341276);
nor I_19928 (I340855,I341132,I341293);
nand I_19929 (I340840,I341149,I341293);
nor I_19930 (I340849,I340895,I341276);
DFFARX1 I_19931 (I341276,I2507,I340869,I340858,);
not I_19932 (I341396,I2514);
DFFARX1 I_19933 (I1322588,I2507,I341396,I341422,);
nand I_19934 (I341430,I1322567,I1322567);
and I_19935 (I341447,I341430,I1322594);
DFFARX1 I_19936 (I341447,I2507,I341396,I341473,);
nor I_19937 (I341364,I341473,I341422);
not I_19938 (I341495,I341473);
DFFARX1 I_19939 (I1322582,I2507,I341396,I341521,);
nand I_19940 (I341529,I341521,I1322585);
not I_19941 (I341546,I341529);
DFFARX1 I_19942 (I341546,I2507,I341396,I341572,);
not I_19943 (I341388,I341572);
nor I_19944 (I341594,I341422,I341529);
nor I_19945 (I341370,I341473,I341594);
DFFARX1 I_19946 (I1322576,I2507,I341396,I341634,);
DFFARX1 I_19947 (I341634,I2507,I341396,I341651,);
not I_19948 (I341659,I341651);
not I_19949 (I341676,I341634);
nand I_19950 (I341373,I341676,I341495);
nand I_19951 (I341707,I1322573,I1322570);
and I_19952 (I341724,I341707,I1322591);
DFFARX1 I_19953 (I341724,I2507,I341396,I341750,);
nor I_19954 (I341758,I341750,I341422);
DFFARX1 I_19955 (I341758,I2507,I341396,I341361,);
DFFARX1 I_19956 (I341750,I2507,I341396,I341379,);
nor I_19957 (I341803,I1322579,I1322570);
not I_19958 (I341820,I341803);
nor I_19959 (I341382,I341659,I341820);
nand I_19960 (I341367,I341676,I341820);
nor I_19961 (I341376,I341422,I341803);
DFFARX1 I_19962 (I341803,I2507,I341396,I341385,);
not I_19963 (I341923,I2514);
DFFARX1 I_19964 (I93861,I2507,I341923,I341949,);
nand I_19965 (I341957,I93873,I93882);
and I_19966 (I341974,I341957,I93861);
DFFARX1 I_19967 (I341974,I2507,I341923,I342000,);
nor I_19968 (I341891,I342000,I341949);
not I_19969 (I342022,I342000);
DFFARX1 I_19970 (I93876,I2507,I341923,I342048,);
nand I_19971 (I342056,I342048,I93864);
not I_19972 (I342073,I342056);
DFFARX1 I_19973 (I342073,I2507,I341923,I342099,);
not I_19974 (I341915,I342099);
nor I_19975 (I342121,I341949,I342056);
nor I_19976 (I341897,I342000,I342121);
DFFARX1 I_19977 (I93867,I2507,I341923,I342161,);
DFFARX1 I_19978 (I342161,I2507,I341923,I342178,);
not I_19979 (I342186,I342178);
not I_19980 (I342203,I342161);
nand I_19981 (I341900,I342203,I342022);
nand I_19982 (I342234,I93858,I93858);
and I_19983 (I342251,I342234,I93870);
DFFARX1 I_19984 (I342251,I2507,I341923,I342277,);
nor I_19985 (I342285,I342277,I341949);
DFFARX1 I_19986 (I342285,I2507,I341923,I341888,);
DFFARX1 I_19987 (I342277,I2507,I341923,I341906,);
nor I_19988 (I342330,I93879,I93858);
not I_19989 (I342347,I342330);
nor I_19990 (I341909,I342186,I342347);
nand I_19991 (I341894,I342203,I342347);
nor I_19992 (I341903,I341949,I342330);
DFFARX1 I_19993 (I342330,I2507,I341923,I341912,);
not I_19994 (I342450,I2514);
DFFARX1 I_19995 (I920520,I2507,I342450,I342476,);
nand I_19996 (I342484,I920517,I920535);
and I_19997 (I342501,I342484,I920526);
DFFARX1 I_19998 (I342501,I2507,I342450,I342527,);
nor I_19999 (I342418,I342527,I342476);
not I_20000 (I342549,I342527);
DFFARX1 I_20001 (I920541,I2507,I342450,I342575,);
nand I_20002 (I342583,I342575,I920523);
not I_20003 (I342600,I342583);
DFFARX1 I_20004 (I342600,I2507,I342450,I342626,);
not I_20005 (I342442,I342626);
nor I_20006 (I342648,I342476,I342583);
nor I_20007 (I342424,I342527,I342648);
DFFARX1 I_20008 (I920529,I2507,I342450,I342688,);
DFFARX1 I_20009 (I342688,I2507,I342450,I342705,);
not I_20010 (I342713,I342705);
not I_20011 (I342730,I342688);
nand I_20012 (I342427,I342730,I342549);
nand I_20013 (I342761,I920517,I920544);
and I_20014 (I342778,I342761,I920532);
DFFARX1 I_20015 (I342778,I2507,I342450,I342804,);
nor I_20016 (I342812,I342804,I342476);
DFFARX1 I_20017 (I342812,I2507,I342450,I342415,);
DFFARX1 I_20018 (I342804,I2507,I342450,I342433,);
nor I_20019 (I342857,I920538,I920544);
not I_20020 (I342874,I342857);
nor I_20021 (I342436,I342713,I342874);
nand I_20022 (I342421,I342730,I342874);
nor I_20023 (I342430,I342476,I342857);
DFFARX1 I_20024 (I342857,I2507,I342450,I342439,);
not I_20025 (I342977,I2514);
DFFARX1 I_20026 (I397915,I2507,I342977,I343003,);
nand I_20027 (I343011,I397927,I397906);
and I_20028 (I343028,I343011,I397930);
DFFARX1 I_20029 (I343028,I2507,I342977,I343054,);
nor I_20030 (I342945,I343054,I343003);
not I_20031 (I343076,I343054);
DFFARX1 I_20032 (I397921,I2507,I342977,I343102,);
nand I_20033 (I343110,I343102,I397903);
not I_20034 (I343127,I343110);
DFFARX1 I_20035 (I343127,I2507,I342977,I343153,);
not I_20036 (I342969,I343153);
nor I_20037 (I343175,I343003,I343110);
nor I_20038 (I342951,I343054,I343175);
DFFARX1 I_20039 (I397918,I2507,I342977,I343215,);
DFFARX1 I_20040 (I343215,I2507,I342977,I343232,);
not I_20041 (I343240,I343232);
not I_20042 (I343257,I343215);
nand I_20043 (I342954,I343257,I343076);
nand I_20044 (I343288,I397903,I397909);
and I_20045 (I343305,I343288,I397912);
DFFARX1 I_20046 (I343305,I2507,I342977,I343331,);
nor I_20047 (I343339,I343331,I343003);
DFFARX1 I_20048 (I343339,I2507,I342977,I342942,);
DFFARX1 I_20049 (I343331,I2507,I342977,I342960,);
nor I_20050 (I343384,I397924,I397909);
not I_20051 (I343401,I343384);
nor I_20052 (I342963,I343240,I343401);
nand I_20053 (I342948,I343257,I343401);
nor I_20054 (I342957,I343003,I343384);
DFFARX1 I_20055 (I343384,I2507,I342977,I342966,);
not I_20056 (I343504,I2514);
DFFARX1 I_20057 (I413691,I2507,I343504,I343530,);
nand I_20058 (I343538,I413703,I413682);
and I_20059 (I343555,I343538,I413706);
DFFARX1 I_20060 (I343555,I2507,I343504,I343581,);
nor I_20061 (I343472,I343581,I343530);
not I_20062 (I343603,I343581);
DFFARX1 I_20063 (I413697,I2507,I343504,I343629,);
nand I_20064 (I343637,I343629,I413679);
not I_20065 (I343654,I343637);
DFFARX1 I_20066 (I343654,I2507,I343504,I343680,);
not I_20067 (I343496,I343680);
nor I_20068 (I343702,I343530,I343637);
nor I_20069 (I343478,I343581,I343702);
DFFARX1 I_20070 (I413694,I2507,I343504,I343742,);
DFFARX1 I_20071 (I343742,I2507,I343504,I343759,);
not I_20072 (I343767,I343759);
not I_20073 (I343784,I343742);
nand I_20074 (I343481,I343784,I343603);
nand I_20075 (I343815,I413679,I413685);
and I_20076 (I343832,I343815,I413688);
DFFARX1 I_20077 (I343832,I2507,I343504,I343858,);
nor I_20078 (I343866,I343858,I343530);
DFFARX1 I_20079 (I343866,I2507,I343504,I343469,);
DFFARX1 I_20080 (I343858,I2507,I343504,I343487,);
nor I_20081 (I343911,I413700,I413685);
not I_20082 (I343928,I343911);
nor I_20083 (I343490,I343767,I343928);
nand I_20084 (I343475,I343784,I343928);
nor I_20085 (I343484,I343530,I343911);
DFFARX1 I_20086 (I343911,I2507,I343504,I343493,);
not I_20087 (I344031,I2514);
DFFARX1 I_20088 (I384315,I2507,I344031,I344057,);
nand I_20089 (I344065,I384327,I384306);
and I_20090 (I344082,I344065,I384330);
DFFARX1 I_20091 (I344082,I2507,I344031,I344108,);
nor I_20092 (I343999,I344108,I344057);
not I_20093 (I344130,I344108);
DFFARX1 I_20094 (I384321,I2507,I344031,I344156,);
nand I_20095 (I344164,I344156,I384303);
not I_20096 (I344181,I344164);
DFFARX1 I_20097 (I344181,I2507,I344031,I344207,);
not I_20098 (I344023,I344207);
nor I_20099 (I344229,I344057,I344164);
nor I_20100 (I344005,I344108,I344229);
DFFARX1 I_20101 (I384318,I2507,I344031,I344269,);
DFFARX1 I_20102 (I344269,I2507,I344031,I344286,);
not I_20103 (I344294,I344286);
not I_20104 (I344311,I344269);
nand I_20105 (I344008,I344311,I344130);
nand I_20106 (I344342,I384303,I384309);
and I_20107 (I344359,I344342,I384312);
DFFARX1 I_20108 (I344359,I2507,I344031,I344385,);
nor I_20109 (I344393,I344385,I344057);
DFFARX1 I_20110 (I344393,I2507,I344031,I343996,);
DFFARX1 I_20111 (I344385,I2507,I344031,I344014,);
nor I_20112 (I344438,I384324,I384309);
not I_20113 (I344455,I344438);
nor I_20114 (I344017,I344294,I344455);
nand I_20115 (I344002,I344311,I344455);
nor I_20116 (I344011,I344057,I344438);
DFFARX1 I_20117 (I344438,I2507,I344031,I344020,);
not I_20118 (I344558,I2514);
DFFARX1 I_20119 (I1101720,I2507,I344558,I344584,);
nand I_20120 (I344592,I1101735,I1101720);
and I_20121 (I344609,I344592,I1101738);
DFFARX1 I_20122 (I344609,I2507,I344558,I344635,);
nor I_20123 (I344526,I344635,I344584);
not I_20124 (I344657,I344635);
DFFARX1 I_20125 (I1101744,I2507,I344558,I344683,);
nand I_20126 (I344691,I344683,I1101726);
not I_20127 (I344708,I344691);
DFFARX1 I_20128 (I344708,I2507,I344558,I344734,);
not I_20129 (I344550,I344734);
nor I_20130 (I344756,I344584,I344691);
nor I_20131 (I344532,I344635,I344756);
DFFARX1 I_20132 (I1101723,I2507,I344558,I344796,);
DFFARX1 I_20133 (I344796,I2507,I344558,I344813,);
not I_20134 (I344821,I344813);
not I_20135 (I344838,I344796);
nand I_20136 (I344535,I344838,I344657);
nand I_20137 (I344869,I1101723,I1101729);
and I_20138 (I344886,I344869,I1101741);
DFFARX1 I_20139 (I344886,I2507,I344558,I344912,);
nor I_20140 (I344920,I344912,I344584);
DFFARX1 I_20141 (I344920,I2507,I344558,I344523,);
DFFARX1 I_20142 (I344912,I2507,I344558,I344541,);
nor I_20143 (I344965,I1101732,I1101729);
not I_20144 (I344982,I344965);
nor I_20145 (I344544,I344821,I344982);
nand I_20146 (I344529,I344838,I344982);
nor I_20147 (I344538,I344584,I344965);
DFFARX1 I_20148 (I344965,I2507,I344558,I344547,);
not I_20149 (I345085,I2514);
DFFARX1 I_20150 (I914706,I2507,I345085,I345111,);
nand I_20151 (I345119,I914703,I914721);
and I_20152 (I345136,I345119,I914712);
DFFARX1 I_20153 (I345136,I2507,I345085,I345162,);
nor I_20154 (I345053,I345162,I345111);
not I_20155 (I345184,I345162);
DFFARX1 I_20156 (I914727,I2507,I345085,I345210,);
nand I_20157 (I345218,I345210,I914709);
not I_20158 (I345235,I345218);
DFFARX1 I_20159 (I345235,I2507,I345085,I345261,);
not I_20160 (I345077,I345261);
nor I_20161 (I345283,I345111,I345218);
nor I_20162 (I345059,I345162,I345283);
DFFARX1 I_20163 (I914715,I2507,I345085,I345323,);
DFFARX1 I_20164 (I345323,I2507,I345085,I345340,);
not I_20165 (I345348,I345340);
not I_20166 (I345365,I345323);
nand I_20167 (I345062,I345365,I345184);
nand I_20168 (I345396,I914703,I914730);
and I_20169 (I345413,I345396,I914718);
DFFARX1 I_20170 (I345413,I2507,I345085,I345439,);
nor I_20171 (I345447,I345439,I345111);
DFFARX1 I_20172 (I345447,I2507,I345085,I345050,);
DFFARX1 I_20173 (I345439,I2507,I345085,I345068,);
nor I_20174 (I345492,I914724,I914730);
not I_20175 (I345509,I345492);
nor I_20176 (I345071,I345348,I345509);
nand I_20177 (I345056,I345365,I345509);
nor I_20178 (I345065,I345111,I345492);
DFFARX1 I_20179 (I345492,I2507,I345085,I345074,);
not I_20180 (I345612,I2514);
DFFARX1 I_20181 (I1303102,I2507,I345612,I345638,);
nand I_20182 (I345646,I1303129,I1303105);
and I_20183 (I345663,I345646,I1303114);
DFFARX1 I_20184 (I345663,I2507,I345612,I345689,);
nor I_20185 (I345580,I345689,I345638);
not I_20186 (I345711,I345689);
DFFARX1 I_20187 (I1303102,I2507,I345612,I345737,);
nand I_20188 (I345745,I345737,I1303126);
not I_20189 (I345762,I345745);
DFFARX1 I_20190 (I345762,I2507,I345612,I345788,);
not I_20191 (I345604,I345788);
nor I_20192 (I345810,I345638,I345745);
nor I_20193 (I345586,I345689,I345810);
DFFARX1 I_20194 (I1303108,I2507,I345612,I345850,);
DFFARX1 I_20195 (I345850,I2507,I345612,I345867,);
not I_20196 (I345875,I345867);
not I_20197 (I345892,I345850);
nand I_20198 (I345589,I345892,I345711);
nand I_20199 (I345923,I1303123,I1303111);
and I_20200 (I345940,I345923,I1303117);
DFFARX1 I_20201 (I345940,I2507,I345612,I345966,);
nor I_20202 (I345974,I345966,I345638);
DFFARX1 I_20203 (I345974,I2507,I345612,I345577,);
DFFARX1 I_20204 (I345966,I2507,I345612,I345595,);
nor I_20205 (I346019,I1303120,I1303111);
not I_20206 (I346036,I346019);
nor I_20207 (I345598,I345875,I346036);
nand I_20208 (I345583,I345892,I346036);
nor I_20209 (I345592,I345638,I346019);
DFFARX1 I_20210 (I346019,I2507,I345612,I345601,);
not I_20211 (I346139,I2514);
DFFARX1 I_20212 (I229365,I2507,I346139,I346165,);
nand I_20213 (I346173,I229365,I229371);
and I_20214 (I346190,I346173,I229389);
DFFARX1 I_20215 (I346190,I2507,I346139,I346216,);
nor I_20216 (I346107,I346216,I346165);
not I_20217 (I346238,I346216);
DFFARX1 I_20218 (I229377,I2507,I346139,I346264,);
nand I_20219 (I346272,I346264,I229374);
not I_20220 (I346289,I346272);
DFFARX1 I_20221 (I346289,I2507,I346139,I346315,);
not I_20222 (I346131,I346315);
nor I_20223 (I346337,I346165,I346272);
nor I_20224 (I346113,I346216,I346337);
DFFARX1 I_20225 (I229383,I2507,I346139,I346377,);
DFFARX1 I_20226 (I346377,I2507,I346139,I346394,);
not I_20227 (I346402,I346394);
not I_20228 (I346419,I346377);
nand I_20229 (I346116,I346419,I346238);
nand I_20230 (I346450,I229368,I229368);
and I_20231 (I346467,I346450,I229380);
DFFARX1 I_20232 (I346467,I2507,I346139,I346493,);
nor I_20233 (I346501,I346493,I346165);
DFFARX1 I_20234 (I346501,I2507,I346139,I346104,);
DFFARX1 I_20235 (I346493,I2507,I346139,I346122,);
nor I_20236 (I346546,I229386,I229368);
not I_20237 (I346563,I346546);
nor I_20238 (I346125,I346402,I346563);
nand I_20239 (I346110,I346419,I346563);
nor I_20240 (I346119,I346165,I346546);
DFFARX1 I_20241 (I346546,I2507,I346139,I346128,);
not I_20242 (I346666,I2514);
DFFARX1 I_20243 (I163320,I2507,I346666,I346692,);
nand I_20244 (I346700,I163320,I163326);
and I_20245 (I346717,I346700,I163344);
DFFARX1 I_20246 (I346717,I2507,I346666,I346743,);
nor I_20247 (I346634,I346743,I346692);
not I_20248 (I346765,I346743);
DFFARX1 I_20249 (I163332,I2507,I346666,I346791,);
nand I_20250 (I346799,I346791,I163329);
not I_20251 (I346816,I346799);
DFFARX1 I_20252 (I346816,I2507,I346666,I346842,);
not I_20253 (I346658,I346842);
nor I_20254 (I346864,I346692,I346799);
nor I_20255 (I346640,I346743,I346864);
DFFARX1 I_20256 (I163338,I2507,I346666,I346904,);
DFFARX1 I_20257 (I346904,I2507,I346666,I346921,);
not I_20258 (I346929,I346921);
not I_20259 (I346946,I346904);
nand I_20260 (I346643,I346946,I346765);
nand I_20261 (I346977,I163323,I163323);
and I_20262 (I346994,I346977,I163335);
DFFARX1 I_20263 (I346994,I2507,I346666,I347020,);
nor I_20264 (I347028,I347020,I346692);
DFFARX1 I_20265 (I347028,I2507,I346666,I346631,);
DFFARX1 I_20266 (I347020,I2507,I346666,I346649,);
nor I_20267 (I347073,I163341,I163323);
not I_20268 (I347090,I347073);
nor I_20269 (I346652,I346929,I347090);
nand I_20270 (I346637,I346946,I347090);
nor I_20271 (I346646,I346692,I347073);
DFFARX1 I_20272 (I347073,I2507,I346666,I346655,);
not I_20273 (I347193,I2514);
DFFARX1 I_20274 (I131805,I2507,I347193,I347219,);
nand I_20275 (I347227,I131817,I131826);
and I_20276 (I347244,I347227,I131805);
DFFARX1 I_20277 (I347244,I2507,I347193,I347270,);
nor I_20278 (I347161,I347270,I347219);
not I_20279 (I347292,I347270);
DFFARX1 I_20280 (I131820,I2507,I347193,I347318,);
nand I_20281 (I347326,I347318,I131808);
not I_20282 (I347343,I347326);
DFFARX1 I_20283 (I347343,I2507,I347193,I347369,);
not I_20284 (I347185,I347369);
nor I_20285 (I347391,I347219,I347326);
nor I_20286 (I347167,I347270,I347391);
DFFARX1 I_20287 (I131811,I2507,I347193,I347431,);
DFFARX1 I_20288 (I347431,I2507,I347193,I347448,);
not I_20289 (I347456,I347448);
not I_20290 (I347473,I347431);
nand I_20291 (I347170,I347473,I347292);
nand I_20292 (I347504,I131802,I131802);
and I_20293 (I347521,I347504,I131814);
DFFARX1 I_20294 (I347521,I2507,I347193,I347547,);
nor I_20295 (I347555,I347547,I347219);
DFFARX1 I_20296 (I347555,I2507,I347193,I347158,);
DFFARX1 I_20297 (I347547,I2507,I347193,I347176,);
nor I_20298 (I347600,I131823,I131802);
not I_20299 (I347617,I347600);
nor I_20300 (I347179,I347456,I347617);
nand I_20301 (I347164,I347473,I347617);
nor I_20302 (I347173,I347219,I347600);
DFFARX1 I_20303 (I347600,I2507,I347193,I347182,);
not I_20304 (I347720,I2514);
DFFARX1 I_20305 (I134440,I2507,I347720,I347746,);
nand I_20306 (I347754,I134452,I134461);
and I_20307 (I347771,I347754,I134440);
DFFARX1 I_20308 (I347771,I2507,I347720,I347797,);
nor I_20309 (I347688,I347797,I347746);
not I_20310 (I347819,I347797);
DFFARX1 I_20311 (I134455,I2507,I347720,I347845,);
nand I_20312 (I347853,I347845,I134443);
not I_20313 (I347870,I347853);
DFFARX1 I_20314 (I347870,I2507,I347720,I347896,);
not I_20315 (I347712,I347896);
nor I_20316 (I347918,I347746,I347853);
nor I_20317 (I347694,I347797,I347918);
DFFARX1 I_20318 (I134446,I2507,I347720,I347958,);
DFFARX1 I_20319 (I347958,I2507,I347720,I347975,);
not I_20320 (I347983,I347975);
not I_20321 (I348000,I347958);
nand I_20322 (I347697,I348000,I347819);
nand I_20323 (I348031,I134437,I134437);
and I_20324 (I348048,I348031,I134449);
DFFARX1 I_20325 (I348048,I2507,I347720,I348074,);
nor I_20326 (I348082,I348074,I347746);
DFFARX1 I_20327 (I348082,I2507,I347720,I347685,);
DFFARX1 I_20328 (I348074,I2507,I347720,I347703,);
nor I_20329 (I348127,I134458,I134437);
not I_20330 (I348144,I348127);
nor I_20331 (I347706,I347983,I348144);
nand I_20332 (I347691,I348000,I348144);
nor I_20333 (I347700,I347746,I348127);
DFFARX1 I_20334 (I348127,I2507,I347720,I347709,);
not I_20335 (I348247,I2514);
DFFARX1 I_20336 (I635354,I2507,I348247,I348273,);
nand I_20337 (I348281,I635345,I635360);
and I_20338 (I348298,I348281,I635366);
DFFARX1 I_20339 (I348298,I2507,I348247,I348324,);
nor I_20340 (I348215,I348324,I348273);
not I_20341 (I348346,I348324);
DFFARX1 I_20342 (I635351,I2507,I348247,I348372,);
nand I_20343 (I348380,I348372,I635345);
not I_20344 (I348397,I348380);
DFFARX1 I_20345 (I348397,I2507,I348247,I348423,);
not I_20346 (I348239,I348423);
nor I_20347 (I348445,I348273,I348380);
nor I_20348 (I348221,I348324,I348445);
DFFARX1 I_20349 (I635348,I2507,I348247,I348485,);
DFFARX1 I_20350 (I348485,I2507,I348247,I348502,);
not I_20351 (I348510,I348502);
not I_20352 (I348527,I348485);
nand I_20353 (I348224,I348527,I348346);
nand I_20354 (I348558,I635342,I635357);
and I_20355 (I348575,I348558,I635342);
DFFARX1 I_20356 (I348575,I2507,I348247,I348601,);
nor I_20357 (I348609,I348601,I348273);
DFFARX1 I_20358 (I348609,I2507,I348247,I348212,);
DFFARX1 I_20359 (I348601,I2507,I348247,I348230,);
nor I_20360 (I348654,I635363,I635357);
not I_20361 (I348671,I348654);
nor I_20362 (I348233,I348510,I348671);
nand I_20363 (I348218,I348527,I348671);
nor I_20364 (I348227,I348273,I348654);
DFFARX1 I_20365 (I348654,I2507,I348247,I348236,);
not I_20366 (I348774,I2514);
DFFARX1 I_20367 (I1002562,I2507,I348774,I348800,);
nand I_20368 (I348808,I1002559,I1002577);
and I_20369 (I348825,I348808,I1002568);
DFFARX1 I_20370 (I348825,I2507,I348774,I348851,);
nor I_20371 (I348742,I348851,I348800);
not I_20372 (I348873,I348851);
DFFARX1 I_20373 (I1002583,I2507,I348774,I348899,);
nand I_20374 (I348907,I348899,I1002565);
not I_20375 (I348924,I348907);
DFFARX1 I_20376 (I348924,I2507,I348774,I348950,);
not I_20377 (I348766,I348950);
nor I_20378 (I348972,I348800,I348907);
nor I_20379 (I348748,I348851,I348972);
DFFARX1 I_20380 (I1002571,I2507,I348774,I349012,);
DFFARX1 I_20381 (I349012,I2507,I348774,I349029,);
not I_20382 (I349037,I349029);
not I_20383 (I349054,I349012);
nand I_20384 (I348751,I349054,I348873);
nand I_20385 (I349085,I1002559,I1002586);
and I_20386 (I349102,I349085,I1002574);
DFFARX1 I_20387 (I349102,I2507,I348774,I349128,);
nor I_20388 (I349136,I349128,I348800);
DFFARX1 I_20389 (I349136,I2507,I348774,I348739,);
DFFARX1 I_20390 (I349128,I2507,I348774,I348757,);
nor I_20391 (I349181,I1002580,I1002586);
not I_20392 (I349198,I349181);
nor I_20393 (I348760,I349037,I349198);
nand I_20394 (I348745,I349054,I349198);
nor I_20395 (I348754,I348800,I349181);
DFFARX1 I_20396 (I349181,I2507,I348774,I348763,);
not I_20397 (I349301,I2514);
DFFARX1 I_20398 (I828074,I2507,I349301,I349327,);
nand I_20399 (I349335,I828077,I828071);
and I_20400 (I349352,I349335,I828083);
DFFARX1 I_20401 (I349352,I2507,I349301,I349378,);
nor I_20402 (I349269,I349378,I349327);
not I_20403 (I349400,I349378);
DFFARX1 I_20404 (I828086,I2507,I349301,I349426,);
nand I_20405 (I349434,I349426,I828077);
not I_20406 (I349451,I349434);
DFFARX1 I_20407 (I349451,I2507,I349301,I349477,);
not I_20408 (I349293,I349477);
nor I_20409 (I349499,I349327,I349434);
nor I_20410 (I349275,I349378,I349499);
DFFARX1 I_20411 (I828089,I2507,I349301,I349539,);
DFFARX1 I_20412 (I349539,I2507,I349301,I349556,);
not I_20413 (I349564,I349556);
not I_20414 (I349581,I349539);
nand I_20415 (I349278,I349581,I349400);
nand I_20416 (I349612,I828071,I828080);
and I_20417 (I349629,I349612,I828074);
DFFARX1 I_20418 (I349629,I2507,I349301,I349655,);
nor I_20419 (I349663,I349655,I349327);
DFFARX1 I_20420 (I349663,I2507,I349301,I349266,);
DFFARX1 I_20421 (I349655,I2507,I349301,I349284,);
nor I_20422 (I349708,I828092,I828080);
not I_20423 (I349725,I349708);
nor I_20424 (I349287,I349564,I349725);
nand I_20425 (I349272,I349581,I349725);
nor I_20426 (I349281,I349327,I349708);
DFFARX1 I_20427 (I349708,I2507,I349301,I349290,);
not I_20428 (I349828,I2514);
DFFARX1 I_20429 (I1078600,I2507,I349828,I349854,);
nand I_20430 (I349862,I1078615,I1078600);
and I_20431 (I349879,I349862,I1078618);
DFFARX1 I_20432 (I349879,I2507,I349828,I349905,);
nor I_20433 (I349796,I349905,I349854);
not I_20434 (I349927,I349905);
DFFARX1 I_20435 (I1078624,I2507,I349828,I349953,);
nand I_20436 (I349961,I349953,I1078606);
not I_20437 (I349978,I349961);
DFFARX1 I_20438 (I349978,I2507,I349828,I350004,);
not I_20439 (I349820,I350004);
nor I_20440 (I350026,I349854,I349961);
nor I_20441 (I349802,I349905,I350026);
DFFARX1 I_20442 (I1078603,I2507,I349828,I350066,);
DFFARX1 I_20443 (I350066,I2507,I349828,I350083,);
not I_20444 (I350091,I350083);
not I_20445 (I350108,I350066);
nand I_20446 (I349805,I350108,I349927);
nand I_20447 (I350139,I1078603,I1078609);
and I_20448 (I350156,I350139,I1078621);
DFFARX1 I_20449 (I350156,I2507,I349828,I350182,);
nor I_20450 (I350190,I350182,I349854);
DFFARX1 I_20451 (I350190,I2507,I349828,I349793,);
DFFARX1 I_20452 (I350182,I2507,I349828,I349811,);
nor I_20453 (I350235,I1078612,I1078609);
not I_20454 (I350252,I350235);
nor I_20455 (I349814,I350091,I350252);
nand I_20456 (I349799,I350108,I350252);
nor I_20457 (I349808,I349854,I350235);
DFFARX1 I_20458 (I350235,I2507,I349828,I349817,);
not I_20459 (I350355,I2514);
DFFARX1 I_20460 (I983182,I2507,I350355,I350381,);
nand I_20461 (I350389,I983179,I983197);
and I_20462 (I350406,I350389,I983188);
DFFARX1 I_20463 (I350406,I2507,I350355,I350432,);
nor I_20464 (I350323,I350432,I350381);
not I_20465 (I350454,I350432);
DFFARX1 I_20466 (I983203,I2507,I350355,I350480,);
nand I_20467 (I350488,I350480,I983185);
not I_20468 (I350505,I350488);
DFFARX1 I_20469 (I350505,I2507,I350355,I350531,);
not I_20470 (I350347,I350531);
nor I_20471 (I350553,I350381,I350488);
nor I_20472 (I350329,I350432,I350553);
DFFARX1 I_20473 (I983191,I2507,I350355,I350593,);
DFFARX1 I_20474 (I350593,I2507,I350355,I350610,);
not I_20475 (I350618,I350610);
not I_20476 (I350635,I350593);
nand I_20477 (I350332,I350635,I350454);
nand I_20478 (I350666,I983179,I983206);
and I_20479 (I350683,I350666,I983194);
DFFARX1 I_20480 (I350683,I2507,I350355,I350709,);
nor I_20481 (I350717,I350709,I350381);
DFFARX1 I_20482 (I350717,I2507,I350355,I350320,);
DFFARX1 I_20483 (I350709,I2507,I350355,I350338,);
nor I_20484 (I350762,I983200,I983206);
not I_20485 (I350779,I350762);
nor I_20486 (I350341,I350618,I350779);
nand I_20487 (I350326,I350635,I350779);
nor I_20488 (I350335,I350381,I350762);
DFFARX1 I_20489 (I350762,I2507,I350355,I350344,);
not I_20490 (I350882,I2514);
DFFARX1 I_20491 (I833344,I2507,I350882,I350908,);
nand I_20492 (I350916,I833347,I833341);
and I_20493 (I350933,I350916,I833353);
DFFARX1 I_20494 (I350933,I2507,I350882,I350959,);
nor I_20495 (I350850,I350959,I350908);
not I_20496 (I350981,I350959);
DFFARX1 I_20497 (I833356,I2507,I350882,I351007,);
nand I_20498 (I351015,I351007,I833347);
not I_20499 (I351032,I351015);
DFFARX1 I_20500 (I351032,I2507,I350882,I351058,);
not I_20501 (I350874,I351058);
nor I_20502 (I351080,I350908,I351015);
nor I_20503 (I350856,I350959,I351080);
DFFARX1 I_20504 (I833359,I2507,I350882,I351120,);
DFFARX1 I_20505 (I351120,I2507,I350882,I351137,);
not I_20506 (I351145,I351137);
not I_20507 (I351162,I351120);
nand I_20508 (I350859,I351162,I350981);
nand I_20509 (I351193,I833341,I833350);
and I_20510 (I351210,I351193,I833344);
DFFARX1 I_20511 (I351210,I2507,I350882,I351236,);
nor I_20512 (I351244,I351236,I350908);
DFFARX1 I_20513 (I351244,I2507,I350882,I350847,);
DFFARX1 I_20514 (I351236,I2507,I350882,I350865,);
nor I_20515 (I351289,I833362,I833350);
not I_20516 (I351306,I351289);
nor I_20517 (I350868,I351145,I351306);
nand I_20518 (I350853,I351162,I351306);
nor I_20519 (I350862,I350908,I351289);
DFFARX1 I_20520 (I351289,I2507,I350882,I350871,);
not I_20521 (I351409,I2514);
DFFARX1 I_20522 (I385947,I2507,I351409,I351435,);
nand I_20523 (I351443,I385959,I385938);
and I_20524 (I351460,I351443,I385962);
DFFARX1 I_20525 (I351460,I2507,I351409,I351486,);
nor I_20526 (I351377,I351486,I351435);
not I_20527 (I351508,I351486);
DFFARX1 I_20528 (I385953,I2507,I351409,I351534,);
nand I_20529 (I351542,I351534,I385935);
not I_20530 (I351559,I351542);
DFFARX1 I_20531 (I351559,I2507,I351409,I351585,);
not I_20532 (I351401,I351585);
nor I_20533 (I351607,I351435,I351542);
nor I_20534 (I351383,I351486,I351607);
DFFARX1 I_20535 (I385950,I2507,I351409,I351647,);
DFFARX1 I_20536 (I351647,I2507,I351409,I351664,);
not I_20537 (I351672,I351664);
not I_20538 (I351689,I351647);
nand I_20539 (I351386,I351689,I351508);
nand I_20540 (I351720,I385935,I385941);
and I_20541 (I351737,I351720,I385944);
DFFARX1 I_20542 (I351737,I2507,I351409,I351763,);
nor I_20543 (I351771,I351763,I351435);
DFFARX1 I_20544 (I351771,I2507,I351409,I351374,);
DFFARX1 I_20545 (I351763,I2507,I351409,I351392,);
nor I_20546 (I351816,I385956,I385941);
not I_20547 (I351833,I351816);
nor I_20548 (I351395,I351672,I351833);
nand I_20549 (I351380,I351689,I351833);
nor I_20550 (I351389,I351435,I351816);
DFFARX1 I_20551 (I351816,I2507,I351409,I351398,);
not I_20552 (I351936,I2514);
DFFARX1 I_20553 (I9077,I2507,I351936,I351962,);
nand I_20554 (I351970,I9068,I9071);
and I_20555 (I351987,I351970,I9062);
DFFARX1 I_20556 (I351987,I2507,I351936,I352013,);
nor I_20557 (I351904,I352013,I351962);
not I_20558 (I352035,I352013);
DFFARX1 I_20559 (I9068,I2507,I351936,I352061,);
nand I_20560 (I352069,I352061,I9074);
not I_20561 (I352086,I352069);
DFFARX1 I_20562 (I352086,I2507,I351936,I352112,);
not I_20563 (I351928,I352112);
nor I_20564 (I352134,I351962,I352069);
nor I_20565 (I351910,I352013,I352134);
DFFARX1 I_20566 (I9065,I2507,I351936,I352174,);
DFFARX1 I_20567 (I352174,I2507,I351936,I352191,);
not I_20568 (I352199,I352191);
not I_20569 (I352216,I352174);
nand I_20570 (I351913,I352216,I352035);
nand I_20571 (I352247,I9065,I9080);
and I_20572 (I352264,I352247,I9062);
DFFARX1 I_20573 (I352264,I2507,I351936,I352290,);
nor I_20574 (I352298,I352290,I351962);
DFFARX1 I_20575 (I352298,I2507,I351936,I351901,);
DFFARX1 I_20576 (I352290,I2507,I351936,I351919,);
nor I_20577 (I352343,I9083,I9080);
not I_20578 (I352360,I352343);
nor I_20579 (I351922,I352199,I352360);
nand I_20580 (I351907,I352216,I352360);
nor I_20581 (I351916,I351962,I352343);
DFFARX1 I_20582 (I352343,I2507,I351936,I351925,);
not I_20583 (I352463,I2514);
DFFARX1 I_20584 (I9672,I2507,I352463,I352489,);
nand I_20585 (I352497,I9663,I9666);
and I_20586 (I352514,I352497,I9657);
DFFARX1 I_20587 (I352514,I2507,I352463,I352540,);
nor I_20588 (I352431,I352540,I352489);
not I_20589 (I352562,I352540);
DFFARX1 I_20590 (I9663,I2507,I352463,I352588,);
nand I_20591 (I352596,I352588,I9669);
not I_20592 (I352613,I352596);
DFFARX1 I_20593 (I352613,I2507,I352463,I352639,);
not I_20594 (I352455,I352639);
nor I_20595 (I352661,I352489,I352596);
nor I_20596 (I352437,I352540,I352661);
DFFARX1 I_20597 (I9660,I2507,I352463,I352701,);
DFFARX1 I_20598 (I352701,I2507,I352463,I352718,);
not I_20599 (I352726,I352718);
not I_20600 (I352743,I352701);
nand I_20601 (I352440,I352743,I352562);
nand I_20602 (I352774,I9660,I9675);
and I_20603 (I352791,I352774,I9657);
DFFARX1 I_20604 (I352791,I2507,I352463,I352817,);
nor I_20605 (I352825,I352817,I352489);
DFFARX1 I_20606 (I352825,I2507,I352463,I352428,);
DFFARX1 I_20607 (I352817,I2507,I352463,I352446,);
nor I_20608 (I352870,I9678,I9675);
not I_20609 (I352887,I352870);
nor I_20610 (I352449,I352726,I352887);
nand I_20611 (I352434,I352743,I352887);
nor I_20612 (I352443,I352489,I352870);
DFFARX1 I_20613 (I352870,I2507,I352463,I352452,);
not I_20614 (I352990,I2514);
DFFARX1 I_20615 (I96496,I2507,I352990,I353016,);
nand I_20616 (I353024,I96508,I96517);
and I_20617 (I353041,I353024,I96496);
DFFARX1 I_20618 (I353041,I2507,I352990,I353067,);
nor I_20619 (I352958,I353067,I353016);
not I_20620 (I353089,I353067);
DFFARX1 I_20621 (I96511,I2507,I352990,I353115,);
nand I_20622 (I353123,I353115,I96499);
not I_20623 (I353140,I353123);
DFFARX1 I_20624 (I353140,I2507,I352990,I353166,);
not I_20625 (I352982,I353166);
nor I_20626 (I353188,I353016,I353123);
nor I_20627 (I352964,I353067,I353188);
DFFARX1 I_20628 (I96502,I2507,I352990,I353228,);
DFFARX1 I_20629 (I353228,I2507,I352990,I353245,);
not I_20630 (I353253,I353245);
not I_20631 (I353270,I353228);
nand I_20632 (I352967,I353270,I353089);
nand I_20633 (I353301,I96493,I96493);
and I_20634 (I353318,I353301,I96505);
DFFARX1 I_20635 (I353318,I2507,I352990,I353344,);
nor I_20636 (I353352,I353344,I353016);
DFFARX1 I_20637 (I353352,I2507,I352990,I352955,);
DFFARX1 I_20638 (I353344,I2507,I352990,I352973,);
nor I_20639 (I353397,I96514,I96493);
not I_20640 (I353414,I353397);
nor I_20641 (I352976,I353253,I353414);
nand I_20642 (I352961,I353270,I353414);
nor I_20643 (I352970,I353016,I353397);
DFFARX1 I_20644 (I353397,I2507,I352990,I352979,);
not I_20645 (I353517,I2514);
DFFARX1 I_20646 (I54863,I2507,I353517,I353543,);
nand I_20647 (I353551,I54875,I54884);
and I_20648 (I353568,I353551,I54863);
DFFARX1 I_20649 (I353568,I2507,I353517,I353594,);
nor I_20650 (I353485,I353594,I353543);
not I_20651 (I353616,I353594);
DFFARX1 I_20652 (I54878,I2507,I353517,I353642,);
nand I_20653 (I353650,I353642,I54866);
not I_20654 (I353667,I353650);
DFFARX1 I_20655 (I353667,I2507,I353517,I353693,);
not I_20656 (I353509,I353693);
nor I_20657 (I353715,I353543,I353650);
nor I_20658 (I353491,I353594,I353715);
DFFARX1 I_20659 (I54869,I2507,I353517,I353755,);
DFFARX1 I_20660 (I353755,I2507,I353517,I353772,);
not I_20661 (I353780,I353772);
not I_20662 (I353797,I353755);
nand I_20663 (I353494,I353797,I353616);
nand I_20664 (I353828,I54860,I54860);
and I_20665 (I353845,I353828,I54872);
DFFARX1 I_20666 (I353845,I2507,I353517,I353871,);
nor I_20667 (I353879,I353871,I353543);
DFFARX1 I_20668 (I353879,I2507,I353517,I353482,);
DFFARX1 I_20669 (I353871,I2507,I353517,I353500,);
nor I_20670 (I353924,I54881,I54860);
not I_20671 (I353941,I353924);
nor I_20672 (I353503,I353780,I353941);
nand I_20673 (I353488,I353797,I353941);
nor I_20674 (I353497,I353543,I353924);
DFFARX1 I_20675 (I353924,I2507,I353517,I353506,);
not I_20676 (I354044,I2514);
DFFARX1 I_20677 (I146089,I2507,I354044,I354070,);
nand I_20678 (I354078,I146074,I146065);
and I_20679 (I354095,I354078,I146080);
DFFARX1 I_20680 (I354095,I2507,I354044,I354121,);
nor I_20681 (I354012,I354121,I354070);
not I_20682 (I354143,I354121);
DFFARX1 I_20683 (I146092,I2507,I354044,I354169,);
nand I_20684 (I354177,I354169,I146083);
not I_20685 (I354194,I354177);
DFFARX1 I_20686 (I354194,I2507,I354044,I354220,);
not I_20687 (I354036,I354220);
nor I_20688 (I354242,I354070,I354177);
nor I_20689 (I354018,I354121,I354242);
DFFARX1 I_20690 (I146071,I2507,I354044,I354282,);
DFFARX1 I_20691 (I354282,I2507,I354044,I354299,);
not I_20692 (I354307,I354299);
not I_20693 (I354324,I354282);
nand I_20694 (I354021,I354324,I354143);
nand I_20695 (I354355,I146077,I146068);
and I_20696 (I354372,I354355,I146065);
DFFARX1 I_20697 (I354372,I2507,I354044,I354398,);
nor I_20698 (I354406,I354398,I354070);
DFFARX1 I_20699 (I354406,I2507,I354044,I354009,);
DFFARX1 I_20700 (I354398,I2507,I354044,I354027,);
nor I_20701 (I354451,I146086,I146068);
not I_20702 (I354468,I354451);
nor I_20703 (I354030,I354307,I354468);
nand I_20704 (I354015,I354324,I354468);
nor I_20705 (I354024,I354070,I354451);
DFFARX1 I_20706 (I354451,I2507,I354044,I354033,);
not I_20707 (I354571,I2514);
DFFARX1 I_20708 (I451771,I2507,I354571,I354597,);
nand I_20709 (I354605,I451783,I451762);
and I_20710 (I354622,I354605,I451786);
DFFARX1 I_20711 (I354622,I2507,I354571,I354648,);
nor I_20712 (I354539,I354648,I354597);
not I_20713 (I354670,I354648);
DFFARX1 I_20714 (I451777,I2507,I354571,I354696,);
nand I_20715 (I354704,I354696,I451759);
not I_20716 (I354721,I354704);
DFFARX1 I_20717 (I354721,I2507,I354571,I354747,);
not I_20718 (I354563,I354747);
nor I_20719 (I354769,I354597,I354704);
nor I_20720 (I354545,I354648,I354769);
DFFARX1 I_20721 (I451774,I2507,I354571,I354809,);
DFFARX1 I_20722 (I354809,I2507,I354571,I354826,);
not I_20723 (I354834,I354826);
not I_20724 (I354851,I354809);
nand I_20725 (I354548,I354851,I354670);
nand I_20726 (I354882,I451759,I451765);
and I_20727 (I354899,I354882,I451768);
DFFARX1 I_20728 (I354899,I2507,I354571,I354925,);
nor I_20729 (I354933,I354925,I354597);
DFFARX1 I_20730 (I354933,I2507,I354571,I354536,);
DFFARX1 I_20731 (I354925,I2507,I354571,I354554,);
nor I_20732 (I354978,I451780,I451765);
not I_20733 (I354995,I354978);
nor I_20734 (I354557,I354834,I354995);
nand I_20735 (I354542,I354851,I354995);
nor I_20736 (I354551,I354597,I354978);
DFFARX1 I_20737 (I354978,I2507,I354571,I354560,);
not I_20738 (I355098,I2514);
DFFARX1 I_20739 (I526817,I2507,I355098,I355124,);
nand I_20740 (I355132,I526817,I526829);
and I_20741 (I355149,I355132,I526814);
DFFARX1 I_20742 (I355149,I2507,I355098,I355175,);
nor I_20743 (I355066,I355175,I355124);
not I_20744 (I355197,I355175);
DFFARX1 I_20745 (I526838,I2507,I355098,I355223,);
nand I_20746 (I355231,I355223,I526835);
not I_20747 (I355248,I355231);
DFFARX1 I_20748 (I355248,I2507,I355098,I355274,);
not I_20749 (I355090,I355274);
nor I_20750 (I355296,I355124,I355231);
nor I_20751 (I355072,I355175,I355296);
DFFARX1 I_20752 (I526826,I2507,I355098,I355336,);
DFFARX1 I_20753 (I355336,I2507,I355098,I355353,);
not I_20754 (I355361,I355353);
not I_20755 (I355378,I355336);
nand I_20756 (I355075,I355378,I355197);
nand I_20757 (I355409,I526814,I526823);
and I_20758 (I355426,I355409,I526832);
DFFARX1 I_20759 (I355426,I2507,I355098,I355452,);
nor I_20760 (I355460,I355452,I355124);
DFFARX1 I_20761 (I355460,I2507,I355098,I355063,);
DFFARX1 I_20762 (I355452,I2507,I355098,I355081,);
nor I_20763 (I355505,I526820,I526823);
not I_20764 (I355522,I355505);
nor I_20765 (I355084,I355361,I355522);
nand I_20766 (I355069,I355378,I355522);
nor I_20767 (I355078,I355124,I355505);
DFFARX1 I_20768 (I355505,I2507,I355098,I355087,);
not I_20769 (I355625,I2514);
DFFARX1 I_20770 (I768872,I2507,I355625,I355651,);
nand I_20771 (I355659,I768863,I768878);
and I_20772 (I355676,I355659,I768884);
DFFARX1 I_20773 (I355676,I2507,I355625,I355702,);
nor I_20774 (I355593,I355702,I355651);
not I_20775 (I355724,I355702);
DFFARX1 I_20776 (I768869,I2507,I355625,I355750,);
nand I_20777 (I355758,I355750,I768863);
not I_20778 (I355775,I355758);
DFFARX1 I_20779 (I355775,I2507,I355625,I355801,);
not I_20780 (I355617,I355801);
nor I_20781 (I355823,I355651,I355758);
nor I_20782 (I355599,I355702,I355823);
DFFARX1 I_20783 (I768866,I2507,I355625,I355863,);
DFFARX1 I_20784 (I355863,I2507,I355625,I355880,);
not I_20785 (I355888,I355880);
not I_20786 (I355905,I355863);
nand I_20787 (I355602,I355905,I355724);
nand I_20788 (I355936,I768860,I768875);
and I_20789 (I355953,I355936,I768860);
DFFARX1 I_20790 (I355953,I2507,I355625,I355979,);
nor I_20791 (I355987,I355979,I355651);
DFFARX1 I_20792 (I355987,I2507,I355625,I355590,);
DFFARX1 I_20793 (I355979,I2507,I355625,I355608,);
nor I_20794 (I356032,I768881,I768875);
not I_20795 (I356049,I356032);
nor I_20796 (I355611,I355888,I356049);
nand I_20797 (I355596,I355905,I356049);
nor I_20798 (I355605,I355651,I356032);
DFFARX1 I_20799 (I356032,I2507,I355625,I355614,);
not I_20800 (I356152,I2514);
DFFARX1 I_20801 (I1126574,I2507,I356152,I356178,);
nand I_20802 (I356186,I1126589,I1126574);
and I_20803 (I356203,I356186,I1126592);
DFFARX1 I_20804 (I356203,I2507,I356152,I356229,);
nor I_20805 (I356120,I356229,I356178);
not I_20806 (I356251,I356229);
DFFARX1 I_20807 (I1126598,I2507,I356152,I356277,);
nand I_20808 (I356285,I356277,I1126580);
not I_20809 (I356302,I356285);
DFFARX1 I_20810 (I356302,I2507,I356152,I356328,);
not I_20811 (I356144,I356328);
nor I_20812 (I356350,I356178,I356285);
nor I_20813 (I356126,I356229,I356350);
DFFARX1 I_20814 (I1126577,I2507,I356152,I356390,);
DFFARX1 I_20815 (I356390,I2507,I356152,I356407,);
not I_20816 (I356415,I356407);
not I_20817 (I356432,I356390);
nand I_20818 (I356129,I356432,I356251);
nand I_20819 (I356463,I1126577,I1126583);
and I_20820 (I356480,I356463,I1126595);
DFFARX1 I_20821 (I356480,I2507,I356152,I356506,);
nor I_20822 (I356514,I356506,I356178);
DFFARX1 I_20823 (I356514,I2507,I356152,I356117,);
DFFARX1 I_20824 (I356506,I2507,I356152,I356135,);
nor I_20825 (I356559,I1126586,I1126583);
not I_20826 (I356576,I356559);
nor I_20827 (I356138,I356415,I356576);
nand I_20828 (I356123,I356432,I356576);
nor I_20829 (I356132,I356178,I356559);
DFFARX1 I_20830 (I356559,I2507,I356152,I356141,);
not I_20831 (I356679,I2514);
DFFARX1 I_20832 (I1244436,I2507,I356679,I356705,);
nand I_20833 (I356713,I1244418,I1244442);
and I_20834 (I356730,I356713,I1244433);
DFFARX1 I_20835 (I356730,I2507,I356679,I356756,);
nor I_20836 (I356647,I356756,I356705);
not I_20837 (I356778,I356756);
DFFARX1 I_20838 (I1244439,I2507,I356679,I356804,);
nand I_20839 (I356812,I356804,I1244427);
not I_20840 (I356829,I356812);
DFFARX1 I_20841 (I356829,I2507,I356679,I356855,);
not I_20842 (I356671,I356855);
nor I_20843 (I356877,I356705,I356812);
nor I_20844 (I356653,I356756,I356877);
DFFARX1 I_20845 (I1244418,I2507,I356679,I356917,);
DFFARX1 I_20846 (I356917,I2507,I356679,I356934,);
not I_20847 (I356942,I356934);
not I_20848 (I356959,I356917);
nand I_20849 (I356656,I356959,I356778);
nand I_20850 (I356990,I1244424,I1244421);
and I_20851 (I357007,I356990,I1244430);
DFFARX1 I_20852 (I357007,I2507,I356679,I357033,);
nor I_20853 (I357041,I357033,I356705);
DFFARX1 I_20854 (I357041,I2507,I356679,I356644,);
DFFARX1 I_20855 (I357033,I2507,I356679,I356662,);
nor I_20856 (I357086,I1244421,I1244421);
not I_20857 (I357103,I357086);
nor I_20858 (I356665,I356942,I357103);
nand I_20859 (I356650,I356959,I357103);
nor I_20860 (I356659,I356705,I357086);
DFFARX1 I_20861 (I357086,I2507,I356679,I356668,);
not I_20862 (I357206,I2514);
DFFARX1 I_20863 (I89645,I2507,I357206,I357232,);
nand I_20864 (I357240,I89657,I89666);
and I_20865 (I357257,I357240,I89645);
DFFARX1 I_20866 (I357257,I2507,I357206,I357283,);
nor I_20867 (I357174,I357283,I357232);
not I_20868 (I357305,I357283);
DFFARX1 I_20869 (I89660,I2507,I357206,I357331,);
nand I_20870 (I357339,I357331,I89648);
not I_20871 (I357356,I357339);
DFFARX1 I_20872 (I357356,I2507,I357206,I357382,);
not I_20873 (I357198,I357382);
nor I_20874 (I357404,I357232,I357339);
nor I_20875 (I357180,I357283,I357404);
DFFARX1 I_20876 (I89651,I2507,I357206,I357444,);
DFFARX1 I_20877 (I357444,I2507,I357206,I357461,);
not I_20878 (I357469,I357461);
not I_20879 (I357486,I357444);
nand I_20880 (I357183,I357486,I357305);
nand I_20881 (I357517,I89642,I89642);
and I_20882 (I357534,I357517,I89654);
DFFARX1 I_20883 (I357534,I2507,I357206,I357560,);
nor I_20884 (I357568,I357560,I357232);
DFFARX1 I_20885 (I357568,I2507,I357206,I357171,);
DFFARX1 I_20886 (I357560,I2507,I357206,I357189,);
nor I_20887 (I357613,I89663,I89642);
not I_20888 (I357630,I357613);
nor I_20889 (I357192,I357469,I357630);
nand I_20890 (I357177,I357486,I357630);
nor I_20891 (I357186,I357232,I357613);
DFFARX1 I_20892 (I357613,I2507,I357206,I357195,);
not I_20893 (I357733,I2514);
DFFARX1 I_20894 (I458299,I2507,I357733,I357759,);
nand I_20895 (I357767,I458311,I458290);
and I_20896 (I357784,I357767,I458314);
DFFARX1 I_20897 (I357784,I2507,I357733,I357810,);
nor I_20898 (I357701,I357810,I357759);
not I_20899 (I357832,I357810);
DFFARX1 I_20900 (I458305,I2507,I357733,I357858,);
nand I_20901 (I357866,I357858,I458287);
not I_20902 (I357883,I357866);
DFFARX1 I_20903 (I357883,I2507,I357733,I357909,);
not I_20904 (I357725,I357909);
nor I_20905 (I357931,I357759,I357866);
nor I_20906 (I357707,I357810,I357931);
DFFARX1 I_20907 (I458302,I2507,I357733,I357971,);
DFFARX1 I_20908 (I357971,I2507,I357733,I357988,);
not I_20909 (I357996,I357988);
not I_20910 (I358013,I357971);
nand I_20911 (I357710,I358013,I357832);
nand I_20912 (I358044,I458287,I458293);
and I_20913 (I358061,I358044,I458296);
DFFARX1 I_20914 (I358061,I2507,I357733,I358087,);
nor I_20915 (I358095,I358087,I357759);
DFFARX1 I_20916 (I358095,I2507,I357733,I357698,);
DFFARX1 I_20917 (I358087,I2507,I357733,I357716,);
nor I_20918 (I358140,I458308,I458293);
not I_20919 (I358157,I358140);
nor I_20920 (I357719,I357996,I358157);
nand I_20921 (I357704,I358013,I358157);
nor I_20922 (I357713,I357759,I358140);
DFFARX1 I_20923 (I358140,I2507,I357733,I357722,);
not I_20924 (I358260,I2514);
DFFARX1 I_20925 (I156180,I2507,I358260,I358286,);
nand I_20926 (I358294,I156180,I156186);
and I_20927 (I358311,I358294,I156204);
DFFARX1 I_20928 (I358311,I2507,I358260,I358337,);
nor I_20929 (I358228,I358337,I358286);
not I_20930 (I358359,I358337);
DFFARX1 I_20931 (I156192,I2507,I358260,I358385,);
nand I_20932 (I358393,I358385,I156189);
not I_20933 (I358410,I358393);
DFFARX1 I_20934 (I358410,I2507,I358260,I358436,);
not I_20935 (I358252,I358436);
nor I_20936 (I358458,I358286,I358393);
nor I_20937 (I358234,I358337,I358458);
DFFARX1 I_20938 (I156198,I2507,I358260,I358498,);
DFFARX1 I_20939 (I358498,I2507,I358260,I358515,);
not I_20940 (I358523,I358515);
not I_20941 (I358540,I358498);
nand I_20942 (I358237,I358540,I358359);
nand I_20943 (I358571,I156183,I156183);
and I_20944 (I358588,I358571,I156195);
DFFARX1 I_20945 (I358588,I2507,I358260,I358614,);
nor I_20946 (I358622,I358614,I358286);
DFFARX1 I_20947 (I358622,I2507,I358260,I358225,);
DFFARX1 I_20948 (I358614,I2507,I358260,I358243,);
nor I_20949 (I358667,I156201,I156183);
not I_20950 (I358684,I358667);
nor I_20951 (I358246,I358523,I358684);
nand I_20952 (I358231,I358540,I358684);
nor I_20953 (I358240,I358286,I358667);
DFFARX1 I_20954 (I358667,I2507,I358260,I358249,);
not I_20955 (I358787,I2514);
DFFARX1 I_20956 (I190095,I2507,I358787,I358813,);
nand I_20957 (I358821,I190095,I190101);
and I_20958 (I358838,I358821,I190119);
DFFARX1 I_20959 (I358838,I2507,I358787,I358864,);
nor I_20960 (I358755,I358864,I358813);
not I_20961 (I358886,I358864);
DFFARX1 I_20962 (I190107,I2507,I358787,I358912,);
nand I_20963 (I358920,I358912,I190104);
not I_20964 (I358937,I358920);
DFFARX1 I_20965 (I358937,I2507,I358787,I358963,);
not I_20966 (I358779,I358963);
nor I_20967 (I358985,I358813,I358920);
nor I_20968 (I358761,I358864,I358985);
DFFARX1 I_20969 (I190113,I2507,I358787,I359025,);
DFFARX1 I_20970 (I359025,I2507,I358787,I359042,);
not I_20971 (I359050,I359042);
not I_20972 (I359067,I359025);
nand I_20973 (I358764,I359067,I358886);
nand I_20974 (I359098,I190098,I190098);
and I_20975 (I359115,I359098,I190110);
DFFARX1 I_20976 (I359115,I2507,I358787,I359141,);
nor I_20977 (I359149,I359141,I358813);
DFFARX1 I_20978 (I359149,I2507,I358787,I358752,);
DFFARX1 I_20979 (I359141,I2507,I358787,I358770,);
nor I_20980 (I359194,I190116,I190098);
not I_20981 (I359211,I359194);
nor I_20982 (I358773,I359050,I359211);
nand I_20983 (I358758,I359067,I359211);
nor I_20984 (I358767,I358813,I359194);
DFFARX1 I_20985 (I359194,I2507,I358787,I358776,);
not I_20986 (I359314,I2514);
DFFARX1 I_20987 (I1347578,I2507,I359314,I359340,);
nand I_20988 (I359348,I1347557,I1347557);
and I_20989 (I359365,I359348,I1347584);
DFFARX1 I_20990 (I359365,I2507,I359314,I359391,);
nor I_20991 (I359282,I359391,I359340);
not I_20992 (I359413,I359391);
DFFARX1 I_20993 (I1347572,I2507,I359314,I359439,);
nand I_20994 (I359447,I359439,I1347575);
not I_20995 (I359464,I359447);
DFFARX1 I_20996 (I359464,I2507,I359314,I359490,);
not I_20997 (I359306,I359490);
nor I_20998 (I359512,I359340,I359447);
nor I_20999 (I359288,I359391,I359512);
DFFARX1 I_21000 (I1347566,I2507,I359314,I359552,);
DFFARX1 I_21001 (I359552,I2507,I359314,I359569,);
not I_21002 (I359577,I359569);
not I_21003 (I359594,I359552);
nand I_21004 (I359291,I359594,I359413);
nand I_21005 (I359625,I1347563,I1347560);
and I_21006 (I359642,I359625,I1347581);
DFFARX1 I_21007 (I359642,I2507,I359314,I359668,);
nor I_21008 (I359676,I359668,I359340);
DFFARX1 I_21009 (I359676,I2507,I359314,I359279,);
DFFARX1 I_21010 (I359668,I2507,I359314,I359297,);
nor I_21011 (I359721,I1347569,I1347560);
not I_21012 (I359738,I359721);
nor I_21013 (I359300,I359577,I359738);
nand I_21014 (I359285,I359594,I359738);
nor I_21015 (I359294,I359340,I359721);
DFFARX1 I_21016 (I359721,I2507,I359314,I359303,);
not I_21017 (I359841,I2514);
DFFARX1 I_21018 (I431643,I2507,I359841,I359867,);
nand I_21019 (I359875,I431655,I431634);
and I_21020 (I359892,I359875,I431658);
DFFARX1 I_21021 (I359892,I2507,I359841,I359918,);
nor I_21022 (I359809,I359918,I359867);
not I_21023 (I359940,I359918);
DFFARX1 I_21024 (I431649,I2507,I359841,I359966,);
nand I_21025 (I359974,I359966,I431631);
not I_21026 (I359991,I359974);
DFFARX1 I_21027 (I359991,I2507,I359841,I360017,);
not I_21028 (I359833,I360017);
nor I_21029 (I360039,I359867,I359974);
nor I_21030 (I359815,I359918,I360039);
DFFARX1 I_21031 (I431646,I2507,I359841,I360079,);
DFFARX1 I_21032 (I360079,I2507,I359841,I360096,);
not I_21033 (I360104,I360096);
not I_21034 (I360121,I360079);
nand I_21035 (I359818,I360121,I359940);
nand I_21036 (I360152,I431631,I431637);
and I_21037 (I360169,I360152,I431640);
DFFARX1 I_21038 (I360169,I2507,I359841,I360195,);
nor I_21039 (I360203,I360195,I359867);
DFFARX1 I_21040 (I360203,I2507,I359841,I359806,);
DFFARX1 I_21041 (I360195,I2507,I359841,I359824,);
nor I_21042 (I360248,I431652,I431637);
not I_21043 (I360265,I360248);
nor I_21044 (I359827,I360104,I360265);
nand I_21045 (I359812,I360121,I360265);
nor I_21046 (I359821,I359867,I360248);
DFFARX1 I_21047 (I360248,I2507,I359841,I359830,);
not I_21048 (I360368,I2514);
DFFARX1 I_21049 (I70146,I2507,I360368,I360394,);
nand I_21050 (I360402,I70158,I70167);
and I_21051 (I360419,I360402,I70146);
DFFARX1 I_21052 (I360419,I2507,I360368,I360445,);
nor I_21053 (I360336,I360445,I360394);
not I_21054 (I360467,I360445);
DFFARX1 I_21055 (I70161,I2507,I360368,I360493,);
nand I_21056 (I360501,I360493,I70149);
not I_21057 (I360518,I360501);
DFFARX1 I_21058 (I360518,I2507,I360368,I360544,);
not I_21059 (I360360,I360544);
nor I_21060 (I360566,I360394,I360501);
nor I_21061 (I360342,I360445,I360566);
DFFARX1 I_21062 (I70152,I2507,I360368,I360606,);
DFFARX1 I_21063 (I360606,I2507,I360368,I360623,);
not I_21064 (I360631,I360623);
not I_21065 (I360648,I360606);
nand I_21066 (I360345,I360648,I360467);
nand I_21067 (I360679,I70143,I70143);
and I_21068 (I360696,I360679,I70155);
DFFARX1 I_21069 (I360696,I2507,I360368,I360722,);
nor I_21070 (I360730,I360722,I360394);
DFFARX1 I_21071 (I360730,I2507,I360368,I360333,);
DFFARX1 I_21072 (I360722,I2507,I360368,I360351,);
nor I_21073 (I360775,I70164,I70143);
not I_21074 (I360792,I360775);
nor I_21075 (I360354,I360631,I360792);
nand I_21076 (I360339,I360648,I360792);
nor I_21077 (I360348,I360394,I360775);
DFFARX1 I_21078 (I360775,I2507,I360368,I360357,);
not I_21079 (I360895,I2514);
DFFARX1 I_21080 (I75416,I2507,I360895,I360921,);
nand I_21081 (I360929,I75428,I75437);
and I_21082 (I360946,I360929,I75416);
DFFARX1 I_21083 (I360946,I2507,I360895,I360972,);
nor I_21084 (I360863,I360972,I360921);
not I_21085 (I360994,I360972);
DFFARX1 I_21086 (I75431,I2507,I360895,I361020,);
nand I_21087 (I361028,I361020,I75419);
not I_21088 (I361045,I361028);
DFFARX1 I_21089 (I361045,I2507,I360895,I361071,);
not I_21090 (I360887,I361071);
nor I_21091 (I361093,I360921,I361028);
nor I_21092 (I360869,I360972,I361093);
DFFARX1 I_21093 (I75422,I2507,I360895,I361133,);
DFFARX1 I_21094 (I361133,I2507,I360895,I361150,);
not I_21095 (I361158,I361150);
not I_21096 (I361175,I361133);
nand I_21097 (I360872,I361175,I360994);
nand I_21098 (I361206,I75413,I75413);
and I_21099 (I361223,I361206,I75425);
DFFARX1 I_21100 (I361223,I2507,I360895,I361249,);
nor I_21101 (I361257,I361249,I360921);
DFFARX1 I_21102 (I361257,I2507,I360895,I360860,);
DFFARX1 I_21103 (I361249,I2507,I360895,I360878,);
nor I_21104 (I361302,I75434,I75413);
not I_21105 (I361319,I361302);
nor I_21106 (I360881,I361158,I361319);
nand I_21107 (I360866,I361175,I361319);
nor I_21108 (I360875,I360921,I361302);
DFFARX1 I_21109 (I361302,I2507,I360895,I360884,);
not I_21110 (I361422,I2514);
DFFARX1 I_21111 (I745174,I2507,I361422,I361448,);
nand I_21112 (I361456,I745165,I745180);
and I_21113 (I361473,I361456,I745186);
DFFARX1 I_21114 (I361473,I2507,I361422,I361499,);
nor I_21115 (I361390,I361499,I361448);
not I_21116 (I361521,I361499);
DFFARX1 I_21117 (I745171,I2507,I361422,I361547,);
nand I_21118 (I361555,I361547,I745165);
not I_21119 (I361572,I361555);
DFFARX1 I_21120 (I361572,I2507,I361422,I361598,);
not I_21121 (I361414,I361598);
nor I_21122 (I361620,I361448,I361555);
nor I_21123 (I361396,I361499,I361620);
DFFARX1 I_21124 (I745168,I2507,I361422,I361660,);
DFFARX1 I_21125 (I361660,I2507,I361422,I361677,);
not I_21126 (I361685,I361677);
not I_21127 (I361702,I361660);
nand I_21128 (I361399,I361702,I361521);
nand I_21129 (I361733,I745162,I745177);
and I_21130 (I361750,I361733,I745162);
DFFARX1 I_21131 (I361750,I2507,I361422,I361776,);
nor I_21132 (I361784,I361776,I361448);
DFFARX1 I_21133 (I361784,I2507,I361422,I361387,);
DFFARX1 I_21134 (I361776,I2507,I361422,I361405,);
nor I_21135 (I361829,I745183,I745177);
not I_21136 (I361846,I361829);
nor I_21137 (I361408,I361685,I361846);
nand I_21138 (I361393,I361702,I361846);
nor I_21139 (I361402,I361448,I361829);
DFFARX1 I_21140 (I361829,I2507,I361422,I361411,);
not I_21141 (I361949,I2514);
DFFARX1 I_21142 (I941192,I2507,I361949,I361975,);
nand I_21143 (I361983,I941189,I941207);
and I_21144 (I362000,I361983,I941198);
DFFARX1 I_21145 (I362000,I2507,I361949,I362026,);
nor I_21146 (I361917,I362026,I361975);
not I_21147 (I362048,I362026);
DFFARX1 I_21148 (I941213,I2507,I361949,I362074,);
nand I_21149 (I362082,I362074,I941195);
not I_21150 (I362099,I362082);
DFFARX1 I_21151 (I362099,I2507,I361949,I362125,);
not I_21152 (I361941,I362125);
nor I_21153 (I362147,I361975,I362082);
nor I_21154 (I361923,I362026,I362147);
DFFARX1 I_21155 (I941201,I2507,I361949,I362187,);
DFFARX1 I_21156 (I362187,I2507,I361949,I362204,);
not I_21157 (I362212,I362204);
not I_21158 (I362229,I362187);
nand I_21159 (I361926,I362229,I362048);
nand I_21160 (I362260,I941189,I941216);
and I_21161 (I362277,I362260,I941204);
DFFARX1 I_21162 (I362277,I2507,I361949,I362303,);
nor I_21163 (I362311,I362303,I361975);
DFFARX1 I_21164 (I362311,I2507,I361949,I361914,);
DFFARX1 I_21165 (I362303,I2507,I361949,I361932,);
nor I_21166 (I362356,I941210,I941216);
not I_21167 (I362373,I362356);
nor I_21168 (I361935,I362212,I362373);
nand I_21169 (I361920,I362229,I362373);
nor I_21170 (I361929,I361975,I362356);
DFFARX1 I_21171 (I362356,I2507,I361949,I361938,);
not I_21172 (I362476,I2514);
DFFARX1 I_21173 (I749798,I2507,I362476,I362502,);
nand I_21174 (I362510,I749789,I749804);
and I_21175 (I362527,I362510,I749810);
DFFARX1 I_21176 (I362527,I2507,I362476,I362553,);
nor I_21177 (I362444,I362553,I362502);
not I_21178 (I362575,I362553);
DFFARX1 I_21179 (I749795,I2507,I362476,I362601,);
nand I_21180 (I362609,I362601,I749789);
not I_21181 (I362626,I362609);
DFFARX1 I_21182 (I362626,I2507,I362476,I362652,);
not I_21183 (I362468,I362652);
nor I_21184 (I362674,I362502,I362609);
nor I_21185 (I362450,I362553,I362674);
DFFARX1 I_21186 (I749792,I2507,I362476,I362714,);
DFFARX1 I_21187 (I362714,I2507,I362476,I362731,);
not I_21188 (I362739,I362731);
not I_21189 (I362756,I362714);
nand I_21190 (I362453,I362756,I362575);
nand I_21191 (I362787,I749786,I749801);
and I_21192 (I362804,I362787,I749786);
DFFARX1 I_21193 (I362804,I2507,I362476,I362830,);
nor I_21194 (I362838,I362830,I362502);
DFFARX1 I_21195 (I362838,I2507,I362476,I362441,);
DFFARX1 I_21196 (I362830,I2507,I362476,I362459,);
nor I_21197 (I362883,I749807,I749801);
not I_21198 (I362900,I362883);
nor I_21199 (I362462,I362739,I362900);
nand I_21200 (I362447,I362756,I362900);
nor I_21201 (I362456,I362502,I362883);
DFFARX1 I_21202 (I362883,I2507,I362476,I362465,);
not I_21203 (I363003,I2514);
DFFARX1 I_21204 (I548079,I2507,I363003,I363029,);
nand I_21205 (I363037,I548064,I548067);
and I_21206 (I363054,I363037,I548082);
DFFARX1 I_21207 (I363054,I2507,I363003,I363080,);
nor I_21208 (I362971,I363080,I363029);
not I_21209 (I363102,I363080);
DFFARX1 I_21210 (I548076,I2507,I363003,I363128,);
nand I_21211 (I363136,I363128,I548067);
not I_21212 (I363153,I363136);
DFFARX1 I_21213 (I363153,I2507,I363003,I363179,);
not I_21214 (I362995,I363179);
nor I_21215 (I363201,I363029,I363136);
nor I_21216 (I362977,I363080,I363201);
DFFARX1 I_21217 (I548073,I2507,I363003,I363241,);
DFFARX1 I_21218 (I363241,I2507,I363003,I363258,);
not I_21219 (I363266,I363258);
not I_21220 (I363283,I363241);
nand I_21221 (I362980,I363283,I363102);
nand I_21222 (I363314,I548088,I548064);
and I_21223 (I363331,I363314,I548085);
DFFARX1 I_21224 (I363331,I2507,I363003,I363357,);
nor I_21225 (I363365,I363357,I363029);
DFFARX1 I_21226 (I363365,I2507,I363003,I362968,);
DFFARX1 I_21227 (I363357,I2507,I363003,I362986,);
nor I_21228 (I363410,I548070,I548064);
not I_21229 (I363427,I363410);
nor I_21230 (I362989,I363266,I363427);
nand I_21231 (I362974,I363283,I363427);
nor I_21232 (I362983,I363029,I363410);
DFFARX1 I_21233 (I363410,I2507,I363003,I362992,);
not I_21234 (I363530,I2514);
DFFARX1 I_21235 (I1108656,I2507,I363530,I363556,);
nand I_21236 (I363564,I1108671,I1108656);
and I_21237 (I363581,I363564,I1108674);
DFFARX1 I_21238 (I363581,I2507,I363530,I363607,);
nor I_21239 (I363498,I363607,I363556);
not I_21240 (I363629,I363607);
DFFARX1 I_21241 (I1108680,I2507,I363530,I363655,);
nand I_21242 (I363663,I363655,I1108662);
not I_21243 (I363680,I363663);
DFFARX1 I_21244 (I363680,I2507,I363530,I363706,);
not I_21245 (I363522,I363706);
nor I_21246 (I363728,I363556,I363663);
nor I_21247 (I363504,I363607,I363728);
DFFARX1 I_21248 (I1108659,I2507,I363530,I363768,);
DFFARX1 I_21249 (I363768,I2507,I363530,I363785,);
not I_21250 (I363793,I363785);
not I_21251 (I363810,I363768);
nand I_21252 (I363507,I363810,I363629);
nand I_21253 (I363841,I1108659,I1108665);
and I_21254 (I363858,I363841,I1108677);
DFFARX1 I_21255 (I363858,I2507,I363530,I363884,);
nor I_21256 (I363892,I363884,I363556);
DFFARX1 I_21257 (I363892,I2507,I363530,I363495,);
DFFARX1 I_21258 (I363884,I2507,I363530,I363513,);
nor I_21259 (I363937,I1108668,I1108665);
not I_21260 (I363954,I363937);
nor I_21261 (I363516,I363793,I363954);
nand I_21262 (I363501,I363810,I363954);
nor I_21263 (I363510,I363556,I363937);
DFFARX1 I_21264 (I363937,I2507,I363530,I363519,);
not I_21265 (I364057,I2514);
DFFARX1 I_21266 (I1062416,I2507,I364057,I364083,);
nand I_21267 (I364091,I1062431,I1062416);
and I_21268 (I364108,I364091,I1062434);
DFFARX1 I_21269 (I364108,I2507,I364057,I364134,);
nor I_21270 (I364025,I364134,I364083);
not I_21271 (I364156,I364134);
DFFARX1 I_21272 (I1062440,I2507,I364057,I364182,);
nand I_21273 (I364190,I364182,I1062422);
not I_21274 (I364207,I364190);
DFFARX1 I_21275 (I364207,I2507,I364057,I364233,);
not I_21276 (I364049,I364233);
nor I_21277 (I364255,I364083,I364190);
nor I_21278 (I364031,I364134,I364255);
DFFARX1 I_21279 (I1062419,I2507,I364057,I364295,);
DFFARX1 I_21280 (I364295,I2507,I364057,I364312,);
not I_21281 (I364320,I364312);
not I_21282 (I364337,I364295);
nand I_21283 (I364034,I364337,I364156);
nand I_21284 (I364368,I1062419,I1062425);
and I_21285 (I364385,I364368,I1062437);
DFFARX1 I_21286 (I364385,I2507,I364057,I364411,);
nor I_21287 (I364419,I364411,I364083);
DFFARX1 I_21288 (I364419,I2507,I364057,I364022,);
DFFARX1 I_21289 (I364411,I2507,I364057,I364040,);
nor I_21290 (I364464,I1062428,I1062425);
not I_21291 (I364481,I364464);
nor I_21292 (I364043,I364320,I364481);
nand I_21293 (I364028,I364337,I364481);
nor I_21294 (I364037,I364083,I364464);
DFFARX1 I_21295 (I364464,I2507,I364057,I364046,);
not I_21296 (I364584,I2514);
DFFARX1 I_21297 (I163915,I2507,I364584,I364610,);
nand I_21298 (I364618,I163915,I163921);
and I_21299 (I364635,I364618,I163939);
DFFARX1 I_21300 (I364635,I2507,I364584,I364661,);
nor I_21301 (I364552,I364661,I364610);
not I_21302 (I364683,I364661);
DFFARX1 I_21303 (I163927,I2507,I364584,I364709,);
nand I_21304 (I364717,I364709,I163924);
not I_21305 (I364734,I364717);
DFFARX1 I_21306 (I364734,I2507,I364584,I364760,);
not I_21307 (I364576,I364760);
nor I_21308 (I364782,I364610,I364717);
nor I_21309 (I364558,I364661,I364782);
DFFARX1 I_21310 (I163933,I2507,I364584,I364822,);
DFFARX1 I_21311 (I364822,I2507,I364584,I364839,);
not I_21312 (I364847,I364839);
not I_21313 (I364864,I364822);
nand I_21314 (I364561,I364864,I364683);
nand I_21315 (I364895,I163918,I163918);
and I_21316 (I364912,I364895,I163930);
DFFARX1 I_21317 (I364912,I2507,I364584,I364938,);
nor I_21318 (I364946,I364938,I364610);
DFFARX1 I_21319 (I364946,I2507,I364584,I364549,);
DFFARX1 I_21320 (I364938,I2507,I364584,I364567,);
nor I_21321 (I364991,I163936,I163918);
not I_21322 (I365008,I364991);
nor I_21323 (I364570,I364847,I365008);
nand I_21324 (I364555,I364864,I365008);
nor I_21325 (I364564,I364610,I364991);
DFFARX1 I_21326 (I364991,I2507,I364584,I364573,);
not I_21327 (I365111,I2514);
DFFARX1 I_21328 (I1386848,I2507,I365111,I365137,);
nand I_21329 (I365145,I1386827,I1386827);
and I_21330 (I365162,I365145,I1386854);
DFFARX1 I_21331 (I365162,I2507,I365111,I365188,);
nor I_21332 (I365079,I365188,I365137);
not I_21333 (I365210,I365188);
DFFARX1 I_21334 (I1386842,I2507,I365111,I365236,);
nand I_21335 (I365244,I365236,I1386845);
not I_21336 (I365261,I365244);
DFFARX1 I_21337 (I365261,I2507,I365111,I365287,);
not I_21338 (I365103,I365287);
nor I_21339 (I365309,I365137,I365244);
nor I_21340 (I365085,I365188,I365309);
DFFARX1 I_21341 (I1386836,I2507,I365111,I365349,);
DFFARX1 I_21342 (I365349,I2507,I365111,I365366,);
not I_21343 (I365374,I365366);
not I_21344 (I365391,I365349);
nand I_21345 (I365088,I365391,I365210);
nand I_21346 (I365422,I1386833,I1386830);
and I_21347 (I365439,I365422,I1386851);
DFFARX1 I_21348 (I365439,I2507,I365111,I365465,);
nor I_21349 (I365473,I365465,I365137);
DFFARX1 I_21350 (I365473,I2507,I365111,I365076,);
DFFARX1 I_21351 (I365465,I2507,I365111,I365094,);
nor I_21352 (I365518,I1386839,I1386830);
not I_21353 (I365535,I365518);
nor I_21354 (I365097,I365374,I365535);
nand I_21355 (I365082,I365391,I365535);
nor I_21356 (I365091,I365137,I365518);
DFFARX1 I_21357 (I365518,I2507,I365111,I365100,);
not I_21358 (I365638,I2514);
DFFARX1 I_21359 (I644602,I2507,I365638,I365664,);
nand I_21360 (I365672,I644593,I644608);
and I_21361 (I365689,I365672,I644614);
DFFARX1 I_21362 (I365689,I2507,I365638,I365715,);
nor I_21363 (I365606,I365715,I365664);
not I_21364 (I365737,I365715);
DFFARX1 I_21365 (I644599,I2507,I365638,I365763,);
nand I_21366 (I365771,I365763,I644593);
not I_21367 (I365788,I365771);
DFFARX1 I_21368 (I365788,I2507,I365638,I365814,);
not I_21369 (I365630,I365814);
nor I_21370 (I365836,I365664,I365771);
nor I_21371 (I365612,I365715,I365836);
DFFARX1 I_21372 (I644596,I2507,I365638,I365876,);
DFFARX1 I_21373 (I365876,I2507,I365638,I365893,);
not I_21374 (I365901,I365893);
not I_21375 (I365918,I365876);
nand I_21376 (I365615,I365918,I365737);
nand I_21377 (I365949,I644590,I644605);
and I_21378 (I365966,I365949,I644590);
DFFARX1 I_21379 (I365966,I2507,I365638,I365992,);
nor I_21380 (I366000,I365992,I365664);
DFFARX1 I_21381 (I366000,I2507,I365638,I365603,);
DFFARX1 I_21382 (I365992,I2507,I365638,I365621,);
nor I_21383 (I366045,I644611,I644605);
not I_21384 (I366062,I366045);
nor I_21385 (I365624,I365901,I366062);
nand I_21386 (I365609,I365918,I366062);
nor I_21387 (I365618,I365664,I366045);
DFFARX1 I_21388 (I366045,I2507,I365638,I365627,);
not I_21389 (I366165,I2514);
DFFARX1 I_21390 (I1184952,I2507,I366165,I366191,);
nand I_21391 (I366199,I1184967,I1184952);
and I_21392 (I366216,I366199,I1184970);
DFFARX1 I_21393 (I366216,I2507,I366165,I366242,);
nor I_21394 (I366133,I366242,I366191);
not I_21395 (I366264,I366242);
DFFARX1 I_21396 (I1184976,I2507,I366165,I366290,);
nand I_21397 (I366298,I366290,I1184958);
not I_21398 (I366315,I366298);
DFFARX1 I_21399 (I366315,I2507,I366165,I366341,);
not I_21400 (I366157,I366341);
nor I_21401 (I366363,I366191,I366298);
nor I_21402 (I366139,I366242,I366363);
DFFARX1 I_21403 (I1184955,I2507,I366165,I366403,);
DFFARX1 I_21404 (I366403,I2507,I366165,I366420,);
not I_21405 (I366428,I366420);
not I_21406 (I366445,I366403);
nand I_21407 (I366142,I366445,I366264);
nand I_21408 (I366476,I1184955,I1184961);
and I_21409 (I366493,I366476,I1184973);
DFFARX1 I_21410 (I366493,I2507,I366165,I366519,);
nor I_21411 (I366527,I366519,I366191);
DFFARX1 I_21412 (I366527,I2507,I366165,I366130,);
DFFARX1 I_21413 (I366519,I2507,I366165,I366148,);
nor I_21414 (I366572,I1184964,I1184961);
not I_21415 (I366589,I366572);
nor I_21416 (I366151,I366428,I366589);
nand I_21417 (I366136,I366445,I366589);
nor I_21418 (I366145,I366191,I366572);
DFFARX1 I_21419 (I366572,I2507,I366165,I366154,);
not I_21420 (I366692,I2514);
DFFARX1 I_21421 (I1208532,I2507,I366692,I366718,);
nand I_21422 (I366726,I1208514,I1208538);
and I_21423 (I366743,I366726,I1208529);
DFFARX1 I_21424 (I366743,I2507,I366692,I366769,);
nor I_21425 (I366660,I366769,I366718);
not I_21426 (I366791,I366769);
DFFARX1 I_21427 (I1208535,I2507,I366692,I366817,);
nand I_21428 (I366825,I366817,I1208523);
not I_21429 (I366842,I366825);
DFFARX1 I_21430 (I366842,I2507,I366692,I366868,);
not I_21431 (I366684,I366868);
nor I_21432 (I366890,I366718,I366825);
nor I_21433 (I366666,I366769,I366890);
DFFARX1 I_21434 (I1208514,I2507,I366692,I366930,);
DFFARX1 I_21435 (I366930,I2507,I366692,I366947,);
not I_21436 (I366955,I366947);
not I_21437 (I366972,I366930);
nand I_21438 (I366669,I366972,I366791);
nand I_21439 (I367003,I1208520,I1208517);
and I_21440 (I367020,I367003,I1208526);
DFFARX1 I_21441 (I367020,I2507,I366692,I367046,);
nor I_21442 (I367054,I367046,I366718);
DFFARX1 I_21443 (I367054,I2507,I366692,I366657,);
DFFARX1 I_21444 (I367046,I2507,I366692,I366675,);
nor I_21445 (I367099,I1208517,I1208517);
not I_21446 (I367116,I367099);
nor I_21447 (I366678,I366955,I367116);
nand I_21448 (I366663,I366972,I367116);
nor I_21449 (I366672,I366718,I367099);
DFFARX1 I_21450 (I367099,I2507,I366692,I366681,);
not I_21451 (I367219,I2514);
DFFARX1 I_21452 (I1195356,I2507,I367219,I367245,);
nand I_21453 (I367253,I1195371,I1195356);
and I_21454 (I367270,I367253,I1195374);
DFFARX1 I_21455 (I367270,I2507,I367219,I367296,);
nor I_21456 (I367187,I367296,I367245);
not I_21457 (I367318,I367296);
DFFARX1 I_21458 (I1195380,I2507,I367219,I367344,);
nand I_21459 (I367352,I367344,I1195362);
not I_21460 (I367369,I367352);
DFFARX1 I_21461 (I367369,I2507,I367219,I367395,);
not I_21462 (I367211,I367395);
nor I_21463 (I367417,I367245,I367352);
nor I_21464 (I367193,I367296,I367417);
DFFARX1 I_21465 (I1195359,I2507,I367219,I367457,);
DFFARX1 I_21466 (I367457,I2507,I367219,I367474,);
not I_21467 (I367482,I367474);
not I_21468 (I367499,I367457);
nand I_21469 (I367196,I367499,I367318);
nand I_21470 (I367530,I1195359,I1195365);
and I_21471 (I367547,I367530,I1195377);
DFFARX1 I_21472 (I367547,I2507,I367219,I367573,);
nor I_21473 (I367581,I367573,I367245);
DFFARX1 I_21474 (I367581,I2507,I367219,I367184,);
DFFARX1 I_21475 (I367573,I2507,I367219,I367202,);
nor I_21476 (I367626,I1195368,I1195365);
not I_21477 (I367643,I367626);
nor I_21478 (I367205,I367482,I367643);
nand I_21479 (I367190,I367499,I367643);
nor I_21480 (I367199,I367245,I367626);
DFFARX1 I_21481 (I367626,I2507,I367219,I367208,);
not I_21482 (I367746,I2514);
DFFARX1 I_21483 (I770606,I2507,I367746,I367772,);
nand I_21484 (I367780,I770597,I770612);
and I_21485 (I367797,I367780,I770618);
DFFARX1 I_21486 (I367797,I2507,I367746,I367823,);
nor I_21487 (I367714,I367823,I367772);
not I_21488 (I367845,I367823);
DFFARX1 I_21489 (I770603,I2507,I367746,I367871,);
nand I_21490 (I367879,I367871,I770597);
not I_21491 (I367896,I367879);
DFFARX1 I_21492 (I367896,I2507,I367746,I367922,);
not I_21493 (I367738,I367922);
nor I_21494 (I367944,I367772,I367879);
nor I_21495 (I367720,I367823,I367944);
DFFARX1 I_21496 (I770600,I2507,I367746,I367984,);
DFFARX1 I_21497 (I367984,I2507,I367746,I368001,);
not I_21498 (I368009,I368001);
not I_21499 (I368026,I367984);
nand I_21500 (I367723,I368026,I367845);
nand I_21501 (I368057,I770594,I770609);
and I_21502 (I368074,I368057,I770594);
DFFARX1 I_21503 (I368074,I2507,I367746,I368100,);
nor I_21504 (I368108,I368100,I367772);
DFFARX1 I_21505 (I368108,I2507,I367746,I367711,);
DFFARX1 I_21506 (I368100,I2507,I367746,I367729,);
nor I_21507 (I368153,I770615,I770609);
not I_21508 (I368170,I368153);
nor I_21509 (I367732,I368009,I368170);
nand I_21510 (I367717,I368026,I368170);
nor I_21511 (I367726,I367772,I368153);
DFFARX1 I_21512 (I368153,I2507,I367746,I367735,);
not I_21513 (I368273,I2514);
DFFARX1 I_21514 (I1123106,I2507,I368273,I368299,);
nand I_21515 (I368307,I1123121,I1123106);
and I_21516 (I368324,I368307,I1123124);
DFFARX1 I_21517 (I368324,I2507,I368273,I368350,);
nor I_21518 (I368241,I368350,I368299);
not I_21519 (I368372,I368350);
DFFARX1 I_21520 (I1123130,I2507,I368273,I368398,);
nand I_21521 (I368406,I368398,I1123112);
not I_21522 (I368423,I368406);
DFFARX1 I_21523 (I368423,I2507,I368273,I368449,);
not I_21524 (I368265,I368449);
nor I_21525 (I368471,I368299,I368406);
nor I_21526 (I368247,I368350,I368471);
DFFARX1 I_21527 (I1123109,I2507,I368273,I368511,);
DFFARX1 I_21528 (I368511,I2507,I368273,I368528,);
not I_21529 (I368536,I368528);
not I_21530 (I368553,I368511);
nand I_21531 (I368250,I368553,I368372);
nand I_21532 (I368584,I1123109,I1123115);
and I_21533 (I368601,I368584,I1123127);
DFFARX1 I_21534 (I368601,I2507,I368273,I368627,);
nor I_21535 (I368635,I368627,I368299);
DFFARX1 I_21536 (I368635,I2507,I368273,I368238,);
DFFARX1 I_21537 (I368627,I2507,I368273,I368256,);
nor I_21538 (I368680,I1123118,I1123115);
not I_21539 (I368697,I368680);
nor I_21540 (I368259,I368536,I368697);
nand I_21541 (I368244,I368553,I368697);
nor I_21542 (I368253,I368299,I368680);
DFFARX1 I_21543 (I368680,I2507,I368273,I368262,);
not I_21544 (I368800,I2514);
DFFARX1 I_21545 (I875504,I2507,I368800,I368826,);
nand I_21546 (I368834,I875507,I875501);
and I_21547 (I368851,I368834,I875513);
DFFARX1 I_21548 (I368851,I2507,I368800,I368877,);
nor I_21549 (I368768,I368877,I368826);
not I_21550 (I368899,I368877);
DFFARX1 I_21551 (I875516,I2507,I368800,I368925,);
nand I_21552 (I368933,I368925,I875507);
not I_21553 (I368950,I368933);
DFFARX1 I_21554 (I368950,I2507,I368800,I368976,);
not I_21555 (I368792,I368976);
nor I_21556 (I368998,I368826,I368933);
nor I_21557 (I368774,I368877,I368998);
DFFARX1 I_21558 (I875519,I2507,I368800,I369038,);
DFFARX1 I_21559 (I369038,I2507,I368800,I369055,);
not I_21560 (I369063,I369055);
not I_21561 (I369080,I369038);
nand I_21562 (I368777,I369080,I368899);
nand I_21563 (I369111,I875501,I875510);
and I_21564 (I369128,I369111,I875504);
DFFARX1 I_21565 (I369128,I2507,I368800,I369154,);
nor I_21566 (I369162,I369154,I368826);
DFFARX1 I_21567 (I369162,I2507,I368800,I368765,);
DFFARX1 I_21568 (I369154,I2507,I368800,I368783,);
nor I_21569 (I369207,I875522,I875510);
not I_21570 (I369224,I369207);
nor I_21571 (I368786,I369063,I369224);
nand I_21572 (I368771,I369080,I369224);
nor I_21573 (I368780,I368826,I369207);
DFFARX1 I_21574 (I369207,I2507,I368800,I368789,);
not I_21575 (I369327,I2514);
DFFARX1 I_21576 (I169270,I2507,I369327,I369353,);
nand I_21577 (I369361,I169270,I169276);
and I_21578 (I369378,I369361,I169294);
DFFARX1 I_21579 (I369378,I2507,I369327,I369404,);
nor I_21580 (I369295,I369404,I369353);
not I_21581 (I369426,I369404);
DFFARX1 I_21582 (I169282,I2507,I369327,I369452,);
nand I_21583 (I369460,I369452,I169279);
not I_21584 (I369477,I369460);
DFFARX1 I_21585 (I369477,I2507,I369327,I369503,);
not I_21586 (I369319,I369503);
nor I_21587 (I369525,I369353,I369460);
nor I_21588 (I369301,I369404,I369525);
DFFARX1 I_21589 (I169288,I2507,I369327,I369565,);
DFFARX1 I_21590 (I369565,I2507,I369327,I369582,);
not I_21591 (I369590,I369582);
not I_21592 (I369607,I369565);
nand I_21593 (I369304,I369607,I369426);
nand I_21594 (I369638,I169273,I169273);
and I_21595 (I369655,I369638,I169285);
DFFARX1 I_21596 (I369655,I2507,I369327,I369681,);
nor I_21597 (I369689,I369681,I369353);
DFFARX1 I_21598 (I369689,I2507,I369327,I369292,);
DFFARX1 I_21599 (I369681,I2507,I369327,I369310,);
nor I_21600 (I369734,I169291,I169273);
not I_21601 (I369751,I369734);
nor I_21602 (I369313,I369590,I369751);
nand I_21603 (I369298,I369607,I369751);
nor I_21604 (I369307,I369353,I369734);
DFFARX1 I_21605 (I369734,I2507,I369327,I369316,);
not I_21606 (I369854,I2514);
DFFARX1 I_21607 (I1069930,I2507,I369854,I369880,);
nand I_21608 (I369888,I1069945,I1069930);
and I_21609 (I369905,I369888,I1069948);
DFFARX1 I_21610 (I369905,I2507,I369854,I369931,);
nor I_21611 (I369822,I369931,I369880);
not I_21612 (I369953,I369931);
DFFARX1 I_21613 (I1069954,I2507,I369854,I369979,);
nand I_21614 (I369987,I369979,I1069936);
not I_21615 (I370004,I369987);
DFFARX1 I_21616 (I370004,I2507,I369854,I370030,);
not I_21617 (I369846,I370030);
nor I_21618 (I370052,I369880,I369987);
nor I_21619 (I369828,I369931,I370052);
DFFARX1 I_21620 (I1069933,I2507,I369854,I370092,);
DFFARX1 I_21621 (I370092,I2507,I369854,I370109,);
not I_21622 (I370117,I370109);
not I_21623 (I370134,I370092);
nand I_21624 (I369831,I370134,I369953);
nand I_21625 (I370165,I1069933,I1069939);
and I_21626 (I370182,I370165,I1069951);
DFFARX1 I_21627 (I370182,I2507,I369854,I370208,);
nor I_21628 (I370216,I370208,I369880);
DFFARX1 I_21629 (I370216,I2507,I369854,I369819,);
DFFARX1 I_21630 (I370208,I2507,I369854,I369837,);
nor I_21631 (I370261,I1069942,I1069939);
not I_21632 (I370278,I370261);
nor I_21633 (I369840,I370117,I370278);
nand I_21634 (I369825,I370134,I370278);
nor I_21635 (I369834,I369880,I370261);
DFFARX1 I_21636 (I370261,I2507,I369854,I369843,);
not I_21637 (I370381,I2514);
DFFARX1 I_21638 (I1055024,I2507,I370381,I370407,);
nand I_21639 (I370415,I1055021,I1055024);
and I_21640 (I370432,I370415,I1055033);
DFFARX1 I_21641 (I370432,I2507,I370381,I370458,);
nor I_21642 (I370349,I370458,I370407);
not I_21643 (I370480,I370458);
DFFARX1 I_21644 (I1055021,I2507,I370381,I370506,);
nand I_21645 (I370514,I370506,I1055039);
not I_21646 (I370531,I370514);
DFFARX1 I_21647 (I370531,I2507,I370381,I370557,);
not I_21648 (I370373,I370557);
nor I_21649 (I370579,I370407,I370514);
nor I_21650 (I370355,I370458,I370579);
DFFARX1 I_21651 (I1055027,I2507,I370381,I370619,);
DFFARX1 I_21652 (I370619,I2507,I370381,I370636,);
not I_21653 (I370644,I370636);
not I_21654 (I370661,I370619);
nand I_21655 (I370358,I370661,I370480);
nand I_21656 (I370692,I1055036,I1055042);
and I_21657 (I370709,I370692,I1055027);
DFFARX1 I_21658 (I370709,I2507,I370381,I370735,);
nor I_21659 (I370743,I370735,I370407);
DFFARX1 I_21660 (I370743,I2507,I370381,I370346,);
DFFARX1 I_21661 (I370735,I2507,I370381,I370364,);
nor I_21662 (I370788,I1055030,I1055042);
not I_21663 (I370805,I370788);
nor I_21664 (I370367,I370644,I370805);
nand I_21665 (I370352,I370661,I370805);
nor I_21666 (I370361,I370407,I370788);
DFFARX1 I_21667 (I370788,I2507,I370381,I370370,);
not I_21668 (I370908,I2514);
DFFARX1 I_21669 (I627840,I2507,I370908,I370934,);
nand I_21670 (I370942,I627831,I627846);
and I_21671 (I370959,I370942,I627852);
DFFARX1 I_21672 (I370959,I2507,I370908,I370985,);
nor I_21673 (I370876,I370985,I370934);
not I_21674 (I371007,I370985);
DFFARX1 I_21675 (I627837,I2507,I370908,I371033,);
nand I_21676 (I371041,I371033,I627831);
not I_21677 (I371058,I371041);
DFFARX1 I_21678 (I371058,I2507,I370908,I371084,);
not I_21679 (I370900,I371084);
nor I_21680 (I371106,I370934,I371041);
nor I_21681 (I370882,I370985,I371106);
DFFARX1 I_21682 (I627834,I2507,I370908,I371146,);
DFFARX1 I_21683 (I371146,I2507,I370908,I371163,);
not I_21684 (I371171,I371163);
not I_21685 (I371188,I371146);
nand I_21686 (I370885,I371188,I371007);
nand I_21687 (I371219,I627828,I627843);
and I_21688 (I371236,I371219,I627828);
DFFARX1 I_21689 (I371236,I2507,I370908,I371262,);
nor I_21690 (I371270,I371262,I370934);
DFFARX1 I_21691 (I371270,I2507,I370908,I370873,);
DFFARX1 I_21692 (I371262,I2507,I370908,I370891,);
nor I_21693 (I371315,I627849,I627843);
not I_21694 (I371332,I371315);
nor I_21695 (I370894,I371171,I371332);
nand I_21696 (I370879,I371188,I371332);
nor I_21697 (I370888,I370934,I371315);
DFFARX1 I_21698 (I371315,I2507,I370908,I370897,);
not I_21699 (I371435,I2514);
DFFARX1 I_21700 (I1198246,I2507,I371435,I371461,);
nand I_21701 (I371469,I1198261,I1198246);
and I_21702 (I371486,I371469,I1198264);
DFFARX1 I_21703 (I371486,I2507,I371435,I371512,);
nor I_21704 (I371403,I371512,I371461);
not I_21705 (I371534,I371512);
DFFARX1 I_21706 (I1198270,I2507,I371435,I371560,);
nand I_21707 (I371568,I371560,I1198252);
not I_21708 (I371585,I371568);
DFFARX1 I_21709 (I371585,I2507,I371435,I371611,);
not I_21710 (I371427,I371611);
nor I_21711 (I371633,I371461,I371568);
nor I_21712 (I371409,I371512,I371633);
DFFARX1 I_21713 (I1198249,I2507,I371435,I371673,);
DFFARX1 I_21714 (I371673,I2507,I371435,I371690,);
not I_21715 (I371698,I371690);
not I_21716 (I371715,I371673);
nand I_21717 (I371412,I371715,I371534);
nand I_21718 (I371746,I1198249,I1198255);
and I_21719 (I371763,I371746,I1198267);
DFFARX1 I_21720 (I371763,I2507,I371435,I371789,);
nor I_21721 (I371797,I371789,I371461);
DFFARX1 I_21722 (I371797,I2507,I371435,I371400,);
DFFARX1 I_21723 (I371789,I2507,I371435,I371418,);
nor I_21724 (I371842,I1198258,I1198255);
not I_21725 (I371859,I371842);
nor I_21726 (I371421,I371698,I371859);
nand I_21727 (I371406,I371715,I371859);
nor I_21728 (I371415,I371461,I371842);
DFFARX1 I_21729 (I371842,I2507,I371435,I371424,);
not I_21730 (I371962,I2514);
DFFARX1 I_21731 (I1298614,I2507,I371962,I371988,);
nand I_21732 (I371996,I1298641,I1298617);
and I_21733 (I372013,I371996,I1298626);
DFFARX1 I_21734 (I372013,I2507,I371962,I372039,);
nor I_21735 (I371930,I372039,I371988);
not I_21736 (I372061,I372039);
DFFARX1 I_21737 (I1298614,I2507,I371962,I372087,);
nand I_21738 (I372095,I372087,I1298638);
not I_21739 (I372112,I372095);
DFFARX1 I_21740 (I372112,I2507,I371962,I372138,);
not I_21741 (I371954,I372138);
nor I_21742 (I372160,I371988,I372095);
nor I_21743 (I371936,I372039,I372160);
DFFARX1 I_21744 (I1298620,I2507,I371962,I372200,);
DFFARX1 I_21745 (I372200,I2507,I371962,I372217,);
not I_21746 (I372225,I372217);
not I_21747 (I372242,I372200);
nand I_21748 (I371939,I372242,I372061);
nand I_21749 (I372273,I1298635,I1298623);
and I_21750 (I372290,I372273,I1298629);
DFFARX1 I_21751 (I372290,I2507,I371962,I372316,);
nor I_21752 (I372324,I372316,I371988);
DFFARX1 I_21753 (I372324,I2507,I371962,I371927,);
DFFARX1 I_21754 (I372316,I2507,I371962,I371945,);
nor I_21755 (I372369,I1298632,I1298623);
not I_21756 (I372386,I372369);
nor I_21757 (I371948,I372225,I372386);
nand I_21758 (I371933,I372242,I372386);
nor I_21759 (I371942,I371988,I372369);
DFFARX1 I_21760 (I372369,I2507,I371962,I371951,);
not I_21761 (I372489,I2514);
DFFARX1 I_21762 (I870234,I2507,I372489,I372515,);
nand I_21763 (I372523,I870237,I870231);
and I_21764 (I372540,I372523,I870243);
DFFARX1 I_21765 (I372540,I2507,I372489,I372566,);
nor I_21766 (I372457,I372566,I372515);
not I_21767 (I372588,I372566);
DFFARX1 I_21768 (I870246,I2507,I372489,I372614,);
nand I_21769 (I372622,I372614,I870237);
not I_21770 (I372639,I372622);
DFFARX1 I_21771 (I372639,I2507,I372489,I372665,);
not I_21772 (I372481,I372665);
nor I_21773 (I372687,I372515,I372622);
nor I_21774 (I372463,I372566,I372687);
DFFARX1 I_21775 (I870249,I2507,I372489,I372727,);
DFFARX1 I_21776 (I372727,I2507,I372489,I372744,);
not I_21777 (I372752,I372744);
not I_21778 (I372769,I372727);
nand I_21779 (I372466,I372769,I372588);
nand I_21780 (I372800,I870231,I870240);
and I_21781 (I372817,I372800,I870234);
DFFARX1 I_21782 (I372817,I2507,I372489,I372843,);
nor I_21783 (I372851,I372843,I372515);
DFFARX1 I_21784 (I372851,I2507,I372489,I372454,);
DFFARX1 I_21785 (I372843,I2507,I372489,I372472,);
nor I_21786 (I372896,I870252,I870240);
not I_21787 (I372913,I372896);
nor I_21788 (I372475,I372752,I372913);
nand I_21789 (I372460,I372769,I372913);
nor I_21790 (I372469,I372515,I372896);
DFFARX1 I_21791 (I372896,I2507,I372489,I372478,);
not I_21792 (I373016,I2514);
DFFARX1 I_21793 (I728412,I2507,I373016,I373042,);
nand I_21794 (I373050,I728403,I728418);
and I_21795 (I373067,I373050,I728424);
DFFARX1 I_21796 (I373067,I2507,I373016,I373093,);
nor I_21797 (I372984,I373093,I373042);
not I_21798 (I373115,I373093);
DFFARX1 I_21799 (I728409,I2507,I373016,I373141,);
nand I_21800 (I373149,I373141,I728403);
not I_21801 (I373166,I373149);
DFFARX1 I_21802 (I373166,I2507,I373016,I373192,);
not I_21803 (I373008,I373192);
nor I_21804 (I373214,I373042,I373149);
nor I_21805 (I372990,I373093,I373214);
DFFARX1 I_21806 (I728406,I2507,I373016,I373254,);
DFFARX1 I_21807 (I373254,I2507,I373016,I373271,);
not I_21808 (I373279,I373271);
not I_21809 (I373296,I373254);
nand I_21810 (I372993,I373296,I373115);
nand I_21811 (I373327,I728400,I728415);
and I_21812 (I373344,I373327,I728400);
DFFARX1 I_21813 (I373344,I2507,I373016,I373370,);
nor I_21814 (I373378,I373370,I373042);
DFFARX1 I_21815 (I373378,I2507,I373016,I372981,);
DFFARX1 I_21816 (I373370,I2507,I373016,I372999,);
nor I_21817 (I373423,I728421,I728415);
not I_21818 (I373440,I373423);
nor I_21819 (I373002,I373279,I373440);
nand I_21820 (I372987,I373296,I373440);
nor I_21821 (I372996,I373042,I373423);
DFFARX1 I_21822 (I373423,I2507,I373016,I373005,);
not I_21823 (I373543,I2514);
DFFARX1 I_21824 (I1037072,I2507,I373543,I373569,);
nand I_21825 (I373577,I1037069,I1037072);
and I_21826 (I373594,I373577,I1037081);
DFFARX1 I_21827 (I373594,I2507,I373543,I373620,);
nor I_21828 (I373511,I373620,I373569);
not I_21829 (I373642,I373620);
DFFARX1 I_21830 (I1037069,I2507,I373543,I373668,);
nand I_21831 (I373676,I373668,I1037087);
not I_21832 (I373693,I373676);
DFFARX1 I_21833 (I373693,I2507,I373543,I373719,);
not I_21834 (I373535,I373719);
nor I_21835 (I373741,I373569,I373676);
nor I_21836 (I373517,I373620,I373741);
DFFARX1 I_21837 (I1037075,I2507,I373543,I373781,);
DFFARX1 I_21838 (I373781,I2507,I373543,I373798,);
not I_21839 (I373806,I373798);
not I_21840 (I373823,I373781);
nand I_21841 (I373520,I373823,I373642);
nand I_21842 (I373854,I1037084,I1037090);
and I_21843 (I373871,I373854,I1037075);
DFFARX1 I_21844 (I373871,I2507,I373543,I373897,);
nor I_21845 (I373905,I373897,I373569);
DFFARX1 I_21846 (I373905,I2507,I373543,I373508,);
DFFARX1 I_21847 (I373897,I2507,I373543,I373526,);
nor I_21848 (I373950,I1037078,I1037090);
not I_21849 (I373967,I373950);
nor I_21850 (I373529,I373806,I373967);
nand I_21851 (I373514,I373823,I373967);
nor I_21852 (I373523,I373569,I373950);
DFFARX1 I_21853 (I373950,I2507,I373543,I373532,);
not I_21854 (I374070,I2514);
DFFARX1 I_21855 (I983828,I2507,I374070,I374096,);
nand I_21856 (I374104,I983825,I983843);
and I_21857 (I374121,I374104,I983834);
DFFARX1 I_21858 (I374121,I2507,I374070,I374147,);
nor I_21859 (I374038,I374147,I374096);
not I_21860 (I374169,I374147);
DFFARX1 I_21861 (I983849,I2507,I374070,I374195,);
nand I_21862 (I374203,I374195,I983831);
not I_21863 (I374220,I374203);
DFFARX1 I_21864 (I374220,I2507,I374070,I374246,);
not I_21865 (I374062,I374246);
nor I_21866 (I374268,I374096,I374203);
nor I_21867 (I374044,I374147,I374268);
DFFARX1 I_21868 (I983837,I2507,I374070,I374308,);
DFFARX1 I_21869 (I374308,I2507,I374070,I374325,);
not I_21870 (I374333,I374325);
not I_21871 (I374350,I374308);
nand I_21872 (I374047,I374350,I374169);
nand I_21873 (I374381,I983825,I983852);
and I_21874 (I374398,I374381,I983840);
DFFARX1 I_21875 (I374398,I2507,I374070,I374424,);
nor I_21876 (I374432,I374424,I374096);
DFFARX1 I_21877 (I374432,I2507,I374070,I374035,);
DFFARX1 I_21878 (I374424,I2507,I374070,I374053,);
nor I_21879 (I374477,I983846,I983852);
not I_21880 (I374494,I374477);
nor I_21881 (I374056,I374333,I374494);
nand I_21882 (I374041,I374350,I374494);
nor I_21883 (I374050,I374096,I374477);
DFFARX1 I_21884 (I374477,I2507,I374070,I374059,);
not I_21885 (I374597,I2514);
DFFARX1 I_21886 (I139544,I2507,I374597,I374623,);
nand I_21887 (I374631,I139529,I139520);
and I_21888 (I374648,I374631,I139535);
DFFARX1 I_21889 (I374648,I2507,I374597,I374674,);
nor I_21890 (I374565,I374674,I374623);
not I_21891 (I374696,I374674);
DFFARX1 I_21892 (I139547,I2507,I374597,I374722,);
nand I_21893 (I374730,I374722,I139538);
not I_21894 (I374747,I374730);
DFFARX1 I_21895 (I374747,I2507,I374597,I374773,);
not I_21896 (I374589,I374773);
nor I_21897 (I374795,I374623,I374730);
nor I_21898 (I374571,I374674,I374795);
DFFARX1 I_21899 (I139526,I2507,I374597,I374835,);
DFFARX1 I_21900 (I374835,I2507,I374597,I374852,);
not I_21901 (I374860,I374852);
not I_21902 (I374877,I374835);
nand I_21903 (I374574,I374877,I374696);
nand I_21904 (I374908,I139532,I139523);
and I_21905 (I374925,I374908,I139520);
DFFARX1 I_21906 (I374925,I2507,I374597,I374951,);
nor I_21907 (I374959,I374951,I374623);
DFFARX1 I_21908 (I374959,I2507,I374597,I374562,);
DFFARX1 I_21909 (I374951,I2507,I374597,I374580,);
nor I_21910 (I375004,I139541,I139523);
not I_21911 (I375021,I375004);
nor I_21912 (I374583,I374860,I375021);
nand I_21913 (I374568,I374877,I375021);
nor I_21914 (I374577,I374623,I375004);
DFFARX1 I_21915 (I375004,I2507,I374597,I374586,);
not I_21916 (I375124,I2514);
DFFARX1 I_21917 (I1308308,I2507,I375124,I375150,);
nand I_21918 (I375158,I1308287,I1308287);
and I_21919 (I375175,I375158,I1308314);
DFFARX1 I_21920 (I375175,I2507,I375124,I375201,);
nor I_21921 (I375092,I375201,I375150);
not I_21922 (I375223,I375201);
DFFARX1 I_21923 (I1308302,I2507,I375124,I375249,);
nand I_21924 (I375257,I375249,I1308305);
not I_21925 (I375274,I375257);
DFFARX1 I_21926 (I375274,I2507,I375124,I375300,);
not I_21927 (I375116,I375300);
nor I_21928 (I375322,I375150,I375257);
nor I_21929 (I375098,I375201,I375322);
DFFARX1 I_21930 (I1308296,I2507,I375124,I375362,);
DFFARX1 I_21931 (I375362,I2507,I375124,I375379,);
not I_21932 (I375387,I375379);
not I_21933 (I375404,I375362);
nand I_21934 (I375101,I375404,I375223);
nand I_21935 (I375435,I1308293,I1308290);
and I_21936 (I375452,I375435,I1308311);
DFFARX1 I_21937 (I375452,I2507,I375124,I375478,);
nor I_21938 (I375486,I375478,I375150);
DFFARX1 I_21939 (I375486,I2507,I375124,I375089,);
DFFARX1 I_21940 (I375478,I2507,I375124,I375107,);
nor I_21941 (I375531,I1308299,I1308290);
not I_21942 (I375548,I375531);
nor I_21943 (I375110,I375387,I375548);
nand I_21944 (I375095,I375404,I375548);
nor I_21945 (I375104,I375150,I375531);
DFFARX1 I_21946 (I375531,I2507,I375124,I375113,);
not I_21947 (I375651,I2514);
DFFARX1 I_21948 (I1124262,I2507,I375651,I375677,);
nand I_21949 (I375685,I1124277,I1124262);
and I_21950 (I375702,I375685,I1124280);
DFFARX1 I_21951 (I375702,I2507,I375651,I375728,);
nor I_21952 (I375619,I375728,I375677);
not I_21953 (I375750,I375728);
DFFARX1 I_21954 (I1124286,I2507,I375651,I375776,);
nand I_21955 (I375784,I375776,I1124268);
not I_21956 (I375801,I375784);
DFFARX1 I_21957 (I375801,I2507,I375651,I375827,);
not I_21958 (I375643,I375827);
nor I_21959 (I375849,I375677,I375784);
nor I_21960 (I375625,I375728,I375849);
DFFARX1 I_21961 (I1124265,I2507,I375651,I375889,);
DFFARX1 I_21962 (I375889,I2507,I375651,I375906,);
not I_21963 (I375914,I375906);
not I_21964 (I375931,I375889);
nand I_21965 (I375628,I375931,I375750);
nand I_21966 (I375962,I1124265,I1124271);
and I_21967 (I375979,I375962,I1124283);
DFFARX1 I_21968 (I375979,I2507,I375651,I376005,);
nor I_21969 (I376013,I376005,I375677);
DFFARX1 I_21970 (I376013,I2507,I375651,I375616,);
DFFARX1 I_21971 (I376005,I2507,I375651,I375634,);
nor I_21972 (I376058,I1124274,I1124271);
not I_21973 (I376075,I376058);
nor I_21974 (I375637,I375914,I376075);
nand I_21975 (I375622,I375931,I376075);
nor I_21976 (I375631,I375677,I376058);
DFFARX1 I_21977 (I376058,I2507,I375651,I375640,);
not I_21978 (I376178,I2514);
DFFARX1 I_21979 (I182369,I2507,I376178,I376204,);
DFFARX1 I_21980 (I376204,I2507,I376178,I376221,);
not I_21981 (I376170,I376221);
not I_21982 (I376243,I376204);
nand I_21983 (I376260,I182381,I182360);
and I_21984 (I376277,I376260,I182363);
DFFARX1 I_21985 (I376277,I2507,I376178,I376303,);
not I_21986 (I376311,I376303);
DFFARX1 I_21987 (I182372,I2507,I376178,I376337,);
and I_21988 (I376345,I376337,I182384);
nand I_21989 (I376362,I376337,I182384);
nand I_21990 (I376149,I376311,I376362);
DFFARX1 I_21991 (I182378,I2507,I376178,I376402,);
nor I_21992 (I376410,I376402,I376345);
DFFARX1 I_21993 (I376410,I2507,I376178,I376143,);
nor I_21994 (I376158,I376402,I376303);
nand I_21995 (I376455,I182366,I182363);
and I_21996 (I376472,I376455,I182375);
DFFARX1 I_21997 (I376472,I2507,I376178,I376498,);
nor I_21998 (I376146,I376498,I376402);
not I_21999 (I376520,I376498);
nor I_22000 (I376537,I376520,I376311);
nor I_22001 (I376554,I376243,I376537);
DFFARX1 I_22002 (I376554,I2507,I376178,I376161,);
nor I_22003 (I376585,I376520,I376402);
nor I_22004 (I376602,I182360,I182363);
nor I_22005 (I376152,I376602,I376585);
not I_22006 (I376633,I376602);
nand I_22007 (I376155,I376362,I376633);
DFFARX1 I_22008 (I376602,I2507,I376178,I376167,);
DFFARX1 I_22009 (I376602,I2507,I376178,I376164,);
not I_22010 (I376722,I2514);
DFFARX1 I_22011 (I961221,I2507,I376722,I376748,);
DFFARX1 I_22012 (I376748,I2507,I376722,I376765,);
not I_22013 (I376714,I376765);
not I_22014 (I376787,I376748);
nand I_22015 (I376804,I961236,I961224);
and I_22016 (I376821,I376804,I961215);
DFFARX1 I_22017 (I376821,I2507,I376722,I376847,);
not I_22018 (I376855,I376847);
DFFARX1 I_22019 (I961227,I2507,I376722,I376881,);
and I_22020 (I376889,I376881,I961218);
nand I_22021 (I376906,I376881,I961218);
nand I_22022 (I376693,I376855,I376906);
DFFARX1 I_22023 (I961233,I2507,I376722,I376946,);
nor I_22024 (I376954,I376946,I376889);
DFFARX1 I_22025 (I376954,I2507,I376722,I376687,);
nor I_22026 (I376702,I376946,I376847);
nand I_22027 (I376999,I961242,I961230);
and I_22028 (I377016,I376999,I961239);
DFFARX1 I_22029 (I377016,I2507,I376722,I377042,);
nor I_22030 (I376690,I377042,I376946);
not I_22031 (I377064,I377042);
nor I_22032 (I377081,I377064,I376855);
nor I_22033 (I377098,I376787,I377081);
DFFARX1 I_22034 (I377098,I2507,I376722,I376705,);
nor I_22035 (I377129,I377064,I376946);
nor I_22036 (I377146,I961215,I961230);
nor I_22037 (I376696,I377146,I377129);
not I_22038 (I377177,I377146);
nand I_22039 (I376699,I376906,I377177);
DFFARX1 I_22040 (I377146,I2507,I376722,I376711,);
DFFARX1 I_22041 (I377146,I2507,I376722,I376708,);
not I_22042 (I377266,I2514);
DFFARX1 I_22043 (I1238437,I2507,I377266,I377292,);
DFFARX1 I_22044 (I377292,I2507,I377266,I377309,);
not I_22045 (I377258,I377309);
not I_22046 (I377331,I377292);
nand I_22047 (I377348,I1238449,I1238452);
and I_22048 (I377365,I377348,I1238455);
DFFARX1 I_22049 (I377365,I2507,I377266,I377391,);
not I_22050 (I377399,I377391);
DFFARX1 I_22051 (I1238440,I2507,I377266,I377425,);
and I_22052 (I377433,I377425,I1238446);
nand I_22053 (I377450,I377425,I1238446);
nand I_22054 (I377237,I377399,I377450);
DFFARX1 I_22055 (I1238434,I2507,I377266,I377490,);
nor I_22056 (I377498,I377490,I377433);
DFFARX1 I_22057 (I377498,I2507,I377266,I377231,);
nor I_22058 (I377246,I377490,I377391);
nand I_22059 (I377543,I1238437,I1238458);
and I_22060 (I377560,I377543,I1238443);
DFFARX1 I_22061 (I377560,I2507,I377266,I377586,);
nor I_22062 (I377234,I377586,I377490);
not I_22063 (I377608,I377586);
nor I_22064 (I377625,I377608,I377399);
nor I_22065 (I377642,I377331,I377625);
DFFARX1 I_22066 (I377642,I2507,I377266,I377249,);
nor I_22067 (I377673,I377608,I377490);
nor I_22068 (I377690,I1238434,I1238458);
nor I_22069 (I377240,I377690,I377673);
not I_22070 (I377721,I377690);
nand I_22071 (I377243,I377450,I377721);
DFFARX1 I_22072 (I377690,I2507,I377266,I377255,);
DFFARX1 I_22073 (I377690,I2507,I377266,I377252,);
not I_22074 (I377810,I2514);
DFFARX1 I_22075 (I578123,I2507,I377810,I377836,);
DFFARX1 I_22076 (I377836,I2507,I377810,I377853,);
not I_22077 (I377802,I377853);
not I_22078 (I377875,I377836);
nand I_22079 (I377892,I578120,I578141);
and I_22080 (I377909,I377892,I578144);
DFFARX1 I_22081 (I377909,I2507,I377810,I377935,);
not I_22082 (I377943,I377935);
DFFARX1 I_22083 (I578129,I2507,I377810,I377969,);
and I_22084 (I377977,I377969,I578132);
nand I_22085 (I377994,I377969,I578132);
nand I_22086 (I377781,I377943,I377994);
DFFARX1 I_22087 (I578135,I2507,I377810,I378034,);
nor I_22088 (I378042,I378034,I377977);
DFFARX1 I_22089 (I378042,I2507,I377810,I377775,);
nor I_22090 (I377790,I378034,I377935);
nand I_22091 (I378087,I578120,I578126);
and I_22092 (I378104,I378087,I578138);
DFFARX1 I_22093 (I378104,I2507,I377810,I378130,);
nor I_22094 (I377778,I378130,I378034);
not I_22095 (I378152,I378130);
nor I_22096 (I378169,I378152,I377943);
nor I_22097 (I378186,I377875,I378169);
DFFARX1 I_22098 (I378186,I2507,I377810,I377793,);
nor I_22099 (I378217,I378152,I378034);
nor I_22100 (I378234,I578123,I578126);
nor I_22101 (I377784,I378234,I378217);
not I_22102 (I378265,I378234);
nand I_22103 (I377787,I377994,I378265);
DFFARX1 I_22104 (I378234,I2507,I377810,I377799,);
DFFARX1 I_22105 (I378234,I2507,I377810,I377796,);
not I_22106 (I378354,I2514);
DFFARX1 I_22107 (I1213957,I2507,I378354,I378380,);
DFFARX1 I_22108 (I378380,I2507,I378354,I378397,);
not I_22109 (I378346,I378397);
not I_22110 (I378419,I378380);
nand I_22111 (I378436,I1213969,I1213972);
and I_22112 (I378453,I378436,I1213975);
DFFARX1 I_22113 (I378453,I2507,I378354,I378479,);
not I_22114 (I378487,I378479);
DFFARX1 I_22115 (I1213960,I2507,I378354,I378513,);
and I_22116 (I378521,I378513,I1213966);
nand I_22117 (I378538,I378513,I1213966);
nand I_22118 (I378325,I378487,I378538);
DFFARX1 I_22119 (I1213954,I2507,I378354,I378578,);
nor I_22120 (I378586,I378578,I378521);
DFFARX1 I_22121 (I378586,I2507,I378354,I378319,);
nor I_22122 (I378334,I378578,I378479);
nand I_22123 (I378631,I1213957,I1213978);
and I_22124 (I378648,I378631,I1213963);
DFFARX1 I_22125 (I378648,I2507,I378354,I378674,);
nor I_22126 (I378322,I378674,I378578);
not I_22127 (I378696,I378674);
nor I_22128 (I378713,I378696,I378487);
nor I_22129 (I378730,I378419,I378713);
DFFARX1 I_22130 (I378730,I2507,I378354,I378337,);
nor I_22131 (I378761,I378696,I378578);
nor I_22132 (I378778,I1213954,I1213978);
nor I_22133 (I378328,I378778,I378761);
not I_22134 (I378809,I378778);
nand I_22135 (I378331,I378538,I378809);
DFFARX1 I_22136 (I378778,I2507,I378354,I378343,);
DFFARX1 I_22137 (I378778,I2507,I378354,I378340,);
not I_22138 (I378898,I2514);
DFFARX1 I_22139 (I863392,I2507,I378898,I378924,);
DFFARX1 I_22140 (I378924,I2507,I378898,I378941,);
not I_22141 (I378890,I378941);
not I_22142 (I378963,I378924);
nand I_22143 (I378980,I863386,I863383);
and I_22144 (I378997,I378980,I863398);
DFFARX1 I_22145 (I378997,I2507,I378898,I379023,);
not I_22146 (I379031,I379023);
DFFARX1 I_22147 (I863386,I2507,I378898,I379057,);
and I_22148 (I379065,I379057,I863380);
nand I_22149 (I379082,I379057,I863380);
nand I_22150 (I378869,I379031,I379082);
DFFARX1 I_22151 (I863380,I2507,I378898,I379122,);
nor I_22152 (I379130,I379122,I379065);
DFFARX1 I_22153 (I379130,I2507,I378898,I378863,);
nor I_22154 (I378878,I379122,I379023);
nand I_22155 (I379175,I863395,I863389);
and I_22156 (I379192,I379175,I863383);
DFFARX1 I_22157 (I379192,I2507,I378898,I379218,);
nor I_22158 (I378866,I379218,I379122);
not I_22159 (I379240,I379218);
nor I_22160 (I379257,I379240,I379031);
nor I_22161 (I379274,I378963,I379257);
DFFARX1 I_22162 (I379274,I2507,I378898,I378881,);
nor I_22163 (I379305,I379240,I379122);
nor I_22164 (I379322,I863401,I863389);
nor I_22165 (I378872,I379322,I379305);
not I_22166 (I379353,I379322);
nand I_22167 (I378875,I379082,I379353);
DFFARX1 I_22168 (I379322,I2507,I378898,I378887,);
DFFARX1 I_22169 (I379322,I2507,I378898,I378884,);
not I_22170 (I379442,I2514);
DFFARX1 I_22171 (I1207973,I2507,I379442,I379468,);
DFFARX1 I_22172 (I379468,I2507,I379442,I379485,);
not I_22173 (I379434,I379485);
not I_22174 (I379507,I379468);
nand I_22175 (I379524,I1207985,I1207988);
and I_22176 (I379541,I379524,I1207991);
DFFARX1 I_22177 (I379541,I2507,I379442,I379567,);
not I_22178 (I379575,I379567);
DFFARX1 I_22179 (I1207976,I2507,I379442,I379601,);
and I_22180 (I379609,I379601,I1207982);
nand I_22181 (I379626,I379601,I1207982);
nand I_22182 (I379413,I379575,I379626);
DFFARX1 I_22183 (I1207970,I2507,I379442,I379666,);
nor I_22184 (I379674,I379666,I379609);
DFFARX1 I_22185 (I379674,I2507,I379442,I379407,);
nor I_22186 (I379422,I379666,I379567);
nand I_22187 (I379719,I1207973,I1207994);
and I_22188 (I379736,I379719,I1207979);
DFFARX1 I_22189 (I379736,I2507,I379442,I379762,);
nor I_22190 (I379410,I379762,I379666);
not I_22191 (I379784,I379762);
nor I_22192 (I379801,I379784,I379575);
nor I_22193 (I379818,I379507,I379801);
DFFARX1 I_22194 (I379818,I2507,I379442,I379425,);
nor I_22195 (I379849,I379784,I379666);
nor I_22196 (I379866,I1207970,I1207994);
nor I_22197 (I379416,I379866,I379849);
not I_22198 (I379897,I379866);
nand I_22199 (I379419,I379626,I379897);
DFFARX1 I_22200 (I379866,I2507,I379442,I379431,);
DFFARX1 I_22201 (I379866,I2507,I379442,I379428,);
not I_22202 (I379986,I2514);
DFFARX1 I_22203 (I175229,I2507,I379986,I380012,);
DFFARX1 I_22204 (I380012,I2507,I379986,I380029,);
not I_22205 (I379978,I380029);
not I_22206 (I380051,I380012);
nand I_22207 (I380068,I175241,I175220);
and I_22208 (I380085,I380068,I175223);
DFFARX1 I_22209 (I380085,I2507,I379986,I380111,);
not I_22210 (I380119,I380111);
DFFARX1 I_22211 (I175232,I2507,I379986,I380145,);
and I_22212 (I380153,I380145,I175244);
nand I_22213 (I380170,I380145,I175244);
nand I_22214 (I379957,I380119,I380170);
DFFARX1 I_22215 (I175238,I2507,I379986,I380210,);
nor I_22216 (I380218,I380210,I380153);
DFFARX1 I_22217 (I380218,I2507,I379986,I379951,);
nor I_22218 (I379966,I380210,I380111);
nand I_22219 (I380263,I175226,I175223);
and I_22220 (I380280,I380263,I175235);
DFFARX1 I_22221 (I380280,I2507,I379986,I380306,);
nor I_22222 (I379954,I380306,I380210);
not I_22223 (I380328,I380306);
nor I_22224 (I380345,I380328,I380119);
nor I_22225 (I380362,I380051,I380345);
DFFARX1 I_22226 (I380362,I2507,I379986,I379969,);
nor I_22227 (I380393,I380328,I380210);
nor I_22228 (I380410,I175220,I175223);
nor I_22229 (I379960,I380410,I380393);
not I_22230 (I380441,I380410);
nand I_22231 (I379963,I380170,I380441);
DFFARX1 I_22232 (I380410,I2507,I379986,I379975,);
DFFARX1 I_22233 (I380410,I2507,I379986,I379972,);
not I_22234 (I380530,I2514);
DFFARX1 I_22235 (I1249861,I2507,I380530,I380556,);
DFFARX1 I_22236 (I380556,I2507,I380530,I380573,);
not I_22237 (I380522,I380573);
not I_22238 (I380595,I380556);
nand I_22239 (I380612,I1249873,I1249876);
and I_22240 (I380629,I380612,I1249879);
DFFARX1 I_22241 (I380629,I2507,I380530,I380655,);
not I_22242 (I380663,I380655);
DFFARX1 I_22243 (I1249864,I2507,I380530,I380689,);
and I_22244 (I380697,I380689,I1249870);
nand I_22245 (I380714,I380689,I1249870);
nand I_22246 (I380501,I380663,I380714);
DFFARX1 I_22247 (I1249858,I2507,I380530,I380754,);
nor I_22248 (I380762,I380754,I380697);
DFFARX1 I_22249 (I380762,I2507,I380530,I380495,);
nor I_22250 (I380510,I380754,I380655);
nand I_22251 (I380807,I1249861,I1249882);
and I_22252 (I380824,I380807,I1249867);
DFFARX1 I_22253 (I380824,I2507,I380530,I380850,);
nor I_22254 (I380498,I380850,I380754);
not I_22255 (I380872,I380850);
nor I_22256 (I380889,I380872,I380663);
nor I_22257 (I380906,I380595,I380889);
DFFARX1 I_22258 (I380906,I2507,I380530,I380513,);
nor I_22259 (I380937,I380872,I380754);
nor I_22260 (I380954,I1249858,I1249882);
nor I_22261 (I380504,I380954,I380937);
not I_22262 (I380985,I380954);
nand I_22263 (I380507,I380714,I380985);
DFFARX1 I_22264 (I380954,I2507,I380530,I380519,);
DFFARX1 I_22265 (I380954,I2507,I380530,I380516,);
not I_22266 (I381074,I2514);
DFFARX1 I_22267 (I1258240,I2507,I381074,I381100,);
DFFARX1 I_22268 (I381100,I2507,I381074,I381117,);
not I_22269 (I381066,I381117);
not I_22270 (I381139,I381100);
nand I_22271 (I381156,I1258237,I1258234);
and I_22272 (I381173,I381156,I1258222);
DFFARX1 I_22273 (I381173,I2507,I381074,I381199,);
not I_22274 (I381207,I381199);
DFFARX1 I_22275 (I1258246,I2507,I381074,I381233,);
and I_22276 (I381241,I381233,I1258231);
nand I_22277 (I381258,I381233,I1258231);
nand I_22278 (I381045,I381207,I381258);
DFFARX1 I_22279 (I1258225,I2507,I381074,I381298,);
nor I_22280 (I381306,I381298,I381241);
DFFARX1 I_22281 (I381306,I2507,I381074,I381039,);
nor I_22282 (I381054,I381298,I381199);
nand I_22283 (I381351,I1258222,I1258228);
and I_22284 (I381368,I381351,I1258243);
DFFARX1 I_22285 (I381368,I2507,I381074,I381394,);
nor I_22286 (I381042,I381394,I381298);
not I_22287 (I381416,I381394);
nor I_22288 (I381433,I381416,I381207);
nor I_22289 (I381450,I381139,I381433);
DFFARX1 I_22290 (I381450,I2507,I381074,I381057,);
nor I_22291 (I381481,I381416,I381298);
nor I_22292 (I381498,I1258225,I1258228);
nor I_22293 (I381048,I381498,I381481);
not I_22294 (I381529,I381498);
nand I_22295 (I381051,I381258,I381529);
DFFARX1 I_22296 (I381498,I2507,I381074,I381063,);
DFFARX1 I_22297 (I381498,I2507,I381074,I381060,);
not I_22298 (I381618,I2514);
DFFARX1 I_22299 (I59082,I2507,I381618,I381644,);
DFFARX1 I_22300 (I381644,I2507,I381618,I381661,);
not I_22301 (I381610,I381661);
not I_22302 (I381683,I381644);
nand I_22303 (I381700,I59097,I59076);
and I_22304 (I381717,I381700,I59079);
DFFARX1 I_22305 (I381717,I2507,I381618,I381743,);
not I_22306 (I381751,I381743);
DFFARX1 I_22307 (I59085,I2507,I381618,I381777,);
and I_22308 (I381785,I381777,I59079);
nand I_22309 (I381802,I381777,I59079);
nand I_22310 (I381589,I381751,I381802);
DFFARX1 I_22311 (I59094,I2507,I381618,I381842,);
nor I_22312 (I381850,I381842,I381785);
DFFARX1 I_22313 (I381850,I2507,I381618,I381583,);
nor I_22314 (I381598,I381842,I381743);
nand I_22315 (I381895,I59076,I59091);
and I_22316 (I381912,I381895,I59088);
DFFARX1 I_22317 (I381912,I2507,I381618,I381938,);
nor I_22318 (I381586,I381938,I381842);
not I_22319 (I381960,I381938);
nor I_22320 (I381977,I381960,I381751);
nor I_22321 (I381994,I381683,I381977);
DFFARX1 I_22322 (I381994,I2507,I381618,I381601,);
nor I_22323 (I382025,I381960,I381842);
nor I_22324 (I382042,I59100,I59091);
nor I_22325 (I381592,I382042,I382025);
not I_22326 (I382073,I382042);
nand I_22327 (I381595,I381802,I382073);
DFFARX1 I_22328 (I382042,I2507,I381618,I381607,);
DFFARX1 I_22329 (I382042,I2507,I381618,I381604,);
not I_22330 (I382162,I2514);
DFFARX1 I_22331 (I545755,I2507,I382162,I382188,);
DFFARX1 I_22332 (I382188,I2507,I382162,I382205,);
not I_22333 (I382154,I382205);
not I_22334 (I382227,I382188);
nand I_22335 (I382244,I545752,I545773);
and I_22336 (I382261,I382244,I545776);
DFFARX1 I_22337 (I382261,I2507,I382162,I382287,);
not I_22338 (I382295,I382287);
DFFARX1 I_22339 (I545761,I2507,I382162,I382321,);
and I_22340 (I382329,I382321,I545764);
nand I_22341 (I382346,I382321,I545764);
nand I_22342 (I382133,I382295,I382346);
DFFARX1 I_22343 (I545767,I2507,I382162,I382386,);
nor I_22344 (I382394,I382386,I382329);
DFFARX1 I_22345 (I382394,I2507,I382162,I382127,);
nor I_22346 (I382142,I382386,I382287);
nand I_22347 (I382439,I545752,I545758);
and I_22348 (I382456,I382439,I545770);
DFFARX1 I_22349 (I382456,I2507,I382162,I382482,);
nor I_22350 (I382130,I382482,I382386);
not I_22351 (I382504,I382482);
nor I_22352 (I382521,I382504,I382295);
nor I_22353 (I382538,I382227,I382521);
DFFARX1 I_22354 (I382538,I2507,I382162,I382145,);
nor I_22355 (I382569,I382504,I382386);
nor I_22356 (I382586,I545755,I545758);
nor I_22357 (I382136,I382586,I382569);
not I_22358 (I382617,I382586);
nand I_22359 (I382139,I382346,I382617);
DFFARX1 I_22360 (I382586,I2507,I382162,I382151,);
DFFARX1 I_22361 (I382586,I2507,I382162,I382148,);
not I_22362 (I382706,I2514);
DFFARX1 I_22363 (I176419,I2507,I382706,I382732,);
DFFARX1 I_22364 (I382732,I2507,I382706,I382749,);
not I_22365 (I382698,I382749);
not I_22366 (I382771,I382732);
nand I_22367 (I382788,I176431,I176410);
and I_22368 (I382805,I382788,I176413);
DFFARX1 I_22369 (I382805,I2507,I382706,I382831,);
not I_22370 (I382839,I382831);
DFFARX1 I_22371 (I176422,I2507,I382706,I382865,);
and I_22372 (I382873,I382865,I176434);
nand I_22373 (I382890,I382865,I176434);
nand I_22374 (I382677,I382839,I382890);
DFFARX1 I_22375 (I176428,I2507,I382706,I382930,);
nor I_22376 (I382938,I382930,I382873);
DFFARX1 I_22377 (I382938,I2507,I382706,I382671,);
nor I_22378 (I382686,I382930,I382831);
nand I_22379 (I382983,I176416,I176413);
and I_22380 (I383000,I382983,I176425);
DFFARX1 I_22381 (I383000,I2507,I382706,I383026,);
nor I_22382 (I382674,I383026,I382930);
not I_22383 (I383048,I383026);
nor I_22384 (I383065,I383048,I382839);
nor I_22385 (I383082,I382771,I383065);
DFFARX1 I_22386 (I383082,I2507,I382706,I382689,);
nor I_22387 (I383113,I383048,I382930);
nor I_22388 (I383130,I176410,I176413);
nor I_22389 (I382680,I383130,I383113);
not I_22390 (I383161,I383130);
nand I_22391 (I382683,I382890,I383161);
DFFARX1 I_22392 (I383130,I2507,I382706,I382695,);
DFFARX1 I_22393 (I383130,I2507,I382706,I382692,);
not I_22394 (I383250,I2514);
DFFARX1 I_22395 (I10865,I2507,I383250,I383276,);
DFFARX1 I_22396 (I383276,I2507,I383250,I383293,);
not I_22397 (I383242,I383293);
not I_22398 (I383315,I383276);
nand I_22399 (I383332,I10868,I10856);
and I_22400 (I383349,I383332,I10862);
DFFARX1 I_22401 (I383349,I2507,I383250,I383375,);
not I_22402 (I383383,I383375);
DFFARX1 I_22403 (I10850,I2507,I383250,I383409,);
and I_22404 (I383417,I383409,I10847);
nand I_22405 (I383434,I383409,I10847);
nand I_22406 (I383221,I383383,I383434);
DFFARX1 I_22407 (I10853,I2507,I383250,I383474,);
nor I_22408 (I383482,I383474,I383417);
DFFARX1 I_22409 (I383482,I2507,I383250,I383215,);
nor I_22410 (I383230,I383474,I383375);
nand I_22411 (I383527,I10853,I10850);
and I_22412 (I383544,I383527,I10847);
DFFARX1 I_22413 (I383544,I2507,I383250,I383570,);
nor I_22414 (I383218,I383570,I383474);
not I_22415 (I383592,I383570);
nor I_22416 (I383609,I383592,I383383);
nor I_22417 (I383626,I383315,I383609);
DFFARX1 I_22418 (I383626,I2507,I383250,I383233,);
nor I_22419 (I383657,I383592,I383474);
nor I_22420 (I383674,I10859,I10850);
nor I_22421 (I383224,I383674,I383657);
not I_22422 (I383705,I383674);
nand I_22423 (I383227,I383434,I383705);
DFFARX1 I_22424 (I383674,I2507,I383250,I383239,);
DFFARX1 I_22425 (I383674,I2507,I383250,I383236,);
not I_22426 (I383794,I2514);
DFFARX1 I_22427 (I1259974,I2507,I383794,I383820,);
DFFARX1 I_22428 (I383820,I2507,I383794,I383837,);
not I_22429 (I383786,I383837);
not I_22430 (I383859,I383820);
nand I_22431 (I383876,I1259971,I1259968);
and I_22432 (I383893,I383876,I1259956);
DFFARX1 I_22433 (I383893,I2507,I383794,I383919,);
not I_22434 (I383927,I383919);
DFFARX1 I_22435 (I1259980,I2507,I383794,I383953,);
and I_22436 (I383961,I383953,I1259965);
nand I_22437 (I383978,I383953,I1259965);
nand I_22438 (I383765,I383927,I383978);
DFFARX1 I_22439 (I1259959,I2507,I383794,I384018,);
nor I_22440 (I384026,I384018,I383961);
DFFARX1 I_22441 (I384026,I2507,I383794,I383759,);
nor I_22442 (I383774,I384018,I383919);
nand I_22443 (I384071,I1259956,I1259962);
and I_22444 (I384088,I384071,I1259977);
DFFARX1 I_22445 (I384088,I2507,I383794,I384114,);
nor I_22446 (I383762,I384114,I384018);
not I_22447 (I384136,I384114);
nor I_22448 (I384153,I384136,I383927);
nor I_22449 (I384170,I383859,I384153);
DFFARX1 I_22450 (I384170,I2507,I383794,I383777,);
nor I_22451 (I384201,I384136,I384018);
nor I_22452 (I384218,I1259959,I1259962);
nor I_22453 (I383768,I384218,I384201);
not I_22454 (I384249,I384218);
nand I_22455 (I383771,I383978,I384249);
DFFARX1 I_22456 (I384218,I2507,I383794,I383783,);
DFFARX1 I_22457 (I384218,I2507,I383794,I383780,);
not I_22458 (I384338,I2514);
DFFARX1 I_22459 (I1108081,I2507,I384338,I384364,);
DFFARX1 I_22460 (I384364,I2507,I384338,I384381,);
not I_22461 (I384330,I384381);
not I_22462 (I384403,I384364);
nand I_22463 (I384420,I1108093,I1108081);
and I_22464 (I384437,I384420,I1108084);
DFFARX1 I_22465 (I384437,I2507,I384338,I384463,);
not I_22466 (I384471,I384463);
DFFARX1 I_22467 (I1108102,I2507,I384338,I384497,);
and I_22468 (I384505,I384497,I1108078);
nand I_22469 (I384522,I384497,I1108078);
nand I_22470 (I384309,I384471,I384522);
DFFARX1 I_22471 (I1108096,I2507,I384338,I384562,);
nor I_22472 (I384570,I384562,I384505);
DFFARX1 I_22473 (I384570,I2507,I384338,I384303,);
nor I_22474 (I384318,I384562,I384463);
nand I_22475 (I384615,I1108090,I1108087);
and I_22476 (I384632,I384615,I1108099);
DFFARX1 I_22477 (I384632,I2507,I384338,I384658,);
nor I_22478 (I384306,I384658,I384562);
not I_22479 (I384680,I384658);
nor I_22480 (I384697,I384680,I384471);
nor I_22481 (I384714,I384403,I384697);
DFFARX1 I_22482 (I384714,I2507,I384338,I384321,);
nor I_22483 (I384745,I384680,I384562);
nor I_22484 (I384762,I1108078,I1108087);
nor I_22485 (I384312,I384762,I384745);
not I_22486 (I384793,I384762);
nand I_22487 (I384315,I384522,I384793);
DFFARX1 I_22488 (I384762,I2507,I384338,I384327,);
DFFARX1 I_22489 (I384762,I2507,I384338,I384324,);
not I_22490 (I384882,I2514);
DFFARX1 I_22491 (I111782,I2507,I384882,I384908,);
DFFARX1 I_22492 (I384908,I2507,I384882,I384925,);
not I_22493 (I384874,I384925);
not I_22494 (I384947,I384908);
nand I_22495 (I384964,I111797,I111776);
and I_22496 (I384981,I384964,I111779);
DFFARX1 I_22497 (I384981,I2507,I384882,I385007,);
not I_22498 (I385015,I385007);
DFFARX1 I_22499 (I111785,I2507,I384882,I385041,);
and I_22500 (I385049,I385041,I111779);
nand I_22501 (I385066,I385041,I111779);
nand I_22502 (I384853,I385015,I385066);
DFFARX1 I_22503 (I111794,I2507,I384882,I385106,);
nor I_22504 (I385114,I385106,I385049);
DFFARX1 I_22505 (I385114,I2507,I384882,I384847,);
nor I_22506 (I384862,I385106,I385007);
nand I_22507 (I385159,I111776,I111791);
and I_22508 (I385176,I385159,I111788);
DFFARX1 I_22509 (I385176,I2507,I384882,I385202,);
nor I_22510 (I384850,I385202,I385106);
not I_22511 (I385224,I385202);
nor I_22512 (I385241,I385224,I385015);
nor I_22513 (I385258,I384947,I385241);
DFFARX1 I_22514 (I385258,I2507,I384882,I384865,);
nor I_22515 (I385289,I385224,I385106);
nor I_22516 (I385306,I111800,I111791);
nor I_22517 (I384856,I385306,I385289);
not I_22518 (I385337,I385306);
nand I_22519 (I384859,I385066,I385337);
DFFARX1 I_22520 (I385306,I2507,I384882,I384871,);
DFFARX1 I_22521 (I385306,I2507,I384882,I384868,);
not I_22522 (I385426,I2514);
DFFARX1 I_22523 (I1363649,I2507,I385426,I385452,);
DFFARX1 I_22524 (I385452,I2507,I385426,I385469,);
not I_22525 (I385418,I385469);
not I_22526 (I385491,I385452);
nand I_22527 (I385508,I1363625,I1363646);
and I_22528 (I385525,I385508,I1363643);
DFFARX1 I_22529 (I385525,I2507,I385426,I385551,);
not I_22530 (I385559,I385551);
DFFARX1 I_22531 (I1363622,I2507,I385426,I385585,);
and I_22532 (I385593,I385585,I1363634);
nand I_22533 (I385610,I385585,I1363634);
nand I_22534 (I385397,I385559,I385610);
DFFARX1 I_22535 (I1363637,I2507,I385426,I385650,);
nor I_22536 (I385658,I385650,I385593);
DFFARX1 I_22537 (I385658,I2507,I385426,I385391,);
nor I_22538 (I385406,I385650,I385551);
nand I_22539 (I385703,I1363640,I1363628);
and I_22540 (I385720,I385703,I1363631);
DFFARX1 I_22541 (I385720,I2507,I385426,I385746,);
nor I_22542 (I385394,I385746,I385650);
not I_22543 (I385768,I385746);
nor I_22544 (I385785,I385768,I385559);
nor I_22545 (I385802,I385491,I385785);
DFFARX1 I_22546 (I385802,I2507,I385426,I385409,);
nor I_22547 (I385833,I385768,I385650);
nor I_22548 (I385850,I1363622,I1363628);
nor I_22549 (I385400,I385850,I385833);
not I_22550 (I385881,I385850);
nand I_22551 (I385403,I385610,I385881);
DFFARX1 I_22552 (I385850,I2507,I385426,I385415,);
DFFARX1 I_22553 (I385850,I2507,I385426,I385412,);
not I_22554 (I385970,I2514);
DFFARX1 I_22555 (I819651,I2507,I385970,I385996,);
DFFARX1 I_22556 (I385996,I2507,I385970,I386013,);
not I_22557 (I385962,I386013);
not I_22558 (I386035,I385996);
nand I_22559 (I386052,I819645,I819642);
and I_22560 (I386069,I386052,I819657);
DFFARX1 I_22561 (I386069,I2507,I385970,I386095,);
not I_22562 (I386103,I386095);
DFFARX1 I_22563 (I819645,I2507,I385970,I386129,);
and I_22564 (I386137,I386129,I819639);
nand I_22565 (I386154,I386129,I819639);
nand I_22566 (I385941,I386103,I386154);
DFFARX1 I_22567 (I819639,I2507,I385970,I386194,);
nor I_22568 (I386202,I386194,I386137);
DFFARX1 I_22569 (I386202,I2507,I385970,I385935,);
nor I_22570 (I385950,I386194,I386095);
nand I_22571 (I386247,I819654,I819648);
and I_22572 (I386264,I386247,I819642);
DFFARX1 I_22573 (I386264,I2507,I385970,I386290,);
nor I_22574 (I385938,I386290,I386194);
not I_22575 (I386312,I386290);
nor I_22576 (I386329,I386312,I386103);
nor I_22577 (I386346,I386035,I386329);
DFFARX1 I_22578 (I386346,I2507,I385970,I385953,);
nor I_22579 (I386377,I386312,I386194);
nor I_22580 (I386394,I819660,I819648);
nor I_22581 (I385944,I386394,I386377);
not I_22582 (I386425,I386394);
nand I_22583 (I385947,I386154,I386425);
DFFARX1 I_22584 (I386394,I2507,I385970,I385959,);
DFFARX1 I_22585 (I386394,I2507,I385970,I385956,);
not I_22586 (I386514,I2514);
DFFARX1 I_22587 (I191889,I2507,I386514,I386540,);
DFFARX1 I_22588 (I386540,I2507,I386514,I386557,);
not I_22589 (I386506,I386557);
not I_22590 (I386579,I386540);
nand I_22591 (I386596,I191901,I191880);
and I_22592 (I386613,I386596,I191883);
DFFARX1 I_22593 (I386613,I2507,I386514,I386639,);
not I_22594 (I386647,I386639);
DFFARX1 I_22595 (I191892,I2507,I386514,I386673,);
and I_22596 (I386681,I386673,I191904);
nand I_22597 (I386698,I386673,I191904);
nand I_22598 (I386485,I386647,I386698);
DFFARX1 I_22599 (I191898,I2507,I386514,I386738,);
nor I_22600 (I386746,I386738,I386681);
DFFARX1 I_22601 (I386746,I2507,I386514,I386479,);
nor I_22602 (I386494,I386738,I386639);
nand I_22603 (I386791,I191886,I191883);
and I_22604 (I386808,I386791,I191895);
DFFARX1 I_22605 (I386808,I2507,I386514,I386834,);
nor I_22606 (I386482,I386834,I386738);
not I_22607 (I386856,I386834);
nor I_22608 (I386873,I386856,I386647);
nor I_22609 (I386890,I386579,I386873);
DFFARX1 I_22610 (I386890,I2507,I386514,I386497,);
nor I_22611 (I386921,I386856,I386738);
nor I_22612 (I386938,I191880,I191883);
nor I_22613 (I386488,I386938,I386921);
not I_22614 (I386969,I386938);
nand I_22615 (I386491,I386698,I386969);
DFFARX1 I_22616 (I386938,I2507,I386514,I386503,);
DFFARX1 I_22617 (I386938,I2507,I386514,I386500,);
not I_22618 (I387058,I2514);
DFFARX1 I_22619 (I1060107,I2507,I387058,I387084,);
DFFARX1 I_22620 (I387084,I2507,I387058,I387101,);
not I_22621 (I387050,I387101);
not I_22622 (I387123,I387084);
nand I_22623 (I387140,I1060119,I1060107);
and I_22624 (I387157,I387140,I1060110);
DFFARX1 I_22625 (I387157,I2507,I387058,I387183,);
not I_22626 (I387191,I387183);
DFFARX1 I_22627 (I1060128,I2507,I387058,I387217,);
and I_22628 (I387225,I387217,I1060104);
nand I_22629 (I387242,I387217,I1060104);
nand I_22630 (I387029,I387191,I387242);
DFFARX1 I_22631 (I1060122,I2507,I387058,I387282,);
nor I_22632 (I387290,I387282,I387225);
DFFARX1 I_22633 (I387290,I2507,I387058,I387023,);
nor I_22634 (I387038,I387282,I387183);
nand I_22635 (I387335,I1060116,I1060113);
and I_22636 (I387352,I387335,I1060125);
DFFARX1 I_22637 (I387352,I2507,I387058,I387378,);
nor I_22638 (I387026,I387378,I387282);
not I_22639 (I387400,I387378);
nor I_22640 (I387417,I387400,I387191);
nor I_22641 (I387434,I387123,I387417);
DFFARX1 I_22642 (I387434,I2507,I387058,I387041,);
nor I_22643 (I387465,I387400,I387282);
nor I_22644 (I387482,I1060104,I1060113);
nor I_22645 (I387032,I387482,I387465);
not I_22646 (I387513,I387482);
nand I_22647 (I387035,I387242,I387513);
DFFARX1 I_22648 (I387482,I2507,I387058,I387047,);
DFFARX1 I_22649 (I387482,I2507,I387058,I387044,);
not I_22650 (I387602,I2514);
DFFARX1 I_22651 (I291844,I2507,I387602,I387628,);
DFFARX1 I_22652 (I387628,I2507,I387602,I387645,);
not I_22653 (I387594,I387645);
not I_22654 (I387667,I387628);
nand I_22655 (I387684,I291823,I291847);
and I_22656 (I387701,I387684,I291850);
DFFARX1 I_22657 (I387701,I2507,I387602,I387727,);
not I_22658 (I387735,I387727);
DFFARX1 I_22659 (I291832,I2507,I387602,I387761,);
and I_22660 (I387769,I387761,I291838);
nand I_22661 (I387786,I387761,I291838);
nand I_22662 (I387573,I387735,I387786);
DFFARX1 I_22663 (I291826,I2507,I387602,I387826,);
nor I_22664 (I387834,I387826,I387769);
DFFARX1 I_22665 (I387834,I2507,I387602,I387567,);
nor I_22666 (I387582,I387826,I387727);
nand I_22667 (I387879,I291835,I291823);
and I_22668 (I387896,I387879,I291829);
DFFARX1 I_22669 (I387896,I2507,I387602,I387922,);
nor I_22670 (I387570,I387922,I387826);
not I_22671 (I387944,I387922);
nor I_22672 (I387961,I387944,I387735);
nor I_22673 (I387978,I387667,I387961);
DFFARX1 I_22674 (I387978,I2507,I387602,I387585,);
nor I_22675 (I388009,I387944,I387826);
nor I_22676 (I388026,I291841,I291823);
nor I_22677 (I387576,I388026,I388009);
not I_22678 (I388057,I388026);
nand I_22679 (I387579,I387786,I388057);
DFFARX1 I_22680 (I388026,I2507,I387602,I387591,);
DFFARX1 I_22681 (I388026,I2507,I387602,I387588,);
not I_22682 (I388146,I2514);
DFFARX1 I_22683 (I1275580,I2507,I388146,I388172,);
DFFARX1 I_22684 (I388172,I2507,I388146,I388189,);
not I_22685 (I388138,I388189);
not I_22686 (I388211,I388172);
nand I_22687 (I388228,I1275577,I1275574);
and I_22688 (I388245,I388228,I1275562);
DFFARX1 I_22689 (I388245,I2507,I388146,I388271,);
not I_22690 (I388279,I388271);
DFFARX1 I_22691 (I1275586,I2507,I388146,I388305,);
and I_22692 (I388313,I388305,I1275571);
nand I_22693 (I388330,I388305,I1275571);
nand I_22694 (I388117,I388279,I388330);
DFFARX1 I_22695 (I1275565,I2507,I388146,I388370,);
nor I_22696 (I388378,I388370,I388313);
DFFARX1 I_22697 (I388378,I2507,I388146,I388111,);
nor I_22698 (I388126,I388370,I388271);
nand I_22699 (I388423,I1275562,I1275568);
and I_22700 (I388440,I388423,I1275583);
DFFARX1 I_22701 (I388440,I2507,I388146,I388466,);
nor I_22702 (I388114,I388466,I388370);
not I_22703 (I388488,I388466);
nor I_22704 (I388505,I388488,I388279);
nor I_22705 (I388522,I388211,I388505);
DFFARX1 I_22706 (I388522,I2507,I388146,I388129,);
nor I_22707 (I388553,I388488,I388370);
nor I_22708 (I388570,I1275565,I1275568);
nor I_22709 (I388120,I388570,I388553);
not I_22710 (I388601,I388570);
nand I_22711 (I388123,I388330,I388601);
DFFARX1 I_22712 (I388570,I2507,I388146,I388135,);
DFFARX1 I_22713 (I388570,I2507,I388146,I388132,);
not I_22714 (I388690,I2514);
DFFARX1 I_22715 (I939257,I2507,I388690,I388716,);
DFFARX1 I_22716 (I388716,I2507,I388690,I388733,);
not I_22717 (I388682,I388733);
not I_22718 (I388755,I388716);
nand I_22719 (I388772,I939272,I939260);
and I_22720 (I388789,I388772,I939251);
DFFARX1 I_22721 (I388789,I2507,I388690,I388815,);
not I_22722 (I388823,I388815);
DFFARX1 I_22723 (I939263,I2507,I388690,I388849,);
and I_22724 (I388857,I388849,I939254);
nand I_22725 (I388874,I388849,I939254);
nand I_22726 (I388661,I388823,I388874);
DFFARX1 I_22727 (I939269,I2507,I388690,I388914,);
nor I_22728 (I388922,I388914,I388857);
DFFARX1 I_22729 (I388922,I2507,I388690,I388655,);
nor I_22730 (I388670,I388914,I388815);
nand I_22731 (I388967,I939278,I939266);
and I_22732 (I388984,I388967,I939275);
DFFARX1 I_22733 (I388984,I2507,I388690,I389010,);
nor I_22734 (I388658,I389010,I388914);
not I_22735 (I389032,I389010);
nor I_22736 (I389049,I389032,I388823);
nor I_22737 (I389066,I388755,I389049);
DFFARX1 I_22738 (I389066,I2507,I388690,I388673,);
nor I_22739 (I389097,I389032,I388914);
nor I_22740 (I389114,I939251,I939266);
nor I_22741 (I388664,I389114,I389097);
not I_22742 (I389145,I389114);
nand I_22743 (I388667,I388874,I389145);
DFFARX1 I_22744 (I389114,I2507,I388690,I388679,);
DFFARX1 I_22745 (I389114,I2507,I388690,I388676,);
not I_22746 (I389234,I2514);
DFFARX1 I_22747 (I348760,I2507,I389234,I389260,);
DFFARX1 I_22748 (I389260,I2507,I389234,I389277,);
not I_22749 (I389226,I389277);
not I_22750 (I389299,I389260);
nand I_22751 (I389316,I348739,I348763);
and I_22752 (I389333,I389316,I348766);
DFFARX1 I_22753 (I389333,I2507,I389234,I389359,);
not I_22754 (I389367,I389359);
DFFARX1 I_22755 (I348748,I2507,I389234,I389393,);
and I_22756 (I389401,I389393,I348754);
nand I_22757 (I389418,I389393,I348754);
nand I_22758 (I389205,I389367,I389418);
DFFARX1 I_22759 (I348742,I2507,I389234,I389458,);
nor I_22760 (I389466,I389458,I389401);
DFFARX1 I_22761 (I389466,I2507,I389234,I389199,);
nor I_22762 (I389214,I389458,I389359);
nand I_22763 (I389511,I348751,I348739);
and I_22764 (I389528,I389511,I348745);
DFFARX1 I_22765 (I389528,I2507,I389234,I389554,);
nor I_22766 (I389202,I389554,I389458);
not I_22767 (I389576,I389554);
nor I_22768 (I389593,I389576,I389367);
nor I_22769 (I389610,I389299,I389593);
DFFARX1 I_22770 (I389610,I2507,I389234,I389217,);
nor I_22771 (I389641,I389576,I389458);
nor I_22772 (I389658,I348757,I348739);
nor I_22773 (I389208,I389658,I389641);
not I_22774 (I389689,I389658);
nand I_22775 (I389211,I389418,I389689);
DFFARX1 I_22776 (I389658,I2507,I389234,I389223,);
DFFARX1 I_22777 (I389658,I2507,I389234,I389220,);
not I_22778 (I389778,I2514);
DFFARX1 I_22779 (I4320,I2507,I389778,I389804,);
DFFARX1 I_22780 (I389804,I2507,I389778,I389821,);
not I_22781 (I389770,I389821);
not I_22782 (I389843,I389804);
nand I_22783 (I389860,I4323,I4311);
and I_22784 (I389877,I389860,I4317);
DFFARX1 I_22785 (I389877,I2507,I389778,I389903,);
not I_22786 (I389911,I389903);
DFFARX1 I_22787 (I4305,I2507,I389778,I389937,);
and I_22788 (I389945,I389937,I4302);
nand I_22789 (I389962,I389937,I4302);
nand I_22790 (I389749,I389911,I389962);
DFFARX1 I_22791 (I4308,I2507,I389778,I390002,);
nor I_22792 (I390010,I390002,I389945);
DFFARX1 I_22793 (I390010,I2507,I389778,I389743,);
nor I_22794 (I389758,I390002,I389903);
nand I_22795 (I390055,I4308,I4305);
and I_22796 (I390072,I390055,I4302);
DFFARX1 I_22797 (I390072,I2507,I389778,I390098,);
nor I_22798 (I389746,I390098,I390002);
not I_22799 (I390120,I390098);
nor I_22800 (I390137,I390120,I389911);
nor I_22801 (I390154,I389843,I390137);
DFFARX1 I_22802 (I390154,I2507,I389778,I389761,);
nor I_22803 (I390185,I390120,I390002);
nor I_22804 (I390202,I4314,I4305);
nor I_22805 (I389752,I390202,I390185);
not I_22806 (I390233,I390202);
nand I_22807 (I389755,I389962,I390233);
DFFARX1 I_22808 (I390202,I2507,I389778,I389767,);
DFFARX1 I_22809 (I390202,I2507,I389778,I389764,);
not I_22810 (I390322,I2514);
DFFARX1 I_22811 (I204384,I2507,I390322,I390348,);
DFFARX1 I_22812 (I390348,I2507,I390322,I390365,);
not I_22813 (I390314,I390365);
not I_22814 (I390387,I390348);
nand I_22815 (I390404,I204396,I204375);
and I_22816 (I390421,I390404,I204378);
DFFARX1 I_22817 (I390421,I2507,I390322,I390447,);
not I_22818 (I390455,I390447);
DFFARX1 I_22819 (I204387,I2507,I390322,I390481,);
and I_22820 (I390489,I390481,I204399);
nand I_22821 (I390506,I390481,I204399);
nand I_22822 (I390293,I390455,I390506);
DFFARX1 I_22823 (I204393,I2507,I390322,I390546,);
nor I_22824 (I390554,I390546,I390489);
DFFARX1 I_22825 (I390554,I2507,I390322,I390287,);
nor I_22826 (I390302,I390546,I390447);
nand I_22827 (I390599,I204381,I204378);
and I_22828 (I390616,I390599,I204390);
DFFARX1 I_22829 (I390616,I2507,I390322,I390642,);
nor I_22830 (I390290,I390642,I390546);
not I_22831 (I390664,I390642);
nor I_22832 (I390681,I390664,I390455);
nor I_22833 (I390698,I390387,I390681);
DFFARX1 I_22834 (I390698,I2507,I390322,I390305,);
nor I_22835 (I390729,I390664,I390546);
nor I_22836 (I390746,I204375,I204378);
nor I_22837 (I390296,I390746,I390729);
not I_22838 (I390777,I390746);
nand I_22839 (I390299,I390506,I390777);
DFFARX1 I_22840 (I390746,I2507,I390322,I390311,);
DFFARX1 I_22841 (I390746,I2507,I390322,I390308,);
not I_22842 (I390866,I2514);
DFFARX1 I_22843 (I912771,I2507,I390866,I390892,);
DFFARX1 I_22844 (I390892,I2507,I390866,I390909,);
not I_22845 (I390858,I390909);
not I_22846 (I390931,I390892);
nand I_22847 (I390948,I912786,I912774);
and I_22848 (I390965,I390948,I912765);
DFFARX1 I_22849 (I390965,I2507,I390866,I390991,);
not I_22850 (I390999,I390991);
DFFARX1 I_22851 (I912777,I2507,I390866,I391025,);
and I_22852 (I391033,I391025,I912768);
nand I_22853 (I391050,I391025,I912768);
nand I_22854 (I390837,I390999,I391050);
DFFARX1 I_22855 (I912783,I2507,I390866,I391090,);
nor I_22856 (I391098,I391090,I391033);
DFFARX1 I_22857 (I391098,I2507,I390866,I390831,);
nor I_22858 (I390846,I391090,I390991);
nand I_22859 (I391143,I912792,I912780);
and I_22860 (I391160,I391143,I912789);
DFFARX1 I_22861 (I391160,I2507,I390866,I391186,);
nor I_22862 (I390834,I391186,I391090);
not I_22863 (I391208,I391186);
nor I_22864 (I391225,I391208,I390999);
nor I_22865 (I391242,I390931,I391225);
DFFARX1 I_22866 (I391242,I2507,I390866,I390849,);
nor I_22867 (I391273,I391208,I391090);
nor I_22868 (I391290,I912765,I912780);
nor I_22869 (I390840,I391290,I391273);
not I_22870 (I391321,I391290);
nand I_22871 (I390843,I391050,I391321);
DFFARX1 I_22872 (I391290,I2507,I390866,I390855,);
DFFARX1 I_22873 (I391290,I2507,I390866,I390852,);
not I_22874 (I391410,I2514);
DFFARX1 I_22875 (I1302556,I2507,I391410,I391436,);
DFFARX1 I_22876 (I391436,I2507,I391410,I391453,);
not I_22877 (I391402,I391453);
not I_22878 (I391475,I391436);
nand I_22879 (I391492,I1302562,I1302565);
and I_22880 (I391509,I391492,I1302541);
DFFARX1 I_22881 (I391509,I2507,I391410,I391535,);
not I_22882 (I391543,I391535);
DFFARX1 I_22883 (I1302568,I2507,I391410,I391569,);
and I_22884 (I391577,I391569,I1302550);
nand I_22885 (I391594,I391569,I1302550);
nand I_22886 (I391381,I391543,I391594);
DFFARX1 I_22887 (I1302547,I2507,I391410,I391634,);
nor I_22888 (I391642,I391634,I391577);
DFFARX1 I_22889 (I391642,I2507,I391410,I391375,);
nor I_22890 (I391390,I391634,I391535);
nand I_22891 (I391687,I1302544,I1302553);
and I_22892 (I391704,I391687,I1302559);
DFFARX1 I_22893 (I391704,I2507,I391410,I391730,);
nor I_22894 (I391378,I391730,I391634);
not I_22895 (I391752,I391730);
nor I_22896 (I391769,I391752,I391543);
nor I_22897 (I391786,I391475,I391769);
DFFARX1 I_22898 (I391786,I2507,I391410,I391393,);
nor I_22899 (I391817,I391752,I391634);
nor I_22900 (I391834,I1302541,I1302553);
nor I_22901 (I391384,I391834,I391817);
not I_22902 (I391865,I391834);
nand I_22903 (I391387,I391594,I391865);
DFFARX1 I_22904 (I391834,I2507,I391410,I391399,);
DFFARX1 I_22905 (I391834,I2507,I391410,I391396,);
not I_22906 (I391954,I2514);
DFFARX1 I_22907 (I745743,I2507,I391954,I391980,);
DFFARX1 I_22908 (I391980,I2507,I391954,I391997,);
not I_22909 (I391946,I391997);
not I_22910 (I392019,I391980);
nand I_22911 (I392036,I745764,I745755);
and I_22912 (I392053,I392036,I745743);
DFFARX1 I_22913 (I392053,I2507,I391954,I392079,);
not I_22914 (I392087,I392079);
DFFARX1 I_22915 (I745749,I2507,I391954,I392113,);
and I_22916 (I392121,I392113,I745746);
nand I_22917 (I392138,I392113,I745746);
nand I_22918 (I391925,I392087,I392138);
DFFARX1 I_22919 (I745740,I2507,I391954,I392178,);
nor I_22920 (I392186,I392178,I392121);
DFFARX1 I_22921 (I392186,I2507,I391954,I391919,);
nor I_22922 (I391934,I392178,I392079);
nand I_22923 (I392231,I745740,I745752);
and I_22924 (I392248,I392231,I745761);
DFFARX1 I_22925 (I392248,I2507,I391954,I392274,);
nor I_22926 (I391922,I392274,I392178);
not I_22927 (I392296,I392274);
nor I_22928 (I392313,I392296,I392087);
nor I_22929 (I392330,I392019,I392313);
DFFARX1 I_22930 (I392330,I2507,I391954,I391937,);
nor I_22931 (I392361,I392296,I392178);
nor I_22932 (I392378,I745758,I745752);
nor I_22933 (I391928,I392378,I392361);
not I_22934 (I392409,I392378);
nand I_22935 (I391931,I392138,I392409);
DFFARX1 I_22936 (I392378,I2507,I391954,I391943,);
DFFARX1 I_22937 (I392378,I2507,I391954,I391940,);
not I_22938 (I392498,I2514);
DFFARX1 I_22939 (I582747,I2507,I392498,I392524,);
DFFARX1 I_22940 (I392524,I2507,I392498,I392541,);
not I_22941 (I392490,I392541);
not I_22942 (I392563,I392524);
nand I_22943 (I392580,I582744,I582765);
and I_22944 (I392597,I392580,I582768);
DFFARX1 I_22945 (I392597,I2507,I392498,I392623,);
not I_22946 (I392631,I392623);
DFFARX1 I_22947 (I582753,I2507,I392498,I392657,);
and I_22948 (I392665,I392657,I582756);
nand I_22949 (I392682,I392657,I582756);
nand I_22950 (I392469,I392631,I392682);
DFFARX1 I_22951 (I582759,I2507,I392498,I392722,);
nor I_22952 (I392730,I392722,I392665);
DFFARX1 I_22953 (I392730,I2507,I392498,I392463,);
nor I_22954 (I392478,I392722,I392623);
nand I_22955 (I392775,I582744,I582750);
and I_22956 (I392792,I392775,I582762);
DFFARX1 I_22957 (I392792,I2507,I392498,I392818,);
nor I_22958 (I392466,I392818,I392722);
not I_22959 (I392840,I392818);
nor I_22960 (I392857,I392840,I392631);
nor I_22961 (I392874,I392563,I392857);
DFFARX1 I_22962 (I392874,I2507,I392498,I392481,);
nor I_22963 (I392905,I392840,I392722);
nor I_22964 (I392922,I582747,I582750);
nor I_22965 (I392472,I392922,I392905);
not I_22966 (I392953,I392922);
nand I_22967 (I392475,I392682,I392953);
DFFARX1 I_22968 (I392922,I2507,I392498,I392487,);
DFFARX1 I_22969 (I392922,I2507,I392498,I392484,);
not I_22970 (I393042,I2514);
DFFARX1 I_22971 (I667135,I2507,I393042,I393068,);
DFFARX1 I_22972 (I393068,I2507,I393042,I393085,);
not I_22973 (I393034,I393085);
not I_22974 (I393107,I393068);
nand I_22975 (I393124,I667156,I667147);
and I_22976 (I393141,I393124,I667135);
DFFARX1 I_22977 (I393141,I2507,I393042,I393167,);
not I_22978 (I393175,I393167);
DFFARX1 I_22979 (I667141,I2507,I393042,I393201,);
and I_22980 (I393209,I393201,I667138);
nand I_22981 (I393226,I393201,I667138);
nand I_22982 (I393013,I393175,I393226);
DFFARX1 I_22983 (I667132,I2507,I393042,I393266,);
nor I_22984 (I393274,I393266,I393209);
DFFARX1 I_22985 (I393274,I2507,I393042,I393007,);
nor I_22986 (I393022,I393266,I393167);
nand I_22987 (I393319,I667132,I667144);
and I_22988 (I393336,I393319,I667153);
DFFARX1 I_22989 (I393336,I2507,I393042,I393362,);
nor I_22990 (I393010,I393362,I393266);
not I_22991 (I393384,I393362);
nor I_22992 (I393401,I393384,I393175);
nor I_22993 (I393418,I393107,I393401);
DFFARX1 I_22994 (I393418,I2507,I393042,I393025,);
nor I_22995 (I393449,I393384,I393266);
nor I_22996 (I393466,I667150,I667144);
nor I_22997 (I393016,I393466,I393449);
not I_22998 (I393497,I393466);
nand I_22999 (I393019,I393226,I393497);
DFFARX1 I_23000 (I393466,I2507,I393042,I393031,);
DFFARX1 I_23001 (I393466,I2507,I393042,I393028,);
not I_23002 (I393586,I2514);
DFFARX1 I_23003 (I1120797,I2507,I393586,I393612,);
DFFARX1 I_23004 (I393612,I2507,I393586,I393629,);
not I_23005 (I393578,I393629);
not I_23006 (I393651,I393612);
nand I_23007 (I393668,I1120809,I1120797);
and I_23008 (I393685,I393668,I1120800);
DFFARX1 I_23009 (I393685,I2507,I393586,I393711,);
not I_23010 (I393719,I393711);
DFFARX1 I_23011 (I1120818,I2507,I393586,I393745,);
and I_23012 (I393753,I393745,I1120794);
nand I_23013 (I393770,I393745,I1120794);
nand I_23014 (I393557,I393719,I393770);
DFFARX1 I_23015 (I1120812,I2507,I393586,I393810,);
nor I_23016 (I393818,I393810,I393753);
DFFARX1 I_23017 (I393818,I2507,I393586,I393551,);
nor I_23018 (I393566,I393810,I393711);
nand I_23019 (I393863,I1120806,I1120803);
and I_23020 (I393880,I393863,I1120815);
DFFARX1 I_23021 (I393880,I2507,I393586,I393906,);
nor I_23022 (I393554,I393906,I393810);
not I_23023 (I393928,I393906);
nor I_23024 (I393945,I393928,I393719);
nor I_23025 (I393962,I393651,I393945);
DFFARX1 I_23026 (I393962,I2507,I393586,I393569,);
nor I_23027 (I393993,I393928,I393810);
nor I_23028 (I394010,I1120794,I1120803);
nor I_23029 (I393560,I394010,I393993);
not I_23030 (I394041,I394010);
nand I_23031 (I393563,I393770,I394041);
DFFARX1 I_23032 (I394010,I2507,I393586,I393575,);
DFFARX1 I_23033 (I394010,I2507,I393586,I393572,);
not I_23034 (I394130,I2514);
DFFARX1 I_23035 (I970265,I2507,I394130,I394156,);
DFFARX1 I_23036 (I394156,I2507,I394130,I394173,);
not I_23037 (I394122,I394173);
not I_23038 (I394195,I394156);
nand I_23039 (I394212,I970280,I970268);
and I_23040 (I394229,I394212,I970259);
DFFARX1 I_23041 (I394229,I2507,I394130,I394255,);
not I_23042 (I394263,I394255);
DFFARX1 I_23043 (I970271,I2507,I394130,I394289,);
and I_23044 (I394297,I394289,I970262);
nand I_23045 (I394314,I394289,I970262);
nand I_23046 (I394101,I394263,I394314);
DFFARX1 I_23047 (I970277,I2507,I394130,I394354,);
nor I_23048 (I394362,I394354,I394297);
DFFARX1 I_23049 (I394362,I2507,I394130,I394095,);
nor I_23050 (I394110,I394354,I394255);
nand I_23051 (I394407,I970286,I970274);
and I_23052 (I394424,I394407,I970283);
DFFARX1 I_23053 (I394424,I2507,I394130,I394450,);
nor I_23054 (I394098,I394450,I394354);
not I_23055 (I394472,I394450);
nor I_23056 (I394489,I394472,I394263);
nor I_23057 (I394506,I394195,I394489);
DFFARX1 I_23058 (I394506,I2507,I394130,I394113,);
nor I_23059 (I394537,I394472,I394354);
nor I_23060 (I394554,I970259,I970274);
nor I_23061 (I394104,I394554,I394537);
not I_23062 (I394585,I394554);
nand I_23063 (I394107,I394314,I394585);
DFFARX1 I_23064 (I394554,I2507,I394130,I394119,);
DFFARX1 I_23065 (I394554,I2507,I394130,I394116,);
not I_23066 (I394674,I2514);
DFFARX1 I_23067 (I1357104,I2507,I394674,I394700,);
DFFARX1 I_23068 (I394700,I2507,I394674,I394717,);
not I_23069 (I394666,I394717);
not I_23070 (I394739,I394700);
nand I_23071 (I394756,I1357080,I1357101);
and I_23072 (I394773,I394756,I1357098);
DFFARX1 I_23073 (I394773,I2507,I394674,I394799,);
not I_23074 (I394807,I394799);
DFFARX1 I_23075 (I1357077,I2507,I394674,I394833,);
and I_23076 (I394841,I394833,I1357089);
nand I_23077 (I394858,I394833,I1357089);
nand I_23078 (I394645,I394807,I394858);
DFFARX1 I_23079 (I1357092,I2507,I394674,I394898,);
nor I_23080 (I394906,I394898,I394841);
DFFARX1 I_23081 (I394906,I2507,I394674,I394639,);
nor I_23082 (I394654,I394898,I394799);
nand I_23083 (I394951,I1357095,I1357083);
and I_23084 (I394968,I394951,I1357086);
DFFARX1 I_23085 (I394968,I2507,I394674,I394994,);
nor I_23086 (I394642,I394994,I394898);
not I_23087 (I395016,I394994);
nor I_23088 (I395033,I395016,I394807);
nor I_23089 (I395050,I394739,I395033);
DFFARX1 I_23090 (I395050,I2507,I394674,I394657,);
nor I_23091 (I395081,I395016,I394898);
nor I_23092 (I395098,I1357077,I1357083);
nor I_23093 (I394648,I395098,I395081);
not I_23094 (I395129,I395098);
nand I_23095 (I394651,I394858,I395129);
DFFARX1 I_23096 (I395098,I2507,I394674,I394663,);
DFFARX1 I_23097 (I395098,I2507,I394674,I394660,);
not I_23098 (I395218,I2514);
DFFARX1 I_23099 (I735339,I2507,I395218,I395244,);
DFFARX1 I_23100 (I395244,I2507,I395218,I395261,);
not I_23101 (I395210,I395261);
not I_23102 (I395283,I395244);
nand I_23103 (I395300,I735360,I735351);
and I_23104 (I395317,I395300,I735339);
DFFARX1 I_23105 (I395317,I2507,I395218,I395343,);
not I_23106 (I395351,I395343);
DFFARX1 I_23107 (I735345,I2507,I395218,I395377,);
and I_23108 (I395385,I395377,I735342);
nand I_23109 (I395402,I395377,I735342);
nand I_23110 (I395189,I395351,I395402);
DFFARX1 I_23111 (I735336,I2507,I395218,I395442,);
nor I_23112 (I395450,I395442,I395385);
DFFARX1 I_23113 (I395450,I2507,I395218,I395183,);
nor I_23114 (I395198,I395442,I395343);
nand I_23115 (I395495,I735336,I735348);
and I_23116 (I395512,I395495,I735357);
DFFARX1 I_23117 (I395512,I2507,I395218,I395538,);
nor I_23118 (I395186,I395538,I395442);
not I_23119 (I395560,I395538);
nor I_23120 (I395577,I395560,I395351);
nor I_23121 (I395594,I395283,I395577);
DFFARX1 I_23122 (I395594,I2507,I395218,I395201,);
nor I_23123 (I395625,I395560,I395442);
nor I_23124 (I395642,I735354,I735348);
nor I_23125 (I395192,I395642,I395625);
not I_23126 (I395673,I395642);
nand I_23127 (I395195,I395402,I395673);
DFFARX1 I_23128 (I395642,I2507,I395218,I395207,);
DFFARX1 I_23129 (I395642,I2507,I395218,I395204,);
not I_23130 (I395762,I2514);
DFFARX1 I_23131 (I939903,I2507,I395762,I395788,);
DFFARX1 I_23132 (I395788,I2507,I395762,I395805,);
not I_23133 (I395754,I395805);
not I_23134 (I395827,I395788);
nand I_23135 (I395844,I939918,I939906);
and I_23136 (I395861,I395844,I939897);
DFFARX1 I_23137 (I395861,I2507,I395762,I395887,);
not I_23138 (I395895,I395887);
DFFARX1 I_23139 (I939909,I2507,I395762,I395921,);
and I_23140 (I395929,I395921,I939900);
nand I_23141 (I395946,I395921,I939900);
nand I_23142 (I395733,I395895,I395946);
DFFARX1 I_23143 (I939915,I2507,I395762,I395986,);
nor I_23144 (I395994,I395986,I395929);
DFFARX1 I_23145 (I395994,I2507,I395762,I395727,);
nor I_23146 (I395742,I395986,I395887);
nand I_23147 (I396039,I939924,I939912);
and I_23148 (I396056,I396039,I939921);
DFFARX1 I_23149 (I396056,I2507,I395762,I396082,);
nor I_23150 (I395730,I396082,I395986);
not I_23151 (I396104,I396082);
nor I_23152 (I396121,I396104,I395895);
nor I_23153 (I396138,I395827,I396121);
DFFARX1 I_23154 (I396138,I2507,I395762,I395745,);
nor I_23155 (I396169,I396104,I395986);
nor I_23156 (I396186,I939897,I939912);
nor I_23157 (I395736,I396186,I396169);
not I_23158 (I396217,I396186);
nand I_23159 (I395739,I395946,I396217);
DFFARX1 I_23160 (I396186,I2507,I395762,I395751,);
DFFARX1 I_23161 (I396186,I2507,I395762,I395748,);
not I_23162 (I396306,I2514);
DFFARX1 I_23163 (I1139871,I2507,I396306,I396332,);
DFFARX1 I_23164 (I396332,I2507,I396306,I396349,);
not I_23165 (I396298,I396349);
not I_23166 (I396371,I396332);
nand I_23167 (I396388,I1139883,I1139871);
and I_23168 (I396405,I396388,I1139874);
DFFARX1 I_23169 (I396405,I2507,I396306,I396431,);
not I_23170 (I396439,I396431);
DFFARX1 I_23171 (I1139892,I2507,I396306,I396465,);
and I_23172 (I396473,I396465,I1139868);
nand I_23173 (I396490,I396465,I1139868);
nand I_23174 (I396277,I396439,I396490);
DFFARX1 I_23175 (I1139886,I2507,I396306,I396530,);
nor I_23176 (I396538,I396530,I396473);
DFFARX1 I_23177 (I396538,I2507,I396306,I396271,);
nor I_23178 (I396286,I396530,I396431);
nand I_23179 (I396583,I1139880,I1139877);
and I_23180 (I396600,I396583,I1139889);
DFFARX1 I_23181 (I396600,I2507,I396306,I396626,);
nor I_23182 (I396274,I396626,I396530);
not I_23183 (I396648,I396626);
nor I_23184 (I396665,I396648,I396439);
nor I_23185 (I396682,I396371,I396665);
DFFARX1 I_23186 (I396682,I2507,I396306,I396289,);
nor I_23187 (I396713,I396648,I396530);
nor I_23188 (I396730,I1139868,I1139877);
nor I_23189 (I396280,I396730,I396713);
not I_23190 (I396761,I396730);
nand I_23191 (I396283,I396490,I396761);
DFFARX1 I_23192 (I396730,I2507,I396306,I396295,);
DFFARX1 I_23193 (I396730,I2507,I396306,I396292,);
not I_23194 (I396850,I2514);
DFFARX1 I_23195 (I985123,I2507,I396850,I396876,);
DFFARX1 I_23196 (I396876,I2507,I396850,I396893,);
not I_23197 (I396842,I396893);
not I_23198 (I396915,I396876);
nand I_23199 (I396932,I985138,I985126);
and I_23200 (I396949,I396932,I985117);
DFFARX1 I_23201 (I396949,I2507,I396850,I396975,);
not I_23202 (I396983,I396975);
DFFARX1 I_23203 (I985129,I2507,I396850,I397009,);
and I_23204 (I397017,I397009,I985120);
nand I_23205 (I397034,I397009,I985120);
nand I_23206 (I396821,I396983,I397034);
DFFARX1 I_23207 (I985135,I2507,I396850,I397074,);
nor I_23208 (I397082,I397074,I397017);
DFFARX1 I_23209 (I397082,I2507,I396850,I396815,);
nor I_23210 (I396830,I397074,I396975);
nand I_23211 (I397127,I985144,I985132);
and I_23212 (I397144,I397127,I985141);
DFFARX1 I_23213 (I397144,I2507,I396850,I397170,);
nor I_23214 (I396818,I397170,I397074);
not I_23215 (I397192,I397170);
nor I_23216 (I397209,I397192,I396983);
nor I_23217 (I397226,I396915,I397209);
DFFARX1 I_23218 (I397226,I2507,I396850,I396833,);
nor I_23219 (I397257,I397192,I397074);
nor I_23220 (I397274,I985117,I985132);
nor I_23221 (I396824,I397274,I397257);
not I_23222 (I397305,I397274);
nand I_23223 (I396827,I397034,I397305);
DFFARX1 I_23224 (I397274,I2507,I396850,I396839,);
DFFARX1 I_23225 (I397274,I2507,I396850,I396836,);
not I_23226 (I397394,I2514);
DFFARX1 I_23227 (I162139,I2507,I397394,I397420,);
DFFARX1 I_23228 (I397420,I2507,I397394,I397437,);
not I_23229 (I397386,I397437);
not I_23230 (I397459,I397420);
nand I_23231 (I397476,I162151,I162130);
and I_23232 (I397493,I397476,I162133);
DFFARX1 I_23233 (I397493,I2507,I397394,I397519,);
not I_23234 (I397527,I397519);
DFFARX1 I_23235 (I162142,I2507,I397394,I397553,);
and I_23236 (I397561,I397553,I162154);
nand I_23237 (I397578,I397553,I162154);
nand I_23238 (I397365,I397527,I397578);
DFFARX1 I_23239 (I162148,I2507,I397394,I397618,);
nor I_23240 (I397626,I397618,I397561);
DFFARX1 I_23241 (I397626,I2507,I397394,I397359,);
nor I_23242 (I397374,I397618,I397519);
nand I_23243 (I397671,I162136,I162133);
and I_23244 (I397688,I397671,I162145);
DFFARX1 I_23245 (I397688,I2507,I397394,I397714,);
nor I_23246 (I397362,I397714,I397618);
not I_23247 (I397736,I397714);
nor I_23248 (I397753,I397736,I397527);
nor I_23249 (I397770,I397459,I397753);
DFFARX1 I_23250 (I397770,I2507,I397394,I397377,);
nor I_23251 (I397801,I397736,I397618);
nor I_23252 (I397818,I162130,I162133);
nor I_23253 (I397368,I397818,I397801);
not I_23254 (I397849,I397818);
nand I_23255 (I397371,I397578,I397849);
DFFARX1 I_23256 (I397818,I2507,I397394,I397383,);
DFFARX1 I_23257 (I397818,I2507,I397394,I397380,);
not I_23258 (I397938,I2514);
DFFARX1 I_23259 (I706439,I2507,I397938,I397964,);
DFFARX1 I_23260 (I397964,I2507,I397938,I397981,);
not I_23261 (I397930,I397981);
not I_23262 (I398003,I397964);
nand I_23263 (I398020,I706460,I706451);
and I_23264 (I398037,I398020,I706439);
DFFARX1 I_23265 (I398037,I2507,I397938,I398063,);
not I_23266 (I398071,I398063);
DFFARX1 I_23267 (I706445,I2507,I397938,I398097,);
and I_23268 (I398105,I398097,I706442);
nand I_23269 (I398122,I398097,I706442);
nand I_23270 (I397909,I398071,I398122);
DFFARX1 I_23271 (I706436,I2507,I397938,I398162,);
nor I_23272 (I398170,I398162,I398105);
DFFARX1 I_23273 (I398170,I2507,I397938,I397903,);
nor I_23274 (I397918,I398162,I398063);
nand I_23275 (I398215,I706436,I706448);
and I_23276 (I398232,I398215,I706457);
DFFARX1 I_23277 (I398232,I2507,I397938,I398258,);
nor I_23278 (I397906,I398258,I398162);
not I_23279 (I398280,I398258);
nor I_23280 (I398297,I398280,I398071);
nor I_23281 (I398314,I398003,I398297);
DFFARX1 I_23282 (I398314,I2507,I397938,I397921,);
nor I_23283 (I398345,I398280,I398162);
nor I_23284 (I398362,I706454,I706448);
nor I_23285 (I397912,I398362,I398345);
not I_23286 (I398393,I398362);
nand I_23287 (I397915,I398122,I398393);
DFFARX1 I_23288 (I398362,I2507,I397938,I397927,);
DFFARX1 I_23289 (I398362,I2507,I397938,I397924,);
not I_23290 (I398482,I2514);
DFFARX1 I_23291 (I1390424,I2507,I398482,I398508,);
DFFARX1 I_23292 (I398508,I2507,I398482,I398525,);
not I_23293 (I398474,I398525);
not I_23294 (I398547,I398508);
nand I_23295 (I398564,I1390400,I1390421);
and I_23296 (I398581,I398564,I1390418);
DFFARX1 I_23297 (I398581,I2507,I398482,I398607,);
not I_23298 (I398615,I398607);
DFFARX1 I_23299 (I1390397,I2507,I398482,I398641,);
and I_23300 (I398649,I398641,I1390409);
nand I_23301 (I398666,I398641,I1390409);
nand I_23302 (I398453,I398615,I398666);
DFFARX1 I_23303 (I1390412,I2507,I398482,I398706,);
nor I_23304 (I398714,I398706,I398649);
DFFARX1 I_23305 (I398714,I2507,I398482,I398447,);
nor I_23306 (I398462,I398706,I398607);
nand I_23307 (I398759,I1390415,I1390403);
and I_23308 (I398776,I398759,I1390406);
DFFARX1 I_23309 (I398776,I2507,I398482,I398802,);
nor I_23310 (I398450,I398802,I398706);
not I_23311 (I398824,I398802);
nor I_23312 (I398841,I398824,I398615);
nor I_23313 (I398858,I398547,I398841);
DFFARX1 I_23314 (I398858,I2507,I398482,I398465,);
nor I_23315 (I398889,I398824,I398706);
nor I_23316 (I398906,I1390397,I1390403);
nor I_23317 (I398456,I398906,I398889);
not I_23318 (I398937,I398906);
nand I_23319 (I398459,I398666,I398937);
DFFARX1 I_23320 (I398906,I2507,I398482,I398471,);
DFFARX1 I_23321 (I398906,I2507,I398482,I398468,);
not I_23322 (I399026,I2514);
DFFARX1 I_23323 (I752679,I2507,I399026,I399052,);
DFFARX1 I_23324 (I399052,I2507,I399026,I399069,);
not I_23325 (I399018,I399069);
not I_23326 (I399091,I399052);
nand I_23327 (I399108,I752700,I752691);
and I_23328 (I399125,I399108,I752679);
DFFARX1 I_23329 (I399125,I2507,I399026,I399151,);
not I_23330 (I399159,I399151);
DFFARX1 I_23331 (I752685,I2507,I399026,I399185,);
and I_23332 (I399193,I399185,I752682);
nand I_23333 (I399210,I399185,I752682);
nand I_23334 (I398997,I399159,I399210);
DFFARX1 I_23335 (I752676,I2507,I399026,I399250,);
nor I_23336 (I399258,I399250,I399193);
DFFARX1 I_23337 (I399258,I2507,I399026,I398991,);
nor I_23338 (I399006,I399250,I399151);
nand I_23339 (I399303,I752676,I752688);
and I_23340 (I399320,I399303,I752697);
DFFARX1 I_23341 (I399320,I2507,I399026,I399346,);
nor I_23342 (I398994,I399346,I399250);
not I_23343 (I399368,I399346);
nor I_23344 (I399385,I399368,I399159);
nor I_23345 (I399402,I399091,I399385);
DFFARX1 I_23346 (I399402,I2507,I399026,I399009,);
nor I_23347 (I399433,I399368,I399250);
nor I_23348 (I399450,I752694,I752688);
nor I_23349 (I399000,I399450,I399433);
not I_23350 (I399481,I399450);
nand I_23351 (I399003,I399210,I399481);
DFFARX1 I_23352 (I399450,I2507,I399026,I399015,);
DFFARX1 I_23353 (I399450,I2507,I399026,I399012,);
not I_23354 (I399570,I2514);
DFFARX1 I_23355 (I881310,I2507,I399570,I399596,);
DFFARX1 I_23356 (I399596,I2507,I399570,I399613,);
not I_23357 (I399562,I399613);
not I_23358 (I399635,I399596);
nand I_23359 (I399652,I881304,I881301);
and I_23360 (I399669,I399652,I881316);
DFFARX1 I_23361 (I399669,I2507,I399570,I399695,);
not I_23362 (I399703,I399695);
DFFARX1 I_23363 (I881304,I2507,I399570,I399729,);
and I_23364 (I399737,I399729,I881298);
nand I_23365 (I399754,I399729,I881298);
nand I_23366 (I399541,I399703,I399754);
DFFARX1 I_23367 (I881298,I2507,I399570,I399794,);
nor I_23368 (I399802,I399794,I399737);
DFFARX1 I_23369 (I399802,I2507,I399570,I399535,);
nor I_23370 (I399550,I399794,I399695);
nand I_23371 (I399847,I881313,I881307);
and I_23372 (I399864,I399847,I881301);
DFFARX1 I_23373 (I399864,I2507,I399570,I399890,);
nor I_23374 (I399538,I399890,I399794);
not I_23375 (I399912,I399890);
nor I_23376 (I399929,I399912,I399703);
nor I_23377 (I399946,I399635,I399929);
DFFARX1 I_23378 (I399946,I2507,I399570,I399553,);
nor I_23379 (I399977,I399912,I399794);
nor I_23380 (I399994,I881319,I881307);
nor I_23381 (I399544,I399994,I399977);
not I_23382 (I400025,I399994);
nand I_23383 (I399547,I399754,I400025);
DFFARX1 I_23384 (I399994,I2507,I399570,I399559,);
DFFARX1 I_23385 (I399994,I2507,I399570,I399556,);
not I_23386 (I400114,I2514);
DFFARX1 I_23387 (I937319,I2507,I400114,I400140,);
DFFARX1 I_23388 (I400140,I2507,I400114,I400157,);
not I_23389 (I400106,I400157);
not I_23390 (I400179,I400140);
nand I_23391 (I400196,I937334,I937322);
and I_23392 (I400213,I400196,I937313);
DFFARX1 I_23393 (I400213,I2507,I400114,I400239,);
not I_23394 (I400247,I400239);
DFFARX1 I_23395 (I937325,I2507,I400114,I400273,);
and I_23396 (I400281,I400273,I937316);
nand I_23397 (I400298,I400273,I937316);
nand I_23398 (I400085,I400247,I400298);
DFFARX1 I_23399 (I937331,I2507,I400114,I400338,);
nor I_23400 (I400346,I400338,I400281);
DFFARX1 I_23401 (I400346,I2507,I400114,I400079,);
nor I_23402 (I400094,I400338,I400239);
nand I_23403 (I400391,I937340,I937328);
and I_23404 (I400408,I400391,I937337);
DFFARX1 I_23405 (I400408,I2507,I400114,I400434,);
nor I_23406 (I400082,I400434,I400338);
not I_23407 (I400456,I400434);
nor I_23408 (I400473,I400456,I400247);
nor I_23409 (I400490,I400179,I400473);
DFFARX1 I_23410 (I400490,I2507,I400114,I400097,);
nor I_23411 (I400521,I400456,I400338);
nor I_23412 (I400538,I937313,I937328);
nor I_23413 (I400088,I400538,I400521);
not I_23414 (I400569,I400538);
nand I_23415 (I400091,I400298,I400569);
DFFARX1 I_23416 (I400538,I2507,I400114,I400103,);
DFFARX1 I_23417 (I400538,I2507,I400114,I400100,);
not I_23418 (I400658,I2514);
DFFARX1 I_23419 (I1029215,I2507,I400658,I400684,);
DFFARX1 I_23420 (I400684,I2507,I400658,I400701,);
not I_23421 (I400650,I400701);
not I_23422 (I400723,I400684);
nand I_23423 (I400740,I1029215,I1029233);
and I_23424 (I400757,I400740,I1029227);
DFFARX1 I_23425 (I400757,I2507,I400658,I400783,);
not I_23426 (I400791,I400783);
DFFARX1 I_23427 (I1029221,I2507,I400658,I400817,);
and I_23428 (I400825,I400817,I1029230);
nand I_23429 (I400842,I400817,I1029230);
nand I_23430 (I400629,I400791,I400842);
DFFARX1 I_23431 (I1029218,I2507,I400658,I400882,);
nor I_23432 (I400890,I400882,I400825);
DFFARX1 I_23433 (I400890,I2507,I400658,I400623,);
nor I_23434 (I400638,I400882,I400783);
nand I_23435 (I400935,I1029218,I1029236);
and I_23436 (I400952,I400935,I1029221);
DFFARX1 I_23437 (I400952,I2507,I400658,I400978,);
nor I_23438 (I400626,I400978,I400882);
not I_23439 (I401000,I400978);
nor I_23440 (I401017,I401000,I400791);
nor I_23441 (I401034,I400723,I401017);
DFFARX1 I_23442 (I401034,I2507,I400658,I400641,);
nor I_23443 (I401065,I401000,I400882);
nor I_23444 (I401082,I1029224,I1029236);
nor I_23445 (I400632,I401082,I401065);
not I_23446 (I401113,I401082);
nand I_23447 (I400635,I400842,I401113);
DFFARX1 I_23448 (I401082,I2507,I400658,I400647,);
DFFARX1 I_23449 (I401082,I2507,I400658,I400644,);
not I_23450 (I401202,I2514);
DFFARX1 I_23451 (I42224,I2507,I401202,I401228,);
DFFARX1 I_23452 (I401228,I2507,I401202,I401245,);
not I_23453 (I401194,I401245);
not I_23454 (I401267,I401228);
nand I_23455 (I401284,I42212,I42227);
and I_23456 (I401301,I401284,I42215);
DFFARX1 I_23457 (I401301,I2507,I401202,I401327,);
not I_23458 (I401335,I401327);
DFFARX1 I_23459 (I42236,I2507,I401202,I401361,);
and I_23460 (I401369,I401361,I42230);
nand I_23461 (I401386,I401361,I42230);
nand I_23462 (I401173,I401335,I401386);
DFFARX1 I_23463 (I42233,I2507,I401202,I401426,);
nor I_23464 (I401434,I401426,I401369);
DFFARX1 I_23465 (I401434,I2507,I401202,I401167,);
nor I_23466 (I401182,I401426,I401327);
nand I_23467 (I401479,I42212,I42215);
and I_23468 (I401496,I401479,I42218);
DFFARX1 I_23469 (I401496,I2507,I401202,I401522,);
nor I_23470 (I401170,I401522,I401426);
not I_23471 (I401544,I401522);
nor I_23472 (I401561,I401544,I401335);
nor I_23473 (I401578,I401267,I401561);
DFFARX1 I_23474 (I401578,I2507,I401202,I401185,);
nor I_23475 (I401609,I401544,I401426);
nor I_23476 (I401626,I42221,I42215);
nor I_23477 (I401176,I401626,I401609);
not I_23478 (I401657,I401626);
nand I_23479 (I401179,I401386,I401657);
DFFARX1 I_23480 (I401626,I2507,I401202,I401191,);
DFFARX1 I_23481 (I401626,I2507,I401202,I401188,);
not I_23482 (I401746,I2514);
DFFARX1 I_23483 (I1201139,I2507,I401746,I401772,);
DFFARX1 I_23484 (I401772,I2507,I401746,I401789,);
not I_23485 (I401738,I401789);
not I_23486 (I401811,I401772);
nand I_23487 (I401828,I1201151,I1201139);
and I_23488 (I401845,I401828,I1201142);
DFFARX1 I_23489 (I401845,I2507,I401746,I401871,);
not I_23490 (I401879,I401871);
DFFARX1 I_23491 (I1201160,I2507,I401746,I401905,);
and I_23492 (I401913,I401905,I1201136);
nand I_23493 (I401930,I401905,I1201136);
nand I_23494 (I401717,I401879,I401930);
DFFARX1 I_23495 (I1201154,I2507,I401746,I401970,);
nor I_23496 (I401978,I401970,I401913);
DFFARX1 I_23497 (I401978,I2507,I401746,I401711,);
nor I_23498 (I401726,I401970,I401871);
nand I_23499 (I402023,I1201148,I1201145);
and I_23500 (I402040,I402023,I1201157);
DFFARX1 I_23501 (I402040,I2507,I401746,I402066,);
nor I_23502 (I401714,I402066,I401970);
not I_23503 (I402088,I402066);
nor I_23504 (I402105,I402088,I401879);
nor I_23505 (I402122,I401811,I402105);
DFFARX1 I_23506 (I402122,I2507,I401746,I401729,);
nor I_23507 (I402153,I402088,I401970);
nor I_23508 (I402170,I1201136,I1201145);
nor I_23509 (I401720,I402170,I402153);
not I_23510 (I402201,I402170);
nand I_23511 (I401723,I401930,I402201);
DFFARX1 I_23512 (I402170,I2507,I401746,I401735,);
DFFARX1 I_23513 (I402170,I2507,I401746,I401732,);
not I_23514 (I402290,I2514);
DFFARX1 I_23515 (I284993,I2507,I402290,I402316,);
DFFARX1 I_23516 (I402316,I2507,I402290,I402333,);
not I_23517 (I402282,I402333);
not I_23518 (I402355,I402316);
nand I_23519 (I402372,I284972,I284996);
and I_23520 (I402389,I402372,I284999);
DFFARX1 I_23521 (I402389,I2507,I402290,I402415,);
not I_23522 (I402423,I402415);
DFFARX1 I_23523 (I284981,I2507,I402290,I402449,);
and I_23524 (I402457,I402449,I284987);
nand I_23525 (I402474,I402449,I284987);
nand I_23526 (I402261,I402423,I402474);
DFFARX1 I_23527 (I284975,I2507,I402290,I402514,);
nor I_23528 (I402522,I402514,I402457);
DFFARX1 I_23529 (I402522,I2507,I402290,I402255,);
nor I_23530 (I402270,I402514,I402415);
nand I_23531 (I402567,I284984,I284972);
and I_23532 (I402584,I402567,I284978);
DFFARX1 I_23533 (I402584,I2507,I402290,I402610,);
nor I_23534 (I402258,I402610,I402514);
not I_23535 (I402632,I402610);
nor I_23536 (I402649,I402632,I402423);
nor I_23537 (I402666,I402355,I402649);
DFFARX1 I_23538 (I402666,I2507,I402290,I402273,);
nor I_23539 (I402697,I402632,I402514);
nor I_23540 (I402714,I284990,I284972);
nor I_23541 (I402264,I402714,I402697);
not I_23542 (I402745,I402714);
nand I_23543 (I402267,I402474,I402745);
DFFARX1 I_23544 (I402714,I2507,I402290,I402279,);
DFFARX1 I_23545 (I402714,I2507,I402290,I402276,);
not I_23546 (I402834,I2514);
DFFARX1 I_23547 (I1217765,I2507,I402834,I402860,);
DFFARX1 I_23548 (I402860,I2507,I402834,I402877,);
not I_23549 (I402826,I402877);
not I_23550 (I402899,I402860);
nand I_23551 (I402916,I1217777,I1217780);
and I_23552 (I402933,I402916,I1217783);
DFFARX1 I_23553 (I402933,I2507,I402834,I402959,);
not I_23554 (I402967,I402959);
DFFARX1 I_23555 (I1217768,I2507,I402834,I402993,);
and I_23556 (I403001,I402993,I1217774);
nand I_23557 (I403018,I402993,I1217774);
nand I_23558 (I402805,I402967,I403018);
DFFARX1 I_23559 (I1217762,I2507,I402834,I403058,);
nor I_23560 (I403066,I403058,I403001);
DFFARX1 I_23561 (I403066,I2507,I402834,I402799,);
nor I_23562 (I402814,I403058,I402959);
nand I_23563 (I403111,I1217765,I1217786);
and I_23564 (I403128,I403111,I1217771);
DFFARX1 I_23565 (I403128,I2507,I402834,I403154,);
nor I_23566 (I402802,I403154,I403058);
not I_23567 (I403176,I403154);
nor I_23568 (I403193,I403176,I402967);
nor I_23569 (I403210,I402899,I403193);
DFFARX1 I_23570 (I403210,I2507,I402834,I402817,);
nor I_23571 (I403241,I403176,I403058);
nor I_23572 (I403258,I1217762,I1217786);
nor I_23573 (I402808,I403258,I403241);
not I_23574 (I403289,I403258);
nand I_23575 (I402811,I403018,I403289);
DFFARX1 I_23576 (I403258,I2507,I402834,I402823,);
DFFARX1 I_23577 (I403258,I2507,I402834,I402820,);
not I_23578 (I403378,I2514);
DFFARX1 I_23579 (I879202,I2507,I403378,I403404,);
DFFARX1 I_23580 (I403404,I2507,I403378,I403421,);
not I_23581 (I403370,I403421);
not I_23582 (I403443,I403404);
nand I_23583 (I403460,I879196,I879193);
and I_23584 (I403477,I403460,I879208);
DFFARX1 I_23585 (I403477,I2507,I403378,I403503,);
not I_23586 (I403511,I403503);
DFFARX1 I_23587 (I879196,I2507,I403378,I403537,);
and I_23588 (I403545,I403537,I879190);
nand I_23589 (I403562,I403537,I879190);
nand I_23590 (I403349,I403511,I403562);
DFFARX1 I_23591 (I879190,I2507,I403378,I403602,);
nor I_23592 (I403610,I403602,I403545);
DFFARX1 I_23593 (I403610,I2507,I403378,I403343,);
nor I_23594 (I403358,I403602,I403503);
nand I_23595 (I403655,I879205,I879199);
and I_23596 (I403672,I403655,I879193);
DFFARX1 I_23597 (I403672,I2507,I403378,I403698,);
nor I_23598 (I403346,I403698,I403602);
not I_23599 (I403720,I403698);
nor I_23600 (I403737,I403720,I403511);
nor I_23601 (I403754,I403443,I403737);
DFFARX1 I_23602 (I403754,I2507,I403378,I403361,);
nor I_23603 (I403785,I403720,I403602);
nor I_23604 (I403802,I879211,I879199);
nor I_23605 (I403352,I403802,I403785);
not I_23606 (I403833,I403802);
nand I_23607 (I403355,I403562,I403833);
DFFARX1 I_23608 (I403802,I2507,I403378,I403367,);
DFFARX1 I_23609 (I403802,I2507,I403378,I403364,);
not I_23610 (I403922,I2514);
DFFARX1 I_23611 (I554425,I2507,I403922,I403948,);
DFFARX1 I_23612 (I403948,I2507,I403922,I403965,);
not I_23613 (I403914,I403965);
not I_23614 (I403987,I403948);
nand I_23615 (I404004,I554422,I554443);
and I_23616 (I404021,I404004,I554446);
DFFARX1 I_23617 (I404021,I2507,I403922,I404047,);
not I_23618 (I404055,I404047);
DFFARX1 I_23619 (I554431,I2507,I403922,I404081,);
and I_23620 (I404089,I404081,I554434);
nand I_23621 (I404106,I404081,I554434);
nand I_23622 (I403893,I404055,I404106);
DFFARX1 I_23623 (I554437,I2507,I403922,I404146,);
nor I_23624 (I404154,I404146,I404089);
DFFARX1 I_23625 (I404154,I2507,I403922,I403887,);
nor I_23626 (I403902,I404146,I404047);
nand I_23627 (I404199,I554422,I554428);
and I_23628 (I404216,I404199,I554440);
DFFARX1 I_23629 (I404216,I2507,I403922,I404242,);
nor I_23630 (I403890,I404242,I404146);
not I_23631 (I404264,I404242);
nor I_23632 (I404281,I404264,I404055);
nor I_23633 (I404298,I403987,I404281);
DFFARX1 I_23634 (I404298,I2507,I403922,I403905,);
nor I_23635 (I404329,I404264,I404146);
nor I_23636 (I404346,I554425,I554428);
nor I_23637 (I403896,I404346,I404329);
not I_23638 (I404377,I404346);
nand I_23639 (I403899,I404106,I404377);
DFFARX1 I_23640 (I404346,I2507,I403922,I403911,);
DFFARX1 I_23641 (I404346,I2507,I403922,I403908,);
not I_23642 (I404466,I2514);
DFFARX1 I_23643 (I947655,I2507,I404466,I404492,);
DFFARX1 I_23644 (I404492,I2507,I404466,I404509,);
not I_23645 (I404458,I404509);
not I_23646 (I404531,I404492);
nand I_23647 (I404548,I947670,I947658);
and I_23648 (I404565,I404548,I947649);
DFFARX1 I_23649 (I404565,I2507,I404466,I404591,);
not I_23650 (I404599,I404591);
DFFARX1 I_23651 (I947661,I2507,I404466,I404625,);
and I_23652 (I404633,I404625,I947652);
nand I_23653 (I404650,I404625,I947652);
nand I_23654 (I404437,I404599,I404650);
DFFARX1 I_23655 (I947667,I2507,I404466,I404690,);
nor I_23656 (I404698,I404690,I404633);
DFFARX1 I_23657 (I404698,I2507,I404466,I404431,);
nor I_23658 (I404446,I404690,I404591);
nand I_23659 (I404743,I947676,I947664);
and I_23660 (I404760,I404743,I947673);
DFFARX1 I_23661 (I404760,I2507,I404466,I404786,);
nor I_23662 (I404434,I404786,I404690);
not I_23663 (I404808,I404786);
nor I_23664 (I404825,I404808,I404599);
nor I_23665 (I404842,I404531,I404825);
DFFARX1 I_23666 (I404842,I2507,I404466,I404449,);
nor I_23667 (I404873,I404808,I404690);
nor I_23668 (I404890,I947649,I947664);
nor I_23669 (I404440,I404890,I404873);
not I_23670 (I404921,I404890);
nand I_23671 (I404443,I404650,I404921);
DFFARX1 I_23672 (I404890,I2507,I404466,I404455,);
DFFARX1 I_23673 (I404890,I2507,I404466,I404452,);
not I_23674 (I405010,I2514);
DFFARX1 I_23675 (I189509,I2507,I405010,I405036,);
DFFARX1 I_23676 (I405036,I2507,I405010,I405053,);
not I_23677 (I405002,I405053);
not I_23678 (I405075,I405036);
nand I_23679 (I405092,I189521,I189500);
and I_23680 (I405109,I405092,I189503);
DFFARX1 I_23681 (I405109,I2507,I405010,I405135,);
not I_23682 (I405143,I405135);
DFFARX1 I_23683 (I189512,I2507,I405010,I405169,);
and I_23684 (I405177,I405169,I189524);
nand I_23685 (I405194,I405169,I189524);
nand I_23686 (I404981,I405143,I405194);
DFFARX1 I_23687 (I189518,I2507,I405010,I405234,);
nor I_23688 (I405242,I405234,I405177);
DFFARX1 I_23689 (I405242,I2507,I405010,I404975,);
nor I_23690 (I404990,I405234,I405135);
nand I_23691 (I405287,I189506,I189503);
and I_23692 (I405304,I405287,I189515);
DFFARX1 I_23693 (I405304,I2507,I405010,I405330,);
nor I_23694 (I404978,I405330,I405234);
not I_23695 (I405352,I405330);
nor I_23696 (I405369,I405352,I405143);
nor I_23697 (I405386,I405075,I405369);
DFFARX1 I_23698 (I405386,I2507,I405010,I404993,);
nor I_23699 (I405417,I405352,I405234);
nor I_23700 (I405434,I189500,I189503);
nor I_23701 (I404984,I405434,I405417);
not I_23702 (I405465,I405434);
nand I_23703 (I404987,I405194,I405465);
DFFARX1 I_23704 (I405434,I2507,I405010,I404999,);
DFFARX1 I_23705 (I405434,I2507,I405010,I404996,);
not I_23706 (I405554,I2514);
DFFARX1 I_23707 (I97553,I2507,I405554,I405580,);
DFFARX1 I_23708 (I405580,I2507,I405554,I405597,);
not I_23709 (I405546,I405597);
not I_23710 (I405619,I405580);
nand I_23711 (I405636,I97568,I97547);
and I_23712 (I405653,I405636,I97550);
DFFARX1 I_23713 (I405653,I2507,I405554,I405679,);
not I_23714 (I405687,I405679);
DFFARX1 I_23715 (I97556,I2507,I405554,I405713,);
and I_23716 (I405721,I405713,I97550);
nand I_23717 (I405738,I405713,I97550);
nand I_23718 (I405525,I405687,I405738);
DFFARX1 I_23719 (I97565,I2507,I405554,I405778,);
nor I_23720 (I405786,I405778,I405721);
DFFARX1 I_23721 (I405786,I2507,I405554,I405519,);
nor I_23722 (I405534,I405778,I405679);
nand I_23723 (I405831,I97547,I97562);
and I_23724 (I405848,I405831,I97559);
DFFARX1 I_23725 (I405848,I2507,I405554,I405874,);
nor I_23726 (I405522,I405874,I405778);
not I_23727 (I405896,I405874);
nor I_23728 (I405913,I405896,I405687);
nor I_23729 (I405930,I405619,I405913);
DFFARX1 I_23730 (I405930,I2507,I405554,I405537,);
nor I_23731 (I405961,I405896,I405778);
nor I_23732 (I405978,I97571,I97562);
nor I_23733 (I405528,I405978,I405961);
not I_23734 (I406009,I405978);
nand I_23735 (I405531,I405738,I406009);
DFFARX1 I_23736 (I405978,I2507,I405554,I405543,);
DFFARX1 I_23737 (I405978,I2507,I405554,I405540,);
not I_23738 (I406098,I2514);
DFFARX1 I_23739 (I683897,I2507,I406098,I406124,);
DFFARX1 I_23740 (I406124,I2507,I406098,I406141,);
not I_23741 (I406090,I406141);
not I_23742 (I406163,I406124);
nand I_23743 (I406180,I683918,I683909);
and I_23744 (I406197,I406180,I683897);
DFFARX1 I_23745 (I406197,I2507,I406098,I406223,);
not I_23746 (I406231,I406223);
DFFARX1 I_23747 (I683903,I2507,I406098,I406257,);
and I_23748 (I406265,I406257,I683900);
nand I_23749 (I406282,I406257,I683900);
nand I_23750 (I406069,I406231,I406282);
DFFARX1 I_23751 (I683894,I2507,I406098,I406322,);
nor I_23752 (I406330,I406322,I406265);
DFFARX1 I_23753 (I406330,I2507,I406098,I406063,);
nor I_23754 (I406078,I406322,I406223);
nand I_23755 (I406375,I683894,I683906);
and I_23756 (I406392,I406375,I683915);
DFFARX1 I_23757 (I406392,I2507,I406098,I406418,);
nor I_23758 (I406066,I406418,I406322);
not I_23759 (I406440,I406418);
nor I_23760 (I406457,I406440,I406231);
nor I_23761 (I406474,I406163,I406457);
DFFARX1 I_23762 (I406474,I2507,I406098,I406081,);
nor I_23763 (I406505,I406440,I406322);
nor I_23764 (I406522,I683912,I683906);
nor I_23765 (I406072,I406522,I406505);
not I_23766 (I406553,I406522);
nand I_23767 (I406075,I406282,I406553);
DFFARX1 I_23768 (I406522,I2507,I406098,I406087,);
DFFARX1 I_23769 (I406522,I2507,I406098,I406084,);
not I_23770 (I406642,I2514);
DFFARX1 I_23771 (I338747,I2507,I406642,I406668,);
DFFARX1 I_23772 (I406668,I2507,I406642,I406685,);
not I_23773 (I406634,I406685);
not I_23774 (I406707,I406668);
nand I_23775 (I406724,I338726,I338750);
and I_23776 (I406741,I406724,I338753);
DFFARX1 I_23777 (I406741,I2507,I406642,I406767,);
not I_23778 (I406775,I406767);
DFFARX1 I_23779 (I338735,I2507,I406642,I406801,);
and I_23780 (I406809,I406801,I338741);
nand I_23781 (I406826,I406801,I338741);
nand I_23782 (I406613,I406775,I406826);
DFFARX1 I_23783 (I338729,I2507,I406642,I406866,);
nor I_23784 (I406874,I406866,I406809);
DFFARX1 I_23785 (I406874,I2507,I406642,I406607,);
nor I_23786 (I406622,I406866,I406767);
nand I_23787 (I406919,I338738,I338726);
and I_23788 (I406936,I406919,I338732);
DFFARX1 I_23789 (I406936,I2507,I406642,I406962,);
nor I_23790 (I406610,I406962,I406866);
not I_23791 (I406984,I406962);
nor I_23792 (I407001,I406984,I406775);
nor I_23793 (I407018,I406707,I407001);
DFFARX1 I_23794 (I407018,I2507,I406642,I406625,);
nor I_23795 (I407049,I406984,I406866);
nor I_23796 (I407066,I338744,I338726);
nor I_23797 (I406616,I407066,I407049);
not I_23798 (I407097,I407066);
nand I_23799 (I406619,I406826,I407097);
DFFARX1 I_23800 (I407066,I2507,I406642,I406631,);
DFFARX1 I_23801 (I407066,I2507,I406642,I406628,);
not I_23802 (I407186,I2514);
DFFARX1 I_23803 (I1080915,I2507,I407186,I407212,);
DFFARX1 I_23804 (I407212,I2507,I407186,I407229,);
not I_23805 (I407178,I407229);
not I_23806 (I407251,I407212);
nand I_23807 (I407268,I1080927,I1080915);
and I_23808 (I407285,I407268,I1080918);
DFFARX1 I_23809 (I407285,I2507,I407186,I407311,);
not I_23810 (I407319,I407311);
DFFARX1 I_23811 (I1080936,I2507,I407186,I407345,);
and I_23812 (I407353,I407345,I1080912);
nand I_23813 (I407370,I407345,I1080912);
nand I_23814 (I407157,I407319,I407370);
DFFARX1 I_23815 (I1080930,I2507,I407186,I407410,);
nor I_23816 (I407418,I407410,I407353);
DFFARX1 I_23817 (I407418,I2507,I407186,I407151,);
nor I_23818 (I407166,I407410,I407311);
nand I_23819 (I407463,I1080924,I1080921);
and I_23820 (I407480,I407463,I1080933);
DFFARX1 I_23821 (I407480,I2507,I407186,I407506,);
nor I_23822 (I407154,I407506,I407410);
not I_23823 (I407528,I407506);
nor I_23824 (I407545,I407528,I407319);
nor I_23825 (I407562,I407251,I407545);
DFFARX1 I_23826 (I407562,I2507,I407186,I407169,);
nor I_23827 (I407593,I407528,I407410);
nor I_23828 (I407610,I1080912,I1080921);
nor I_23829 (I407160,I407610,I407593);
not I_23830 (I407641,I407610);
nand I_23831 (I407163,I407370,I407641);
DFFARX1 I_23832 (I407610,I2507,I407186,I407175,);
DFFARX1 I_23833 (I407610,I2507,I407186,I407172,);
not I_23834 (I407730,I2514);
DFFARX1 I_23835 (I517892,I2507,I407730,I407756,);
DFFARX1 I_23836 (I407756,I2507,I407730,I407773,);
not I_23837 (I407722,I407773);
not I_23838 (I407795,I407756);
nand I_23839 (I407812,I517895,I517913);
and I_23840 (I407829,I407812,I517901);
DFFARX1 I_23841 (I407829,I2507,I407730,I407855,);
not I_23842 (I407863,I407855);
DFFARX1 I_23843 (I517892,I2507,I407730,I407889,);
and I_23844 (I407897,I407889,I517910);
nand I_23845 (I407914,I407889,I517910);
nand I_23846 (I407701,I407863,I407914);
DFFARX1 I_23847 (I517904,I2507,I407730,I407954,);
nor I_23848 (I407962,I407954,I407897);
DFFARX1 I_23849 (I407962,I2507,I407730,I407695,);
nor I_23850 (I407710,I407954,I407855);
nand I_23851 (I408007,I517907,I517889);
and I_23852 (I408024,I408007,I517898);
DFFARX1 I_23853 (I408024,I2507,I407730,I408050,);
nor I_23854 (I407698,I408050,I407954);
not I_23855 (I408072,I408050);
nor I_23856 (I408089,I408072,I407863);
nor I_23857 (I408106,I407795,I408089);
DFFARX1 I_23858 (I408106,I2507,I407730,I407713,);
nor I_23859 (I408137,I408072,I407954);
nor I_23860 (I408154,I517889,I517889);
nor I_23861 (I407704,I408154,I408137);
not I_23862 (I408185,I408154);
nand I_23863 (I407707,I407914,I408185);
DFFARX1 I_23864 (I408154,I2507,I407730,I407719,);
DFFARX1 I_23865 (I408154,I2507,I407730,I407716,);
not I_23866 (I408274,I2514);
DFFARX1 I_23867 (I1380309,I2507,I408274,I408300,);
DFFARX1 I_23868 (I408300,I2507,I408274,I408317,);
not I_23869 (I408266,I408317);
not I_23870 (I408339,I408300);
nand I_23871 (I408356,I1380285,I1380306);
and I_23872 (I408373,I408356,I1380303);
DFFARX1 I_23873 (I408373,I2507,I408274,I408399,);
not I_23874 (I408407,I408399);
DFFARX1 I_23875 (I1380282,I2507,I408274,I408433,);
and I_23876 (I408441,I408433,I1380294);
nand I_23877 (I408458,I408433,I1380294);
nand I_23878 (I408245,I408407,I408458);
DFFARX1 I_23879 (I1380297,I2507,I408274,I408498,);
nor I_23880 (I408506,I408498,I408441);
DFFARX1 I_23881 (I408506,I2507,I408274,I408239,);
nor I_23882 (I408254,I408498,I408399);
nand I_23883 (I408551,I1380300,I1380288);
and I_23884 (I408568,I408551,I1380291);
DFFARX1 I_23885 (I408568,I2507,I408274,I408594,);
nor I_23886 (I408242,I408594,I408498);
not I_23887 (I408616,I408594);
nor I_23888 (I408633,I408616,I408407);
nor I_23889 (I408650,I408339,I408633);
DFFARX1 I_23890 (I408650,I2507,I408274,I408257,);
nor I_23891 (I408681,I408616,I408498);
nor I_23892 (I408698,I1380282,I1380288);
nor I_23893 (I408248,I408698,I408681);
not I_23894 (I408729,I408698);
nand I_23895 (I408251,I408458,I408729);
DFFARX1 I_23896 (I408698,I2507,I408274,I408263,);
DFFARX1 I_23897 (I408698,I2507,I408274,I408260,);
not I_23898 (I408818,I2514);
DFFARX1 I_23899 (I149644,I2507,I408818,I408844,);
DFFARX1 I_23900 (I408844,I2507,I408818,I408861,);
not I_23901 (I408810,I408861);
not I_23902 (I408883,I408844);
nand I_23903 (I408900,I149656,I149635);
and I_23904 (I408917,I408900,I149638);
DFFARX1 I_23905 (I408917,I2507,I408818,I408943,);
not I_23906 (I408951,I408943);
DFFARX1 I_23907 (I149647,I2507,I408818,I408977,);
and I_23908 (I408985,I408977,I149659);
nand I_23909 (I409002,I408977,I149659);
nand I_23910 (I408789,I408951,I409002);
DFFARX1 I_23911 (I149653,I2507,I408818,I409042,);
nor I_23912 (I409050,I409042,I408985);
DFFARX1 I_23913 (I409050,I2507,I408818,I408783,);
nor I_23914 (I408798,I409042,I408943);
nand I_23915 (I409095,I149641,I149638);
and I_23916 (I409112,I409095,I149650);
DFFARX1 I_23917 (I409112,I2507,I408818,I409138,);
nor I_23918 (I408786,I409138,I409042);
not I_23919 (I409160,I409138);
nor I_23920 (I409177,I409160,I408951);
nor I_23921 (I409194,I408883,I409177);
DFFARX1 I_23922 (I409194,I2507,I408818,I408801,);
nor I_23923 (I409225,I409160,I409042);
nor I_23924 (I409242,I149635,I149638);
nor I_23925 (I408792,I409242,I409225);
not I_23926 (I409273,I409242);
nand I_23927 (I408795,I409002,I409273);
DFFARX1 I_23928 (I409242,I2507,I408818,I408807,);
DFFARX1 I_23929 (I409242,I2507,I408818,I408804,);
not I_23930 (I409362,I2514);
DFFARX1 I_23931 (I801206,I2507,I409362,I409388,);
DFFARX1 I_23932 (I409388,I2507,I409362,I409405,);
not I_23933 (I409354,I409405);
not I_23934 (I409427,I409388);
nand I_23935 (I409444,I801200,I801197);
and I_23936 (I409461,I409444,I801212);
DFFARX1 I_23937 (I409461,I2507,I409362,I409487,);
not I_23938 (I409495,I409487);
DFFARX1 I_23939 (I801200,I2507,I409362,I409521,);
and I_23940 (I409529,I409521,I801194);
nand I_23941 (I409546,I409521,I801194);
nand I_23942 (I409333,I409495,I409546);
DFFARX1 I_23943 (I801194,I2507,I409362,I409586,);
nor I_23944 (I409594,I409586,I409529);
DFFARX1 I_23945 (I409594,I2507,I409362,I409327,);
nor I_23946 (I409342,I409586,I409487);
nand I_23947 (I409639,I801209,I801203);
and I_23948 (I409656,I409639,I801197);
DFFARX1 I_23949 (I409656,I2507,I409362,I409682,);
nor I_23950 (I409330,I409682,I409586);
not I_23951 (I409704,I409682);
nor I_23952 (I409721,I409704,I409495);
nor I_23953 (I409738,I409427,I409721);
DFFARX1 I_23954 (I409738,I2507,I409362,I409345,);
nor I_23955 (I409769,I409704,I409586);
nor I_23956 (I409786,I801215,I801203);
nor I_23957 (I409336,I409786,I409769);
not I_23958 (I409817,I409786);
nand I_23959 (I409339,I409546,I409817);
DFFARX1 I_23960 (I409786,I2507,I409362,I409351,);
DFFARX1 I_23961 (I409786,I2507,I409362,I409348,);
not I_23962 (I409906,I2514);
DFFARX1 I_23963 (I138342,I2507,I409906,I409932,);
DFFARX1 I_23964 (I409932,I2507,I409906,I409949,);
not I_23965 (I409898,I409949);
not I_23966 (I409971,I409932);
nand I_23967 (I409988,I138351,I138354);
and I_23968 (I410005,I409988,I138333);
DFFARX1 I_23969 (I410005,I2507,I409906,I410031,);
not I_23970 (I410039,I410031);
DFFARX1 I_23971 (I138348,I2507,I409906,I410065,);
and I_23972 (I410073,I410065,I138336);
nand I_23973 (I410090,I410065,I138336);
nand I_23974 (I409877,I410039,I410090);
DFFARX1 I_23975 (I138330,I2507,I409906,I410130,);
nor I_23976 (I410138,I410130,I410073);
DFFARX1 I_23977 (I410138,I2507,I409906,I409871,);
nor I_23978 (I409886,I410130,I410031);
nand I_23979 (I410183,I138345,I138339);
and I_23980 (I410200,I410183,I138330);
DFFARX1 I_23981 (I410200,I2507,I409906,I410226,);
nor I_23982 (I409874,I410226,I410130);
not I_23983 (I410248,I410226);
nor I_23984 (I410265,I410248,I410039);
nor I_23985 (I410282,I409971,I410265);
DFFARX1 I_23986 (I410282,I2507,I409906,I409889,);
nor I_23987 (I410313,I410248,I410130);
nor I_23988 (I410330,I138357,I138339);
nor I_23989 (I409880,I410330,I410313);
not I_23990 (I410361,I410330);
nand I_23991 (I409883,I410090,I410361);
DFFARX1 I_23992 (I410330,I2507,I409906,I409895,);
DFFARX1 I_23993 (I410330,I2507,I409906,I409892,);
not I_23994 (I410450,I2514);
DFFARX1 I_23995 (I1234629,I2507,I410450,I410476,);
DFFARX1 I_23996 (I410476,I2507,I410450,I410493,);
not I_23997 (I410442,I410493);
not I_23998 (I410515,I410476);
nand I_23999 (I410532,I1234641,I1234644);
and I_24000 (I410549,I410532,I1234647);
DFFARX1 I_24001 (I410549,I2507,I410450,I410575,);
not I_24002 (I410583,I410575);
DFFARX1 I_24003 (I1234632,I2507,I410450,I410609,);
and I_24004 (I410617,I410609,I1234638);
nand I_24005 (I410634,I410609,I1234638);
nand I_24006 (I410421,I410583,I410634);
DFFARX1 I_24007 (I1234626,I2507,I410450,I410674,);
nor I_24008 (I410682,I410674,I410617);
DFFARX1 I_24009 (I410682,I2507,I410450,I410415,);
nor I_24010 (I410430,I410674,I410575);
nand I_24011 (I410727,I1234629,I1234650);
and I_24012 (I410744,I410727,I1234635);
DFFARX1 I_24013 (I410744,I2507,I410450,I410770,);
nor I_24014 (I410418,I410770,I410674);
not I_24015 (I410792,I410770);
nor I_24016 (I410809,I410792,I410583);
nor I_24017 (I410826,I410515,I410809);
DFFARX1 I_24018 (I410826,I2507,I410450,I410433,);
nor I_24019 (I410857,I410792,I410674);
nor I_24020 (I410874,I1234626,I1234650);
nor I_24021 (I410424,I410874,I410857);
not I_24022 (I410905,I410874);
nand I_24023 (I410427,I410634,I410905);
DFFARX1 I_24024 (I410874,I2507,I410450,I410439,);
DFFARX1 I_24025 (I410874,I2507,I410450,I410436,);
not I_24026 (I410994,I2514);
DFFARX1 I_24027 (I1143917,I2507,I410994,I411020,);
DFFARX1 I_24028 (I411020,I2507,I410994,I411037,);
not I_24029 (I410986,I411037);
not I_24030 (I411059,I411020);
nand I_24031 (I411076,I1143929,I1143917);
and I_24032 (I411093,I411076,I1143920);
DFFARX1 I_24033 (I411093,I2507,I410994,I411119,);
not I_24034 (I411127,I411119);
DFFARX1 I_24035 (I1143938,I2507,I410994,I411153,);
and I_24036 (I411161,I411153,I1143914);
nand I_24037 (I411178,I411153,I1143914);
nand I_24038 (I410965,I411127,I411178);
DFFARX1 I_24039 (I1143932,I2507,I410994,I411218,);
nor I_24040 (I411226,I411218,I411161);
DFFARX1 I_24041 (I411226,I2507,I410994,I410959,);
nor I_24042 (I410974,I411218,I411119);
nand I_24043 (I411271,I1143926,I1143923);
and I_24044 (I411288,I411271,I1143935);
DFFARX1 I_24045 (I411288,I2507,I410994,I411314,);
nor I_24046 (I410962,I411314,I411218);
not I_24047 (I411336,I411314);
nor I_24048 (I411353,I411336,I411127);
nor I_24049 (I411370,I411059,I411353);
DFFARX1 I_24050 (I411370,I2507,I410994,I410977,);
nor I_24051 (I411401,I411336,I411218);
nor I_24052 (I411418,I1143914,I1143923);
nor I_24053 (I410968,I411418,I411401);
not I_24054 (I411449,I411418);
nand I_24055 (I410971,I411178,I411449);
DFFARX1 I_24056 (I411418,I2507,I410994,I410983,);
DFFARX1 I_24057 (I411418,I2507,I410994,I410980,);
not I_24058 (I411538,I2514);
DFFARX1 I_24059 (I1101145,I2507,I411538,I411564,);
DFFARX1 I_24060 (I411564,I2507,I411538,I411581,);
not I_24061 (I411530,I411581);
not I_24062 (I411603,I411564);
nand I_24063 (I411620,I1101157,I1101145);
and I_24064 (I411637,I411620,I1101148);
DFFARX1 I_24065 (I411637,I2507,I411538,I411663,);
not I_24066 (I411671,I411663);
DFFARX1 I_24067 (I1101166,I2507,I411538,I411697,);
and I_24068 (I411705,I411697,I1101142);
nand I_24069 (I411722,I411697,I1101142);
nand I_24070 (I411509,I411671,I411722);
DFFARX1 I_24071 (I1101160,I2507,I411538,I411762,);
nor I_24072 (I411770,I411762,I411705);
DFFARX1 I_24073 (I411770,I2507,I411538,I411503,);
nor I_24074 (I411518,I411762,I411663);
nand I_24075 (I411815,I1101154,I1101151);
and I_24076 (I411832,I411815,I1101163);
DFFARX1 I_24077 (I411832,I2507,I411538,I411858,);
nor I_24078 (I411506,I411858,I411762);
not I_24079 (I411880,I411858);
nor I_24080 (I411897,I411880,I411671);
nor I_24081 (I411914,I411603,I411897);
DFFARX1 I_24082 (I411914,I2507,I411538,I411521,);
nor I_24083 (I411945,I411880,I411762);
nor I_24084 (I411962,I1101142,I1101151);
nor I_24085 (I411512,I411962,I411945);
not I_24086 (I411993,I411962);
nand I_24087 (I411515,I411722,I411993);
DFFARX1 I_24088 (I411962,I2507,I411538,I411527,);
DFFARX1 I_24089 (I411962,I2507,I411538,I411524,);
not I_24090 (I412082,I2514);
DFFARX1 I_24091 (I360354,I2507,I412082,I412108,);
DFFARX1 I_24092 (I412108,I2507,I412082,I412125,);
not I_24093 (I412074,I412125);
not I_24094 (I412147,I412108);
nand I_24095 (I412164,I360333,I360357);
and I_24096 (I412181,I412164,I360360);
DFFARX1 I_24097 (I412181,I2507,I412082,I412207,);
not I_24098 (I412215,I412207);
DFFARX1 I_24099 (I360342,I2507,I412082,I412241,);
and I_24100 (I412249,I412241,I360348);
nand I_24101 (I412266,I412241,I360348);
nand I_24102 (I412053,I412215,I412266);
DFFARX1 I_24103 (I360336,I2507,I412082,I412306,);
nor I_24104 (I412314,I412306,I412249);
DFFARX1 I_24105 (I412314,I2507,I412082,I412047,);
nor I_24106 (I412062,I412306,I412207);
nand I_24107 (I412359,I360345,I360333);
and I_24108 (I412376,I412359,I360339);
DFFARX1 I_24109 (I412376,I2507,I412082,I412402,);
nor I_24110 (I412050,I412402,I412306);
not I_24111 (I412424,I412402);
nor I_24112 (I412441,I412424,I412215);
nor I_24113 (I412458,I412147,I412441);
DFFARX1 I_24114 (I412458,I2507,I412082,I412065,);
nor I_24115 (I412489,I412424,I412306);
nor I_24116 (I412506,I360351,I360333);
nor I_24117 (I412056,I412506,I412489);
not I_24118 (I412537,I412506);
nand I_24119 (I412059,I412266,I412537);
DFFARX1 I_24120 (I412506,I2507,I412082,I412071,);
DFFARX1 I_24121 (I412506,I2507,I412082,I412068,);
not I_24122 (I412626,I2514);
DFFARX1 I_24123 (I150834,I2507,I412626,I412652,);
DFFARX1 I_24124 (I412652,I2507,I412626,I412669,);
not I_24125 (I412618,I412669);
not I_24126 (I412691,I412652);
nand I_24127 (I412708,I150846,I150825);
and I_24128 (I412725,I412708,I150828);
DFFARX1 I_24129 (I412725,I2507,I412626,I412751,);
not I_24130 (I412759,I412751);
DFFARX1 I_24131 (I150837,I2507,I412626,I412785,);
and I_24132 (I412793,I412785,I150849);
nand I_24133 (I412810,I412785,I150849);
nand I_24134 (I412597,I412759,I412810);
DFFARX1 I_24135 (I150843,I2507,I412626,I412850,);
nor I_24136 (I412858,I412850,I412793);
DFFARX1 I_24137 (I412858,I2507,I412626,I412591,);
nor I_24138 (I412606,I412850,I412751);
nand I_24139 (I412903,I150831,I150828);
and I_24140 (I412920,I412903,I150840);
DFFARX1 I_24141 (I412920,I2507,I412626,I412946,);
nor I_24142 (I412594,I412946,I412850);
not I_24143 (I412968,I412946);
nor I_24144 (I412985,I412968,I412759);
nor I_24145 (I413002,I412691,I412985);
DFFARX1 I_24146 (I413002,I2507,I412626,I412609,);
nor I_24147 (I413033,I412968,I412850);
nor I_24148 (I413050,I150825,I150828);
nor I_24149 (I412600,I413050,I413033);
not I_24150 (I413081,I413050);
nand I_24151 (I412603,I412810,I413081);
DFFARX1 I_24152 (I413050,I2507,I412626,I412615,);
DFFARX1 I_24153 (I413050,I2507,I412626,I412612,);
not I_24154 (I413170,I2514);
DFFARX1 I_24155 (I1255350,I2507,I413170,I413196,);
DFFARX1 I_24156 (I413196,I2507,I413170,I413213,);
not I_24157 (I413162,I413213);
not I_24158 (I413235,I413196);
nand I_24159 (I413252,I1255347,I1255344);
and I_24160 (I413269,I413252,I1255332);
DFFARX1 I_24161 (I413269,I2507,I413170,I413295,);
not I_24162 (I413303,I413295);
DFFARX1 I_24163 (I1255356,I2507,I413170,I413329,);
and I_24164 (I413337,I413329,I1255341);
nand I_24165 (I413354,I413329,I1255341);
nand I_24166 (I413141,I413303,I413354);
DFFARX1 I_24167 (I1255335,I2507,I413170,I413394,);
nor I_24168 (I413402,I413394,I413337);
DFFARX1 I_24169 (I413402,I2507,I413170,I413135,);
nor I_24170 (I413150,I413394,I413295);
nand I_24171 (I413447,I1255332,I1255338);
and I_24172 (I413464,I413447,I1255353);
DFFARX1 I_24173 (I413464,I2507,I413170,I413490,);
nor I_24174 (I413138,I413490,I413394);
not I_24175 (I413512,I413490);
nor I_24176 (I413529,I413512,I413303);
nor I_24177 (I413546,I413235,I413529);
DFFARX1 I_24178 (I413546,I2507,I413170,I413153,);
nor I_24179 (I413577,I413512,I413394);
nor I_24180 (I413594,I1255335,I1255338);
nor I_24181 (I413144,I413594,I413577);
not I_24182 (I413625,I413594);
nand I_24183 (I413147,I413354,I413625);
DFFARX1 I_24184 (I413594,I2507,I413170,I413159,);
DFFARX1 I_24185 (I413594,I2507,I413170,I413156,);
not I_24186 (I413714,I2514);
DFFARX1 I_24187 (I1373764,I2507,I413714,I413740,);
DFFARX1 I_24188 (I413740,I2507,I413714,I413757,);
not I_24189 (I413706,I413757);
not I_24190 (I413779,I413740);
nand I_24191 (I413796,I1373740,I1373761);
and I_24192 (I413813,I413796,I1373758);
DFFARX1 I_24193 (I413813,I2507,I413714,I413839,);
not I_24194 (I413847,I413839);
DFFARX1 I_24195 (I1373737,I2507,I413714,I413873,);
and I_24196 (I413881,I413873,I1373749);
nand I_24197 (I413898,I413873,I1373749);
nand I_24198 (I413685,I413847,I413898);
DFFARX1 I_24199 (I1373752,I2507,I413714,I413938,);
nor I_24200 (I413946,I413938,I413881);
DFFARX1 I_24201 (I413946,I2507,I413714,I413679,);
nor I_24202 (I413694,I413938,I413839);
nand I_24203 (I413991,I1373755,I1373743);
and I_24204 (I414008,I413991,I1373746);
DFFARX1 I_24205 (I414008,I2507,I413714,I414034,);
nor I_24206 (I413682,I414034,I413938);
not I_24207 (I414056,I414034);
nor I_24208 (I414073,I414056,I413847);
nor I_24209 (I414090,I413779,I414073);
DFFARX1 I_24210 (I414090,I2507,I413714,I413697,);
nor I_24211 (I414121,I414056,I413938);
nor I_24212 (I414138,I1373737,I1373743);
nor I_24213 (I413688,I414138,I414121);
not I_24214 (I414169,I414138);
nand I_24215 (I413691,I413898,I414169);
DFFARX1 I_24216 (I414138,I2507,I413714,I413703,);
DFFARX1 I_24217 (I414138,I2507,I413714,I413700,);
not I_24218 (I414258,I2514);
DFFARX1 I_24219 (I364570,I2507,I414258,I414284,);
DFFARX1 I_24220 (I414284,I2507,I414258,I414301,);
not I_24221 (I414250,I414301);
not I_24222 (I414323,I414284);
nand I_24223 (I414340,I364549,I364573);
and I_24224 (I414357,I414340,I364576);
DFFARX1 I_24225 (I414357,I2507,I414258,I414383,);
not I_24226 (I414391,I414383);
DFFARX1 I_24227 (I364558,I2507,I414258,I414417,);
and I_24228 (I414425,I414417,I364564);
nand I_24229 (I414442,I414417,I364564);
nand I_24230 (I414229,I414391,I414442);
DFFARX1 I_24231 (I364552,I2507,I414258,I414482,);
nor I_24232 (I414490,I414482,I414425);
DFFARX1 I_24233 (I414490,I2507,I414258,I414223,);
nor I_24234 (I414238,I414482,I414383);
nand I_24235 (I414535,I364561,I364549);
and I_24236 (I414552,I414535,I364555);
DFFARX1 I_24237 (I414552,I2507,I414258,I414578,);
nor I_24238 (I414226,I414578,I414482);
not I_24239 (I414600,I414578);
nor I_24240 (I414617,I414600,I414391);
nor I_24241 (I414634,I414323,I414617);
DFFARX1 I_24242 (I414634,I2507,I414258,I414241,);
nor I_24243 (I414665,I414600,I414482);
nor I_24244 (I414682,I364567,I364549);
nor I_24245 (I414232,I414682,I414665);
not I_24246 (I414713,I414682);
nand I_24247 (I414235,I414442,I414713);
DFFARX1 I_24248 (I414682,I2507,I414258,I414247,);
DFFARX1 I_24249 (I414682,I2507,I414258,I414244,);
not I_24250 (I414802,I2514);
DFFARX1 I_24251 (I1106347,I2507,I414802,I414828,);
DFFARX1 I_24252 (I414828,I2507,I414802,I414845,);
not I_24253 (I414794,I414845);
not I_24254 (I414867,I414828);
nand I_24255 (I414884,I1106359,I1106347);
and I_24256 (I414901,I414884,I1106350);
DFFARX1 I_24257 (I414901,I2507,I414802,I414927,);
not I_24258 (I414935,I414927);
DFFARX1 I_24259 (I1106368,I2507,I414802,I414961,);
and I_24260 (I414969,I414961,I1106344);
nand I_24261 (I414986,I414961,I1106344);
nand I_24262 (I414773,I414935,I414986);
DFFARX1 I_24263 (I1106362,I2507,I414802,I415026,);
nor I_24264 (I415034,I415026,I414969);
DFFARX1 I_24265 (I415034,I2507,I414802,I414767,);
nor I_24266 (I414782,I415026,I414927);
nand I_24267 (I415079,I1106356,I1106353);
and I_24268 (I415096,I415079,I1106365);
DFFARX1 I_24269 (I415096,I2507,I414802,I415122,);
nor I_24270 (I414770,I415122,I415026);
not I_24271 (I415144,I415122);
nor I_24272 (I415161,I415144,I414935);
nor I_24273 (I415178,I414867,I415161);
DFFARX1 I_24274 (I415178,I2507,I414802,I414785,);
nor I_24275 (I415209,I415144,I415026);
nor I_24276 (I415226,I1106344,I1106353);
nor I_24277 (I414776,I415226,I415209);
not I_24278 (I415257,I415226);
nand I_24279 (I414779,I414986,I415257);
DFFARX1 I_24280 (I415226,I2507,I414802,I414791,);
DFFARX1 I_24281 (I415226,I2507,I414802,I414788,);
not I_24282 (I415346,I2514);
DFFARX1 I_24283 (I1237893,I2507,I415346,I415372,);
DFFARX1 I_24284 (I415372,I2507,I415346,I415389,);
not I_24285 (I415338,I415389);
not I_24286 (I415411,I415372);
nand I_24287 (I415428,I1237905,I1237908);
and I_24288 (I415445,I415428,I1237911);
DFFARX1 I_24289 (I415445,I2507,I415346,I415471,);
not I_24290 (I415479,I415471);
DFFARX1 I_24291 (I1237896,I2507,I415346,I415505,);
and I_24292 (I415513,I415505,I1237902);
nand I_24293 (I415530,I415505,I1237902);
nand I_24294 (I415317,I415479,I415530);
DFFARX1 I_24295 (I1237890,I2507,I415346,I415570,);
nor I_24296 (I415578,I415570,I415513);
DFFARX1 I_24297 (I415578,I2507,I415346,I415311,);
nor I_24298 (I415326,I415570,I415471);
nand I_24299 (I415623,I1237893,I1237914);
and I_24300 (I415640,I415623,I1237899);
DFFARX1 I_24301 (I415640,I2507,I415346,I415666,);
nor I_24302 (I415314,I415666,I415570);
not I_24303 (I415688,I415666);
nor I_24304 (I415705,I415688,I415479);
nor I_24305 (I415722,I415411,I415705);
DFFARX1 I_24306 (I415722,I2507,I415346,I415329,);
nor I_24307 (I415753,I415688,I415570);
nor I_24308 (I415770,I1237890,I1237914);
nor I_24309 (I415320,I415770,I415753);
not I_24310 (I415801,I415770);
nand I_24311 (I415323,I415530,I415801);
DFFARX1 I_24312 (I415770,I2507,I415346,I415335,);
DFFARX1 I_24313 (I415770,I2507,I415346,I415332,);
not I_24314 (I415890,I2514);
DFFARX1 I_24315 (I860757,I2507,I415890,I415916,);
DFFARX1 I_24316 (I415916,I2507,I415890,I415933,);
not I_24317 (I415882,I415933);
not I_24318 (I415955,I415916);
nand I_24319 (I415972,I860751,I860748);
and I_24320 (I415989,I415972,I860763);
DFFARX1 I_24321 (I415989,I2507,I415890,I416015,);
not I_24322 (I416023,I416015);
DFFARX1 I_24323 (I860751,I2507,I415890,I416049,);
and I_24324 (I416057,I416049,I860745);
nand I_24325 (I416074,I416049,I860745);
nand I_24326 (I415861,I416023,I416074);
DFFARX1 I_24327 (I860745,I2507,I415890,I416114,);
nor I_24328 (I416122,I416114,I416057);
DFFARX1 I_24329 (I416122,I2507,I415890,I415855,);
nor I_24330 (I415870,I416114,I416015);
nand I_24331 (I416167,I860760,I860754);
and I_24332 (I416184,I416167,I860748);
DFFARX1 I_24333 (I416184,I2507,I415890,I416210,);
nor I_24334 (I415858,I416210,I416114);
not I_24335 (I416232,I416210);
nor I_24336 (I416249,I416232,I416023);
nor I_24337 (I416266,I415955,I416249);
DFFARX1 I_24338 (I416266,I2507,I415890,I415873,);
nor I_24339 (I416297,I416232,I416114);
nor I_24340 (I416314,I860766,I860754);
nor I_24341 (I415864,I416314,I416297);
not I_24342 (I416345,I416314);
nand I_24343 (I415867,I416074,I416345);
DFFARX1 I_24344 (I416314,I2507,I415890,I415879,);
DFFARX1 I_24345 (I416314,I2507,I415890,I415876,);
not I_24346 (I416434,I2514);
DFFARX1 I_24347 (I685631,I2507,I416434,I416460,);
DFFARX1 I_24348 (I416460,I2507,I416434,I416477,);
not I_24349 (I416426,I416477);
not I_24350 (I416499,I416460);
nand I_24351 (I416516,I685652,I685643);
and I_24352 (I416533,I416516,I685631);
DFFARX1 I_24353 (I416533,I2507,I416434,I416559,);
not I_24354 (I416567,I416559);
DFFARX1 I_24355 (I685637,I2507,I416434,I416593,);
and I_24356 (I416601,I416593,I685634);
nand I_24357 (I416618,I416593,I685634);
nand I_24358 (I416405,I416567,I416618);
DFFARX1 I_24359 (I685628,I2507,I416434,I416658,);
nor I_24360 (I416666,I416658,I416601);
DFFARX1 I_24361 (I416666,I2507,I416434,I416399,);
nor I_24362 (I416414,I416658,I416559);
nand I_24363 (I416711,I685628,I685640);
and I_24364 (I416728,I416711,I685649);
DFFARX1 I_24365 (I416728,I2507,I416434,I416754,);
nor I_24366 (I416402,I416754,I416658);
not I_24367 (I416776,I416754);
nor I_24368 (I416793,I416776,I416567);
nor I_24369 (I416810,I416499,I416793);
DFFARX1 I_24370 (I416810,I2507,I416434,I416417,);
nor I_24371 (I416841,I416776,I416658);
nor I_24372 (I416858,I685646,I685640);
nor I_24373 (I416408,I416858,I416841);
not I_24374 (I416889,I416858);
nand I_24375 (I416411,I416618,I416889);
DFFARX1 I_24376 (I416858,I2507,I416434,I416423,);
DFFARX1 I_24377 (I416858,I2507,I416434,I416420,);
not I_24378 (I416978,I2514);
DFFARX1 I_24379 (I1374954,I2507,I416978,I417004,);
DFFARX1 I_24380 (I417004,I2507,I416978,I417021,);
not I_24381 (I416970,I417021);
not I_24382 (I417043,I417004);
nand I_24383 (I417060,I1374930,I1374951);
and I_24384 (I417077,I417060,I1374948);
DFFARX1 I_24385 (I417077,I2507,I416978,I417103,);
not I_24386 (I417111,I417103);
DFFARX1 I_24387 (I1374927,I2507,I416978,I417137,);
and I_24388 (I417145,I417137,I1374939);
nand I_24389 (I417162,I417137,I1374939);
nand I_24390 (I416949,I417111,I417162);
DFFARX1 I_24391 (I1374942,I2507,I416978,I417202,);
nor I_24392 (I417210,I417202,I417145);
DFFARX1 I_24393 (I417210,I2507,I416978,I416943,);
nor I_24394 (I416958,I417202,I417103);
nand I_24395 (I417255,I1374945,I1374933);
and I_24396 (I417272,I417255,I1374936);
DFFARX1 I_24397 (I417272,I2507,I416978,I417298,);
nor I_24398 (I416946,I417298,I417202);
not I_24399 (I417320,I417298);
nor I_24400 (I417337,I417320,I417111);
nor I_24401 (I417354,I417043,I417337);
DFFARX1 I_24402 (I417354,I2507,I416978,I416961,);
nor I_24403 (I417385,I417320,I417202);
nor I_24404 (I417402,I1374927,I1374933);
nor I_24405 (I416952,I417402,I417385);
not I_24406 (I417433,I417402);
nand I_24407 (I416955,I417162,I417433);
DFFARX1 I_24408 (I417402,I2507,I416978,I416967,);
DFFARX1 I_24409 (I417402,I2507,I416978,I416964,);
not I_24410 (I417522,I2514);
DFFARX1 I_24411 (I736495,I2507,I417522,I417548,);
DFFARX1 I_24412 (I417548,I2507,I417522,I417565,);
not I_24413 (I417514,I417565);
not I_24414 (I417587,I417548);
nand I_24415 (I417604,I736516,I736507);
and I_24416 (I417621,I417604,I736495);
DFFARX1 I_24417 (I417621,I2507,I417522,I417647,);
not I_24418 (I417655,I417647);
DFFARX1 I_24419 (I736501,I2507,I417522,I417681,);
and I_24420 (I417689,I417681,I736498);
nand I_24421 (I417706,I417681,I736498);
nand I_24422 (I417493,I417655,I417706);
DFFARX1 I_24423 (I736492,I2507,I417522,I417746,);
nor I_24424 (I417754,I417746,I417689);
DFFARX1 I_24425 (I417754,I2507,I417522,I417487,);
nor I_24426 (I417502,I417746,I417647);
nand I_24427 (I417799,I736492,I736504);
and I_24428 (I417816,I417799,I736513);
DFFARX1 I_24429 (I417816,I2507,I417522,I417842,);
nor I_24430 (I417490,I417842,I417746);
not I_24431 (I417864,I417842);
nor I_24432 (I417881,I417864,I417655);
nor I_24433 (I417898,I417587,I417881);
DFFARX1 I_24434 (I417898,I2507,I417522,I417505,);
nor I_24435 (I417929,I417864,I417746);
nor I_24436 (I417946,I736510,I736504);
nor I_24437 (I417496,I417946,I417929);
not I_24438 (I417977,I417946);
nand I_24439 (I417499,I417706,I417977);
DFFARX1 I_24440 (I417946,I2507,I417522,I417511,);
DFFARX1 I_24441 (I417946,I2507,I417522,I417508,);
not I_24442 (I418066,I2514);
DFFARX1 I_24443 (I815962,I2507,I418066,I418092,);
DFFARX1 I_24444 (I418092,I2507,I418066,I418109,);
not I_24445 (I418058,I418109);
not I_24446 (I418131,I418092);
nand I_24447 (I418148,I815956,I815953);
and I_24448 (I418165,I418148,I815968);
DFFARX1 I_24449 (I418165,I2507,I418066,I418191,);
not I_24450 (I418199,I418191);
DFFARX1 I_24451 (I815956,I2507,I418066,I418225,);
and I_24452 (I418233,I418225,I815950);
nand I_24453 (I418250,I418225,I815950);
nand I_24454 (I418037,I418199,I418250);
DFFARX1 I_24455 (I815950,I2507,I418066,I418290,);
nor I_24456 (I418298,I418290,I418233);
DFFARX1 I_24457 (I418298,I2507,I418066,I418031,);
nor I_24458 (I418046,I418290,I418191);
nand I_24459 (I418343,I815965,I815959);
and I_24460 (I418360,I418343,I815953);
DFFARX1 I_24461 (I418360,I2507,I418066,I418386,);
nor I_24462 (I418034,I418386,I418290);
not I_24463 (I418408,I418386);
nor I_24464 (I418425,I418408,I418199);
nor I_24465 (I418442,I418131,I418425);
DFFARX1 I_24466 (I418442,I2507,I418066,I418049,);
nor I_24467 (I418473,I418408,I418290);
nor I_24468 (I418490,I815971,I815959);
nor I_24469 (I418040,I418490,I418473);
not I_24470 (I418521,I418490);
nand I_24471 (I418043,I418250,I418521);
DFFARX1 I_24472 (I418490,I2507,I418066,I418055,);
DFFARX1 I_24473 (I418490,I2507,I418066,I418052,);
not I_24474 (I418610,I2514);
DFFARX1 I_24475 (I81216,I2507,I418610,I418636,);
DFFARX1 I_24476 (I418636,I2507,I418610,I418653,);
not I_24477 (I418602,I418653);
not I_24478 (I418675,I418636);
nand I_24479 (I418692,I81231,I81210);
and I_24480 (I418709,I418692,I81213);
DFFARX1 I_24481 (I418709,I2507,I418610,I418735,);
not I_24482 (I418743,I418735);
DFFARX1 I_24483 (I81219,I2507,I418610,I418769,);
and I_24484 (I418777,I418769,I81213);
nand I_24485 (I418794,I418769,I81213);
nand I_24486 (I418581,I418743,I418794);
DFFARX1 I_24487 (I81228,I2507,I418610,I418834,);
nor I_24488 (I418842,I418834,I418777);
DFFARX1 I_24489 (I418842,I2507,I418610,I418575,);
nor I_24490 (I418590,I418834,I418735);
nand I_24491 (I418887,I81210,I81225);
and I_24492 (I418904,I418887,I81222);
DFFARX1 I_24493 (I418904,I2507,I418610,I418930,);
nor I_24494 (I418578,I418930,I418834);
not I_24495 (I418952,I418930);
nor I_24496 (I418969,I418952,I418743);
nor I_24497 (I418986,I418675,I418969);
DFFARX1 I_24498 (I418986,I2507,I418610,I418593,);
nor I_24499 (I419017,I418952,I418834);
nor I_24500 (I419034,I81234,I81225);
nor I_24501 (I418584,I419034,I419017);
not I_24502 (I419065,I419034);
nand I_24503 (I418587,I418794,I419065);
DFFARX1 I_24504 (I419034,I2507,I418610,I418599,);
DFFARX1 I_24505 (I419034,I2507,I418610,I418596,);
not I_24506 (I419154,I2514);
DFFARX1 I_24507 (I1023605,I2507,I419154,I419180,);
DFFARX1 I_24508 (I419180,I2507,I419154,I419197,);
not I_24509 (I419146,I419197);
not I_24510 (I419219,I419180);
nand I_24511 (I419236,I1023605,I1023623);
and I_24512 (I419253,I419236,I1023617);
DFFARX1 I_24513 (I419253,I2507,I419154,I419279,);
not I_24514 (I419287,I419279);
DFFARX1 I_24515 (I1023611,I2507,I419154,I419313,);
and I_24516 (I419321,I419313,I1023620);
nand I_24517 (I419338,I419313,I1023620);
nand I_24518 (I419125,I419287,I419338);
DFFARX1 I_24519 (I1023608,I2507,I419154,I419378,);
nor I_24520 (I419386,I419378,I419321);
DFFARX1 I_24521 (I419386,I2507,I419154,I419119,);
nor I_24522 (I419134,I419378,I419279);
nand I_24523 (I419431,I1023608,I1023626);
and I_24524 (I419448,I419431,I1023611);
DFFARX1 I_24525 (I419448,I2507,I419154,I419474,);
nor I_24526 (I419122,I419474,I419378);
not I_24527 (I419496,I419474);
nor I_24528 (I419513,I419496,I419287);
nor I_24529 (I419530,I419219,I419513);
DFFARX1 I_24530 (I419530,I2507,I419154,I419137,);
nor I_24531 (I419561,I419496,I419378);
nor I_24532 (I419578,I1023614,I1023626);
nor I_24533 (I419128,I419578,I419561);
not I_24534 (I419609,I419578);
nand I_24535 (I419131,I419338,I419609);
DFFARX1 I_24536 (I419578,I2507,I419154,I419143,);
DFFARX1 I_24537 (I419578,I2507,I419154,I419140,);
not I_24538 (I419698,I2514);
DFFARX1 I_24539 (I597197,I2507,I419698,I419724,);
DFFARX1 I_24540 (I419724,I2507,I419698,I419741,);
not I_24541 (I419690,I419741);
not I_24542 (I419763,I419724);
nand I_24543 (I419780,I597194,I597215);
and I_24544 (I419797,I419780,I597218);
DFFARX1 I_24545 (I419797,I2507,I419698,I419823,);
not I_24546 (I419831,I419823);
DFFARX1 I_24547 (I597203,I2507,I419698,I419857,);
and I_24548 (I419865,I419857,I597206);
nand I_24549 (I419882,I419857,I597206);
nand I_24550 (I419669,I419831,I419882);
DFFARX1 I_24551 (I597209,I2507,I419698,I419922,);
nor I_24552 (I419930,I419922,I419865);
DFFARX1 I_24553 (I419930,I2507,I419698,I419663,);
nor I_24554 (I419678,I419922,I419823);
nand I_24555 (I419975,I597194,I597200);
and I_24556 (I419992,I419975,I597212);
DFFARX1 I_24557 (I419992,I2507,I419698,I420018,);
nor I_24558 (I419666,I420018,I419922);
not I_24559 (I420040,I420018);
nor I_24560 (I420057,I420040,I419831);
nor I_24561 (I420074,I419763,I420057);
DFFARX1 I_24562 (I420074,I2507,I419698,I419681,);
nor I_24563 (I420105,I420040,I419922);
nor I_24564 (I420122,I597197,I597200);
nor I_24565 (I419672,I420122,I420105);
not I_24566 (I420153,I420122);
nand I_24567 (I419675,I419882,I420153);
DFFARX1 I_24568 (I420122,I2507,I419698,I419687,);
DFFARX1 I_24569 (I420122,I2507,I419698,I419684,);
not I_24570 (I420242,I2514);
DFFARX1 I_24571 (I1154321,I2507,I420242,I420268,);
DFFARX1 I_24572 (I420268,I2507,I420242,I420285,);
not I_24573 (I420234,I420285);
not I_24574 (I420307,I420268);
nand I_24575 (I420324,I1154333,I1154321);
and I_24576 (I420341,I420324,I1154324);
DFFARX1 I_24577 (I420341,I2507,I420242,I420367,);
not I_24578 (I420375,I420367);
DFFARX1 I_24579 (I1154342,I2507,I420242,I420401,);
and I_24580 (I420409,I420401,I1154318);
nand I_24581 (I420426,I420401,I1154318);
nand I_24582 (I420213,I420375,I420426);
DFFARX1 I_24583 (I1154336,I2507,I420242,I420466,);
nor I_24584 (I420474,I420466,I420409);
DFFARX1 I_24585 (I420474,I2507,I420242,I420207,);
nor I_24586 (I420222,I420466,I420367);
nand I_24587 (I420519,I1154330,I1154327);
and I_24588 (I420536,I420519,I1154339);
DFFARX1 I_24589 (I420536,I2507,I420242,I420562,);
nor I_24590 (I420210,I420562,I420466);
not I_24591 (I420584,I420562);
nor I_24592 (I420601,I420584,I420375);
nor I_24593 (I420618,I420307,I420601);
DFFARX1 I_24594 (I420618,I2507,I420242,I420225,);
nor I_24595 (I420649,I420584,I420466);
nor I_24596 (I420666,I1154318,I1154327);
nor I_24597 (I420216,I420666,I420649);
not I_24598 (I420697,I420666);
nand I_24599 (I420219,I420426,I420697);
DFFARX1 I_24600 (I420666,I2507,I420242,I420231,);
DFFARX1 I_24601 (I420666,I2507,I420242,I420228,);
not I_24602 (I420786,I2514);
DFFARX1 I_24603 (I119687,I2507,I420786,I420812,);
DFFARX1 I_24604 (I420812,I2507,I420786,I420829,);
not I_24605 (I420778,I420829);
not I_24606 (I420851,I420812);
nand I_24607 (I420868,I119702,I119681);
and I_24608 (I420885,I420868,I119684);
DFFARX1 I_24609 (I420885,I2507,I420786,I420911,);
not I_24610 (I420919,I420911);
DFFARX1 I_24611 (I119690,I2507,I420786,I420945,);
and I_24612 (I420953,I420945,I119684);
nand I_24613 (I420970,I420945,I119684);
nand I_24614 (I420757,I420919,I420970);
DFFARX1 I_24615 (I119699,I2507,I420786,I421010,);
nor I_24616 (I421018,I421010,I420953);
DFFARX1 I_24617 (I421018,I2507,I420786,I420751,);
nor I_24618 (I420766,I421010,I420911);
nand I_24619 (I421063,I119681,I119696);
and I_24620 (I421080,I421063,I119693);
DFFARX1 I_24621 (I421080,I2507,I420786,I421106,);
nor I_24622 (I420754,I421106,I421010);
not I_24623 (I421128,I421106);
nor I_24624 (I421145,I421128,I420919);
nor I_24625 (I421162,I420851,I421145);
DFFARX1 I_24626 (I421162,I2507,I420786,I420769,);
nor I_24627 (I421193,I421128,I421010);
nor I_24628 (I421210,I119705,I119696);
nor I_24629 (I420760,I421210,I421193);
not I_24630 (I421241,I421210);
nand I_24631 (I420763,I420970,I421241);
DFFARX1 I_24632 (I421210,I2507,I420786,I420775,);
DFFARX1 I_24633 (I421210,I2507,I420786,I420772,);
not I_24634 (I421330,I2514);
DFFARX1 I_24635 (I855487,I2507,I421330,I421356,);
DFFARX1 I_24636 (I421356,I2507,I421330,I421373,);
not I_24637 (I421322,I421373);
not I_24638 (I421395,I421356);
nand I_24639 (I421412,I855481,I855478);
and I_24640 (I421429,I421412,I855493);
DFFARX1 I_24641 (I421429,I2507,I421330,I421455,);
not I_24642 (I421463,I421455);
DFFARX1 I_24643 (I855481,I2507,I421330,I421489,);
and I_24644 (I421497,I421489,I855475);
nand I_24645 (I421514,I421489,I855475);
nand I_24646 (I421301,I421463,I421514);
DFFARX1 I_24647 (I855475,I2507,I421330,I421554,);
nor I_24648 (I421562,I421554,I421497);
DFFARX1 I_24649 (I421562,I2507,I421330,I421295,);
nor I_24650 (I421310,I421554,I421455);
nand I_24651 (I421607,I855490,I855484);
and I_24652 (I421624,I421607,I855478);
DFFARX1 I_24653 (I421624,I2507,I421330,I421650,);
nor I_24654 (I421298,I421650,I421554);
not I_24655 (I421672,I421650);
nor I_24656 (I421689,I421672,I421463);
nor I_24657 (I421706,I421395,I421689);
DFFARX1 I_24658 (I421706,I2507,I421330,I421313,);
nor I_24659 (I421737,I421672,I421554);
nor I_24660 (I421754,I855496,I855484);
nor I_24661 (I421304,I421754,I421737);
not I_24662 (I421785,I421754);
nand I_24663 (I421307,I421514,I421785);
DFFARX1 I_24664 (I421754,I2507,I421330,I421319,);
DFFARX1 I_24665 (I421754,I2507,I421330,I421316,);
not I_24666 (I421874,I2514);
DFFARX1 I_24667 (I117052,I2507,I421874,I421900,);
DFFARX1 I_24668 (I421900,I2507,I421874,I421917,);
not I_24669 (I421866,I421917);
not I_24670 (I421939,I421900);
nand I_24671 (I421956,I117067,I117046);
and I_24672 (I421973,I421956,I117049);
DFFARX1 I_24673 (I421973,I2507,I421874,I421999,);
not I_24674 (I422007,I421999);
DFFARX1 I_24675 (I117055,I2507,I421874,I422033,);
and I_24676 (I422041,I422033,I117049);
nand I_24677 (I422058,I422033,I117049);
nand I_24678 (I421845,I422007,I422058);
DFFARX1 I_24679 (I117064,I2507,I421874,I422098,);
nor I_24680 (I422106,I422098,I422041);
DFFARX1 I_24681 (I422106,I2507,I421874,I421839,);
nor I_24682 (I421854,I422098,I421999);
nand I_24683 (I422151,I117046,I117061);
and I_24684 (I422168,I422151,I117058);
DFFARX1 I_24685 (I422168,I2507,I421874,I422194,);
nor I_24686 (I421842,I422194,I422098);
not I_24687 (I422216,I422194);
nor I_24688 (I422233,I422216,I422007);
nor I_24689 (I422250,I421939,I422233);
DFFARX1 I_24690 (I422250,I2507,I421874,I421857,);
nor I_24691 (I422281,I422216,I422098);
nor I_24692 (I422298,I117070,I117061);
nor I_24693 (I421848,I422298,I422281);
not I_24694 (I422329,I422298);
nand I_24695 (I421851,I422058,I422329);
DFFARX1 I_24696 (I422298,I2507,I421874,I421863,);
DFFARX1 I_24697 (I422298,I2507,I421874,I421860,);
not I_24698 (I422418,I2514);
DFFARX1 I_24699 (I602399,I2507,I422418,I422444,);
DFFARX1 I_24700 (I422444,I2507,I422418,I422461,);
not I_24701 (I422410,I422461);
not I_24702 (I422483,I422444);
nand I_24703 (I422500,I602396,I602417);
and I_24704 (I422517,I422500,I602420);
DFFARX1 I_24705 (I422517,I2507,I422418,I422543,);
not I_24706 (I422551,I422543);
DFFARX1 I_24707 (I602405,I2507,I422418,I422577,);
and I_24708 (I422585,I422577,I602408);
nand I_24709 (I422602,I422577,I602408);
nand I_24710 (I422389,I422551,I422602);
DFFARX1 I_24711 (I602411,I2507,I422418,I422642,);
nor I_24712 (I422650,I422642,I422585);
DFFARX1 I_24713 (I422650,I2507,I422418,I422383,);
nor I_24714 (I422398,I422642,I422543);
nand I_24715 (I422695,I602396,I602402);
and I_24716 (I422712,I422695,I602414);
DFFARX1 I_24717 (I422712,I2507,I422418,I422738,);
nor I_24718 (I422386,I422738,I422642);
not I_24719 (I422760,I422738);
nor I_24720 (I422777,I422760,I422551);
nor I_24721 (I422794,I422483,I422777);
DFFARX1 I_24722 (I422794,I2507,I422418,I422401,);
nor I_24723 (I422825,I422760,I422642);
nor I_24724 (I422842,I602399,I602402);
nor I_24725 (I422392,I422842,I422825);
not I_24726 (I422873,I422842);
nand I_24727 (I422395,I422602,I422873);
DFFARX1 I_24728 (I422842,I2507,I422418,I422407,);
DFFARX1 I_24729 (I422842,I2507,I422418,I422404,);
not I_24730 (I422962,I2514);
DFFARX1 I_24731 (I1076291,I2507,I422962,I422988,);
DFFARX1 I_24732 (I422988,I2507,I422962,I423005,);
not I_24733 (I422954,I423005);
not I_24734 (I423027,I422988);
nand I_24735 (I423044,I1076303,I1076291);
and I_24736 (I423061,I423044,I1076294);
DFFARX1 I_24737 (I423061,I2507,I422962,I423087,);
not I_24738 (I423095,I423087);
DFFARX1 I_24739 (I1076312,I2507,I422962,I423121,);
and I_24740 (I423129,I423121,I1076288);
nand I_24741 (I423146,I423121,I1076288);
nand I_24742 (I422933,I423095,I423146);
DFFARX1 I_24743 (I1076306,I2507,I422962,I423186,);
nor I_24744 (I423194,I423186,I423129);
DFFARX1 I_24745 (I423194,I2507,I422962,I422927,);
nor I_24746 (I422942,I423186,I423087);
nand I_24747 (I423239,I1076300,I1076297);
and I_24748 (I423256,I423239,I1076309);
DFFARX1 I_24749 (I423256,I2507,I422962,I423282,);
nor I_24750 (I422930,I423282,I423186);
not I_24751 (I423304,I423282);
nor I_24752 (I423321,I423304,I423095);
nor I_24753 (I423338,I423027,I423321);
DFFARX1 I_24754 (I423338,I2507,I422962,I422945,);
nor I_24755 (I423369,I423304,I423186);
nor I_24756 (I423386,I1076288,I1076297);
nor I_24757 (I422936,I423386,I423369);
not I_24758 (I423417,I423386);
nand I_24759 (I422939,I423146,I423417);
DFFARX1 I_24760 (I423386,I2507,I422962,I422951,);
DFFARX1 I_24761 (I423386,I2507,I422962,I422948,);
not I_24762 (I423506,I2514);
DFFARX1 I_24763 (I581591,I2507,I423506,I423532,);
DFFARX1 I_24764 (I423532,I2507,I423506,I423549,);
not I_24765 (I423498,I423549);
not I_24766 (I423571,I423532);
nand I_24767 (I423588,I581588,I581609);
and I_24768 (I423605,I423588,I581612);
DFFARX1 I_24769 (I423605,I2507,I423506,I423631,);
not I_24770 (I423639,I423631);
DFFARX1 I_24771 (I581597,I2507,I423506,I423665,);
and I_24772 (I423673,I423665,I581600);
nand I_24773 (I423690,I423665,I581600);
nand I_24774 (I423477,I423639,I423690);
DFFARX1 I_24775 (I581603,I2507,I423506,I423730,);
nor I_24776 (I423738,I423730,I423673);
DFFARX1 I_24777 (I423738,I2507,I423506,I423471,);
nor I_24778 (I423486,I423730,I423631);
nand I_24779 (I423783,I581588,I581594);
and I_24780 (I423800,I423783,I581606);
DFFARX1 I_24781 (I423800,I2507,I423506,I423826,);
nor I_24782 (I423474,I423826,I423730);
not I_24783 (I423848,I423826);
nor I_24784 (I423865,I423848,I423639);
nor I_24785 (I423882,I423571,I423865);
DFFARX1 I_24786 (I423882,I2507,I423506,I423489,);
nor I_24787 (I423913,I423848,I423730);
nor I_24788 (I423930,I581591,I581594);
nor I_24789 (I423480,I423930,I423913);
not I_24790 (I423961,I423930);
nand I_24791 (I423483,I423690,I423961);
DFFARX1 I_24792 (I423930,I2507,I423506,I423495,);
DFFARX1 I_24793 (I423930,I2507,I423506,I423492,);
not I_24794 (I424050,I2514);
DFFARX1 I_24795 (I1355319,I2507,I424050,I424076,);
DFFARX1 I_24796 (I424076,I2507,I424050,I424093,);
not I_24797 (I424042,I424093);
not I_24798 (I424115,I424076);
nand I_24799 (I424132,I1355295,I1355316);
and I_24800 (I424149,I424132,I1355313);
DFFARX1 I_24801 (I424149,I2507,I424050,I424175,);
not I_24802 (I424183,I424175);
DFFARX1 I_24803 (I1355292,I2507,I424050,I424209,);
and I_24804 (I424217,I424209,I1355304);
nand I_24805 (I424234,I424209,I1355304);
nand I_24806 (I424021,I424183,I424234);
DFFARX1 I_24807 (I1355307,I2507,I424050,I424274,);
nor I_24808 (I424282,I424274,I424217);
DFFARX1 I_24809 (I424282,I2507,I424050,I424015,);
nor I_24810 (I424030,I424274,I424175);
nand I_24811 (I424327,I1355310,I1355298);
and I_24812 (I424344,I424327,I1355301);
DFFARX1 I_24813 (I424344,I2507,I424050,I424370,);
nor I_24814 (I424018,I424370,I424274);
not I_24815 (I424392,I424370);
nor I_24816 (I424409,I424392,I424183);
nor I_24817 (I424426,I424115,I424409);
DFFARX1 I_24818 (I424426,I2507,I424050,I424033,);
nor I_24819 (I424457,I424392,I424274);
nor I_24820 (I424474,I1355292,I1355298);
nor I_24821 (I424024,I424474,I424457);
not I_24822 (I424505,I424474);
nand I_24823 (I424027,I424234,I424505);
DFFARX1 I_24824 (I424474,I2507,I424050,I424039,);
DFFARX1 I_24825 (I424474,I2507,I424050,I424036,);
not I_24826 (I424594,I2514);
DFFARX1 I_24827 (I1221573,I2507,I424594,I424620,);
DFFARX1 I_24828 (I424620,I2507,I424594,I424637,);
not I_24829 (I424586,I424637);
not I_24830 (I424659,I424620);
nand I_24831 (I424676,I1221585,I1221588);
and I_24832 (I424693,I424676,I1221591);
DFFARX1 I_24833 (I424693,I2507,I424594,I424719,);
not I_24834 (I424727,I424719);
DFFARX1 I_24835 (I1221576,I2507,I424594,I424753,);
and I_24836 (I424761,I424753,I1221582);
nand I_24837 (I424778,I424753,I1221582);
nand I_24838 (I424565,I424727,I424778);
DFFARX1 I_24839 (I1221570,I2507,I424594,I424818,);
nor I_24840 (I424826,I424818,I424761);
DFFARX1 I_24841 (I424826,I2507,I424594,I424559,);
nor I_24842 (I424574,I424818,I424719);
nand I_24843 (I424871,I1221573,I1221594);
and I_24844 (I424888,I424871,I1221579);
DFFARX1 I_24845 (I424888,I2507,I424594,I424914,);
nor I_24846 (I424562,I424914,I424818);
not I_24847 (I424936,I424914);
nor I_24848 (I424953,I424936,I424727);
nor I_24849 (I424970,I424659,I424953);
DFFARX1 I_24850 (I424970,I2507,I424594,I424577,);
nor I_24851 (I425001,I424936,I424818);
nor I_24852 (I425018,I1221570,I1221594);
nor I_24853 (I424568,I425018,I425001);
not I_24854 (I425049,I425018);
nand I_24855 (I424571,I424778,I425049);
DFFARX1 I_24856 (I425018,I2507,I424594,I424583,);
DFFARX1 I_24857 (I425018,I2507,I424594,I424580,);
not I_24858 (I425138,I2514);
DFFARX1 I_24859 (I856014,I2507,I425138,I425164,);
DFFARX1 I_24860 (I425164,I2507,I425138,I425181,);
not I_24861 (I425130,I425181);
not I_24862 (I425203,I425164);
nand I_24863 (I425220,I856008,I856005);
and I_24864 (I425237,I425220,I856020);
DFFARX1 I_24865 (I425237,I2507,I425138,I425263,);
not I_24866 (I425271,I425263);
DFFARX1 I_24867 (I856008,I2507,I425138,I425297,);
and I_24868 (I425305,I425297,I856002);
nand I_24869 (I425322,I425297,I856002);
nand I_24870 (I425109,I425271,I425322);
DFFARX1 I_24871 (I856002,I2507,I425138,I425362,);
nor I_24872 (I425370,I425362,I425305);
DFFARX1 I_24873 (I425370,I2507,I425138,I425103,);
nor I_24874 (I425118,I425362,I425263);
nand I_24875 (I425415,I856017,I856011);
and I_24876 (I425432,I425415,I856005);
DFFARX1 I_24877 (I425432,I2507,I425138,I425458,);
nor I_24878 (I425106,I425458,I425362);
not I_24879 (I425480,I425458);
nor I_24880 (I425497,I425480,I425271);
nor I_24881 (I425514,I425203,I425497);
DFFARX1 I_24882 (I425514,I2507,I425138,I425121,);
nor I_24883 (I425545,I425480,I425362);
nor I_24884 (I425562,I856023,I856011);
nor I_24885 (I425112,I425562,I425545);
not I_24886 (I425593,I425562);
nand I_24887 (I425115,I425322,I425593);
DFFARX1 I_24888 (I425562,I2507,I425138,I425127,);
DFFARX1 I_24889 (I425562,I2507,I425138,I425124,);
not I_24890 (I425682,I2514);
DFFARX1 I_24891 (I716265,I2507,I425682,I425708,);
DFFARX1 I_24892 (I425708,I2507,I425682,I425725,);
not I_24893 (I425674,I425725);
not I_24894 (I425747,I425708);
nand I_24895 (I425764,I716286,I716277);
and I_24896 (I425781,I425764,I716265);
DFFARX1 I_24897 (I425781,I2507,I425682,I425807,);
not I_24898 (I425815,I425807);
DFFARX1 I_24899 (I716271,I2507,I425682,I425841,);
and I_24900 (I425849,I425841,I716268);
nand I_24901 (I425866,I425841,I716268);
nand I_24902 (I425653,I425815,I425866);
DFFARX1 I_24903 (I716262,I2507,I425682,I425906,);
nor I_24904 (I425914,I425906,I425849);
DFFARX1 I_24905 (I425914,I2507,I425682,I425647,);
nor I_24906 (I425662,I425906,I425807);
nand I_24907 (I425959,I716262,I716274);
and I_24908 (I425976,I425959,I716283);
DFFARX1 I_24909 (I425976,I2507,I425682,I426002,);
nor I_24910 (I425650,I426002,I425906);
not I_24911 (I426024,I426002);
nor I_24912 (I426041,I426024,I425815);
nor I_24913 (I426058,I425747,I426041);
DFFARX1 I_24914 (I426058,I2507,I425682,I425665,);
nor I_24915 (I426089,I426024,I425906);
nor I_24916 (I426106,I716280,I716274);
nor I_24917 (I425656,I426106,I426089);
not I_24918 (I426137,I426106);
nand I_24919 (I425659,I425866,I426137);
DFFARX1 I_24920 (I426106,I2507,I425682,I425671,);
DFFARX1 I_24921 (I426106,I2507,I425682,I425668,);
not I_24922 (I426226,I2514);
DFFARX1 I_24923 (I759615,I2507,I426226,I426252,);
DFFARX1 I_24924 (I426252,I2507,I426226,I426269,);
not I_24925 (I426218,I426269);
not I_24926 (I426291,I426252);
nand I_24927 (I426308,I759636,I759627);
and I_24928 (I426325,I426308,I759615);
DFFARX1 I_24929 (I426325,I2507,I426226,I426351,);
not I_24930 (I426359,I426351);
DFFARX1 I_24931 (I759621,I2507,I426226,I426385,);
and I_24932 (I426393,I426385,I759618);
nand I_24933 (I426410,I426385,I759618);
nand I_24934 (I426197,I426359,I426410);
DFFARX1 I_24935 (I759612,I2507,I426226,I426450,);
nor I_24936 (I426458,I426450,I426393);
DFFARX1 I_24937 (I426458,I2507,I426226,I426191,);
nor I_24938 (I426206,I426450,I426351);
nand I_24939 (I426503,I759612,I759624);
and I_24940 (I426520,I426503,I759633);
DFFARX1 I_24941 (I426520,I2507,I426226,I426546,);
nor I_24942 (I426194,I426546,I426450);
not I_24943 (I426568,I426546);
nor I_24944 (I426585,I426568,I426359);
nor I_24945 (I426602,I426291,I426585);
DFFARX1 I_24946 (I426602,I2507,I426226,I426209,);
nor I_24947 (I426633,I426568,I426450);
nor I_24948 (I426650,I759630,I759624);
nor I_24949 (I426200,I426650,I426633);
not I_24950 (I426681,I426650);
nand I_24951 (I426203,I426410,I426681);
DFFARX1 I_24952 (I426650,I2507,I426226,I426215,);
DFFARX1 I_24953 (I426650,I2507,I426226,I426212,);
not I_24954 (I426770,I2514);
DFFARX1 I_24955 (I85959,I2507,I426770,I426796,);
DFFARX1 I_24956 (I426796,I2507,I426770,I426813,);
not I_24957 (I426762,I426813);
not I_24958 (I426835,I426796);
nand I_24959 (I426852,I85974,I85953);
and I_24960 (I426869,I426852,I85956);
DFFARX1 I_24961 (I426869,I2507,I426770,I426895,);
not I_24962 (I426903,I426895);
DFFARX1 I_24963 (I85962,I2507,I426770,I426929,);
and I_24964 (I426937,I426929,I85956);
nand I_24965 (I426954,I426929,I85956);
nand I_24966 (I426741,I426903,I426954);
DFFARX1 I_24967 (I85971,I2507,I426770,I426994,);
nor I_24968 (I427002,I426994,I426937);
DFFARX1 I_24969 (I427002,I2507,I426770,I426735,);
nor I_24970 (I426750,I426994,I426895);
nand I_24971 (I427047,I85953,I85968);
and I_24972 (I427064,I427047,I85965);
DFFARX1 I_24973 (I427064,I2507,I426770,I427090,);
nor I_24974 (I426738,I427090,I426994);
not I_24975 (I427112,I427090);
nor I_24976 (I427129,I427112,I426903);
nor I_24977 (I427146,I426835,I427129);
DFFARX1 I_24978 (I427146,I2507,I426770,I426753,);
nor I_24979 (I427177,I427112,I426994);
nor I_24980 (I427194,I85977,I85968);
nor I_24981 (I426744,I427194,I427177);
not I_24982 (I427225,I427194);
nand I_24983 (I426747,I426954,I427225);
DFFARX1 I_24984 (I427194,I2507,I426770,I426759,);
DFFARX1 I_24985 (I427194,I2507,I426770,I426756,);
not I_24986 (I427314,I2514);
DFFARX1 I_24987 (I1366029,I2507,I427314,I427340,);
DFFARX1 I_24988 (I427340,I2507,I427314,I427357,);
not I_24989 (I427306,I427357);
not I_24990 (I427379,I427340);
nand I_24991 (I427396,I1366005,I1366026);
and I_24992 (I427413,I427396,I1366023);
DFFARX1 I_24993 (I427413,I2507,I427314,I427439,);
not I_24994 (I427447,I427439);
DFFARX1 I_24995 (I1366002,I2507,I427314,I427473,);
and I_24996 (I427481,I427473,I1366014);
nand I_24997 (I427498,I427473,I1366014);
nand I_24998 (I427285,I427447,I427498);
DFFARX1 I_24999 (I1366017,I2507,I427314,I427538,);
nor I_25000 (I427546,I427538,I427481);
DFFARX1 I_25001 (I427546,I2507,I427314,I427279,);
nor I_25002 (I427294,I427538,I427439);
nand I_25003 (I427591,I1366020,I1366008);
and I_25004 (I427608,I427591,I1366011);
DFFARX1 I_25005 (I427608,I2507,I427314,I427634,);
nor I_25006 (I427282,I427634,I427538);
not I_25007 (I427656,I427634);
nor I_25008 (I427673,I427656,I427447);
nor I_25009 (I427690,I427379,I427673);
DFFARX1 I_25010 (I427690,I2507,I427314,I427297,);
nor I_25011 (I427721,I427656,I427538);
nor I_25012 (I427738,I1366002,I1366008);
nor I_25013 (I427288,I427738,I427721);
not I_25014 (I427769,I427738);
nand I_25015 (I427291,I427498,I427769);
DFFARX1 I_25016 (I427738,I2507,I427314,I427303,);
DFFARX1 I_25017 (I427738,I2507,I427314,I427300,);
not I_25018 (I427858,I2514);
DFFARX1 I_25019 (I210334,I2507,I427858,I427884,);
DFFARX1 I_25020 (I427884,I2507,I427858,I427901,);
not I_25021 (I427850,I427901);
not I_25022 (I427923,I427884);
nand I_25023 (I427940,I210346,I210325);
and I_25024 (I427957,I427940,I210328);
DFFARX1 I_25025 (I427957,I2507,I427858,I427983,);
not I_25026 (I427991,I427983);
DFFARX1 I_25027 (I210337,I2507,I427858,I428017,);
and I_25028 (I428025,I428017,I210349);
nand I_25029 (I428042,I428017,I210349);
nand I_25030 (I427829,I427991,I428042);
DFFARX1 I_25031 (I210343,I2507,I427858,I428082,);
nor I_25032 (I428090,I428082,I428025);
DFFARX1 I_25033 (I428090,I2507,I427858,I427823,);
nor I_25034 (I427838,I428082,I427983);
nand I_25035 (I428135,I210331,I210328);
and I_25036 (I428152,I428135,I210340);
DFFARX1 I_25037 (I428152,I2507,I427858,I428178,);
nor I_25038 (I427826,I428178,I428082);
not I_25039 (I428200,I428178);
nor I_25040 (I428217,I428200,I427991);
nor I_25041 (I428234,I427923,I428217);
DFFARX1 I_25042 (I428234,I2507,I427858,I427841,);
nor I_25043 (I428265,I428200,I428082);
nor I_25044 (I428282,I210325,I210328);
nor I_25045 (I427832,I428282,I428265);
not I_25046 (I428313,I428282);
nand I_25047 (I427835,I428042,I428313);
DFFARX1 I_25048 (I428282,I2507,I427858,I427847,);
DFFARX1 I_25049 (I428282,I2507,I427858,I427844,);
not I_25050 (I428402,I2514);
DFFARX1 I_25051 (I245439,I2507,I428402,I428428,);
DFFARX1 I_25052 (I428428,I2507,I428402,I428445,);
not I_25053 (I428394,I428445);
not I_25054 (I428467,I428428);
nand I_25055 (I428484,I245451,I245430);
and I_25056 (I428501,I428484,I245433);
DFFARX1 I_25057 (I428501,I2507,I428402,I428527,);
not I_25058 (I428535,I428527);
DFFARX1 I_25059 (I245442,I2507,I428402,I428561,);
and I_25060 (I428569,I428561,I245454);
nand I_25061 (I428586,I428561,I245454);
nand I_25062 (I428373,I428535,I428586);
DFFARX1 I_25063 (I245448,I2507,I428402,I428626,);
nor I_25064 (I428634,I428626,I428569);
DFFARX1 I_25065 (I428634,I2507,I428402,I428367,);
nor I_25066 (I428382,I428626,I428527);
nand I_25067 (I428679,I245436,I245433);
and I_25068 (I428696,I428679,I245445);
DFFARX1 I_25069 (I428696,I2507,I428402,I428722,);
nor I_25070 (I428370,I428722,I428626);
not I_25071 (I428744,I428722);
nor I_25072 (I428761,I428744,I428535);
nor I_25073 (I428778,I428467,I428761);
DFFARX1 I_25074 (I428778,I2507,I428402,I428385,);
nor I_25075 (I428809,I428744,I428626);
nor I_25076 (I428826,I245430,I245433);
nor I_25077 (I428376,I428826,I428809);
not I_25078 (I428857,I428826);
nand I_25079 (I428379,I428586,I428857);
DFFARX1 I_25080 (I428826,I2507,I428402,I428391,);
DFFARX1 I_25081 (I428826,I2507,I428402,I428388,);
not I_25082 (I428946,I2514);
DFFARX1 I_25083 (I746899,I2507,I428946,I428972,);
DFFARX1 I_25084 (I428972,I2507,I428946,I428989,);
not I_25085 (I428938,I428989);
not I_25086 (I429011,I428972);
nand I_25087 (I429028,I746920,I746911);
and I_25088 (I429045,I429028,I746899);
DFFARX1 I_25089 (I429045,I2507,I428946,I429071,);
not I_25090 (I429079,I429071);
DFFARX1 I_25091 (I746905,I2507,I428946,I429105,);
and I_25092 (I429113,I429105,I746902);
nand I_25093 (I429130,I429105,I746902);
nand I_25094 (I428917,I429079,I429130);
DFFARX1 I_25095 (I746896,I2507,I428946,I429170,);
nor I_25096 (I429178,I429170,I429113);
DFFARX1 I_25097 (I429178,I2507,I428946,I428911,);
nor I_25098 (I428926,I429170,I429071);
nand I_25099 (I429223,I746896,I746908);
and I_25100 (I429240,I429223,I746917);
DFFARX1 I_25101 (I429240,I2507,I428946,I429266,);
nor I_25102 (I428914,I429266,I429170);
not I_25103 (I429288,I429266);
nor I_25104 (I429305,I429288,I429079);
nor I_25105 (I429322,I429011,I429305);
DFFARX1 I_25106 (I429322,I2507,I428946,I428929,);
nor I_25107 (I429353,I429288,I429170);
nor I_25108 (I429370,I746914,I746908);
nor I_25109 (I428920,I429370,I429353);
not I_25110 (I429401,I429370);
nand I_25111 (I428923,I429130,I429401);
DFFARX1 I_25112 (I429370,I2507,I428946,I428935,);
DFFARX1 I_25113 (I429370,I2507,I428946,I428932,);
not I_25114 (I429490,I2514);
DFFARX1 I_25115 (I1354724,I2507,I429490,I429516,);
DFFARX1 I_25116 (I429516,I2507,I429490,I429533,);
not I_25117 (I429482,I429533);
not I_25118 (I429555,I429516);
nand I_25119 (I429572,I1354700,I1354721);
and I_25120 (I429589,I429572,I1354718);
DFFARX1 I_25121 (I429589,I2507,I429490,I429615,);
not I_25122 (I429623,I429615);
DFFARX1 I_25123 (I1354697,I2507,I429490,I429649,);
and I_25124 (I429657,I429649,I1354709);
nand I_25125 (I429674,I429649,I1354709);
nand I_25126 (I429461,I429623,I429674);
DFFARX1 I_25127 (I1354712,I2507,I429490,I429714,);
nor I_25128 (I429722,I429714,I429657);
DFFARX1 I_25129 (I429722,I2507,I429490,I429455,);
nor I_25130 (I429470,I429714,I429615);
nand I_25131 (I429767,I1354715,I1354703);
and I_25132 (I429784,I429767,I1354706);
DFFARX1 I_25133 (I429784,I2507,I429490,I429810,);
nor I_25134 (I429458,I429810,I429714);
not I_25135 (I429832,I429810);
nor I_25136 (I429849,I429832,I429623);
nor I_25137 (I429866,I429555,I429849);
DFFARX1 I_25138 (I429866,I2507,I429490,I429473,);
nor I_25139 (I429897,I429832,I429714);
nor I_25140 (I429914,I1354697,I1354703);
nor I_25141 (I429464,I429914,I429897);
not I_25142 (I429945,I429914);
nand I_25143 (I429467,I429674,I429945);
DFFARX1 I_25144 (I429914,I2507,I429490,I429479,);
DFFARX1 I_25145 (I429914,I2507,I429490,I429476,);
not I_25146 (I430034,I2514);
DFFARX1 I_25147 (I560783,I2507,I430034,I430060,);
DFFARX1 I_25148 (I430060,I2507,I430034,I430077,);
not I_25149 (I430026,I430077);
not I_25150 (I430099,I430060);
nand I_25151 (I430116,I560780,I560801);
and I_25152 (I430133,I430116,I560804);
DFFARX1 I_25153 (I430133,I2507,I430034,I430159,);
not I_25154 (I430167,I430159);
DFFARX1 I_25155 (I560789,I2507,I430034,I430193,);
and I_25156 (I430201,I430193,I560792);
nand I_25157 (I430218,I430193,I560792);
nand I_25158 (I430005,I430167,I430218);
DFFARX1 I_25159 (I560795,I2507,I430034,I430258,);
nor I_25160 (I430266,I430258,I430201);
DFFARX1 I_25161 (I430266,I2507,I430034,I429999,);
nor I_25162 (I430014,I430258,I430159);
nand I_25163 (I430311,I560780,I560786);
and I_25164 (I430328,I430311,I560798);
DFFARX1 I_25165 (I430328,I2507,I430034,I430354,);
nor I_25166 (I430002,I430354,I430258);
not I_25167 (I430376,I430354);
nor I_25168 (I430393,I430376,I430167);
nor I_25169 (I430410,I430099,I430393);
DFFARX1 I_25170 (I430410,I2507,I430034,I430017,);
nor I_25171 (I430441,I430376,I430258);
nor I_25172 (I430458,I560783,I560786);
nor I_25173 (I430008,I430458,I430441);
not I_25174 (I430489,I430458);
nand I_25175 (I430011,I430218,I430489);
DFFARX1 I_25176 (I430458,I2507,I430034,I430023,);
DFFARX1 I_25177 (I430458,I2507,I430034,I430020,);
not I_25178 (I430578,I2514);
DFFARX1 I_25179 (I717999,I2507,I430578,I430604,);
DFFARX1 I_25180 (I430604,I2507,I430578,I430621,);
not I_25181 (I430570,I430621);
not I_25182 (I430643,I430604);
nand I_25183 (I430660,I718020,I718011);
and I_25184 (I430677,I430660,I717999);
DFFARX1 I_25185 (I430677,I2507,I430578,I430703,);
not I_25186 (I430711,I430703);
DFFARX1 I_25187 (I718005,I2507,I430578,I430737,);
and I_25188 (I430745,I430737,I718002);
nand I_25189 (I430762,I430737,I718002);
nand I_25190 (I430549,I430711,I430762);
DFFARX1 I_25191 (I717996,I2507,I430578,I430802,);
nor I_25192 (I430810,I430802,I430745);
DFFARX1 I_25193 (I430810,I2507,I430578,I430543,);
nor I_25194 (I430558,I430802,I430703);
nand I_25195 (I430855,I717996,I718008);
and I_25196 (I430872,I430855,I718017);
DFFARX1 I_25197 (I430872,I2507,I430578,I430898,);
nor I_25198 (I430546,I430898,I430802);
not I_25199 (I430920,I430898);
nor I_25200 (I430937,I430920,I430711);
nor I_25201 (I430954,I430643,I430937);
DFFARX1 I_25202 (I430954,I2507,I430578,I430561,);
nor I_25203 (I430985,I430920,I430802);
nor I_25204 (I431002,I718014,I718008);
nor I_25205 (I430552,I431002,I430985);
not I_25206 (I431033,I431002);
nand I_25207 (I430555,I430762,I431033);
DFFARX1 I_25208 (I431002,I2507,I430578,I430567,);
DFFARX1 I_25209 (I431002,I2507,I430578,I430564,);
not I_25210 (I431122,I2514);
DFFARX1 I_25211 (I1158367,I2507,I431122,I431148,);
DFFARX1 I_25212 (I431148,I2507,I431122,I431165,);
not I_25213 (I431114,I431165);
not I_25214 (I431187,I431148);
nand I_25215 (I431204,I1158379,I1158367);
and I_25216 (I431221,I431204,I1158370);
DFFARX1 I_25217 (I431221,I2507,I431122,I431247,);
not I_25218 (I431255,I431247);
DFFARX1 I_25219 (I1158388,I2507,I431122,I431281,);
and I_25220 (I431289,I431281,I1158364);
nand I_25221 (I431306,I431281,I1158364);
nand I_25222 (I431093,I431255,I431306);
DFFARX1 I_25223 (I1158382,I2507,I431122,I431346,);
nor I_25224 (I431354,I431346,I431289);
DFFARX1 I_25225 (I431354,I2507,I431122,I431087,);
nor I_25226 (I431102,I431346,I431247);
nand I_25227 (I431399,I1158376,I1158373);
and I_25228 (I431416,I431399,I1158385);
DFFARX1 I_25229 (I431416,I2507,I431122,I431442,);
nor I_25230 (I431090,I431442,I431346);
not I_25231 (I431464,I431442);
nor I_25232 (I431481,I431464,I431255);
nor I_25233 (I431498,I431187,I431481);
DFFARX1 I_25234 (I431498,I2507,I431122,I431105,);
nor I_25235 (I431529,I431464,I431346);
nor I_25236 (I431546,I1158364,I1158373);
nor I_25237 (I431096,I431546,I431529);
not I_25238 (I431577,I431546);
nand I_25239 (I431099,I431306,I431577);
DFFARX1 I_25240 (I431546,I2507,I431122,I431111,);
DFFARX1 I_25241 (I431546,I2507,I431122,I431108,);
not I_25242 (I431666,I2514);
DFFARX1 I_25243 (I230564,I2507,I431666,I431692,);
DFFARX1 I_25244 (I431692,I2507,I431666,I431709,);
not I_25245 (I431658,I431709);
not I_25246 (I431731,I431692);
nand I_25247 (I431748,I230576,I230555);
and I_25248 (I431765,I431748,I230558);
DFFARX1 I_25249 (I431765,I2507,I431666,I431791,);
not I_25250 (I431799,I431791);
DFFARX1 I_25251 (I230567,I2507,I431666,I431825,);
and I_25252 (I431833,I431825,I230579);
nand I_25253 (I431850,I431825,I230579);
nand I_25254 (I431637,I431799,I431850);
DFFARX1 I_25255 (I230573,I2507,I431666,I431890,);
nor I_25256 (I431898,I431890,I431833);
DFFARX1 I_25257 (I431898,I2507,I431666,I431631,);
nor I_25258 (I431646,I431890,I431791);
nand I_25259 (I431943,I230561,I230558);
and I_25260 (I431960,I431943,I230570);
DFFARX1 I_25261 (I431960,I2507,I431666,I431986,);
nor I_25262 (I431634,I431986,I431890);
not I_25263 (I432008,I431986);
nor I_25264 (I432025,I432008,I431799);
nor I_25265 (I432042,I431731,I432025);
DFFARX1 I_25266 (I432042,I2507,I431666,I431649,);
nor I_25267 (I432073,I432008,I431890);
nor I_25268 (I432090,I230555,I230558);
nor I_25269 (I431640,I432090,I432073);
not I_25270 (I432121,I432090);
nand I_25271 (I431643,I431850,I432121);
DFFARX1 I_25272 (I432090,I2507,I431666,I431655,);
DFFARX1 I_25273 (I432090,I2507,I431666,I431652,);
not I_25274 (I432210,I2514);
DFFARX1 I_25275 (I103350,I2507,I432210,I432236,);
DFFARX1 I_25276 (I432236,I2507,I432210,I432253,);
not I_25277 (I432202,I432253);
not I_25278 (I432275,I432236);
nand I_25279 (I432292,I103365,I103344);
and I_25280 (I432309,I432292,I103347);
DFFARX1 I_25281 (I432309,I2507,I432210,I432335,);
not I_25282 (I432343,I432335);
DFFARX1 I_25283 (I103353,I2507,I432210,I432369,);
and I_25284 (I432377,I432369,I103347);
nand I_25285 (I432394,I432369,I103347);
nand I_25286 (I432181,I432343,I432394);
DFFARX1 I_25287 (I103362,I2507,I432210,I432434,);
nor I_25288 (I432442,I432434,I432377);
DFFARX1 I_25289 (I432442,I2507,I432210,I432175,);
nor I_25290 (I432190,I432434,I432335);
nand I_25291 (I432487,I103344,I103359);
and I_25292 (I432504,I432487,I103356);
DFFARX1 I_25293 (I432504,I2507,I432210,I432530,);
nor I_25294 (I432178,I432530,I432434);
not I_25295 (I432552,I432530);
nor I_25296 (I432569,I432552,I432343);
nor I_25297 (I432586,I432275,I432569);
DFFARX1 I_25298 (I432586,I2507,I432210,I432193,);
nor I_25299 (I432617,I432552,I432434);
nor I_25300 (I432634,I103368,I103359);
nor I_25301 (I432184,I432634,I432617);
not I_25302 (I432665,I432634);
nand I_25303 (I432187,I432394,I432665);
DFFARX1 I_25304 (I432634,I2507,I432210,I432199,);
DFFARX1 I_25305 (I432634,I2507,I432210,I432196,);
not I_25306 (I432754,I2514);
DFFARX1 I_25307 (I1125999,I2507,I432754,I432780,);
DFFARX1 I_25308 (I432780,I2507,I432754,I432797,);
not I_25309 (I432746,I432797);
not I_25310 (I432819,I432780);
nand I_25311 (I432836,I1126011,I1125999);
and I_25312 (I432853,I432836,I1126002);
DFFARX1 I_25313 (I432853,I2507,I432754,I432879,);
not I_25314 (I432887,I432879);
DFFARX1 I_25315 (I1126020,I2507,I432754,I432913,);
and I_25316 (I432921,I432913,I1125996);
nand I_25317 (I432938,I432913,I1125996);
nand I_25318 (I432725,I432887,I432938);
DFFARX1 I_25319 (I1126014,I2507,I432754,I432978,);
nor I_25320 (I432986,I432978,I432921);
DFFARX1 I_25321 (I432986,I2507,I432754,I432719,);
nor I_25322 (I432734,I432978,I432879);
nand I_25323 (I433031,I1126008,I1126005);
and I_25324 (I433048,I433031,I1126017);
DFFARX1 I_25325 (I433048,I2507,I432754,I433074,);
nor I_25326 (I432722,I433074,I432978);
not I_25327 (I433096,I433074);
nor I_25328 (I433113,I433096,I432887);
nor I_25329 (I433130,I432819,I433113);
DFFARX1 I_25330 (I433130,I2507,I432754,I432737,);
nor I_25331 (I433161,I433096,I432978);
nor I_25332 (I433178,I1125996,I1126005);
nor I_25333 (I432728,I433178,I433161);
not I_25334 (I433209,I433178);
nand I_25335 (I432731,I432938,I433209);
DFFARX1 I_25336 (I433178,I2507,I432754,I432743,);
DFFARX1 I_25337 (I433178,I2507,I432754,I432740,);
not I_25338 (I433298,I2514);
DFFARX1 I_25339 (I782761,I2507,I433298,I433324,);
DFFARX1 I_25340 (I433324,I2507,I433298,I433341,);
not I_25341 (I433290,I433341);
not I_25342 (I433363,I433324);
nand I_25343 (I433380,I782755,I782752);
and I_25344 (I433397,I433380,I782767);
DFFARX1 I_25345 (I433397,I2507,I433298,I433423,);
not I_25346 (I433431,I433423);
DFFARX1 I_25347 (I782755,I2507,I433298,I433457,);
and I_25348 (I433465,I433457,I782749);
nand I_25349 (I433482,I433457,I782749);
nand I_25350 (I433269,I433431,I433482);
DFFARX1 I_25351 (I782749,I2507,I433298,I433522,);
nor I_25352 (I433530,I433522,I433465);
DFFARX1 I_25353 (I433530,I2507,I433298,I433263,);
nor I_25354 (I433278,I433522,I433423);
nand I_25355 (I433575,I782764,I782758);
and I_25356 (I433592,I433575,I782752);
DFFARX1 I_25357 (I433592,I2507,I433298,I433618,);
nor I_25358 (I433266,I433618,I433522);
not I_25359 (I433640,I433618);
nor I_25360 (I433657,I433640,I433431);
nor I_25361 (I433674,I433363,I433657);
DFFARX1 I_25362 (I433674,I2507,I433298,I433281,);
nor I_25363 (I433705,I433640,I433522);
nor I_25364 (I433722,I782770,I782758);
nor I_25365 (I433272,I433722,I433705);
not I_25366 (I433753,I433722);
nand I_25367 (I433275,I433482,I433753);
DFFARX1 I_25368 (I433722,I2507,I433298,I433287,);
DFFARX1 I_25369 (I433722,I2507,I433298,I433284,);
not I_25370 (I433842,I2514);
DFFARX1 I_25371 (I1307124,I2507,I433842,I433868,);
DFFARX1 I_25372 (I433868,I2507,I433842,I433885,);
not I_25373 (I433834,I433885);
not I_25374 (I433907,I433868);
nand I_25375 (I433924,I1307100,I1307121);
and I_25376 (I433941,I433924,I1307118);
DFFARX1 I_25377 (I433941,I2507,I433842,I433967,);
not I_25378 (I433975,I433967);
DFFARX1 I_25379 (I1307097,I2507,I433842,I434001,);
and I_25380 (I434009,I434001,I1307109);
nand I_25381 (I434026,I434001,I1307109);
nand I_25382 (I433813,I433975,I434026);
DFFARX1 I_25383 (I1307112,I2507,I433842,I434066,);
nor I_25384 (I434074,I434066,I434009);
DFFARX1 I_25385 (I434074,I2507,I433842,I433807,);
nor I_25386 (I433822,I434066,I433967);
nand I_25387 (I434119,I1307115,I1307103);
and I_25388 (I434136,I434119,I1307106);
DFFARX1 I_25389 (I434136,I2507,I433842,I434162,);
nor I_25390 (I433810,I434162,I434066);
not I_25391 (I434184,I434162);
nor I_25392 (I434201,I434184,I433975);
nor I_25393 (I434218,I433907,I434201);
DFFARX1 I_25394 (I434218,I2507,I433842,I433825,);
nor I_25395 (I434249,I434184,I434066);
nor I_25396 (I434266,I1307097,I1307103);
nor I_25397 (I433816,I434266,I434249);
not I_25398 (I434297,I434266);
nand I_25399 (I433819,I434026,I434297);
DFFARX1 I_25400 (I434266,I2507,I433842,I433831,);
DFFARX1 I_25401 (I434266,I2507,I433842,I433828,);
not I_25402 (I434386,I2514);
DFFARX1 I_25403 (I342963,I2507,I434386,I434412,);
DFFARX1 I_25404 (I434412,I2507,I434386,I434429,);
not I_25405 (I434378,I434429);
not I_25406 (I434451,I434412);
nand I_25407 (I434468,I342942,I342966);
and I_25408 (I434485,I434468,I342969);
DFFARX1 I_25409 (I434485,I2507,I434386,I434511,);
not I_25410 (I434519,I434511);
DFFARX1 I_25411 (I342951,I2507,I434386,I434545,);
and I_25412 (I434553,I434545,I342957);
nand I_25413 (I434570,I434545,I342957);
nand I_25414 (I434357,I434519,I434570);
DFFARX1 I_25415 (I342945,I2507,I434386,I434610,);
nor I_25416 (I434618,I434610,I434553);
DFFARX1 I_25417 (I434618,I2507,I434386,I434351,);
nor I_25418 (I434366,I434610,I434511);
nand I_25419 (I434663,I342954,I342942);
and I_25420 (I434680,I434663,I342948);
DFFARX1 I_25421 (I434680,I2507,I434386,I434706,);
nor I_25422 (I434354,I434706,I434610);
not I_25423 (I434728,I434706);
nor I_25424 (I434745,I434728,I434519);
nor I_25425 (I434762,I434451,I434745);
DFFARX1 I_25426 (I434762,I2507,I434386,I434369,);
nor I_25427 (I434793,I434728,I434610);
nor I_25428 (I434810,I342960,I342942);
nor I_25429 (I434360,I434810,I434793);
not I_25430 (I434841,I434810);
nand I_25431 (I434363,I434570,I434841);
DFFARX1 I_25432 (I434810,I2507,I434386,I434375,);
DFFARX1 I_25433 (I434810,I2507,I434386,I434372,);
not I_25434 (I434930,I2514);
DFFARX1 I_25435 (I967035,I2507,I434930,I434956,);
DFFARX1 I_25436 (I434956,I2507,I434930,I434973,);
not I_25437 (I434922,I434973);
not I_25438 (I434995,I434956);
nand I_25439 (I435012,I967050,I967038);
and I_25440 (I435029,I435012,I967029);
DFFARX1 I_25441 (I435029,I2507,I434930,I435055,);
not I_25442 (I435063,I435055);
DFFARX1 I_25443 (I967041,I2507,I434930,I435089,);
and I_25444 (I435097,I435089,I967032);
nand I_25445 (I435114,I435089,I967032);
nand I_25446 (I434901,I435063,I435114);
DFFARX1 I_25447 (I967047,I2507,I434930,I435154,);
nor I_25448 (I435162,I435154,I435097);
DFFARX1 I_25449 (I435162,I2507,I434930,I434895,);
nor I_25450 (I434910,I435154,I435055);
nand I_25451 (I435207,I967056,I967044);
and I_25452 (I435224,I435207,I967053);
DFFARX1 I_25453 (I435224,I2507,I434930,I435250,);
nor I_25454 (I434898,I435250,I435154);
not I_25455 (I435272,I435250);
nor I_25456 (I435289,I435272,I435063);
nor I_25457 (I435306,I434995,I435289);
DFFARX1 I_25458 (I435306,I2507,I434930,I434913,);
nor I_25459 (I435337,I435272,I435154);
nor I_25460 (I435354,I967029,I967044);
nor I_25461 (I434904,I435354,I435337);
not I_25462 (I435385,I435354);
nand I_25463 (I434907,I435114,I435385);
DFFARX1 I_25464 (I435354,I2507,I434930,I434919,);
DFFARX1 I_25465 (I435354,I2507,I434930,I434916,);
not I_25466 (I435474,I2514);
DFFARX1 I_25467 (I1223205,I2507,I435474,I435500,);
DFFARX1 I_25468 (I435500,I2507,I435474,I435517,);
not I_25469 (I435466,I435517);
not I_25470 (I435539,I435500);
nand I_25471 (I435556,I1223217,I1223220);
and I_25472 (I435573,I435556,I1223223);
DFFARX1 I_25473 (I435573,I2507,I435474,I435599,);
not I_25474 (I435607,I435599);
DFFARX1 I_25475 (I1223208,I2507,I435474,I435633,);
and I_25476 (I435641,I435633,I1223214);
nand I_25477 (I435658,I435633,I1223214);
nand I_25478 (I435445,I435607,I435658);
DFFARX1 I_25479 (I1223202,I2507,I435474,I435698,);
nor I_25480 (I435706,I435698,I435641);
DFFARX1 I_25481 (I435706,I2507,I435474,I435439,);
nor I_25482 (I435454,I435698,I435599);
nand I_25483 (I435751,I1223205,I1223226);
and I_25484 (I435768,I435751,I1223211);
DFFARX1 I_25485 (I435768,I2507,I435474,I435794,);
nor I_25486 (I435442,I435794,I435698);
not I_25487 (I435816,I435794);
nor I_25488 (I435833,I435816,I435607);
nor I_25489 (I435850,I435539,I435833);
DFFARX1 I_25490 (I435850,I2507,I435474,I435457,);
nor I_25491 (I435881,I435816,I435698);
nor I_25492 (I435898,I1223202,I1223226);
nor I_25493 (I435448,I435898,I435881);
not I_25494 (I435929,I435898);
nand I_25495 (I435451,I435658,I435929);
DFFARX1 I_25496 (I435898,I2507,I435474,I435463,);
DFFARX1 I_25497 (I435898,I2507,I435474,I435460,);
not I_25498 (I436018,I2514);
DFFARX1 I_25499 (I1389829,I2507,I436018,I436044,);
DFFARX1 I_25500 (I436044,I2507,I436018,I436061,);
not I_25501 (I436010,I436061);
not I_25502 (I436083,I436044);
nand I_25503 (I436100,I1389805,I1389826);
and I_25504 (I436117,I436100,I1389823);
DFFARX1 I_25505 (I436117,I2507,I436018,I436143,);
not I_25506 (I436151,I436143);
DFFARX1 I_25507 (I1389802,I2507,I436018,I436177,);
and I_25508 (I436185,I436177,I1389814);
nand I_25509 (I436202,I436177,I1389814);
nand I_25510 (I435989,I436151,I436202);
DFFARX1 I_25511 (I1389817,I2507,I436018,I436242,);
nor I_25512 (I436250,I436242,I436185);
DFFARX1 I_25513 (I436250,I2507,I436018,I435983,);
nor I_25514 (I435998,I436242,I436143);
nand I_25515 (I436295,I1389820,I1389808);
and I_25516 (I436312,I436295,I1389811);
DFFARX1 I_25517 (I436312,I2507,I436018,I436338,);
nor I_25518 (I435986,I436338,I436242);
not I_25519 (I436360,I436338);
nor I_25520 (I436377,I436360,I436151);
nor I_25521 (I436394,I436083,I436377);
DFFARX1 I_25522 (I436394,I2507,I436018,I436001,);
nor I_25523 (I436425,I436360,I436242);
nor I_25524 (I436442,I1389802,I1389808);
nor I_25525 (I435992,I436442,I436425);
not I_25526 (I436473,I436442);
nand I_25527 (I435995,I436202,I436473);
DFFARX1 I_25528 (I436442,I2507,I436018,I436007,);
DFFARX1 I_25529 (I436442,I2507,I436018,I436004,);
not I_25530 (I436562,I2514);
DFFARX1 I_25531 (I1194781,I2507,I436562,I436588,);
DFFARX1 I_25532 (I436588,I2507,I436562,I436605,);
not I_25533 (I436554,I436605);
not I_25534 (I436627,I436588);
nand I_25535 (I436644,I1194793,I1194781);
and I_25536 (I436661,I436644,I1194784);
DFFARX1 I_25537 (I436661,I2507,I436562,I436687,);
not I_25538 (I436695,I436687);
DFFARX1 I_25539 (I1194802,I2507,I436562,I436721,);
and I_25540 (I436729,I436721,I1194778);
nand I_25541 (I436746,I436721,I1194778);
nand I_25542 (I436533,I436695,I436746);
DFFARX1 I_25543 (I1194796,I2507,I436562,I436786,);
nor I_25544 (I436794,I436786,I436729);
DFFARX1 I_25545 (I436794,I2507,I436562,I436527,);
nor I_25546 (I436542,I436786,I436687);
nand I_25547 (I436839,I1194790,I1194787);
and I_25548 (I436856,I436839,I1194799);
DFFARX1 I_25549 (I436856,I2507,I436562,I436882,);
nor I_25550 (I436530,I436882,I436786);
not I_25551 (I436904,I436882);
nor I_25552 (I436921,I436904,I436695);
nor I_25553 (I436938,I436627,I436921);
DFFARX1 I_25554 (I436938,I2507,I436562,I436545,);
nor I_25555 (I436969,I436904,I436786);
nor I_25556 (I436986,I1194778,I1194787);
nor I_25557 (I436536,I436986,I436969);
not I_25558 (I437017,I436986);
nand I_25559 (I436539,I436746,I437017);
DFFARX1 I_25560 (I436986,I2507,I436562,I436551,);
DFFARX1 I_25561 (I436986,I2507,I436562,I436548,);
not I_25562 (I437106,I2514);
DFFARX1 I_25563 (I332950,I2507,I437106,I437132,);
DFFARX1 I_25564 (I437132,I2507,I437106,I437149,);
not I_25565 (I437098,I437149);
not I_25566 (I437171,I437132);
nand I_25567 (I437188,I332929,I332953);
and I_25568 (I437205,I437188,I332956);
DFFARX1 I_25569 (I437205,I2507,I437106,I437231,);
not I_25570 (I437239,I437231);
DFFARX1 I_25571 (I332938,I2507,I437106,I437265,);
and I_25572 (I437273,I437265,I332944);
nand I_25573 (I437290,I437265,I332944);
nand I_25574 (I437077,I437239,I437290);
DFFARX1 I_25575 (I332932,I2507,I437106,I437330,);
nor I_25576 (I437338,I437330,I437273);
DFFARX1 I_25577 (I437338,I2507,I437106,I437071,);
nor I_25578 (I437086,I437330,I437231);
nand I_25579 (I437383,I332941,I332929);
and I_25580 (I437400,I437383,I332935);
DFFARX1 I_25581 (I437400,I2507,I437106,I437426,);
nor I_25582 (I437074,I437426,I437330);
not I_25583 (I437448,I437426);
nor I_25584 (I437465,I437448,I437239);
nor I_25585 (I437482,I437171,I437465);
DFFARX1 I_25586 (I437482,I2507,I437106,I437089,);
nor I_25587 (I437513,I437448,I437330);
nor I_25588 (I437530,I332947,I332929);
nor I_25589 (I437080,I437530,I437513);
not I_25590 (I437561,I437530);
nand I_25591 (I437083,I437290,I437561);
DFFARX1 I_25592 (I437530,I2507,I437106,I437095,);
DFFARX1 I_25593 (I437530,I2507,I437106,I437092,);
not I_25594 (I437650,I2514);
DFFARX1 I_25595 (I781707,I2507,I437650,I437676,);
DFFARX1 I_25596 (I437676,I2507,I437650,I437693,);
not I_25597 (I437642,I437693);
not I_25598 (I437715,I437676);
nand I_25599 (I437732,I781701,I781698);
and I_25600 (I437749,I437732,I781713);
DFFARX1 I_25601 (I437749,I2507,I437650,I437775,);
not I_25602 (I437783,I437775);
DFFARX1 I_25603 (I781701,I2507,I437650,I437809,);
and I_25604 (I437817,I437809,I781695);
nand I_25605 (I437834,I437809,I781695);
nand I_25606 (I437621,I437783,I437834);
DFFARX1 I_25607 (I781695,I2507,I437650,I437874,);
nor I_25608 (I437882,I437874,I437817);
DFFARX1 I_25609 (I437882,I2507,I437650,I437615,);
nor I_25610 (I437630,I437874,I437775);
nand I_25611 (I437927,I781710,I781704);
and I_25612 (I437944,I437927,I781698);
DFFARX1 I_25613 (I437944,I2507,I437650,I437970,);
nor I_25614 (I437618,I437970,I437874);
not I_25615 (I437992,I437970);
nor I_25616 (I438009,I437992,I437783);
nor I_25617 (I438026,I437715,I438009);
DFFARX1 I_25618 (I438026,I2507,I437650,I437633,);
nor I_25619 (I438057,I437992,I437874);
nor I_25620 (I438074,I781716,I781704);
nor I_25621 (I437624,I438074,I438057);
not I_25622 (I438105,I438074);
nand I_25623 (I437627,I437834,I438105);
DFFARX1 I_25624 (I438074,I2507,I437650,I437639,);
DFFARX1 I_25625 (I438074,I2507,I437650,I437636,);
not I_25626 (I438194,I2514);
DFFARX1 I_25627 (I976079,I2507,I438194,I438220,);
DFFARX1 I_25628 (I438220,I2507,I438194,I438237,);
not I_25629 (I438186,I438237);
not I_25630 (I438259,I438220);
nand I_25631 (I438276,I976094,I976082);
and I_25632 (I438293,I438276,I976073);
DFFARX1 I_25633 (I438293,I2507,I438194,I438319,);
not I_25634 (I438327,I438319);
DFFARX1 I_25635 (I976085,I2507,I438194,I438353,);
and I_25636 (I438361,I438353,I976076);
nand I_25637 (I438378,I438353,I976076);
nand I_25638 (I438165,I438327,I438378);
DFFARX1 I_25639 (I976091,I2507,I438194,I438418,);
nor I_25640 (I438426,I438418,I438361);
DFFARX1 I_25641 (I438426,I2507,I438194,I438159,);
nor I_25642 (I438174,I438418,I438319);
nand I_25643 (I438471,I976100,I976088);
and I_25644 (I438488,I438471,I976097);
DFFARX1 I_25645 (I438488,I2507,I438194,I438514,);
nor I_25646 (I438162,I438514,I438418);
not I_25647 (I438536,I438514);
nor I_25648 (I438553,I438536,I438327);
nor I_25649 (I438570,I438259,I438553);
DFFARX1 I_25650 (I438570,I2507,I438194,I438177,);
nor I_25651 (I438601,I438536,I438418);
nor I_25652 (I438618,I976073,I976088);
nor I_25653 (I438168,I438618,I438601);
not I_25654 (I438649,I438618);
nand I_25655 (I438171,I438378,I438649);
DFFARX1 I_25656 (I438618,I2507,I438194,I438183,);
DFFARX1 I_25657 (I438618,I2507,I438194,I438180,);
not I_25658 (I438738,I2514);
DFFARX1 I_25659 (I74365,I2507,I438738,I438764,);
DFFARX1 I_25660 (I438764,I2507,I438738,I438781,);
not I_25661 (I438730,I438781);
not I_25662 (I438803,I438764);
nand I_25663 (I438820,I74380,I74359);
and I_25664 (I438837,I438820,I74362);
DFFARX1 I_25665 (I438837,I2507,I438738,I438863,);
not I_25666 (I438871,I438863);
DFFARX1 I_25667 (I74368,I2507,I438738,I438897,);
and I_25668 (I438905,I438897,I74362);
nand I_25669 (I438922,I438897,I74362);
nand I_25670 (I438709,I438871,I438922);
DFFARX1 I_25671 (I74377,I2507,I438738,I438962,);
nor I_25672 (I438970,I438962,I438905);
DFFARX1 I_25673 (I438970,I2507,I438738,I438703,);
nor I_25674 (I438718,I438962,I438863);
nand I_25675 (I439015,I74359,I74374);
and I_25676 (I439032,I439015,I74371);
DFFARX1 I_25677 (I439032,I2507,I438738,I439058,);
nor I_25678 (I438706,I439058,I438962);
not I_25679 (I439080,I439058);
nor I_25680 (I439097,I439080,I438871);
nor I_25681 (I439114,I438803,I439097);
DFFARX1 I_25682 (I439114,I2507,I438738,I438721,);
nor I_25683 (I439145,I439080,I438962);
nor I_25684 (I439162,I74383,I74374);
nor I_25685 (I438712,I439162,I439145);
not I_25686 (I439193,I439162);
nand I_25687 (I438715,I438922,I439193);
DFFARX1 I_25688 (I439162,I2507,I438738,I438727,);
DFFARX1 I_25689 (I439162,I2507,I438738,I438724,);
not I_25690 (I439282,I2514);
DFFARX1 I_25691 (I782234,I2507,I439282,I439308,);
DFFARX1 I_25692 (I439308,I2507,I439282,I439325,);
not I_25693 (I439274,I439325);
not I_25694 (I439347,I439308);
nand I_25695 (I439364,I782228,I782225);
and I_25696 (I439381,I439364,I782240);
DFFARX1 I_25697 (I439381,I2507,I439282,I439407,);
not I_25698 (I439415,I439407);
DFFARX1 I_25699 (I782228,I2507,I439282,I439441,);
and I_25700 (I439449,I439441,I782222);
nand I_25701 (I439466,I439441,I782222);
nand I_25702 (I439253,I439415,I439466);
DFFARX1 I_25703 (I782222,I2507,I439282,I439506,);
nor I_25704 (I439514,I439506,I439449);
DFFARX1 I_25705 (I439514,I2507,I439282,I439247,);
nor I_25706 (I439262,I439506,I439407);
nand I_25707 (I439559,I782237,I782231);
and I_25708 (I439576,I439559,I782225);
DFFARX1 I_25709 (I439576,I2507,I439282,I439602,);
nor I_25710 (I439250,I439602,I439506);
not I_25711 (I439624,I439602);
nor I_25712 (I439641,I439624,I439415);
nor I_25713 (I439658,I439347,I439641);
DFFARX1 I_25714 (I439658,I2507,I439282,I439265,);
nor I_25715 (I439689,I439624,I439506);
nor I_25716 (I439706,I782243,I782231);
nor I_25717 (I439256,I439706,I439689);
not I_25718 (I439737,I439706);
nand I_25719 (I439259,I439466,I439737);
DFFARX1 I_25720 (I439706,I2507,I439282,I439271,);
DFFARX1 I_25721 (I439706,I2507,I439282,I439268,);
not I_25722 (I439826,I2514);
DFFARX1 I_25723 (I884993,I2507,I439826,I439852,);
DFFARX1 I_25724 (I439852,I2507,I439826,I439869,);
not I_25725 (I439818,I439869);
not I_25726 (I439891,I439852);
nand I_25727 (I439908,I885008,I884996);
and I_25728 (I439925,I439908,I884987);
DFFARX1 I_25729 (I439925,I2507,I439826,I439951,);
not I_25730 (I439959,I439951);
DFFARX1 I_25731 (I884999,I2507,I439826,I439985,);
and I_25732 (I439993,I439985,I884990);
nand I_25733 (I440010,I439985,I884990);
nand I_25734 (I439797,I439959,I440010);
DFFARX1 I_25735 (I885005,I2507,I439826,I440050,);
nor I_25736 (I440058,I440050,I439993);
DFFARX1 I_25737 (I440058,I2507,I439826,I439791,);
nor I_25738 (I439806,I440050,I439951);
nand I_25739 (I440103,I885014,I885002);
and I_25740 (I440120,I440103,I885011);
DFFARX1 I_25741 (I440120,I2507,I439826,I440146,);
nor I_25742 (I439794,I440146,I440050);
not I_25743 (I440168,I440146);
nor I_25744 (I440185,I440168,I439959);
nor I_25745 (I440202,I439891,I440185);
DFFARX1 I_25746 (I440202,I2507,I439826,I439809,);
nor I_25747 (I440233,I440168,I440050);
nor I_25748 (I440250,I884987,I885002);
nor I_25749 (I439800,I440250,I440233);
not I_25750 (I440281,I440250);
nand I_25751 (I439803,I440010,I440281);
DFFARX1 I_25752 (I440250,I2507,I439826,I439815,);
DFFARX1 I_25753 (I440250,I2507,I439826,I439812,);
not I_25754 (I440370,I2514);
DFFARX1 I_25755 (I283939,I2507,I440370,I440396,);
DFFARX1 I_25756 (I440396,I2507,I440370,I440413,);
not I_25757 (I440362,I440413);
not I_25758 (I440435,I440396);
nand I_25759 (I440452,I283918,I283942);
and I_25760 (I440469,I440452,I283945);
DFFARX1 I_25761 (I440469,I2507,I440370,I440495,);
not I_25762 (I440503,I440495);
DFFARX1 I_25763 (I283927,I2507,I440370,I440529,);
and I_25764 (I440537,I440529,I283933);
nand I_25765 (I440554,I440529,I283933);
nand I_25766 (I440341,I440503,I440554);
DFFARX1 I_25767 (I283921,I2507,I440370,I440594,);
nor I_25768 (I440602,I440594,I440537);
DFFARX1 I_25769 (I440602,I2507,I440370,I440335,);
nor I_25770 (I440350,I440594,I440495);
nand I_25771 (I440647,I283930,I283918);
and I_25772 (I440664,I440647,I283924);
DFFARX1 I_25773 (I440664,I2507,I440370,I440690,);
nor I_25774 (I440338,I440690,I440594);
not I_25775 (I440712,I440690);
nor I_25776 (I440729,I440712,I440503);
nor I_25777 (I440746,I440435,I440729);
DFFARX1 I_25778 (I440746,I2507,I440370,I440353,);
nor I_25779 (I440777,I440712,I440594);
nor I_25780 (I440794,I283936,I283918);
nor I_25781 (I440344,I440794,I440777);
not I_25782 (I440825,I440794);
nand I_25783 (I440347,I440554,I440825);
DFFARX1 I_25784 (I440794,I2507,I440370,I440359,);
DFFARX1 I_25785 (I440794,I2507,I440370,I440356,);
not I_25786 (I440914,I2514);
DFFARX1 I_25787 (I1177441,I2507,I440914,I440940,);
DFFARX1 I_25788 (I440940,I2507,I440914,I440957,);
not I_25789 (I440906,I440957);
not I_25790 (I440979,I440940);
nand I_25791 (I440996,I1177453,I1177441);
and I_25792 (I441013,I440996,I1177444);
DFFARX1 I_25793 (I441013,I2507,I440914,I441039,);
not I_25794 (I441047,I441039);
DFFARX1 I_25795 (I1177462,I2507,I440914,I441073,);
and I_25796 (I441081,I441073,I1177438);
nand I_25797 (I441098,I441073,I1177438);
nand I_25798 (I440885,I441047,I441098);
DFFARX1 I_25799 (I1177456,I2507,I440914,I441138,);
nor I_25800 (I441146,I441138,I441081);
DFFARX1 I_25801 (I441146,I2507,I440914,I440879,);
nor I_25802 (I440894,I441138,I441039);
nand I_25803 (I441191,I1177450,I1177447);
and I_25804 (I441208,I441191,I1177459);
DFFARX1 I_25805 (I441208,I2507,I440914,I441234,);
nor I_25806 (I440882,I441234,I441138);
not I_25807 (I441256,I441234);
nor I_25808 (I441273,I441256,I441047);
nor I_25809 (I441290,I440979,I441273);
DFFARX1 I_25810 (I441290,I2507,I440914,I440897,);
nor I_25811 (I441321,I441256,I441138);
nor I_25812 (I441338,I1177438,I1177447);
nor I_25813 (I440888,I441338,I441321);
not I_25814 (I441369,I441338);
nand I_25815 (I440891,I441098,I441369);
DFFARX1 I_25816 (I441338,I2507,I440914,I440903,);
DFFARX1 I_25817 (I441338,I2507,I440914,I440900,);
not I_25818 (I441458,I2514);
DFFARX1 I_25819 (I755569,I2507,I441458,I441484,);
DFFARX1 I_25820 (I441484,I2507,I441458,I441501,);
not I_25821 (I441450,I441501);
not I_25822 (I441523,I441484);
nand I_25823 (I441540,I755590,I755581);
and I_25824 (I441557,I441540,I755569);
DFFARX1 I_25825 (I441557,I2507,I441458,I441583,);
not I_25826 (I441591,I441583);
DFFARX1 I_25827 (I755575,I2507,I441458,I441617,);
and I_25828 (I441625,I441617,I755572);
nand I_25829 (I441642,I441617,I755572);
nand I_25830 (I441429,I441591,I441642);
DFFARX1 I_25831 (I755566,I2507,I441458,I441682,);
nor I_25832 (I441690,I441682,I441625);
DFFARX1 I_25833 (I441690,I2507,I441458,I441423,);
nor I_25834 (I441438,I441682,I441583);
nand I_25835 (I441735,I755566,I755578);
and I_25836 (I441752,I441735,I755587);
DFFARX1 I_25837 (I441752,I2507,I441458,I441778,);
nor I_25838 (I441426,I441778,I441682);
not I_25839 (I441800,I441778);
nor I_25840 (I441817,I441800,I441591);
nor I_25841 (I441834,I441523,I441817);
DFFARX1 I_25842 (I441834,I2507,I441458,I441441,);
nor I_25843 (I441865,I441800,I441682);
nor I_25844 (I441882,I755584,I755578);
nor I_25845 (I441432,I441882,I441865);
not I_25846 (I441913,I441882);
nand I_25847 (I441435,I441642,I441913);
DFFARX1 I_25848 (I441882,I2507,I441458,I441447,);
DFFARX1 I_25849 (I441882,I2507,I441458,I441444,);
not I_25850 (I442002,I2514);
DFFARX1 I_25851 (I1166459,I2507,I442002,I442028,);
DFFARX1 I_25852 (I442028,I2507,I442002,I442045,);
not I_25853 (I441994,I442045);
not I_25854 (I442067,I442028);
nand I_25855 (I442084,I1166471,I1166459);
and I_25856 (I442101,I442084,I1166462);
DFFARX1 I_25857 (I442101,I2507,I442002,I442127,);
not I_25858 (I442135,I442127);
DFFARX1 I_25859 (I1166480,I2507,I442002,I442161,);
and I_25860 (I442169,I442161,I1166456);
nand I_25861 (I442186,I442161,I1166456);
nand I_25862 (I441973,I442135,I442186);
DFFARX1 I_25863 (I1166474,I2507,I442002,I442226,);
nor I_25864 (I442234,I442226,I442169);
DFFARX1 I_25865 (I442234,I2507,I442002,I441967,);
nor I_25866 (I441982,I442226,I442127);
nand I_25867 (I442279,I1166468,I1166465);
and I_25868 (I442296,I442279,I1166477);
DFFARX1 I_25869 (I442296,I2507,I442002,I442322,);
nor I_25870 (I441970,I442322,I442226);
not I_25871 (I442344,I442322);
nor I_25872 (I442361,I442344,I442135);
nor I_25873 (I442378,I442067,I442361);
DFFARX1 I_25874 (I442378,I2507,I442002,I441985,);
nor I_25875 (I442409,I442344,I442226);
nor I_25876 (I442426,I1166456,I1166465);
nor I_25877 (I441976,I442426,I442409);
not I_25878 (I442457,I442426);
nand I_25879 (I441979,I442186,I442457);
DFFARX1 I_25880 (I442426,I2507,I442002,I441991,);
DFFARX1 I_25881 (I442426,I2507,I442002,I441988,);
not I_25882 (I442546,I2514);
DFFARX1 I_25883 (I650951,I2507,I442546,I442572,);
DFFARX1 I_25884 (I442572,I2507,I442546,I442589,);
not I_25885 (I442538,I442589);
not I_25886 (I442611,I442572);
nand I_25887 (I442628,I650972,I650963);
and I_25888 (I442645,I442628,I650951);
DFFARX1 I_25889 (I442645,I2507,I442546,I442671,);
not I_25890 (I442679,I442671);
DFFARX1 I_25891 (I650957,I2507,I442546,I442705,);
and I_25892 (I442713,I442705,I650954);
nand I_25893 (I442730,I442705,I650954);
nand I_25894 (I442517,I442679,I442730);
DFFARX1 I_25895 (I650948,I2507,I442546,I442770,);
nor I_25896 (I442778,I442770,I442713);
DFFARX1 I_25897 (I442778,I2507,I442546,I442511,);
nor I_25898 (I442526,I442770,I442671);
nand I_25899 (I442823,I650948,I650960);
and I_25900 (I442840,I442823,I650969);
DFFARX1 I_25901 (I442840,I2507,I442546,I442866,);
nor I_25902 (I442514,I442866,I442770);
not I_25903 (I442888,I442866);
nor I_25904 (I442905,I442888,I442679);
nor I_25905 (I442922,I442611,I442905);
DFFARX1 I_25906 (I442922,I2507,I442546,I442529,);
nor I_25907 (I442953,I442888,I442770);
nor I_25908 (I442970,I650966,I650960);
nor I_25909 (I442520,I442970,I442953);
not I_25910 (I443001,I442970);
nand I_25911 (I442523,I442730,I443001);
DFFARX1 I_25912 (I442970,I2507,I442546,I442535,);
DFFARX1 I_25913 (I442970,I2507,I442546,I442532,);
not I_25914 (I443090,I2514);
DFFARX1 I_25915 (I899851,I2507,I443090,I443116,);
DFFARX1 I_25916 (I443116,I2507,I443090,I443133,);
not I_25917 (I443082,I443133);
not I_25918 (I443155,I443116);
nand I_25919 (I443172,I899866,I899854);
and I_25920 (I443189,I443172,I899845);
DFFARX1 I_25921 (I443189,I2507,I443090,I443215,);
not I_25922 (I443223,I443215);
DFFARX1 I_25923 (I899857,I2507,I443090,I443249,);
and I_25924 (I443257,I443249,I899848);
nand I_25925 (I443274,I443249,I899848);
nand I_25926 (I443061,I443223,I443274);
DFFARX1 I_25927 (I899863,I2507,I443090,I443314,);
nor I_25928 (I443322,I443314,I443257);
DFFARX1 I_25929 (I443322,I2507,I443090,I443055,);
nor I_25930 (I443070,I443314,I443215);
nand I_25931 (I443367,I899872,I899860);
and I_25932 (I443384,I443367,I899869);
DFFARX1 I_25933 (I443384,I2507,I443090,I443410,);
nor I_25934 (I443058,I443410,I443314);
not I_25935 (I443432,I443410);
nor I_25936 (I443449,I443432,I443223);
nor I_25937 (I443466,I443155,I443449);
DFFARX1 I_25938 (I443466,I2507,I443090,I443073,);
nor I_25939 (I443497,I443432,I443314);
nor I_25940 (I443514,I899845,I899860);
nor I_25941 (I443064,I443514,I443497);
not I_25942 (I443545,I443514);
nand I_25943 (I443067,I443274,I443545);
DFFARX1 I_25944 (I443514,I2507,I443090,I443079,);
DFFARX1 I_25945 (I443514,I2507,I443090,I443076,);
not I_25946 (I443634,I2514);
DFFARX1 I_25947 (I707017,I2507,I443634,I443660,);
DFFARX1 I_25948 (I443660,I2507,I443634,I443677,);
not I_25949 (I443626,I443677);
not I_25950 (I443699,I443660);
nand I_25951 (I443716,I707038,I707029);
and I_25952 (I443733,I443716,I707017);
DFFARX1 I_25953 (I443733,I2507,I443634,I443759,);
not I_25954 (I443767,I443759);
DFFARX1 I_25955 (I707023,I2507,I443634,I443793,);
and I_25956 (I443801,I443793,I707020);
nand I_25957 (I443818,I443793,I707020);
nand I_25958 (I443605,I443767,I443818);
DFFARX1 I_25959 (I707014,I2507,I443634,I443858,);
nor I_25960 (I443866,I443858,I443801);
DFFARX1 I_25961 (I443866,I2507,I443634,I443599,);
nor I_25962 (I443614,I443858,I443759);
nand I_25963 (I443911,I707014,I707026);
and I_25964 (I443928,I443911,I707035);
DFFARX1 I_25965 (I443928,I2507,I443634,I443954,);
nor I_25966 (I443602,I443954,I443858);
not I_25967 (I443976,I443954);
nor I_25968 (I443993,I443976,I443767);
nor I_25969 (I444010,I443699,I443993);
DFFARX1 I_25970 (I444010,I2507,I443634,I443617,);
nor I_25971 (I444041,I443976,I443858);
nor I_25972 (I444058,I707032,I707026);
nor I_25973 (I443608,I444058,I444041);
not I_25974 (I444089,I444058);
nand I_25975 (I443611,I443818,I444089);
DFFARX1 I_25976 (I444058,I2507,I443634,I443623,);
DFFARX1 I_25977 (I444058,I2507,I443634,I443620,);
not I_25978 (I444178,I2514);
DFFARX1 I_25979 (I162734,I2507,I444178,I444204,);
DFFARX1 I_25980 (I444204,I2507,I444178,I444221,);
not I_25981 (I444170,I444221);
not I_25982 (I444243,I444204);
nand I_25983 (I444260,I162746,I162725);
and I_25984 (I444277,I444260,I162728);
DFFARX1 I_25985 (I444277,I2507,I444178,I444303,);
not I_25986 (I444311,I444303);
DFFARX1 I_25987 (I162737,I2507,I444178,I444337,);
and I_25988 (I444345,I444337,I162749);
nand I_25989 (I444362,I444337,I162749);
nand I_25990 (I444149,I444311,I444362);
DFFARX1 I_25991 (I162743,I2507,I444178,I444402,);
nor I_25992 (I444410,I444402,I444345);
DFFARX1 I_25993 (I444410,I2507,I444178,I444143,);
nor I_25994 (I444158,I444402,I444303);
nand I_25995 (I444455,I162731,I162728);
and I_25996 (I444472,I444455,I162740);
DFFARX1 I_25997 (I444472,I2507,I444178,I444498,);
nor I_25998 (I444146,I444498,I444402);
not I_25999 (I444520,I444498);
nor I_26000 (I444537,I444520,I444311);
nor I_26001 (I444554,I444243,I444537);
DFFARX1 I_26002 (I444554,I2507,I444178,I444161,);
nor I_26003 (I444585,I444520,I444402);
nor I_26004 (I444602,I162725,I162728);
nor I_26005 (I444152,I444602,I444585);
not I_26006 (I444633,I444602);
nand I_26007 (I444155,I444362,I444633);
DFFARX1 I_26008 (I444602,I2507,I444178,I444167,);
DFFARX1 I_26009 (I444602,I2507,I444178,I444164,);
not I_26010 (I444722,I2514);
DFFARX1 I_26011 (I1242789,I2507,I444722,I444748,);
DFFARX1 I_26012 (I444748,I2507,I444722,I444765,);
not I_26013 (I444714,I444765);
not I_26014 (I444787,I444748);
nand I_26015 (I444804,I1242801,I1242804);
and I_26016 (I444821,I444804,I1242807);
DFFARX1 I_26017 (I444821,I2507,I444722,I444847,);
not I_26018 (I444855,I444847);
DFFARX1 I_26019 (I1242792,I2507,I444722,I444881,);
and I_26020 (I444889,I444881,I1242798);
nand I_26021 (I444906,I444881,I1242798);
nand I_26022 (I444693,I444855,I444906);
DFFARX1 I_26023 (I1242786,I2507,I444722,I444946,);
nor I_26024 (I444954,I444946,I444889);
DFFARX1 I_26025 (I444954,I2507,I444722,I444687,);
nor I_26026 (I444702,I444946,I444847);
nand I_26027 (I444999,I1242789,I1242810);
and I_26028 (I445016,I444999,I1242795);
DFFARX1 I_26029 (I445016,I2507,I444722,I445042,);
nor I_26030 (I444690,I445042,I444946);
not I_26031 (I445064,I445042);
nor I_26032 (I445081,I445064,I444855);
nor I_26033 (I445098,I444787,I445081);
DFFARX1 I_26034 (I445098,I2507,I444722,I444705,);
nor I_26035 (I445129,I445064,I444946);
nor I_26036 (I445146,I1242786,I1242810);
nor I_26037 (I444696,I445146,I445129);
not I_26038 (I445177,I445146);
nand I_26039 (I444699,I444906,I445177);
DFFARX1 I_26040 (I445146,I2507,I444722,I444711,);
DFFARX1 I_26041 (I445146,I2507,I444722,I444708,);
not I_26042 (I445266,I2514);
DFFARX1 I_26043 (I851271,I2507,I445266,I445292,);
DFFARX1 I_26044 (I445292,I2507,I445266,I445309,);
not I_26045 (I445258,I445309);
not I_26046 (I445331,I445292);
nand I_26047 (I445348,I851265,I851262);
and I_26048 (I445365,I445348,I851277);
DFFARX1 I_26049 (I445365,I2507,I445266,I445391,);
not I_26050 (I445399,I445391);
DFFARX1 I_26051 (I851265,I2507,I445266,I445425,);
and I_26052 (I445433,I445425,I851259);
nand I_26053 (I445450,I445425,I851259);
nand I_26054 (I445237,I445399,I445450);
DFFARX1 I_26055 (I851259,I2507,I445266,I445490,);
nor I_26056 (I445498,I445490,I445433);
DFFARX1 I_26057 (I445498,I2507,I445266,I445231,);
nor I_26058 (I445246,I445490,I445391);
nand I_26059 (I445543,I851274,I851268);
and I_26060 (I445560,I445543,I851262);
DFFARX1 I_26061 (I445560,I2507,I445266,I445586,);
nor I_26062 (I445234,I445586,I445490);
not I_26063 (I445608,I445586);
nor I_26064 (I445625,I445608,I445399);
nor I_26065 (I445642,I445331,I445625);
DFFARX1 I_26066 (I445642,I2507,I445266,I445249,);
nor I_26067 (I445673,I445608,I445490);
nor I_26068 (I445690,I851280,I851268);
nor I_26069 (I445240,I445690,I445673);
not I_26070 (I445721,I445690);
nand I_26071 (I445243,I445450,I445721);
DFFARX1 I_26072 (I445690,I2507,I445266,I445255,);
DFFARX1 I_26073 (I445690,I2507,I445266,I445252,);
not I_26074 (I445810,I2514);
DFFARX1 I_26075 (I734183,I2507,I445810,I445836,);
DFFARX1 I_26076 (I445836,I2507,I445810,I445853,);
not I_26077 (I445802,I445853);
not I_26078 (I445875,I445836);
nand I_26079 (I445892,I734204,I734195);
and I_26080 (I445909,I445892,I734183);
DFFARX1 I_26081 (I445909,I2507,I445810,I445935,);
not I_26082 (I445943,I445935);
DFFARX1 I_26083 (I734189,I2507,I445810,I445969,);
and I_26084 (I445977,I445969,I734186);
nand I_26085 (I445994,I445969,I734186);
nand I_26086 (I445781,I445943,I445994);
DFFARX1 I_26087 (I734180,I2507,I445810,I446034,);
nor I_26088 (I446042,I446034,I445977);
DFFARX1 I_26089 (I446042,I2507,I445810,I445775,);
nor I_26090 (I445790,I446034,I445935);
nand I_26091 (I446087,I734180,I734192);
and I_26092 (I446104,I446087,I734201);
DFFARX1 I_26093 (I446104,I2507,I445810,I446130,);
nor I_26094 (I445778,I446130,I446034);
not I_26095 (I446152,I446130);
nor I_26096 (I446169,I446152,I445943);
nor I_26097 (I446186,I445875,I446169);
DFFARX1 I_26098 (I446186,I2507,I445810,I445793,);
nor I_26099 (I446217,I446152,I446034);
nor I_26100 (I446234,I734198,I734192);
nor I_26101 (I445784,I446234,I446217);
not I_26102 (I446265,I446234);
nand I_26103 (I445787,I445994,I446265);
DFFARX1 I_26104 (I446234,I2507,I445810,I445799,);
DFFARX1 I_26105 (I446234,I2507,I445810,I445796,);
not I_26106 (I446354,I2514);
DFFARX1 I_26107 (I237704,I2507,I446354,I446380,);
DFFARX1 I_26108 (I446380,I2507,I446354,I446397,);
not I_26109 (I446346,I446397);
not I_26110 (I446419,I446380);
nand I_26111 (I446436,I237716,I237695);
and I_26112 (I446453,I446436,I237698);
DFFARX1 I_26113 (I446453,I2507,I446354,I446479,);
not I_26114 (I446487,I446479);
DFFARX1 I_26115 (I237707,I2507,I446354,I446513,);
and I_26116 (I446521,I446513,I237719);
nand I_26117 (I446538,I446513,I237719);
nand I_26118 (I446325,I446487,I446538);
DFFARX1 I_26119 (I237713,I2507,I446354,I446578,);
nor I_26120 (I446586,I446578,I446521);
DFFARX1 I_26121 (I446586,I2507,I446354,I446319,);
nor I_26122 (I446334,I446578,I446479);
nand I_26123 (I446631,I237701,I237698);
and I_26124 (I446648,I446631,I237710);
DFFARX1 I_26125 (I446648,I2507,I446354,I446674,);
nor I_26126 (I446322,I446674,I446578);
not I_26127 (I446696,I446674);
nor I_26128 (I446713,I446696,I446487);
nor I_26129 (I446730,I446419,I446713);
DFFARX1 I_26130 (I446730,I2507,I446354,I446337,);
nor I_26131 (I446761,I446696,I446578);
nor I_26132 (I446778,I237695,I237698);
nor I_26133 (I446328,I446778,I446761);
not I_26134 (I446809,I446778);
nand I_26135 (I446331,I446538,I446809);
DFFARX1 I_26136 (I446778,I2507,I446354,I446343,);
DFFARX1 I_26137 (I446778,I2507,I446354,I446340,);
not I_26138 (I446898,I2514);
DFFARX1 I_26139 (I564251,I2507,I446898,I446924,);
DFFARX1 I_26140 (I446924,I2507,I446898,I446941,);
not I_26141 (I446890,I446941);
not I_26142 (I446963,I446924);
nand I_26143 (I446980,I564248,I564269);
and I_26144 (I446997,I446980,I564272);
DFFARX1 I_26145 (I446997,I2507,I446898,I447023,);
not I_26146 (I447031,I447023);
DFFARX1 I_26147 (I564257,I2507,I446898,I447057,);
and I_26148 (I447065,I447057,I564260);
nand I_26149 (I447082,I447057,I564260);
nand I_26150 (I446869,I447031,I447082);
DFFARX1 I_26151 (I564263,I2507,I446898,I447122,);
nor I_26152 (I447130,I447122,I447065);
DFFARX1 I_26153 (I447130,I2507,I446898,I446863,);
nor I_26154 (I446878,I447122,I447023);
nand I_26155 (I447175,I564248,I564254);
and I_26156 (I447192,I447175,I564266);
DFFARX1 I_26157 (I447192,I2507,I446898,I447218,);
nor I_26158 (I446866,I447218,I447122);
not I_26159 (I447240,I447218);
nor I_26160 (I447257,I447240,I447031);
nor I_26161 (I447274,I446963,I447257);
DFFARX1 I_26162 (I447274,I2507,I446898,I446881,);
nor I_26163 (I447305,I447240,I447122);
nor I_26164 (I447322,I564251,I564254);
nor I_26165 (I446872,I447322,I447305);
not I_26166 (I447353,I447322);
nand I_26167 (I446875,I447082,I447353);
DFFARX1 I_26168 (I447322,I2507,I446898,I446887,);
DFFARX1 I_26169 (I447322,I2507,I446898,I446884,);
not I_26170 (I447442,I2514);
DFFARX1 I_26171 (I810165,I2507,I447442,I447468,);
DFFARX1 I_26172 (I447468,I2507,I447442,I447485,);
not I_26173 (I447434,I447485);
not I_26174 (I447507,I447468);
nand I_26175 (I447524,I810159,I810156);
and I_26176 (I447541,I447524,I810171);
DFFARX1 I_26177 (I447541,I2507,I447442,I447567,);
not I_26178 (I447575,I447567);
DFFARX1 I_26179 (I810159,I2507,I447442,I447601,);
and I_26180 (I447609,I447601,I810153);
nand I_26181 (I447626,I447601,I810153);
nand I_26182 (I447413,I447575,I447626);
DFFARX1 I_26183 (I810153,I2507,I447442,I447666,);
nor I_26184 (I447674,I447666,I447609);
DFFARX1 I_26185 (I447674,I2507,I447442,I447407,);
nor I_26186 (I447422,I447666,I447567);
nand I_26187 (I447719,I810168,I810162);
and I_26188 (I447736,I447719,I810156);
DFFARX1 I_26189 (I447736,I2507,I447442,I447762,);
nor I_26190 (I447410,I447762,I447666);
not I_26191 (I447784,I447762);
nor I_26192 (I447801,I447784,I447575);
nor I_26193 (I447818,I447507,I447801);
DFFARX1 I_26194 (I447818,I2507,I447442,I447425,);
nor I_26195 (I447849,I447784,I447666);
nor I_26196 (I447866,I810174,I810162);
nor I_26197 (I447416,I447866,I447849);
not I_26198 (I447897,I447866);
nand I_26199 (I447419,I447626,I447897);
DFFARX1 I_26200 (I447866,I2507,I447442,I447431,);
DFFARX1 I_26201 (I447866,I2507,I447442,I447428,);
not I_26202 (I447986,I2514);
DFFARX1 I_26203 (I921815,I2507,I447986,I448012,);
DFFARX1 I_26204 (I448012,I2507,I447986,I448029,);
not I_26205 (I447978,I448029);
not I_26206 (I448051,I448012);
nand I_26207 (I448068,I921830,I921818);
and I_26208 (I448085,I448068,I921809);
DFFARX1 I_26209 (I448085,I2507,I447986,I448111,);
not I_26210 (I448119,I448111);
DFFARX1 I_26211 (I921821,I2507,I447986,I448145,);
and I_26212 (I448153,I448145,I921812);
nand I_26213 (I448170,I448145,I921812);
nand I_26214 (I447957,I448119,I448170);
DFFARX1 I_26215 (I921827,I2507,I447986,I448210,);
nor I_26216 (I448218,I448210,I448153);
DFFARX1 I_26217 (I448218,I2507,I447986,I447951,);
nor I_26218 (I447966,I448210,I448111);
nand I_26219 (I448263,I921836,I921824);
and I_26220 (I448280,I448263,I921833);
DFFARX1 I_26221 (I448280,I2507,I447986,I448306,);
nor I_26222 (I447954,I448306,I448210);
not I_26223 (I448328,I448306);
nor I_26224 (I448345,I448328,I448119);
nor I_26225 (I448362,I448051,I448345);
DFFARX1 I_26226 (I448362,I2507,I447986,I447969,);
nor I_26227 (I448393,I448328,I448210);
nor I_26228 (I448410,I921809,I921824);
nor I_26229 (I447960,I448410,I448393);
not I_26230 (I448441,I448410);
nand I_26231 (I447963,I448170,I448441);
DFFARX1 I_26232 (I448410,I2507,I447986,I447975,);
DFFARX1 I_26233 (I448410,I2507,I447986,I447972,);
not I_26234 (I448530,I2514);
DFFARX1 I_26235 (I525627,I2507,I448530,I448556,);
DFFARX1 I_26236 (I448556,I2507,I448530,I448573,);
not I_26237 (I448522,I448573);
not I_26238 (I448595,I448556);
nand I_26239 (I448612,I525630,I525648);
and I_26240 (I448629,I448612,I525636);
DFFARX1 I_26241 (I448629,I2507,I448530,I448655,);
not I_26242 (I448663,I448655);
DFFARX1 I_26243 (I525627,I2507,I448530,I448689,);
and I_26244 (I448697,I448689,I525645);
nand I_26245 (I448714,I448689,I525645);
nand I_26246 (I448501,I448663,I448714);
DFFARX1 I_26247 (I525639,I2507,I448530,I448754,);
nor I_26248 (I448762,I448754,I448697);
DFFARX1 I_26249 (I448762,I2507,I448530,I448495,);
nor I_26250 (I448510,I448754,I448655);
nand I_26251 (I448807,I525642,I525624);
and I_26252 (I448824,I448807,I525633);
DFFARX1 I_26253 (I448824,I2507,I448530,I448850,);
nor I_26254 (I448498,I448850,I448754);
not I_26255 (I448872,I448850);
nor I_26256 (I448889,I448872,I448663);
nor I_26257 (I448906,I448595,I448889);
DFFARX1 I_26258 (I448906,I2507,I448530,I448513,);
nor I_26259 (I448937,I448872,I448754);
nor I_26260 (I448954,I525624,I525624);
nor I_26261 (I448504,I448954,I448937);
not I_26262 (I448985,I448954);
nand I_26263 (I448507,I448714,I448985);
DFFARX1 I_26264 (I448954,I2507,I448530,I448519,);
DFFARX1 I_26265 (I448954,I2507,I448530,I448516,);
not I_26266 (I449074,I2514);
DFFARX1 I_26267 (I168684,I2507,I449074,I449100,);
DFFARX1 I_26268 (I449100,I2507,I449074,I449117,);
not I_26269 (I449066,I449117);
not I_26270 (I449139,I449100);
nand I_26271 (I449156,I168696,I168675);
and I_26272 (I449173,I449156,I168678);
DFFARX1 I_26273 (I449173,I2507,I449074,I449199,);
not I_26274 (I449207,I449199);
DFFARX1 I_26275 (I168687,I2507,I449074,I449233,);
and I_26276 (I449241,I449233,I168699);
nand I_26277 (I449258,I449233,I168699);
nand I_26278 (I449045,I449207,I449258);
DFFARX1 I_26279 (I168693,I2507,I449074,I449298,);
nor I_26280 (I449306,I449298,I449241);
DFFARX1 I_26281 (I449306,I2507,I449074,I449039,);
nor I_26282 (I449054,I449298,I449199);
nand I_26283 (I449351,I168681,I168678);
and I_26284 (I449368,I449351,I168690);
DFFARX1 I_26285 (I449368,I2507,I449074,I449394,);
nor I_26286 (I449042,I449394,I449298);
not I_26287 (I449416,I449394);
nor I_26288 (I449433,I449416,I449207);
nor I_26289 (I449450,I449139,I449433);
DFFARX1 I_26290 (I449450,I2507,I449074,I449057,);
nor I_26291 (I449481,I449416,I449298);
nor I_26292 (I449498,I168675,I168678);
nor I_26293 (I449048,I449498,I449481);
not I_26294 (I449529,I449498);
nand I_26295 (I449051,I449258,I449529);
DFFARX1 I_26296 (I449498,I2507,I449074,I449063,);
DFFARX1 I_26297 (I449498,I2507,I449074,I449060,);
not I_26298 (I449618,I2514);
DFFARX1 I_26299 (I946363,I2507,I449618,I449644,);
DFFARX1 I_26300 (I449644,I2507,I449618,I449661,);
not I_26301 (I449610,I449661);
not I_26302 (I449683,I449644);
nand I_26303 (I449700,I946378,I946366);
and I_26304 (I449717,I449700,I946357);
DFFARX1 I_26305 (I449717,I2507,I449618,I449743,);
not I_26306 (I449751,I449743);
DFFARX1 I_26307 (I946369,I2507,I449618,I449777,);
and I_26308 (I449785,I449777,I946360);
nand I_26309 (I449802,I449777,I946360);
nand I_26310 (I449589,I449751,I449802);
DFFARX1 I_26311 (I946375,I2507,I449618,I449842,);
nor I_26312 (I449850,I449842,I449785);
DFFARX1 I_26313 (I449850,I2507,I449618,I449583,);
nor I_26314 (I449598,I449842,I449743);
nand I_26315 (I449895,I946384,I946372);
and I_26316 (I449912,I449895,I946381);
DFFARX1 I_26317 (I449912,I2507,I449618,I449938,);
nor I_26318 (I449586,I449938,I449842);
not I_26319 (I449960,I449938);
nor I_26320 (I449977,I449960,I449751);
nor I_26321 (I449994,I449683,I449977);
DFFARX1 I_26322 (I449994,I2507,I449618,I449601,);
nor I_26323 (I450025,I449960,I449842);
nor I_26324 (I450042,I946357,I946372);
nor I_26325 (I449592,I450042,I450025);
not I_26326 (I450073,I450042);
nand I_26327 (I449595,I449802,I450073);
DFFARX1 I_26328 (I450042,I2507,I449618,I449607,);
DFFARX1 I_26329 (I450042,I2507,I449618,I449604,);
not I_26330 (I450162,I2514);
DFFARX1 I_26331 (I720311,I2507,I450162,I450188,);
DFFARX1 I_26332 (I450188,I2507,I450162,I450205,);
not I_26333 (I450154,I450205);
not I_26334 (I450227,I450188);
nand I_26335 (I450244,I720332,I720323);
and I_26336 (I450261,I450244,I720311);
DFFARX1 I_26337 (I450261,I2507,I450162,I450287,);
not I_26338 (I450295,I450287);
DFFARX1 I_26339 (I720317,I2507,I450162,I450321,);
and I_26340 (I450329,I450321,I720314);
nand I_26341 (I450346,I450321,I720314);
nand I_26342 (I450133,I450295,I450346);
DFFARX1 I_26343 (I720308,I2507,I450162,I450386,);
nor I_26344 (I450394,I450386,I450329);
DFFARX1 I_26345 (I450394,I2507,I450162,I450127,);
nor I_26346 (I450142,I450386,I450287);
nand I_26347 (I450439,I720308,I720320);
and I_26348 (I450456,I450439,I720329);
DFFARX1 I_26349 (I450456,I2507,I450162,I450482,);
nor I_26350 (I450130,I450482,I450386);
not I_26351 (I450504,I450482);
nor I_26352 (I450521,I450504,I450295);
nor I_26353 (I450538,I450227,I450521);
DFFARX1 I_26354 (I450538,I2507,I450162,I450145,);
nor I_26355 (I450569,I450504,I450386);
nor I_26356 (I450586,I720326,I720320);
nor I_26357 (I450136,I450586,I450569);
not I_26358 (I450617,I450586);
nand I_26359 (I450139,I450346,I450617);
DFFARX1 I_26360 (I450586,I2507,I450162,I450151,);
DFFARX1 I_26361 (I450586,I2507,I450162,I450148,);
not I_26362 (I450706,I2514);
DFFARX1 I_26363 (I744009,I2507,I450706,I450732,);
DFFARX1 I_26364 (I450732,I2507,I450706,I450749,);
not I_26365 (I450698,I450749);
not I_26366 (I450771,I450732);
nand I_26367 (I450788,I744030,I744021);
and I_26368 (I450805,I450788,I744009);
DFFARX1 I_26369 (I450805,I2507,I450706,I450831,);
not I_26370 (I450839,I450831);
DFFARX1 I_26371 (I744015,I2507,I450706,I450865,);
and I_26372 (I450873,I450865,I744012);
nand I_26373 (I450890,I450865,I744012);
nand I_26374 (I450677,I450839,I450890);
DFFARX1 I_26375 (I744006,I2507,I450706,I450930,);
nor I_26376 (I450938,I450930,I450873);
DFFARX1 I_26377 (I450938,I2507,I450706,I450671,);
nor I_26378 (I450686,I450930,I450831);
nand I_26379 (I450983,I744006,I744018);
and I_26380 (I451000,I450983,I744027);
DFFARX1 I_26381 (I451000,I2507,I450706,I451026,);
nor I_26382 (I450674,I451026,I450930);
not I_26383 (I451048,I451026);
nor I_26384 (I451065,I451048,I450839);
nor I_26385 (I451082,I450771,I451065);
DFFARX1 I_26386 (I451082,I2507,I450706,I450689,);
nor I_26387 (I451113,I451048,I450930);
nor I_26388 (I451130,I744024,I744018);
nor I_26389 (I450680,I451130,I451113);
not I_26390 (I451161,I451130);
nand I_26391 (I450683,I450890,I451161);
DFFARX1 I_26392 (I451130,I2507,I450706,I450695,);
DFFARX1 I_26393 (I451130,I2507,I450706,I450692,);
not I_26394 (I451250,I2514);
DFFARX1 I_26395 (I922461,I2507,I451250,I451276,);
DFFARX1 I_26396 (I451276,I2507,I451250,I451293,);
not I_26397 (I451242,I451293);
not I_26398 (I451315,I451276);
nand I_26399 (I451332,I922476,I922464);
and I_26400 (I451349,I451332,I922455);
DFFARX1 I_26401 (I451349,I2507,I451250,I451375,);
not I_26402 (I451383,I451375);
DFFARX1 I_26403 (I922467,I2507,I451250,I451409,);
and I_26404 (I451417,I451409,I922458);
nand I_26405 (I451434,I451409,I922458);
nand I_26406 (I451221,I451383,I451434);
DFFARX1 I_26407 (I922473,I2507,I451250,I451474,);
nor I_26408 (I451482,I451474,I451417);
DFFARX1 I_26409 (I451482,I2507,I451250,I451215,);
nor I_26410 (I451230,I451474,I451375);
nand I_26411 (I451527,I922482,I922470);
and I_26412 (I451544,I451527,I922479);
DFFARX1 I_26413 (I451544,I2507,I451250,I451570,);
nor I_26414 (I451218,I451570,I451474);
not I_26415 (I451592,I451570);
nor I_26416 (I451609,I451592,I451383);
nor I_26417 (I451626,I451315,I451609);
DFFARX1 I_26418 (I451626,I2507,I451250,I451233,);
nor I_26419 (I451657,I451592,I451474);
nor I_26420 (I451674,I922455,I922470);
nor I_26421 (I451224,I451674,I451657);
not I_26422 (I451705,I451674);
nand I_26423 (I451227,I451434,I451705);
DFFARX1 I_26424 (I451674,I2507,I451250,I451239,);
DFFARX1 I_26425 (I451674,I2507,I451250,I451236,);
not I_26426 (I451794,I2514);
DFFARX1 I_26427 (I1241157,I2507,I451794,I451820,);
DFFARX1 I_26428 (I451820,I2507,I451794,I451837,);
not I_26429 (I451786,I451837);
not I_26430 (I451859,I451820);
nand I_26431 (I451876,I1241169,I1241172);
and I_26432 (I451893,I451876,I1241175);
DFFARX1 I_26433 (I451893,I2507,I451794,I451919,);
not I_26434 (I451927,I451919);
DFFARX1 I_26435 (I1241160,I2507,I451794,I451953,);
and I_26436 (I451961,I451953,I1241166);
nand I_26437 (I451978,I451953,I1241166);
nand I_26438 (I451765,I451927,I451978);
DFFARX1 I_26439 (I1241154,I2507,I451794,I452018,);
nor I_26440 (I452026,I452018,I451961);
DFFARX1 I_26441 (I452026,I2507,I451794,I451759,);
nor I_26442 (I451774,I452018,I451919);
nand I_26443 (I452071,I1241157,I1241178);
and I_26444 (I452088,I452071,I1241163);
DFFARX1 I_26445 (I452088,I2507,I451794,I452114,);
nor I_26446 (I451762,I452114,I452018);
not I_26447 (I452136,I452114);
nor I_26448 (I452153,I452136,I451927);
nor I_26449 (I452170,I451859,I452153);
DFFARX1 I_26450 (I452170,I2507,I451794,I451777,);
nor I_26451 (I452201,I452136,I452018);
nor I_26452 (I452218,I1241154,I1241178);
nor I_26453 (I451768,I452218,I452201);
not I_26454 (I452249,I452218);
nand I_26455 (I451771,I451978,I452249);
DFFARX1 I_26456 (I452218,I2507,I451794,I451783,);
DFFARX1 I_26457 (I452218,I2507,I451794,I451780,);
not I_26458 (I452338,I2514);
DFFARX1 I_26459 (I1116751,I2507,I452338,I452364,);
DFFARX1 I_26460 (I452364,I2507,I452338,I452381,);
not I_26461 (I452330,I452381);
not I_26462 (I452403,I452364);
nand I_26463 (I452420,I1116763,I1116751);
and I_26464 (I452437,I452420,I1116754);
DFFARX1 I_26465 (I452437,I2507,I452338,I452463,);
not I_26466 (I452471,I452463);
DFFARX1 I_26467 (I1116772,I2507,I452338,I452497,);
and I_26468 (I452505,I452497,I1116748);
nand I_26469 (I452522,I452497,I1116748);
nand I_26470 (I452309,I452471,I452522);
DFFARX1 I_26471 (I1116766,I2507,I452338,I452562,);
nor I_26472 (I452570,I452562,I452505);
DFFARX1 I_26473 (I452570,I2507,I452338,I452303,);
nor I_26474 (I452318,I452562,I452463);
nand I_26475 (I452615,I1116760,I1116757);
and I_26476 (I452632,I452615,I1116769);
DFFARX1 I_26477 (I452632,I2507,I452338,I452658,);
nor I_26478 (I452306,I452658,I452562);
not I_26479 (I452680,I452658);
nor I_26480 (I452697,I452680,I452471);
nor I_26481 (I452714,I452403,I452697);
DFFARX1 I_26482 (I452714,I2507,I452338,I452321,);
nor I_26483 (I452745,I452680,I452562);
nor I_26484 (I452762,I1116748,I1116757);
nor I_26485 (I452312,I452762,I452745);
not I_26486 (I452793,I452762);
nand I_26487 (I452315,I452522,I452793);
DFFARX1 I_26488 (I452762,I2507,I452338,I452327,);
DFFARX1 I_26489 (I452762,I2507,I452338,I452324,);
not I_26490 (I452882,I2514);
DFFARX1 I_26491 (I347179,I2507,I452882,I452908,);
DFFARX1 I_26492 (I452908,I2507,I452882,I452925,);
not I_26493 (I452874,I452925);
not I_26494 (I452947,I452908);
nand I_26495 (I452964,I347158,I347182);
and I_26496 (I452981,I452964,I347185);
DFFARX1 I_26497 (I452981,I2507,I452882,I453007,);
not I_26498 (I453015,I453007);
DFFARX1 I_26499 (I347167,I2507,I452882,I453041,);
and I_26500 (I453049,I453041,I347173);
nand I_26501 (I453066,I453041,I347173);
nand I_26502 (I452853,I453015,I453066);
DFFARX1 I_26503 (I347161,I2507,I452882,I453106,);
nor I_26504 (I453114,I453106,I453049);
DFFARX1 I_26505 (I453114,I2507,I452882,I452847,);
nor I_26506 (I452862,I453106,I453007);
nand I_26507 (I453159,I347170,I347158);
and I_26508 (I453176,I453159,I347164);
DFFARX1 I_26509 (I453176,I2507,I452882,I453202,);
nor I_26510 (I452850,I453202,I453106);
not I_26511 (I453224,I453202);
nor I_26512 (I453241,I453224,I453015);
nor I_26513 (I453258,I452947,I453241);
DFFARX1 I_26514 (I453258,I2507,I452882,I452865,);
nor I_26515 (I453289,I453224,I453106);
nor I_26516 (I453306,I347176,I347158);
nor I_26517 (I452856,I453306,I453289);
not I_26518 (I453337,I453306);
nand I_26519 (I452859,I453066,I453337);
DFFARX1 I_26520 (I453306,I2507,I452882,I452871,);
DFFARX1 I_26521 (I453306,I2507,I452882,I452868,);
not I_26522 (I453426,I2514);
DFFARX1 I_26523 (I1228645,I2507,I453426,I453452,);
DFFARX1 I_26524 (I453452,I2507,I453426,I453469,);
not I_26525 (I453418,I453469);
not I_26526 (I453491,I453452);
nand I_26527 (I453508,I1228657,I1228660);
and I_26528 (I453525,I453508,I1228663);
DFFARX1 I_26529 (I453525,I2507,I453426,I453551,);
not I_26530 (I453559,I453551);
DFFARX1 I_26531 (I1228648,I2507,I453426,I453585,);
and I_26532 (I453593,I453585,I1228654);
nand I_26533 (I453610,I453585,I1228654);
nand I_26534 (I453397,I453559,I453610);
DFFARX1 I_26535 (I1228642,I2507,I453426,I453650,);
nor I_26536 (I453658,I453650,I453593);
DFFARX1 I_26537 (I453658,I2507,I453426,I453391,);
nor I_26538 (I453406,I453650,I453551);
nand I_26539 (I453703,I1228645,I1228666);
and I_26540 (I453720,I453703,I1228651);
DFFARX1 I_26541 (I453720,I2507,I453426,I453746,);
nor I_26542 (I453394,I453746,I453650);
not I_26543 (I453768,I453746);
nor I_26544 (I453785,I453768,I453559);
nor I_26545 (I453802,I453491,I453785);
DFFARX1 I_26546 (I453802,I2507,I453426,I453409,);
nor I_26547 (I453833,I453768,I453650);
nor I_26548 (I453850,I1228642,I1228666);
nor I_26549 (I453400,I453850,I453833);
not I_26550 (I453881,I453850);
nand I_26551 (I453403,I453610,I453881);
DFFARX1 I_26552 (I453850,I2507,I453426,I453415,);
DFFARX1 I_26553 (I453850,I2507,I453426,I453412,);
not I_26554 (I453970,I2514);
DFFARX1 I_26555 (I722045,I2507,I453970,I453996,);
DFFARX1 I_26556 (I453996,I2507,I453970,I454013,);
not I_26557 (I453962,I454013);
not I_26558 (I454035,I453996);
nand I_26559 (I454052,I722066,I722057);
and I_26560 (I454069,I454052,I722045);
DFFARX1 I_26561 (I454069,I2507,I453970,I454095,);
not I_26562 (I454103,I454095);
DFFARX1 I_26563 (I722051,I2507,I453970,I454129,);
and I_26564 (I454137,I454129,I722048);
nand I_26565 (I454154,I454129,I722048);
nand I_26566 (I453941,I454103,I454154);
DFFARX1 I_26567 (I722042,I2507,I453970,I454194,);
nor I_26568 (I454202,I454194,I454137);
DFFARX1 I_26569 (I454202,I2507,I453970,I453935,);
nor I_26570 (I453950,I454194,I454095);
nand I_26571 (I454247,I722042,I722054);
and I_26572 (I454264,I454247,I722063);
DFFARX1 I_26573 (I454264,I2507,I453970,I454290,);
nor I_26574 (I453938,I454290,I454194);
not I_26575 (I454312,I454290);
nor I_26576 (I454329,I454312,I454103);
nor I_26577 (I454346,I454035,I454329);
DFFARX1 I_26578 (I454346,I2507,I453970,I453953,);
nor I_26579 (I454377,I454312,I454194);
nor I_26580 (I454394,I722060,I722054);
nor I_26581 (I453944,I454394,I454377);
not I_26582 (I454425,I454394);
nand I_26583 (I453947,I454154,I454425);
DFFARX1 I_26584 (I454394,I2507,I453970,I453959,);
DFFARX1 I_26585 (I454394,I2507,I453970,I453956,);
not I_26586 (I454514,I2514);
DFFARX1 I_26587 (I13239,I2507,I454514,I454540,);
DFFARX1 I_26588 (I454540,I2507,I454514,I454557,);
not I_26589 (I454506,I454557);
not I_26590 (I454579,I454540);
nand I_26591 (I454596,I13227,I13242);
and I_26592 (I454613,I454596,I13230);
DFFARX1 I_26593 (I454613,I2507,I454514,I454639,);
not I_26594 (I454647,I454639);
DFFARX1 I_26595 (I13251,I2507,I454514,I454673,);
and I_26596 (I454681,I454673,I13245);
nand I_26597 (I454698,I454673,I13245);
nand I_26598 (I454485,I454647,I454698);
DFFARX1 I_26599 (I13248,I2507,I454514,I454738,);
nor I_26600 (I454746,I454738,I454681);
DFFARX1 I_26601 (I454746,I2507,I454514,I454479,);
nor I_26602 (I454494,I454738,I454639);
nand I_26603 (I454791,I13227,I13230);
and I_26604 (I454808,I454791,I13233);
DFFARX1 I_26605 (I454808,I2507,I454514,I454834,);
nor I_26606 (I454482,I454834,I454738);
not I_26607 (I454856,I454834);
nor I_26608 (I454873,I454856,I454647);
nor I_26609 (I454890,I454579,I454873);
DFFARX1 I_26610 (I454890,I2507,I454514,I454497,);
nor I_26611 (I454921,I454856,I454738);
nor I_26612 (I454938,I13236,I13230);
nor I_26613 (I454488,I454938,I454921);
not I_26614 (I454969,I454938);
nand I_26615 (I454491,I454698,I454969);
DFFARX1 I_26616 (I454938,I2507,I454514,I454503,);
DFFARX1 I_26617 (I454938,I2507,I454514,I454500,);
not I_26618 (I455058,I2514);
DFFARX1 I_26619 (I1274424,I2507,I455058,I455084,);
DFFARX1 I_26620 (I455084,I2507,I455058,I455101,);
not I_26621 (I455050,I455101);
not I_26622 (I455123,I455084);
nand I_26623 (I455140,I1274421,I1274418);
and I_26624 (I455157,I455140,I1274406);
DFFARX1 I_26625 (I455157,I2507,I455058,I455183,);
not I_26626 (I455191,I455183);
DFFARX1 I_26627 (I1274430,I2507,I455058,I455217,);
and I_26628 (I455225,I455217,I1274415);
nand I_26629 (I455242,I455217,I1274415);
nand I_26630 (I455029,I455191,I455242);
DFFARX1 I_26631 (I1274409,I2507,I455058,I455282,);
nor I_26632 (I455290,I455282,I455225);
DFFARX1 I_26633 (I455290,I2507,I455058,I455023,);
nor I_26634 (I455038,I455282,I455183);
nand I_26635 (I455335,I1274406,I1274412);
and I_26636 (I455352,I455335,I1274427);
DFFARX1 I_26637 (I455352,I2507,I455058,I455378,);
nor I_26638 (I455026,I455378,I455282);
not I_26639 (I455400,I455378);
nor I_26640 (I455417,I455400,I455191);
nor I_26641 (I455434,I455123,I455417);
DFFARX1 I_26642 (I455434,I2507,I455058,I455041,);
nor I_26643 (I455465,I455400,I455282);
nor I_26644 (I455482,I1274409,I1274412);
nor I_26645 (I455032,I455482,I455465);
not I_26646 (I455513,I455482);
nand I_26647 (I455035,I455242,I455513);
DFFARX1 I_26648 (I455482,I2507,I455058,I455047,);
DFFARX1 I_26649 (I455482,I2507,I455058,I455044,);
not I_26650 (I455602,I2514);
DFFARX1 I_26651 (I570031,I2507,I455602,I455628,);
DFFARX1 I_26652 (I455628,I2507,I455602,I455645,);
not I_26653 (I455594,I455645);
not I_26654 (I455667,I455628);
nand I_26655 (I455684,I570028,I570049);
and I_26656 (I455701,I455684,I570052);
DFFARX1 I_26657 (I455701,I2507,I455602,I455727,);
not I_26658 (I455735,I455727);
DFFARX1 I_26659 (I570037,I2507,I455602,I455761,);
and I_26660 (I455769,I455761,I570040);
nand I_26661 (I455786,I455761,I570040);
nand I_26662 (I455573,I455735,I455786);
DFFARX1 I_26663 (I570043,I2507,I455602,I455826,);
nor I_26664 (I455834,I455826,I455769);
DFFARX1 I_26665 (I455834,I2507,I455602,I455567,);
nor I_26666 (I455582,I455826,I455727);
nand I_26667 (I455879,I570028,I570034);
and I_26668 (I455896,I455879,I570046);
DFFARX1 I_26669 (I455896,I2507,I455602,I455922,);
nor I_26670 (I455570,I455922,I455826);
not I_26671 (I455944,I455922);
nor I_26672 (I455961,I455944,I455735);
nor I_26673 (I455978,I455667,I455961);
DFFARX1 I_26674 (I455978,I2507,I455602,I455585,);
nor I_26675 (I456009,I455944,I455826);
nor I_26676 (I456026,I570031,I570034);
nor I_26677 (I455576,I456026,I456009);
not I_26678 (I456057,I456026);
nand I_26679 (I455579,I455786,I456057);
DFFARX1 I_26680 (I456026,I2507,I455602,I455591,);
DFFARX1 I_26681 (I456026,I2507,I455602,I455588,);
not I_26682 (I456146,I2514);
DFFARX1 I_26683 (I764817,I2507,I456146,I456172,);
DFFARX1 I_26684 (I456172,I2507,I456146,I456189,);
not I_26685 (I456138,I456189);
not I_26686 (I456211,I456172);
nand I_26687 (I456228,I764838,I764829);
and I_26688 (I456245,I456228,I764817);
DFFARX1 I_26689 (I456245,I2507,I456146,I456271,);
not I_26690 (I456279,I456271);
DFFARX1 I_26691 (I764823,I2507,I456146,I456305,);
and I_26692 (I456313,I456305,I764820);
nand I_26693 (I456330,I456305,I764820);
nand I_26694 (I456117,I456279,I456330);
DFFARX1 I_26695 (I764814,I2507,I456146,I456370,);
nor I_26696 (I456378,I456370,I456313);
DFFARX1 I_26697 (I456378,I2507,I456146,I456111,);
nor I_26698 (I456126,I456370,I456271);
nand I_26699 (I456423,I764814,I764826);
and I_26700 (I456440,I456423,I764835);
DFFARX1 I_26701 (I456440,I2507,I456146,I456466,);
nor I_26702 (I456114,I456466,I456370);
not I_26703 (I456488,I456466);
nor I_26704 (I456505,I456488,I456279);
nor I_26705 (I456522,I456211,I456505);
DFFARX1 I_26706 (I456522,I2507,I456146,I456129,);
nor I_26707 (I456553,I456488,I456370);
nor I_26708 (I456570,I764832,I764826);
nor I_26709 (I456120,I456570,I456553);
not I_26710 (I456601,I456570);
nand I_26711 (I456123,I456330,I456601);
DFFARX1 I_26712 (I456570,I2507,I456146,I456135,);
DFFARX1 I_26713 (I456570,I2507,I456146,I456132,);
not I_26714 (I456690,I2514);
DFFARX1 I_26715 (I752101,I2507,I456690,I456716,);
DFFARX1 I_26716 (I456716,I2507,I456690,I456733,);
not I_26717 (I456682,I456733);
not I_26718 (I456755,I456716);
nand I_26719 (I456772,I752122,I752113);
and I_26720 (I456789,I456772,I752101);
DFFARX1 I_26721 (I456789,I2507,I456690,I456815,);
not I_26722 (I456823,I456815);
DFFARX1 I_26723 (I752107,I2507,I456690,I456849,);
and I_26724 (I456857,I456849,I752104);
nand I_26725 (I456874,I456849,I752104);
nand I_26726 (I456661,I456823,I456874);
DFFARX1 I_26727 (I752098,I2507,I456690,I456914,);
nor I_26728 (I456922,I456914,I456857);
DFFARX1 I_26729 (I456922,I2507,I456690,I456655,);
nor I_26730 (I456670,I456914,I456815);
nand I_26731 (I456967,I752098,I752110);
and I_26732 (I456984,I456967,I752119);
DFFARX1 I_26733 (I456984,I2507,I456690,I457010,);
nor I_26734 (I456658,I457010,I456914);
not I_26735 (I457032,I457010);
nor I_26736 (I457049,I457032,I456823);
nor I_26737 (I457066,I456755,I457049);
DFFARX1 I_26738 (I457066,I2507,I456690,I456673,);
nor I_26739 (I457097,I457032,I456914);
nor I_26740 (I457114,I752116,I752110);
nor I_26741 (I456664,I457114,I457097);
not I_26742 (I457145,I457114);
nand I_26743 (I456667,I456874,I457145);
DFFARX1 I_26744 (I457114,I2507,I456690,I456679,);
DFFARX1 I_26745 (I457114,I2507,I456690,I456676,);
not I_26746 (I457234,I2514);
DFFARX1 I_26747 (I691411,I2507,I457234,I457260,);
DFFARX1 I_26748 (I457260,I2507,I457234,I457277,);
not I_26749 (I457226,I457277);
not I_26750 (I457299,I457260);
nand I_26751 (I457316,I691432,I691423);
and I_26752 (I457333,I457316,I691411);
DFFARX1 I_26753 (I457333,I2507,I457234,I457359,);
not I_26754 (I457367,I457359);
DFFARX1 I_26755 (I691417,I2507,I457234,I457393,);
and I_26756 (I457401,I457393,I691414);
nand I_26757 (I457418,I457393,I691414);
nand I_26758 (I457205,I457367,I457418);
DFFARX1 I_26759 (I691408,I2507,I457234,I457458,);
nor I_26760 (I457466,I457458,I457401);
DFFARX1 I_26761 (I457466,I2507,I457234,I457199,);
nor I_26762 (I457214,I457458,I457359);
nand I_26763 (I457511,I691408,I691420);
and I_26764 (I457528,I457511,I691429);
DFFARX1 I_26765 (I457528,I2507,I457234,I457554,);
nor I_26766 (I457202,I457554,I457458);
not I_26767 (I457576,I457554);
nor I_26768 (I457593,I457576,I457367);
nor I_26769 (I457610,I457299,I457593);
DFFARX1 I_26770 (I457610,I2507,I457234,I457217,);
nor I_26771 (I457641,I457576,I457458);
nor I_26772 (I457658,I691426,I691420);
nor I_26773 (I457208,I457658,I457641);
not I_26774 (I457689,I457658);
nand I_26775 (I457211,I457418,I457689);
DFFARX1 I_26776 (I457658,I2507,I457234,I457223,);
DFFARX1 I_26777 (I457658,I2507,I457234,I457220,);
not I_26778 (I457778,I2514);
DFFARX1 I_26779 (I1089585,I2507,I457778,I457804,);
DFFARX1 I_26780 (I457804,I2507,I457778,I457821,);
not I_26781 (I457770,I457821);
not I_26782 (I457843,I457804);
nand I_26783 (I457860,I1089597,I1089585);
and I_26784 (I457877,I457860,I1089588);
DFFARX1 I_26785 (I457877,I2507,I457778,I457903,);
not I_26786 (I457911,I457903);
DFFARX1 I_26787 (I1089606,I2507,I457778,I457937,);
and I_26788 (I457945,I457937,I1089582);
nand I_26789 (I457962,I457937,I1089582);
nand I_26790 (I457749,I457911,I457962);
DFFARX1 I_26791 (I1089600,I2507,I457778,I458002,);
nor I_26792 (I458010,I458002,I457945);
DFFARX1 I_26793 (I458010,I2507,I457778,I457743,);
nor I_26794 (I457758,I458002,I457903);
nand I_26795 (I458055,I1089594,I1089591);
and I_26796 (I458072,I458055,I1089603);
DFFARX1 I_26797 (I458072,I2507,I457778,I458098,);
nor I_26798 (I457746,I458098,I458002);
not I_26799 (I458120,I458098);
nor I_26800 (I458137,I458120,I457911);
nor I_26801 (I458154,I457843,I458137);
DFFARX1 I_26802 (I458154,I2507,I457778,I457761,);
nor I_26803 (I458185,I458120,I458002);
nor I_26804 (I458202,I1089582,I1089591);
nor I_26805 (I457752,I458202,I458185);
not I_26806 (I458233,I458202);
nand I_26807 (I457755,I457962,I458233);
DFFARX1 I_26808 (I458202,I2507,I457778,I457767,);
DFFARX1 I_26809 (I458202,I2507,I457778,I457764,);
not I_26810 (I458322,I2514);
DFFARX1 I_26811 (I590839,I2507,I458322,I458348,);
DFFARX1 I_26812 (I458348,I2507,I458322,I458365,);
not I_26813 (I458314,I458365);
not I_26814 (I458387,I458348);
nand I_26815 (I458404,I590836,I590857);
and I_26816 (I458421,I458404,I590860);
DFFARX1 I_26817 (I458421,I2507,I458322,I458447,);
not I_26818 (I458455,I458447);
DFFARX1 I_26819 (I590845,I2507,I458322,I458481,);
and I_26820 (I458489,I458481,I590848);
nand I_26821 (I458506,I458481,I590848);
nand I_26822 (I458293,I458455,I458506);
DFFARX1 I_26823 (I590851,I2507,I458322,I458546,);
nor I_26824 (I458554,I458546,I458489);
DFFARX1 I_26825 (I458554,I2507,I458322,I458287,);
nor I_26826 (I458302,I458546,I458447);
nand I_26827 (I458599,I590836,I590842);
and I_26828 (I458616,I458599,I590854);
DFFARX1 I_26829 (I458616,I2507,I458322,I458642,);
nor I_26830 (I458290,I458642,I458546);
not I_26831 (I458664,I458642);
nor I_26832 (I458681,I458664,I458455);
nor I_26833 (I458698,I458387,I458681);
DFFARX1 I_26834 (I458698,I2507,I458322,I458305,);
nor I_26835 (I458729,I458664,I458546);
nor I_26836 (I458746,I590839,I590842);
nor I_26837 (I458296,I458746,I458729);
not I_26838 (I458777,I458746);
nand I_26839 (I458299,I458506,I458777);
DFFARX1 I_26840 (I458746,I2507,I458322,I458311,);
DFFARX1 I_26841 (I458746,I2507,I458322,I458308,);
not I_26842 (I458866,I2514);
DFFARX1 I_26843 (I1171083,I2507,I458866,I458892,);
DFFARX1 I_26844 (I458892,I2507,I458866,I458909,);
not I_26845 (I458858,I458909);
not I_26846 (I458931,I458892);
nand I_26847 (I458948,I1171095,I1171083);
and I_26848 (I458965,I458948,I1171086);
DFFARX1 I_26849 (I458965,I2507,I458866,I458991,);
not I_26850 (I458999,I458991);
DFFARX1 I_26851 (I1171104,I2507,I458866,I459025,);
and I_26852 (I459033,I459025,I1171080);
nand I_26853 (I459050,I459025,I1171080);
nand I_26854 (I458837,I458999,I459050);
DFFARX1 I_26855 (I1171098,I2507,I458866,I459090,);
nor I_26856 (I459098,I459090,I459033);
DFFARX1 I_26857 (I459098,I2507,I458866,I458831,);
nor I_26858 (I458846,I459090,I458991);
nand I_26859 (I459143,I1171092,I1171089);
and I_26860 (I459160,I459143,I1171101);
DFFARX1 I_26861 (I459160,I2507,I458866,I459186,);
nor I_26862 (I458834,I459186,I459090);
not I_26863 (I459208,I459186);
nor I_26864 (I459225,I459208,I458999);
nor I_26865 (I459242,I458931,I459225);
DFFARX1 I_26866 (I459242,I2507,I458866,I458849,);
nor I_26867 (I459273,I459208,I459090);
nor I_26868 (I459290,I1171080,I1171089);
nor I_26869 (I458840,I459290,I459273);
not I_26870 (I459321,I459290);
nand I_26871 (I458843,I459050,I459321);
DFFARX1 I_26872 (I459290,I2507,I458866,I458855,);
DFFARX1 I_26873 (I459290,I2507,I458866,I458852,);
not I_26874 (I459410,I2514);
DFFARX1 I_26875 (I1061263,I2507,I459410,I459436,);
DFFARX1 I_26876 (I459436,I2507,I459410,I459453,);
not I_26877 (I459402,I459453);
not I_26878 (I459475,I459436);
nand I_26879 (I459492,I1061275,I1061263);
and I_26880 (I459509,I459492,I1061266);
DFFARX1 I_26881 (I459509,I2507,I459410,I459535,);
not I_26882 (I459543,I459535);
DFFARX1 I_26883 (I1061284,I2507,I459410,I459569,);
and I_26884 (I459577,I459569,I1061260);
nand I_26885 (I459594,I459569,I1061260);
nand I_26886 (I459381,I459543,I459594);
DFFARX1 I_26887 (I1061278,I2507,I459410,I459634,);
nor I_26888 (I459642,I459634,I459577);
DFFARX1 I_26889 (I459642,I2507,I459410,I459375,);
nor I_26890 (I459390,I459634,I459535);
nand I_26891 (I459687,I1061272,I1061269);
and I_26892 (I459704,I459687,I1061281);
DFFARX1 I_26893 (I459704,I2507,I459410,I459730,);
nor I_26894 (I459378,I459730,I459634);
not I_26895 (I459752,I459730);
nor I_26896 (I459769,I459752,I459543);
nor I_26897 (I459786,I459475,I459769);
DFFARX1 I_26898 (I459786,I2507,I459410,I459393,);
nor I_26899 (I459817,I459752,I459634);
nor I_26900 (I459834,I1061260,I1061269);
nor I_26901 (I459384,I459834,I459817);
not I_26902 (I459865,I459834);
nand I_26903 (I459387,I459594,I459865);
DFFARX1 I_26904 (I459834,I2507,I459410,I459399,);
DFFARX1 I_26905 (I459834,I2507,I459410,I459396,);
not I_26906 (I459954,I2514);
DFFARX1 I_26907 (I504207,I2507,I459954,I459980,);
DFFARX1 I_26908 (I459980,I2507,I459954,I459997,);
not I_26909 (I459946,I459997);
not I_26910 (I460019,I459980);
nand I_26911 (I460036,I504210,I504228);
and I_26912 (I460053,I460036,I504216);
DFFARX1 I_26913 (I460053,I2507,I459954,I460079,);
not I_26914 (I460087,I460079);
DFFARX1 I_26915 (I504207,I2507,I459954,I460113,);
and I_26916 (I460121,I460113,I504225);
nand I_26917 (I460138,I460113,I504225);
nand I_26918 (I459925,I460087,I460138);
DFFARX1 I_26919 (I504219,I2507,I459954,I460178,);
nor I_26920 (I460186,I460178,I460121);
DFFARX1 I_26921 (I460186,I2507,I459954,I459919,);
nor I_26922 (I459934,I460178,I460079);
nand I_26923 (I460231,I504222,I504204);
and I_26924 (I460248,I460231,I504213);
DFFARX1 I_26925 (I460248,I2507,I459954,I460274,);
nor I_26926 (I459922,I460274,I460178);
not I_26927 (I460296,I460274);
nor I_26928 (I460313,I460296,I460087);
nor I_26929 (I460330,I460019,I460313);
DFFARX1 I_26930 (I460330,I2507,I459954,I459937,);
nor I_26931 (I460361,I460296,I460178);
nor I_26932 (I460378,I504204,I504204);
nor I_26933 (I459928,I460378,I460361);
not I_26934 (I460409,I460378);
nand I_26935 (I459931,I460138,I460409);
DFFARX1 I_26936 (I460378,I2507,I459954,I459943,);
DFFARX1 I_26937 (I460378,I2507,I459954,I459940,);
not I_26938 (I460498,I2514);
DFFARX1 I_26939 (I1003211,I2507,I460498,I460524,);
DFFARX1 I_26940 (I460524,I2507,I460498,I460541,);
not I_26941 (I460490,I460541);
not I_26942 (I460563,I460524);
nand I_26943 (I460580,I1003226,I1003214);
and I_26944 (I460597,I460580,I1003205);
DFFARX1 I_26945 (I460597,I2507,I460498,I460623,);
not I_26946 (I460631,I460623);
DFFARX1 I_26947 (I1003217,I2507,I460498,I460657,);
and I_26948 (I460665,I460657,I1003208);
nand I_26949 (I460682,I460657,I1003208);
nand I_26950 (I460469,I460631,I460682);
DFFARX1 I_26951 (I1003223,I2507,I460498,I460722,);
nor I_26952 (I460730,I460722,I460665);
DFFARX1 I_26953 (I460730,I2507,I460498,I460463,);
nor I_26954 (I460478,I460722,I460623);
nand I_26955 (I460775,I1003232,I1003220);
and I_26956 (I460792,I460775,I1003229);
DFFARX1 I_26957 (I460792,I2507,I460498,I460818,);
nor I_26958 (I460466,I460818,I460722);
not I_26959 (I460840,I460818);
nor I_26960 (I460857,I460840,I460631);
nor I_26961 (I460874,I460563,I460857);
DFFARX1 I_26962 (I460874,I2507,I460498,I460481,);
nor I_26963 (I460905,I460840,I460722);
nor I_26964 (I460922,I1003205,I1003220);
nor I_26965 (I460472,I460922,I460905);
not I_26966 (I460953,I460922);
nand I_26967 (I460475,I460682,I460953);
DFFARX1 I_26968 (I460922,I2507,I460498,I460487,);
DFFARX1 I_26969 (I460922,I2507,I460498,I460484,);
not I_26970 (I461042,I2514);
DFFARX1 I_26971 (I2484,I2507,I461042,I461068,);
DFFARX1 I_26972 (I461068,I2507,I461042,I461085,);
not I_26973 (I461034,I461085);
not I_26974 (I461107,I461068);
nand I_26975 (I461124,I1676,I1612);
and I_26976 (I461141,I461124,I1876);
DFFARX1 I_26977 (I461141,I2507,I461042,I461167,);
not I_26978 (I461175,I461167);
DFFARX1 I_26979 (I1996,I2507,I461042,I461201,);
and I_26980 (I461209,I461201,I1884);
nand I_26981 (I461226,I461201,I1884);
nand I_26982 (I461013,I461175,I461226);
DFFARX1 I_26983 (I2148,I2507,I461042,I461266,);
nor I_26984 (I461274,I461266,I461209);
DFFARX1 I_26985 (I461274,I2507,I461042,I461007,);
nor I_26986 (I461022,I461266,I461167);
nand I_26987 (I461319,I1780,I1908);
and I_26988 (I461336,I461319,I1796);
DFFARX1 I_26989 (I461336,I2507,I461042,I461362,);
nor I_26990 (I461010,I461362,I461266);
not I_26991 (I461384,I461362);
nor I_26992 (I461401,I461384,I461175);
nor I_26993 (I461418,I461107,I461401);
DFFARX1 I_26994 (I461418,I2507,I461042,I461025,);
nor I_26995 (I461449,I461384,I461266);
nor I_26996 (I461466,I2140,I1908);
nor I_26997 (I461016,I461466,I461449);
not I_26998 (I461497,I461466);
nand I_26999 (I461019,I461226,I461497);
DFFARX1 I_27000 (I461466,I2507,I461042,I461031,);
DFFARX1 I_27001 (I461466,I2507,I461042,I461028,);
not I_27002 (I461586,I2514);
DFFARX1 I_27003 (I1168193,I2507,I461586,I461612,);
DFFARX1 I_27004 (I461612,I2507,I461586,I461629,);
not I_27005 (I461578,I461629);
not I_27006 (I461651,I461612);
nand I_27007 (I461668,I1168205,I1168193);
and I_27008 (I461685,I461668,I1168196);
DFFARX1 I_27009 (I461685,I2507,I461586,I461711,);
not I_27010 (I461719,I461711);
DFFARX1 I_27011 (I1168214,I2507,I461586,I461745,);
and I_27012 (I461753,I461745,I1168190);
nand I_27013 (I461770,I461745,I1168190);
nand I_27014 (I461557,I461719,I461770);
DFFARX1 I_27015 (I1168208,I2507,I461586,I461810,);
nor I_27016 (I461818,I461810,I461753);
DFFARX1 I_27017 (I461818,I2507,I461586,I461551,);
nor I_27018 (I461566,I461810,I461711);
nand I_27019 (I461863,I1168202,I1168199);
and I_27020 (I461880,I461863,I1168211);
DFFARX1 I_27021 (I461880,I2507,I461586,I461906,);
nor I_27022 (I461554,I461906,I461810);
not I_27023 (I461928,I461906);
nor I_27024 (I461945,I461928,I461719);
nor I_27025 (I461962,I461651,I461945);
DFFARX1 I_27026 (I461962,I2507,I461586,I461569,);
nor I_27027 (I461993,I461928,I461810);
nor I_27028 (I462010,I1168190,I1168199);
nor I_27029 (I461560,I462010,I461993);
not I_27030 (I462041,I462010);
nand I_27031 (I461563,I461770,I462041);
DFFARX1 I_27032 (I462010,I2507,I461586,I461575,);
DFFARX1 I_27033 (I462010,I2507,I461586,I461572,);
not I_27034 (I462130,I2514);
DFFARX1 I_27035 (I816489,I2507,I462130,I462156,);
DFFARX1 I_27036 (I462156,I2507,I462130,I462173,);
not I_27037 (I462122,I462173);
not I_27038 (I462195,I462156);
nand I_27039 (I462212,I816483,I816480);
and I_27040 (I462229,I462212,I816495);
DFFARX1 I_27041 (I462229,I2507,I462130,I462255,);
not I_27042 (I462263,I462255);
DFFARX1 I_27043 (I816483,I2507,I462130,I462289,);
and I_27044 (I462297,I462289,I816477);
nand I_27045 (I462314,I462289,I816477);
nand I_27046 (I462101,I462263,I462314);
DFFARX1 I_27047 (I816477,I2507,I462130,I462354,);
nor I_27048 (I462362,I462354,I462297);
DFFARX1 I_27049 (I462362,I2507,I462130,I462095,);
nor I_27050 (I462110,I462354,I462255);
nand I_27051 (I462407,I816492,I816486);
and I_27052 (I462424,I462407,I816480);
DFFARX1 I_27053 (I462424,I2507,I462130,I462450,);
nor I_27054 (I462098,I462450,I462354);
not I_27055 (I462472,I462450);
nor I_27056 (I462489,I462472,I462263);
nor I_27057 (I462506,I462195,I462489);
DFFARX1 I_27058 (I462506,I2507,I462130,I462113,);
nor I_27059 (I462537,I462472,I462354);
nor I_27060 (I462554,I816498,I816486);
nor I_27061 (I462104,I462554,I462537);
not I_27062 (I462585,I462554);
nand I_27063 (I462107,I462314,I462585);
DFFARX1 I_27064 (I462554,I2507,I462130,I462119,);
DFFARX1 I_27065 (I462554,I2507,I462130,I462116,);
not I_27066 (I462674,I2514);
DFFARX1 I_27067 (I523842,I2507,I462674,I462700,);
DFFARX1 I_27068 (I462700,I2507,I462674,I462717,);
not I_27069 (I462666,I462717);
not I_27070 (I462739,I462700);
nand I_27071 (I462756,I523845,I523863);
and I_27072 (I462773,I462756,I523851);
DFFARX1 I_27073 (I462773,I2507,I462674,I462799,);
not I_27074 (I462807,I462799);
DFFARX1 I_27075 (I523842,I2507,I462674,I462833,);
and I_27076 (I462841,I462833,I523860);
nand I_27077 (I462858,I462833,I523860);
nand I_27078 (I462645,I462807,I462858);
DFFARX1 I_27079 (I523854,I2507,I462674,I462898,);
nor I_27080 (I462906,I462898,I462841);
DFFARX1 I_27081 (I462906,I2507,I462674,I462639,);
nor I_27082 (I462654,I462898,I462799);
nand I_27083 (I462951,I523857,I523839);
and I_27084 (I462968,I462951,I523848);
DFFARX1 I_27085 (I462968,I2507,I462674,I462994,);
nor I_27086 (I462642,I462994,I462898);
not I_27087 (I463016,I462994);
nor I_27088 (I463033,I463016,I462807);
nor I_27089 (I463050,I462739,I463033);
DFFARX1 I_27090 (I463050,I2507,I462674,I462657,);
nor I_27091 (I463081,I463016,I462898);
nor I_27092 (I463098,I523839,I523839);
nor I_27093 (I462648,I463098,I463081);
not I_27094 (I463129,I463098);
nand I_27095 (I462651,I462858,I463129);
DFFARX1 I_27096 (I463098,I2507,I462674,I462663,);
DFFARX1 I_27097 (I463098,I2507,I462674,I462660,);
not I_27098 (I463218,I2514);
DFFARX1 I_27099 (I963805,I2507,I463218,I463244,);
DFFARX1 I_27100 (I463244,I2507,I463218,I463261,);
not I_27101 (I463210,I463261);
not I_27102 (I463283,I463244);
nand I_27103 (I463300,I963820,I963808);
and I_27104 (I463317,I463300,I963799);
DFFARX1 I_27105 (I463317,I2507,I463218,I463343,);
not I_27106 (I463351,I463343);
DFFARX1 I_27107 (I963811,I2507,I463218,I463377,);
and I_27108 (I463385,I463377,I963802);
nand I_27109 (I463402,I463377,I963802);
nand I_27110 (I463189,I463351,I463402);
DFFARX1 I_27111 (I963817,I2507,I463218,I463442,);
nor I_27112 (I463450,I463442,I463385);
DFFARX1 I_27113 (I463450,I2507,I463218,I463183,);
nor I_27114 (I463198,I463442,I463343);
nand I_27115 (I463495,I963826,I963814);
and I_27116 (I463512,I463495,I963823);
DFFARX1 I_27117 (I463512,I2507,I463218,I463538,);
nor I_27118 (I463186,I463538,I463442);
not I_27119 (I463560,I463538);
nor I_27120 (I463577,I463560,I463351);
nor I_27121 (I463594,I463283,I463577);
DFFARX1 I_27122 (I463594,I2507,I463218,I463201,);
nor I_27123 (I463625,I463560,I463442);
nor I_27124 (I463642,I963799,I963814);
nor I_27125 (I463192,I463642,I463625);
not I_27126 (I463673,I463642);
nand I_27127 (I463195,I463402,I463673);
DFFARX1 I_27128 (I463642,I2507,I463218,I463207,);
DFFARX1 I_27129 (I463642,I2507,I463218,I463204,);
not I_27130 (I463762,I2514);
DFFARX1 I_27131 (I69095,I2507,I463762,I463788,);
DFFARX1 I_27132 (I463788,I2507,I463762,I463805,);
not I_27133 (I463754,I463805);
not I_27134 (I463827,I463788);
nand I_27135 (I463844,I69110,I69089);
and I_27136 (I463861,I463844,I69092);
DFFARX1 I_27137 (I463861,I2507,I463762,I463887,);
not I_27138 (I463895,I463887);
DFFARX1 I_27139 (I69098,I2507,I463762,I463921,);
and I_27140 (I463929,I463921,I69092);
nand I_27141 (I463946,I463921,I69092);
nand I_27142 (I463733,I463895,I463946);
DFFARX1 I_27143 (I69107,I2507,I463762,I463986,);
nor I_27144 (I463994,I463986,I463929);
DFFARX1 I_27145 (I463994,I2507,I463762,I463727,);
nor I_27146 (I463742,I463986,I463887);
nand I_27147 (I464039,I69089,I69104);
and I_27148 (I464056,I464039,I69101);
DFFARX1 I_27149 (I464056,I2507,I463762,I464082,);
nor I_27150 (I463730,I464082,I463986);
not I_27151 (I464104,I464082);
nor I_27152 (I464121,I464104,I463895);
nor I_27153 (I464138,I463827,I464121);
DFFARX1 I_27154 (I464138,I2507,I463762,I463745,);
nor I_27155 (I464169,I464104,I463986);
nor I_27156 (I464186,I69113,I69104);
nor I_27157 (I463736,I464186,I464169);
not I_27158 (I464217,I464186);
nand I_27159 (I463739,I463946,I464217);
DFFARX1 I_27160 (I464186,I2507,I463762,I463751,);
DFFARX1 I_27161 (I464186,I2507,I463762,I463748,);
not I_27162 (I464306,I2514);
DFFARX1 I_27163 (I100188,I2507,I464306,I464332,);
DFFARX1 I_27164 (I464332,I2507,I464306,I464349,);
not I_27165 (I464298,I464349);
not I_27166 (I464371,I464332);
nand I_27167 (I464388,I100203,I100182);
and I_27168 (I464405,I464388,I100185);
DFFARX1 I_27169 (I464405,I2507,I464306,I464431,);
not I_27170 (I464439,I464431);
DFFARX1 I_27171 (I100191,I2507,I464306,I464465,);
and I_27172 (I464473,I464465,I100185);
nand I_27173 (I464490,I464465,I100185);
nand I_27174 (I464277,I464439,I464490);
DFFARX1 I_27175 (I100200,I2507,I464306,I464530,);
nor I_27176 (I464538,I464530,I464473);
DFFARX1 I_27177 (I464538,I2507,I464306,I464271,);
nor I_27178 (I464286,I464530,I464431);
nand I_27179 (I464583,I100182,I100197);
and I_27180 (I464600,I464583,I100194);
DFFARX1 I_27181 (I464600,I2507,I464306,I464626,);
nor I_27182 (I464274,I464626,I464530);
not I_27183 (I464648,I464626);
nor I_27184 (I464665,I464648,I464439);
nor I_27185 (I464682,I464371,I464665);
DFFARX1 I_27186 (I464682,I2507,I464306,I464289,);
nor I_27187 (I464713,I464648,I464530);
nor I_27188 (I464730,I100206,I100197);
nor I_27189 (I464280,I464730,I464713);
not I_27190 (I464761,I464730);
nand I_27191 (I464283,I464490,I464761);
DFFARX1 I_27192 (I464730,I2507,I464306,I464295,);
DFFARX1 I_27193 (I464730,I2507,I464306,I464292,);
not I_27194 (I464850,I2514);
DFFARX1 I_27195 (I769441,I2507,I464850,I464876,);
DFFARX1 I_27196 (I464876,I2507,I464850,I464893,);
not I_27197 (I464842,I464893);
not I_27198 (I464915,I464876);
nand I_27199 (I464932,I769462,I769453);
and I_27200 (I464949,I464932,I769441);
DFFARX1 I_27201 (I464949,I2507,I464850,I464975,);
not I_27202 (I464983,I464975);
DFFARX1 I_27203 (I769447,I2507,I464850,I465009,);
and I_27204 (I465017,I465009,I769444);
nand I_27205 (I465034,I465009,I769444);
nand I_27206 (I464821,I464983,I465034);
DFFARX1 I_27207 (I769438,I2507,I464850,I465074,);
nor I_27208 (I465082,I465074,I465017);
DFFARX1 I_27209 (I465082,I2507,I464850,I464815,);
nor I_27210 (I464830,I465074,I464975);
nand I_27211 (I465127,I769438,I769450);
and I_27212 (I465144,I465127,I769459);
DFFARX1 I_27213 (I465144,I2507,I464850,I465170,);
nor I_27214 (I464818,I465170,I465074);
not I_27215 (I465192,I465170);
nor I_27216 (I465209,I465192,I464983);
nor I_27217 (I465226,I464915,I465209);
DFFARX1 I_27218 (I465226,I2507,I464850,I464833,);
nor I_27219 (I465257,I465192,I465074);
nor I_27220 (I465274,I769456,I769450);
nor I_27221 (I464824,I465274,I465257);
not I_27222 (I465305,I465274);
nand I_27223 (I464827,I465034,I465305);
DFFARX1 I_27224 (I465274,I2507,I464850,I464839,);
DFFARX1 I_27225 (I465274,I2507,I464850,I464836,);
not I_27226 (I465394,I2514);
DFFARX1 I_27227 (I959283,I2507,I465394,I465420,);
DFFARX1 I_27228 (I465420,I2507,I465394,I465437,);
not I_27229 (I465386,I465437);
not I_27230 (I465459,I465420);
nand I_27231 (I465476,I959298,I959286);
and I_27232 (I465493,I465476,I959277);
DFFARX1 I_27233 (I465493,I2507,I465394,I465519,);
not I_27234 (I465527,I465519);
DFFARX1 I_27235 (I959289,I2507,I465394,I465553,);
and I_27236 (I465561,I465553,I959280);
nand I_27237 (I465578,I465553,I959280);
nand I_27238 (I465365,I465527,I465578);
DFFARX1 I_27239 (I959295,I2507,I465394,I465618,);
nor I_27240 (I465626,I465618,I465561);
DFFARX1 I_27241 (I465626,I2507,I465394,I465359,);
nor I_27242 (I465374,I465618,I465519);
nand I_27243 (I465671,I959304,I959292);
and I_27244 (I465688,I465671,I959301);
DFFARX1 I_27245 (I465688,I2507,I465394,I465714,);
nor I_27246 (I465362,I465714,I465618);
not I_27247 (I465736,I465714);
nor I_27248 (I465753,I465736,I465527);
nor I_27249 (I465770,I465459,I465753);
DFFARX1 I_27250 (I465770,I2507,I465394,I465377,);
nor I_27251 (I465801,I465736,I465618);
nor I_27252 (I465818,I959277,I959292);
nor I_27253 (I465368,I465818,I465801);
not I_27254 (I465849,I465818);
nand I_27255 (I465371,I465578,I465849);
DFFARX1 I_27256 (I465818,I2507,I465394,I465383,);
DFFARX1 I_27257 (I465818,I2507,I465394,I465380,);
not I_27258 (I465938,I2514);
DFFARX1 I_27259 (I877621,I2507,I465938,I465964,);
DFFARX1 I_27260 (I465964,I2507,I465938,I465981,);
not I_27261 (I465930,I465981);
not I_27262 (I466003,I465964);
nand I_27263 (I466020,I877615,I877612);
and I_27264 (I466037,I466020,I877627);
DFFARX1 I_27265 (I466037,I2507,I465938,I466063,);
not I_27266 (I466071,I466063);
DFFARX1 I_27267 (I877615,I2507,I465938,I466097,);
and I_27268 (I466105,I466097,I877609);
nand I_27269 (I466122,I466097,I877609);
nand I_27270 (I465909,I466071,I466122);
DFFARX1 I_27271 (I877609,I2507,I465938,I466162,);
nor I_27272 (I466170,I466162,I466105);
DFFARX1 I_27273 (I466170,I2507,I465938,I465903,);
nor I_27274 (I465918,I466162,I466063);
nand I_27275 (I466215,I877624,I877618);
and I_27276 (I466232,I466215,I877612);
DFFARX1 I_27277 (I466232,I2507,I465938,I466258,);
nor I_27278 (I465906,I466258,I466162);
not I_27279 (I466280,I466258);
nor I_27280 (I466297,I466280,I466071);
nor I_27281 (I466314,I466003,I466297);
DFFARX1 I_27282 (I466314,I2507,I465938,I465921,);
nor I_27283 (I466345,I466280,I466162);
nor I_27284 (I466362,I877630,I877618);
nor I_27285 (I465912,I466362,I466345);
not I_27286 (I466393,I466362);
nand I_27287 (I465915,I466122,I466393);
DFFARX1 I_27288 (I466362,I2507,I465938,I465927,);
DFFARX1 I_27289 (I466362,I2507,I465938,I465924,);
not I_27290 (I466482,I2514);
DFFARX1 I_27291 (I323991,I2507,I466482,I466508,);
DFFARX1 I_27292 (I466508,I2507,I466482,I466525,);
not I_27293 (I466474,I466525);
not I_27294 (I466547,I466508);
nand I_27295 (I466564,I323970,I323994);
and I_27296 (I466581,I466564,I323997);
DFFARX1 I_27297 (I466581,I2507,I466482,I466607,);
not I_27298 (I466615,I466607);
DFFARX1 I_27299 (I323979,I2507,I466482,I466641,);
and I_27300 (I466649,I466641,I323985);
nand I_27301 (I466666,I466641,I323985);
nand I_27302 (I466453,I466615,I466666);
DFFARX1 I_27303 (I323973,I2507,I466482,I466706,);
nor I_27304 (I466714,I466706,I466649);
DFFARX1 I_27305 (I466714,I2507,I466482,I466447,);
nor I_27306 (I466462,I466706,I466607);
nand I_27307 (I466759,I323982,I323970);
and I_27308 (I466776,I466759,I323976);
DFFARX1 I_27309 (I466776,I2507,I466482,I466802,);
nor I_27310 (I466450,I466802,I466706);
not I_27311 (I466824,I466802);
nor I_27312 (I466841,I466824,I466615);
nor I_27313 (I466858,I466547,I466841);
DFFARX1 I_27314 (I466858,I2507,I466482,I466465,);
nor I_27315 (I466889,I466824,I466706);
nor I_27316 (I466906,I323988,I323970);
nor I_27317 (I466456,I466906,I466889);
not I_27318 (I466937,I466906);
nand I_27319 (I466459,I466666,I466937);
DFFARX1 I_27320 (I466906,I2507,I466482,I466471,);
DFFARX1 I_27321 (I466906,I2507,I466482,I466468,);
not I_27322 (I467026,I2514);
DFFARX1 I_27323 (I934089,I2507,I467026,I467052,);
DFFARX1 I_27324 (I467052,I2507,I467026,I467069,);
not I_27325 (I467018,I467069);
not I_27326 (I467091,I467052);
nand I_27327 (I467108,I934104,I934092);
and I_27328 (I467125,I467108,I934083);
DFFARX1 I_27329 (I467125,I2507,I467026,I467151,);
not I_27330 (I467159,I467151);
DFFARX1 I_27331 (I934095,I2507,I467026,I467185,);
and I_27332 (I467193,I467185,I934086);
nand I_27333 (I467210,I467185,I934086);
nand I_27334 (I466997,I467159,I467210);
DFFARX1 I_27335 (I934101,I2507,I467026,I467250,);
nor I_27336 (I467258,I467250,I467193);
DFFARX1 I_27337 (I467258,I2507,I467026,I466991,);
nor I_27338 (I467006,I467250,I467151);
nand I_27339 (I467303,I934110,I934098);
and I_27340 (I467320,I467303,I934107);
DFFARX1 I_27341 (I467320,I2507,I467026,I467346,);
nor I_27342 (I466994,I467346,I467250);
not I_27343 (I467368,I467346);
nor I_27344 (I467385,I467368,I467159);
nor I_27345 (I467402,I467091,I467385);
DFFARX1 I_27346 (I467402,I2507,I467026,I467009,);
nor I_27347 (I467433,I467368,I467250);
nor I_27348 (I467450,I934083,I934098);
nor I_27349 (I467000,I467450,I467433);
not I_27350 (I467481,I467450);
nand I_27351 (I467003,I467210,I467481);
DFFARX1 I_27352 (I467450,I2507,I467026,I467015,);
DFFARX1 I_27353 (I467450,I2507,I467026,I467012,);
not I_27354 (I467570,I2514);
DFFARX1 I_27355 (I602977,I2507,I467570,I467596,);
DFFARX1 I_27356 (I467596,I2507,I467570,I467613,);
not I_27357 (I467562,I467613);
not I_27358 (I467635,I467596);
nand I_27359 (I467652,I602974,I602995);
and I_27360 (I467669,I467652,I602998);
DFFARX1 I_27361 (I467669,I2507,I467570,I467695,);
not I_27362 (I467703,I467695);
DFFARX1 I_27363 (I602983,I2507,I467570,I467729,);
and I_27364 (I467737,I467729,I602986);
nand I_27365 (I467754,I467729,I602986);
nand I_27366 (I467541,I467703,I467754);
DFFARX1 I_27367 (I602989,I2507,I467570,I467794,);
nor I_27368 (I467802,I467794,I467737);
DFFARX1 I_27369 (I467802,I2507,I467570,I467535,);
nor I_27370 (I467550,I467794,I467695);
nand I_27371 (I467847,I602974,I602980);
and I_27372 (I467864,I467847,I602992);
DFFARX1 I_27373 (I467864,I2507,I467570,I467890,);
nor I_27374 (I467538,I467890,I467794);
not I_27375 (I467912,I467890);
nor I_27376 (I467929,I467912,I467703);
nor I_27377 (I467946,I467635,I467929);
DFFARX1 I_27378 (I467946,I2507,I467570,I467553,);
nor I_27379 (I467977,I467912,I467794);
nor I_27380 (I467994,I602977,I602980);
nor I_27381 (I467544,I467994,I467977);
not I_27382 (I468025,I467994);
nand I_27383 (I467547,I467754,I468025);
DFFARX1 I_27384 (I467994,I2507,I467570,I467559,);
DFFARX1 I_27385 (I467994,I2507,I467570,I467556,);
not I_27386 (I468114,I2514);
DFFARX1 I_27387 (I1008379,I2507,I468114,I468140,);
DFFARX1 I_27388 (I468140,I2507,I468114,I468157,);
not I_27389 (I468106,I468157);
not I_27390 (I468179,I468140);
nand I_27391 (I468196,I1008394,I1008382);
and I_27392 (I468213,I468196,I1008373);
DFFARX1 I_27393 (I468213,I2507,I468114,I468239,);
not I_27394 (I468247,I468239);
DFFARX1 I_27395 (I1008385,I2507,I468114,I468273,);
and I_27396 (I468281,I468273,I1008376);
nand I_27397 (I468298,I468273,I1008376);
nand I_27398 (I468085,I468247,I468298);
DFFARX1 I_27399 (I1008391,I2507,I468114,I468338,);
nor I_27400 (I468346,I468338,I468281);
DFFARX1 I_27401 (I468346,I2507,I468114,I468079,);
nor I_27402 (I468094,I468338,I468239);
nand I_27403 (I468391,I1008400,I1008388);
and I_27404 (I468408,I468391,I1008397);
DFFARX1 I_27405 (I468408,I2507,I468114,I468434,);
nor I_27406 (I468082,I468434,I468338);
not I_27407 (I468456,I468434);
nor I_27408 (I468473,I468456,I468247);
nor I_27409 (I468490,I468179,I468473);
DFFARX1 I_27410 (I468490,I2507,I468114,I468097,);
nor I_27411 (I468521,I468456,I468338);
nor I_27412 (I468538,I1008373,I1008388);
nor I_27413 (I468088,I468538,I468521);
not I_27414 (I468569,I468538);
nand I_27415 (I468091,I468298,I468569);
DFFARX1 I_27416 (I468538,I2507,I468114,I468103,);
DFFARX1 I_27417 (I468538,I2507,I468114,I468100,);
not I_27418 (I468658,I2514);
DFFARX1 I_27419 (I967681,I2507,I468658,I468684,);
DFFARX1 I_27420 (I468684,I2507,I468658,I468701,);
not I_27421 (I468650,I468701);
not I_27422 (I468723,I468684);
nand I_27423 (I468740,I967696,I967684);
and I_27424 (I468757,I468740,I967675);
DFFARX1 I_27425 (I468757,I2507,I468658,I468783,);
not I_27426 (I468791,I468783);
DFFARX1 I_27427 (I967687,I2507,I468658,I468817,);
and I_27428 (I468825,I468817,I967678);
nand I_27429 (I468842,I468817,I967678);
nand I_27430 (I468629,I468791,I468842);
DFFARX1 I_27431 (I967693,I2507,I468658,I468882,);
nor I_27432 (I468890,I468882,I468825);
DFFARX1 I_27433 (I468890,I2507,I468658,I468623,);
nor I_27434 (I468638,I468882,I468783);
nand I_27435 (I468935,I967702,I967690);
and I_27436 (I468952,I468935,I967699);
DFFARX1 I_27437 (I468952,I2507,I468658,I468978,);
nor I_27438 (I468626,I468978,I468882);
not I_27439 (I469000,I468978);
nor I_27440 (I469017,I469000,I468791);
nor I_27441 (I469034,I468723,I469017);
DFFARX1 I_27442 (I469034,I2507,I468658,I468641,);
nor I_27443 (I469065,I469000,I468882);
nor I_27444 (I469082,I967675,I967690);
nor I_27445 (I468632,I469082,I469065);
not I_27446 (I469113,I469082);
nand I_27447 (I468635,I468842,I469113);
DFFARX1 I_27448 (I469082,I2507,I468658,I468647,);
DFFARX1 I_27449 (I469082,I2507,I468658,I468644,);
not I_27450 (I469202,I2514);
DFFARX1 I_27451 (I95972,I2507,I469202,I469228,);
DFFARX1 I_27452 (I469228,I2507,I469202,I469245,);
not I_27453 (I469194,I469245);
not I_27454 (I469267,I469228);
nand I_27455 (I469284,I95987,I95966);
and I_27456 (I469301,I469284,I95969);
DFFARX1 I_27457 (I469301,I2507,I469202,I469327,);
not I_27458 (I469335,I469327);
DFFARX1 I_27459 (I95975,I2507,I469202,I469361,);
and I_27460 (I469369,I469361,I95969);
nand I_27461 (I469386,I469361,I95969);
nand I_27462 (I469173,I469335,I469386);
DFFARX1 I_27463 (I95984,I2507,I469202,I469426,);
nor I_27464 (I469434,I469426,I469369);
DFFARX1 I_27465 (I469434,I2507,I469202,I469167,);
nor I_27466 (I469182,I469426,I469327);
nand I_27467 (I469479,I95966,I95981);
and I_27468 (I469496,I469479,I95978);
DFFARX1 I_27469 (I469496,I2507,I469202,I469522,);
nor I_27470 (I469170,I469522,I469426);
not I_27471 (I469544,I469522);
nor I_27472 (I469561,I469544,I469335);
nor I_27473 (I469578,I469267,I469561);
DFFARX1 I_27474 (I469578,I2507,I469202,I469185,);
nor I_27475 (I469609,I469544,I469426);
nor I_27476 (I469626,I95990,I95981);
nor I_27477 (I469176,I469626,I469609);
not I_27478 (I469657,I469626);
nand I_27479 (I469179,I469386,I469657);
DFFARX1 I_27480 (I469626,I2507,I469202,I469191,);
DFFARX1 I_27481 (I469626,I2507,I469202,I469188,);
not I_27482 (I469746,I2514);
DFFARX1 I_27483 (I319248,I2507,I469746,I469772,);
DFFARX1 I_27484 (I469772,I2507,I469746,I469789,);
not I_27485 (I469738,I469789);
not I_27486 (I469811,I469772);
nand I_27487 (I469828,I319227,I319251);
and I_27488 (I469845,I469828,I319254);
DFFARX1 I_27489 (I469845,I2507,I469746,I469871,);
not I_27490 (I469879,I469871);
DFFARX1 I_27491 (I319236,I2507,I469746,I469905,);
and I_27492 (I469913,I469905,I319242);
nand I_27493 (I469930,I469905,I319242);
nand I_27494 (I469717,I469879,I469930);
DFFARX1 I_27495 (I319230,I2507,I469746,I469970,);
nor I_27496 (I469978,I469970,I469913);
DFFARX1 I_27497 (I469978,I2507,I469746,I469711,);
nor I_27498 (I469726,I469970,I469871);
nand I_27499 (I470023,I319239,I319227);
and I_27500 (I470040,I470023,I319233);
DFFARX1 I_27501 (I470040,I2507,I469746,I470066,);
nor I_27502 (I469714,I470066,I469970);
not I_27503 (I470088,I470066);
nor I_27504 (I470105,I470088,I469879);
nor I_27505 (I470122,I469811,I470105);
DFFARX1 I_27506 (I470122,I2507,I469746,I469729,);
nor I_27507 (I470153,I470088,I469970);
nor I_27508 (I470170,I319245,I319227);
nor I_27509 (I469720,I470170,I470153);
not I_27510 (I470201,I470170);
nand I_27511 (I469723,I469930,I470201);
DFFARX1 I_27512 (I470170,I2507,I469746,I469735,);
DFFARX1 I_27513 (I470170,I2507,I469746,I469732,);
not I_27514 (I470290,I2514);
DFFARX1 I_27515 (I31684,I2507,I470290,I470316,);
DFFARX1 I_27516 (I470316,I2507,I470290,I470333,);
not I_27517 (I470282,I470333);
not I_27518 (I470355,I470316);
nand I_27519 (I470372,I31672,I31687);
and I_27520 (I470389,I470372,I31675);
DFFARX1 I_27521 (I470389,I2507,I470290,I470415,);
not I_27522 (I470423,I470415);
DFFARX1 I_27523 (I31696,I2507,I470290,I470449,);
and I_27524 (I470457,I470449,I31690);
nand I_27525 (I470474,I470449,I31690);
nand I_27526 (I470261,I470423,I470474);
DFFARX1 I_27527 (I31693,I2507,I470290,I470514,);
nor I_27528 (I470522,I470514,I470457);
DFFARX1 I_27529 (I470522,I2507,I470290,I470255,);
nor I_27530 (I470270,I470514,I470415);
nand I_27531 (I470567,I31672,I31675);
and I_27532 (I470584,I470567,I31678);
DFFARX1 I_27533 (I470584,I2507,I470290,I470610,);
nor I_27534 (I470258,I470610,I470514);
not I_27535 (I470632,I470610);
nor I_27536 (I470649,I470632,I470423);
nor I_27537 (I470666,I470355,I470649);
DFFARX1 I_27538 (I470666,I2507,I470290,I470273,);
nor I_27539 (I470697,I470632,I470514);
nor I_27540 (I470714,I31681,I31675);
nor I_27541 (I470264,I470714,I470697);
not I_27542 (I470745,I470714);
nand I_27543 (I470267,I470474,I470745);
DFFARX1 I_27544 (I470714,I2507,I470290,I470279,);
DFFARX1 I_27545 (I470714,I2507,I470290,I470276,);
not I_27546 (I470834,I2514);
DFFARX1 I_27547 (I33792,I2507,I470834,I470860,);
DFFARX1 I_27548 (I470860,I2507,I470834,I470877,);
not I_27549 (I470826,I470877);
not I_27550 (I470899,I470860);
nand I_27551 (I470916,I33780,I33795);
and I_27552 (I470933,I470916,I33783);
DFFARX1 I_27553 (I470933,I2507,I470834,I470959,);
not I_27554 (I470967,I470959);
DFFARX1 I_27555 (I33804,I2507,I470834,I470993,);
and I_27556 (I471001,I470993,I33798);
nand I_27557 (I471018,I470993,I33798);
nand I_27558 (I470805,I470967,I471018);
DFFARX1 I_27559 (I33801,I2507,I470834,I471058,);
nor I_27560 (I471066,I471058,I471001);
DFFARX1 I_27561 (I471066,I2507,I470834,I470799,);
nor I_27562 (I470814,I471058,I470959);
nand I_27563 (I471111,I33780,I33783);
and I_27564 (I471128,I471111,I33786);
DFFARX1 I_27565 (I471128,I2507,I470834,I471154,);
nor I_27566 (I470802,I471154,I471058);
not I_27567 (I471176,I471154);
nor I_27568 (I471193,I471176,I470967);
nor I_27569 (I471210,I470899,I471193);
DFFARX1 I_27570 (I471210,I2507,I470834,I470817,);
nor I_27571 (I471241,I471176,I471058);
nor I_27572 (I471258,I33789,I33783);
nor I_27573 (I470808,I471258,I471241);
not I_27574 (I471289,I471258);
nand I_27575 (I470811,I471018,I471289);
DFFARX1 I_27576 (I471258,I2507,I470834,I470823,);
DFFARX1 I_27577 (I471258,I2507,I470834,I470820,);
not I_27578 (I471378,I2514);
DFFARX1 I_27579 (I687365,I2507,I471378,I471404,);
DFFARX1 I_27580 (I471404,I2507,I471378,I471421,);
not I_27581 (I471370,I471421);
not I_27582 (I471443,I471404);
nand I_27583 (I471460,I687386,I687377);
and I_27584 (I471477,I471460,I687365);
DFFARX1 I_27585 (I471477,I2507,I471378,I471503,);
not I_27586 (I471511,I471503);
DFFARX1 I_27587 (I687371,I2507,I471378,I471537,);
and I_27588 (I471545,I471537,I687368);
nand I_27589 (I471562,I471537,I687368);
nand I_27590 (I471349,I471511,I471562);
DFFARX1 I_27591 (I687362,I2507,I471378,I471602,);
nor I_27592 (I471610,I471602,I471545);
DFFARX1 I_27593 (I471610,I2507,I471378,I471343,);
nor I_27594 (I471358,I471602,I471503);
nand I_27595 (I471655,I687362,I687374);
and I_27596 (I471672,I471655,I687383);
DFFARX1 I_27597 (I471672,I2507,I471378,I471698,);
nor I_27598 (I471346,I471698,I471602);
not I_27599 (I471720,I471698);
nor I_27600 (I471737,I471720,I471511);
nor I_27601 (I471754,I471443,I471737);
DFFARX1 I_27602 (I471754,I2507,I471378,I471361,);
nor I_27603 (I471785,I471720,I471602);
nor I_27604 (I471802,I687380,I687374);
nor I_27605 (I471352,I471802,I471785);
not I_27606 (I471833,I471802);
nand I_27607 (I471355,I471562,I471833);
DFFARX1 I_27608 (I471802,I2507,I471378,I471367,);
DFFARX1 I_27609 (I471802,I2507,I471378,I471364,);
not I_27610 (I471922,I2514);
DFFARX1 I_27611 (I263386,I2507,I471922,I471948,);
DFFARX1 I_27612 (I471948,I2507,I471922,I471965,);
not I_27613 (I471914,I471965);
not I_27614 (I471987,I471948);
nand I_27615 (I472004,I263365,I263389);
and I_27616 (I472021,I472004,I263392);
DFFARX1 I_27617 (I472021,I2507,I471922,I472047,);
not I_27618 (I472055,I472047);
DFFARX1 I_27619 (I263374,I2507,I471922,I472081,);
and I_27620 (I472089,I472081,I263380);
nand I_27621 (I472106,I472081,I263380);
nand I_27622 (I471893,I472055,I472106);
DFFARX1 I_27623 (I263368,I2507,I471922,I472146,);
nor I_27624 (I472154,I472146,I472089);
DFFARX1 I_27625 (I472154,I2507,I471922,I471887,);
nor I_27626 (I471902,I472146,I472047);
nand I_27627 (I472199,I263377,I263365);
and I_27628 (I472216,I472199,I263371);
DFFARX1 I_27629 (I472216,I2507,I471922,I472242,);
nor I_27630 (I471890,I472242,I472146);
not I_27631 (I472264,I472242);
nor I_27632 (I472281,I472264,I472055);
nor I_27633 (I472298,I471987,I472281);
DFFARX1 I_27634 (I472298,I2507,I471922,I471905,);
nor I_27635 (I472329,I472264,I472146);
nor I_27636 (I472346,I263383,I263365);
nor I_27637 (I471896,I472346,I472329);
not I_27638 (I472377,I472346);
nand I_27639 (I471899,I472106,I472377);
DFFARX1 I_27640 (I472346,I2507,I471922,I471911,);
DFFARX1 I_27641 (I472346,I2507,I471922,I471908,);
not I_27642 (I472466,I2514);
DFFARX1 I_27643 (I1283094,I2507,I472466,I472492,);
DFFARX1 I_27644 (I472492,I2507,I472466,I472509,);
not I_27645 (I472458,I472509);
not I_27646 (I472531,I472492);
nand I_27647 (I472548,I1283091,I1283088);
and I_27648 (I472565,I472548,I1283076);
DFFARX1 I_27649 (I472565,I2507,I472466,I472591,);
not I_27650 (I472599,I472591);
DFFARX1 I_27651 (I1283100,I2507,I472466,I472625,);
and I_27652 (I472633,I472625,I1283085);
nand I_27653 (I472650,I472625,I1283085);
nand I_27654 (I472437,I472599,I472650);
DFFARX1 I_27655 (I1283079,I2507,I472466,I472690,);
nor I_27656 (I472698,I472690,I472633);
DFFARX1 I_27657 (I472698,I2507,I472466,I472431,);
nor I_27658 (I472446,I472690,I472591);
nand I_27659 (I472743,I1283076,I1283082);
and I_27660 (I472760,I472743,I1283097);
DFFARX1 I_27661 (I472760,I2507,I472466,I472786,);
nor I_27662 (I472434,I472786,I472690);
not I_27663 (I472808,I472786);
nor I_27664 (I472825,I472808,I472599);
nor I_27665 (I472842,I472531,I472825);
DFFARX1 I_27666 (I472842,I2507,I472466,I472449,);
nor I_27667 (I472873,I472808,I472690);
nor I_27668 (I472890,I1283079,I1283082);
nor I_27669 (I472440,I472890,I472873);
not I_27670 (I472921,I472890);
nand I_27671 (I472443,I472650,I472921);
DFFARX1 I_27672 (I472890,I2507,I472466,I472455,);
DFFARX1 I_27673 (I472890,I2507,I472466,I472452,);
not I_27674 (I473010,I2514);
DFFARX1 I_27675 (I996105,I2507,I473010,I473036,);
DFFARX1 I_27676 (I473036,I2507,I473010,I473053,);
not I_27677 (I473002,I473053);
not I_27678 (I473075,I473036);
nand I_27679 (I473092,I996120,I996108);
and I_27680 (I473109,I473092,I996099);
DFFARX1 I_27681 (I473109,I2507,I473010,I473135,);
not I_27682 (I473143,I473135);
DFFARX1 I_27683 (I996111,I2507,I473010,I473169,);
and I_27684 (I473177,I473169,I996102);
nand I_27685 (I473194,I473169,I996102);
nand I_27686 (I472981,I473143,I473194);
DFFARX1 I_27687 (I996117,I2507,I473010,I473234,);
nor I_27688 (I473242,I473234,I473177);
DFFARX1 I_27689 (I473242,I2507,I473010,I472975,);
nor I_27690 (I472990,I473234,I473135);
nand I_27691 (I473287,I996126,I996114);
and I_27692 (I473304,I473287,I996123);
DFFARX1 I_27693 (I473304,I2507,I473010,I473330,);
nor I_27694 (I472978,I473330,I473234);
not I_27695 (I473352,I473330);
nor I_27696 (I473369,I473352,I473143);
nor I_27697 (I473386,I473075,I473369);
DFFARX1 I_27698 (I473386,I2507,I473010,I472993,);
nor I_27699 (I473417,I473352,I473234);
nor I_27700 (I473434,I996099,I996114);
nor I_27701 (I472984,I473434,I473417);
not I_27702 (I473465,I473434);
nand I_27703 (I472987,I473194,I473465);
DFFARX1 I_27704 (I473434,I2507,I473010,I472999,);
DFFARX1 I_27705 (I473434,I2507,I473010,I472996,);
not I_27706 (I473554,I2514);
DFFARX1 I_27707 (I934735,I2507,I473554,I473580,);
DFFARX1 I_27708 (I473580,I2507,I473554,I473597,);
not I_27709 (I473546,I473597);
not I_27710 (I473619,I473580);
nand I_27711 (I473636,I934750,I934738);
and I_27712 (I473653,I473636,I934729);
DFFARX1 I_27713 (I473653,I2507,I473554,I473679,);
not I_27714 (I473687,I473679);
DFFARX1 I_27715 (I934741,I2507,I473554,I473713,);
and I_27716 (I473721,I473713,I934732);
nand I_27717 (I473738,I473713,I934732);
nand I_27718 (I473525,I473687,I473738);
DFFARX1 I_27719 (I934747,I2507,I473554,I473778,);
nor I_27720 (I473786,I473778,I473721);
DFFARX1 I_27721 (I473786,I2507,I473554,I473519,);
nor I_27722 (I473534,I473778,I473679);
nand I_27723 (I473831,I934756,I934744);
and I_27724 (I473848,I473831,I934753);
DFFARX1 I_27725 (I473848,I2507,I473554,I473874,);
nor I_27726 (I473522,I473874,I473778);
not I_27727 (I473896,I473874);
nor I_27728 (I473913,I473896,I473687);
nor I_27729 (I473930,I473619,I473913);
DFFARX1 I_27730 (I473930,I2507,I473554,I473537,);
nor I_27731 (I473961,I473896,I473778);
nor I_27732 (I473978,I934729,I934744);
nor I_27733 (I473528,I473978,I473961);
not I_27734 (I474009,I473978);
nand I_27735 (I473531,I473738,I474009);
DFFARX1 I_27736 (I473978,I2507,I473554,I473543,);
DFFARX1 I_27737 (I473978,I2507,I473554,I473540,);
not I_27738 (I474098,I2514);
DFFARX1 I_27739 (I267075,I2507,I474098,I474124,);
DFFARX1 I_27740 (I474124,I2507,I474098,I474141,);
not I_27741 (I474090,I474141);
not I_27742 (I474163,I474124);
nand I_27743 (I474180,I267054,I267078);
and I_27744 (I474197,I474180,I267081);
DFFARX1 I_27745 (I474197,I2507,I474098,I474223,);
not I_27746 (I474231,I474223);
DFFARX1 I_27747 (I267063,I2507,I474098,I474257,);
and I_27748 (I474265,I474257,I267069);
nand I_27749 (I474282,I474257,I267069);
nand I_27750 (I474069,I474231,I474282);
DFFARX1 I_27751 (I267057,I2507,I474098,I474322,);
nor I_27752 (I474330,I474322,I474265);
DFFARX1 I_27753 (I474330,I2507,I474098,I474063,);
nor I_27754 (I474078,I474322,I474223);
nand I_27755 (I474375,I267066,I267054);
and I_27756 (I474392,I474375,I267060);
DFFARX1 I_27757 (I474392,I2507,I474098,I474418,);
nor I_27758 (I474066,I474418,I474322);
not I_27759 (I474440,I474418);
nor I_27760 (I474457,I474440,I474231);
nor I_27761 (I474474,I474163,I474457);
DFFARX1 I_27762 (I474474,I2507,I474098,I474081,);
nor I_27763 (I474505,I474440,I474322);
nor I_27764 (I474522,I267072,I267054);
nor I_27765 (I474072,I474522,I474505);
not I_27766 (I474553,I474522);
nand I_27767 (I474075,I474282,I474553);
DFFARX1 I_27768 (I474522,I2507,I474098,I474087,);
DFFARX1 I_27769 (I474522,I2507,I474098,I474084,);
not I_27770 (I474642,I2514);
DFFARX1 I_27771 (I1096521,I2507,I474642,I474668,);
DFFARX1 I_27772 (I474668,I2507,I474642,I474685,);
not I_27773 (I474634,I474685);
not I_27774 (I474707,I474668);
nand I_27775 (I474724,I1096533,I1096521);
and I_27776 (I474741,I474724,I1096524);
DFFARX1 I_27777 (I474741,I2507,I474642,I474767,);
not I_27778 (I474775,I474767);
DFFARX1 I_27779 (I1096542,I2507,I474642,I474801,);
and I_27780 (I474809,I474801,I1096518);
nand I_27781 (I474826,I474801,I1096518);
nand I_27782 (I474613,I474775,I474826);
DFFARX1 I_27783 (I1096536,I2507,I474642,I474866,);
nor I_27784 (I474874,I474866,I474809);
DFFARX1 I_27785 (I474874,I2507,I474642,I474607,);
nor I_27786 (I474622,I474866,I474767);
nand I_27787 (I474919,I1096530,I1096527);
and I_27788 (I474936,I474919,I1096539);
DFFARX1 I_27789 (I474936,I2507,I474642,I474962,);
nor I_27790 (I474610,I474962,I474866);
not I_27791 (I474984,I474962);
nor I_27792 (I475001,I474984,I474775);
nor I_27793 (I475018,I474707,I475001);
DFFARX1 I_27794 (I475018,I2507,I474642,I474625,);
nor I_27795 (I475049,I474984,I474866);
nor I_27796 (I475066,I1096518,I1096527);
nor I_27797 (I474616,I475066,I475049);
not I_27798 (I475097,I475066);
nand I_27799 (I474619,I474826,I475097);
DFFARX1 I_27800 (I475066,I2507,I474642,I474631,);
DFFARX1 I_27801 (I475066,I2507,I474642,I474628,);
not I_27802 (I475186,I2514);
DFFARX1 I_27803 (I1230821,I2507,I475186,I475212,);
DFFARX1 I_27804 (I475212,I2507,I475186,I475229,);
not I_27805 (I475178,I475229);
not I_27806 (I475251,I475212);
nand I_27807 (I475268,I1230833,I1230836);
and I_27808 (I475285,I475268,I1230839);
DFFARX1 I_27809 (I475285,I2507,I475186,I475311,);
not I_27810 (I475319,I475311);
DFFARX1 I_27811 (I1230824,I2507,I475186,I475345,);
and I_27812 (I475353,I475345,I1230830);
nand I_27813 (I475370,I475345,I1230830);
nand I_27814 (I475157,I475319,I475370);
DFFARX1 I_27815 (I1230818,I2507,I475186,I475410,);
nor I_27816 (I475418,I475410,I475353);
DFFARX1 I_27817 (I475418,I2507,I475186,I475151,);
nor I_27818 (I475166,I475410,I475311);
nand I_27819 (I475463,I1230821,I1230842);
and I_27820 (I475480,I475463,I1230827);
DFFARX1 I_27821 (I475480,I2507,I475186,I475506,);
nor I_27822 (I475154,I475506,I475410);
not I_27823 (I475528,I475506);
nor I_27824 (I475545,I475528,I475319);
nor I_27825 (I475562,I475251,I475545);
DFFARX1 I_27826 (I475562,I2507,I475186,I475169,);
nor I_27827 (I475593,I475528,I475410);
nor I_27828 (I475610,I1230818,I1230842);
nor I_27829 (I475160,I475610,I475593);
not I_27830 (I475641,I475610);
nand I_27831 (I475163,I475370,I475641);
DFFARX1 I_27832 (I475610,I2507,I475186,I475175,);
DFFARX1 I_27833 (I475610,I2507,I475186,I475172,);
not I_27834 (I475730,I2514);
DFFARX1 I_27835 (I78581,I2507,I475730,I475756,);
DFFARX1 I_27836 (I475756,I2507,I475730,I475773,);
not I_27837 (I475722,I475773);
not I_27838 (I475795,I475756);
nand I_27839 (I475812,I78596,I78575);
and I_27840 (I475829,I475812,I78578);
DFFARX1 I_27841 (I475829,I2507,I475730,I475855,);
not I_27842 (I475863,I475855);
DFFARX1 I_27843 (I78584,I2507,I475730,I475889,);
and I_27844 (I475897,I475889,I78578);
nand I_27845 (I475914,I475889,I78578);
nand I_27846 (I475701,I475863,I475914);
DFFARX1 I_27847 (I78593,I2507,I475730,I475954,);
nor I_27848 (I475962,I475954,I475897);
DFFARX1 I_27849 (I475962,I2507,I475730,I475695,);
nor I_27850 (I475710,I475954,I475855);
nand I_27851 (I476007,I78575,I78590);
and I_27852 (I476024,I476007,I78587);
DFFARX1 I_27853 (I476024,I2507,I475730,I476050,);
nor I_27854 (I475698,I476050,I475954);
not I_27855 (I476072,I476050);
nor I_27856 (I476089,I476072,I475863);
nor I_27857 (I476106,I475795,I476089);
DFFARX1 I_27858 (I476106,I2507,I475730,I475713,);
nor I_27859 (I476137,I476072,I475954);
nor I_27860 (I476154,I78599,I78590);
nor I_27861 (I475704,I476154,I476137);
not I_27862 (I476185,I476154);
nand I_27863 (I475707,I475914,I476185);
DFFARX1 I_27864 (I476154,I2507,I475730,I475719,);
DFFARX1 I_27865 (I476154,I2507,I475730,I475716,);
not I_27866 (I476274,I2514);
DFFARX1 I_27867 (I1287718,I2507,I476274,I476300,);
DFFARX1 I_27868 (I476300,I2507,I476274,I476317,);
not I_27869 (I476266,I476317);
not I_27870 (I476339,I476300);
nand I_27871 (I476356,I1287715,I1287712);
and I_27872 (I476373,I476356,I1287700);
DFFARX1 I_27873 (I476373,I2507,I476274,I476399,);
not I_27874 (I476407,I476399);
DFFARX1 I_27875 (I1287724,I2507,I476274,I476433,);
and I_27876 (I476441,I476433,I1287709);
nand I_27877 (I476458,I476433,I1287709);
nand I_27878 (I476245,I476407,I476458);
DFFARX1 I_27879 (I1287703,I2507,I476274,I476498,);
nor I_27880 (I476506,I476498,I476441);
DFFARX1 I_27881 (I476506,I2507,I476274,I476239,);
nor I_27882 (I476254,I476498,I476399);
nand I_27883 (I476551,I1287700,I1287706);
and I_27884 (I476568,I476551,I1287721);
DFFARX1 I_27885 (I476568,I2507,I476274,I476594,);
nor I_27886 (I476242,I476594,I476498);
not I_27887 (I476616,I476594);
nor I_27888 (I476633,I476616,I476407);
nor I_27889 (I476650,I476339,I476633);
DFFARX1 I_27890 (I476650,I2507,I476274,I476257,);
nor I_27891 (I476681,I476616,I476498);
nor I_27892 (I476698,I1287703,I1287706);
nor I_27893 (I476248,I476698,I476681);
not I_27894 (I476729,I476698);
nand I_27895 (I476251,I476458,I476729);
DFFARX1 I_27896 (I476698,I2507,I476274,I476263,);
DFFARX1 I_27897 (I476698,I2507,I476274,I476260,);
not I_27898 (I476818,I2514);
DFFARX1 I_27899 (I352976,I2507,I476818,I476844,);
DFFARX1 I_27900 (I476844,I2507,I476818,I476861,);
not I_27901 (I476810,I476861);
not I_27902 (I476883,I476844);
nand I_27903 (I476900,I352955,I352979);
and I_27904 (I476917,I476900,I352982);
DFFARX1 I_27905 (I476917,I2507,I476818,I476943,);
not I_27906 (I476951,I476943);
DFFARX1 I_27907 (I352964,I2507,I476818,I476977,);
and I_27908 (I476985,I476977,I352970);
nand I_27909 (I477002,I476977,I352970);
nand I_27910 (I476789,I476951,I477002);
DFFARX1 I_27911 (I352958,I2507,I476818,I477042,);
nor I_27912 (I477050,I477042,I476985);
DFFARX1 I_27913 (I477050,I2507,I476818,I476783,);
nor I_27914 (I476798,I477042,I476943);
nand I_27915 (I477095,I352967,I352955);
and I_27916 (I477112,I477095,I352961);
DFFARX1 I_27917 (I477112,I2507,I476818,I477138,);
nor I_27918 (I476786,I477138,I477042);
not I_27919 (I477160,I477138);
nor I_27920 (I477177,I477160,I476951);
nor I_27921 (I477194,I476883,I477177);
DFFARX1 I_27922 (I477194,I2507,I476818,I476801,);
nor I_27923 (I477225,I477160,I477042);
nor I_27924 (I477242,I352973,I352955);
nor I_27925 (I476792,I477242,I477225);
not I_27926 (I477273,I477242);
nand I_27927 (I476795,I477002,I477273);
DFFARX1 I_27928 (I477242,I2507,I476818,I476807,);
DFFARX1 I_27929 (I477242,I2507,I476818,I476804,);
not I_27930 (I477362,I2514);
DFFARX1 I_27931 (I287628,I2507,I477362,I477388,);
DFFARX1 I_27932 (I477388,I2507,I477362,I477405,);
not I_27933 (I477354,I477405);
not I_27934 (I477427,I477388);
nand I_27935 (I477444,I287607,I287631);
and I_27936 (I477461,I477444,I287634);
DFFARX1 I_27937 (I477461,I2507,I477362,I477487,);
not I_27938 (I477495,I477487);
DFFARX1 I_27939 (I287616,I2507,I477362,I477521,);
and I_27940 (I477529,I477521,I287622);
nand I_27941 (I477546,I477521,I287622);
nand I_27942 (I477333,I477495,I477546);
DFFARX1 I_27943 (I287610,I2507,I477362,I477586,);
nor I_27944 (I477594,I477586,I477529);
DFFARX1 I_27945 (I477594,I2507,I477362,I477327,);
nor I_27946 (I477342,I477586,I477487);
nand I_27947 (I477639,I287619,I287607);
and I_27948 (I477656,I477639,I287613);
DFFARX1 I_27949 (I477656,I2507,I477362,I477682,);
nor I_27950 (I477330,I477682,I477586);
not I_27951 (I477704,I477682);
nor I_27952 (I477721,I477704,I477495);
nor I_27953 (I477738,I477427,I477721);
DFFARX1 I_27954 (I477738,I2507,I477362,I477345,);
nor I_27955 (I477769,I477704,I477586);
nor I_27956 (I477786,I287625,I287607);
nor I_27957 (I477336,I477786,I477769);
not I_27958 (I477817,I477786);
nand I_27959 (I477339,I477546,I477817);
DFFARX1 I_27960 (I477786,I2507,I477362,I477351,);
DFFARX1 I_27961 (I477786,I2507,I477362,I477348,);
not I_27962 (I477906,I2514);
DFFARX1 I_27963 (I829664,I2507,I477906,I477932,);
DFFARX1 I_27964 (I477932,I2507,I477906,I477949,);
not I_27965 (I477898,I477949);
not I_27966 (I477971,I477932);
nand I_27967 (I477988,I829658,I829655);
and I_27968 (I478005,I477988,I829670);
DFFARX1 I_27969 (I478005,I2507,I477906,I478031,);
not I_27970 (I478039,I478031);
DFFARX1 I_27971 (I829658,I2507,I477906,I478065,);
and I_27972 (I478073,I478065,I829652);
nand I_27973 (I478090,I478065,I829652);
nand I_27974 (I477877,I478039,I478090);
DFFARX1 I_27975 (I829652,I2507,I477906,I478130,);
nor I_27976 (I478138,I478130,I478073);
DFFARX1 I_27977 (I478138,I2507,I477906,I477871,);
nor I_27978 (I477886,I478130,I478031);
nand I_27979 (I478183,I829667,I829661);
and I_27980 (I478200,I478183,I829655);
DFFARX1 I_27981 (I478200,I2507,I477906,I478226,);
nor I_27982 (I477874,I478226,I478130);
not I_27983 (I478248,I478226);
nor I_27984 (I478265,I478248,I478039);
nor I_27985 (I478282,I477971,I478265);
DFFARX1 I_27986 (I478282,I2507,I477906,I477889,);
nor I_27987 (I478313,I478248,I478130);
nor I_27988 (I478330,I829673,I829661);
nor I_27989 (I477880,I478330,I478313);
not I_27990 (I478361,I478330);
nand I_27991 (I477883,I478090,I478361);
DFFARX1 I_27992 (I478330,I2507,I477906,I477895,);
DFFARX1 I_27993 (I478330,I2507,I477906,I477892,);
not I_27994 (I478450,I2514);
DFFARX1 I_27995 (I1106925,I2507,I478450,I478476,);
DFFARX1 I_27996 (I478476,I2507,I478450,I478493,);
not I_27997 (I478442,I478493);
not I_27998 (I478515,I478476);
nand I_27999 (I478532,I1106937,I1106925);
and I_28000 (I478549,I478532,I1106928);
DFFARX1 I_28001 (I478549,I2507,I478450,I478575,);
not I_28002 (I478583,I478575);
DFFARX1 I_28003 (I1106946,I2507,I478450,I478609,);
and I_28004 (I478617,I478609,I1106922);
nand I_28005 (I478634,I478609,I1106922);
nand I_28006 (I478421,I478583,I478634);
DFFARX1 I_28007 (I1106940,I2507,I478450,I478674,);
nor I_28008 (I478682,I478674,I478617);
DFFARX1 I_28009 (I478682,I2507,I478450,I478415,);
nor I_28010 (I478430,I478674,I478575);
nand I_28011 (I478727,I1106934,I1106931);
and I_28012 (I478744,I478727,I1106943);
DFFARX1 I_28013 (I478744,I2507,I478450,I478770,);
nor I_28014 (I478418,I478770,I478674);
not I_28015 (I478792,I478770);
nor I_28016 (I478809,I478792,I478583);
nor I_28017 (I478826,I478515,I478809);
DFFARX1 I_28018 (I478826,I2507,I478450,I478433,);
nor I_28019 (I478857,I478792,I478674);
nor I_28020 (I478874,I1106922,I1106931);
nor I_28021 (I478424,I478874,I478857);
not I_28022 (I478905,I478874);
nand I_28023 (I478427,I478634,I478905);
DFFARX1 I_28024 (I478874,I2507,I478450,I478439,);
DFFARX1 I_28025 (I478874,I2507,I478450,I478436,);
not I_28026 (I478994,I2514);
DFFARX1 I_28027 (I1120219,I2507,I478994,I479020,);
DFFARX1 I_28028 (I479020,I2507,I478994,I479037,);
not I_28029 (I478986,I479037);
not I_28030 (I479059,I479020);
nand I_28031 (I479076,I1120231,I1120219);
and I_28032 (I479093,I479076,I1120222);
DFFARX1 I_28033 (I479093,I2507,I478994,I479119,);
not I_28034 (I479127,I479119);
DFFARX1 I_28035 (I1120240,I2507,I478994,I479153,);
and I_28036 (I479161,I479153,I1120216);
nand I_28037 (I479178,I479153,I1120216);
nand I_28038 (I478965,I479127,I479178);
DFFARX1 I_28039 (I1120234,I2507,I478994,I479218,);
nor I_28040 (I479226,I479218,I479161);
DFFARX1 I_28041 (I479226,I2507,I478994,I478959,);
nor I_28042 (I478974,I479218,I479119);
nand I_28043 (I479271,I1120228,I1120225);
and I_28044 (I479288,I479271,I1120237);
DFFARX1 I_28045 (I479288,I2507,I478994,I479314,);
nor I_28046 (I478962,I479314,I479218);
not I_28047 (I479336,I479314);
nor I_28048 (I479353,I479336,I479127);
nor I_28049 (I479370,I479059,I479353);
DFFARX1 I_28050 (I479370,I2507,I478994,I478977,);
nor I_28051 (I479401,I479336,I479218);
nor I_28052 (I479418,I1120216,I1120225);
nor I_28053 (I478968,I479418,I479401);
not I_28054 (I479449,I479418);
nand I_28055 (I478971,I479178,I479449);
DFFARX1 I_28056 (I479418,I2507,I478994,I478983,);
DFFARX1 I_28057 (I479418,I2507,I478994,I478980,);
not I_28058 (I479538,I2514);
DFFARX1 I_28059 (I16928,I2507,I479538,I479564,);
DFFARX1 I_28060 (I479564,I2507,I479538,I479581,);
not I_28061 (I479530,I479581);
not I_28062 (I479603,I479564);
nand I_28063 (I479620,I16916,I16931);
and I_28064 (I479637,I479620,I16919);
DFFARX1 I_28065 (I479637,I2507,I479538,I479663,);
not I_28066 (I479671,I479663);
DFFARX1 I_28067 (I16940,I2507,I479538,I479697,);
and I_28068 (I479705,I479697,I16934);
nand I_28069 (I479722,I479697,I16934);
nand I_28070 (I479509,I479671,I479722);
DFFARX1 I_28071 (I16937,I2507,I479538,I479762,);
nor I_28072 (I479770,I479762,I479705);
DFFARX1 I_28073 (I479770,I2507,I479538,I479503,);
nor I_28074 (I479518,I479762,I479663);
nand I_28075 (I479815,I16916,I16919);
and I_28076 (I479832,I479815,I16922);
DFFARX1 I_28077 (I479832,I2507,I479538,I479858,);
nor I_28078 (I479506,I479858,I479762);
not I_28079 (I479880,I479858);
nor I_28080 (I479897,I479880,I479671);
nor I_28081 (I479914,I479603,I479897);
DFFARX1 I_28082 (I479914,I2507,I479538,I479521,);
nor I_28083 (I479945,I479880,I479762);
nor I_28084 (I479962,I16925,I16919);
nor I_28085 (I479512,I479962,I479945);
not I_28086 (I479993,I479962);
nand I_28087 (I479515,I479722,I479993);
DFFARX1 I_28088 (I479962,I2507,I479538,I479527,);
DFFARX1 I_28089 (I479962,I2507,I479538,I479524,);
not I_28090 (I480082,I2514);
DFFARX1 I_28091 (I542287,I2507,I480082,I480108,);
DFFARX1 I_28092 (I480108,I2507,I480082,I480125,);
not I_28093 (I480074,I480125);
not I_28094 (I480147,I480108);
nand I_28095 (I480164,I542284,I542305);
and I_28096 (I480181,I480164,I542308);
DFFARX1 I_28097 (I480181,I2507,I480082,I480207,);
not I_28098 (I480215,I480207);
DFFARX1 I_28099 (I542293,I2507,I480082,I480241,);
and I_28100 (I480249,I480241,I542296);
nand I_28101 (I480266,I480241,I542296);
nand I_28102 (I480053,I480215,I480266);
DFFARX1 I_28103 (I542299,I2507,I480082,I480306,);
nor I_28104 (I480314,I480306,I480249);
DFFARX1 I_28105 (I480314,I2507,I480082,I480047,);
nor I_28106 (I480062,I480306,I480207);
nand I_28107 (I480359,I542284,I542290);
and I_28108 (I480376,I480359,I542302);
DFFARX1 I_28109 (I480376,I2507,I480082,I480402,);
nor I_28110 (I480050,I480402,I480306);
not I_28111 (I480424,I480402);
nor I_28112 (I480441,I480424,I480215);
nor I_28113 (I480458,I480147,I480441);
DFFARX1 I_28114 (I480458,I2507,I480082,I480065,);
nor I_28115 (I480489,I480424,I480306);
nor I_28116 (I480506,I542287,I542290);
nor I_28117 (I480056,I480506,I480489);
not I_28118 (I480537,I480506);
nand I_28119 (I480059,I480266,I480537);
DFFARX1 I_28120 (I480506,I2507,I480082,I480071,);
DFFARX1 I_28121 (I480506,I2507,I480082,I480068,);
not I_28122 (I480626,I2514);
DFFARX1 I_28123 (I916647,I2507,I480626,I480652,);
DFFARX1 I_28124 (I480652,I2507,I480626,I480669,);
not I_28125 (I480618,I480669);
not I_28126 (I480691,I480652);
nand I_28127 (I480708,I916662,I916650);
and I_28128 (I480725,I480708,I916641);
DFFARX1 I_28129 (I480725,I2507,I480626,I480751,);
not I_28130 (I480759,I480751);
DFFARX1 I_28131 (I916653,I2507,I480626,I480785,);
and I_28132 (I480793,I480785,I916644);
nand I_28133 (I480810,I480785,I916644);
nand I_28134 (I480597,I480759,I480810);
DFFARX1 I_28135 (I916659,I2507,I480626,I480850,);
nor I_28136 (I480858,I480850,I480793);
DFFARX1 I_28137 (I480858,I2507,I480626,I480591,);
nor I_28138 (I480606,I480850,I480751);
nand I_28139 (I480903,I916668,I916656);
and I_28140 (I480920,I480903,I916665);
DFFARX1 I_28141 (I480920,I2507,I480626,I480946,);
nor I_28142 (I480594,I480946,I480850);
not I_28143 (I480968,I480946);
nor I_28144 (I480985,I480968,I480759);
nor I_28145 (I481002,I480691,I480985);
DFFARX1 I_28146 (I481002,I2507,I480626,I480609,);
nor I_28147 (I481033,I480968,I480850);
nor I_28148 (I481050,I916641,I916656);
nor I_28149 (I480600,I481050,I481033);
not I_28150 (I481081,I481050);
nand I_28151 (I480603,I480810,I481081);
DFFARX1 I_28152 (I481050,I2507,I480626,I480615,);
DFFARX1 I_28153 (I481050,I2507,I480626,I480612,);
not I_28154 (I481170,I2514);
DFFARX1 I_28155 (I963159,I2507,I481170,I481196,);
DFFARX1 I_28156 (I481196,I2507,I481170,I481213,);
not I_28157 (I481162,I481213);
not I_28158 (I481235,I481196);
nand I_28159 (I481252,I963174,I963162);
and I_28160 (I481269,I481252,I963153);
DFFARX1 I_28161 (I481269,I2507,I481170,I481295,);
not I_28162 (I481303,I481295);
DFFARX1 I_28163 (I963165,I2507,I481170,I481329,);
and I_28164 (I481337,I481329,I963156);
nand I_28165 (I481354,I481329,I963156);
nand I_28166 (I481141,I481303,I481354);
DFFARX1 I_28167 (I963171,I2507,I481170,I481394,);
nor I_28168 (I481402,I481394,I481337);
DFFARX1 I_28169 (I481402,I2507,I481170,I481135,);
nor I_28170 (I481150,I481394,I481295);
nand I_28171 (I481447,I963180,I963168);
and I_28172 (I481464,I481447,I963177);
DFFARX1 I_28173 (I481464,I2507,I481170,I481490,);
nor I_28174 (I481138,I481490,I481394);
not I_28175 (I481512,I481490);
nor I_28176 (I481529,I481512,I481303);
nor I_28177 (I481546,I481235,I481529);
DFFARX1 I_28178 (I481546,I2507,I481170,I481153,);
nor I_28179 (I481577,I481512,I481394);
nor I_28180 (I481594,I963153,I963168);
nor I_28181 (I481144,I481594,I481577);
not I_28182 (I481625,I481594);
nand I_28183 (I481147,I481354,I481625);
DFFARX1 I_28184 (I481594,I2507,I481170,I481159,);
DFFARX1 I_28185 (I481594,I2507,I481170,I481156,);
not I_28186 (I481714,I2514);
DFFARX1 I_28187 (I1260552,I2507,I481714,I481740,);
DFFARX1 I_28188 (I481740,I2507,I481714,I481757,);
not I_28189 (I481706,I481757);
not I_28190 (I481779,I481740);
nand I_28191 (I481796,I1260549,I1260546);
and I_28192 (I481813,I481796,I1260534);
DFFARX1 I_28193 (I481813,I2507,I481714,I481839,);
not I_28194 (I481847,I481839);
DFFARX1 I_28195 (I1260558,I2507,I481714,I481873,);
and I_28196 (I481881,I481873,I1260543);
nand I_28197 (I481898,I481873,I1260543);
nand I_28198 (I481685,I481847,I481898);
DFFARX1 I_28199 (I1260537,I2507,I481714,I481938,);
nor I_28200 (I481946,I481938,I481881);
DFFARX1 I_28201 (I481946,I2507,I481714,I481679,);
nor I_28202 (I481694,I481938,I481839);
nand I_28203 (I481991,I1260534,I1260540);
and I_28204 (I482008,I481991,I1260555);
DFFARX1 I_28205 (I482008,I2507,I481714,I482034,);
nor I_28206 (I481682,I482034,I481938);
not I_28207 (I482056,I482034);
nor I_28208 (I482073,I482056,I481847);
nor I_28209 (I482090,I481779,I482073);
DFFARX1 I_28210 (I482090,I2507,I481714,I481697,);
nor I_28211 (I482121,I482056,I481938);
nor I_28212 (I482138,I1260537,I1260540);
nor I_28213 (I481688,I482138,I482121);
not I_28214 (I482169,I482138);
nand I_28215 (I481691,I481898,I482169);
DFFARX1 I_28216 (I482138,I2507,I481714,I481703,);
DFFARX1 I_28217 (I482138,I2507,I481714,I481700,);
not I_28218 (I482258,I2514);
DFFARX1 I_28219 (I301330,I2507,I482258,I482284,);
DFFARX1 I_28220 (I482284,I2507,I482258,I482301,);
not I_28221 (I482250,I482301);
not I_28222 (I482323,I482284);
nand I_28223 (I482340,I301309,I301333);
and I_28224 (I482357,I482340,I301336);
DFFARX1 I_28225 (I482357,I2507,I482258,I482383,);
not I_28226 (I482391,I482383);
DFFARX1 I_28227 (I301318,I2507,I482258,I482417,);
and I_28228 (I482425,I482417,I301324);
nand I_28229 (I482442,I482417,I301324);
nand I_28230 (I482229,I482391,I482442);
DFFARX1 I_28231 (I301312,I2507,I482258,I482482,);
nor I_28232 (I482490,I482482,I482425);
DFFARX1 I_28233 (I482490,I2507,I482258,I482223,);
nor I_28234 (I482238,I482482,I482383);
nand I_28235 (I482535,I301321,I301309);
and I_28236 (I482552,I482535,I301315);
DFFARX1 I_28237 (I482552,I2507,I482258,I482578,);
nor I_28238 (I482226,I482578,I482482);
not I_28239 (I482600,I482578);
nor I_28240 (I482617,I482600,I482391);
nor I_28241 (I482634,I482323,I482617);
DFFARX1 I_28242 (I482634,I2507,I482258,I482241,);
nor I_28243 (I482665,I482600,I482482);
nor I_28244 (I482682,I301327,I301309);
nor I_28245 (I482232,I482682,I482665);
not I_28246 (I482713,I482682);
nand I_28247 (I482235,I482442,I482713);
DFFARX1 I_28248 (I482682,I2507,I482258,I482247,);
DFFARX1 I_28249 (I482682,I2507,I482258,I482244,);
not I_28250 (I482802,I2514);
DFFARX1 I_28251 (I945717,I2507,I482802,I482828,);
DFFARX1 I_28252 (I482828,I2507,I482802,I482845,);
not I_28253 (I482794,I482845);
not I_28254 (I482867,I482828);
nand I_28255 (I482884,I945732,I945720);
and I_28256 (I482901,I482884,I945711);
DFFARX1 I_28257 (I482901,I2507,I482802,I482927,);
not I_28258 (I482935,I482927);
DFFARX1 I_28259 (I945723,I2507,I482802,I482961,);
and I_28260 (I482969,I482961,I945714);
nand I_28261 (I482986,I482961,I945714);
nand I_28262 (I482773,I482935,I482986);
DFFARX1 I_28263 (I945729,I2507,I482802,I483026,);
nor I_28264 (I483034,I483026,I482969);
DFFARX1 I_28265 (I483034,I2507,I482802,I482767,);
nor I_28266 (I482782,I483026,I482927);
nand I_28267 (I483079,I945738,I945726);
and I_28268 (I483096,I483079,I945735);
DFFARX1 I_28269 (I483096,I2507,I482802,I483122,);
nor I_28270 (I482770,I483122,I483026);
not I_28271 (I483144,I483122);
nor I_28272 (I483161,I483144,I482935);
nor I_28273 (I483178,I482867,I483161);
DFFARX1 I_28274 (I483178,I2507,I482802,I482785,);
nor I_28275 (I483209,I483144,I483026);
nor I_28276 (I483226,I945711,I945726);
nor I_28277 (I482776,I483226,I483209);
not I_28278 (I483257,I483226);
nand I_28279 (I482779,I482986,I483257);
DFFARX1 I_28280 (I483226,I2507,I482802,I482791,);
DFFARX1 I_28281 (I483226,I2507,I482802,I482788,);
not I_28282 (I483346,I2514);
DFFARX1 I_28283 (I1005795,I2507,I483346,I483372,);
DFFARX1 I_28284 (I483372,I2507,I483346,I483389,);
not I_28285 (I483338,I483389);
not I_28286 (I483411,I483372);
nand I_28287 (I483428,I1005810,I1005798);
and I_28288 (I483445,I483428,I1005789);
DFFARX1 I_28289 (I483445,I2507,I483346,I483471,);
not I_28290 (I483479,I483471);
DFFARX1 I_28291 (I1005801,I2507,I483346,I483505,);
and I_28292 (I483513,I483505,I1005792);
nand I_28293 (I483530,I483505,I1005792);
nand I_28294 (I483317,I483479,I483530);
DFFARX1 I_28295 (I1005807,I2507,I483346,I483570,);
nor I_28296 (I483578,I483570,I483513);
DFFARX1 I_28297 (I483578,I2507,I483346,I483311,);
nor I_28298 (I483326,I483570,I483471);
nand I_28299 (I483623,I1005816,I1005804);
and I_28300 (I483640,I483623,I1005813);
DFFARX1 I_28301 (I483640,I2507,I483346,I483666,);
nor I_28302 (I483314,I483666,I483570);
not I_28303 (I483688,I483666);
nor I_28304 (I483705,I483688,I483479);
nor I_28305 (I483722,I483411,I483705);
DFFARX1 I_28306 (I483722,I2507,I483346,I483329,);
nor I_28307 (I483753,I483688,I483570);
nor I_28308 (I483770,I1005789,I1005804);
nor I_28309 (I483320,I483770,I483753);
not I_28310 (I483801,I483770);
nand I_28311 (I483323,I483530,I483801);
DFFARX1 I_28312 (I483770,I2507,I483346,I483335,);
DFFARX1 I_28313 (I483770,I2507,I483346,I483332,);
not I_28314 (I483890,I2514);
DFFARX1 I_28315 (I1343419,I2507,I483890,I483916,);
DFFARX1 I_28316 (I483916,I2507,I483890,I483933,);
not I_28317 (I483882,I483933);
not I_28318 (I483955,I483916);
nand I_28319 (I483972,I1343395,I1343416);
and I_28320 (I483989,I483972,I1343413);
DFFARX1 I_28321 (I483989,I2507,I483890,I484015,);
not I_28322 (I484023,I484015);
DFFARX1 I_28323 (I1343392,I2507,I483890,I484049,);
and I_28324 (I484057,I484049,I1343404);
nand I_28325 (I484074,I484049,I1343404);
nand I_28326 (I483861,I484023,I484074);
DFFARX1 I_28327 (I1343407,I2507,I483890,I484114,);
nor I_28328 (I484122,I484114,I484057);
DFFARX1 I_28329 (I484122,I2507,I483890,I483855,);
nor I_28330 (I483870,I484114,I484015);
nand I_28331 (I484167,I1343410,I1343398);
and I_28332 (I484184,I484167,I1343401);
DFFARX1 I_28333 (I484184,I2507,I483890,I484210,);
nor I_28334 (I483858,I484210,I484114);
not I_28335 (I484232,I484210);
nor I_28336 (I484249,I484232,I484023);
nor I_28337 (I484266,I483955,I484249);
DFFARX1 I_28338 (I484266,I2507,I483890,I483873,);
nor I_28339 (I484297,I484232,I484114);
nor I_28340 (I484314,I1343392,I1343398);
nor I_28341 (I483864,I484314,I484297);
not I_28342 (I484345,I484314);
nand I_28343 (I483867,I484074,I484345);
DFFARX1 I_28344 (I484314,I2507,I483890,I483879,);
DFFARX1 I_28345 (I484314,I2507,I483890,I483876,);
not I_28346 (I484434,I2514);
DFFARX1 I_28347 (I1083227,I2507,I484434,I484460,);
DFFARX1 I_28348 (I484460,I2507,I484434,I484477,);
not I_28349 (I484426,I484477);
not I_28350 (I484499,I484460);
nand I_28351 (I484516,I1083239,I1083227);
and I_28352 (I484533,I484516,I1083230);
DFFARX1 I_28353 (I484533,I2507,I484434,I484559,);
not I_28354 (I484567,I484559);
DFFARX1 I_28355 (I1083248,I2507,I484434,I484593,);
and I_28356 (I484601,I484593,I1083224);
nand I_28357 (I484618,I484593,I1083224);
nand I_28358 (I484405,I484567,I484618);
DFFARX1 I_28359 (I1083242,I2507,I484434,I484658,);
nor I_28360 (I484666,I484658,I484601);
DFFARX1 I_28361 (I484666,I2507,I484434,I484399,);
nor I_28362 (I484414,I484658,I484559);
nand I_28363 (I484711,I1083236,I1083233);
and I_28364 (I484728,I484711,I1083245);
DFFARX1 I_28365 (I484728,I2507,I484434,I484754,);
nor I_28366 (I484402,I484754,I484658);
not I_28367 (I484776,I484754);
nor I_28368 (I484793,I484776,I484567);
nor I_28369 (I484810,I484499,I484793);
DFFARX1 I_28370 (I484810,I2507,I484434,I484417,);
nor I_28371 (I484841,I484776,I484658);
nor I_28372 (I484858,I1083224,I1083233);
nor I_28373 (I484408,I484858,I484841);
not I_28374 (I484889,I484858);
nand I_28375 (I484411,I484618,I484889);
DFFARX1 I_28376 (I484858,I2507,I484434,I484423,);
DFFARX1 I_28377 (I484858,I2507,I484434,I484420,);
not I_28378 (I484978,I2514);
DFFARX1 I_28379 (I870770,I2507,I484978,I485004,);
DFFARX1 I_28380 (I485004,I2507,I484978,I485021,);
not I_28381 (I484970,I485021);
not I_28382 (I485043,I485004);
nand I_28383 (I485060,I870764,I870761);
and I_28384 (I485077,I485060,I870776);
DFFARX1 I_28385 (I485077,I2507,I484978,I485103,);
not I_28386 (I485111,I485103);
DFFARX1 I_28387 (I870764,I2507,I484978,I485137,);
and I_28388 (I485145,I485137,I870758);
nand I_28389 (I485162,I485137,I870758);
nand I_28390 (I484949,I485111,I485162);
DFFARX1 I_28391 (I870758,I2507,I484978,I485202,);
nor I_28392 (I485210,I485202,I485145);
DFFARX1 I_28393 (I485210,I2507,I484978,I484943,);
nor I_28394 (I484958,I485202,I485103);
nand I_28395 (I485255,I870773,I870767);
and I_28396 (I485272,I485255,I870761);
DFFARX1 I_28397 (I485272,I2507,I484978,I485298,);
nor I_28398 (I484946,I485298,I485202);
not I_28399 (I485320,I485298);
nor I_28400 (I485337,I485320,I485111);
nor I_28401 (I485354,I485043,I485337);
DFFARX1 I_28402 (I485354,I2507,I484978,I484961,);
nor I_28403 (I485385,I485320,I485202);
nor I_28404 (I485402,I870779,I870767);
nor I_28405 (I484952,I485402,I485385);
not I_28406 (I485433,I485402);
nand I_28407 (I484955,I485162,I485433);
DFFARX1 I_28408 (I485402,I2507,I484978,I484967,);
DFFARX1 I_28409 (I485402,I2507,I484978,I484964,);
not I_28410 (I485522,I2514);
DFFARX1 I_28411 (I1021922,I2507,I485522,I485548,);
DFFARX1 I_28412 (I485548,I2507,I485522,I485565,);
not I_28413 (I485514,I485565);
not I_28414 (I485587,I485548);
nand I_28415 (I485604,I1021922,I1021940);
and I_28416 (I485621,I485604,I1021934);
DFFARX1 I_28417 (I485621,I2507,I485522,I485647,);
not I_28418 (I485655,I485647);
DFFARX1 I_28419 (I1021928,I2507,I485522,I485681,);
and I_28420 (I485689,I485681,I1021937);
nand I_28421 (I485706,I485681,I1021937);
nand I_28422 (I485493,I485655,I485706);
DFFARX1 I_28423 (I1021925,I2507,I485522,I485746,);
nor I_28424 (I485754,I485746,I485689);
DFFARX1 I_28425 (I485754,I2507,I485522,I485487,);
nor I_28426 (I485502,I485746,I485647);
nand I_28427 (I485799,I1021925,I1021943);
and I_28428 (I485816,I485799,I1021928);
DFFARX1 I_28429 (I485816,I2507,I485522,I485842,);
nor I_28430 (I485490,I485842,I485746);
not I_28431 (I485864,I485842);
nor I_28432 (I485881,I485864,I485655);
nor I_28433 (I485898,I485587,I485881);
DFFARX1 I_28434 (I485898,I2507,I485522,I485505,);
nor I_28435 (I485929,I485864,I485746);
nor I_28436 (I485946,I1021931,I1021943);
nor I_28437 (I485496,I485946,I485929);
not I_28438 (I485977,I485946);
nand I_28439 (I485499,I485706,I485977);
DFFARX1 I_28440 (I485946,I2507,I485522,I485511,);
DFFARX1 I_28441 (I485946,I2507,I485522,I485508,);
not I_28442 (I486066,I2514);
DFFARX1 I_28443 (I676961,I2507,I486066,I486092,);
DFFARX1 I_28444 (I486092,I2507,I486066,I486109,);
not I_28445 (I486058,I486109);
not I_28446 (I486131,I486092);
nand I_28447 (I486148,I676982,I676973);
and I_28448 (I486165,I486148,I676961);
DFFARX1 I_28449 (I486165,I2507,I486066,I486191,);
not I_28450 (I486199,I486191);
DFFARX1 I_28451 (I676967,I2507,I486066,I486225,);
and I_28452 (I486233,I486225,I676964);
nand I_28453 (I486250,I486225,I676964);
nand I_28454 (I486037,I486199,I486250);
DFFARX1 I_28455 (I676958,I2507,I486066,I486290,);
nor I_28456 (I486298,I486290,I486233);
DFFARX1 I_28457 (I486298,I2507,I486066,I486031,);
nor I_28458 (I486046,I486290,I486191);
nand I_28459 (I486343,I676958,I676970);
and I_28460 (I486360,I486343,I676979);
DFFARX1 I_28461 (I486360,I2507,I486066,I486386,);
nor I_28462 (I486034,I486386,I486290);
not I_28463 (I486408,I486386);
nor I_28464 (I486425,I486408,I486199);
nor I_28465 (I486442,I486131,I486425);
DFFARX1 I_28466 (I486442,I2507,I486066,I486049,);
nor I_28467 (I486473,I486408,I486290);
nor I_28468 (I486490,I676976,I676970);
nor I_28469 (I486040,I486490,I486473);
not I_28470 (I486521,I486490);
nand I_28471 (I486043,I486250,I486521);
DFFARX1 I_28472 (I486490,I2507,I486066,I486055,);
DFFARX1 I_28473 (I486490,I2507,I486066,I486052,);
not I_28474 (I486610,I2514);
DFFARX1 I_28475 (I943779,I2507,I486610,I486636,);
DFFARX1 I_28476 (I486636,I2507,I486610,I486653,);
not I_28477 (I486602,I486653);
not I_28478 (I486675,I486636);
nand I_28479 (I486692,I943794,I943782);
and I_28480 (I486709,I486692,I943773);
DFFARX1 I_28481 (I486709,I2507,I486610,I486735,);
not I_28482 (I486743,I486735);
DFFARX1 I_28483 (I943785,I2507,I486610,I486769,);
and I_28484 (I486777,I486769,I943776);
nand I_28485 (I486794,I486769,I943776);
nand I_28486 (I486581,I486743,I486794);
DFFARX1 I_28487 (I943791,I2507,I486610,I486834,);
nor I_28488 (I486842,I486834,I486777);
DFFARX1 I_28489 (I486842,I2507,I486610,I486575,);
nor I_28490 (I486590,I486834,I486735);
nand I_28491 (I486887,I943800,I943788);
and I_28492 (I486904,I486887,I943797);
DFFARX1 I_28493 (I486904,I2507,I486610,I486930,);
nor I_28494 (I486578,I486930,I486834);
not I_28495 (I486952,I486930);
nor I_28496 (I486969,I486952,I486743);
nor I_28497 (I486986,I486675,I486969);
DFFARX1 I_28498 (I486986,I2507,I486610,I486593,);
nor I_28499 (I487017,I486952,I486834);
nor I_28500 (I487034,I943773,I943788);
nor I_28501 (I486584,I487034,I487017);
not I_28502 (I487065,I487034);
nand I_28503 (I486587,I486794,I487065);
DFFARX1 I_28504 (I487034,I2507,I486610,I486599,);
DFFARX1 I_28505 (I487034,I2507,I486610,I486596,);
not I_28506 (I487154,I2514);
DFFARX1 I_28507 (I17455,I2507,I487154,I487180,);
DFFARX1 I_28508 (I487180,I2507,I487154,I487197,);
not I_28509 (I487146,I487197);
not I_28510 (I487219,I487180);
nand I_28511 (I487236,I17443,I17458);
and I_28512 (I487253,I487236,I17446);
DFFARX1 I_28513 (I487253,I2507,I487154,I487279,);
not I_28514 (I487287,I487279);
DFFARX1 I_28515 (I17467,I2507,I487154,I487313,);
and I_28516 (I487321,I487313,I17461);
nand I_28517 (I487338,I487313,I17461);
nand I_28518 (I487125,I487287,I487338);
DFFARX1 I_28519 (I17464,I2507,I487154,I487378,);
nor I_28520 (I487386,I487378,I487321);
DFFARX1 I_28521 (I487386,I2507,I487154,I487119,);
nor I_28522 (I487134,I487378,I487279);
nand I_28523 (I487431,I17443,I17446);
and I_28524 (I487448,I487431,I17449);
DFFARX1 I_28525 (I487448,I2507,I487154,I487474,);
nor I_28526 (I487122,I487474,I487378);
not I_28527 (I487496,I487474);
nor I_28528 (I487513,I487496,I487287);
nor I_28529 (I487530,I487219,I487513);
DFFARX1 I_28530 (I487530,I2507,I487154,I487137,);
nor I_28531 (I487561,I487496,I487378);
nor I_28532 (I487578,I17452,I17446);
nor I_28533 (I487128,I487578,I487561);
not I_28534 (I487609,I487578);
nand I_28535 (I487131,I487338,I487609);
DFFARX1 I_28536 (I487578,I2507,I487154,I487143,);
DFFARX1 I_28537 (I487578,I2507,I487154,I487140,);
not I_28538 (I487698,I2514);
DFFARX1 I_28539 (I965097,I2507,I487698,I487724,);
DFFARX1 I_28540 (I487724,I2507,I487698,I487741,);
not I_28541 (I487690,I487741);
not I_28542 (I487763,I487724);
nand I_28543 (I487780,I965112,I965100);
and I_28544 (I487797,I487780,I965091);
DFFARX1 I_28545 (I487797,I2507,I487698,I487823,);
not I_28546 (I487831,I487823);
DFFARX1 I_28547 (I965103,I2507,I487698,I487857,);
and I_28548 (I487865,I487857,I965094);
nand I_28549 (I487882,I487857,I965094);
nand I_28550 (I487669,I487831,I487882);
DFFARX1 I_28551 (I965109,I2507,I487698,I487922,);
nor I_28552 (I487930,I487922,I487865);
DFFARX1 I_28553 (I487930,I2507,I487698,I487663,);
nor I_28554 (I487678,I487922,I487823);
nand I_28555 (I487975,I965118,I965106);
and I_28556 (I487992,I487975,I965115);
DFFARX1 I_28557 (I487992,I2507,I487698,I488018,);
nor I_28558 (I487666,I488018,I487922);
not I_28559 (I488040,I488018);
nor I_28560 (I488057,I488040,I487831);
nor I_28561 (I488074,I487763,I488057);
DFFARX1 I_28562 (I488074,I2507,I487698,I487681,);
nor I_28563 (I488105,I488040,I487922);
nor I_28564 (I488122,I965091,I965106);
nor I_28565 (I487672,I488122,I488105);
not I_28566 (I488153,I488122);
nand I_28567 (I487675,I487882,I488153);
DFFARX1 I_28568 (I488122,I2507,I487698,I487687,);
DFFARX1 I_28569 (I488122,I2507,I487698,I487684,);
not I_28570 (I488242,I2514);
DFFARX1 I_28571 (I1001919,I2507,I488242,I488268,);
DFFARX1 I_28572 (I488268,I2507,I488242,I488285,);
not I_28573 (I488234,I488285);
not I_28574 (I488307,I488268);
nand I_28575 (I488324,I1001934,I1001922);
and I_28576 (I488341,I488324,I1001913);
DFFARX1 I_28577 (I488341,I2507,I488242,I488367,);
not I_28578 (I488375,I488367);
DFFARX1 I_28579 (I1001925,I2507,I488242,I488401,);
and I_28580 (I488409,I488401,I1001916);
nand I_28581 (I488426,I488401,I1001916);
nand I_28582 (I488213,I488375,I488426);
DFFARX1 I_28583 (I1001931,I2507,I488242,I488466,);
nor I_28584 (I488474,I488466,I488409);
DFFARX1 I_28585 (I488474,I2507,I488242,I488207,);
nor I_28586 (I488222,I488466,I488367);
nand I_28587 (I488519,I1001940,I1001928);
and I_28588 (I488536,I488519,I1001937);
DFFARX1 I_28589 (I488536,I2507,I488242,I488562,);
nor I_28590 (I488210,I488562,I488466);
not I_28591 (I488584,I488562);
nor I_28592 (I488601,I488584,I488375);
nor I_28593 (I488618,I488307,I488601);
DFFARX1 I_28594 (I488618,I2507,I488242,I488225,);
nor I_28595 (I488649,I488584,I488466);
nor I_28596 (I488666,I1001913,I1001928);
nor I_28597 (I488216,I488666,I488649);
not I_28598 (I488697,I488666);
nand I_28599 (I488219,I488426,I488697);
DFFARX1 I_28600 (I488666,I2507,I488242,I488231,);
DFFARX1 I_28601 (I488666,I2507,I488242,I488228,);
not I_28602 (I488786,I2514);
DFFARX1 I_28603 (I536932,I2507,I488786,I488812,);
DFFARX1 I_28604 (I488812,I2507,I488786,I488829,);
not I_28605 (I488778,I488829);
not I_28606 (I488851,I488812);
nand I_28607 (I488868,I536935,I536953);
and I_28608 (I488885,I488868,I536941);
DFFARX1 I_28609 (I488885,I2507,I488786,I488911,);
not I_28610 (I488919,I488911);
DFFARX1 I_28611 (I536932,I2507,I488786,I488945,);
and I_28612 (I488953,I488945,I536950);
nand I_28613 (I488970,I488945,I536950);
nand I_28614 (I488757,I488919,I488970);
DFFARX1 I_28615 (I536944,I2507,I488786,I489010,);
nor I_28616 (I489018,I489010,I488953);
DFFARX1 I_28617 (I489018,I2507,I488786,I488751,);
nor I_28618 (I488766,I489010,I488911);
nand I_28619 (I489063,I536947,I536929);
and I_28620 (I489080,I489063,I536938);
DFFARX1 I_28621 (I489080,I2507,I488786,I489106,);
nor I_28622 (I488754,I489106,I489010);
not I_28623 (I489128,I489106);
nor I_28624 (I489145,I489128,I488919);
nor I_28625 (I489162,I488851,I489145);
DFFARX1 I_28626 (I489162,I2507,I488786,I488769,);
nor I_28627 (I489193,I489128,I489010);
nor I_28628 (I489210,I536929,I536929);
nor I_28629 (I488760,I489210,I489193);
not I_28630 (I489241,I489210);
nand I_28631 (I488763,I488970,I489241);
DFFARX1 I_28632 (I489210,I2507,I488786,I488775,);
DFFARX1 I_28633 (I489210,I2507,I488786,I488772,);
not I_28634 (I489330,I2514);
DFFARX1 I_28635 (I652685,I2507,I489330,I489356,);
DFFARX1 I_28636 (I489356,I2507,I489330,I489373,);
not I_28637 (I489322,I489373);
not I_28638 (I489395,I489356);
nand I_28639 (I489412,I652706,I652697);
and I_28640 (I489429,I489412,I652685);
DFFARX1 I_28641 (I489429,I2507,I489330,I489455,);
not I_28642 (I489463,I489455);
DFFARX1 I_28643 (I652691,I2507,I489330,I489489,);
and I_28644 (I489497,I489489,I652688);
nand I_28645 (I489514,I489489,I652688);
nand I_28646 (I489301,I489463,I489514);
DFFARX1 I_28647 (I652682,I2507,I489330,I489554,);
nor I_28648 (I489562,I489554,I489497);
DFFARX1 I_28649 (I489562,I2507,I489330,I489295,);
nor I_28650 (I489310,I489554,I489455);
nand I_28651 (I489607,I652682,I652694);
and I_28652 (I489624,I489607,I652703);
DFFARX1 I_28653 (I489624,I2507,I489330,I489650,);
nor I_28654 (I489298,I489650,I489554);
not I_28655 (I489672,I489650);
nor I_28656 (I489689,I489672,I489463);
nor I_28657 (I489706,I489395,I489689);
DFFARX1 I_28658 (I489706,I2507,I489330,I489313,);
nor I_28659 (I489737,I489672,I489554);
nor I_28660 (I489754,I652700,I652694);
nor I_28661 (I489304,I489754,I489737);
not I_28662 (I489785,I489754);
nand I_28663 (I489307,I489514,I489785);
DFFARX1 I_28664 (I489754,I2507,I489330,I489319,);
DFFARX1 I_28665 (I489754,I2507,I489330,I489316,);
not I_28666 (I489874,I2514);
DFFARX1 I_28667 (I20090,I2507,I489874,I489900,);
DFFARX1 I_28668 (I489900,I2507,I489874,I489917,);
not I_28669 (I489866,I489917);
not I_28670 (I489939,I489900);
nand I_28671 (I489956,I20078,I20093);
and I_28672 (I489973,I489956,I20081);
DFFARX1 I_28673 (I489973,I2507,I489874,I489999,);
not I_28674 (I490007,I489999);
DFFARX1 I_28675 (I20102,I2507,I489874,I490033,);
and I_28676 (I490041,I490033,I20096);
nand I_28677 (I490058,I490033,I20096);
nand I_28678 (I489845,I490007,I490058);
DFFARX1 I_28679 (I20099,I2507,I489874,I490098,);
nor I_28680 (I490106,I490098,I490041);
DFFARX1 I_28681 (I490106,I2507,I489874,I489839,);
nor I_28682 (I489854,I490098,I489999);
nand I_28683 (I490151,I20078,I20081);
and I_28684 (I490168,I490151,I20084);
DFFARX1 I_28685 (I490168,I2507,I489874,I490194,);
nor I_28686 (I489842,I490194,I490098);
not I_28687 (I490216,I490194);
nor I_28688 (I490233,I490216,I490007);
nor I_28689 (I490250,I489939,I490233);
DFFARX1 I_28690 (I490250,I2507,I489874,I489857,);
nor I_28691 (I490281,I490216,I490098);
nor I_28692 (I490298,I20087,I20081);
nor I_28693 (I489848,I490298,I490281);
not I_28694 (I490329,I490298);
nand I_28695 (I489851,I490058,I490329);
DFFARX1 I_28696 (I490298,I2507,I489874,I489863,);
DFFARX1 I_28697 (I490298,I2507,I489874,I489860,);
not I_28698 (I490418,I2514);
DFFARX1 I_28699 (I213309,I2507,I490418,I490444,);
DFFARX1 I_28700 (I490444,I2507,I490418,I490461,);
not I_28701 (I490410,I490461);
not I_28702 (I490483,I490444);
nand I_28703 (I490500,I213321,I213300);
and I_28704 (I490517,I490500,I213303);
DFFARX1 I_28705 (I490517,I2507,I490418,I490543,);
not I_28706 (I490551,I490543);
DFFARX1 I_28707 (I213312,I2507,I490418,I490577,);
and I_28708 (I490585,I490577,I213324);
nand I_28709 (I490602,I490577,I213324);
nand I_28710 (I490389,I490551,I490602);
DFFARX1 I_28711 (I213318,I2507,I490418,I490642,);
nor I_28712 (I490650,I490642,I490585);
DFFARX1 I_28713 (I490650,I2507,I490418,I490383,);
nor I_28714 (I490398,I490642,I490543);
nand I_28715 (I490695,I213306,I213303);
and I_28716 (I490712,I490695,I213315);
DFFARX1 I_28717 (I490712,I2507,I490418,I490738,);
nor I_28718 (I490386,I490738,I490642);
not I_28719 (I490760,I490738);
nor I_28720 (I490777,I490760,I490551);
nor I_28721 (I490794,I490483,I490777);
DFFARX1 I_28722 (I490794,I2507,I490418,I490401,);
nor I_28723 (I490825,I490760,I490642);
nor I_28724 (I490842,I213300,I213303);
nor I_28725 (I490392,I490842,I490825);
not I_28726 (I490873,I490842);
nand I_28727 (I490395,I490602,I490873);
DFFARX1 I_28728 (I490842,I2507,I490418,I490407,);
DFFARX1 I_28729 (I490842,I2507,I490418,I490404,);
not I_28730 (I490962,I2514);
DFFARX1 I_28731 (I1138137,I2507,I490962,I490988,);
DFFARX1 I_28732 (I490988,I2507,I490962,I491005,);
not I_28733 (I490954,I491005);
not I_28734 (I491027,I490988);
nand I_28735 (I491044,I1138149,I1138137);
and I_28736 (I491061,I491044,I1138140);
DFFARX1 I_28737 (I491061,I2507,I490962,I491087,);
not I_28738 (I491095,I491087);
DFFARX1 I_28739 (I1138158,I2507,I490962,I491121,);
and I_28740 (I491129,I491121,I1138134);
nand I_28741 (I491146,I491121,I1138134);
nand I_28742 (I490933,I491095,I491146);
DFFARX1 I_28743 (I1138152,I2507,I490962,I491186,);
nor I_28744 (I491194,I491186,I491129);
DFFARX1 I_28745 (I491194,I2507,I490962,I490927,);
nor I_28746 (I490942,I491186,I491087);
nand I_28747 (I491239,I1138146,I1138143);
and I_28748 (I491256,I491239,I1138155);
DFFARX1 I_28749 (I491256,I2507,I490962,I491282,);
nor I_28750 (I490930,I491282,I491186);
not I_28751 (I491304,I491282);
nor I_28752 (I491321,I491304,I491095);
nor I_28753 (I491338,I491027,I491321);
DFFARX1 I_28754 (I491338,I2507,I490962,I490945,);
nor I_28755 (I491369,I491304,I491186);
nor I_28756 (I491386,I1138134,I1138143);
nor I_28757 (I490936,I491386,I491369);
not I_28758 (I491417,I491386);
nand I_28759 (I490939,I491146,I491417);
DFFARX1 I_28760 (I491386,I2507,I490962,I490951,);
DFFARX1 I_28761 (I491386,I2507,I490962,I490948,);
not I_28762 (I491506,I2514);
DFFARX1 I_28763 (I783288,I2507,I491506,I491532,);
DFFARX1 I_28764 (I491532,I2507,I491506,I491549,);
not I_28765 (I491498,I491549);
not I_28766 (I491571,I491532);
nand I_28767 (I491588,I783282,I783279);
and I_28768 (I491605,I491588,I783294);
DFFARX1 I_28769 (I491605,I2507,I491506,I491631,);
not I_28770 (I491639,I491631);
DFFARX1 I_28771 (I783282,I2507,I491506,I491665,);
and I_28772 (I491673,I491665,I783276);
nand I_28773 (I491690,I491665,I783276);
nand I_28774 (I491477,I491639,I491690);
DFFARX1 I_28775 (I783276,I2507,I491506,I491730,);
nor I_28776 (I491738,I491730,I491673);
DFFARX1 I_28777 (I491738,I2507,I491506,I491471,);
nor I_28778 (I491486,I491730,I491631);
nand I_28779 (I491783,I783291,I783285);
and I_28780 (I491800,I491783,I783279);
DFFARX1 I_28781 (I491800,I2507,I491506,I491826,);
nor I_28782 (I491474,I491826,I491730);
not I_28783 (I491848,I491826);
nor I_28784 (I491865,I491848,I491639);
nor I_28785 (I491882,I491571,I491865);
DFFARX1 I_28786 (I491882,I2507,I491506,I491489,);
nor I_28787 (I491913,I491848,I491730);
nor I_28788 (I491930,I783297,I783285);
nor I_28789 (I491480,I491930,I491913);
not I_28790 (I491961,I491930);
nand I_28791 (I491483,I491690,I491961);
DFFARX1 I_28792 (I491930,I2507,I491506,I491495,);
DFFARX1 I_28793 (I491930,I2507,I491506,I491492,);
not I_28794 (I492050,I2514);
DFFARX1 I_28795 (I648061,I2507,I492050,I492076,);
DFFARX1 I_28796 (I492076,I2507,I492050,I492093,);
not I_28797 (I492042,I492093);
not I_28798 (I492115,I492076);
nand I_28799 (I492132,I648082,I648073);
and I_28800 (I492149,I492132,I648061);
DFFARX1 I_28801 (I492149,I2507,I492050,I492175,);
not I_28802 (I492183,I492175);
DFFARX1 I_28803 (I648067,I2507,I492050,I492209,);
and I_28804 (I492217,I492209,I648064);
nand I_28805 (I492234,I492209,I648064);
nand I_28806 (I492021,I492183,I492234);
DFFARX1 I_28807 (I648058,I2507,I492050,I492274,);
nor I_28808 (I492282,I492274,I492217);
DFFARX1 I_28809 (I492282,I2507,I492050,I492015,);
nor I_28810 (I492030,I492274,I492175);
nand I_28811 (I492327,I648058,I648070);
and I_28812 (I492344,I492327,I648079);
DFFARX1 I_28813 (I492344,I2507,I492050,I492370,);
nor I_28814 (I492018,I492370,I492274);
not I_28815 (I492392,I492370);
nor I_28816 (I492409,I492392,I492183);
nor I_28817 (I492426,I492115,I492409);
DFFARX1 I_28818 (I492426,I2507,I492050,I492033,);
nor I_28819 (I492457,I492392,I492274);
nor I_28820 (I492474,I648076,I648070);
nor I_28821 (I492024,I492474,I492457);
not I_28822 (I492505,I492474);
nand I_28823 (I492027,I492234,I492505);
DFFARX1 I_28824 (I492474,I2507,I492050,I492039,);
DFFARX1 I_28825 (I492474,I2507,I492050,I492036,);
not I_28826 (I492594,I2514);
DFFARX1 I_28827 (I1348179,I2507,I492594,I492620,);
DFFARX1 I_28828 (I492620,I2507,I492594,I492637,);
not I_28829 (I492586,I492637);
not I_28830 (I492659,I492620);
nand I_28831 (I492676,I1348155,I1348176);
and I_28832 (I492693,I492676,I1348173);
DFFARX1 I_28833 (I492693,I2507,I492594,I492719,);
not I_28834 (I492727,I492719);
DFFARX1 I_28835 (I1348152,I2507,I492594,I492753,);
and I_28836 (I492761,I492753,I1348164);
nand I_28837 (I492778,I492753,I1348164);
nand I_28838 (I492565,I492727,I492778);
DFFARX1 I_28839 (I1348167,I2507,I492594,I492818,);
nor I_28840 (I492826,I492818,I492761);
DFFARX1 I_28841 (I492826,I2507,I492594,I492559,);
nor I_28842 (I492574,I492818,I492719);
nand I_28843 (I492871,I1348170,I1348158);
and I_28844 (I492888,I492871,I1348161);
DFFARX1 I_28845 (I492888,I2507,I492594,I492914,);
nor I_28846 (I492562,I492914,I492818);
not I_28847 (I492936,I492914);
nor I_28848 (I492953,I492936,I492727);
nor I_28849 (I492970,I492659,I492953);
DFFARX1 I_28850 (I492970,I2507,I492594,I492577,);
nor I_28851 (I493001,I492936,I492818);
nor I_28852 (I493018,I1348152,I1348158);
nor I_28853 (I492568,I493018,I493001);
not I_28854 (I493049,I493018);
nand I_28855 (I492571,I492778,I493049);
DFFARX1 I_28856 (I493018,I2507,I492594,I492583,);
DFFARX1 I_28857 (I493018,I2507,I492594,I492580,);
not I_28858 (I493138,I2514);
DFFARX1 I_28859 (I1229733,I2507,I493138,I493164,);
DFFARX1 I_28860 (I493164,I2507,I493138,I493181,);
not I_28861 (I493130,I493181);
not I_28862 (I493203,I493164);
nand I_28863 (I493220,I1229745,I1229748);
and I_28864 (I493237,I493220,I1229751);
DFFARX1 I_28865 (I493237,I2507,I493138,I493263,);
not I_28866 (I493271,I493263);
DFFARX1 I_28867 (I1229736,I2507,I493138,I493297,);
and I_28868 (I493305,I493297,I1229742);
nand I_28869 (I493322,I493297,I1229742);
nand I_28870 (I493109,I493271,I493322);
DFFARX1 I_28871 (I1229730,I2507,I493138,I493362,);
nor I_28872 (I493370,I493362,I493305);
DFFARX1 I_28873 (I493370,I2507,I493138,I493103,);
nor I_28874 (I493118,I493362,I493263);
nand I_28875 (I493415,I1229733,I1229754);
and I_28876 (I493432,I493415,I1229739);
DFFARX1 I_28877 (I493432,I2507,I493138,I493458,);
nor I_28878 (I493106,I493458,I493362);
not I_28879 (I493480,I493458);
nor I_28880 (I493497,I493480,I493271);
nor I_28881 (I493514,I493203,I493497);
DFFARX1 I_28882 (I493514,I2507,I493138,I493121,);
nor I_28883 (I493545,I493480,I493362);
nor I_28884 (I493562,I1229730,I1229754);
nor I_28885 (I493112,I493562,I493545);
not I_28886 (I493593,I493562);
nand I_28887 (I493115,I493322,I493593);
DFFARX1 I_28888 (I493562,I2507,I493138,I493127,);
DFFARX1 I_28889 (I493562,I2507,I493138,I493124,);
not I_28890 (I493682,I2514);
DFFARX1 I_28891 (I1373169,I2507,I493682,I493708,);
DFFARX1 I_28892 (I493708,I2507,I493682,I493725,);
not I_28893 (I493674,I493725);
not I_28894 (I493747,I493708);
nand I_28895 (I493764,I1373145,I1373166);
and I_28896 (I493781,I493764,I1373163);
DFFARX1 I_28897 (I493781,I2507,I493682,I493807,);
not I_28898 (I493815,I493807);
DFFARX1 I_28899 (I1373142,I2507,I493682,I493841,);
and I_28900 (I493849,I493841,I1373154);
nand I_28901 (I493866,I493841,I1373154);
nand I_28902 (I493653,I493815,I493866);
DFFARX1 I_28903 (I1373157,I2507,I493682,I493906,);
nor I_28904 (I493914,I493906,I493849);
DFFARX1 I_28905 (I493914,I2507,I493682,I493647,);
nor I_28906 (I493662,I493906,I493807);
nand I_28907 (I493959,I1373160,I1373148);
and I_28908 (I493976,I493959,I1373151);
DFFARX1 I_28909 (I493976,I2507,I493682,I494002,);
nor I_28910 (I493650,I494002,I493906);
not I_28911 (I494024,I494002);
nor I_28912 (I494041,I494024,I493815);
nor I_28913 (I494058,I493747,I494041);
DFFARX1 I_28914 (I494058,I2507,I493682,I493665,);
nor I_28915 (I494089,I494024,I493906);
nor I_28916 (I494106,I1373142,I1373148);
nor I_28917 (I493656,I494106,I494089);
not I_28918 (I494137,I494106);
nand I_28919 (I493659,I493866,I494137);
DFFARX1 I_28920 (I494106,I2507,I493682,I493671,);
DFFARX1 I_28921 (I494106,I2507,I493682,I493668,);
not I_28922 (I494226,I2514);
DFFARX1 I_28923 (I1344609,I2507,I494226,I494252,);
DFFARX1 I_28924 (I494252,I2507,I494226,I494269,);
not I_28925 (I494218,I494269);
not I_28926 (I494291,I494252);
nand I_28927 (I494308,I1344585,I1344606);
and I_28928 (I494325,I494308,I1344603);
DFFARX1 I_28929 (I494325,I2507,I494226,I494351,);
not I_28930 (I494359,I494351);
DFFARX1 I_28931 (I1344582,I2507,I494226,I494385,);
and I_28932 (I494393,I494385,I1344594);
nand I_28933 (I494410,I494385,I1344594);
nand I_28934 (I494197,I494359,I494410);
DFFARX1 I_28935 (I1344597,I2507,I494226,I494450,);
nor I_28936 (I494458,I494450,I494393);
DFFARX1 I_28937 (I494458,I2507,I494226,I494191,);
nor I_28938 (I494206,I494450,I494351);
nand I_28939 (I494503,I1344600,I1344588);
and I_28940 (I494520,I494503,I1344591);
DFFARX1 I_28941 (I494520,I2507,I494226,I494546,);
nor I_28942 (I494194,I494546,I494450);
not I_28943 (I494568,I494546);
nor I_28944 (I494585,I494568,I494359);
nor I_28945 (I494602,I494291,I494585);
DFFARX1 I_28946 (I494602,I2507,I494226,I494209,);
nor I_28947 (I494633,I494568,I494450);
nor I_28948 (I494650,I1344582,I1344588);
nor I_28949 (I494200,I494650,I494633);
not I_28950 (I494681,I494650);
nand I_28951 (I494203,I494410,I494681);
DFFARX1 I_28952 (I494650,I2507,I494226,I494215,);
DFFARX1 I_28953 (I494650,I2507,I494226,I494212,);
not I_28954 (I494770,I2514);
DFFARX1 I_28955 (I73311,I2507,I494770,I494796,);
DFFARX1 I_28956 (I494796,I2507,I494770,I494813,);
not I_28957 (I494762,I494813);
not I_28958 (I494835,I494796);
nand I_28959 (I494852,I73326,I73305);
and I_28960 (I494869,I494852,I73308);
DFFARX1 I_28961 (I494869,I2507,I494770,I494895,);
not I_28962 (I494903,I494895);
DFFARX1 I_28963 (I73314,I2507,I494770,I494929,);
and I_28964 (I494937,I494929,I73308);
nand I_28965 (I494954,I494929,I73308);
nand I_28966 (I494741,I494903,I494954);
DFFARX1 I_28967 (I73323,I2507,I494770,I494994,);
nor I_28968 (I495002,I494994,I494937);
DFFARX1 I_28969 (I495002,I2507,I494770,I494735,);
nor I_28970 (I494750,I494994,I494895);
nand I_28971 (I495047,I73305,I73320);
and I_28972 (I495064,I495047,I73317);
DFFARX1 I_28973 (I495064,I2507,I494770,I495090,);
nor I_28974 (I494738,I495090,I494994);
not I_28975 (I495112,I495090);
nor I_28976 (I495129,I495112,I494903);
nor I_28977 (I495146,I494835,I495129);
DFFARX1 I_28978 (I495146,I2507,I494770,I494753,);
nor I_28979 (I495177,I495112,I494994);
nor I_28980 (I495194,I73329,I73320);
nor I_28981 (I494744,I495194,I495177);
not I_28982 (I495225,I495194);
nand I_28983 (I494747,I494954,I495225);
DFFARX1 I_28984 (I495194,I2507,I494770,I494759,);
DFFARX1 I_28985 (I495194,I2507,I494770,I494756,);
not I_28986 (I495311,I2514);
DFFARX1 I_28987 (I932160,I2507,I495311,I495337,);
DFFARX1 I_28988 (I495337,I2507,I495311,I495354,);
not I_28989 (I495303,I495354);
DFFARX1 I_28990 (I932148,I2507,I495311,I495385,);
not I_28991 (I495393,I932145);
nor I_28992 (I495410,I495337,I495393);
not I_28993 (I495427,I932157);
not I_28994 (I495444,I932154);
nand I_28995 (I495461,I495444,I932157);
nor I_28996 (I495478,I495393,I495461);
nor I_28997 (I495495,I495385,I495478);
DFFARX1 I_28998 (I495444,I2507,I495311,I495300,);
nor I_28999 (I495526,I932154,I932163);
nand I_29000 (I495543,I495526,I932166);
nor I_29001 (I495560,I495543,I495427);
nand I_29002 (I495285,I495560,I932145);
DFFARX1 I_29003 (I495543,I2507,I495311,I495297,);
nand I_29004 (I495605,I495427,I932154);
nor I_29005 (I495622,I495427,I932154);
nand I_29006 (I495291,I495410,I495622);
not I_29007 (I495653,I932169);
nor I_29008 (I495670,I495653,I495605);
DFFARX1 I_29009 (I495670,I2507,I495311,I495279,);
nor I_29010 (I495701,I495653,I932172);
and I_29011 (I495718,I495701,I932151);
or I_29012 (I495735,I495718,I932145);
DFFARX1 I_29013 (I495735,I2507,I495311,I495761,);
nor I_29014 (I495769,I495761,I495385);
nor I_29015 (I495288,I495337,I495769);
not I_29016 (I495800,I495761);
nor I_29017 (I495817,I495800,I495495);
DFFARX1 I_29018 (I495817,I2507,I495311,I495294,);
nand I_29019 (I495848,I495800,I495427);
nor I_29020 (I495282,I495653,I495848);
not I_29021 (I495906,I2514);
DFFARX1 I_29022 (I1097692,I2507,I495906,I495932,);
DFFARX1 I_29023 (I495932,I2507,I495906,I495949,);
not I_29024 (I495898,I495949);
DFFARX1 I_29025 (I1097674,I2507,I495906,I495980,);
not I_29026 (I495988,I1097680);
nor I_29027 (I496005,I495932,I495988);
not I_29028 (I496022,I1097695);
not I_29029 (I496039,I1097686);
nand I_29030 (I496056,I496039,I1097695);
nor I_29031 (I496073,I495988,I496056);
nor I_29032 (I496090,I495980,I496073);
DFFARX1 I_29033 (I496039,I2507,I495906,I495895,);
nor I_29034 (I496121,I1097686,I1097698);
nand I_29035 (I496138,I496121,I1097677);
nor I_29036 (I496155,I496138,I496022);
nand I_29037 (I495880,I496155,I1097680);
DFFARX1 I_29038 (I496138,I2507,I495906,I495892,);
nand I_29039 (I496200,I496022,I1097686);
nor I_29040 (I496217,I496022,I1097686);
nand I_29041 (I495886,I496005,I496217);
not I_29042 (I496248,I1097683);
nor I_29043 (I496265,I496248,I496200);
DFFARX1 I_29044 (I496265,I2507,I495906,I495874,);
nor I_29045 (I496296,I496248,I1097689);
and I_29046 (I496313,I496296,I1097674);
or I_29047 (I496330,I496313,I1097677);
DFFARX1 I_29048 (I496330,I2507,I495906,I496356,);
nor I_29049 (I496364,I496356,I495980);
nor I_29050 (I495883,I495932,I496364);
not I_29051 (I496395,I496356);
nor I_29052 (I496412,I496395,I496090);
DFFARX1 I_29053 (I496412,I2507,I495906,I495889,);
nand I_29054 (I496443,I496395,I496022);
nor I_29055 (I495877,I496248,I496443);
not I_29056 (I496501,I2514);
DFFARX1 I_29057 (I864970,I2507,I496501,I496527,);
DFFARX1 I_29058 (I496527,I2507,I496501,I496544,);
not I_29059 (I496493,I496544);
DFFARX1 I_29060 (I864967,I2507,I496501,I496575,);
not I_29061 (I496583,I864967);
nor I_29062 (I496600,I496527,I496583);
not I_29063 (I496617,I864964);
not I_29064 (I496634,I864979);
nand I_29065 (I496651,I496634,I864964);
nor I_29066 (I496668,I496583,I496651);
nor I_29067 (I496685,I496575,I496668);
DFFARX1 I_29068 (I496634,I2507,I496501,I496490,);
nor I_29069 (I496716,I864979,I864973);
nand I_29070 (I496733,I496716,I864961);
nor I_29071 (I496750,I496733,I496617);
nand I_29072 (I496475,I496750,I864967);
DFFARX1 I_29073 (I496733,I2507,I496501,I496487,);
nand I_29074 (I496795,I496617,I864979);
nor I_29075 (I496812,I496617,I864979);
nand I_29076 (I496481,I496600,I496812);
not I_29077 (I496843,I864982);
nor I_29078 (I496860,I496843,I496795);
DFFARX1 I_29079 (I496860,I2507,I496501,I496469,);
nor I_29080 (I496891,I496843,I864961);
and I_29081 (I496908,I496891,I864976);
or I_29082 (I496925,I496908,I864964);
DFFARX1 I_29083 (I496925,I2507,I496501,I496951,);
nor I_29084 (I496959,I496951,I496575);
nor I_29085 (I496478,I496527,I496959);
not I_29086 (I496990,I496951);
nor I_29087 (I497007,I496990,I496685);
DFFARX1 I_29088 (I497007,I2507,I496501,I496484,);
nand I_29089 (I497038,I496990,I496617);
nor I_29090 (I496472,I496843,I497038);
not I_29091 (I497096,I2514);
DFFARX1 I_29092 (I1067636,I2507,I497096,I497122,);
DFFARX1 I_29093 (I497122,I2507,I497096,I497139,);
not I_29094 (I497088,I497139);
DFFARX1 I_29095 (I1067618,I2507,I497096,I497170,);
not I_29096 (I497178,I1067624);
nor I_29097 (I497195,I497122,I497178);
not I_29098 (I497212,I1067639);
not I_29099 (I497229,I1067630);
nand I_29100 (I497246,I497229,I1067639);
nor I_29101 (I497263,I497178,I497246);
nor I_29102 (I497280,I497170,I497263);
DFFARX1 I_29103 (I497229,I2507,I497096,I497085,);
nor I_29104 (I497311,I1067630,I1067642);
nand I_29105 (I497328,I497311,I1067621);
nor I_29106 (I497345,I497328,I497212);
nand I_29107 (I497070,I497345,I1067624);
DFFARX1 I_29108 (I497328,I2507,I497096,I497082,);
nand I_29109 (I497390,I497212,I1067630);
nor I_29110 (I497407,I497212,I1067630);
nand I_29111 (I497076,I497195,I497407);
not I_29112 (I497438,I1067627);
nor I_29113 (I497455,I497438,I497390);
DFFARX1 I_29114 (I497455,I2507,I497096,I497064,);
nor I_29115 (I497486,I497438,I1067633);
and I_29116 (I497503,I497486,I1067618);
or I_29117 (I497520,I497503,I1067621);
DFFARX1 I_29118 (I497520,I2507,I497096,I497546,);
nor I_29119 (I497554,I497546,I497170);
nor I_29120 (I497073,I497122,I497554);
not I_29121 (I497585,I497546);
nor I_29122 (I497602,I497585,I497280);
DFFARX1 I_29123 (I497602,I2507,I497096,I497079,);
nand I_29124 (I497633,I497585,I497212);
nor I_29125 (I497067,I497438,I497633);
not I_29126 (I497691,I2514);
DFFARX1 I_29127 (I792771,I2507,I497691,I497717,);
DFFARX1 I_29128 (I497717,I2507,I497691,I497734,);
not I_29129 (I497683,I497734);
DFFARX1 I_29130 (I792768,I2507,I497691,I497765,);
not I_29131 (I497773,I792768);
nor I_29132 (I497790,I497717,I497773);
not I_29133 (I497807,I792765);
not I_29134 (I497824,I792780);
nand I_29135 (I497841,I497824,I792765);
nor I_29136 (I497858,I497773,I497841);
nor I_29137 (I497875,I497765,I497858);
DFFARX1 I_29138 (I497824,I2507,I497691,I497680,);
nor I_29139 (I497906,I792780,I792774);
nand I_29140 (I497923,I497906,I792762);
nor I_29141 (I497940,I497923,I497807);
nand I_29142 (I497665,I497940,I792768);
DFFARX1 I_29143 (I497923,I2507,I497691,I497677,);
nand I_29144 (I497985,I497807,I792780);
nor I_29145 (I498002,I497807,I792780);
nand I_29146 (I497671,I497790,I498002);
not I_29147 (I498033,I792783);
nor I_29148 (I498050,I498033,I497985);
DFFARX1 I_29149 (I498050,I2507,I497691,I497659,);
nor I_29150 (I498081,I498033,I792762);
and I_29151 (I498098,I498081,I792777);
or I_29152 (I498115,I498098,I792765);
DFFARX1 I_29153 (I498115,I2507,I497691,I498141,);
nor I_29154 (I498149,I498141,I497765);
nor I_29155 (I497668,I497717,I498149);
not I_29156 (I498180,I498141);
nor I_29157 (I498197,I498180,I497875);
DFFARX1 I_29158 (I498197,I2507,I497691,I497674,);
nand I_29159 (I498228,I498180,I497807);
nor I_29160 (I497662,I498033,I498228);
not I_29161 (I498286,I2514);
DFFARX1 I_29162 (I956708,I2507,I498286,I498312,);
DFFARX1 I_29163 (I498312,I2507,I498286,I498329,);
not I_29164 (I498278,I498329);
DFFARX1 I_29165 (I956696,I2507,I498286,I498360,);
not I_29166 (I498368,I956693);
nor I_29167 (I498385,I498312,I498368);
not I_29168 (I498402,I956705);
not I_29169 (I498419,I956702);
nand I_29170 (I498436,I498419,I956705);
nor I_29171 (I498453,I498368,I498436);
nor I_29172 (I498470,I498360,I498453);
DFFARX1 I_29173 (I498419,I2507,I498286,I498275,);
nor I_29174 (I498501,I956702,I956711);
nand I_29175 (I498518,I498501,I956714);
nor I_29176 (I498535,I498518,I498402);
nand I_29177 (I498260,I498535,I956693);
DFFARX1 I_29178 (I498518,I2507,I498286,I498272,);
nand I_29179 (I498580,I498402,I956702);
nor I_29180 (I498597,I498402,I956702);
nand I_29181 (I498266,I498385,I498597);
not I_29182 (I498628,I956717);
nor I_29183 (I498645,I498628,I498580);
DFFARX1 I_29184 (I498645,I2507,I498286,I498254,);
nor I_29185 (I498676,I498628,I956720);
and I_29186 (I498693,I498676,I956699);
or I_29187 (I498710,I498693,I956693);
DFFARX1 I_29188 (I498710,I2507,I498286,I498736,);
nor I_29189 (I498744,I498736,I498360);
nor I_29190 (I498263,I498312,I498744);
not I_29191 (I498775,I498736);
nor I_29192 (I498792,I498775,I498470);
DFFARX1 I_29193 (I498792,I2507,I498286,I498269,);
nand I_29194 (I498823,I498775,I498402);
nor I_29195 (I498257,I498628,I498823);
not I_29196 (I498881,I2514);
DFFARX1 I_29197 (I1113298,I2507,I498881,I498907,);
DFFARX1 I_29198 (I498907,I2507,I498881,I498924,);
not I_29199 (I498873,I498924);
DFFARX1 I_29200 (I1113280,I2507,I498881,I498955,);
not I_29201 (I498963,I1113286);
nor I_29202 (I498980,I498907,I498963);
not I_29203 (I498997,I1113301);
not I_29204 (I499014,I1113292);
nand I_29205 (I499031,I499014,I1113301);
nor I_29206 (I499048,I498963,I499031);
nor I_29207 (I499065,I498955,I499048);
DFFARX1 I_29208 (I499014,I2507,I498881,I498870,);
nor I_29209 (I499096,I1113292,I1113304);
nand I_29210 (I499113,I499096,I1113283);
nor I_29211 (I499130,I499113,I498997);
nand I_29212 (I498855,I499130,I1113286);
DFFARX1 I_29213 (I499113,I2507,I498881,I498867,);
nand I_29214 (I499175,I498997,I1113292);
nor I_29215 (I499192,I498997,I1113292);
nand I_29216 (I498861,I498980,I499192);
not I_29217 (I499223,I1113289);
nor I_29218 (I499240,I499223,I499175);
DFFARX1 I_29219 (I499240,I2507,I498881,I498849,);
nor I_29220 (I499271,I499223,I1113295);
and I_29221 (I499288,I499271,I1113280);
or I_29222 (I499305,I499288,I1113283);
DFFARX1 I_29223 (I499305,I2507,I498881,I499331,);
nor I_29224 (I499339,I499331,I498955);
nor I_29225 (I498858,I498907,I499339);
not I_29226 (I499370,I499331);
nor I_29227 (I499387,I499370,I499065);
DFFARX1 I_29228 (I499387,I2507,I498881,I498864,);
nand I_29229 (I499418,I499370,I498997);
nor I_29230 (I498852,I499223,I499418);
not I_29231 (I499476,I2514);
DFFARX1 I_29232 (I998052,I2507,I499476,I499502,);
DFFARX1 I_29233 (I499502,I2507,I499476,I499519,);
not I_29234 (I499468,I499519);
DFFARX1 I_29235 (I998040,I2507,I499476,I499550,);
not I_29236 (I499558,I998037);
nor I_29237 (I499575,I499502,I499558);
not I_29238 (I499592,I998049);
not I_29239 (I499609,I998046);
nand I_29240 (I499626,I499609,I998049);
nor I_29241 (I499643,I499558,I499626);
nor I_29242 (I499660,I499550,I499643);
DFFARX1 I_29243 (I499609,I2507,I499476,I499465,);
nor I_29244 (I499691,I998046,I998055);
nand I_29245 (I499708,I499691,I998058);
nor I_29246 (I499725,I499708,I499592);
nand I_29247 (I499450,I499725,I998037);
DFFARX1 I_29248 (I499708,I2507,I499476,I499462,);
nand I_29249 (I499770,I499592,I998046);
nor I_29250 (I499787,I499592,I998046);
nand I_29251 (I499456,I499575,I499787);
not I_29252 (I499818,I998061);
nor I_29253 (I499835,I499818,I499770);
DFFARX1 I_29254 (I499835,I2507,I499476,I499444,);
nor I_29255 (I499866,I499818,I998064);
and I_29256 (I499883,I499866,I998043);
or I_29257 (I499900,I499883,I998037);
DFFARX1 I_29258 (I499900,I2507,I499476,I499926,);
nor I_29259 (I499934,I499926,I499550);
nor I_29260 (I499453,I499502,I499934);
not I_29261 (I499965,I499926);
nor I_29262 (I499982,I499965,I499660);
DFFARX1 I_29263 (I499982,I2507,I499476,I499459,);
nand I_29264 (I500013,I499965,I499592);
nor I_29265 (I499447,I499818,I500013);
not I_29266 (I500071,I2514);
DFFARX1 I_29267 (I289203,I2507,I500071,I500097,);
DFFARX1 I_29268 (I500097,I2507,I500071,I500114,);
not I_29269 (I500063,I500114);
DFFARX1 I_29270 (I289191,I2507,I500071,I500145,);
not I_29271 (I500153,I289194);
nor I_29272 (I500170,I500097,I500153);
not I_29273 (I500187,I289197);
not I_29274 (I500204,I289209);
nand I_29275 (I500221,I500204,I289197);
nor I_29276 (I500238,I500153,I500221);
nor I_29277 (I500255,I500145,I500238);
DFFARX1 I_29278 (I500204,I2507,I500071,I500060,);
nor I_29279 (I500286,I289209,I289200);
nand I_29280 (I500303,I500286,I289188);
nor I_29281 (I500320,I500303,I500187);
nand I_29282 (I500045,I500320,I289194);
DFFARX1 I_29283 (I500303,I2507,I500071,I500057,);
nand I_29284 (I500365,I500187,I289209);
nor I_29285 (I500382,I500187,I289209);
nand I_29286 (I500051,I500170,I500382);
not I_29287 (I500413,I289206);
nor I_29288 (I500430,I500413,I500365);
DFFARX1 I_29289 (I500430,I2507,I500071,I500039,);
nor I_29290 (I500461,I500413,I289212);
and I_29291 (I500478,I500461,I289215);
or I_29292 (I500495,I500478,I289188);
DFFARX1 I_29293 (I500495,I2507,I500071,I500521,);
nor I_29294 (I500529,I500521,I500145);
nor I_29295 (I500048,I500097,I500529);
not I_29296 (I500560,I500521);
nor I_29297 (I500577,I500560,I500255);
DFFARX1 I_29298 (I500577,I2507,I500071,I500054,);
nand I_29299 (I500608,I500560,I500187);
nor I_29300 (I500042,I500413,I500608);
not I_29301 (I500666,I2514);
DFFARX1 I_29302 (I489295,I2507,I500666,I500692,);
DFFARX1 I_29303 (I500692,I2507,I500666,I500709,);
not I_29304 (I500658,I500709);
DFFARX1 I_29305 (I489319,I2507,I500666,I500740,);
not I_29306 (I500748,I489298);
nor I_29307 (I500765,I500692,I500748);
not I_29308 (I500782,I489304);
not I_29309 (I500799,I489310);
nand I_29310 (I500816,I500799,I489304);
nor I_29311 (I500833,I500748,I500816);
nor I_29312 (I500850,I500740,I500833);
DFFARX1 I_29313 (I500799,I2507,I500666,I500655,);
nor I_29314 (I500881,I489310,I489322);
nand I_29315 (I500898,I500881,I489316);
nor I_29316 (I500915,I500898,I500782);
nand I_29317 (I500640,I500915,I489298);
DFFARX1 I_29318 (I500898,I2507,I500666,I500652,);
nand I_29319 (I500960,I500782,I489310);
nor I_29320 (I500977,I500782,I489310);
nand I_29321 (I500646,I500765,I500977);
not I_29322 (I501008,I489301);
nor I_29323 (I501025,I501008,I500960);
DFFARX1 I_29324 (I501025,I2507,I500666,I500634,);
nor I_29325 (I501056,I501008,I489295);
and I_29326 (I501073,I501056,I489313);
or I_29327 (I501090,I501073,I489307);
DFFARX1 I_29328 (I501090,I2507,I500666,I501116,);
nor I_29329 (I501124,I501116,I500740);
nor I_29330 (I500643,I500692,I501124);
not I_29331 (I501155,I501116);
nor I_29332 (I501172,I501155,I500850);
DFFARX1 I_29333 (I501172,I2507,I500666,I500649,);
nand I_29334 (I501203,I501155,I500782);
nor I_29335 (I500637,I501008,I501203);
not I_29336 (I501261,I2514);
DFFARX1 I_29337 (I563673,I2507,I501261,I501287,);
DFFARX1 I_29338 (I501287,I2507,I501261,I501304,);
not I_29339 (I501253,I501304);
DFFARX1 I_29340 (I563685,I2507,I501261,I501335,);
not I_29341 (I501343,I563670);
nor I_29342 (I501360,I501287,I501343);
not I_29343 (I501377,I563688);
not I_29344 (I501394,I563679);
nand I_29345 (I501411,I501394,I563688);
nor I_29346 (I501428,I501343,I501411);
nor I_29347 (I501445,I501335,I501428);
DFFARX1 I_29348 (I501394,I2507,I501261,I501250,);
nor I_29349 (I501476,I563679,I563691);
nand I_29350 (I501493,I501476,I563694);
nor I_29351 (I501510,I501493,I501377);
nand I_29352 (I501235,I501510,I563670);
DFFARX1 I_29353 (I501493,I2507,I501261,I501247,);
nand I_29354 (I501555,I501377,I563679);
nor I_29355 (I501572,I501377,I563679);
nand I_29356 (I501241,I501360,I501572);
not I_29357 (I501603,I563670);
nor I_29358 (I501620,I501603,I501555);
DFFARX1 I_29359 (I501620,I2507,I501261,I501229,);
nor I_29360 (I501651,I501603,I563682);
and I_29361 (I501668,I501651,I563676);
or I_29362 (I501685,I501668,I563673);
DFFARX1 I_29363 (I501685,I2507,I501261,I501711,);
nor I_29364 (I501719,I501711,I501335);
nor I_29365 (I501238,I501287,I501719);
not I_29366 (I501750,I501711);
nor I_29367 (I501767,I501750,I501445);
DFFARX1 I_29368 (I501767,I2507,I501261,I501244,);
nand I_29369 (I501798,I501750,I501377);
nor I_29370 (I501232,I501603,I501798);
not I_29371 (I501856,I2514);
DFFARX1 I_29372 (I1225922,I2507,I501856,I501882,);
DFFARX1 I_29373 (I501882,I2507,I501856,I501899,);
not I_29374 (I501848,I501899);
DFFARX1 I_29375 (I1225937,I2507,I501856,I501930,);
not I_29376 (I501938,I1225946);
nor I_29377 (I501955,I501882,I501938);
not I_29378 (I501972,I1225925);
not I_29379 (I501989,I1225931);
nand I_29380 (I502006,I501989,I1225925);
nor I_29381 (I502023,I501938,I502006);
nor I_29382 (I502040,I501930,I502023);
DFFARX1 I_29383 (I501989,I2507,I501856,I501845,);
nor I_29384 (I502071,I1225931,I1225943);
nand I_29385 (I502088,I502071,I1225940);
nor I_29386 (I502105,I502088,I501972);
nand I_29387 (I501830,I502105,I1225946);
DFFARX1 I_29388 (I502088,I2507,I501856,I501842,);
nand I_29389 (I502150,I501972,I1225931);
nor I_29390 (I502167,I501972,I1225931);
nand I_29391 (I501836,I501955,I502167);
not I_29392 (I502198,I1225922);
nor I_29393 (I502215,I502198,I502150);
DFFARX1 I_29394 (I502215,I2507,I501856,I501824,);
nor I_29395 (I502246,I502198,I1225934);
and I_29396 (I502263,I502246,I1225928);
or I_29397 (I502280,I502263,I1225925);
DFFARX1 I_29398 (I502280,I2507,I501856,I502306,);
nor I_29399 (I502314,I502306,I501930);
nor I_29400 (I501833,I501882,I502314);
not I_29401 (I502345,I502306);
nor I_29402 (I502362,I502345,I502040);
DFFARX1 I_29403 (I502362,I2507,I501856,I501839,);
nand I_29404 (I502393,I502345,I501972);
nor I_29405 (I501827,I502198,I502393);
not I_29406 (I502451,I2514);
DFFARX1 I_29407 (I656737,I2507,I502451,I502477,);
DFFARX1 I_29408 (I502477,I2507,I502451,I502494,);
not I_29409 (I502443,I502494);
DFFARX1 I_29410 (I656731,I2507,I502451,I502525,);
not I_29411 (I502533,I656728);
nor I_29412 (I502550,I502477,I502533);
not I_29413 (I502567,I656740);
not I_29414 (I502584,I656743);
nand I_29415 (I502601,I502584,I656740);
nor I_29416 (I502618,I502533,I502601);
nor I_29417 (I502635,I502525,I502618);
DFFARX1 I_29418 (I502584,I2507,I502451,I502440,);
nor I_29419 (I502666,I656743,I656752);
nand I_29420 (I502683,I502666,I656746);
nor I_29421 (I502700,I502683,I502567);
nand I_29422 (I502425,I502700,I656728);
DFFARX1 I_29423 (I502683,I2507,I502451,I502437,);
nand I_29424 (I502745,I502567,I656743);
nor I_29425 (I502762,I502567,I656743);
nand I_29426 (I502431,I502550,I502762);
not I_29427 (I502793,I656734);
nor I_29428 (I502810,I502793,I502745);
DFFARX1 I_29429 (I502810,I2507,I502451,I502419,);
nor I_29430 (I502841,I502793,I656749);
and I_29431 (I502858,I502841,I656728);
or I_29432 (I502875,I502858,I656731);
DFFARX1 I_29433 (I502875,I2507,I502451,I502901,);
nor I_29434 (I502909,I502901,I502525);
nor I_29435 (I502428,I502477,I502909);
not I_29436 (I502940,I502901);
nor I_29437 (I502957,I502940,I502635);
DFFARX1 I_29438 (I502957,I2507,I502451,I502434,);
nand I_29439 (I502988,I502940,I502567);
nor I_29440 (I502422,I502793,I502988);
not I_29441 (I503046,I2514);
DFFARX1 I_29442 (I393007,I2507,I503046,I503072,);
DFFARX1 I_29443 (I503072,I2507,I503046,I503089,);
not I_29444 (I503038,I503089);
DFFARX1 I_29445 (I393031,I2507,I503046,I503120,);
not I_29446 (I503128,I393010);
nor I_29447 (I503145,I503072,I503128);
not I_29448 (I503162,I393016);
not I_29449 (I503179,I393022);
nand I_29450 (I503196,I503179,I393016);
nor I_29451 (I503213,I503128,I503196);
nor I_29452 (I503230,I503120,I503213);
DFFARX1 I_29453 (I503179,I2507,I503046,I503035,);
nor I_29454 (I503261,I393022,I393034);
nand I_29455 (I503278,I503261,I393028);
nor I_29456 (I503295,I503278,I503162);
nand I_29457 (I503020,I503295,I393010);
DFFARX1 I_29458 (I503278,I2507,I503046,I503032,);
nand I_29459 (I503340,I503162,I393022);
nor I_29460 (I503357,I503162,I393022);
nand I_29461 (I503026,I503145,I503357);
not I_29462 (I503388,I393013);
nor I_29463 (I503405,I503388,I503340);
DFFARX1 I_29464 (I503405,I2507,I503046,I503014,);
nor I_29465 (I503436,I503388,I393007);
and I_29466 (I503453,I503436,I393025);
or I_29467 (I503470,I503453,I393019);
DFFARX1 I_29468 (I503470,I2507,I503046,I503496,);
nor I_29469 (I503504,I503496,I503120);
nor I_29470 (I503023,I503072,I503504);
not I_29471 (I503535,I503496);
nor I_29472 (I503552,I503535,I503230);
DFFARX1 I_29473 (I503552,I2507,I503046,I503029,);
nand I_29474 (I503583,I503535,I503162);
nor I_29475 (I503017,I503388,I503583);
not I_29476 (I503641,I2514);
DFFARX1 I_29477 (I308702,I2507,I503641,I503667,);
DFFARX1 I_29478 (I503667,I2507,I503641,I503684,);
not I_29479 (I503633,I503684);
DFFARX1 I_29480 (I308690,I2507,I503641,I503715,);
not I_29481 (I503723,I308693);
nor I_29482 (I503740,I503667,I503723);
not I_29483 (I503757,I308696);
not I_29484 (I503774,I308708);
nand I_29485 (I503791,I503774,I308696);
nor I_29486 (I503808,I503723,I503791);
nor I_29487 (I503825,I503715,I503808);
DFFARX1 I_29488 (I503774,I2507,I503641,I503630,);
nor I_29489 (I503856,I308708,I308699);
nand I_29490 (I503873,I503856,I308687);
nor I_29491 (I503890,I503873,I503757);
nand I_29492 (I503615,I503890,I308693);
DFFARX1 I_29493 (I503873,I2507,I503641,I503627,);
nand I_29494 (I503935,I503757,I308708);
nor I_29495 (I503952,I503757,I308708);
nand I_29496 (I503621,I503740,I503952);
not I_29497 (I503983,I308705);
nor I_29498 (I504000,I503983,I503935);
DFFARX1 I_29499 (I504000,I2507,I503641,I503609,);
nor I_29500 (I504031,I503983,I308711);
and I_29501 (I504048,I504031,I308714);
or I_29502 (I504065,I504048,I308687);
DFFARX1 I_29503 (I504065,I2507,I503641,I504091,);
nor I_29504 (I504099,I504091,I503715);
nor I_29505 (I503618,I503667,I504099);
not I_29506 (I504130,I504091);
nor I_29507 (I504147,I504130,I503825);
DFFARX1 I_29508 (I504147,I2507,I503641,I503624,);
nand I_29509 (I504178,I504130,I503757);
nor I_29510 (I503612,I503983,I504178);
not I_29511 (I504236,I2514);
DFFARX1 I_29512 (I820175,I2507,I504236,I504262,);
DFFARX1 I_29513 (I504262,I2507,I504236,I504279,);
not I_29514 (I504228,I504279);
DFFARX1 I_29515 (I820172,I2507,I504236,I504310,);
not I_29516 (I504318,I820172);
nor I_29517 (I504335,I504262,I504318);
not I_29518 (I504352,I820169);
not I_29519 (I504369,I820184);
nand I_29520 (I504386,I504369,I820169);
nor I_29521 (I504403,I504318,I504386);
nor I_29522 (I504420,I504310,I504403);
DFFARX1 I_29523 (I504369,I2507,I504236,I504225,);
nor I_29524 (I504451,I820184,I820178);
nand I_29525 (I504468,I504451,I820166);
nor I_29526 (I504485,I504468,I504352);
nand I_29527 (I504210,I504485,I820172);
DFFARX1 I_29528 (I504468,I2507,I504236,I504222,);
nand I_29529 (I504530,I504352,I820184);
nor I_29530 (I504547,I504352,I820184);
nand I_29531 (I504216,I504335,I504547);
not I_29532 (I504578,I820187);
nor I_29533 (I504595,I504578,I504530);
DFFARX1 I_29534 (I504595,I2507,I504236,I504204,);
nor I_29535 (I504626,I504578,I820166);
and I_29536 (I504643,I504626,I820181);
or I_29537 (I504660,I504643,I820169);
DFFARX1 I_29538 (I504660,I2507,I504236,I504686,);
nor I_29539 (I504694,I504686,I504310);
nor I_29540 (I504213,I504262,I504694);
not I_29541 (I504725,I504686);
nor I_29542 (I504742,I504725,I504420);
DFFARX1 I_29543 (I504742,I2507,I504236,I504219,);
nand I_29544 (I504773,I504725,I504352);
nor I_29545 (I504207,I504578,I504773);
not I_29546 (I504831,I2514);
DFFARX1 I_29547 (I1310072,I2507,I504831,I504857,);
DFFARX1 I_29548 (I504857,I2507,I504831,I504874,);
not I_29549 (I504823,I504874);
DFFARX1 I_29550 (I1310078,I2507,I504831,I504905,);
not I_29551 (I504913,I1310093);
nor I_29552 (I504930,I504857,I504913);
not I_29553 (I504947,I1310084);
not I_29554 (I504964,I1310081);
nand I_29555 (I504981,I504964,I1310084);
nor I_29556 (I504998,I504913,I504981);
nor I_29557 (I505015,I504905,I504998);
DFFARX1 I_29558 (I504964,I2507,I504831,I504820,);
nor I_29559 (I505046,I1310081,I1310072);
nand I_29560 (I505063,I505046,I1310096);
nor I_29561 (I505080,I505063,I504947);
nand I_29562 (I504805,I505080,I1310093);
DFFARX1 I_29563 (I505063,I2507,I504831,I504817,);
nand I_29564 (I505125,I504947,I1310081);
nor I_29565 (I505142,I504947,I1310081);
nand I_29566 (I504811,I504930,I505142);
not I_29567 (I505173,I1310090);
nor I_29568 (I505190,I505173,I505125);
DFFARX1 I_29569 (I505190,I2507,I504831,I504799,);
nor I_29570 (I505221,I505173,I1310075);
and I_29571 (I505238,I505221,I1310087);
or I_29572 (I505255,I505238,I1310099);
DFFARX1 I_29573 (I505255,I2507,I504831,I505281,);
nor I_29574 (I505289,I505281,I504905);
nor I_29575 (I504808,I504857,I505289);
not I_29576 (I505320,I505281);
nor I_29577 (I505337,I505320,I505015);
DFFARX1 I_29578 (I505337,I2507,I504831,I504814,);
nand I_29579 (I505368,I505320,I504947);
nor I_29580 (I504802,I505173,I505368);
not I_29581 (I505426,I2514);
DFFARX1 I_29582 (I425647,I2507,I505426,I505452,);
DFFARX1 I_29583 (I505452,I2507,I505426,I505469,);
not I_29584 (I505418,I505469);
DFFARX1 I_29585 (I425671,I2507,I505426,I505500,);
not I_29586 (I505508,I425650);
nor I_29587 (I505525,I505452,I505508);
not I_29588 (I505542,I425656);
not I_29589 (I505559,I425662);
nand I_29590 (I505576,I505559,I425656);
nor I_29591 (I505593,I505508,I505576);
nor I_29592 (I505610,I505500,I505593);
DFFARX1 I_29593 (I505559,I2507,I505426,I505415,);
nor I_29594 (I505641,I425662,I425674);
nand I_29595 (I505658,I505641,I425668);
nor I_29596 (I505675,I505658,I505542);
nand I_29597 (I505400,I505675,I425650);
DFFARX1 I_29598 (I505658,I2507,I505426,I505412,);
nand I_29599 (I505720,I505542,I425662);
nor I_29600 (I505737,I505542,I425662);
nand I_29601 (I505406,I505525,I505737);
not I_29602 (I505768,I425653);
nor I_29603 (I505785,I505768,I505720);
DFFARX1 I_29604 (I505785,I2507,I505426,I505394,);
nor I_29605 (I505816,I505768,I425647);
and I_29606 (I505833,I505816,I425665);
or I_29607 (I505850,I505833,I425659);
DFFARX1 I_29608 (I505850,I2507,I505426,I505876,);
nor I_29609 (I505884,I505876,I505500);
nor I_29610 (I505403,I505452,I505884);
not I_29611 (I505915,I505876);
nor I_29612 (I505932,I505915,I505610);
DFFARX1 I_29613 (I505932,I2507,I505426,I505409,);
nand I_29614 (I505963,I505915,I505542);
nor I_29615 (I505397,I505768,I505963);
not I_29616 (I506021,I2514);
DFFARX1 I_29617 (I899214,I2507,I506021,I506047,);
DFFARX1 I_29618 (I506047,I2507,I506021,I506064,);
not I_29619 (I506013,I506064);
DFFARX1 I_29620 (I899202,I2507,I506021,I506095,);
not I_29621 (I506103,I899199);
nor I_29622 (I506120,I506047,I506103);
not I_29623 (I506137,I899211);
not I_29624 (I506154,I899208);
nand I_29625 (I506171,I506154,I899211);
nor I_29626 (I506188,I506103,I506171);
nor I_29627 (I506205,I506095,I506188);
DFFARX1 I_29628 (I506154,I2507,I506021,I506010,);
nor I_29629 (I506236,I899208,I899217);
nand I_29630 (I506253,I506236,I899220);
nor I_29631 (I506270,I506253,I506137);
nand I_29632 (I505995,I506270,I899199);
DFFARX1 I_29633 (I506253,I2507,I506021,I506007,);
nand I_29634 (I506315,I506137,I899208);
nor I_29635 (I506332,I506137,I899208);
nand I_29636 (I506001,I506120,I506332);
not I_29637 (I506363,I899223);
nor I_29638 (I506380,I506363,I506315);
DFFARX1 I_29639 (I506380,I2507,I506021,I505989,);
nor I_29640 (I506411,I506363,I899226);
and I_29641 (I506428,I506411,I899205);
or I_29642 (I506445,I506428,I899199);
DFFARX1 I_29643 (I506445,I2507,I506021,I506471,);
nor I_29644 (I506479,I506471,I506095);
nor I_29645 (I505998,I506047,I506479);
not I_29646 (I506510,I506471);
nor I_29647 (I506527,I506510,I506205);
DFFARX1 I_29648 (I506527,I2507,I506021,I506004,);
nand I_29649 (I506558,I506510,I506137);
nor I_29650 (I505992,I506363,I506558);
not I_29651 (I506616,I2514);
DFFARX1 I_29652 (I135500,I2507,I506616,I506642,);
DFFARX1 I_29653 (I506642,I2507,I506616,I506659,);
not I_29654 (I506608,I506659);
DFFARX1 I_29655 (I135512,I2507,I506616,I506690,);
not I_29656 (I506698,I135503);
nor I_29657 (I506715,I506642,I506698);
not I_29658 (I506732,I135494);
not I_29659 (I506749,I135491);
nand I_29660 (I506766,I506749,I135494);
nor I_29661 (I506783,I506698,I506766);
nor I_29662 (I506800,I506690,I506783);
DFFARX1 I_29663 (I506749,I2507,I506616,I506605,);
nor I_29664 (I506831,I135491,I135491);
nand I_29665 (I506848,I506831,I135509);
nor I_29666 (I506865,I506848,I506732);
nand I_29667 (I506590,I506865,I135503);
DFFARX1 I_29668 (I506848,I2507,I506616,I506602,);
nand I_29669 (I506910,I506732,I135491);
nor I_29670 (I506927,I506732,I135491);
nand I_29671 (I506596,I506715,I506927);
not I_29672 (I506958,I135515);
nor I_29673 (I506975,I506958,I506910);
DFFARX1 I_29674 (I506975,I2507,I506616,I506584,);
nor I_29675 (I507006,I506958,I135494);
and I_29676 (I507023,I507006,I135497);
or I_29677 (I507040,I507023,I135506);
DFFARX1 I_29678 (I507040,I2507,I506616,I507066,);
nor I_29679 (I507074,I507066,I506690);
nor I_29680 (I506593,I506642,I507074);
not I_29681 (I507105,I507066);
nor I_29682 (I507122,I507105,I506800);
DFFARX1 I_29683 (I507122,I2507,I506616,I506599,);
nand I_29684 (I507153,I507105,I506732);
nor I_29685 (I506587,I506958,I507153);
not I_29686 (I507211,I2514);
DFFARX1 I_29687 (I1025288,I2507,I507211,I507237,);
DFFARX1 I_29688 (I507237,I2507,I507211,I507254,);
not I_29689 (I507203,I507254);
DFFARX1 I_29690 (I1025291,I2507,I507211,I507285,);
not I_29691 (I507293,I1025294);
nor I_29692 (I507310,I507237,I507293);
not I_29693 (I507327,I1025306);
not I_29694 (I507344,I1025297);
nand I_29695 (I507361,I507344,I1025306);
nor I_29696 (I507378,I507293,I507361);
nor I_29697 (I507395,I507285,I507378);
DFFARX1 I_29698 (I507344,I2507,I507211,I507200,);
nor I_29699 (I507426,I1025297,I1025303);
nand I_29700 (I507443,I507426,I1025291);
nor I_29701 (I507460,I507443,I507327);
nand I_29702 (I507185,I507460,I1025294);
DFFARX1 I_29703 (I507443,I2507,I507211,I507197,);
nand I_29704 (I507505,I507327,I1025297);
nor I_29705 (I507522,I507327,I1025297);
nand I_29706 (I507191,I507310,I507522);
not I_29707 (I507553,I1025294);
nor I_29708 (I507570,I507553,I507505);
DFFARX1 I_29709 (I507570,I2507,I507211,I507179,);
nor I_29710 (I507601,I507553,I1025300);
and I_29711 (I507618,I507601,I1025288);
or I_29712 (I507635,I507618,I1025309);
DFFARX1 I_29713 (I507635,I2507,I507211,I507661,);
nor I_29714 (I507669,I507661,I507285);
nor I_29715 (I507188,I507237,I507669);
not I_29716 (I507700,I507661);
nor I_29717 (I507717,I507700,I507395);
DFFARX1 I_29718 (I507717,I2507,I507211,I507194,);
nand I_29719 (I507748,I507700,I507327);
nor I_29720 (I507182,I507553,I507748);
not I_29721 (I507806,I2514);
DFFARX1 I_29722 (I1257075,I2507,I507806,I507832,);
DFFARX1 I_29723 (I507832,I2507,I507806,I507849,);
not I_29724 (I507798,I507849);
DFFARX1 I_29725 (I1257081,I2507,I507806,I507880,);
not I_29726 (I507888,I1257069);
nor I_29727 (I507905,I507832,I507888);
not I_29728 (I507922,I1257072);
not I_29729 (I507939,I1257078);
nand I_29730 (I507956,I507939,I1257072);
nor I_29731 (I507973,I507888,I507956);
nor I_29732 (I507990,I507880,I507973);
DFFARX1 I_29733 (I507939,I2507,I507806,I507795,);
nor I_29734 (I508021,I1257078,I1257069);
nand I_29735 (I508038,I508021,I1257087);
nor I_29736 (I508055,I508038,I507922);
nand I_29737 (I507780,I508055,I1257069);
DFFARX1 I_29738 (I508038,I2507,I507806,I507792,);
nand I_29739 (I508100,I507922,I1257078);
nor I_29740 (I508117,I507922,I1257078);
nand I_29741 (I507786,I507905,I508117);
not I_29742 (I508148,I1257066);
nor I_29743 (I508165,I508148,I508100);
DFFARX1 I_29744 (I508165,I2507,I507806,I507774,);
nor I_29745 (I508196,I508148,I1257090);
and I_29746 (I508213,I508196,I1257066);
or I_29747 (I508230,I508213,I1257084);
DFFARX1 I_29748 (I508230,I2507,I507806,I508256,);
nor I_29749 (I508264,I508256,I507880);
nor I_29750 (I507783,I507832,I508264);
not I_29751 (I508295,I508256);
nor I_29752 (I508312,I508295,I507990);
DFFARX1 I_29753 (I508312,I2507,I507806,I507789,);
nand I_29754 (I508343,I508295,I507922);
nor I_29755 (I507777,I508148,I508343);
not I_29756 (I508401,I2514);
DFFARX1 I_29757 (I586793,I2507,I508401,I508427,);
DFFARX1 I_29758 (I508427,I2507,I508401,I508444,);
not I_29759 (I508393,I508444);
DFFARX1 I_29760 (I586805,I2507,I508401,I508475,);
not I_29761 (I508483,I586790);
nor I_29762 (I508500,I508427,I508483);
not I_29763 (I508517,I586808);
not I_29764 (I508534,I586799);
nand I_29765 (I508551,I508534,I586808);
nor I_29766 (I508568,I508483,I508551);
nor I_29767 (I508585,I508475,I508568);
DFFARX1 I_29768 (I508534,I2507,I508401,I508390,);
nor I_29769 (I508616,I586799,I586811);
nand I_29770 (I508633,I508616,I586814);
nor I_29771 (I508650,I508633,I508517);
nand I_29772 (I508375,I508650,I586790);
DFFARX1 I_29773 (I508633,I2507,I508401,I508387,);
nand I_29774 (I508695,I508517,I586799);
nor I_29775 (I508712,I508517,I586799);
nand I_29776 (I508381,I508500,I508712);
not I_29777 (I508743,I586790);
nor I_29778 (I508760,I508743,I508695);
DFFARX1 I_29779 (I508760,I2507,I508401,I508369,);
nor I_29780 (I508791,I508743,I586802);
and I_29781 (I508808,I508791,I586796);
or I_29782 (I508825,I508808,I586793);
DFFARX1 I_29783 (I508825,I2507,I508401,I508851,);
nor I_29784 (I508859,I508851,I508475);
nor I_29785 (I508378,I508427,I508859);
not I_29786 (I508890,I508851);
nor I_29787 (I508907,I508890,I508585);
DFFARX1 I_29788 (I508907,I2507,I508401,I508384,);
nand I_29789 (I508938,I508890,I508517);
nor I_29790 (I508372,I508743,I508938);
not I_29791 (I508996,I2514);
DFFARX1 I_29792 (I1178034,I2507,I508996,I509022,);
DFFARX1 I_29793 (I509022,I2507,I508996,I509039,);
not I_29794 (I508988,I509039);
DFFARX1 I_29795 (I1178016,I2507,I508996,I509070,);
not I_29796 (I509078,I1178022);
nor I_29797 (I509095,I509022,I509078);
not I_29798 (I509112,I1178037);
not I_29799 (I509129,I1178028);
nand I_29800 (I509146,I509129,I1178037);
nor I_29801 (I509163,I509078,I509146);
nor I_29802 (I509180,I509070,I509163);
DFFARX1 I_29803 (I509129,I2507,I508996,I508985,);
nor I_29804 (I509211,I1178028,I1178040);
nand I_29805 (I509228,I509211,I1178019);
nor I_29806 (I509245,I509228,I509112);
nand I_29807 (I508970,I509245,I1178022);
DFFARX1 I_29808 (I509228,I2507,I508996,I508982,);
nand I_29809 (I509290,I509112,I1178028);
nor I_29810 (I509307,I509112,I1178028);
nand I_29811 (I508976,I509095,I509307);
not I_29812 (I509338,I1178025);
nor I_29813 (I509355,I509338,I509290);
DFFARX1 I_29814 (I509355,I2507,I508996,I508964,);
nor I_29815 (I509386,I509338,I1178031);
and I_29816 (I509403,I509386,I1178016);
or I_29817 (I509420,I509403,I1178019);
DFFARX1 I_29818 (I509420,I2507,I508996,I509446,);
nor I_29819 (I509454,I509446,I509070);
nor I_29820 (I508973,I509022,I509454);
not I_29821 (I509485,I509446);
nor I_29822 (I509502,I509485,I509180);
DFFARX1 I_29823 (I509502,I2507,I508996,I508979,);
nand I_29824 (I509533,I509485,I509112);
nor I_29825 (I508967,I509338,I509533);
not I_29826 (I509591,I2514);
DFFARX1 I_29827 (I406607,I2507,I509591,I509617,);
DFFARX1 I_29828 (I509617,I2507,I509591,I509634,);
not I_29829 (I509583,I509634);
DFFARX1 I_29830 (I406631,I2507,I509591,I509665,);
not I_29831 (I509673,I406610);
nor I_29832 (I509690,I509617,I509673);
not I_29833 (I509707,I406616);
not I_29834 (I509724,I406622);
nand I_29835 (I509741,I509724,I406616);
nor I_29836 (I509758,I509673,I509741);
nor I_29837 (I509775,I509665,I509758);
DFFARX1 I_29838 (I509724,I2507,I509591,I509580,);
nor I_29839 (I509806,I406622,I406634);
nand I_29840 (I509823,I509806,I406628);
nor I_29841 (I509840,I509823,I509707);
nand I_29842 (I509565,I509840,I406610);
DFFARX1 I_29843 (I509823,I2507,I509591,I509577,);
nand I_29844 (I509885,I509707,I406622);
nor I_29845 (I509902,I509707,I406622);
nand I_29846 (I509571,I509690,I509902);
not I_29847 (I509933,I406613);
nor I_29848 (I509950,I509933,I509885);
DFFARX1 I_29849 (I509950,I2507,I509591,I509559,);
nor I_29850 (I509981,I509933,I406607);
and I_29851 (I509998,I509981,I406625);
or I_29852 (I510015,I509998,I406619);
DFFARX1 I_29853 (I510015,I2507,I509591,I510041,);
nor I_29854 (I510049,I510041,I509665);
nor I_29855 (I509568,I509617,I510049);
not I_29856 (I510080,I510041);
nor I_29857 (I510097,I510080,I509775);
DFFARX1 I_29858 (I510097,I2507,I509591,I509574,);
nand I_29859 (I510128,I510080,I509707);
nor I_29860 (I509562,I509933,I510128);
not I_29861 (I510186,I2514);
DFFARX1 I_29862 (I252840,I2507,I510186,I510212,);
DFFARX1 I_29863 (I510212,I2507,I510186,I510229,);
not I_29864 (I510178,I510229);
DFFARX1 I_29865 (I252828,I2507,I510186,I510260,);
not I_29866 (I510268,I252831);
nor I_29867 (I510285,I510212,I510268);
not I_29868 (I510302,I252834);
not I_29869 (I510319,I252846);
nand I_29870 (I510336,I510319,I252834);
nor I_29871 (I510353,I510268,I510336);
nor I_29872 (I510370,I510260,I510353);
DFFARX1 I_29873 (I510319,I2507,I510186,I510175,);
nor I_29874 (I510401,I252846,I252837);
nand I_29875 (I510418,I510401,I252825);
nor I_29876 (I510435,I510418,I510302);
nand I_29877 (I510160,I510435,I252831);
DFFARX1 I_29878 (I510418,I2507,I510186,I510172,);
nand I_29879 (I510480,I510302,I252846);
nor I_29880 (I510497,I510302,I252846);
nand I_29881 (I510166,I510285,I510497);
not I_29882 (I510528,I252843);
nor I_29883 (I510545,I510528,I510480);
DFFARX1 I_29884 (I510545,I2507,I510186,I510154,);
nor I_29885 (I510576,I510528,I252849);
and I_29886 (I510593,I510576,I252852);
or I_29887 (I510610,I510593,I252825);
DFFARX1 I_29888 (I510610,I2507,I510186,I510636,);
nor I_29889 (I510644,I510636,I510260);
nor I_29890 (I510163,I510212,I510644);
not I_29891 (I510675,I510636);
nor I_29892 (I510692,I510675,I510370);
DFFARX1 I_29893 (I510692,I2507,I510186,I510169,);
nand I_29894 (I510723,I510675,I510302);
nor I_29895 (I510157,I510528,I510723);
not I_29896 (I510781,I2514);
DFFARX1 I_29897 (I239480,I2507,I510781,I510807,);
DFFARX1 I_29898 (I510807,I2507,I510781,I510824,);
not I_29899 (I510773,I510824);
DFFARX1 I_29900 (I239504,I2507,I510781,I510855,);
not I_29901 (I510863,I239498);
nor I_29902 (I510880,I510807,I510863);
not I_29903 (I510897,I239492);
not I_29904 (I510914,I239489);
nand I_29905 (I510931,I510914,I239492);
nor I_29906 (I510948,I510863,I510931);
nor I_29907 (I510965,I510855,I510948);
DFFARX1 I_29908 (I510914,I2507,I510781,I510770,);
nor I_29909 (I510996,I239489,I239483);
nand I_29910 (I511013,I510996,I239501);
nor I_29911 (I511030,I511013,I510897);
nand I_29912 (I510755,I511030,I239498);
DFFARX1 I_29913 (I511013,I2507,I510781,I510767,);
nand I_29914 (I511075,I510897,I239489);
nor I_29915 (I511092,I510897,I239489);
nand I_29916 (I510761,I510880,I511092);
not I_29917 (I511123,I239495);
nor I_29918 (I511140,I511123,I511075);
DFFARX1 I_29919 (I511140,I2507,I510781,I510749,);
nor I_29920 (I511171,I511123,I239480);
and I_29921 (I511188,I511171,I239486);
or I_29922 (I511205,I511188,I239483);
DFFARX1 I_29923 (I511205,I2507,I510781,I511231,);
nor I_29924 (I511239,I511231,I510855);
nor I_29925 (I510758,I510807,I511239);
not I_29926 (I511270,I511231);
nor I_29927 (I511287,I511270,I510965);
DFFARX1 I_29928 (I511287,I2507,I510781,I510764,);
nand I_29929 (I511318,I511270,I510897);
nor I_29930 (I510752,I511123,I511318);
not I_29931 (I511376,I2514);
DFFARX1 I_29932 (I297635,I2507,I511376,I511402,);
DFFARX1 I_29933 (I511402,I2507,I511376,I511419,);
not I_29934 (I511368,I511419);
DFFARX1 I_29935 (I297623,I2507,I511376,I511450,);
not I_29936 (I511458,I297626);
nor I_29937 (I511475,I511402,I511458);
not I_29938 (I511492,I297629);
not I_29939 (I511509,I297641);
nand I_29940 (I511526,I511509,I297629);
nor I_29941 (I511543,I511458,I511526);
nor I_29942 (I511560,I511450,I511543);
DFFARX1 I_29943 (I511509,I2507,I511376,I511365,);
nor I_29944 (I511591,I297641,I297632);
nand I_29945 (I511608,I511591,I297620);
nor I_29946 (I511625,I511608,I511492);
nand I_29947 (I511350,I511625,I297626);
DFFARX1 I_29948 (I511608,I2507,I511376,I511362,);
nand I_29949 (I511670,I511492,I297641);
nor I_29950 (I511687,I511492,I297641);
nand I_29951 (I511356,I511475,I511687);
not I_29952 (I511718,I297638);
nor I_29953 (I511735,I511718,I511670);
DFFARX1 I_29954 (I511735,I2507,I511376,I511344,);
nor I_29955 (I511766,I511718,I297644);
and I_29956 (I511783,I511766,I297647);
or I_29957 (I511800,I511783,I297620);
DFFARX1 I_29958 (I511800,I2507,I511376,I511826,);
nor I_29959 (I511834,I511826,I511450);
nor I_29960 (I511353,I511402,I511834);
not I_29961 (I511865,I511826);
nor I_29962 (I511882,I511865,I511560);
DFFARX1 I_29963 (I511882,I2507,I511376,I511359,);
nand I_29964 (I511913,I511865,I511492);
nor I_29965 (I511347,I511718,I511913);
not I_29966 (I511971,I2514);
DFFARX1 I_29967 (I296054,I2507,I511971,I511997,);
DFFARX1 I_29968 (I511997,I2507,I511971,I512014,);
not I_29969 (I511963,I512014);
DFFARX1 I_29970 (I296042,I2507,I511971,I512045,);
not I_29971 (I512053,I296045);
nor I_29972 (I512070,I511997,I512053);
not I_29973 (I512087,I296048);
not I_29974 (I512104,I296060);
nand I_29975 (I512121,I512104,I296048);
nor I_29976 (I512138,I512053,I512121);
nor I_29977 (I512155,I512045,I512138);
DFFARX1 I_29978 (I512104,I2507,I511971,I511960,);
nor I_29979 (I512186,I296060,I296051);
nand I_29980 (I512203,I512186,I296039);
nor I_29981 (I512220,I512203,I512087);
nand I_29982 (I511945,I512220,I296045);
DFFARX1 I_29983 (I512203,I2507,I511971,I511957,);
nand I_29984 (I512265,I512087,I296060);
nor I_29985 (I512282,I512087,I296060);
nand I_29986 (I511951,I512070,I512282);
not I_29987 (I512313,I296057);
nor I_29988 (I512330,I512313,I512265);
DFFARX1 I_29989 (I512330,I2507,I511971,I511939,);
nor I_29990 (I512361,I512313,I296063);
and I_29991 (I512378,I512361,I296066);
or I_29992 (I512395,I512378,I296039);
DFFARX1 I_29993 (I512395,I2507,I511971,I512421,);
nor I_29994 (I512429,I512421,I512045);
nor I_29995 (I511948,I511997,I512429);
not I_29996 (I512460,I512421);
nor I_29997 (I512477,I512460,I512155);
DFFARX1 I_29998 (I512477,I2507,I511971,I511954,);
nand I_29999 (I512508,I512460,I512087);
nor I_30000 (I511942,I512313,I512508);
not I_30001 (I512566,I2514);
DFFARX1 I_30002 (I1213410,I2507,I512566,I512592,);
DFFARX1 I_30003 (I512592,I2507,I512566,I512609,);
not I_30004 (I512558,I512609);
DFFARX1 I_30005 (I1213425,I2507,I512566,I512640,);
not I_30006 (I512648,I1213434);
nor I_30007 (I512665,I512592,I512648);
not I_30008 (I512682,I1213413);
not I_30009 (I512699,I1213419);
nand I_30010 (I512716,I512699,I1213413);
nor I_30011 (I512733,I512648,I512716);
nor I_30012 (I512750,I512640,I512733);
DFFARX1 I_30013 (I512699,I2507,I512566,I512555,);
nor I_30014 (I512781,I1213419,I1213431);
nand I_30015 (I512798,I512781,I1213428);
nor I_30016 (I512815,I512798,I512682);
nand I_30017 (I512540,I512815,I1213434);
DFFARX1 I_30018 (I512798,I2507,I512566,I512552,);
nand I_30019 (I512860,I512682,I1213419);
nor I_30020 (I512877,I512682,I1213419);
nand I_30021 (I512546,I512665,I512877);
not I_30022 (I512908,I1213410);
nor I_30023 (I512925,I512908,I512860);
DFFARX1 I_30024 (I512925,I2507,I512566,I512534,);
nor I_30025 (I512956,I512908,I1213422);
and I_30026 (I512973,I512956,I1213416);
or I_30027 (I512990,I512973,I1213413);
DFFARX1 I_30028 (I512990,I2507,I512566,I513016,);
nor I_30029 (I513024,I513016,I512640);
nor I_30030 (I512543,I512592,I513024);
not I_30031 (I513055,I513016);
nor I_30032 (I513072,I513055,I512750);
DFFARX1 I_30033 (I513072,I2507,I512566,I512549,);
nand I_30034 (I513103,I513055,I512682);
nor I_30035 (I512537,I512908,I513103);
not I_30036 (I513161,I2514);
DFFARX1 I_30037 (I268650,I2507,I513161,I513187,);
DFFARX1 I_30038 (I513187,I2507,I513161,I513204,);
not I_30039 (I513153,I513204);
DFFARX1 I_30040 (I268638,I2507,I513161,I513235,);
not I_30041 (I513243,I268641);
nor I_30042 (I513260,I513187,I513243);
not I_30043 (I513277,I268644);
not I_30044 (I513294,I268656);
nand I_30045 (I513311,I513294,I268644);
nor I_30046 (I513328,I513243,I513311);
nor I_30047 (I513345,I513235,I513328);
DFFARX1 I_30048 (I513294,I2507,I513161,I513150,);
nor I_30049 (I513376,I268656,I268647);
nand I_30050 (I513393,I513376,I268635);
nor I_30051 (I513410,I513393,I513277);
nand I_30052 (I513135,I513410,I268641);
DFFARX1 I_30053 (I513393,I2507,I513161,I513147,);
nand I_30054 (I513455,I513277,I268656);
nor I_30055 (I513472,I513277,I268656);
nand I_30056 (I513141,I513260,I513472);
not I_30057 (I513503,I268653);
nor I_30058 (I513520,I513503,I513455);
DFFARX1 I_30059 (I513520,I2507,I513161,I513129,);
nor I_30060 (I513551,I513503,I268659);
and I_30061 (I513568,I513551,I268662);
or I_30062 (I513585,I513568,I268635);
DFFARX1 I_30063 (I513585,I2507,I513161,I513611,);
nor I_30064 (I513619,I513611,I513235);
nor I_30065 (I513138,I513187,I513619);
not I_30066 (I513650,I513611);
nor I_30067 (I513667,I513650,I513345);
DFFARX1 I_30068 (I513667,I2507,I513161,I513144,);
nand I_30069 (I513698,I513650,I513277);
nor I_30070 (I513132,I513503,I513698);
not I_30071 (I513756,I2514);
DFFARX1 I_30072 (I1377902,I2507,I513756,I513782,);
DFFARX1 I_30073 (I513782,I2507,I513756,I513799,);
not I_30074 (I513748,I513799);
DFFARX1 I_30075 (I1377908,I2507,I513756,I513830,);
not I_30076 (I513838,I1377923);
nor I_30077 (I513855,I513782,I513838);
not I_30078 (I513872,I1377914);
not I_30079 (I513889,I1377911);
nand I_30080 (I513906,I513889,I1377914);
nor I_30081 (I513923,I513838,I513906);
nor I_30082 (I513940,I513830,I513923);
DFFARX1 I_30083 (I513889,I2507,I513756,I513745,);
nor I_30084 (I513971,I1377911,I1377902);
nand I_30085 (I513988,I513971,I1377926);
nor I_30086 (I514005,I513988,I513872);
nand I_30087 (I513730,I514005,I1377923);
DFFARX1 I_30088 (I513988,I2507,I513756,I513742,);
nand I_30089 (I514050,I513872,I1377911);
nor I_30090 (I514067,I513872,I1377911);
nand I_30091 (I513736,I513855,I514067);
not I_30092 (I514098,I1377920);
nor I_30093 (I514115,I514098,I514050);
DFFARX1 I_30094 (I514115,I2507,I513756,I513724,);
nor I_30095 (I514146,I514098,I1377905);
and I_30096 (I514163,I514146,I1377917);
or I_30097 (I514180,I514163,I1377929);
DFFARX1 I_30098 (I514180,I2507,I513756,I514206,);
nor I_30099 (I514214,I514206,I513830);
nor I_30100 (I513733,I513782,I514214);
not I_30101 (I514245,I514206);
nor I_30102 (I514262,I514245,I513940);
DFFARX1 I_30103 (I514262,I2507,I513756,I513739,);
nand I_30104 (I514293,I514245,I513872);
nor I_30105 (I513727,I514098,I514293);
not I_30106 (I514351,I2514);
DFFARX1 I_30107 (I28510,I2507,I514351,I514377,);
DFFARX1 I_30108 (I514377,I2507,I514351,I514394,);
not I_30109 (I514343,I514394);
DFFARX1 I_30110 (I28510,I2507,I514351,I514425,);
not I_30111 (I514433,I28525);
nor I_30112 (I514450,I514377,I514433);
not I_30113 (I514467,I28528);
not I_30114 (I514484,I28519);
nand I_30115 (I514501,I514484,I28528);
nor I_30116 (I514518,I514433,I514501);
nor I_30117 (I514535,I514425,I514518);
DFFARX1 I_30118 (I514484,I2507,I514351,I514340,);
nor I_30119 (I514566,I28519,I28531);
nand I_30120 (I514583,I514566,I28513);
nor I_30121 (I514600,I514583,I514467);
nand I_30122 (I514325,I514600,I28525);
DFFARX1 I_30123 (I514583,I2507,I514351,I514337,);
nand I_30124 (I514645,I514467,I28519);
nor I_30125 (I514662,I514467,I28519);
nand I_30126 (I514331,I514450,I514662);
not I_30127 (I514693,I28513);
nor I_30128 (I514710,I514693,I514645);
DFFARX1 I_30129 (I514710,I2507,I514351,I514319,);
nor I_30130 (I514741,I514693,I28522);
and I_30131 (I514758,I514741,I28516);
or I_30132 (I514775,I514758,I28534);
DFFARX1 I_30133 (I514775,I2507,I514351,I514801,);
nor I_30134 (I514809,I514801,I514425);
nor I_30135 (I514328,I514377,I514809);
not I_30136 (I514840,I514801);
nor I_30137 (I514857,I514840,I514535);
DFFARX1 I_30138 (I514857,I2507,I514351,I514334,);
nand I_30139 (I514888,I514840,I514467);
nor I_30140 (I514322,I514693,I514888);
not I_30141 (I514946,I2514);
DFFARX1 I_30142 (I318715,I2507,I514946,I514972,);
DFFARX1 I_30143 (I514972,I2507,I514946,I514989,);
not I_30144 (I514938,I514989);
DFFARX1 I_30145 (I318703,I2507,I514946,I515020,);
not I_30146 (I515028,I318706);
nor I_30147 (I515045,I514972,I515028);
not I_30148 (I515062,I318709);
not I_30149 (I515079,I318721);
nand I_30150 (I515096,I515079,I318709);
nor I_30151 (I515113,I515028,I515096);
nor I_30152 (I515130,I515020,I515113);
DFFARX1 I_30153 (I515079,I2507,I514946,I514935,);
nor I_30154 (I515161,I318721,I318712);
nand I_30155 (I515178,I515161,I318700);
nor I_30156 (I515195,I515178,I515062);
nand I_30157 (I514920,I515195,I318706);
DFFARX1 I_30158 (I515178,I2507,I514946,I514932,);
nand I_30159 (I515240,I515062,I318721);
nor I_30160 (I515257,I515062,I318721);
nand I_30161 (I514926,I515045,I515257);
not I_30162 (I515288,I318718);
nor I_30163 (I515305,I515288,I515240);
DFFARX1 I_30164 (I515305,I2507,I514946,I514914,);
nor I_30165 (I515336,I515288,I318724);
and I_30166 (I515353,I515336,I318727);
or I_30167 (I515370,I515353,I318700);
DFFARX1 I_30168 (I515370,I2507,I514946,I515396,);
nor I_30169 (I515404,I515396,I515020);
nor I_30170 (I514923,I514972,I515404);
not I_30171 (I515435,I515396);
nor I_30172 (I515452,I515435,I515130);
DFFARX1 I_30173 (I515452,I2507,I514946,I514929,);
nand I_30174 (I515483,I515435,I515062);
nor I_30175 (I514917,I515288,I515483);
not I_30176 (I515541,I2514);
DFFARX1 I_30177 (I682169,I2507,I515541,I515567,);
DFFARX1 I_30178 (I515567,I2507,I515541,I515584,);
not I_30179 (I515533,I515584);
DFFARX1 I_30180 (I682163,I2507,I515541,I515615,);
not I_30181 (I515623,I682160);
nor I_30182 (I515640,I515567,I515623);
not I_30183 (I515657,I682172);
not I_30184 (I515674,I682175);
nand I_30185 (I515691,I515674,I682172);
nor I_30186 (I515708,I515623,I515691);
nor I_30187 (I515725,I515615,I515708);
DFFARX1 I_30188 (I515674,I2507,I515541,I515530,);
nor I_30189 (I515756,I682175,I682184);
nand I_30190 (I515773,I515756,I682178);
nor I_30191 (I515790,I515773,I515657);
nand I_30192 (I515515,I515790,I682160);
DFFARX1 I_30193 (I515773,I2507,I515541,I515527,);
nand I_30194 (I515835,I515657,I682175);
nor I_30195 (I515852,I515657,I682175);
nand I_30196 (I515521,I515640,I515852);
not I_30197 (I515883,I682166);
nor I_30198 (I515900,I515883,I515835);
DFFARX1 I_30199 (I515900,I2507,I515541,I515509,);
nor I_30200 (I515931,I515883,I682181);
and I_30201 (I515948,I515931,I682160);
or I_30202 (I515965,I515948,I682163);
DFFARX1 I_30203 (I515965,I2507,I515541,I515991,);
nor I_30204 (I515999,I515991,I515615);
nor I_30205 (I515518,I515567,I515999);
not I_30206 (I516030,I515991);
nor I_30207 (I516047,I516030,I515725);
DFFARX1 I_30208 (I516047,I2507,I515541,I515524,);
nand I_30209 (I516078,I516030,I515657);
nor I_30210 (I515512,I515883,I516078);
not I_30211 (I516136,I2514);
DFFARX1 I_30212 (I910842,I2507,I516136,I516162,);
DFFARX1 I_30213 (I516162,I2507,I516136,I516179,);
not I_30214 (I516128,I516179);
DFFARX1 I_30215 (I910830,I2507,I516136,I516210,);
not I_30216 (I516218,I910827);
nor I_30217 (I516235,I516162,I516218);
not I_30218 (I516252,I910839);
not I_30219 (I516269,I910836);
nand I_30220 (I516286,I516269,I910839);
nor I_30221 (I516303,I516218,I516286);
nor I_30222 (I516320,I516210,I516303);
DFFARX1 I_30223 (I516269,I2507,I516136,I516125,);
nor I_30224 (I516351,I910836,I910845);
nand I_30225 (I516368,I516351,I910848);
nor I_30226 (I516385,I516368,I516252);
nand I_30227 (I516110,I516385,I910827);
DFFARX1 I_30228 (I516368,I2507,I516136,I516122,);
nand I_30229 (I516430,I516252,I910836);
nor I_30230 (I516447,I516252,I910836);
nand I_30231 (I516116,I516235,I516447);
not I_30232 (I516478,I910851);
nor I_30233 (I516495,I516478,I516430);
DFFARX1 I_30234 (I516495,I2507,I516136,I516104,);
nor I_30235 (I516526,I516478,I910854);
and I_30236 (I516543,I516526,I910833);
or I_30237 (I516560,I516543,I910827);
DFFARX1 I_30238 (I516560,I2507,I516136,I516586,);
nor I_30239 (I516594,I516586,I516210);
nor I_30240 (I516113,I516162,I516594);
not I_30241 (I516625,I516586);
nor I_30242 (I516642,I516625,I516320);
DFFARX1 I_30243 (I516642,I2507,I516136,I516119,);
nand I_30244 (I516673,I516625,I516252);
nor I_30245 (I516107,I516478,I516673);
not I_30246 (I516731,I2514);
DFFARX1 I_30247 (I1327327,I2507,I516731,I516757,);
DFFARX1 I_30248 (I516757,I2507,I516731,I516774,);
not I_30249 (I516723,I516774);
DFFARX1 I_30250 (I1327333,I2507,I516731,I516805,);
not I_30251 (I516813,I1327348);
nor I_30252 (I516830,I516757,I516813);
not I_30253 (I516847,I1327339);
not I_30254 (I516864,I1327336);
nand I_30255 (I516881,I516864,I1327339);
nor I_30256 (I516898,I516813,I516881);
nor I_30257 (I516915,I516805,I516898);
DFFARX1 I_30258 (I516864,I2507,I516731,I516720,);
nor I_30259 (I516946,I1327336,I1327327);
nand I_30260 (I516963,I516946,I1327351);
nor I_30261 (I516980,I516963,I516847);
nand I_30262 (I516705,I516980,I1327348);
DFFARX1 I_30263 (I516963,I2507,I516731,I516717,);
nand I_30264 (I517025,I516847,I1327336);
nor I_30265 (I517042,I516847,I1327336);
nand I_30266 (I516711,I516830,I517042);
not I_30267 (I517073,I1327345);
nor I_30268 (I517090,I517073,I517025);
DFFARX1 I_30269 (I517090,I2507,I516731,I516699,);
nor I_30270 (I517121,I517073,I1327330);
and I_30271 (I517138,I517121,I1327342);
or I_30272 (I517155,I517138,I1327354);
DFFARX1 I_30273 (I517155,I2507,I516731,I517181,);
nor I_30274 (I517189,I517181,I516805);
nor I_30275 (I516708,I516757,I517189);
not I_30276 (I517220,I517181);
nor I_30277 (I517237,I517220,I516915);
DFFARX1 I_30278 (I517237,I2507,I516731,I516714,);
nand I_30279 (I517268,I517220,I516847);
nor I_30280 (I516702,I517073,I517268);
not I_30281 (I517326,I2514);
DFFARX1 I_30282 (I1318402,I2507,I517326,I517352,);
DFFARX1 I_30283 (I517352,I2507,I517326,I517369,);
not I_30284 (I517318,I517369);
DFFARX1 I_30285 (I1318408,I2507,I517326,I517400,);
not I_30286 (I517408,I1318423);
nor I_30287 (I517425,I517352,I517408);
not I_30288 (I517442,I1318414);
not I_30289 (I517459,I1318411);
nand I_30290 (I517476,I517459,I1318414);
nor I_30291 (I517493,I517408,I517476);
nor I_30292 (I517510,I517400,I517493);
DFFARX1 I_30293 (I517459,I2507,I517326,I517315,);
nor I_30294 (I517541,I1318411,I1318402);
nand I_30295 (I517558,I517541,I1318426);
nor I_30296 (I517575,I517558,I517442);
nand I_30297 (I517300,I517575,I1318423);
DFFARX1 I_30298 (I517558,I2507,I517326,I517312,);
nand I_30299 (I517620,I517442,I1318411);
nor I_30300 (I517637,I517442,I1318411);
nand I_30301 (I517306,I517425,I517637);
not I_30302 (I517668,I1318420);
nor I_30303 (I517685,I517668,I517620);
DFFARX1 I_30304 (I517685,I2507,I517326,I517294,);
nor I_30305 (I517716,I517668,I1318405);
and I_30306 (I517733,I517716,I1318417);
or I_30307 (I517750,I517733,I1318429);
DFFARX1 I_30308 (I517750,I2507,I517326,I517776,);
nor I_30309 (I517784,I517776,I517400);
nor I_30310 (I517303,I517352,I517784);
not I_30311 (I517815,I517776);
nor I_30312 (I517832,I517815,I517510);
DFFARX1 I_30313 (I517832,I2507,I517326,I517309,);
nand I_30314 (I517863,I517815,I517442);
nor I_30315 (I517297,I517668,I517863);
not I_30316 (I517921,I2514);
DFFARX1 I_30317 (I1183814,I2507,I517921,I517947,);
DFFARX1 I_30318 (I517947,I2507,I517921,I517964,);
not I_30319 (I517913,I517964);
DFFARX1 I_30320 (I1183796,I2507,I517921,I517995,);
not I_30321 (I518003,I1183802);
nor I_30322 (I518020,I517947,I518003);
not I_30323 (I518037,I1183817);
not I_30324 (I518054,I1183808);
nand I_30325 (I518071,I518054,I1183817);
nor I_30326 (I518088,I518003,I518071);
nor I_30327 (I518105,I517995,I518088);
DFFARX1 I_30328 (I518054,I2507,I517921,I517910,);
nor I_30329 (I518136,I1183808,I1183820);
nand I_30330 (I518153,I518136,I1183799);
nor I_30331 (I518170,I518153,I518037);
nand I_30332 (I517895,I518170,I1183802);
DFFARX1 I_30333 (I518153,I2507,I517921,I517907,);
nand I_30334 (I518215,I518037,I1183808);
nor I_30335 (I518232,I518037,I1183808);
nand I_30336 (I517901,I518020,I518232);
not I_30337 (I518263,I1183805);
nor I_30338 (I518280,I518263,I518215);
DFFARX1 I_30339 (I518280,I2507,I517921,I517889,);
nor I_30340 (I518311,I518263,I1183811);
and I_30341 (I518328,I518311,I1183796);
or I_30342 (I518345,I518328,I1183799);
DFFARX1 I_30343 (I518345,I2507,I517921,I518371,);
nor I_30344 (I518379,I518371,I517995);
nor I_30345 (I517898,I517947,I518379);
not I_30346 (I518410,I518371);
nor I_30347 (I518427,I518410,I518105);
DFFARX1 I_30348 (I518427,I2507,I517921,I517904,);
nand I_30349 (I518458,I518410,I518037);
nor I_30350 (I517892,I518263,I518458);
not I_30351 (I518516,I2514);
DFFARX1 I_30352 (I1237346,I2507,I518516,I518542,);
DFFARX1 I_30353 (I518542,I2507,I518516,I518559,);
not I_30354 (I518508,I518559);
DFFARX1 I_30355 (I1237361,I2507,I518516,I518590,);
not I_30356 (I518598,I1237370);
nor I_30357 (I518615,I518542,I518598);
not I_30358 (I518632,I1237349);
not I_30359 (I518649,I1237355);
nand I_30360 (I518666,I518649,I1237349);
nor I_30361 (I518683,I518598,I518666);
nor I_30362 (I518700,I518590,I518683);
DFFARX1 I_30363 (I518649,I2507,I518516,I518505,);
nor I_30364 (I518731,I1237355,I1237367);
nand I_30365 (I518748,I518731,I1237364);
nor I_30366 (I518765,I518748,I518632);
nand I_30367 (I518490,I518765,I1237370);
DFFARX1 I_30368 (I518748,I2507,I518516,I518502,);
nand I_30369 (I518810,I518632,I1237355);
nor I_30370 (I518827,I518632,I1237355);
nand I_30371 (I518496,I518615,I518827);
not I_30372 (I518858,I1237346);
nor I_30373 (I518875,I518858,I518810);
DFFARX1 I_30374 (I518875,I2507,I518516,I518484,);
nor I_30375 (I518906,I518858,I1237358);
and I_30376 (I518923,I518906,I1237352);
or I_30377 (I518940,I518923,I1237349);
DFFARX1 I_30378 (I518940,I2507,I518516,I518966,);
nor I_30379 (I518974,I518966,I518590);
nor I_30380 (I518493,I518542,I518974);
not I_30381 (I519005,I518966);
nor I_30382 (I519022,I519005,I518700);
DFFARX1 I_30383 (I519022,I2507,I518516,I518499,);
nand I_30384 (I519053,I519005,I518632);
nor I_30385 (I518487,I518858,I519053);
not I_30386 (I519111,I2514);
DFFARX1 I_30387 (I218655,I2507,I519111,I519137,);
DFFARX1 I_30388 (I519137,I2507,I519111,I519154,);
not I_30389 (I519103,I519154);
DFFARX1 I_30390 (I218679,I2507,I519111,I519185,);
not I_30391 (I519193,I218673);
nor I_30392 (I519210,I519137,I519193);
not I_30393 (I519227,I218667);
not I_30394 (I519244,I218664);
nand I_30395 (I519261,I519244,I218667);
nor I_30396 (I519278,I519193,I519261);
nor I_30397 (I519295,I519185,I519278);
DFFARX1 I_30398 (I519244,I2507,I519111,I519100,);
nor I_30399 (I519326,I218664,I218658);
nand I_30400 (I519343,I519326,I218676);
nor I_30401 (I519360,I519343,I519227);
nand I_30402 (I519085,I519360,I218673);
DFFARX1 I_30403 (I519343,I2507,I519111,I519097,);
nand I_30404 (I519405,I519227,I218664);
nor I_30405 (I519422,I519227,I218664);
nand I_30406 (I519091,I519210,I519422);
not I_30407 (I519453,I218670);
nor I_30408 (I519470,I519453,I519405);
DFFARX1 I_30409 (I519470,I2507,I519111,I519079,);
nor I_30410 (I519501,I519453,I218655);
and I_30411 (I519518,I519501,I218661);
or I_30412 (I519535,I519518,I218658);
DFFARX1 I_30413 (I519535,I2507,I519111,I519561,);
nor I_30414 (I519569,I519561,I519185);
nor I_30415 (I519088,I519137,I519569);
not I_30416 (I519600,I519561);
nor I_30417 (I519617,I519600,I519295);
DFFARX1 I_30418 (I519617,I2507,I519111,I519094,);
nand I_30419 (I519648,I519600,I519227);
nor I_30420 (I519082,I519453,I519648);
not I_30421 (I519706,I2514);
DFFARX1 I_30422 (I665407,I2507,I519706,I519732,);
DFFARX1 I_30423 (I519732,I2507,I519706,I519749,);
not I_30424 (I519698,I519749);
DFFARX1 I_30425 (I665401,I2507,I519706,I519780,);
not I_30426 (I519788,I665398);
nor I_30427 (I519805,I519732,I519788);
not I_30428 (I519822,I665410);
not I_30429 (I519839,I665413);
nand I_30430 (I519856,I519839,I665410);
nor I_30431 (I519873,I519788,I519856);
nor I_30432 (I519890,I519780,I519873);
DFFARX1 I_30433 (I519839,I2507,I519706,I519695,);
nor I_30434 (I519921,I665413,I665422);
nand I_30435 (I519938,I519921,I665416);
nor I_30436 (I519955,I519938,I519822);
nand I_30437 (I519680,I519955,I665398);
DFFARX1 I_30438 (I519938,I2507,I519706,I519692,);
nand I_30439 (I520000,I519822,I665413);
nor I_30440 (I520017,I519822,I665413);
nand I_30441 (I519686,I519805,I520017);
not I_30442 (I520048,I665404);
nor I_30443 (I520065,I520048,I520000);
DFFARX1 I_30444 (I520065,I2507,I519706,I519674,);
nor I_30445 (I520096,I520048,I665419);
and I_30446 (I520113,I520096,I665398);
or I_30447 (I520130,I520113,I665401);
DFFARX1 I_30448 (I520130,I2507,I519706,I520156,);
nor I_30449 (I520164,I520156,I519780);
nor I_30450 (I519683,I519732,I520164);
not I_30451 (I520195,I520156);
nor I_30452 (I520212,I520195,I519890);
DFFARX1 I_30453 (I520212,I2507,I519706,I519689,);
nand I_30454 (I520243,I520195,I519822);
nor I_30455 (I519677,I520048,I520243);
not I_30456 (I520301,I2514);
DFFARX1 I_30457 (I421295,I2507,I520301,I520327,);
DFFARX1 I_30458 (I520327,I2507,I520301,I520344,);
not I_30459 (I520293,I520344);
DFFARX1 I_30460 (I421319,I2507,I520301,I520375,);
not I_30461 (I520383,I421298);
nor I_30462 (I520400,I520327,I520383);
not I_30463 (I520417,I421304);
not I_30464 (I520434,I421310);
nand I_30465 (I520451,I520434,I421304);
nor I_30466 (I520468,I520383,I520451);
nor I_30467 (I520485,I520375,I520468);
DFFARX1 I_30468 (I520434,I2507,I520301,I520290,);
nor I_30469 (I520516,I421310,I421322);
nand I_30470 (I520533,I520516,I421316);
nor I_30471 (I520550,I520533,I520417);
nand I_30472 (I520275,I520550,I421298);
DFFARX1 I_30473 (I520533,I2507,I520301,I520287,);
nand I_30474 (I520595,I520417,I421310);
nor I_30475 (I520612,I520417,I421310);
nand I_30476 (I520281,I520400,I520612);
not I_30477 (I520643,I421301);
nor I_30478 (I520660,I520643,I520595);
DFFARX1 I_30479 (I520660,I2507,I520301,I520269,);
nor I_30480 (I520691,I520643,I421295);
and I_30481 (I520708,I520691,I421313);
or I_30482 (I520725,I520708,I421307);
DFFARX1 I_30483 (I520725,I2507,I520301,I520751,);
nor I_30484 (I520759,I520751,I520375);
nor I_30485 (I520278,I520327,I520759);
not I_30486 (I520790,I520751);
nor I_30487 (I520807,I520790,I520485);
DFFARX1 I_30488 (I520807,I2507,I520301,I520284,);
nand I_30489 (I520838,I520790,I520417);
nor I_30490 (I520272,I520643,I520838);
not I_30491 (I520896,I2514);
DFFARX1 I_30492 (I120217,I2507,I520896,I520922,);
DFFARX1 I_30493 (I520922,I2507,I520896,I520939,);
not I_30494 (I520888,I520939);
DFFARX1 I_30495 (I120229,I2507,I520896,I520970,);
not I_30496 (I520978,I120220);
nor I_30497 (I520995,I520922,I520978);
not I_30498 (I521012,I120211);
not I_30499 (I521029,I120208);
nand I_30500 (I521046,I521029,I120211);
nor I_30501 (I521063,I520978,I521046);
nor I_30502 (I521080,I520970,I521063);
DFFARX1 I_30503 (I521029,I2507,I520896,I520885,);
nor I_30504 (I521111,I120208,I120208);
nand I_30505 (I521128,I521111,I120226);
nor I_30506 (I521145,I521128,I521012);
nand I_30507 (I520870,I521145,I120220);
DFFARX1 I_30508 (I521128,I2507,I520896,I520882,);
nand I_30509 (I521190,I521012,I120208);
nor I_30510 (I521207,I521012,I120208);
nand I_30511 (I520876,I520995,I521207);
not I_30512 (I521238,I120232);
nor I_30513 (I521255,I521238,I521190);
DFFARX1 I_30514 (I521255,I2507,I520896,I520864,);
nor I_30515 (I521286,I521238,I120211);
and I_30516 (I521303,I521286,I120214);
or I_30517 (I521320,I521303,I120223);
DFFARX1 I_30518 (I521320,I2507,I520896,I521346,);
nor I_30519 (I521354,I521346,I520970);
nor I_30520 (I520873,I520922,I521354);
not I_30521 (I521385,I521346);
nor I_30522 (I521402,I521385,I521080);
DFFARX1 I_30523 (I521402,I2507,I520896,I520879,);
nand I_30524 (I521433,I521385,I521012);
nor I_30525 (I520867,I521238,I521433);
not I_30526 (I521491,I2514);
DFFARX1 I_30527 (I112839,I2507,I521491,I521517,);
DFFARX1 I_30528 (I521517,I2507,I521491,I521534,);
not I_30529 (I521483,I521534);
DFFARX1 I_30530 (I112851,I2507,I521491,I521565,);
not I_30531 (I521573,I112842);
nor I_30532 (I521590,I521517,I521573);
not I_30533 (I521607,I112833);
not I_30534 (I521624,I112830);
nand I_30535 (I521641,I521624,I112833);
nor I_30536 (I521658,I521573,I521641);
nor I_30537 (I521675,I521565,I521658);
DFFARX1 I_30538 (I521624,I2507,I521491,I521480,);
nor I_30539 (I521706,I112830,I112830);
nand I_30540 (I521723,I521706,I112848);
nor I_30541 (I521740,I521723,I521607);
nand I_30542 (I521465,I521740,I112842);
DFFARX1 I_30543 (I521723,I2507,I521491,I521477,);
nand I_30544 (I521785,I521607,I112830);
nor I_30545 (I521802,I521607,I112830);
nand I_30546 (I521471,I521590,I521802);
not I_30547 (I521833,I112854);
nor I_30548 (I521850,I521833,I521785);
DFFARX1 I_30549 (I521850,I2507,I521491,I521459,);
nor I_30550 (I521881,I521833,I112833);
and I_30551 (I521898,I521881,I112836);
or I_30552 (I521915,I521898,I112845);
DFFARX1 I_30553 (I521915,I2507,I521491,I521941,);
nor I_30554 (I521949,I521941,I521565);
nor I_30555 (I521468,I521517,I521949);
not I_30556 (I521980,I521941);
nor I_30557 (I521997,I521980,I521675);
DFFARX1 I_30558 (I521997,I2507,I521491,I521474,);
nand I_30559 (I522028,I521980,I521607);
nor I_30560 (I521462,I521833,I522028);
not I_30561 (I522086,I2514);
DFFARX1 I_30562 (I6096,I2507,I522086,I522112,);
DFFARX1 I_30563 (I522112,I2507,I522086,I522129,);
not I_30564 (I522078,I522129);
DFFARX1 I_30565 (I6087,I2507,I522086,I522160,);
not I_30566 (I522168,I6090);
nor I_30567 (I522185,I522112,I522168);
not I_30568 (I522202,I6102);
not I_30569 (I522219,I6087);
nand I_30570 (I522236,I522219,I6102);
nor I_30571 (I522253,I522168,I522236);
nor I_30572 (I522270,I522160,I522253);
DFFARX1 I_30573 (I522219,I2507,I522086,I522075,);
nor I_30574 (I522301,I6087,I6093);
nand I_30575 (I522318,I522301,I6105);
nor I_30576 (I522335,I522318,I522202);
nand I_30577 (I522060,I522335,I6090);
DFFARX1 I_30578 (I522318,I2507,I522086,I522072,);
nand I_30579 (I522380,I522202,I6087);
nor I_30580 (I522397,I522202,I6087);
nand I_30581 (I522066,I522185,I522397);
not I_30582 (I522428,I6108);
nor I_30583 (I522445,I522428,I522380);
DFFARX1 I_30584 (I522445,I2507,I522086,I522054,);
nor I_30585 (I522476,I522428,I6090);
and I_30586 (I522493,I522476,I6099);
or I_30587 (I522510,I522493,I6093);
DFFARX1 I_30588 (I522510,I2507,I522086,I522536,);
nor I_30589 (I522544,I522536,I522160);
nor I_30590 (I522063,I522112,I522544);
not I_30591 (I522575,I522536);
nor I_30592 (I522592,I522575,I522270);
DFFARX1 I_30593 (I522592,I2507,I522086,I522069,);
nand I_30594 (I522623,I522575,I522202);
nor I_30595 (I522057,I522428,I522623);
not I_30596 (I522681,I2514);
DFFARX1 I_30597 (I116528,I2507,I522681,I522707,);
DFFARX1 I_30598 (I522707,I2507,I522681,I522724,);
not I_30599 (I522673,I522724);
DFFARX1 I_30600 (I116540,I2507,I522681,I522755,);
not I_30601 (I522763,I116531);
nor I_30602 (I522780,I522707,I522763);
not I_30603 (I522797,I116522);
not I_30604 (I522814,I116519);
nand I_30605 (I522831,I522814,I116522);
nor I_30606 (I522848,I522763,I522831);
nor I_30607 (I522865,I522755,I522848);
DFFARX1 I_30608 (I522814,I2507,I522681,I522670,);
nor I_30609 (I522896,I116519,I116519);
nand I_30610 (I522913,I522896,I116537);
nor I_30611 (I522930,I522913,I522797);
nand I_30612 (I522655,I522930,I116531);
DFFARX1 I_30613 (I522913,I2507,I522681,I522667,);
nand I_30614 (I522975,I522797,I116519);
nor I_30615 (I522992,I522797,I116519);
nand I_30616 (I522661,I522780,I522992);
not I_30617 (I523023,I116543);
nor I_30618 (I523040,I523023,I522975);
DFFARX1 I_30619 (I523040,I2507,I522681,I522649,);
nor I_30620 (I523071,I523023,I116522);
and I_30621 (I523088,I523071,I116525);
or I_30622 (I523105,I523088,I116534);
DFFARX1 I_30623 (I523105,I2507,I522681,I523131,);
nor I_30624 (I523139,I523131,I522755);
nor I_30625 (I522658,I522707,I523139);
not I_30626 (I523170,I523131);
nor I_30627 (I523187,I523170,I522865);
DFFARX1 I_30628 (I523187,I2507,I522681,I522664,);
nand I_30629 (I523218,I523170,I522797);
nor I_30630 (I522652,I523023,I523218);
not I_30631 (I523276,I2514);
DFFARX1 I_30632 (I714537,I2507,I523276,I523302,);
DFFARX1 I_30633 (I523302,I2507,I523276,I523319,);
not I_30634 (I523268,I523319);
DFFARX1 I_30635 (I714531,I2507,I523276,I523350,);
not I_30636 (I523358,I714528);
nor I_30637 (I523375,I523302,I523358);
not I_30638 (I523392,I714540);
not I_30639 (I523409,I714543);
nand I_30640 (I523426,I523409,I714540);
nor I_30641 (I523443,I523358,I523426);
nor I_30642 (I523460,I523350,I523443);
DFFARX1 I_30643 (I523409,I2507,I523276,I523265,);
nor I_30644 (I523491,I714543,I714552);
nand I_30645 (I523508,I523491,I714546);
nor I_30646 (I523525,I523508,I523392);
nand I_30647 (I523250,I523525,I714528);
DFFARX1 I_30648 (I523508,I2507,I523276,I523262,);
nand I_30649 (I523570,I523392,I714543);
nor I_30650 (I523587,I523392,I714543);
nand I_30651 (I523256,I523375,I523587);
not I_30652 (I523618,I714534);
nor I_30653 (I523635,I523618,I523570);
DFFARX1 I_30654 (I523635,I2507,I523276,I523244,);
nor I_30655 (I523666,I523618,I714549);
and I_30656 (I523683,I523666,I714528);
or I_30657 (I523700,I523683,I714531);
DFFARX1 I_30658 (I523700,I2507,I523276,I523726,);
nor I_30659 (I523734,I523726,I523350);
nor I_30660 (I523253,I523302,I523734);
not I_30661 (I523765,I523726);
nor I_30662 (I523782,I523765,I523460);
DFFARX1 I_30663 (I523782,I2507,I523276,I523259,);
nand I_30664 (I523813,I523765,I523392);
nor I_30665 (I523247,I523618,I523813);
not I_30666 (I523871,I2514);
DFFARX1 I_30667 (I547489,I2507,I523871,I523897,);
DFFARX1 I_30668 (I523897,I2507,I523871,I523914,);
not I_30669 (I523863,I523914);
DFFARX1 I_30670 (I547501,I2507,I523871,I523945,);
not I_30671 (I523953,I547486);
nor I_30672 (I523970,I523897,I523953);
not I_30673 (I523987,I547504);
not I_30674 (I524004,I547495);
nand I_30675 (I524021,I524004,I547504);
nor I_30676 (I524038,I523953,I524021);
nor I_30677 (I524055,I523945,I524038);
DFFARX1 I_30678 (I524004,I2507,I523871,I523860,);
nor I_30679 (I524086,I547495,I547507);
nand I_30680 (I524103,I524086,I547510);
nor I_30681 (I524120,I524103,I523987);
nand I_30682 (I523845,I524120,I547486);
DFFARX1 I_30683 (I524103,I2507,I523871,I523857,);
nand I_30684 (I524165,I523987,I547495);
nor I_30685 (I524182,I523987,I547495);
nand I_30686 (I523851,I523970,I524182);
not I_30687 (I524213,I547486);
nor I_30688 (I524230,I524213,I524165);
DFFARX1 I_30689 (I524230,I2507,I523871,I523839,);
nor I_30690 (I524261,I524213,I547498);
and I_30691 (I524278,I524261,I547492);
or I_30692 (I524295,I524278,I547489);
DFFARX1 I_30693 (I524295,I2507,I523871,I524321,);
nor I_30694 (I524329,I524321,I523945);
nor I_30695 (I523848,I523897,I524329);
not I_30696 (I524360,I524321);
nor I_30697 (I524377,I524360,I524055);
DFFARX1 I_30698 (I524377,I2507,I523871,I523854,);
nand I_30699 (I524408,I524360,I523987);
nor I_30700 (I523842,I524213,I524408);
not I_30701 (I524466,I2514);
DFFARX1 I_30702 (I67517,I2507,I524466,I524492,);
DFFARX1 I_30703 (I524492,I2507,I524466,I524509,);
not I_30704 (I524458,I524509);
DFFARX1 I_30705 (I67529,I2507,I524466,I524540,);
not I_30706 (I524548,I67520);
nor I_30707 (I524565,I524492,I524548);
not I_30708 (I524582,I67511);
not I_30709 (I524599,I67508);
nand I_30710 (I524616,I524599,I67511);
nor I_30711 (I524633,I524548,I524616);
nor I_30712 (I524650,I524540,I524633);
DFFARX1 I_30713 (I524599,I2507,I524466,I524455,);
nor I_30714 (I524681,I67508,I67508);
nand I_30715 (I524698,I524681,I67526);
nor I_30716 (I524715,I524698,I524582);
nand I_30717 (I524440,I524715,I67520);
DFFARX1 I_30718 (I524698,I2507,I524466,I524452,);
nand I_30719 (I524760,I524582,I67508);
nor I_30720 (I524777,I524582,I67508);
nand I_30721 (I524446,I524565,I524777);
not I_30722 (I524808,I67532);
nor I_30723 (I524825,I524808,I524760);
DFFARX1 I_30724 (I524825,I2507,I524466,I524434,);
nor I_30725 (I524856,I524808,I67511);
and I_30726 (I524873,I524856,I67514);
or I_30727 (I524890,I524873,I67523);
DFFARX1 I_30728 (I524890,I2507,I524466,I524916,);
nor I_30729 (I524924,I524916,I524540);
nor I_30730 (I524443,I524492,I524924);
not I_30731 (I524955,I524916);
nor I_30732 (I524972,I524955,I524650);
DFFARX1 I_30733 (I524972,I2507,I524466,I524449,);
nand I_30734 (I525003,I524955,I524582);
nor I_30735 (I524437,I524808,I525003);
not I_30736 (I525061,I2514);
DFFARX1 I_30737 (I678701,I2507,I525061,I525087,);
DFFARX1 I_30738 (I525087,I2507,I525061,I525104,);
not I_30739 (I525053,I525104);
DFFARX1 I_30740 (I678695,I2507,I525061,I525135,);
not I_30741 (I525143,I678692);
nor I_30742 (I525160,I525087,I525143);
not I_30743 (I525177,I678704);
not I_30744 (I525194,I678707);
nand I_30745 (I525211,I525194,I678704);
nor I_30746 (I525228,I525143,I525211);
nor I_30747 (I525245,I525135,I525228);
DFFARX1 I_30748 (I525194,I2507,I525061,I525050,);
nor I_30749 (I525276,I678707,I678716);
nand I_30750 (I525293,I525276,I678710);
nor I_30751 (I525310,I525293,I525177);
nand I_30752 (I525035,I525310,I678692);
DFFARX1 I_30753 (I525293,I2507,I525061,I525047,);
nand I_30754 (I525355,I525177,I678707);
nor I_30755 (I525372,I525177,I678707);
nand I_30756 (I525041,I525160,I525372);
not I_30757 (I525403,I678698);
nor I_30758 (I525420,I525403,I525355);
DFFARX1 I_30759 (I525420,I2507,I525061,I525029,);
nor I_30760 (I525451,I525403,I678713);
and I_30761 (I525468,I525451,I678692);
or I_30762 (I525485,I525468,I678695);
DFFARX1 I_30763 (I525485,I2507,I525061,I525511,);
nor I_30764 (I525519,I525511,I525135);
nor I_30765 (I525038,I525087,I525519);
not I_30766 (I525550,I525511);
nor I_30767 (I525567,I525550,I525245);
DFFARX1 I_30768 (I525567,I2507,I525061,I525044,);
nand I_30769 (I525598,I525550,I525177);
nor I_30770 (I525032,I525403,I525598);
not I_30771 (I525656,I2514);
DFFARX1 I_30772 (I1048850,I2507,I525656,I525682,);
DFFARX1 I_30773 (I525682,I2507,I525656,I525699,);
not I_30774 (I525648,I525699);
DFFARX1 I_30775 (I1048853,I2507,I525656,I525730,);
not I_30776 (I525738,I1048856);
nor I_30777 (I525755,I525682,I525738);
not I_30778 (I525772,I1048868);
not I_30779 (I525789,I1048859);
nand I_30780 (I525806,I525789,I1048868);
nor I_30781 (I525823,I525738,I525806);
nor I_30782 (I525840,I525730,I525823);
DFFARX1 I_30783 (I525789,I2507,I525656,I525645,);
nor I_30784 (I525871,I1048859,I1048865);
nand I_30785 (I525888,I525871,I1048853);
nor I_30786 (I525905,I525888,I525772);
nand I_30787 (I525630,I525905,I1048856);
DFFARX1 I_30788 (I525888,I2507,I525656,I525642,);
nand I_30789 (I525950,I525772,I1048859);
nor I_30790 (I525967,I525772,I1048859);
nand I_30791 (I525636,I525755,I525967);
not I_30792 (I525998,I1048856);
nor I_30793 (I526015,I525998,I525950);
DFFARX1 I_30794 (I526015,I2507,I525656,I525624,);
nor I_30795 (I526046,I525998,I1048862);
and I_30796 (I526063,I526046,I1048850);
or I_30797 (I526080,I526063,I1048871);
DFFARX1 I_30798 (I526080,I2507,I525656,I526106,);
nor I_30799 (I526114,I526106,I525730);
nor I_30800 (I525633,I525682,I526114);
not I_30801 (I526145,I526106);
nor I_30802 (I526162,I526145,I525840);
DFFARX1 I_30803 (I526162,I2507,I525656,I525639,);
nand I_30804 (I526193,I526145,I525772);
nor I_30805 (I525627,I525998,I526193);
not I_30806 (I526251,I2514);
DFFARX1 I_30807 (I201400,I2507,I526251,I526277,);
DFFARX1 I_30808 (I526277,I2507,I526251,I526294,);
not I_30809 (I526243,I526294);
DFFARX1 I_30810 (I201424,I2507,I526251,I526325,);
not I_30811 (I526333,I201418);
nor I_30812 (I526350,I526277,I526333);
not I_30813 (I526367,I201412);
not I_30814 (I526384,I201409);
nand I_30815 (I526401,I526384,I201412);
nor I_30816 (I526418,I526333,I526401);
nor I_30817 (I526435,I526325,I526418);
DFFARX1 I_30818 (I526384,I2507,I526251,I526240,);
nor I_30819 (I526466,I201409,I201403);
nand I_30820 (I526483,I526466,I201421);
nor I_30821 (I526500,I526483,I526367);
nand I_30822 (I526225,I526500,I201418);
DFFARX1 I_30823 (I526483,I2507,I526251,I526237,);
nand I_30824 (I526545,I526367,I201409);
nor I_30825 (I526562,I526367,I201409);
nand I_30826 (I526231,I526350,I526562);
not I_30827 (I526593,I201415);
nor I_30828 (I526610,I526593,I526545);
DFFARX1 I_30829 (I526610,I2507,I526251,I526219,);
nor I_30830 (I526641,I526593,I201400);
and I_30831 (I526658,I526641,I201406);
or I_30832 (I526675,I526658,I201403);
DFFARX1 I_30833 (I526675,I2507,I526251,I526701,);
nor I_30834 (I526709,I526701,I526325);
nor I_30835 (I526228,I526277,I526709);
not I_30836 (I526740,I526701);
nor I_30837 (I526757,I526740,I526435);
DFFARX1 I_30838 (I526757,I2507,I526251,I526234,);
nand I_30839 (I526788,I526740,I526367);
nor I_30840 (I526222,I526593,I526788);
not I_30841 (I526846,I2514);
DFFARX1 I_30842 (I350862,I2507,I526846,I526872,);
DFFARX1 I_30843 (I526872,I2507,I526846,I526889,);
not I_30844 (I526838,I526889);
DFFARX1 I_30845 (I350850,I2507,I526846,I526920,);
not I_30846 (I526928,I350853);
nor I_30847 (I526945,I526872,I526928);
not I_30848 (I526962,I350856);
not I_30849 (I526979,I350868);
nand I_30850 (I526996,I526979,I350856);
nor I_30851 (I527013,I526928,I526996);
nor I_30852 (I527030,I526920,I527013);
DFFARX1 I_30853 (I526979,I2507,I526846,I526835,);
nor I_30854 (I527061,I350868,I350859);
nand I_30855 (I527078,I527061,I350847);
nor I_30856 (I527095,I527078,I526962);
nand I_30857 (I526820,I527095,I350853);
DFFARX1 I_30858 (I527078,I2507,I526846,I526832,);
nand I_30859 (I527140,I526962,I350868);
nor I_30860 (I527157,I526962,I350868);
nand I_30861 (I526826,I526945,I527157);
not I_30862 (I527188,I350865);
nor I_30863 (I527205,I527188,I527140);
DFFARX1 I_30864 (I527205,I2507,I526846,I526814,);
nor I_30865 (I527236,I527188,I350871);
and I_30866 (I527253,I527236,I350874);
or I_30867 (I527270,I527253,I350847);
DFFARX1 I_30868 (I527270,I2507,I526846,I527296,);
nor I_30869 (I527304,I527296,I526920);
nor I_30870 (I526823,I526872,I527304);
not I_30871 (I527335,I527296);
nor I_30872 (I527352,I527335,I527030);
DFFARX1 I_30873 (I527352,I2507,I526846,I526829,);
nand I_30874 (I527383,I527335,I526962);
nor I_30875 (I526817,I527188,I527383);
not I_30876 (I527441,I2514);
DFFARX1 I_30877 (I327674,I2507,I527441,I527467,);
DFFARX1 I_30878 (I527467,I2507,I527441,I527484,);
not I_30879 (I527433,I527484);
DFFARX1 I_30880 (I327662,I2507,I527441,I527515,);
not I_30881 (I527523,I327665);
nor I_30882 (I527540,I527467,I527523);
not I_30883 (I527557,I327668);
not I_30884 (I527574,I327680);
nand I_30885 (I527591,I527574,I327668);
nor I_30886 (I527608,I527523,I527591);
nor I_30887 (I527625,I527515,I527608);
DFFARX1 I_30888 (I527574,I2507,I527441,I527430,);
nor I_30889 (I527656,I327680,I327671);
nand I_30890 (I527673,I527656,I327659);
nor I_30891 (I527690,I527673,I527557);
nand I_30892 (I527415,I527690,I327665);
DFFARX1 I_30893 (I527673,I2507,I527441,I527427,);
nand I_30894 (I527735,I527557,I327680);
nor I_30895 (I527752,I527557,I327680);
nand I_30896 (I527421,I527540,I527752);
not I_30897 (I527783,I327677);
nor I_30898 (I527800,I527783,I527735);
DFFARX1 I_30899 (I527800,I2507,I527441,I527409,);
nor I_30900 (I527831,I527783,I327683);
and I_30901 (I527848,I527831,I327686);
or I_30902 (I527865,I527848,I327659);
DFFARX1 I_30903 (I527865,I2507,I527441,I527891,);
nor I_30904 (I527899,I527891,I527515);
nor I_30905 (I527418,I527467,I527899);
not I_30906 (I527930,I527891);
nor I_30907 (I527947,I527930,I527625);
DFFARX1 I_30908 (I527947,I2507,I527441,I527424,);
nand I_30909 (I527978,I527930,I527557);
nor I_30910 (I527412,I527783,I527978);
not I_30911 (I528036,I2514);
DFFARX1 I_30912 (I1019117,I2507,I528036,I528062,);
DFFARX1 I_30913 (I528062,I2507,I528036,I528079,);
not I_30914 (I528028,I528079);
DFFARX1 I_30915 (I1019120,I2507,I528036,I528110,);
not I_30916 (I528118,I1019123);
nor I_30917 (I528135,I528062,I528118);
not I_30918 (I528152,I1019135);
not I_30919 (I528169,I1019126);
nand I_30920 (I528186,I528169,I1019135);
nor I_30921 (I528203,I528118,I528186);
nor I_30922 (I528220,I528110,I528203);
DFFARX1 I_30923 (I528169,I2507,I528036,I528025,);
nor I_30924 (I528251,I1019126,I1019132);
nand I_30925 (I528268,I528251,I1019120);
nor I_30926 (I528285,I528268,I528152);
nand I_30927 (I528010,I528285,I1019123);
DFFARX1 I_30928 (I528268,I2507,I528036,I528022,);
nand I_30929 (I528330,I528152,I1019126);
nor I_30930 (I528347,I528152,I1019126);
nand I_30931 (I528016,I528135,I528347);
not I_30932 (I528378,I1019123);
nor I_30933 (I528395,I528378,I528330);
DFFARX1 I_30934 (I528395,I2507,I528036,I528004,);
nor I_30935 (I528426,I528378,I1019129);
and I_30936 (I528443,I528426,I1019117);
or I_30937 (I528460,I528443,I1019138);
DFFARX1 I_30938 (I528460,I2507,I528036,I528486,);
nor I_30939 (I528494,I528486,I528110);
nor I_30940 (I528013,I528062,I528494);
not I_30941 (I528525,I528486);
nor I_30942 (I528542,I528525,I528220);
DFFARX1 I_30943 (I528542,I2507,I528036,I528019,);
nand I_30944 (I528573,I528525,I528152);
nor I_30945 (I528007,I528378,I528573);
not I_30946 (I528631,I2514);
DFFARX1 I_30947 (I1948,I2507,I528631,I528657,);
DFFARX1 I_30948 (I528657,I2507,I528631,I528674,);
not I_30949 (I528623,I528674);
DFFARX1 I_30950 (I1532,I2507,I528631,I528705,);
not I_30951 (I528713,I2196);
nor I_30952 (I528730,I528657,I528713);
not I_30953 (I528747,I2060);
not I_30954 (I528764,I2276);
nand I_30955 (I528781,I528764,I2060);
nor I_30956 (I528798,I528713,I528781);
nor I_30957 (I528815,I528705,I528798);
DFFARX1 I_30958 (I528764,I2507,I528631,I528620,);
nor I_30959 (I528846,I2276,I1460);
nand I_30960 (I528863,I528846,I1508);
nor I_30961 (I528880,I528863,I528747);
nand I_30962 (I528605,I528880,I2196);
DFFARX1 I_30963 (I528863,I2507,I528631,I528617,);
nand I_30964 (I528925,I528747,I2276);
nor I_30965 (I528942,I528747,I2276);
nand I_30966 (I528611,I528730,I528942);
not I_30967 (I528973,I2444);
nor I_30968 (I528990,I528973,I528925);
DFFARX1 I_30969 (I528990,I2507,I528631,I528599,);
nor I_30970 (I529021,I528973,I2076);
and I_30971 (I529038,I529021,I2364);
or I_30972 (I529055,I529038,I2172);
DFFARX1 I_30973 (I529055,I2507,I528631,I529081,);
nor I_30974 (I529089,I529081,I528705);
nor I_30975 (I528608,I528657,I529089);
not I_30976 (I529120,I529081);
nor I_30977 (I529137,I529120,I528815);
DFFARX1 I_30978 (I529137,I2507,I528631,I528614,);
nand I_30979 (I529168,I529120,I528747);
nor I_30980 (I528602,I528973,I529168);
not I_30981 (I529226,I2514);
DFFARX1 I_30982 (I1235714,I2507,I529226,I529252,);
DFFARX1 I_30983 (I529252,I2507,I529226,I529269,);
not I_30984 (I529218,I529269);
DFFARX1 I_30985 (I1235729,I2507,I529226,I529300,);
not I_30986 (I529308,I1235738);
nor I_30987 (I529325,I529252,I529308);
not I_30988 (I529342,I1235717);
not I_30989 (I529359,I1235723);
nand I_30990 (I529376,I529359,I1235717);
nor I_30991 (I529393,I529308,I529376);
nor I_30992 (I529410,I529300,I529393);
DFFARX1 I_30993 (I529359,I2507,I529226,I529215,);
nor I_30994 (I529441,I1235723,I1235735);
nand I_30995 (I529458,I529441,I1235732);
nor I_30996 (I529475,I529458,I529342);
nand I_30997 (I529200,I529475,I1235738);
DFFARX1 I_30998 (I529458,I2507,I529226,I529212,);
nand I_30999 (I529520,I529342,I1235723);
nor I_31000 (I529537,I529342,I1235723);
nand I_31001 (I529206,I529325,I529537);
not I_31002 (I529568,I1235714);
nor I_31003 (I529585,I529568,I529520);
DFFARX1 I_31004 (I529585,I2507,I529226,I529194,);
nor I_31005 (I529616,I529568,I1235726);
and I_31006 (I529633,I529616,I1235720);
or I_31007 (I529650,I529633,I1235717);
DFFARX1 I_31008 (I529650,I2507,I529226,I529676,);
nor I_31009 (I529684,I529676,I529300);
nor I_31010 (I529203,I529252,I529684);
not I_31011 (I529715,I529676);
nor I_31012 (I529732,I529715,I529410);
DFFARX1 I_31013 (I529732,I2507,I529226,I529209,);
nand I_31014 (I529763,I529715,I529342);
nor I_31015 (I529197,I529568,I529763);
not I_31016 (I529821,I2514);
DFFARX1 I_31017 (I26929,I2507,I529821,I529847,);
DFFARX1 I_31018 (I529847,I2507,I529821,I529864,);
not I_31019 (I529813,I529864);
DFFARX1 I_31020 (I26929,I2507,I529821,I529895,);
not I_31021 (I529903,I26944);
nor I_31022 (I529920,I529847,I529903);
not I_31023 (I529937,I26947);
not I_31024 (I529954,I26938);
nand I_31025 (I529971,I529954,I26947);
nor I_31026 (I529988,I529903,I529971);
nor I_31027 (I530005,I529895,I529988);
DFFARX1 I_31028 (I529954,I2507,I529821,I529810,);
nor I_31029 (I530036,I26938,I26950);
nand I_31030 (I530053,I530036,I26932);
nor I_31031 (I530070,I530053,I529937);
nand I_31032 (I529795,I530070,I26944);
DFFARX1 I_31033 (I530053,I2507,I529821,I529807,);
nand I_31034 (I530115,I529937,I26938);
nor I_31035 (I530132,I529937,I26938);
nand I_31036 (I529801,I529920,I530132);
not I_31037 (I530163,I26932);
nor I_31038 (I530180,I530163,I530115);
DFFARX1 I_31039 (I530180,I2507,I529821,I529789,);
nor I_31040 (I530211,I530163,I26941);
and I_31041 (I530228,I530211,I26935);
or I_31042 (I530245,I530228,I26953);
DFFARX1 I_31043 (I530245,I2507,I529821,I530271,);
nor I_31044 (I530279,I530271,I529895);
nor I_31045 (I529798,I529847,I530279);
not I_31046 (I530310,I530271);
nor I_31047 (I530327,I530310,I530005);
DFFARX1 I_31048 (I530327,I2507,I529821,I529804,);
nand I_31049 (I530358,I530310,I529937);
nor I_31050 (I529792,I530163,I530358);
not I_31051 (I530416,I2514);
DFFARX1 I_31052 (I1176878,I2507,I530416,I530442,);
DFFARX1 I_31053 (I530442,I2507,I530416,I530459,);
not I_31054 (I530408,I530459);
DFFARX1 I_31055 (I1176860,I2507,I530416,I530490,);
not I_31056 (I530498,I1176866);
nor I_31057 (I530515,I530442,I530498);
not I_31058 (I530532,I1176881);
not I_31059 (I530549,I1176872);
nand I_31060 (I530566,I530549,I1176881);
nor I_31061 (I530583,I530498,I530566);
nor I_31062 (I530600,I530490,I530583);
DFFARX1 I_31063 (I530549,I2507,I530416,I530405,);
nor I_31064 (I530631,I1176872,I1176884);
nand I_31065 (I530648,I530631,I1176863);
nor I_31066 (I530665,I530648,I530532);
nand I_31067 (I530390,I530665,I1176866);
DFFARX1 I_31068 (I530648,I2507,I530416,I530402,);
nand I_31069 (I530710,I530532,I1176872);
nor I_31070 (I530727,I530532,I1176872);
nand I_31071 (I530396,I530515,I530727);
not I_31072 (I530758,I1176869);
nor I_31073 (I530775,I530758,I530710);
DFFARX1 I_31074 (I530775,I2507,I530416,I530384,);
nor I_31075 (I530806,I530758,I1176875);
and I_31076 (I530823,I530806,I1176860);
or I_31077 (I530840,I530823,I1176863);
DFFARX1 I_31078 (I530840,I2507,I530416,I530866,);
nor I_31079 (I530874,I530866,I530490);
nor I_31080 (I530393,I530442,I530874);
not I_31081 (I530905,I530866);
nor I_31082 (I530922,I530905,I530600);
DFFARX1 I_31083 (I530922,I2507,I530416,I530399,);
nand I_31084 (I530953,I530905,I530532);
nor I_31085 (I530387,I530758,I530953);
not I_31086 (I531011,I2514);
DFFARX1 I_31087 (I1057265,I2507,I531011,I531037,);
DFFARX1 I_31088 (I531037,I2507,I531011,I531054,);
not I_31089 (I531003,I531054);
DFFARX1 I_31090 (I1057268,I2507,I531011,I531085,);
not I_31091 (I531093,I1057271);
nor I_31092 (I531110,I531037,I531093);
not I_31093 (I531127,I1057283);
not I_31094 (I531144,I1057274);
nand I_31095 (I531161,I531144,I1057283);
nor I_31096 (I531178,I531093,I531161);
nor I_31097 (I531195,I531085,I531178);
DFFARX1 I_31098 (I531144,I2507,I531011,I531000,);
nor I_31099 (I531226,I1057274,I1057280);
nand I_31100 (I531243,I531226,I1057268);
nor I_31101 (I531260,I531243,I531127);
nand I_31102 (I530985,I531260,I1057271);
DFFARX1 I_31103 (I531243,I2507,I531011,I530997,);
nand I_31104 (I531305,I531127,I1057274);
nor I_31105 (I531322,I531127,I1057274);
nand I_31106 (I530991,I531110,I531322);
not I_31107 (I531353,I1057271);
nor I_31108 (I531370,I531353,I531305);
DFFARX1 I_31109 (I531370,I2507,I531011,I530979,);
nor I_31110 (I531401,I531353,I1057277);
and I_31111 (I531418,I531401,I1057265);
or I_31112 (I531435,I531418,I1057286);
DFFARX1 I_31113 (I531435,I2507,I531011,I531461,);
nor I_31114 (I531469,I531461,I531085);
nor I_31115 (I530988,I531037,I531469);
not I_31116 (I531500,I531461);
nor I_31117 (I531517,I531500,I531195);
DFFARX1 I_31118 (I531517,I2507,I531011,I530994,);
nand I_31119 (I531548,I531500,I531127);
nor I_31120 (I530982,I531353,I531548);
not I_31121 (I531606,I2514);
DFFARX1 I_31122 (I1047167,I2507,I531606,I531632,);
DFFARX1 I_31123 (I531632,I2507,I531606,I531649,);
not I_31124 (I531598,I531649);
DFFARX1 I_31125 (I1047170,I2507,I531606,I531680,);
not I_31126 (I531688,I1047173);
nor I_31127 (I531705,I531632,I531688);
not I_31128 (I531722,I1047185);
not I_31129 (I531739,I1047176);
nand I_31130 (I531756,I531739,I1047185);
nor I_31131 (I531773,I531688,I531756);
nor I_31132 (I531790,I531680,I531773);
DFFARX1 I_31133 (I531739,I2507,I531606,I531595,);
nor I_31134 (I531821,I1047176,I1047182);
nand I_31135 (I531838,I531821,I1047170);
nor I_31136 (I531855,I531838,I531722);
nand I_31137 (I531580,I531855,I1047173);
DFFARX1 I_31138 (I531838,I2507,I531606,I531592,);
nand I_31139 (I531900,I531722,I1047176);
nor I_31140 (I531917,I531722,I1047176);
nand I_31141 (I531586,I531705,I531917);
not I_31142 (I531948,I1047173);
nor I_31143 (I531965,I531948,I531900);
DFFARX1 I_31144 (I531965,I2507,I531606,I531574,);
nor I_31145 (I531996,I531948,I1047179);
and I_31146 (I532013,I531996,I1047167);
or I_31147 (I532030,I532013,I1047188);
DFFARX1 I_31148 (I532030,I2507,I531606,I532056,);
nor I_31149 (I532064,I532056,I531680);
nor I_31150 (I531583,I531632,I532064);
not I_31151 (I532095,I532056);
nor I_31152 (I532112,I532095,I531790);
DFFARX1 I_31153 (I532112,I2507,I531606,I531589,);
nand I_31154 (I532143,I532095,I531722);
nor I_31155 (I531577,I531948,I532143);
not I_31156 (I532201,I2514);
DFFARX1 I_31157 (I1391587,I2507,I532201,I532227,);
DFFARX1 I_31158 (I532227,I2507,I532201,I532244,);
not I_31159 (I532193,I532244);
DFFARX1 I_31160 (I1391593,I2507,I532201,I532275,);
not I_31161 (I532283,I1391608);
nor I_31162 (I532300,I532227,I532283);
not I_31163 (I532317,I1391599);
not I_31164 (I532334,I1391596);
nand I_31165 (I532351,I532334,I1391599);
nor I_31166 (I532368,I532283,I532351);
nor I_31167 (I532385,I532275,I532368);
DFFARX1 I_31168 (I532334,I2507,I532201,I532190,);
nor I_31169 (I532416,I1391596,I1391587);
nand I_31170 (I532433,I532416,I1391611);
nor I_31171 (I532450,I532433,I532317);
nand I_31172 (I532175,I532450,I1391608);
DFFARX1 I_31173 (I532433,I2507,I532201,I532187,);
nand I_31174 (I532495,I532317,I1391596);
nor I_31175 (I532512,I532317,I1391596);
nand I_31176 (I532181,I532300,I532512);
not I_31177 (I532543,I1391605);
nor I_31178 (I532560,I532543,I532495);
DFFARX1 I_31179 (I532560,I2507,I532201,I532169,);
nor I_31180 (I532591,I532543,I1391590);
and I_31181 (I532608,I532591,I1391602);
or I_31182 (I532625,I532608,I1391614);
DFFARX1 I_31183 (I532625,I2507,I532201,I532651,);
nor I_31184 (I532659,I532651,I532275);
nor I_31185 (I532178,I532227,I532659);
not I_31186 (I532690,I532651);
nor I_31187 (I532707,I532690,I532385);
DFFARX1 I_31188 (I532707,I2507,I532201,I532184,);
nand I_31189 (I532738,I532690,I532317);
nor I_31190 (I532172,I532543,I532738);
not I_31191 (I532796,I2514);
DFFARX1 I_31192 (I361402,I2507,I532796,I532822,);
DFFARX1 I_31193 (I532822,I2507,I532796,I532839,);
not I_31194 (I532788,I532839);
DFFARX1 I_31195 (I361390,I2507,I532796,I532870,);
not I_31196 (I532878,I361393);
nor I_31197 (I532895,I532822,I532878);
not I_31198 (I532912,I361396);
not I_31199 (I532929,I361408);
nand I_31200 (I532946,I532929,I361396);
nor I_31201 (I532963,I532878,I532946);
nor I_31202 (I532980,I532870,I532963);
DFFARX1 I_31203 (I532929,I2507,I532796,I532785,);
nor I_31204 (I533011,I361408,I361399);
nand I_31205 (I533028,I533011,I361387);
nor I_31206 (I533045,I533028,I532912);
nand I_31207 (I532770,I533045,I361393);
DFFARX1 I_31208 (I533028,I2507,I532796,I532782,);
nand I_31209 (I533090,I532912,I361408);
nor I_31210 (I533107,I532912,I361408);
nand I_31211 (I532776,I532895,I533107);
not I_31212 (I533138,I361405);
nor I_31213 (I533155,I533138,I533090);
DFFARX1 I_31214 (I533155,I2507,I532796,I532764,);
nor I_31215 (I533186,I533138,I361411);
and I_31216 (I533203,I533186,I361414);
or I_31217 (I533220,I533203,I361387);
DFFARX1 I_31218 (I533220,I2507,I532796,I533246,);
nor I_31219 (I533254,I533246,I532870);
nor I_31220 (I532773,I532822,I533254);
not I_31221 (I533285,I533246);
nor I_31222 (I533302,I533285,I532980);
DFFARX1 I_31223 (I533302,I2507,I532796,I532779,);
nand I_31224 (I533333,I533285,I532912);
nor I_31225 (I532767,I533138,I533333);
not I_31226 (I533391,I2514);
DFFARX1 I_31227 (I22713,I2507,I533391,I533417,);
DFFARX1 I_31228 (I533417,I2507,I533391,I533434,);
not I_31229 (I533383,I533434);
DFFARX1 I_31230 (I22713,I2507,I533391,I533465,);
not I_31231 (I533473,I22728);
nor I_31232 (I533490,I533417,I533473);
not I_31233 (I533507,I22731);
not I_31234 (I533524,I22722);
nand I_31235 (I533541,I533524,I22731);
nor I_31236 (I533558,I533473,I533541);
nor I_31237 (I533575,I533465,I533558);
DFFARX1 I_31238 (I533524,I2507,I533391,I533380,);
nor I_31239 (I533606,I22722,I22734);
nand I_31240 (I533623,I533606,I22716);
nor I_31241 (I533640,I533623,I533507);
nand I_31242 (I533365,I533640,I22728);
DFFARX1 I_31243 (I533623,I2507,I533391,I533377,);
nand I_31244 (I533685,I533507,I22722);
nor I_31245 (I533702,I533507,I22722);
nand I_31246 (I533371,I533490,I533702);
not I_31247 (I533733,I22716);
nor I_31248 (I533750,I533733,I533685);
DFFARX1 I_31249 (I533750,I2507,I533391,I533359,);
nor I_31250 (I533781,I533733,I22725);
and I_31251 (I533798,I533781,I22719);
or I_31252 (I533815,I533798,I22737);
DFFARX1 I_31253 (I533815,I2507,I533391,I533841,);
nor I_31254 (I533849,I533841,I533465);
nor I_31255 (I533368,I533417,I533849);
not I_31256 (I533880,I533841);
nor I_31257 (I533897,I533880,I533575);
DFFARX1 I_31258 (I533897,I2507,I533391,I533374,);
nand I_31259 (I533928,I533880,I533507);
nor I_31260 (I533362,I533733,I533928);
not I_31261 (I533986,I2514);
DFFARX1 I_31262 (I46955,I2507,I533986,I534012,);
DFFARX1 I_31263 (I534012,I2507,I533986,I534029,);
not I_31264 (I533978,I534029);
DFFARX1 I_31265 (I46955,I2507,I533986,I534060,);
not I_31266 (I534068,I46970);
nor I_31267 (I534085,I534012,I534068);
not I_31268 (I534102,I46973);
not I_31269 (I534119,I46964);
nand I_31270 (I534136,I534119,I46973);
nor I_31271 (I534153,I534068,I534136);
nor I_31272 (I534170,I534060,I534153);
DFFARX1 I_31273 (I534119,I2507,I533986,I533975,);
nor I_31274 (I534201,I46964,I46976);
nand I_31275 (I534218,I534201,I46958);
nor I_31276 (I534235,I534218,I534102);
nand I_31277 (I533960,I534235,I46970);
DFFARX1 I_31278 (I534218,I2507,I533986,I533972,);
nand I_31279 (I534280,I534102,I46964);
nor I_31280 (I534297,I534102,I46964);
nand I_31281 (I533966,I534085,I534297);
not I_31282 (I534328,I46958);
nor I_31283 (I534345,I534328,I534280);
DFFARX1 I_31284 (I534345,I2507,I533986,I533954,);
nor I_31285 (I534376,I534328,I46967);
and I_31286 (I534393,I534376,I46961);
or I_31287 (I534410,I534393,I46979);
DFFARX1 I_31288 (I534410,I2507,I533986,I534436,);
nor I_31289 (I534444,I534436,I534060);
nor I_31290 (I533963,I534012,I534444);
not I_31291 (I534475,I534436);
nor I_31292 (I534492,I534475,I534170);
DFFARX1 I_31293 (I534492,I2507,I533986,I533969,);
nand I_31294 (I534523,I534475,I534102);
nor I_31295 (I533957,I534328,I534523);
not I_31296 (I534581,I2514);
DFFARX1 I_31297 (I620895,I2507,I534581,I534607,);
DFFARX1 I_31298 (I534607,I2507,I534581,I534624,);
not I_31299 (I534573,I534624);
DFFARX1 I_31300 (I620907,I2507,I534581,I534655,);
not I_31301 (I534663,I620892);
nor I_31302 (I534680,I534607,I534663);
not I_31303 (I534697,I620910);
not I_31304 (I534714,I620901);
nand I_31305 (I534731,I534714,I620910);
nor I_31306 (I534748,I534663,I534731);
nor I_31307 (I534765,I534655,I534748);
DFFARX1 I_31308 (I534714,I2507,I534581,I534570,);
nor I_31309 (I534796,I620901,I620913);
nand I_31310 (I534813,I534796,I620916);
nor I_31311 (I534830,I534813,I534697);
nand I_31312 (I534555,I534830,I620892);
DFFARX1 I_31313 (I534813,I2507,I534581,I534567,);
nand I_31314 (I534875,I534697,I620901);
nor I_31315 (I534892,I534697,I620901);
nand I_31316 (I534561,I534680,I534892);
not I_31317 (I534923,I620892);
nor I_31318 (I534940,I534923,I534875);
DFFARX1 I_31319 (I534940,I2507,I534581,I534549,);
nor I_31320 (I534971,I534923,I620904);
and I_31321 (I534988,I534971,I620898);
or I_31322 (I535005,I534988,I620895);
DFFARX1 I_31323 (I535005,I2507,I534581,I535031,);
nor I_31324 (I535039,I535031,I534655);
nor I_31325 (I534558,I534607,I535039);
not I_31326 (I535070,I535031);
nor I_31327 (I535087,I535070,I534765);
DFFARX1 I_31328 (I535087,I2507,I534581,I534564,);
nand I_31329 (I535118,I535070,I534697);
nor I_31330 (I534552,I534923,I535118);
not I_31331 (I535176,I2514);
DFFARX1 I_31332 (I633617,I2507,I535176,I535202,);
DFFARX1 I_31333 (I535202,I2507,I535176,I535219,);
not I_31334 (I535168,I535219);
DFFARX1 I_31335 (I633611,I2507,I535176,I535250,);
not I_31336 (I535258,I633608);
nor I_31337 (I535275,I535202,I535258);
not I_31338 (I535292,I633620);
not I_31339 (I535309,I633623);
nand I_31340 (I535326,I535309,I633620);
nor I_31341 (I535343,I535258,I535326);
nor I_31342 (I535360,I535250,I535343);
DFFARX1 I_31343 (I535309,I2507,I535176,I535165,);
nor I_31344 (I535391,I633623,I633632);
nand I_31345 (I535408,I535391,I633626);
nor I_31346 (I535425,I535408,I535292);
nand I_31347 (I535150,I535425,I633608);
DFFARX1 I_31348 (I535408,I2507,I535176,I535162,);
nand I_31349 (I535470,I535292,I633623);
nor I_31350 (I535487,I535292,I633623);
nand I_31351 (I535156,I535275,I535487);
not I_31352 (I535518,I633614);
nor I_31353 (I535535,I535518,I535470);
DFFARX1 I_31354 (I535535,I2507,I535176,I535144,);
nor I_31355 (I535566,I535518,I633629);
and I_31356 (I535583,I535566,I633608);
or I_31357 (I535600,I535583,I633611);
DFFARX1 I_31358 (I535600,I2507,I535176,I535626,);
nor I_31359 (I535634,I535626,I535250);
nor I_31360 (I535153,I535202,I535634);
not I_31361 (I535665,I535626);
nor I_31362 (I535682,I535665,I535360);
DFFARX1 I_31363 (I535682,I2507,I535176,I535159,);
nand I_31364 (I535713,I535665,I535292);
nor I_31365 (I535147,I535518,I535713);
not I_31366 (I535771,I2514);
DFFARX1 I_31367 (I1016312,I2507,I535771,I535797,);
DFFARX1 I_31368 (I535797,I2507,I535771,I535814,);
not I_31369 (I535763,I535814);
DFFARX1 I_31370 (I1016315,I2507,I535771,I535845,);
not I_31371 (I535853,I1016318);
nor I_31372 (I535870,I535797,I535853);
not I_31373 (I535887,I1016330);
not I_31374 (I535904,I1016321);
nand I_31375 (I535921,I535904,I1016330);
nor I_31376 (I535938,I535853,I535921);
nor I_31377 (I535955,I535845,I535938);
DFFARX1 I_31378 (I535904,I2507,I535771,I535760,);
nor I_31379 (I535986,I1016321,I1016327);
nand I_31380 (I536003,I535986,I1016315);
nor I_31381 (I536020,I536003,I535887);
nand I_31382 (I535745,I536020,I1016318);
DFFARX1 I_31383 (I536003,I2507,I535771,I535757,);
nand I_31384 (I536065,I535887,I1016321);
nor I_31385 (I536082,I535887,I1016321);
nand I_31386 (I535751,I535870,I536082);
not I_31387 (I536113,I1016318);
nor I_31388 (I536130,I536113,I536065);
DFFARX1 I_31389 (I536130,I2507,I535771,I535739,);
nor I_31390 (I536161,I536113,I1016324);
and I_31391 (I536178,I536161,I1016312);
or I_31392 (I536195,I536178,I1016333);
DFFARX1 I_31393 (I536195,I2507,I535771,I536221,);
nor I_31394 (I536229,I536221,I535845);
nor I_31395 (I535748,I535797,I536229);
not I_31396 (I536260,I536221);
nor I_31397 (I536277,I536260,I535955);
DFFARX1 I_31398 (I536277,I2507,I535771,I535754,);
nand I_31399 (I536308,I536260,I535887);
nor I_31400 (I535742,I536113,I536308);
not I_31401 (I536366,I2514);
DFFARX1 I_31402 (I359821,I2507,I536366,I536392,);
DFFARX1 I_31403 (I536392,I2507,I536366,I536409,);
not I_31404 (I536358,I536409);
DFFARX1 I_31405 (I359809,I2507,I536366,I536440,);
not I_31406 (I536448,I359812);
nor I_31407 (I536465,I536392,I536448);
not I_31408 (I536482,I359815);
not I_31409 (I536499,I359827);
nand I_31410 (I536516,I536499,I359815);
nor I_31411 (I536533,I536448,I536516);
nor I_31412 (I536550,I536440,I536533);
DFFARX1 I_31413 (I536499,I2507,I536366,I536355,);
nor I_31414 (I536581,I359827,I359818);
nand I_31415 (I536598,I536581,I359806);
nor I_31416 (I536615,I536598,I536482);
nand I_31417 (I536340,I536615,I359812);
DFFARX1 I_31418 (I536598,I2507,I536366,I536352,);
nand I_31419 (I536660,I536482,I359827);
nor I_31420 (I536677,I536482,I359827);
nand I_31421 (I536346,I536465,I536677);
not I_31422 (I536708,I359824);
nor I_31423 (I536725,I536708,I536660);
DFFARX1 I_31424 (I536725,I2507,I536366,I536334,);
nor I_31425 (I536756,I536708,I359830);
and I_31426 (I536773,I536756,I359833);
or I_31427 (I536790,I536773,I359806);
DFFARX1 I_31428 (I536790,I2507,I536366,I536816,);
nor I_31429 (I536824,I536816,I536440);
nor I_31430 (I536343,I536392,I536824);
not I_31431 (I536855,I536816);
nor I_31432 (I536872,I536855,I536550);
DFFARX1 I_31433 (I536872,I2507,I536366,I536349,);
nand I_31434 (I536903,I536855,I536482);
nor I_31435 (I536337,I536708,I536903);
not I_31436 (I536961,I2514);
DFFARX1 I_31437 (I1019678,I2507,I536961,I536987,);
DFFARX1 I_31438 (I536987,I2507,I536961,I537004,);
not I_31439 (I536953,I537004);
DFFARX1 I_31440 (I1019681,I2507,I536961,I537035,);
not I_31441 (I537043,I1019684);
nor I_31442 (I537060,I536987,I537043);
not I_31443 (I537077,I1019696);
not I_31444 (I537094,I1019687);
nand I_31445 (I537111,I537094,I1019696);
nor I_31446 (I537128,I537043,I537111);
nor I_31447 (I537145,I537035,I537128);
DFFARX1 I_31448 (I537094,I2507,I536961,I536950,);
nor I_31449 (I537176,I1019687,I1019693);
nand I_31450 (I537193,I537176,I1019681);
nor I_31451 (I537210,I537193,I537077);
nand I_31452 (I536935,I537210,I1019684);
DFFARX1 I_31453 (I537193,I2507,I536961,I536947,);
nand I_31454 (I537255,I537077,I1019687);
nor I_31455 (I537272,I537077,I1019687);
nand I_31456 (I536941,I537060,I537272);
not I_31457 (I537303,I1019684);
nor I_31458 (I537320,I537303,I537255);
DFFARX1 I_31459 (I537320,I2507,I536961,I536929,);
nor I_31460 (I537351,I537303,I1019690);
and I_31461 (I537368,I537351,I1019678);
or I_31462 (I537385,I537368,I1019699);
DFFARX1 I_31463 (I537385,I2507,I536961,I537411,);
nor I_31464 (I537419,I537411,I537035);
nor I_31465 (I536938,I536987,I537419);
not I_31466 (I537450,I537411);
nor I_31467 (I537467,I537450,I537145);
DFFARX1 I_31468 (I537467,I2507,I536961,I536944,);
nand I_31469 (I537498,I537450,I537077);
nor I_31470 (I536932,I537303,I537498);
not I_31471 (I537556,I2514);
DFFARX1 I_31472 (I309756,I2507,I537556,I537582,);
DFFARX1 I_31473 (I537582,I2507,I537556,I537599,);
not I_31474 (I537548,I537599);
DFFARX1 I_31475 (I309744,I2507,I537556,I537630,);
not I_31476 (I537638,I309747);
nor I_31477 (I537655,I537582,I537638);
not I_31478 (I537672,I309750);
not I_31479 (I537689,I309762);
nand I_31480 (I537706,I537689,I309750);
nor I_31481 (I537723,I537638,I537706);
nor I_31482 (I537740,I537630,I537723);
DFFARX1 I_31483 (I537689,I2507,I537556,I537545,);
nor I_31484 (I537771,I309762,I309753);
nand I_31485 (I537788,I537771,I309741);
nor I_31486 (I537805,I537788,I537672);
nand I_31487 (I537530,I537805,I309747);
DFFARX1 I_31488 (I537788,I2507,I537556,I537542,);
nand I_31489 (I537850,I537672,I309762);
nor I_31490 (I537867,I537672,I309762);
nand I_31491 (I537536,I537655,I537867);
not I_31492 (I537898,I309759);
nor I_31493 (I537915,I537898,I537850);
DFFARX1 I_31494 (I537915,I2507,I537556,I537524,);
nor I_31495 (I537946,I537898,I309765);
and I_31496 (I537963,I537946,I309768);
or I_31497 (I537980,I537963,I309741);
DFFARX1 I_31498 (I537980,I2507,I537556,I538006,);
nor I_31499 (I538014,I538006,I537630);
nor I_31500 (I537533,I537582,I538014);
not I_31501 (I538045,I538006);
nor I_31502 (I538062,I538045,I537740);
DFFARX1 I_31503 (I538062,I2507,I537556,I537539,);
nand I_31504 (I538093,I538045,I537672);
nor I_31505 (I537527,I537898,I538093);
not I_31506 (I538151,I2514);
DFFARX1 I_31507 (I1115032,I2507,I538151,I538177,);
DFFARX1 I_31508 (I538177,I2507,I538151,I538194,);
not I_31509 (I538143,I538194);
DFFARX1 I_31510 (I1115014,I2507,I538151,I538225,);
not I_31511 (I538233,I1115020);
nor I_31512 (I538250,I538177,I538233);
not I_31513 (I538267,I1115035);
not I_31514 (I538284,I1115026);
nand I_31515 (I538301,I538284,I1115035);
nor I_31516 (I538318,I538233,I538301);
nor I_31517 (I538335,I538225,I538318);
DFFARX1 I_31518 (I538284,I2507,I538151,I538140,);
nor I_31519 (I538366,I1115026,I1115038);
nand I_31520 (I538383,I538366,I1115017);
nor I_31521 (I538400,I538383,I538267);
nand I_31522 (I538125,I538400,I1115020);
DFFARX1 I_31523 (I538383,I2507,I538151,I538137,);
nand I_31524 (I538445,I538267,I1115026);
nor I_31525 (I538462,I538267,I1115026);
nand I_31526 (I538131,I538250,I538462);
not I_31527 (I538493,I1115023);
nor I_31528 (I538510,I538493,I538445);
DFFARX1 I_31529 (I538510,I2507,I538151,I538119,);
nor I_31530 (I538541,I538493,I1115029);
and I_31531 (I538558,I538541,I1115014);
or I_31532 (I538575,I538558,I1115017);
DFFARX1 I_31533 (I538575,I2507,I538151,I538601,);
nor I_31534 (I538609,I538601,I538225);
nor I_31535 (I538128,I538177,I538609);
not I_31536 (I538640,I538601);
nor I_31537 (I538657,I538640,I538335);
DFFARX1 I_31538 (I538657,I2507,I538151,I538134,);
nand I_31539 (I538688,I538640,I538267);
nor I_31540 (I538122,I538493,I538688);
not I_31541 (I538746,I2514);
DFFARX1 I_31542 (I371942,I2507,I538746,I538772,);
DFFARX1 I_31543 (I538772,I2507,I538746,I538789,);
not I_31544 (I538738,I538789);
DFFARX1 I_31545 (I371930,I2507,I538746,I538820,);
not I_31546 (I538828,I371933);
nor I_31547 (I538845,I538772,I538828);
not I_31548 (I538862,I371936);
not I_31549 (I538879,I371948);
nand I_31550 (I538896,I538879,I371936);
nor I_31551 (I538913,I538828,I538896);
nor I_31552 (I538930,I538820,I538913);
DFFARX1 I_31553 (I538879,I2507,I538746,I538735,);
nor I_31554 (I538961,I371948,I371939);
nand I_31555 (I538978,I538961,I371927);
nor I_31556 (I538995,I538978,I538862);
nand I_31557 (I538720,I538995,I371933);
DFFARX1 I_31558 (I538978,I2507,I538746,I538732,);
nand I_31559 (I539040,I538862,I371948);
nor I_31560 (I539057,I538862,I371948);
nand I_31561 (I538726,I538845,I539057);
not I_31562 (I539088,I371945);
nor I_31563 (I539105,I539088,I539040);
DFFARX1 I_31564 (I539105,I2507,I538746,I538714,);
nor I_31565 (I539136,I539088,I371951);
and I_31566 (I539153,I539136,I371954);
or I_31567 (I539170,I539153,I371927);
DFFARX1 I_31568 (I539170,I2507,I538746,I539196,);
nor I_31569 (I539204,I539196,I538820);
nor I_31570 (I538723,I538772,I539204);
not I_31571 (I539235,I539196);
nor I_31572 (I539252,I539235,I538930);
DFFARX1 I_31573 (I539252,I2507,I538746,I538729,);
nand I_31574 (I539283,I539235,I538862);
nor I_31575 (I538717,I539088,I539283);
not I_31576 (I539341,I2514);
DFFARX1 I_31577 (I1254210,I2507,I539341,I539367,);
DFFARX1 I_31578 (I539367,I2507,I539341,I539384,);
not I_31579 (I539333,I539384);
DFFARX1 I_31580 (I1254225,I2507,I539341,I539415,);
not I_31581 (I539423,I1254234);
nor I_31582 (I539440,I539367,I539423);
not I_31583 (I539457,I1254213);
not I_31584 (I539474,I1254219);
nand I_31585 (I539491,I539474,I1254213);
nor I_31586 (I539508,I539423,I539491);
nor I_31587 (I539525,I539415,I539508);
DFFARX1 I_31588 (I539474,I2507,I539341,I539330,);
nor I_31589 (I539556,I1254219,I1254231);
nand I_31590 (I539573,I539556,I1254228);
nor I_31591 (I539590,I539573,I539457);
nand I_31592 (I539315,I539590,I1254234);
DFFARX1 I_31593 (I539573,I2507,I539341,I539327,);
nand I_31594 (I539635,I539457,I1254219);
nor I_31595 (I539652,I539457,I1254219);
nand I_31596 (I539321,I539440,I539652);
not I_31597 (I539683,I1254210);
nor I_31598 (I539700,I539683,I539635);
DFFARX1 I_31599 (I539700,I2507,I539341,I539309,);
nor I_31600 (I539731,I539683,I1254222);
and I_31601 (I539748,I539731,I1254216);
or I_31602 (I539765,I539748,I1254213);
DFFARX1 I_31603 (I539765,I2507,I539341,I539791,);
nor I_31604 (I539799,I539791,I539415);
nor I_31605 (I539318,I539367,I539799);
not I_31606 (I539830,I539791);
nor I_31607 (I539847,I539830,I539525);
DFFARX1 I_31608 (I539847,I2507,I539341,I539324,);
nand I_31609 (I539878,I539830,I539457);
nor I_31610 (I539312,I539683,I539878);
not I_31611 (I539936,I2514);
DFFARX1 I_31612 (I87016,I2507,I539936,I539962,);
DFFARX1 I_31613 (I539962,I2507,I539936,I539979,);
not I_31614 (I539928,I539979);
DFFARX1 I_31615 (I87028,I2507,I539936,I540010,);
not I_31616 (I540018,I87019);
nor I_31617 (I540035,I539962,I540018);
not I_31618 (I540052,I87010);
not I_31619 (I540069,I87007);
nand I_31620 (I540086,I540069,I87010);
nor I_31621 (I540103,I540018,I540086);
nor I_31622 (I540120,I540010,I540103);
DFFARX1 I_31623 (I540069,I2507,I539936,I539925,);
nor I_31624 (I540151,I87007,I87007);
nand I_31625 (I540168,I540151,I87025);
nor I_31626 (I540185,I540168,I540052);
nand I_31627 (I539910,I540185,I87019);
DFFARX1 I_31628 (I540168,I2507,I539936,I539922,);
nand I_31629 (I540230,I540052,I87007);
nor I_31630 (I540247,I540052,I87007);
nand I_31631 (I539916,I540035,I540247);
not I_31632 (I540278,I87031);
nor I_31633 (I540295,I540278,I540230);
DFFARX1 I_31634 (I540295,I2507,I539936,I539904,);
nor I_31635 (I540326,I540278,I87010);
and I_31636 (I540343,I540326,I87013);
or I_31637 (I540360,I540343,I87022);
DFFARX1 I_31638 (I540360,I2507,I539936,I540386,);
nor I_31639 (I540394,I540386,I540010);
nor I_31640 (I539913,I539962,I540394);
not I_31641 (I540425,I540386);
nor I_31642 (I540442,I540425,I540120);
DFFARX1 I_31643 (I540442,I2507,I539936,I539919,);
nand I_31644 (I540473,I540425,I540052);
nor I_31645 (I539907,I540278,I540473);
not I_31646 (I540531,I2514);
DFFARX1 I_31647 (I1020239,I2507,I540531,I540557,);
DFFARX1 I_31648 (I540557,I2507,I540531,I540574,);
not I_31649 (I540523,I540574);
DFFARX1 I_31650 (I1020242,I2507,I540531,I540605,);
not I_31651 (I540613,I1020245);
nor I_31652 (I540630,I540557,I540613);
not I_31653 (I540647,I1020257);
not I_31654 (I540664,I1020248);
nand I_31655 (I540681,I540664,I1020257);
nor I_31656 (I540698,I540613,I540681);
nor I_31657 (I540715,I540605,I540698);
DFFARX1 I_31658 (I540664,I2507,I540531,I540520,);
nor I_31659 (I540746,I1020248,I1020254);
nand I_31660 (I540763,I540746,I1020242);
nor I_31661 (I540780,I540763,I540647);
nand I_31662 (I540505,I540780,I1020245);
DFFARX1 I_31663 (I540763,I2507,I540531,I540517,);
nand I_31664 (I540825,I540647,I1020248);
nor I_31665 (I540842,I540647,I1020248);
nand I_31666 (I540511,I540630,I540842);
not I_31667 (I540873,I1020245);
nor I_31668 (I540890,I540873,I540825);
DFFARX1 I_31669 (I540890,I2507,I540531,I540499,);
nor I_31670 (I540921,I540873,I1020251);
and I_31671 (I540938,I540921,I1020239);
or I_31672 (I540955,I540938,I1020260);
DFFARX1 I_31673 (I540955,I2507,I540531,I540981,);
nor I_31674 (I540989,I540981,I540605);
nor I_31675 (I540508,I540557,I540989);
not I_31676 (I541020,I540981);
nor I_31677 (I541037,I541020,I540715);
DFFARX1 I_31678 (I541037,I2507,I540531,I540514,);
nand I_31679 (I541068,I541020,I540647);
nor I_31680 (I540502,I540873,I541068);
not I_31681 (I541126,I2514);
DFFARX1 I_31682 (I841255,I2507,I541126,I541152,);
DFFARX1 I_31683 (I541152,I2507,I541126,I541169,);
not I_31684 (I541118,I541169);
DFFARX1 I_31685 (I841252,I2507,I541126,I541200,);
not I_31686 (I541208,I841252);
nor I_31687 (I541225,I541152,I541208);
not I_31688 (I541242,I841249);
not I_31689 (I541259,I841264);
nand I_31690 (I541276,I541259,I841249);
nor I_31691 (I541293,I541208,I541276);
nor I_31692 (I541310,I541200,I541293);
DFFARX1 I_31693 (I541259,I2507,I541126,I541115,);
nor I_31694 (I541341,I841264,I841258);
nand I_31695 (I541358,I541341,I841246);
nor I_31696 (I541375,I541358,I541242);
nand I_31697 (I541100,I541375,I841252);
DFFARX1 I_31698 (I541358,I2507,I541126,I541112,);
nand I_31699 (I541420,I541242,I841264);
nor I_31700 (I541437,I541242,I841264);
nand I_31701 (I541106,I541225,I541437);
not I_31702 (I541468,I841267);
nor I_31703 (I541485,I541468,I541420);
DFFARX1 I_31704 (I541485,I2507,I541126,I541094,);
nor I_31705 (I541516,I541468,I841246);
and I_31706 (I541533,I541516,I841261);
or I_31707 (I541550,I541533,I841249);
DFFARX1 I_31708 (I541550,I2507,I541126,I541576,);
nor I_31709 (I541584,I541576,I541200);
nor I_31710 (I541103,I541152,I541584);
not I_31711 (I541615,I541576);
nor I_31712 (I541632,I541615,I541310);
DFFARX1 I_31713 (I541632,I2507,I541126,I541109,);
nand I_31714 (I541663,I541615,I541242);
nor I_31715 (I541097,I541468,I541663);
not I_31716 (I541721,I2514);
DFFARX1 I_31717 (I609913,I2507,I541721,I541747,);
DFFARX1 I_31718 (I541747,I2507,I541721,I541764,);
not I_31719 (I541713,I541764);
DFFARX1 I_31720 (I609925,I2507,I541721,I541795,);
not I_31721 (I541803,I609910);
nor I_31722 (I541820,I541747,I541803);
not I_31723 (I541837,I609928);
not I_31724 (I541854,I609919);
nand I_31725 (I541871,I541854,I609928);
nor I_31726 (I541888,I541803,I541871);
nor I_31727 (I541905,I541795,I541888);
DFFARX1 I_31728 (I541854,I2507,I541721,I541710,);
nor I_31729 (I541936,I609919,I609931);
nand I_31730 (I541953,I541936,I609934);
nor I_31731 (I541970,I541953,I541837);
nand I_31732 (I541695,I541970,I609910);
DFFARX1 I_31733 (I541953,I2507,I541721,I541707,);
nand I_31734 (I542015,I541837,I609919);
nor I_31735 (I542032,I541837,I609919);
nand I_31736 (I541701,I541820,I542032);
not I_31737 (I542063,I609910);
nor I_31738 (I542080,I542063,I542015);
DFFARX1 I_31739 (I542080,I2507,I541721,I541689,);
nor I_31740 (I542111,I542063,I609922);
and I_31741 (I542128,I542111,I609916);
or I_31742 (I542145,I542128,I609913);
DFFARX1 I_31743 (I542145,I2507,I541721,I542171,);
nor I_31744 (I542179,I542171,I541795);
nor I_31745 (I541698,I541747,I542179);
not I_31746 (I542210,I542171);
nor I_31747 (I542227,I542210,I541905);
DFFARX1 I_31748 (I542227,I2507,I541721,I541704,);
nand I_31749 (I542258,I542210,I541837);
nor I_31750 (I541692,I542063,I542258);
not I_31751 (I542316,I2514);
DFFARX1 I_31752 (I936027,I2507,I542316,I542342,);
not I_31753 (I542350,I542342);
DFFARX1 I_31754 (I936024,I2507,I542316,I542376,);
not I_31755 (I542384,I936021);
nand I_31756 (I542401,I542384,I936048);
not I_31757 (I542418,I542401);
nor I_31758 (I542435,I542418,I936036);
nor I_31759 (I542452,I542350,I542435);
DFFARX1 I_31760 (I542452,I2507,I542316,I542302,);
not I_31761 (I542483,I936036);
nand I_31762 (I542500,I542483,I542418);
and I_31763 (I542517,I542483,I936042);
nand I_31764 (I542534,I542517,I936033);
nor I_31765 (I542299,I542534,I542483);
and I_31766 (I542290,I542376,I542534);
not I_31767 (I542579,I542534);
nand I_31768 (I542293,I542376,I542579);
nor I_31769 (I542287,I542342,I542534);
not I_31770 (I542624,I936030);
nor I_31771 (I542641,I542624,I936042);
nand I_31772 (I542658,I542641,I542483);
nor I_31773 (I542296,I542401,I542658);
nor I_31774 (I542689,I542624,I936045);
and I_31775 (I542706,I542689,I936039);
or I_31776 (I542723,I542706,I936021);
DFFARX1 I_31777 (I542723,I2507,I542316,I542749,);
nor I_31778 (I542757,I542749,I542500);
DFFARX1 I_31779 (I542757,I2507,I542316,I542284,);
DFFARX1 I_31780 (I542749,I2507,I542316,I542308,);
not I_31781 (I542802,I542749);
nor I_31782 (I542819,I542802,I542376);
nor I_31783 (I542836,I542641,I542819);
DFFARX1 I_31784 (I542836,I2507,I542316,I542305,);
not I_31785 (I542894,I2514);
DFFARX1 I_31786 (I362974,I2507,I542894,I542920,);
not I_31787 (I542928,I542920);
DFFARX1 I_31788 (I362989,I2507,I542894,I542954,);
not I_31789 (I542962,I362992);
nand I_31790 (I542979,I542962,I362971);
not I_31791 (I542996,I542979);
nor I_31792 (I543013,I542996,I362995);
nor I_31793 (I543030,I542928,I543013);
DFFARX1 I_31794 (I543030,I2507,I542894,I542880,);
not I_31795 (I543061,I362995);
nand I_31796 (I543078,I543061,I542996);
and I_31797 (I543095,I543061,I362977);
nand I_31798 (I543112,I543095,I362968);
nor I_31799 (I542877,I543112,I543061);
and I_31800 (I542868,I542954,I543112);
not I_31801 (I543157,I543112);
nand I_31802 (I542871,I542954,I543157);
nor I_31803 (I542865,I542920,I543112);
not I_31804 (I543202,I362968);
nor I_31805 (I543219,I543202,I362977);
nand I_31806 (I543236,I543219,I543061);
nor I_31807 (I542874,I542979,I543236);
nor I_31808 (I543267,I543202,I362983);
and I_31809 (I543284,I543267,I362986);
or I_31810 (I543301,I543284,I362980);
DFFARX1 I_31811 (I543301,I2507,I542894,I543327,);
nor I_31812 (I543335,I543327,I543078);
DFFARX1 I_31813 (I543335,I2507,I542894,I542862,);
DFFARX1 I_31814 (I543327,I2507,I542894,I542886,);
not I_31815 (I543380,I543327);
nor I_31816 (I543397,I543380,I542954);
nor I_31817 (I543414,I543219,I543397);
DFFARX1 I_31818 (I543414,I2507,I542894,I542883,);
not I_31819 (I543472,I2514);
DFFARX1 I_31820 (I1117904,I2507,I543472,I543498,);
not I_31821 (I543506,I543498);
DFFARX1 I_31822 (I1117910,I2507,I543472,I543532,);
not I_31823 (I543540,I1117904);
nand I_31824 (I543557,I543540,I1117907);
not I_31825 (I543574,I543557);
nor I_31826 (I543591,I543574,I1117925);
nor I_31827 (I543608,I543506,I543591);
DFFARX1 I_31828 (I543608,I2507,I543472,I543458,);
not I_31829 (I543639,I1117925);
nand I_31830 (I543656,I543639,I543574);
and I_31831 (I543673,I543639,I1117928);
nand I_31832 (I543690,I543673,I1117907);
nor I_31833 (I543455,I543690,I543639);
and I_31834 (I543446,I543532,I543690);
not I_31835 (I543735,I543690);
nand I_31836 (I543449,I543532,I543735);
nor I_31837 (I543443,I543498,I543690);
not I_31838 (I543780,I1117913);
nor I_31839 (I543797,I543780,I1117928);
nand I_31840 (I543814,I543797,I543639);
nor I_31841 (I543452,I543557,I543814);
nor I_31842 (I543845,I543780,I1117919);
and I_31843 (I543862,I543845,I1117916);
or I_31844 (I543879,I543862,I1117922);
DFFARX1 I_31845 (I543879,I2507,I543472,I543905,);
nor I_31846 (I543913,I543905,I543656);
DFFARX1 I_31847 (I543913,I2507,I543472,I543440,);
DFFARX1 I_31848 (I543905,I2507,I543472,I543464,);
not I_31849 (I543958,I543905);
nor I_31850 (I543975,I543958,I543532);
nor I_31851 (I543992,I543797,I543975);
DFFARX1 I_31852 (I543992,I2507,I543472,I543461,);
not I_31853 (I544050,I2514);
DFFARX1 I_31854 (I1169346,I2507,I544050,I544076,);
not I_31855 (I544084,I544076);
DFFARX1 I_31856 (I1169352,I2507,I544050,I544110,);
not I_31857 (I544118,I1169346);
nand I_31858 (I544135,I544118,I1169349);
not I_31859 (I544152,I544135);
nor I_31860 (I544169,I544152,I1169367);
nor I_31861 (I544186,I544084,I544169);
DFFARX1 I_31862 (I544186,I2507,I544050,I544036,);
not I_31863 (I544217,I1169367);
nand I_31864 (I544234,I544217,I544152);
and I_31865 (I544251,I544217,I1169370);
nand I_31866 (I544268,I544251,I1169349);
nor I_31867 (I544033,I544268,I544217);
and I_31868 (I544024,I544110,I544268);
not I_31869 (I544313,I544268);
nand I_31870 (I544027,I544110,I544313);
nor I_31871 (I544021,I544076,I544268);
not I_31872 (I544358,I1169355);
nor I_31873 (I544375,I544358,I1169370);
nand I_31874 (I544392,I544375,I544217);
nor I_31875 (I544030,I544135,I544392);
nor I_31876 (I544423,I544358,I1169361);
and I_31877 (I544440,I544423,I1169358);
or I_31878 (I544457,I544440,I1169364);
DFFARX1 I_31879 (I544457,I2507,I544050,I544483,);
nor I_31880 (I544491,I544483,I544234);
DFFARX1 I_31881 (I544491,I2507,I544050,I544018,);
DFFARX1 I_31882 (I544483,I2507,I544050,I544042,);
not I_31883 (I544536,I544483);
nor I_31884 (I544553,I544536,I544110);
nor I_31885 (I544570,I544375,I544553);
DFFARX1 I_31886 (I544570,I2507,I544050,I544039,);
not I_31887 (I544628,I2514);
DFFARX1 I_31888 (I1082068,I2507,I544628,I544654,);
not I_31889 (I544662,I544654);
DFFARX1 I_31890 (I1082074,I2507,I544628,I544688,);
not I_31891 (I544696,I1082068);
nand I_31892 (I544713,I544696,I1082071);
not I_31893 (I544730,I544713);
nor I_31894 (I544747,I544730,I1082089);
nor I_31895 (I544764,I544662,I544747);
DFFARX1 I_31896 (I544764,I2507,I544628,I544614,);
not I_31897 (I544795,I1082089);
nand I_31898 (I544812,I544795,I544730);
and I_31899 (I544829,I544795,I1082092);
nand I_31900 (I544846,I544829,I1082071);
nor I_31901 (I544611,I544846,I544795);
and I_31902 (I544602,I544688,I544846);
not I_31903 (I544891,I544846);
nand I_31904 (I544605,I544688,I544891);
nor I_31905 (I544599,I544654,I544846);
not I_31906 (I544936,I1082077);
nor I_31907 (I544953,I544936,I1082092);
nand I_31908 (I544970,I544953,I544795);
nor I_31909 (I544608,I544713,I544970);
nor I_31910 (I545001,I544936,I1082083);
and I_31911 (I545018,I545001,I1082080);
or I_31912 (I545035,I545018,I1082086);
DFFARX1 I_31913 (I545035,I2507,I544628,I545061,);
nor I_31914 (I545069,I545061,I544812);
DFFARX1 I_31915 (I545069,I2507,I544628,I544596,);
DFFARX1 I_31916 (I545061,I2507,I544628,I544620,);
not I_31917 (I545114,I545061);
nor I_31918 (I545131,I545114,I544688);
nor I_31919 (I545148,I544953,I545131);
DFFARX1 I_31920 (I545148,I2507,I544628,I544617,);
not I_31921 (I545206,I2514);
DFFARX1 I_31922 (I639388,I2507,I545206,I545232,);
not I_31923 (I545240,I545232);
DFFARX1 I_31924 (I639400,I2507,I545206,I545266,);
not I_31925 (I545274,I639391);
nand I_31926 (I545291,I545274,I639394);
not I_31927 (I545308,I545291);
nor I_31928 (I545325,I545308,I639397);
nor I_31929 (I545342,I545240,I545325);
DFFARX1 I_31930 (I545342,I2507,I545206,I545192,);
not I_31931 (I545373,I639397);
nand I_31932 (I545390,I545373,I545308);
and I_31933 (I545407,I545373,I639391);
nand I_31934 (I545424,I545407,I639403);
nor I_31935 (I545189,I545424,I545373);
and I_31936 (I545180,I545266,I545424);
not I_31937 (I545469,I545424);
nand I_31938 (I545183,I545266,I545469);
nor I_31939 (I545177,I545232,I545424);
not I_31940 (I545514,I639409);
nor I_31941 (I545531,I545514,I639391);
nand I_31942 (I545548,I545531,I545373);
nor I_31943 (I545186,I545291,I545548);
nor I_31944 (I545579,I545514,I639388);
and I_31945 (I545596,I545579,I639406);
or I_31946 (I545613,I545596,I639412);
DFFARX1 I_31947 (I545613,I2507,I545206,I545639,);
nor I_31948 (I545647,I545639,I545390);
DFFARX1 I_31949 (I545647,I2507,I545206,I545174,);
DFFARX1 I_31950 (I545639,I2507,I545206,I545198,);
not I_31951 (I545692,I545639);
nor I_31952 (I545709,I545692,I545266);
nor I_31953 (I545726,I545531,I545709);
DFFARX1 I_31954 (I545726,I2507,I545206,I545195,);
not I_31955 (I545784,I2514);
DFFARX1 I_31956 (I414235,I2507,I545784,I545810,);
not I_31957 (I545818,I545810);
DFFARX1 I_31958 (I414247,I2507,I545784,I545844,);
not I_31959 (I545852,I414223);
nand I_31960 (I545869,I545852,I414250);
not I_31961 (I545886,I545869);
nor I_31962 (I545903,I545886,I414238);
nor I_31963 (I545920,I545818,I545903);
DFFARX1 I_31964 (I545920,I2507,I545784,I545770,);
not I_31965 (I545951,I414238);
nand I_31966 (I545968,I545951,I545886);
and I_31967 (I545985,I545951,I414223);
nand I_31968 (I546002,I545985,I414226);
nor I_31969 (I545767,I546002,I545951);
and I_31970 (I545758,I545844,I546002);
not I_31971 (I546047,I546002);
nand I_31972 (I545761,I545844,I546047);
nor I_31973 (I545755,I545810,I546002);
not I_31974 (I546092,I414232);
nor I_31975 (I546109,I546092,I414223);
nand I_31976 (I546126,I546109,I545951);
nor I_31977 (I545764,I545869,I546126);
nor I_31978 (I546157,I546092,I414241);
and I_31979 (I546174,I546157,I414229);
or I_31980 (I546191,I546174,I414244);
DFFARX1 I_31981 (I546191,I2507,I545784,I546217,);
nor I_31982 (I546225,I546217,I545968);
DFFARX1 I_31983 (I546225,I2507,I545784,I545752,);
DFFARX1 I_31984 (I546217,I2507,I545784,I545776,);
not I_31985 (I546270,I546217);
nor I_31986 (I546287,I546270,I545844);
nor I_31987 (I546304,I546109,I546287);
DFFARX1 I_31988 (I546304,I2507,I545784,I545773,);
not I_31989 (I546362,I2514);
DFFARX1 I_31990 (I710482,I2507,I546362,I546388,);
not I_31991 (I546396,I546388);
DFFARX1 I_31992 (I710494,I2507,I546362,I546422,);
not I_31993 (I546430,I710485);
nand I_31994 (I546447,I546430,I710488);
not I_31995 (I546464,I546447);
nor I_31996 (I546481,I546464,I710491);
nor I_31997 (I546498,I546396,I546481);
DFFARX1 I_31998 (I546498,I2507,I546362,I546348,);
not I_31999 (I546529,I710491);
nand I_32000 (I546546,I546529,I546464);
and I_32001 (I546563,I546529,I710485);
nand I_32002 (I546580,I546563,I710497);
nor I_32003 (I546345,I546580,I546529);
and I_32004 (I546336,I546422,I546580);
not I_32005 (I546625,I546580);
nand I_32006 (I546339,I546422,I546625);
nor I_32007 (I546333,I546388,I546580);
not I_32008 (I546670,I710503);
nor I_32009 (I546687,I546670,I710485);
nand I_32010 (I546704,I546687,I546529);
nor I_32011 (I546342,I546447,I546704);
nor I_32012 (I546735,I546670,I710482);
and I_32013 (I546752,I546735,I710500);
or I_32014 (I546769,I546752,I710506);
DFFARX1 I_32015 (I546769,I2507,I546362,I546795,);
nor I_32016 (I546803,I546795,I546546);
DFFARX1 I_32017 (I546803,I2507,I546362,I546330,);
DFFARX1 I_32018 (I546795,I2507,I546362,I546354,);
not I_32019 (I546848,I546795);
nor I_32020 (I546865,I546848,I546422);
nor I_32021 (I546882,I546687,I546865);
DFFARX1 I_32022 (I546882,I2507,I546362,I546351,);
not I_32023 (I546940,I2514);
DFFARX1 I_32024 (I1292336,I2507,I546940,I546966,);
not I_32025 (I546974,I546966);
DFFARX1 I_32026 (I1292348,I2507,I546940,I547000,);
not I_32027 (I547008,I1292339);
nand I_32028 (I547025,I547008,I1292327);
not I_32029 (I547042,I547025);
nor I_32030 (I547059,I547042,I1292324);
nor I_32031 (I547076,I546974,I547059);
DFFARX1 I_32032 (I547076,I2507,I546940,I546926,);
not I_32033 (I547107,I1292324);
nand I_32034 (I547124,I547107,I547042);
and I_32035 (I547141,I547107,I1292330);
nand I_32036 (I547158,I547141,I1292327);
nor I_32037 (I546923,I547158,I547107);
and I_32038 (I546914,I547000,I547158);
not I_32039 (I547203,I547158);
nand I_32040 (I546917,I547000,I547203);
nor I_32041 (I546911,I546966,I547158);
not I_32042 (I547248,I1292345);
nor I_32043 (I547265,I547248,I1292330);
nand I_32044 (I547282,I547265,I547107);
nor I_32045 (I546920,I547025,I547282);
nor I_32046 (I547313,I547248,I1292333);
and I_32047 (I547330,I547313,I1292324);
or I_32048 (I547347,I547330,I1292342);
DFFARX1 I_32049 (I547347,I2507,I546940,I547373,);
nor I_32050 (I547381,I547373,I547124);
DFFARX1 I_32051 (I547381,I2507,I546940,I546908,);
DFFARX1 I_32052 (I547373,I2507,I546940,I546932,);
not I_32053 (I547426,I547373);
nor I_32054 (I547443,I547426,I547000);
nor I_32055 (I547460,I547265,I547443);
DFFARX1 I_32056 (I547460,I2507,I546940,I546929,);
not I_32057 (I547518,I2514);
DFFARX1 I_32058 (I1262280,I2507,I547518,I547544,);
not I_32059 (I547552,I547544);
DFFARX1 I_32060 (I1262292,I2507,I547518,I547578,);
not I_32061 (I547586,I1262283);
nand I_32062 (I547603,I547586,I1262271);
not I_32063 (I547620,I547603);
nor I_32064 (I547637,I547620,I1262268);
nor I_32065 (I547654,I547552,I547637);
DFFARX1 I_32066 (I547654,I2507,I547518,I547504,);
not I_32067 (I547685,I1262268);
nand I_32068 (I547702,I547685,I547620);
and I_32069 (I547719,I547685,I1262274);
nand I_32070 (I547736,I547719,I1262271);
nor I_32071 (I547501,I547736,I547685);
and I_32072 (I547492,I547578,I547736);
not I_32073 (I547781,I547736);
nand I_32074 (I547495,I547578,I547781);
nor I_32075 (I547489,I547544,I547736);
not I_32076 (I547826,I1262289);
nor I_32077 (I547843,I547826,I1262274);
nand I_32078 (I547860,I547843,I547685);
nor I_32079 (I547498,I547603,I547860);
nor I_32080 (I547891,I547826,I1262277);
and I_32081 (I547908,I547891,I1262268);
or I_32082 (I547925,I547908,I1262286);
DFFARX1 I_32083 (I547925,I2507,I547518,I547951,);
nor I_32084 (I547959,I547951,I547702);
DFFARX1 I_32085 (I547959,I2507,I547518,I547486,);
DFFARX1 I_32086 (I547951,I2507,I547518,I547510,);
not I_32087 (I548004,I547951);
nor I_32088 (I548021,I548004,I547578);
nor I_32089 (I548038,I547843,I548021);
DFFARX1 I_32090 (I548038,I2507,I547518,I547507,);
not I_32091 (I548096,I2514);
DFFARX1 I_32092 (I776374,I2507,I548096,I548122,);
not I_32093 (I548130,I548122);
DFFARX1 I_32094 (I776386,I2507,I548096,I548156,);
not I_32095 (I548164,I776377);
nand I_32096 (I548181,I548164,I776380);
not I_32097 (I548198,I548181);
nor I_32098 (I548215,I548198,I776383);
nor I_32099 (I548232,I548130,I548215);
DFFARX1 I_32100 (I548232,I2507,I548096,I548082,);
not I_32101 (I548263,I776383);
nand I_32102 (I548280,I548263,I548198);
and I_32103 (I548297,I548263,I776377);
nand I_32104 (I548314,I548297,I776389);
nor I_32105 (I548079,I548314,I548263);
and I_32106 (I548070,I548156,I548314);
not I_32107 (I548359,I548314);
nand I_32108 (I548073,I548156,I548359);
nor I_32109 (I548067,I548122,I548314);
not I_32110 (I548404,I776395);
nor I_32111 (I548421,I548404,I776377);
nand I_32112 (I548438,I548421,I548263);
nor I_32113 (I548076,I548181,I548438);
nor I_32114 (I548469,I548404,I776374);
and I_32115 (I548486,I548469,I776392);
or I_32116 (I548503,I548486,I776398);
DFFARX1 I_32117 (I548503,I2507,I548096,I548529,);
nor I_32118 (I548537,I548529,I548280);
DFFARX1 I_32119 (I548537,I2507,I548096,I548064,);
DFFARX1 I_32120 (I548529,I2507,I548096,I548088,);
not I_32121 (I548582,I548529);
nor I_32122 (I548599,I548582,I548156);
nor I_32123 (I548616,I548421,I548599);
DFFARX1 I_32124 (I548616,I2507,I548096,I548085,);
not I_32125 (I548674,I2514);
DFFARX1 I_32126 (I299734,I2507,I548674,I548700,);
not I_32127 (I548708,I548700);
DFFARX1 I_32128 (I299749,I2507,I548674,I548734,);
not I_32129 (I548742,I299752);
nand I_32130 (I548759,I548742,I299731);
not I_32131 (I548776,I548759);
nor I_32132 (I548793,I548776,I299755);
nor I_32133 (I548810,I548708,I548793);
DFFARX1 I_32134 (I548810,I2507,I548674,I548660,);
not I_32135 (I548841,I299755);
nand I_32136 (I548858,I548841,I548776);
and I_32137 (I548875,I548841,I299737);
nand I_32138 (I548892,I548875,I299728);
nor I_32139 (I548657,I548892,I548841);
and I_32140 (I548648,I548734,I548892);
not I_32141 (I548937,I548892);
nand I_32142 (I548651,I548734,I548937);
nor I_32143 (I548645,I548700,I548892);
not I_32144 (I548982,I299728);
nor I_32145 (I548999,I548982,I299737);
nand I_32146 (I549016,I548999,I548841);
nor I_32147 (I548654,I548759,I549016);
nor I_32148 (I549047,I548982,I299743);
and I_32149 (I549064,I549047,I299746);
or I_32150 (I549081,I549064,I299740);
DFFARX1 I_32151 (I549081,I2507,I548674,I549107,);
nor I_32152 (I549115,I549107,I548858);
DFFARX1 I_32153 (I549115,I2507,I548674,I548642,);
DFFARX1 I_32154 (I549107,I2507,I548674,I548666,);
not I_32155 (I549160,I549107);
nor I_32156 (I549177,I549160,I548734);
nor I_32157 (I549194,I548999,I549177);
DFFARX1 I_32158 (I549194,I2507,I548674,I548663,);
not I_32159 (I549252,I2514);
DFFARX1 I_32160 (I834401,I2507,I549252,I549278,);
not I_32161 (I549286,I549278);
DFFARX1 I_32162 (I834401,I2507,I549252,I549312,);
not I_32163 (I549320,I834398);
nand I_32164 (I549337,I549320,I834413);
not I_32165 (I549354,I549337);
nor I_32166 (I549371,I549354,I834407);
nor I_32167 (I549388,I549286,I549371);
DFFARX1 I_32168 (I549388,I2507,I549252,I549238,);
not I_32169 (I549419,I834407);
nand I_32170 (I549436,I549419,I549354);
and I_32171 (I549453,I549419,I834404);
nand I_32172 (I549470,I549453,I834395);
nor I_32173 (I549235,I549470,I549419);
and I_32174 (I549226,I549312,I549470);
not I_32175 (I549515,I549470);
nand I_32176 (I549229,I549312,I549515);
nor I_32177 (I549223,I549278,I549470);
not I_32178 (I549560,I834416);
nor I_32179 (I549577,I549560,I834404);
nand I_32180 (I549594,I549577,I549419);
nor I_32181 (I549232,I549337,I549594);
nor I_32182 (I549625,I549560,I834395);
and I_32183 (I549642,I549625,I834398);
or I_32184 (I549659,I549642,I834410);
DFFARX1 I_32185 (I549659,I2507,I549252,I549685,);
nor I_32186 (I549693,I549685,I549436);
DFFARX1 I_32187 (I549693,I2507,I549252,I549220,);
DFFARX1 I_32188 (I549685,I2507,I549252,I549244,);
not I_32189 (I549738,I549685);
nor I_32190 (I549755,I549738,I549312);
nor I_32191 (I549772,I549577,I549755);
DFFARX1 I_32192 (I549772,I2507,I549252,I549241,);
not I_32193 (I549830,I2514);
DFFARX1 I_32194 (I641122,I2507,I549830,I549856,);
not I_32195 (I549864,I549856);
DFFARX1 I_32196 (I641134,I2507,I549830,I549890,);
not I_32197 (I549898,I641125);
nand I_32198 (I549915,I549898,I641128);
not I_32199 (I549932,I549915);
nor I_32200 (I549949,I549932,I641131);
nor I_32201 (I549966,I549864,I549949);
DFFARX1 I_32202 (I549966,I2507,I549830,I549816,);
not I_32203 (I549997,I641131);
nand I_32204 (I550014,I549997,I549932);
and I_32205 (I550031,I549997,I641125);
nand I_32206 (I550048,I550031,I641137);
nor I_32207 (I549813,I550048,I549997);
and I_32208 (I549804,I549890,I550048);
not I_32209 (I550093,I550048);
nand I_32210 (I549807,I549890,I550093);
nor I_32211 (I549801,I549856,I550048);
not I_32212 (I550138,I641143);
nor I_32213 (I550155,I550138,I641125);
nand I_32214 (I550172,I550155,I549997);
nor I_32215 (I549810,I549915,I550172);
nor I_32216 (I550203,I550138,I641122);
and I_32217 (I550220,I550203,I641140);
or I_32218 (I550237,I550220,I641146);
DFFARX1 I_32219 (I550237,I2507,I549830,I550263,);
nor I_32220 (I550271,I550263,I550014);
DFFARX1 I_32221 (I550271,I2507,I549830,I549798,);
DFFARX1 I_32222 (I550263,I2507,I549830,I549822,);
not I_32223 (I550316,I550263);
nor I_32224 (I550333,I550316,I549890);
nor I_32225 (I550350,I550155,I550333);
DFFARX1 I_32226 (I550350,I2507,I549830,I549819,);
not I_32227 (I550408,I2514);
DFFARX1 I_32228 (I1039334,I2507,I550408,I550434,);
not I_32229 (I550442,I550434);
DFFARX1 I_32230 (I1039325,I2507,I550408,I550468,);
not I_32231 (I550476,I1039319);
nand I_32232 (I550493,I550476,I1039331);
not I_32233 (I550510,I550493);
nor I_32234 (I550527,I550510,I1039322);
nor I_32235 (I550544,I550442,I550527);
DFFARX1 I_32236 (I550544,I2507,I550408,I550394,);
not I_32237 (I550575,I1039322);
nand I_32238 (I550592,I550575,I550510);
and I_32239 (I550609,I550575,I1039328);
nand I_32240 (I550626,I550609,I1039313);
nor I_32241 (I550391,I550626,I550575);
and I_32242 (I550382,I550468,I550626);
not I_32243 (I550671,I550626);
nand I_32244 (I550385,I550468,I550671);
nor I_32245 (I550379,I550434,I550626);
not I_32246 (I550716,I1039313);
nor I_32247 (I550733,I550716,I1039328);
nand I_32248 (I550750,I550733,I550575);
nor I_32249 (I550388,I550493,I550750);
nor I_32250 (I550781,I550716,I1039316);
and I_32251 (I550798,I550781,I1039319);
or I_32252 (I550815,I550798,I1039316);
DFFARX1 I_32253 (I550815,I2507,I550408,I550841,);
nor I_32254 (I550849,I550841,I550592);
DFFARX1 I_32255 (I550849,I2507,I550408,I550376,);
DFFARX1 I_32256 (I550841,I2507,I550408,I550400,);
not I_32257 (I550894,I550841);
nor I_32258 (I550911,I550894,I550468);
nor I_32259 (I550928,I550733,I550911);
DFFARX1 I_32260 (I550928,I2507,I550408,I550397,);
not I_32261 (I550986,I2514);
DFFARX1 I_32262 (I1004503,I2507,I550986,I551012,);
not I_32263 (I551020,I551012);
DFFARX1 I_32264 (I1004500,I2507,I550986,I551046,);
not I_32265 (I551054,I1004497);
nand I_32266 (I551071,I551054,I1004524);
not I_32267 (I551088,I551071);
nor I_32268 (I551105,I551088,I1004512);
nor I_32269 (I551122,I551020,I551105);
DFFARX1 I_32270 (I551122,I2507,I550986,I550972,);
not I_32271 (I551153,I1004512);
nand I_32272 (I551170,I551153,I551088);
and I_32273 (I551187,I551153,I1004518);
nand I_32274 (I551204,I551187,I1004509);
nor I_32275 (I550969,I551204,I551153);
and I_32276 (I550960,I551046,I551204);
not I_32277 (I551249,I551204);
nand I_32278 (I550963,I551046,I551249);
nor I_32279 (I550957,I551012,I551204);
not I_32280 (I551294,I1004506);
nor I_32281 (I551311,I551294,I1004518);
nand I_32282 (I551328,I551311,I551153);
nor I_32283 (I550966,I551071,I551328);
nor I_32284 (I551359,I551294,I1004521);
and I_32285 (I551376,I551359,I1004515);
or I_32286 (I551393,I551376,I1004497);
DFFARX1 I_32287 (I551393,I2507,I550986,I551419,);
nor I_32288 (I551427,I551419,I551170);
DFFARX1 I_32289 (I551427,I2507,I550986,I550954,);
DFFARX1 I_32290 (I551419,I2507,I550986,I550978,);
not I_32291 (I551472,I551419);
nor I_32292 (I551489,I551472,I551046);
nor I_32293 (I551506,I551311,I551489);
DFFARX1 I_32294 (I551506,I2507,I550986,I550975,);
not I_32295 (I551564,I2514);
DFFARX1 I_32296 (I405531,I2507,I551564,I551590,);
not I_32297 (I551598,I551590);
DFFARX1 I_32298 (I405543,I2507,I551564,I551624,);
not I_32299 (I551632,I405519);
nand I_32300 (I551649,I551632,I405546);
not I_32301 (I551666,I551649);
nor I_32302 (I551683,I551666,I405534);
nor I_32303 (I551700,I551598,I551683);
DFFARX1 I_32304 (I551700,I2507,I551564,I551550,);
not I_32305 (I551731,I405534);
nand I_32306 (I551748,I551731,I551666);
and I_32307 (I551765,I551731,I405519);
nand I_32308 (I551782,I551765,I405522);
nor I_32309 (I551547,I551782,I551731);
and I_32310 (I551538,I551624,I551782);
not I_32311 (I551827,I551782);
nand I_32312 (I551541,I551624,I551827);
nor I_32313 (I551535,I551590,I551782);
not I_32314 (I551872,I405528);
nor I_32315 (I551889,I551872,I405519);
nand I_32316 (I551906,I551889,I551731);
nor I_32317 (I551544,I551649,I551906);
nor I_32318 (I551937,I551872,I405537);
and I_32319 (I551954,I551937,I405525);
or I_32320 (I551971,I551954,I405540);
DFFARX1 I_32321 (I551971,I2507,I551564,I551997,);
nor I_32322 (I552005,I551997,I551748);
DFFARX1 I_32323 (I552005,I2507,I551564,I551532,);
DFFARX1 I_32324 (I551997,I2507,I551564,I551556,);
not I_32325 (I552050,I551997);
nor I_32326 (I552067,I552050,I551624);
nor I_32327 (I552084,I551889,I552067);
DFFARX1 I_32328 (I552084,I2507,I551564,I551553,);
not I_32329 (I552142,I2514);
DFFARX1 I_32330 (I737070,I2507,I552142,I552168,);
not I_32331 (I552176,I552168);
DFFARX1 I_32332 (I737082,I2507,I552142,I552202,);
not I_32333 (I552210,I737073);
nand I_32334 (I552227,I552210,I737076);
not I_32335 (I552244,I552227);
nor I_32336 (I552261,I552244,I737079);
nor I_32337 (I552278,I552176,I552261);
DFFARX1 I_32338 (I552278,I2507,I552142,I552128,);
not I_32339 (I552309,I737079);
nand I_32340 (I552326,I552309,I552244);
and I_32341 (I552343,I552309,I737073);
nand I_32342 (I552360,I552343,I737085);
nor I_32343 (I552125,I552360,I552309);
and I_32344 (I552116,I552202,I552360);
not I_32345 (I552405,I552360);
nand I_32346 (I552119,I552202,I552405);
nor I_32347 (I552113,I552168,I552360);
not I_32348 (I552450,I737091);
nor I_32349 (I552467,I552450,I737073);
nand I_32350 (I552484,I552467,I552309);
nor I_32351 (I552122,I552227,I552484);
nor I_32352 (I552515,I552450,I737070);
and I_32353 (I552532,I552515,I737088);
or I_32354 (I552549,I552532,I737094);
DFFARX1 I_32355 (I552549,I2507,I552142,I552575,);
nor I_32356 (I552583,I552575,I552326);
DFFARX1 I_32357 (I552583,I2507,I552142,I552110,);
DFFARX1 I_32358 (I552575,I2507,I552142,I552134,);
not I_32359 (I552628,I552575);
nor I_32360 (I552645,I552628,I552202);
nor I_32361 (I552662,I552467,I552645);
DFFARX1 I_32362 (I552662,I2507,I552142,I552131,);
not I_32363 (I552720,I2514);
DFFARX1 I_32364 (I25351,I2507,I552720,I552746,);
not I_32365 (I552754,I552746);
DFFARX1 I_32366 (I25354,I2507,I552720,I552780,);
not I_32367 (I552788,I25348);
nand I_32368 (I552805,I552788,I25372);
not I_32369 (I552822,I552805);
nor I_32370 (I552839,I552822,I25351);
nor I_32371 (I552856,I552754,I552839);
DFFARX1 I_32372 (I552856,I2507,I552720,I552706,);
not I_32373 (I552887,I25351);
nand I_32374 (I552904,I552887,I552822);
and I_32375 (I552921,I552887,I25366);
nand I_32376 (I552938,I552921,I25360);
nor I_32377 (I552703,I552938,I552887);
and I_32378 (I552694,I552780,I552938);
not I_32379 (I552983,I552938);
nand I_32380 (I552697,I552780,I552983);
nor I_32381 (I552691,I552746,I552938);
not I_32382 (I553028,I25369);
nor I_32383 (I553045,I553028,I25366);
nand I_32384 (I553062,I553045,I552887);
nor I_32385 (I552700,I552805,I553062);
nor I_32386 (I553093,I553028,I25348);
and I_32387 (I553110,I553093,I25357);
or I_32388 (I553127,I553110,I25363);
DFFARX1 I_32389 (I553127,I2507,I552720,I553153,);
nor I_32390 (I553161,I553153,I552904);
DFFARX1 I_32391 (I553161,I2507,I552720,I552688,);
DFFARX1 I_32392 (I553153,I2507,I552720,I552712,);
not I_32393 (I553206,I553153);
nor I_32394 (I553223,I553206,I552780);
nor I_32395 (I553240,I553045,I553223);
DFFARX1 I_32396 (I553240,I2507,I552720,I552709,);
not I_32397 (I553298,I2514);
DFFARX1 I_32398 (I103895,I2507,I553298,I553324,);
not I_32399 (I553332,I553324);
DFFARX1 I_32400 (I103874,I2507,I553298,I553358,);
not I_32401 (I553366,I103871);
nand I_32402 (I553383,I553366,I103886);
not I_32403 (I553400,I553383);
nor I_32404 (I553417,I553400,I103874);
nor I_32405 (I553434,I553332,I553417);
DFFARX1 I_32406 (I553434,I2507,I553298,I553284,);
not I_32407 (I553465,I103874);
nand I_32408 (I553482,I553465,I553400);
and I_32409 (I553499,I553465,I103877);
nand I_32410 (I553516,I553499,I103892);
nor I_32411 (I553281,I553516,I553465);
and I_32412 (I553272,I553358,I553516);
not I_32413 (I553561,I553516);
nand I_32414 (I553275,I553358,I553561);
nor I_32415 (I553269,I553324,I553516);
not I_32416 (I553606,I103883);
nor I_32417 (I553623,I553606,I103877);
nand I_32418 (I553640,I553623,I553465);
nor I_32419 (I553278,I553383,I553640);
nor I_32420 (I553671,I553606,I103871);
and I_32421 (I553688,I553671,I103880);
or I_32422 (I553705,I553688,I103889);
DFFARX1 I_32423 (I553705,I2507,I553298,I553731,);
nor I_32424 (I553739,I553731,I553482);
DFFARX1 I_32425 (I553739,I2507,I553298,I553266,);
DFFARX1 I_32426 (I553731,I2507,I553298,I553290,);
not I_32427 (I553784,I553731);
nor I_32428 (I553801,I553784,I553358);
nor I_32429 (I553818,I553623,I553801);
DFFARX1 I_32430 (I553818,I2507,I553298,I553287,);
not I_32431 (I553876,I2514);
DFFARX1 I_32432 (I1170502,I2507,I553876,I553902,);
not I_32433 (I553910,I553902);
DFFARX1 I_32434 (I1170508,I2507,I553876,I553936,);
not I_32435 (I553944,I1170502);
nand I_32436 (I553961,I553944,I1170505);
not I_32437 (I553978,I553961);
nor I_32438 (I553995,I553978,I1170523);
nor I_32439 (I554012,I553910,I553995);
DFFARX1 I_32440 (I554012,I2507,I553876,I553862,);
not I_32441 (I554043,I1170523);
nand I_32442 (I554060,I554043,I553978);
and I_32443 (I554077,I554043,I1170526);
nand I_32444 (I554094,I554077,I1170505);
nor I_32445 (I553859,I554094,I554043);
and I_32446 (I553850,I553936,I554094);
not I_32447 (I554139,I554094);
nand I_32448 (I553853,I553936,I554139);
nor I_32449 (I553847,I553902,I554094);
not I_32450 (I554184,I1170511);
nor I_32451 (I554201,I554184,I1170526);
nand I_32452 (I554218,I554201,I554043);
nor I_32453 (I553856,I553961,I554218);
nor I_32454 (I554249,I554184,I1170517);
and I_32455 (I554266,I554249,I1170514);
or I_32456 (I554283,I554266,I1170520);
DFFARX1 I_32457 (I554283,I2507,I553876,I554309,);
nor I_32458 (I554317,I554309,I554060);
DFFARX1 I_32459 (I554317,I2507,I553876,I553844,);
DFFARX1 I_32460 (I554309,I2507,I553876,I553868,);
not I_32461 (I554362,I554309);
nor I_32462 (I554379,I554362,I553936);
nor I_32463 (I554396,I554201,I554379);
DFFARX1 I_32464 (I554396,I2507,I553876,I553865,);
not I_32465 (I554454,I2514);
DFFARX1 I_32466 (I1125418,I2507,I554454,I554480,);
not I_32467 (I554488,I554480);
DFFARX1 I_32468 (I1125424,I2507,I554454,I554514,);
not I_32469 (I554522,I1125418);
nand I_32470 (I554539,I554522,I1125421);
not I_32471 (I554556,I554539);
nor I_32472 (I554573,I554556,I1125439);
nor I_32473 (I554590,I554488,I554573);
DFFARX1 I_32474 (I554590,I2507,I554454,I554440,);
not I_32475 (I554621,I1125439);
nand I_32476 (I554638,I554621,I554556);
and I_32477 (I554655,I554621,I1125442);
nand I_32478 (I554672,I554655,I1125421);
nor I_32479 (I554437,I554672,I554621);
and I_32480 (I554428,I554514,I554672);
not I_32481 (I554717,I554672);
nand I_32482 (I554431,I554514,I554717);
nor I_32483 (I554425,I554480,I554672);
not I_32484 (I554762,I1125427);
nor I_32485 (I554779,I554762,I1125442);
nand I_32486 (I554796,I554779,I554621);
nor I_32487 (I554434,I554539,I554796);
nor I_32488 (I554827,I554762,I1125433);
and I_32489 (I554844,I554827,I1125430);
or I_32490 (I554861,I554844,I1125436);
DFFARX1 I_32491 (I554861,I2507,I554454,I554887,);
nor I_32492 (I554895,I554887,I554638);
DFFARX1 I_32493 (I554895,I2507,I554454,I554422,);
DFFARX1 I_32494 (I554887,I2507,I554454,I554446,);
not I_32495 (I554940,I554887);
nor I_32496 (I554957,I554940,I554514);
nor I_32497 (I554974,I554779,I554957);
DFFARX1 I_32498 (I554974,I2507,I554454,I554443,);
not I_32499 (I555032,I2514);
DFFARX1 I_32500 (I1045505,I2507,I555032,I555058,);
not I_32501 (I555066,I555058);
DFFARX1 I_32502 (I1045496,I2507,I555032,I555092,);
not I_32503 (I555100,I1045490);
nand I_32504 (I555117,I555100,I1045502);
not I_32505 (I555134,I555117);
nor I_32506 (I555151,I555134,I1045493);
nor I_32507 (I555168,I555066,I555151);
DFFARX1 I_32508 (I555168,I2507,I555032,I555018,);
not I_32509 (I555199,I1045493);
nand I_32510 (I555216,I555199,I555134);
and I_32511 (I555233,I555199,I1045499);
nand I_32512 (I555250,I555233,I1045484);
nor I_32513 (I555015,I555250,I555199);
and I_32514 (I555006,I555092,I555250);
not I_32515 (I555295,I555250);
nand I_32516 (I555009,I555092,I555295);
nor I_32517 (I555003,I555058,I555250);
not I_32518 (I555340,I1045484);
nor I_32519 (I555357,I555340,I1045499);
nand I_32520 (I555374,I555357,I555199);
nor I_32521 (I555012,I555117,I555374);
nor I_32522 (I555405,I555340,I1045487);
and I_32523 (I555422,I555405,I1045490);
or I_32524 (I555439,I555422,I1045487);
DFFARX1 I_32525 (I555439,I2507,I555032,I555465,);
nor I_32526 (I555473,I555465,I555216);
DFFARX1 I_32527 (I555473,I2507,I555032,I555000,);
DFFARX1 I_32528 (I555465,I2507,I555032,I555024,);
not I_32529 (I555518,I555465);
nor I_32530 (I555535,I555518,I555092);
nor I_32531 (I555552,I555357,I555535);
DFFARX1 I_32532 (I555552,I2507,I555032,I555021,);
not I_32533 (I555610,I2514);
DFFARX1 I_32534 (I1122528,I2507,I555610,I555636,);
not I_32535 (I555644,I555636);
DFFARX1 I_32536 (I1122534,I2507,I555610,I555670,);
not I_32537 (I555678,I1122528);
nand I_32538 (I555695,I555678,I1122531);
not I_32539 (I555712,I555695);
nor I_32540 (I555729,I555712,I1122549);
nor I_32541 (I555746,I555644,I555729);
DFFARX1 I_32542 (I555746,I2507,I555610,I555596,);
not I_32543 (I555777,I1122549);
nand I_32544 (I555794,I555777,I555712);
and I_32545 (I555811,I555777,I1122552);
nand I_32546 (I555828,I555811,I1122531);
nor I_32547 (I555593,I555828,I555777);
and I_32548 (I555584,I555670,I555828);
not I_32549 (I555873,I555828);
nand I_32550 (I555587,I555670,I555873);
nor I_32551 (I555581,I555636,I555828);
not I_32552 (I555918,I1122537);
nor I_32553 (I555935,I555918,I1122552);
nand I_32554 (I555952,I555935,I555777);
nor I_32555 (I555590,I555695,I555952);
nor I_32556 (I555983,I555918,I1122543);
and I_32557 (I556000,I555983,I1122540);
or I_32558 (I556017,I556000,I1122546);
DFFARX1 I_32559 (I556017,I2507,I555610,I556043,);
nor I_32560 (I556051,I556043,I555794);
DFFARX1 I_32561 (I556051,I2507,I555610,I555578,);
DFFARX1 I_32562 (I556043,I2507,I555610,I555602,);
not I_32563 (I556096,I556043);
nor I_32564 (I556113,I556096,I555670);
nor I_32565 (I556130,I555935,I556113);
DFFARX1 I_32566 (I556130,I2507,I555610,I555599,);
not I_32567 (I556188,I2514);
DFFARX1 I_32568 (I1211796,I2507,I556188,I556214,);
not I_32569 (I556222,I556214);
DFFARX1 I_32570 (I1211790,I2507,I556188,I556248,);
not I_32571 (I556256,I1211799);
nand I_32572 (I556273,I556256,I1211778);
not I_32573 (I556290,I556273);
nor I_32574 (I556307,I556290,I1211787);
nor I_32575 (I556324,I556222,I556307);
DFFARX1 I_32576 (I556324,I2507,I556188,I556174,);
not I_32577 (I556355,I1211787);
nand I_32578 (I556372,I556355,I556290);
and I_32579 (I556389,I556355,I1211802);
nand I_32580 (I556406,I556389,I1211781);
nor I_32581 (I556171,I556406,I556355);
and I_32582 (I556162,I556248,I556406);
not I_32583 (I556451,I556406);
nand I_32584 (I556165,I556248,I556451);
nor I_32585 (I556159,I556214,I556406);
not I_32586 (I556496,I1211784);
nor I_32587 (I556513,I556496,I1211802);
nand I_32588 (I556530,I556513,I556355);
nor I_32589 (I556168,I556273,I556530);
nor I_32590 (I556561,I556496,I1211793);
and I_32591 (I556578,I556561,I1211781);
or I_32592 (I556595,I556578,I1211778);
DFFARX1 I_32593 (I556595,I2507,I556188,I556621,);
nor I_32594 (I556629,I556621,I556372);
DFFARX1 I_32595 (I556629,I2507,I556188,I556156,);
DFFARX1 I_32596 (I556621,I2507,I556188,I556180,);
not I_32597 (I556674,I556621);
nor I_32598 (I556691,I556674,I556248);
nor I_32599 (I556708,I556513,I556691);
DFFARX1 I_32600 (I556708,I2507,I556188,I556177,);
not I_32601 (I556766,I2514);
DFFARX1 I_32602 (I303423,I2507,I556766,I556792,);
not I_32603 (I556800,I556792);
DFFARX1 I_32604 (I303438,I2507,I556766,I556826,);
not I_32605 (I556834,I303441);
nand I_32606 (I556851,I556834,I303420);
not I_32607 (I556868,I556851);
nor I_32608 (I556885,I556868,I303444);
nor I_32609 (I556902,I556800,I556885);
DFFARX1 I_32610 (I556902,I2507,I556766,I556752,);
not I_32611 (I556933,I303444);
nand I_32612 (I556950,I556933,I556868);
and I_32613 (I556967,I556933,I303426);
nand I_32614 (I556984,I556967,I303417);
nor I_32615 (I556749,I556984,I556933);
and I_32616 (I556740,I556826,I556984);
not I_32617 (I557029,I556984);
nand I_32618 (I556743,I556826,I557029);
nor I_32619 (I556737,I556792,I556984);
not I_32620 (I557074,I303417);
nor I_32621 (I557091,I557074,I303426);
nand I_32622 (I557108,I557091,I556933);
nor I_32623 (I556746,I556851,I557108);
nor I_32624 (I557139,I557074,I303432);
and I_32625 (I557156,I557139,I303435);
or I_32626 (I557173,I557156,I303429);
DFFARX1 I_32627 (I557173,I2507,I556766,I557199,);
nor I_32628 (I557207,I557199,I556950);
DFFARX1 I_32629 (I557207,I2507,I556766,I556734,);
DFFARX1 I_32630 (I557199,I2507,I556766,I556758,);
not I_32631 (I557252,I557199);
nor I_32632 (I557269,I557252,I556826);
nor I_32633 (I557286,I557091,I557269);
DFFARX1 I_32634 (I557286,I2507,I556766,I556755,);
not I_32635 (I557344,I2514);
DFFARX1 I_32636 (I82815,I2507,I557344,I557370,);
not I_32637 (I557378,I557370);
DFFARX1 I_32638 (I82794,I2507,I557344,I557404,);
not I_32639 (I557412,I82791);
nand I_32640 (I557429,I557412,I82806);
not I_32641 (I557446,I557429);
nor I_32642 (I557463,I557446,I82794);
nor I_32643 (I557480,I557378,I557463);
DFFARX1 I_32644 (I557480,I2507,I557344,I557330,);
not I_32645 (I557511,I82794);
nand I_32646 (I557528,I557511,I557446);
and I_32647 (I557545,I557511,I82797);
nand I_32648 (I557562,I557545,I82812);
nor I_32649 (I557327,I557562,I557511);
and I_32650 (I557318,I557404,I557562);
not I_32651 (I557607,I557562);
nand I_32652 (I557321,I557404,I557607);
nor I_32653 (I557315,I557370,I557562);
not I_32654 (I557652,I82803);
nor I_32655 (I557669,I557652,I82797);
nand I_32656 (I557686,I557669,I557511);
nor I_32657 (I557324,I557429,I557686);
nor I_32658 (I557717,I557652,I82791);
and I_32659 (I557734,I557717,I82800);
or I_32660 (I557751,I557734,I82809);
DFFARX1 I_32661 (I557751,I2507,I557344,I557777,);
nor I_32662 (I557785,I557777,I557528);
DFFARX1 I_32663 (I557785,I2507,I557344,I557312,);
DFFARX1 I_32664 (I557777,I2507,I557344,I557336,);
not I_32665 (I557830,I557777);
nor I_32666 (I557847,I557830,I557404);
nor I_32667 (I557864,I557669,I557847);
DFFARX1 I_32668 (I557864,I2507,I557344,I557333,);
not I_32669 (I557922,I2514);
DFFARX1 I_32670 (I313963,I2507,I557922,I557948,);
not I_32671 (I557956,I557948);
DFFARX1 I_32672 (I313978,I2507,I557922,I557982,);
not I_32673 (I557990,I313981);
nand I_32674 (I558007,I557990,I313960);
not I_32675 (I558024,I558007);
nor I_32676 (I558041,I558024,I313984);
nor I_32677 (I558058,I557956,I558041);
DFFARX1 I_32678 (I558058,I2507,I557922,I557908,);
not I_32679 (I558089,I313984);
nand I_32680 (I558106,I558089,I558024);
and I_32681 (I558123,I558089,I313966);
nand I_32682 (I558140,I558123,I313957);
nor I_32683 (I557905,I558140,I558089);
and I_32684 (I557896,I557982,I558140);
not I_32685 (I558185,I558140);
nand I_32686 (I557899,I557982,I558185);
nor I_32687 (I557893,I557948,I558140);
not I_32688 (I558230,I313957);
nor I_32689 (I558247,I558230,I313966);
nand I_32690 (I558264,I558247,I558089);
nor I_32691 (I557902,I558007,I558264);
nor I_32692 (I558295,I558230,I313972);
and I_32693 (I558312,I558295,I313975);
or I_32694 (I558329,I558312,I313969);
DFFARX1 I_32695 (I558329,I2507,I557922,I558355,);
nor I_32696 (I558363,I558355,I558106);
DFFARX1 I_32697 (I558363,I2507,I557922,I557890,);
DFFARX1 I_32698 (I558355,I2507,I557922,I557914,);
not I_32699 (I558408,I558355);
nor I_32700 (I558425,I558408,I557982);
nor I_32701 (I558442,I558247,I558425);
DFFARX1 I_32702 (I558442,I2507,I557922,I557911,);
not I_32703 (I558500,I2514);
DFFARX1 I_32704 (I762502,I2507,I558500,I558526,);
not I_32705 (I558534,I558526);
DFFARX1 I_32706 (I762514,I2507,I558500,I558560,);
not I_32707 (I558568,I762505);
nand I_32708 (I558585,I558568,I762508);
not I_32709 (I558602,I558585);
nor I_32710 (I558619,I558602,I762511);
nor I_32711 (I558636,I558534,I558619);
DFFARX1 I_32712 (I558636,I2507,I558500,I558486,);
not I_32713 (I558667,I762511);
nand I_32714 (I558684,I558667,I558602);
and I_32715 (I558701,I558667,I762505);
nand I_32716 (I558718,I558701,I762517);
nor I_32717 (I558483,I558718,I558667);
and I_32718 (I558474,I558560,I558718);
not I_32719 (I558763,I558718);
nand I_32720 (I558477,I558560,I558763);
nor I_32721 (I558471,I558526,I558718);
not I_32722 (I558808,I762523);
nor I_32723 (I558825,I558808,I762505);
nand I_32724 (I558842,I558825,I558667);
nor I_32725 (I558480,I558585,I558842);
nor I_32726 (I558873,I558808,I762502);
and I_32727 (I558890,I558873,I762520);
or I_32728 (I558907,I558890,I762526);
DFFARX1 I_32729 (I558907,I2507,I558500,I558933,);
nor I_32730 (I558941,I558933,I558684);
DFFARX1 I_32731 (I558941,I2507,I558500,I558468,);
DFFARX1 I_32732 (I558933,I2507,I558500,I558492,);
not I_32733 (I558986,I558933);
nor I_32734 (I559003,I558986,I558560);
nor I_32735 (I559020,I558825,I559003);
DFFARX1 I_32736 (I559020,I2507,I558500,I558489,);
not I_32737 (I559078,I2514);
DFFARX1 I_32738 (I367717,I2507,I559078,I559104,);
not I_32739 (I559112,I559104);
DFFARX1 I_32740 (I367732,I2507,I559078,I559138,);
not I_32741 (I559146,I367735);
nand I_32742 (I559163,I559146,I367714);
not I_32743 (I559180,I559163);
nor I_32744 (I559197,I559180,I367738);
nor I_32745 (I559214,I559112,I559197);
DFFARX1 I_32746 (I559214,I2507,I559078,I559064,);
not I_32747 (I559245,I367738);
nand I_32748 (I559262,I559245,I559180);
and I_32749 (I559279,I559245,I367720);
nand I_32750 (I559296,I559279,I367711);
nor I_32751 (I559061,I559296,I559245);
and I_32752 (I559052,I559138,I559296);
not I_32753 (I559341,I559296);
nand I_32754 (I559055,I559138,I559341);
nor I_32755 (I559049,I559104,I559296);
not I_32756 (I559386,I367711);
nor I_32757 (I559403,I559386,I367720);
nand I_32758 (I559420,I559403,I559245);
nor I_32759 (I559058,I559163,I559420);
nor I_32760 (I559451,I559386,I367726);
and I_32761 (I559468,I559451,I367729);
or I_32762 (I559485,I559468,I367723);
DFFARX1 I_32763 (I559485,I2507,I559078,I559511,);
nor I_32764 (I559519,I559511,I559262);
DFFARX1 I_32765 (I559519,I2507,I559078,I559046,);
DFFARX1 I_32766 (I559511,I2507,I559078,I559070,);
not I_32767 (I559564,I559511);
nor I_32768 (I559581,I559564,I559138);
nor I_32769 (I559598,I559403,I559581);
DFFARX1 I_32770 (I559598,I2507,I559078,I559067,);
not I_32771 (I559656,I2514);
DFFARX1 I_32772 (I211530,I2507,I559656,I559682,);
not I_32773 (I559690,I559682);
DFFARX1 I_32774 (I211515,I2507,I559656,I559716,);
not I_32775 (I559724,I211533);
nand I_32776 (I559741,I559724,I211518);
not I_32777 (I559758,I559741);
nor I_32778 (I559775,I559758,I211515);
nor I_32779 (I559792,I559690,I559775);
DFFARX1 I_32780 (I559792,I2507,I559656,I559642,);
not I_32781 (I559823,I211515);
nand I_32782 (I559840,I559823,I559758);
and I_32783 (I559857,I559823,I211518);
nand I_32784 (I559874,I559857,I211539);
nor I_32785 (I559639,I559874,I559823);
and I_32786 (I559630,I559716,I559874);
not I_32787 (I559919,I559874);
nand I_32788 (I559633,I559716,I559919);
nor I_32789 (I559627,I559682,I559874);
not I_32790 (I559964,I211527);
nor I_32791 (I559981,I559964,I211518);
nand I_32792 (I559998,I559981,I559823);
nor I_32793 (I559636,I559741,I559998);
nor I_32794 (I560029,I559964,I211521);
and I_32795 (I560046,I560029,I211536);
or I_32796 (I560063,I560046,I211524);
DFFARX1 I_32797 (I560063,I2507,I559656,I560089,);
nor I_32798 (I560097,I560089,I559840);
DFFARX1 I_32799 (I560097,I2507,I559656,I559624,);
DFFARX1 I_32800 (I560089,I2507,I559656,I559648,);
not I_32801 (I560142,I560089);
nor I_32802 (I560159,I560142,I559716);
nor I_32803 (I560176,I559981,I560159);
DFFARX1 I_32804 (I560176,I2507,I559656,I559645,);
not I_32805 (I560234,I2514);
DFFARX1 I_32806 (I793295,I2507,I560234,I560260,);
not I_32807 (I560268,I560260);
DFFARX1 I_32808 (I793295,I2507,I560234,I560294,);
not I_32809 (I560302,I793292);
nand I_32810 (I560319,I560302,I793307);
not I_32811 (I560336,I560319);
nor I_32812 (I560353,I560336,I793301);
nor I_32813 (I560370,I560268,I560353);
DFFARX1 I_32814 (I560370,I2507,I560234,I560220,);
not I_32815 (I560401,I793301);
nand I_32816 (I560418,I560401,I560336);
and I_32817 (I560435,I560401,I793298);
nand I_32818 (I560452,I560435,I793289);
nor I_32819 (I560217,I560452,I560401);
and I_32820 (I560208,I560294,I560452);
not I_32821 (I560497,I560452);
nand I_32822 (I560211,I560294,I560497);
nor I_32823 (I560205,I560260,I560452);
not I_32824 (I560542,I793310);
nor I_32825 (I560559,I560542,I793298);
nand I_32826 (I560576,I560559,I560401);
nor I_32827 (I560214,I560319,I560576);
nor I_32828 (I560607,I560542,I793289);
and I_32829 (I560624,I560607,I793292);
or I_32830 (I560641,I560624,I793304);
DFFARX1 I_32831 (I560641,I2507,I560234,I560667,);
nor I_32832 (I560675,I560667,I560418);
DFFARX1 I_32833 (I560675,I2507,I560234,I560202,);
DFFARX1 I_32834 (I560667,I2507,I560234,I560226,);
not I_32835 (I560720,I560667);
nor I_32836 (I560737,I560720,I560294);
nor I_32837 (I560754,I560559,I560737);
DFFARX1 I_32838 (I560754,I2507,I560234,I560223,);
not I_32839 (I560812,I2514);
DFFARX1 I_32840 (I262844,I2507,I560812,I560838,);
not I_32841 (I560846,I560838);
DFFARX1 I_32842 (I262859,I2507,I560812,I560872,);
not I_32843 (I560880,I262862);
nand I_32844 (I560897,I560880,I262841);
not I_32845 (I560914,I560897);
nor I_32846 (I560931,I560914,I262865);
nor I_32847 (I560948,I560846,I560931);
DFFARX1 I_32848 (I560948,I2507,I560812,I560798,);
not I_32849 (I560979,I262865);
nand I_32850 (I560996,I560979,I560914);
and I_32851 (I561013,I560979,I262847);
nand I_32852 (I561030,I561013,I262838);
nor I_32853 (I560795,I561030,I560979);
and I_32854 (I560786,I560872,I561030);
not I_32855 (I561075,I561030);
nand I_32856 (I560789,I560872,I561075);
nor I_32857 (I560783,I560838,I561030);
not I_32858 (I561120,I262838);
nor I_32859 (I561137,I561120,I262847);
nand I_32860 (I561154,I561137,I560979);
nor I_32861 (I560792,I560897,I561154);
nor I_32862 (I561185,I561120,I262853);
and I_32863 (I561202,I561185,I262856);
or I_32864 (I561219,I561202,I262850);
DFFARX1 I_32865 (I561219,I2507,I560812,I561245,);
nor I_32866 (I561253,I561245,I560996);
DFFARX1 I_32867 (I561253,I2507,I560812,I560780,);
DFFARX1 I_32868 (I561245,I2507,I560812,I560804,);
not I_32869 (I561298,I561245);
nor I_32870 (I561315,I561298,I560872);
nor I_32871 (I561332,I561137,I561315);
DFFARX1 I_32872 (I561332,I2507,I560812,I560801,);
not I_32873 (I561390,I2514);
DFFARX1 I_32874 (I307112,I2507,I561390,I561416,);
not I_32875 (I561424,I561416);
DFFARX1 I_32876 (I307127,I2507,I561390,I561450,);
not I_32877 (I561458,I307130);
nand I_32878 (I561475,I561458,I307109);
not I_32879 (I561492,I561475);
nor I_32880 (I561509,I561492,I307133);
nor I_32881 (I561526,I561424,I561509);
DFFARX1 I_32882 (I561526,I2507,I561390,I561376,);
not I_32883 (I561557,I307133);
nand I_32884 (I561574,I561557,I561492);
and I_32885 (I561591,I561557,I307115);
nand I_32886 (I561608,I561591,I307106);
nor I_32887 (I561373,I561608,I561557);
and I_32888 (I561364,I561450,I561608);
not I_32889 (I561653,I561608);
nand I_32890 (I561367,I561450,I561653);
nor I_32891 (I561361,I561416,I561608);
not I_32892 (I561698,I307106);
nor I_32893 (I561715,I561698,I307115);
nand I_32894 (I561732,I561715,I561557);
nor I_32895 (I561370,I561475,I561732);
nor I_32896 (I561763,I561698,I307121);
and I_32897 (I561780,I561763,I307124);
or I_32898 (I561797,I561780,I307118);
DFFARX1 I_32899 (I561797,I2507,I561390,I561823,);
nor I_32900 (I561831,I561823,I561574);
DFFARX1 I_32901 (I561831,I2507,I561390,I561358,);
DFFARX1 I_32902 (I561823,I2507,I561390,I561382,);
not I_32903 (I561876,I561823);
nor I_32904 (I561893,I561876,I561450);
nor I_32905 (I561910,I561715,I561893);
DFFARX1 I_32906 (I561910,I2507,I561390,I561379,);
not I_32907 (I561968,I2514);
DFFARX1 I_32908 (I253885,I2507,I561968,I561994,);
not I_32909 (I562002,I561994);
DFFARX1 I_32910 (I253900,I2507,I561968,I562028,);
not I_32911 (I562036,I253903);
nand I_32912 (I562053,I562036,I253882);
not I_32913 (I562070,I562053);
nor I_32914 (I562087,I562070,I253906);
nor I_32915 (I562104,I562002,I562087);
DFFARX1 I_32916 (I562104,I2507,I561968,I561954,);
not I_32917 (I562135,I253906);
nand I_32918 (I562152,I562135,I562070);
and I_32919 (I562169,I562135,I253888);
nand I_32920 (I562186,I562169,I253879);
nor I_32921 (I561951,I562186,I562135);
and I_32922 (I561942,I562028,I562186);
not I_32923 (I562231,I562186);
nand I_32924 (I561945,I562028,I562231);
nor I_32925 (I561939,I561994,I562186);
not I_32926 (I562276,I253879);
nor I_32927 (I562293,I562276,I253888);
nand I_32928 (I562310,I562293,I562135);
nor I_32929 (I561948,I562053,I562310);
nor I_32930 (I562341,I562276,I253894);
and I_32931 (I562358,I562341,I253897);
or I_32932 (I562375,I562358,I253891);
DFFARX1 I_32933 (I562375,I2507,I561968,I562401,);
nor I_32934 (I562409,I562401,I562152);
DFFARX1 I_32935 (I562409,I2507,I561968,I561936,);
DFFARX1 I_32936 (I562401,I2507,I561968,I561960,);
not I_32937 (I562454,I562401);
nor I_32938 (I562471,I562454,I562028);
nor I_32939 (I562488,I562293,I562471);
DFFARX1 I_32940 (I562488,I2507,I561968,I561957,);
not I_32941 (I562546,I2514);
DFFARX1 I_32942 (I881831,I2507,I562546,I562572,);
not I_32943 (I562580,I562572);
DFFARX1 I_32944 (I881831,I2507,I562546,I562606,);
not I_32945 (I562614,I881828);
nand I_32946 (I562631,I562614,I881843);
not I_32947 (I562648,I562631);
nor I_32948 (I562665,I562648,I881837);
nor I_32949 (I562682,I562580,I562665);
DFFARX1 I_32950 (I562682,I2507,I562546,I562532,);
not I_32951 (I562713,I881837);
nand I_32952 (I562730,I562713,I562648);
and I_32953 (I562747,I562713,I881834);
nand I_32954 (I562764,I562747,I881825);
nor I_32955 (I562529,I562764,I562713);
and I_32956 (I562520,I562606,I562764);
not I_32957 (I562809,I562764);
nand I_32958 (I562523,I562606,I562809);
nor I_32959 (I562517,I562572,I562764);
not I_32960 (I562854,I881846);
nor I_32961 (I562871,I562854,I881834);
nand I_32962 (I562888,I562871,I562713);
nor I_32963 (I562526,I562631,I562888);
nor I_32964 (I562919,I562854,I881825);
and I_32965 (I562936,I562919,I881828);
or I_32966 (I562953,I562936,I881840);
DFFARX1 I_32967 (I562953,I2507,I562546,I562979,);
nor I_32968 (I562987,I562979,I562730);
DFFARX1 I_32969 (I562987,I2507,I562546,I562514,);
DFFARX1 I_32970 (I562979,I2507,I562546,I562538,);
not I_32971 (I563032,I562979);
nor I_32972 (I563049,I563032,I562606);
nor I_32973 (I563066,I562871,I563049);
DFFARX1 I_32974 (I563066,I2507,I562546,I562535,);
not I_32975 (I563124,I2514);
DFFARX1 I_32976 (I3124,I2507,I563124,I563150,);
not I_32977 (I563158,I563150);
DFFARX1 I_32978 (I3112,I2507,I563124,I563184,);
not I_32979 (I563192,I3121);
nand I_32980 (I563209,I563192,I3118);
not I_32981 (I563226,I563209);
nor I_32982 (I563243,I563226,I3127);
nor I_32983 (I563260,I563158,I563243);
DFFARX1 I_32984 (I563260,I2507,I563124,I563110,);
not I_32985 (I563291,I3127);
nand I_32986 (I563308,I563291,I563226);
and I_32987 (I563325,I563291,I3115);
nand I_32988 (I563342,I563325,I3118);
nor I_32989 (I563107,I563342,I563291);
and I_32990 (I563098,I563184,I563342);
not I_32991 (I563387,I563342);
nand I_32992 (I563101,I563184,I563387);
nor I_32993 (I563095,I563150,I563342);
not I_32994 (I563432,I3133);
nor I_32995 (I563449,I563432,I3115);
nand I_32996 (I563466,I563449,I563291);
nor I_32997 (I563104,I563209,I563466);
nor I_32998 (I563497,I563432,I3115);
and I_32999 (I563514,I563497,I3130);
or I_33000 (I563531,I563514,I3112);
DFFARX1 I_33001 (I563531,I2507,I563124,I563557,);
nor I_33002 (I563565,I563557,I563308);
DFFARX1 I_33003 (I563565,I2507,I563124,I563092,);
DFFARX1 I_33004 (I563557,I2507,I563124,I563116,);
not I_33005 (I563610,I563557);
nor I_33006 (I563627,I563610,I563184);
nor I_33007 (I563644,I563449,I563627);
DFFARX1 I_33008 (I563644,I2507,I563124,I563113,);
not I_33009 (I563702,I2514);
DFFARX1 I_33010 (I734758,I2507,I563702,I563728,);
not I_33011 (I563736,I563728);
DFFARX1 I_33012 (I734770,I2507,I563702,I563762,);
not I_33013 (I563770,I734761);
nand I_33014 (I563787,I563770,I734764);
not I_33015 (I563804,I563787);
nor I_33016 (I563821,I563804,I734767);
nor I_33017 (I563838,I563736,I563821);
DFFARX1 I_33018 (I563838,I2507,I563702,I563688,);
not I_33019 (I563869,I734767);
nand I_33020 (I563886,I563869,I563804);
and I_33021 (I563903,I563869,I734761);
nand I_33022 (I563920,I563903,I734773);
nor I_33023 (I563685,I563920,I563869);
and I_33024 (I563676,I563762,I563920);
not I_33025 (I563965,I563920);
nand I_33026 (I563679,I563762,I563965);
nor I_33027 (I563673,I563728,I563920);
not I_33028 (I564010,I734779);
nor I_33029 (I564027,I564010,I734761);
nand I_33030 (I564044,I564027,I563869);
nor I_33031 (I563682,I563787,I564044);
nor I_33032 (I564075,I564010,I734758);
and I_33033 (I564092,I564075,I734776);
or I_33034 (I564109,I564092,I734782);
DFFARX1 I_33035 (I564109,I2507,I563702,I564135,);
nor I_33036 (I564143,I564135,I563886);
DFFARX1 I_33037 (I564143,I2507,I563702,I563670,);
DFFARX1 I_33038 (I564135,I2507,I563702,I563694,);
not I_33039 (I564188,I564135);
nor I_33040 (I564205,I564188,I563762);
nor I_33041 (I564222,I564027,I564205);
DFFARX1 I_33042 (I564222,I2507,I563702,I563691,);
not I_33043 (I564280,I2514);
DFFARX1 I_33044 (I1098252,I2507,I564280,I564306,);
not I_33045 (I564314,I564306);
DFFARX1 I_33046 (I1098258,I2507,I564280,I564340,);
not I_33047 (I564348,I1098252);
nand I_33048 (I564365,I564348,I1098255);
not I_33049 (I564382,I564365);
nor I_33050 (I564399,I564382,I1098273);
nor I_33051 (I564416,I564314,I564399);
DFFARX1 I_33052 (I564416,I2507,I564280,I564266,);
not I_33053 (I564447,I1098273);
nand I_33054 (I564464,I564447,I564382);
and I_33055 (I564481,I564447,I1098276);
nand I_33056 (I564498,I564481,I1098255);
nor I_33057 (I564263,I564498,I564447);
and I_33058 (I564254,I564340,I564498);
not I_33059 (I564543,I564498);
nand I_33060 (I564257,I564340,I564543);
nor I_33061 (I564251,I564306,I564498);
not I_33062 (I564588,I1098261);
nor I_33063 (I564605,I564588,I1098276);
nand I_33064 (I564622,I564605,I564447);
nor I_33065 (I564260,I564365,I564622);
nor I_33066 (I564653,I564588,I1098267);
and I_33067 (I564670,I564653,I1098264);
or I_33068 (I564687,I564670,I1098270);
DFFARX1 I_33069 (I564687,I2507,I564280,I564713,);
nor I_33070 (I564721,I564713,I564464);
DFFARX1 I_33071 (I564721,I2507,I564280,I564248,);
DFFARX1 I_33072 (I564713,I2507,I564280,I564272,);
not I_33073 (I564766,I564713);
nor I_33074 (I564783,I564766,I564340);
nor I_33075 (I564800,I564605,I564783);
DFFARX1 I_33076 (I564800,I2507,I564280,I564269,);
not I_33077 (I564858,I2514);
DFFARX1 I_33078 (I377787,I2507,I564858,I564884,);
not I_33079 (I564892,I564884);
DFFARX1 I_33080 (I377799,I2507,I564858,I564918,);
not I_33081 (I564926,I377775);
nand I_33082 (I564943,I564926,I377802);
not I_33083 (I564960,I564943);
nor I_33084 (I564977,I564960,I377790);
nor I_33085 (I564994,I564892,I564977);
DFFARX1 I_33086 (I564994,I2507,I564858,I564844,);
not I_33087 (I565025,I377790);
nand I_33088 (I565042,I565025,I564960);
and I_33089 (I565059,I565025,I377775);
nand I_33090 (I565076,I565059,I377778);
nor I_33091 (I564841,I565076,I565025);
and I_33092 (I564832,I564918,I565076);
not I_33093 (I565121,I565076);
nand I_33094 (I564835,I564918,I565121);
nor I_33095 (I564829,I564884,I565076);
not I_33096 (I565166,I377784);
nor I_33097 (I565183,I565166,I377775);
nand I_33098 (I565200,I565183,I565025);
nor I_33099 (I564838,I564943,I565200);
nor I_33100 (I565231,I565166,I377793);
and I_33101 (I565248,I565231,I377781);
or I_33102 (I565265,I565248,I377796);
DFFARX1 I_33103 (I565265,I2507,I564858,I565291,);
nor I_33104 (I565299,I565291,I565042);
DFFARX1 I_33105 (I565299,I2507,I564858,I564826,);
DFFARX1 I_33106 (I565291,I2507,I564858,I564850,);
not I_33107 (I565344,I565291);
nor I_33108 (I565361,I565344,I564918);
nor I_33109 (I565378,I565183,I565361);
DFFARX1 I_33110 (I565378,I2507,I564858,I564847,);
not I_33111 (I565436,I2514);
DFFARX1 I_33112 (I698344,I2507,I565436,I565462,);
not I_33113 (I565470,I565462);
DFFARX1 I_33114 (I698356,I2507,I565436,I565496,);
not I_33115 (I565504,I698347);
nand I_33116 (I565521,I565504,I698350);
not I_33117 (I565538,I565521);
nor I_33118 (I565555,I565538,I698353);
nor I_33119 (I565572,I565470,I565555);
DFFARX1 I_33120 (I565572,I2507,I565436,I565422,);
not I_33121 (I565603,I698353);
nand I_33122 (I565620,I565603,I565538);
and I_33123 (I565637,I565603,I698347);
nand I_33124 (I565654,I565637,I698359);
nor I_33125 (I565419,I565654,I565603);
and I_33126 (I565410,I565496,I565654);
not I_33127 (I565699,I565654);
nand I_33128 (I565413,I565496,I565699);
nor I_33129 (I565407,I565462,I565654);
not I_33130 (I565744,I698365);
nor I_33131 (I565761,I565744,I698347);
nand I_33132 (I565778,I565761,I565603);
nor I_33133 (I565416,I565521,I565778);
nor I_33134 (I565809,I565744,I698344);
and I_33135 (I565826,I565809,I698362);
or I_33136 (I565843,I565826,I698368);
DFFARX1 I_33137 (I565843,I2507,I565436,I565869,);
nor I_33138 (I565877,I565869,I565620);
DFFARX1 I_33139 (I565877,I2507,I565436,I565404,);
DFFARX1 I_33140 (I565869,I2507,I565436,I565428,);
not I_33141 (I565922,I565869);
nor I_33142 (I565939,I565922,I565496);
nor I_33143 (I565956,I565761,I565939);
DFFARX1 I_33144 (I565956,I2507,I565436,I565425,);
not I_33145 (I566014,I2514);
DFFARX1 I_33146 (I914063,I2507,I566014,I566040,);
not I_33147 (I566048,I566040);
DFFARX1 I_33148 (I914060,I2507,I566014,I566074,);
not I_33149 (I566082,I914057);
nand I_33150 (I566099,I566082,I914084);
not I_33151 (I566116,I566099);
nor I_33152 (I566133,I566116,I914072);
nor I_33153 (I566150,I566048,I566133);
DFFARX1 I_33154 (I566150,I2507,I566014,I566000,);
not I_33155 (I566181,I914072);
nand I_33156 (I566198,I566181,I566116);
and I_33157 (I566215,I566181,I914078);
nand I_33158 (I566232,I566215,I914069);
nor I_33159 (I565997,I566232,I566181);
and I_33160 (I565988,I566074,I566232);
not I_33161 (I566277,I566232);
nand I_33162 (I565991,I566074,I566277);
nor I_33163 (I565985,I566040,I566232);
not I_33164 (I566322,I914066);
nor I_33165 (I566339,I566322,I914078);
nand I_33166 (I566356,I566339,I566181);
nor I_33167 (I565994,I566099,I566356);
nor I_33168 (I566387,I566322,I914081);
and I_33169 (I566404,I566387,I914075);
or I_33170 (I566421,I566404,I914057);
DFFARX1 I_33171 (I566421,I2507,I566014,I566447,);
nor I_33172 (I566455,I566447,I566198);
DFFARX1 I_33173 (I566455,I2507,I566014,I565982,);
DFFARX1 I_33174 (I566447,I2507,I566014,I566006,);
not I_33175 (I566500,I566447);
nor I_33176 (I566517,I566500,I566074);
nor I_33177 (I566534,I566339,I566517);
DFFARX1 I_33178 (I566534,I2507,I566014,I566003,);
not I_33179 (I566592,I2514);
DFFARX1 I_33180 (I886931,I2507,I566592,I566618,);
not I_33181 (I566626,I566618);
DFFARX1 I_33182 (I886928,I2507,I566592,I566652,);
not I_33183 (I566660,I886925);
nand I_33184 (I566677,I566660,I886952);
not I_33185 (I566694,I566677);
nor I_33186 (I566711,I566694,I886940);
nor I_33187 (I566728,I566626,I566711);
DFFARX1 I_33188 (I566728,I2507,I566592,I566578,);
not I_33189 (I566759,I886940);
nand I_33190 (I566776,I566759,I566694);
and I_33191 (I566793,I566759,I886946);
nand I_33192 (I566810,I566793,I886937);
nor I_33193 (I566575,I566810,I566759);
and I_33194 (I566566,I566652,I566810);
not I_33195 (I566855,I566810);
nand I_33196 (I566569,I566652,I566855);
nor I_33197 (I566563,I566618,I566810);
not I_33198 (I566900,I886934);
nor I_33199 (I566917,I566900,I886946);
nand I_33200 (I566934,I566917,I566759);
nor I_33201 (I566572,I566677,I566934);
nor I_33202 (I566965,I566900,I886949);
and I_33203 (I566982,I566965,I886943);
or I_33204 (I566999,I566982,I886925);
DFFARX1 I_33205 (I566999,I2507,I566592,I567025,);
nor I_33206 (I567033,I567025,I566776);
DFFARX1 I_33207 (I567033,I2507,I566592,I566560,);
DFFARX1 I_33208 (I567025,I2507,I566592,I566584,);
not I_33209 (I567078,I567025);
nor I_33210 (I567095,I567078,I566652);
nor I_33211 (I567112,I566917,I567095);
DFFARX1 I_33212 (I567112,I2507,I566592,I566581,);
not I_33213 (I567170,I2514);
DFFARX1 I_33214 (I1295804,I2507,I567170,I567196,);
not I_33215 (I567204,I567196);
DFFARX1 I_33216 (I1295816,I2507,I567170,I567230,);
not I_33217 (I567238,I1295807);
nand I_33218 (I567255,I567238,I1295795);
not I_33219 (I567272,I567255);
nor I_33220 (I567289,I567272,I1295792);
nor I_33221 (I567306,I567204,I567289);
DFFARX1 I_33222 (I567306,I2507,I567170,I567156,);
not I_33223 (I567337,I1295792);
nand I_33224 (I567354,I567337,I567272);
and I_33225 (I567371,I567337,I1295798);
nand I_33226 (I567388,I567371,I1295795);
nor I_33227 (I567153,I567388,I567337);
and I_33228 (I567144,I567230,I567388);
not I_33229 (I567433,I567388);
nand I_33230 (I567147,I567230,I567433);
nor I_33231 (I567141,I567196,I567388);
not I_33232 (I567478,I1295813);
nor I_33233 (I567495,I567478,I1295798);
nand I_33234 (I567512,I567495,I567337);
nor I_33235 (I567150,I567255,I567512);
nor I_33236 (I567543,I567478,I1295801);
and I_33237 (I567560,I567543,I1295792);
or I_33238 (I567577,I567560,I1295810);
DFFARX1 I_33239 (I567577,I2507,I567170,I567603,);
nor I_33240 (I567611,I567603,I567354);
DFFARX1 I_33241 (I567611,I2507,I567170,I567138,);
DFFARX1 I_33242 (I567603,I2507,I567170,I567162,);
not I_33243 (I567656,I567603);
nor I_33244 (I567673,I567656,I567230);
nor I_33245 (I567690,I567495,I567673);
DFFARX1 I_33246 (I567690,I2507,I567170,I567159,);
not I_33247 (I567748,I2514);
DFFARX1 I_33248 (I1050554,I2507,I567748,I567774,);
not I_33249 (I567782,I567774);
DFFARX1 I_33250 (I1050545,I2507,I567748,I567808,);
not I_33251 (I567816,I1050539);
nand I_33252 (I567833,I567816,I1050551);
not I_33253 (I567850,I567833);
nor I_33254 (I567867,I567850,I1050542);
nor I_33255 (I567884,I567782,I567867);
DFFARX1 I_33256 (I567884,I2507,I567748,I567734,);
not I_33257 (I567915,I1050542);
nand I_33258 (I567932,I567915,I567850);
and I_33259 (I567949,I567915,I1050548);
nand I_33260 (I567966,I567949,I1050533);
nor I_33261 (I567731,I567966,I567915);
and I_33262 (I567722,I567808,I567966);
not I_33263 (I568011,I567966);
nand I_33264 (I567725,I567808,I568011);
nor I_33265 (I567719,I567774,I567966);
not I_33266 (I568056,I1050533);
nor I_33267 (I568073,I568056,I1050548);
nand I_33268 (I568090,I568073,I567915);
nor I_33269 (I567728,I567833,I568090);
nor I_33270 (I568121,I568056,I1050536);
and I_33271 (I568138,I568121,I1050539);
or I_33272 (I568155,I568138,I1050536);
DFFARX1 I_33273 (I568155,I2507,I567748,I568181,);
nor I_33274 (I568189,I568181,I567932);
DFFARX1 I_33275 (I568189,I2507,I567748,I567716,);
DFFARX1 I_33276 (I568181,I2507,I567748,I567740,);
not I_33277 (I568234,I568181);
nor I_33278 (I568251,I568234,I567808);
nor I_33279 (I568268,I568073,I568251);
DFFARX1 I_33280 (I568268,I2507,I567748,I567737,);
not I_33281 (I568326,I2514);
DFFARX1 I_33282 (I913417,I2507,I568326,I568352,);
not I_33283 (I568360,I568352);
DFFARX1 I_33284 (I913414,I2507,I568326,I568386,);
not I_33285 (I568394,I913411);
nand I_33286 (I568411,I568394,I913438);
not I_33287 (I568428,I568411);
nor I_33288 (I568445,I568428,I913426);
nor I_33289 (I568462,I568360,I568445);
DFFARX1 I_33290 (I568462,I2507,I568326,I568312,);
not I_33291 (I568493,I913426);
nand I_33292 (I568510,I568493,I568428);
and I_33293 (I568527,I568493,I913432);
nand I_33294 (I568544,I568527,I913423);
nor I_33295 (I568309,I568544,I568493);
and I_33296 (I568300,I568386,I568544);
not I_33297 (I568589,I568544);
nand I_33298 (I568303,I568386,I568589);
nor I_33299 (I568297,I568352,I568544);
not I_33300 (I568634,I913420);
nor I_33301 (I568651,I568634,I913432);
nand I_33302 (I568668,I568651,I568493);
nor I_33303 (I568306,I568411,I568668);
nor I_33304 (I568699,I568634,I913435);
and I_33305 (I568716,I568699,I913429);
or I_33306 (I568733,I568716,I913411);
DFFARX1 I_33307 (I568733,I2507,I568326,I568759,);
nor I_33308 (I568767,I568759,I568510);
DFFARX1 I_33309 (I568767,I2507,I568326,I568294,);
DFFARX1 I_33310 (I568759,I2507,I568326,I568318,);
not I_33311 (I568812,I568759);
nor I_33312 (I568829,I568812,I568386);
nor I_33313 (I568846,I568651,I568829);
DFFARX1 I_33314 (I568846,I2507,I568326,I568315,);
not I_33315 (I568904,I2514);
DFFARX1 I_33316 (I342421,I2507,I568904,I568930,);
not I_33317 (I568938,I568930);
DFFARX1 I_33318 (I342436,I2507,I568904,I568964,);
not I_33319 (I568972,I342439);
nand I_33320 (I568989,I568972,I342418);
not I_33321 (I569006,I568989);
nor I_33322 (I569023,I569006,I342442);
nor I_33323 (I569040,I568938,I569023);
DFFARX1 I_33324 (I569040,I2507,I568904,I568890,);
not I_33325 (I569071,I342442);
nand I_33326 (I569088,I569071,I569006);
and I_33327 (I569105,I569071,I342424);
nand I_33328 (I569122,I569105,I342415);
nor I_33329 (I568887,I569122,I569071);
and I_33330 (I568878,I568964,I569122);
not I_33331 (I569167,I569122);
nand I_33332 (I568881,I568964,I569167);
nor I_33333 (I568875,I568930,I569122);
not I_33334 (I569212,I342415);
nor I_33335 (I569229,I569212,I342424);
nand I_33336 (I569246,I569229,I569071);
nor I_33337 (I568884,I568989,I569246);
nor I_33338 (I569277,I569212,I342430);
and I_33339 (I569294,I569277,I342433);
or I_33340 (I569311,I569294,I342427);
DFFARX1 I_33341 (I569311,I2507,I568904,I569337,);
nor I_33342 (I569345,I569337,I569088);
DFFARX1 I_33343 (I569345,I2507,I568904,I568872,);
DFFARX1 I_33344 (I569337,I2507,I568904,I568896,);
not I_33345 (I569390,I569337);
nor I_33346 (I569407,I569390,I568964);
nor I_33347 (I569424,I569229,I569407);
DFFARX1 I_33348 (I569424,I2507,I568904,I568893,);
not I_33349 (I569482,I2514);
DFFARX1 I_33350 (I472443,I2507,I569482,I569508,);
not I_33351 (I569516,I569508);
DFFARX1 I_33352 (I472455,I2507,I569482,I569542,);
not I_33353 (I569550,I472431);
nand I_33354 (I569567,I569550,I472458);
not I_33355 (I569584,I569567);
nor I_33356 (I569601,I569584,I472446);
nor I_33357 (I569618,I569516,I569601);
DFFARX1 I_33358 (I569618,I2507,I569482,I569468,);
not I_33359 (I569649,I472446);
nand I_33360 (I569666,I569649,I569584);
and I_33361 (I569683,I569649,I472431);
nand I_33362 (I569700,I569683,I472434);
nor I_33363 (I569465,I569700,I569649);
and I_33364 (I569456,I569542,I569700);
not I_33365 (I569745,I569700);
nand I_33366 (I569459,I569542,I569745);
nor I_33367 (I569453,I569508,I569700);
not I_33368 (I569790,I472440);
nor I_33369 (I569807,I569790,I472431);
nand I_33370 (I569824,I569807,I569649);
nor I_33371 (I569462,I569567,I569824);
nor I_33372 (I569855,I569790,I472449);
and I_33373 (I569872,I569855,I472437);
or I_33374 (I569889,I569872,I472452);
DFFARX1 I_33375 (I569889,I2507,I569482,I569915,);
nor I_33376 (I569923,I569915,I569666);
DFFARX1 I_33377 (I569923,I2507,I569482,I569450,);
DFFARX1 I_33378 (I569915,I2507,I569482,I569474,);
not I_33379 (I569968,I569915);
nor I_33380 (I569985,I569968,I569542);
nor I_33381 (I570002,I569807,I569985);
DFFARX1 I_33382 (I570002,I2507,I569482,I569471,);
not I_33383 (I570060,I2514);
DFFARX1 I_33384 (I322395,I2507,I570060,I570086,);
not I_33385 (I570094,I570086);
DFFARX1 I_33386 (I322410,I2507,I570060,I570120,);
not I_33387 (I570128,I322413);
nand I_33388 (I570145,I570128,I322392);
not I_33389 (I570162,I570145);
nor I_33390 (I570179,I570162,I322416);
nor I_33391 (I570196,I570094,I570179);
DFFARX1 I_33392 (I570196,I2507,I570060,I570046,);
not I_33393 (I570227,I322416);
nand I_33394 (I570244,I570227,I570162);
and I_33395 (I570261,I570227,I322398);
nand I_33396 (I570278,I570261,I322389);
nor I_33397 (I570043,I570278,I570227);
and I_33398 (I570034,I570120,I570278);
not I_33399 (I570323,I570278);
nand I_33400 (I570037,I570120,I570323);
nor I_33401 (I570031,I570086,I570278);
not I_33402 (I570368,I322389);
nor I_33403 (I570385,I570368,I322398);
nand I_33404 (I570402,I570385,I570227);
nor I_33405 (I570040,I570145,I570402);
nor I_33406 (I570433,I570368,I322404);
and I_33407 (I570450,I570433,I322407);
or I_33408 (I570467,I570450,I322401);
DFFARX1 I_33409 (I570467,I2507,I570060,I570493,);
nor I_33410 (I570501,I570493,I570244);
DFFARX1 I_33411 (I570501,I2507,I570060,I570028,);
DFFARX1 I_33412 (I570493,I2507,I570060,I570052,);
not I_33413 (I570546,I570493);
nor I_33414 (I570563,I570546,I570120);
nor I_33415 (I570580,I570385,I570563);
DFFARX1 I_33416 (I570580,I2507,I570060,I570049,);
not I_33417 (I570638,I2514);
DFFARX1 I_33418 (I254412,I2507,I570638,I570664,);
not I_33419 (I570672,I570664);
DFFARX1 I_33420 (I254427,I2507,I570638,I570698,);
not I_33421 (I570706,I254430);
nand I_33422 (I570723,I570706,I254409);
not I_33423 (I570740,I570723);
nor I_33424 (I570757,I570740,I254433);
nor I_33425 (I570774,I570672,I570757);
DFFARX1 I_33426 (I570774,I2507,I570638,I570624,);
not I_33427 (I570805,I254433);
nand I_33428 (I570822,I570805,I570740);
and I_33429 (I570839,I570805,I254415);
nand I_33430 (I570856,I570839,I254406);
nor I_33431 (I570621,I570856,I570805);
and I_33432 (I570612,I570698,I570856);
not I_33433 (I570901,I570856);
nand I_33434 (I570615,I570698,I570901);
nor I_33435 (I570609,I570664,I570856);
not I_33436 (I570946,I254406);
nor I_33437 (I570963,I570946,I254415);
nand I_33438 (I570980,I570963,I570805);
nor I_33439 (I570618,I570723,I570980);
nor I_33440 (I571011,I570946,I254421);
and I_33441 (I571028,I571011,I254424);
or I_33442 (I571045,I571028,I254418);
DFFARX1 I_33443 (I571045,I2507,I570638,I571071,);
nor I_33444 (I571079,I571071,I570822);
DFFARX1 I_33445 (I571079,I2507,I570638,I570606,);
DFFARX1 I_33446 (I571071,I2507,I570638,I570630,);
not I_33447 (I571124,I571071);
nor I_33448 (I571141,I571124,I570698);
nor I_33449 (I571158,I570963,I571141);
DFFARX1 I_33450 (I571158,I2507,I570638,I570627,);
not I_33451 (I571216,I2514);
DFFARX1 I_33452 (I274965,I2507,I571216,I571242,);
not I_33453 (I571250,I571242);
DFFARX1 I_33454 (I274980,I2507,I571216,I571276,);
not I_33455 (I571284,I274983);
nand I_33456 (I571301,I571284,I274962);
not I_33457 (I571318,I571301);
nor I_33458 (I571335,I571318,I274986);
nor I_33459 (I571352,I571250,I571335);
DFFARX1 I_33460 (I571352,I2507,I571216,I571202,);
not I_33461 (I571383,I274986);
nand I_33462 (I571400,I571383,I571318);
and I_33463 (I571417,I571383,I274968);
nand I_33464 (I571434,I571417,I274959);
nor I_33465 (I571199,I571434,I571383);
and I_33466 (I571190,I571276,I571434);
not I_33467 (I571479,I571434);
nand I_33468 (I571193,I571276,I571479);
nor I_33469 (I571187,I571242,I571434);
not I_33470 (I571524,I274959);
nor I_33471 (I571541,I571524,I274968);
nand I_33472 (I571558,I571541,I571383);
nor I_33473 (I571196,I571301,I571558);
nor I_33474 (I571589,I571524,I274974);
and I_33475 (I571606,I571589,I274977);
or I_33476 (I571623,I571606,I274971);
DFFARX1 I_33477 (I571623,I2507,I571216,I571649,);
nor I_33478 (I571657,I571649,I571400);
DFFARX1 I_33479 (I571657,I2507,I571216,I571184,);
DFFARX1 I_33480 (I571649,I2507,I571216,I571208,);
not I_33481 (I571702,I571649);
nor I_33482 (I571719,I571702,I571276);
nor I_33483 (I571736,I571541,I571719);
DFFARX1 I_33484 (I571736,I2507,I571216,I571205,);
not I_33485 (I571794,I2514);
DFFARX1 I_33486 (I811740,I2507,I571794,I571820,);
not I_33487 (I571828,I571820);
DFFARX1 I_33488 (I811740,I2507,I571794,I571854,);
not I_33489 (I571862,I811737);
nand I_33490 (I571879,I571862,I811752);
not I_33491 (I571896,I571879);
nor I_33492 (I571913,I571896,I811746);
nor I_33493 (I571930,I571828,I571913);
DFFARX1 I_33494 (I571930,I2507,I571794,I571780,);
not I_33495 (I571961,I811746);
nand I_33496 (I571978,I571961,I571896);
and I_33497 (I571995,I571961,I811743);
nand I_33498 (I572012,I571995,I811734);
nor I_33499 (I571777,I572012,I571961);
and I_33500 (I571768,I571854,I572012);
not I_33501 (I572057,I572012);
nand I_33502 (I571771,I571854,I572057);
nor I_33503 (I571765,I571820,I572012);
not I_33504 (I572102,I811755);
nor I_33505 (I572119,I572102,I811743);
nand I_33506 (I572136,I572119,I571961);
nor I_33507 (I571774,I571879,I572136);
nor I_33508 (I572167,I572102,I811734);
and I_33509 (I572184,I572167,I811737);
or I_33510 (I572201,I572184,I811749);
DFFARX1 I_33511 (I572201,I2507,I571794,I572227,);
nor I_33512 (I572235,I572227,I571978);
DFFARX1 I_33513 (I572235,I2507,I571794,I571762,);
DFFARX1 I_33514 (I572227,I2507,I571794,I571786,);
not I_33515 (I572280,I572227);
nor I_33516 (I572297,I572280,I571854);
nor I_33517 (I572314,I572119,I572297);
DFFARX1 I_33518 (I572314,I2507,I571794,I571783,);
not I_33519 (I572372,I2514);
DFFARX1 I_33520 (I1363027,I2507,I572372,I572398,);
not I_33521 (I572406,I572398);
DFFARX1 I_33522 (I1363027,I2507,I572372,I572432,);
not I_33523 (I572440,I1363051);
nand I_33524 (I572457,I572440,I1363033);
not I_33525 (I572474,I572457);
nor I_33526 (I572491,I572474,I1363048);
nor I_33527 (I572508,I572406,I572491);
DFFARX1 I_33528 (I572508,I2507,I572372,I572358,);
not I_33529 (I572539,I1363048);
nand I_33530 (I572556,I572539,I572474);
and I_33531 (I572573,I572539,I1363030);
nand I_33532 (I572590,I572573,I1363039);
nor I_33533 (I572355,I572590,I572539);
and I_33534 (I572346,I572432,I572590);
not I_33535 (I572635,I572590);
nand I_33536 (I572349,I572432,I572635);
nor I_33537 (I572343,I572398,I572590);
not I_33538 (I572680,I1363036);
nor I_33539 (I572697,I572680,I1363030);
nand I_33540 (I572714,I572697,I572539);
nor I_33541 (I572352,I572457,I572714);
nor I_33542 (I572745,I572680,I1363045);
and I_33543 (I572762,I572745,I1363054);
or I_33544 (I572779,I572762,I1363042);
DFFARX1 I_33545 (I572779,I2507,I572372,I572805,);
nor I_33546 (I572813,I572805,I572556);
DFFARX1 I_33547 (I572813,I2507,I572372,I572340,);
DFFARX1 I_33548 (I572805,I2507,I572372,I572364,);
not I_33549 (I572858,I572805);
nor I_33550 (I572875,I572858,I572432);
nor I_33551 (I572892,I572697,I572875);
DFFARX1 I_33552 (I572892,I2507,I572372,I572361,);
not I_33553 (I572950,I2514);
DFFARX1 I_33554 (I393563,I2507,I572950,I572976,);
not I_33555 (I572984,I572976);
DFFARX1 I_33556 (I393575,I2507,I572950,I573010,);
not I_33557 (I573018,I393551);
nand I_33558 (I573035,I573018,I393578);
not I_33559 (I573052,I573035);
nor I_33560 (I573069,I573052,I393566);
nor I_33561 (I573086,I572984,I573069);
DFFARX1 I_33562 (I573086,I2507,I572950,I572936,);
not I_33563 (I573117,I393566);
nand I_33564 (I573134,I573117,I573052);
and I_33565 (I573151,I573117,I393551);
nand I_33566 (I573168,I573151,I393554);
nor I_33567 (I572933,I573168,I573117);
and I_33568 (I572924,I573010,I573168);
not I_33569 (I573213,I573168);
nand I_33570 (I572927,I573010,I573213);
nor I_33571 (I572921,I572976,I573168);
not I_33572 (I573258,I393560);
nor I_33573 (I573275,I573258,I393551);
nand I_33574 (I573292,I573275,I573117);
nor I_33575 (I572930,I573035,I573292);
nor I_33576 (I573323,I573258,I393569);
and I_33577 (I573340,I573323,I393557);
or I_33578 (I573357,I573340,I393572);
DFFARX1 I_33579 (I573357,I2507,I572950,I573383,);
nor I_33580 (I573391,I573383,I573134);
DFFARX1 I_33581 (I573391,I2507,I572950,I572918,);
DFFARX1 I_33582 (I573383,I2507,I572950,I572942,);
not I_33583 (I573436,I573383);
nor I_33584 (I573453,I573436,I573010);
nor I_33585 (I573470,I573275,I573453);
DFFARX1 I_33586 (I573470,I2507,I572950,I572939,);
not I_33587 (I573528,I2514);
DFFARX1 I_33588 (I84396,I2507,I573528,I573554,);
not I_33589 (I573562,I573554);
DFFARX1 I_33590 (I84375,I2507,I573528,I573588,);
not I_33591 (I573596,I84372);
nand I_33592 (I573613,I573596,I84387);
not I_33593 (I573630,I573613);
nor I_33594 (I573647,I573630,I84375);
nor I_33595 (I573664,I573562,I573647);
DFFARX1 I_33596 (I573664,I2507,I573528,I573514,);
not I_33597 (I573695,I84375);
nand I_33598 (I573712,I573695,I573630);
and I_33599 (I573729,I573695,I84378);
nand I_33600 (I573746,I573729,I84393);
nor I_33601 (I573511,I573746,I573695);
and I_33602 (I573502,I573588,I573746);
not I_33603 (I573791,I573746);
nand I_33604 (I573505,I573588,I573791);
nor I_33605 (I573499,I573554,I573746);
not I_33606 (I573836,I84384);
nor I_33607 (I573853,I573836,I84378);
nand I_33608 (I573870,I573853,I573695);
nor I_33609 (I573508,I573613,I573870);
nor I_33610 (I573901,I573836,I84372);
and I_33611 (I573918,I573901,I84381);
or I_33612 (I573935,I573918,I84390);
DFFARX1 I_33613 (I573935,I2507,I573528,I573961,);
nor I_33614 (I573969,I573961,I573712);
DFFARX1 I_33615 (I573969,I2507,I573528,I573496,);
DFFARX1 I_33616 (I573961,I2507,I573528,I573520,);
not I_33617 (I574014,I573961);
nor I_33618 (I574031,I574014,I573588);
nor I_33619 (I574048,I573853,I574031);
DFFARX1 I_33620 (I574048,I2507,I573528,I573517,);
not I_33621 (I574106,I2514);
DFFARX1 I_33622 (I1387422,I2507,I574106,I574132,);
not I_33623 (I574140,I574132);
DFFARX1 I_33624 (I1387422,I2507,I574106,I574166,);
not I_33625 (I574174,I1387446);
nand I_33626 (I574191,I574174,I1387428);
not I_33627 (I574208,I574191);
nor I_33628 (I574225,I574208,I1387443);
nor I_33629 (I574242,I574140,I574225);
DFFARX1 I_33630 (I574242,I2507,I574106,I574092,);
not I_33631 (I574273,I1387443);
nand I_33632 (I574290,I574273,I574208);
and I_33633 (I574307,I574273,I1387425);
nand I_33634 (I574324,I574307,I1387434);
nor I_33635 (I574089,I574324,I574273);
and I_33636 (I574080,I574166,I574324);
not I_33637 (I574369,I574324);
nand I_33638 (I574083,I574166,I574369);
nor I_33639 (I574077,I574132,I574324);
not I_33640 (I574414,I1387431);
nor I_33641 (I574431,I574414,I1387425);
nand I_33642 (I574448,I574431,I574273);
nor I_33643 (I574086,I574191,I574448);
nor I_33644 (I574479,I574414,I1387440);
and I_33645 (I574496,I574479,I1387449);
or I_33646 (I574513,I574496,I1387437);
DFFARX1 I_33647 (I574513,I2507,I574106,I574539,);
nor I_33648 (I574547,I574539,I574290);
DFFARX1 I_33649 (I574547,I2507,I574106,I574074,);
DFFARX1 I_33650 (I574539,I2507,I574106,I574098,);
not I_33651 (I574592,I574539);
nor I_33652 (I574609,I574592,I574166);
nor I_33653 (I574626,I574431,I574609);
DFFARX1 I_33654 (I574626,I2507,I574106,I574095,);
not I_33655 (I574684,I2514);
DFFARX1 I_33656 (I1091316,I2507,I574684,I574710,);
not I_33657 (I574718,I574710);
DFFARX1 I_33658 (I1091322,I2507,I574684,I574744,);
not I_33659 (I574752,I1091316);
nand I_33660 (I574769,I574752,I1091319);
not I_33661 (I574786,I574769);
nor I_33662 (I574803,I574786,I1091337);
nor I_33663 (I574820,I574718,I574803);
DFFARX1 I_33664 (I574820,I2507,I574684,I574670,);
not I_33665 (I574851,I1091337);
nand I_33666 (I574868,I574851,I574786);
and I_33667 (I574885,I574851,I1091340);
nand I_33668 (I574902,I574885,I1091319);
nor I_33669 (I574667,I574902,I574851);
and I_33670 (I574658,I574744,I574902);
not I_33671 (I574947,I574902);
nand I_33672 (I574661,I574744,I574947);
nor I_33673 (I574655,I574710,I574902);
not I_33674 (I574992,I1091325);
nor I_33675 (I575009,I574992,I1091340);
nand I_33676 (I575026,I575009,I574851);
nor I_33677 (I574664,I574769,I575026);
nor I_33678 (I575057,I574992,I1091331);
and I_33679 (I575074,I575057,I1091328);
or I_33680 (I575091,I575074,I1091334);
DFFARX1 I_33681 (I575091,I2507,I574684,I575117,);
nor I_33682 (I575125,I575117,I574868);
DFFARX1 I_33683 (I575125,I2507,I574684,I574652,);
DFFARX1 I_33684 (I575117,I2507,I574684,I574676,);
not I_33685 (I575170,I575117);
nor I_33686 (I575187,I575170,I574744);
nor I_33687 (I575204,I575009,I575187);
DFFARX1 I_33688 (I575204,I2507,I574684,I574673,);
not I_33689 (I575262,I2514);
DFFARX1 I_33690 (I23243,I2507,I575262,I575288,);
not I_33691 (I575296,I575288);
DFFARX1 I_33692 (I23246,I2507,I575262,I575322,);
not I_33693 (I575330,I23240);
nand I_33694 (I575347,I575330,I23264);
not I_33695 (I575364,I575347);
nor I_33696 (I575381,I575364,I23243);
nor I_33697 (I575398,I575296,I575381);
DFFARX1 I_33698 (I575398,I2507,I575262,I575248,);
not I_33699 (I575429,I23243);
nand I_33700 (I575446,I575429,I575364);
and I_33701 (I575463,I575429,I23258);
nand I_33702 (I575480,I575463,I23252);
nor I_33703 (I575245,I575480,I575429);
and I_33704 (I575236,I575322,I575480);
not I_33705 (I575525,I575480);
nand I_33706 (I575239,I575322,I575525);
nor I_33707 (I575233,I575288,I575480);
not I_33708 (I575570,I23261);
nor I_33709 (I575587,I575570,I23258);
nand I_33710 (I575604,I575587,I575429);
nor I_33711 (I575242,I575347,I575604);
nor I_33712 (I575635,I575570,I23240);
and I_33713 (I575652,I575635,I23249);
or I_33714 (I575669,I575652,I23255);
DFFARX1 I_33715 (I575669,I2507,I575262,I575695,);
nor I_33716 (I575703,I575695,I575446);
DFFARX1 I_33717 (I575703,I2507,I575262,I575230,);
DFFARX1 I_33718 (I575695,I2507,I575262,I575254,);
not I_33719 (I575748,I575695);
nor I_33720 (I575765,I575748,I575322);
nor I_33721 (I575782,I575587,I575765);
DFFARX1 I_33722 (I575782,I2507,I575262,I575251,);
not I_33723 (I575840,I2514);
DFFARX1 I_33724 (I1205760,I2507,I575840,I575866,);
not I_33725 (I575874,I575866);
DFFARX1 I_33726 (I1205766,I2507,I575840,I575900,);
not I_33727 (I575908,I1205760);
nand I_33728 (I575925,I575908,I1205763);
not I_33729 (I575942,I575925);
nor I_33730 (I575959,I575942,I1205781);
nor I_33731 (I575976,I575874,I575959);
DFFARX1 I_33732 (I575976,I2507,I575840,I575826,);
not I_33733 (I576007,I1205781);
nand I_33734 (I576024,I576007,I575942);
and I_33735 (I576041,I576007,I1205784);
nand I_33736 (I576058,I576041,I1205763);
nor I_33737 (I575823,I576058,I576007);
and I_33738 (I575814,I575900,I576058);
not I_33739 (I576103,I576058);
nand I_33740 (I575817,I575900,I576103);
nor I_33741 (I575811,I575866,I576058);
not I_33742 (I576148,I1205769);
nor I_33743 (I576165,I576148,I1205784);
nand I_33744 (I576182,I576165,I576007);
nor I_33745 (I575820,I575925,I576182);
nor I_33746 (I576213,I576148,I1205775);
and I_33747 (I576230,I576213,I1205772);
or I_33748 (I576247,I576230,I1205778);
DFFARX1 I_33749 (I576247,I2507,I575840,I576273,);
nor I_33750 (I576281,I576273,I576024);
DFFARX1 I_33751 (I576281,I2507,I575840,I575808,);
DFFARX1 I_33752 (I576273,I2507,I575840,I575832,);
not I_33753 (I576326,I576273);
nor I_33754 (I576343,I576326,I575900);
nor I_33755 (I576360,I576165,I576343);
DFFARX1 I_33756 (I576360,I2507,I575840,I575829,);
not I_33757 (I576418,I2514);
DFFARX1 I_33758 (I286559,I2507,I576418,I576444,);
not I_33759 (I576452,I576444);
DFFARX1 I_33760 (I286574,I2507,I576418,I576478,);
not I_33761 (I576486,I286577);
nand I_33762 (I576503,I576486,I286556);
not I_33763 (I576520,I576503);
nor I_33764 (I576537,I576520,I286580);
nor I_33765 (I576554,I576452,I576537);
DFFARX1 I_33766 (I576554,I2507,I576418,I576404,);
not I_33767 (I576585,I286580);
nand I_33768 (I576602,I576585,I576520);
and I_33769 (I576619,I576585,I286562);
nand I_33770 (I576636,I576619,I286553);
nor I_33771 (I576401,I576636,I576585);
and I_33772 (I576392,I576478,I576636);
not I_33773 (I576681,I576636);
nand I_33774 (I576395,I576478,I576681);
nor I_33775 (I576389,I576444,I576636);
not I_33776 (I576726,I286553);
nor I_33777 (I576743,I576726,I286562);
nand I_33778 (I576760,I576743,I576585);
nor I_33779 (I576398,I576503,I576760);
nor I_33780 (I576791,I576726,I286568);
and I_33781 (I576808,I576791,I286571);
or I_33782 (I576825,I576808,I286565);
DFFARX1 I_33783 (I576825,I2507,I576418,I576851,);
nor I_33784 (I576859,I576851,I576602);
DFFARX1 I_33785 (I576859,I2507,I576418,I576386,);
DFFARX1 I_33786 (I576851,I2507,I576418,I576410,);
not I_33787 (I576904,I576851);
nor I_33788 (I576921,I576904,I576478);
nor I_33789 (I576938,I576743,I576921);
DFFARX1 I_33790 (I576938,I2507,I576418,I576407,);
not I_33791 (I576996,I2514);
DFFARX1 I_33792 (I7884,I2507,I576996,I577022,);
not I_33793 (I577030,I577022);
DFFARX1 I_33794 (I7872,I2507,I576996,I577056,);
not I_33795 (I577064,I7881);
nand I_33796 (I577081,I577064,I7878);
not I_33797 (I577098,I577081);
nor I_33798 (I577115,I577098,I7887);
nor I_33799 (I577132,I577030,I577115);
DFFARX1 I_33800 (I577132,I2507,I576996,I576982,);
not I_33801 (I577163,I7887);
nand I_33802 (I577180,I577163,I577098);
and I_33803 (I577197,I577163,I7875);
nand I_33804 (I577214,I577197,I7878);
nor I_33805 (I576979,I577214,I577163);
and I_33806 (I576970,I577056,I577214);
not I_33807 (I577259,I577214);
nand I_33808 (I576973,I577056,I577259);
nor I_33809 (I576967,I577022,I577214);
not I_33810 (I577304,I7893);
nor I_33811 (I577321,I577304,I7875);
nand I_33812 (I577338,I577321,I577163);
nor I_33813 (I576976,I577081,I577338);
nor I_33814 (I577369,I577304,I7875);
and I_33815 (I577386,I577369,I7890);
or I_33816 (I577403,I577386,I7872);
DFFARX1 I_33817 (I577403,I2507,I576996,I577429,);
nor I_33818 (I577437,I577429,I577180);
DFFARX1 I_33819 (I577437,I2507,I576996,I576964,);
DFFARX1 I_33820 (I577429,I2507,I576996,I576988,);
not I_33821 (I577482,I577429);
nor I_33822 (I577499,I577482,I577056);
nor I_33823 (I577516,I577321,I577499);
DFFARX1 I_33824 (I577516,I2507,I576996,I576985,);
not I_33825 (I577574,I2514);
DFFARX1 I_33826 (I200225,I2507,I577574,I577600,);
not I_33827 (I577608,I577600);
DFFARX1 I_33828 (I200210,I2507,I577574,I577634,);
not I_33829 (I577642,I200228);
nand I_33830 (I577659,I577642,I200213);
not I_33831 (I577676,I577659);
nor I_33832 (I577693,I577676,I200210);
nor I_33833 (I577710,I577608,I577693);
DFFARX1 I_33834 (I577710,I2507,I577574,I577560,);
not I_33835 (I577741,I200210);
nand I_33836 (I577758,I577741,I577676);
and I_33837 (I577775,I577741,I200213);
nand I_33838 (I577792,I577775,I200234);
nor I_33839 (I577557,I577792,I577741);
and I_33840 (I577548,I577634,I577792);
not I_33841 (I577837,I577792);
nand I_33842 (I577551,I577634,I577837);
nor I_33843 (I577545,I577600,I577792);
not I_33844 (I577882,I200222);
nor I_33845 (I577899,I577882,I200213);
nand I_33846 (I577916,I577899,I577741);
nor I_33847 (I577554,I577659,I577916);
nor I_33848 (I577947,I577882,I200216);
and I_33849 (I577964,I577947,I200231);
or I_33850 (I577981,I577964,I200219);
DFFARX1 I_33851 (I577981,I2507,I577574,I578007,);
nor I_33852 (I578015,I578007,I577758);
DFFARX1 I_33853 (I578015,I2507,I577574,I577542,);
DFFARX1 I_33854 (I578007,I2507,I577574,I577566,);
not I_33855 (I578060,I578007);
nor I_33856 (I578077,I578060,I577634);
nor I_33857 (I578094,I577899,I578077);
DFFARX1 I_33858 (I578094,I2507,I577574,I577563,);
not I_33859 (I578152,I2514);
DFFARX1 I_33860 (I1200558,I2507,I578152,I578178,);
not I_33861 (I578186,I578178);
DFFARX1 I_33862 (I1200564,I2507,I578152,I578212,);
not I_33863 (I578220,I1200558);
nand I_33864 (I578237,I578220,I1200561);
not I_33865 (I578254,I578237);
nor I_33866 (I578271,I578254,I1200579);
nor I_33867 (I578288,I578186,I578271);
DFFARX1 I_33868 (I578288,I2507,I578152,I578138,);
not I_33869 (I578319,I1200579);
nand I_33870 (I578336,I578319,I578254);
and I_33871 (I578353,I578319,I1200582);
nand I_33872 (I578370,I578353,I1200561);
nor I_33873 (I578135,I578370,I578319);
and I_33874 (I578126,I578212,I578370);
not I_33875 (I578415,I578370);
nand I_33876 (I578129,I578212,I578415);
nor I_33877 (I578123,I578178,I578370);
not I_33878 (I578460,I1200567);
nor I_33879 (I578477,I578460,I1200582);
nand I_33880 (I578494,I578477,I578319);
nor I_33881 (I578132,I578237,I578494);
nor I_33882 (I578525,I578460,I1200573);
and I_33883 (I578542,I578525,I1200570);
or I_33884 (I578559,I578542,I1200576);
DFFARX1 I_33885 (I578559,I2507,I578152,I578585,);
nor I_33886 (I578593,I578585,I578336);
DFFARX1 I_33887 (I578593,I2507,I578152,I578120,);
DFFARX1 I_33888 (I578585,I2507,I578152,I578144,);
not I_33889 (I578638,I578585);
nor I_33890 (I578655,I578638,I578212);
nor I_33891 (I578672,I578477,I578655);
DFFARX1 I_33892 (I578672,I2507,I578152,I578141,);
not I_33893 (I578730,I2514);
DFFARX1 I_33894 (I653260,I2507,I578730,I578756,);
not I_33895 (I578764,I578756);
DFFARX1 I_33896 (I653272,I2507,I578730,I578790,);
not I_33897 (I578798,I653263);
nand I_33898 (I578815,I578798,I653266);
not I_33899 (I578832,I578815);
nor I_33900 (I578849,I578832,I653269);
nor I_33901 (I578866,I578764,I578849);
DFFARX1 I_33902 (I578866,I2507,I578730,I578716,);
not I_33903 (I578897,I653269);
nand I_33904 (I578914,I578897,I578832);
and I_33905 (I578931,I578897,I653263);
nand I_33906 (I578948,I578931,I653275);
nor I_33907 (I578713,I578948,I578897);
and I_33908 (I578704,I578790,I578948);
not I_33909 (I578993,I578948);
nand I_33910 (I578707,I578790,I578993);
nor I_33911 (I578701,I578756,I578948);
not I_33912 (I579038,I653281);
nor I_33913 (I579055,I579038,I653263);
nand I_33914 (I579072,I579055,I578897);
nor I_33915 (I578710,I578815,I579072);
nor I_33916 (I579103,I579038,I653260);
and I_33917 (I579120,I579103,I653278);
or I_33918 (I579137,I579120,I653284);
DFFARX1 I_33919 (I579137,I2507,I578730,I579163,);
nor I_33920 (I579171,I579163,I578914);
DFFARX1 I_33921 (I579171,I2507,I578730,I578698,);
DFFARX1 I_33922 (I579163,I2507,I578730,I578722,);
not I_33923 (I579216,I579163);
nor I_33924 (I579233,I579216,I578790);
nor I_33925 (I579250,I579055,I579233);
DFFARX1 I_33926 (I579250,I2507,I578730,I578719,);
not I_33927 (I579308,I2514);
DFFARX1 I_33928 (I121813,I2507,I579308,I579334,);
not I_33929 (I579342,I579334);
DFFARX1 I_33930 (I121792,I2507,I579308,I579368,);
not I_33931 (I579376,I121789);
nand I_33932 (I579393,I579376,I121804);
not I_33933 (I579410,I579393);
nor I_33934 (I579427,I579410,I121792);
nor I_33935 (I579444,I579342,I579427);
DFFARX1 I_33936 (I579444,I2507,I579308,I579294,);
not I_33937 (I579475,I121792);
nand I_33938 (I579492,I579475,I579410);
and I_33939 (I579509,I579475,I121795);
nand I_33940 (I579526,I579509,I121810);
nor I_33941 (I579291,I579526,I579475);
and I_33942 (I579282,I579368,I579526);
not I_33943 (I579571,I579526);
nand I_33944 (I579285,I579368,I579571);
nor I_33945 (I579279,I579334,I579526);
not I_33946 (I579616,I121801);
nor I_33947 (I579633,I579616,I121795);
nand I_33948 (I579650,I579633,I579475);
nor I_33949 (I579288,I579393,I579650);
nor I_33950 (I579681,I579616,I121789);
and I_33951 (I579698,I579681,I121798);
or I_33952 (I579715,I579698,I121807);
DFFARX1 I_33953 (I579715,I2507,I579308,I579741,);
nor I_33954 (I579749,I579741,I579492);
DFFARX1 I_33955 (I579749,I2507,I579308,I579276,);
DFFARX1 I_33956 (I579741,I2507,I579308,I579300,);
not I_33957 (I579794,I579741);
nor I_33958 (I579811,I579794,I579368);
nor I_33959 (I579828,I579633,I579811);
DFFARX1 I_33960 (I579828,I2507,I579308,I579297,);
not I_33961 (I579886,I2514);
DFFARX1 I_33962 (I475707,I2507,I579886,I579912,);
not I_33963 (I579920,I579912);
DFFARX1 I_33964 (I475719,I2507,I579886,I579946,);
not I_33965 (I579954,I475695);
nand I_33966 (I579971,I579954,I475722);
not I_33967 (I579988,I579971);
nor I_33968 (I580005,I579988,I475710);
nor I_33969 (I580022,I579920,I580005);
DFFARX1 I_33970 (I580022,I2507,I579886,I579872,);
not I_33971 (I580053,I475710);
nand I_33972 (I580070,I580053,I579988);
and I_33973 (I580087,I580053,I475695);
nand I_33974 (I580104,I580087,I475698);
nor I_33975 (I579869,I580104,I580053);
and I_33976 (I579860,I579946,I580104);
not I_33977 (I580149,I580104);
nand I_33978 (I579863,I579946,I580149);
nor I_33979 (I579857,I579912,I580104);
not I_33980 (I580194,I475704);
nor I_33981 (I580211,I580194,I475695);
nand I_33982 (I580228,I580211,I580053);
nor I_33983 (I579866,I579971,I580228);
nor I_33984 (I580259,I580194,I475713);
and I_33985 (I580276,I580259,I475701);
or I_33986 (I580293,I580276,I475716);
DFFARX1 I_33987 (I580293,I2507,I579886,I580319,);
nor I_33988 (I580327,I580319,I580070);
DFFARX1 I_33989 (I580327,I2507,I579886,I579854,);
DFFARX1 I_33990 (I580319,I2507,I579886,I579878,);
not I_33991 (I580372,I580319);
nor I_33992 (I580389,I580372,I579946);
nor I_33993 (I580406,I580211,I580389);
DFFARX1 I_33994 (I580406,I2507,I579886,I579875,);
not I_33995 (I580464,I2514);
DFFARX1 I_33996 (I147276,I2507,I580464,I580490,);
not I_33997 (I580498,I580490);
DFFARX1 I_33998 (I147255,I2507,I580464,I580524,);
not I_33999 (I580532,I147255);
nand I_34000 (I580549,I580532,I147282);
not I_34001 (I580566,I580549);
nor I_34002 (I580583,I580566,I147258);
nor I_34003 (I580600,I580498,I580583);
DFFARX1 I_34004 (I580600,I2507,I580464,I580450,);
not I_34005 (I580631,I147258);
nand I_34006 (I580648,I580631,I580566);
and I_34007 (I580665,I580631,I147279);
nand I_34008 (I580682,I580665,I147261);
nor I_34009 (I580447,I580682,I580631);
and I_34010 (I580438,I580524,I580682);
not I_34011 (I580727,I580682);
nand I_34012 (I580441,I580524,I580727);
nor I_34013 (I580435,I580490,I580682);
not I_34014 (I580772,I147264);
nor I_34015 (I580789,I580772,I147279);
nand I_34016 (I580806,I580789,I580631);
nor I_34017 (I580444,I580549,I580806);
nor I_34018 (I580837,I580772,I147270);
and I_34019 (I580854,I580837,I147267);
or I_34020 (I580871,I580854,I147273);
DFFARX1 I_34021 (I580871,I2507,I580464,I580897,);
nor I_34022 (I580905,I580897,I580648);
DFFARX1 I_34023 (I580905,I2507,I580464,I580432,);
DFFARX1 I_34024 (I580897,I2507,I580464,I580456,);
not I_34025 (I580950,I580897);
nor I_34026 (I580967,I580950,I580524);
nor I_34027 (I580984,I580789,I580967);
DFFARX1 I_34028 (I580984,I2507,I580464,I580453,);
not I_34029 (I581042,I2514);
DFFARX1 I_34030 (I160360,I2507,I581042,I581068,);
not I_34031 (I581076,I581068);
DFFARX1 I_34032 (I160345,I2507,I581042,I581102,);
not I_34033 (I581110,I160363);
nand I_34034 (I581127,I581110,I160348);
not I_34035 (I581144,I581127);
nor I_34036 (I581161,I581144,I160345);
nor I_34037 (I581178,I581076,I581161);
DFFARX1 I_34038 (I581178,I2507,I581042,I581028,);
not I_34039 (I581209,I160345);
nand I_34040 (I581226,I581209,I581144);
and I_34041 (I581243,I581209,I160348);
nand I_34042 (I581260,I581243,I160369);
nor I_34043 (I581025,I581260,I581209);
and I_34044 (I581016,I581102,I581260);
not I_34045 (I581305,I581260);
nand I_34046 (I581019,I581102,I581305);
nor I_34047 (I581013,I581068,I581260);
not I_34048 (I581350,I160357);
nor I_34049 (I581367,I581350,I160348);
nand I_34050 (I581384,I581367,I581209);
nor I_34051 (I581022,I581127,I581384);
nor I_34052 (I581415,I581350,I160351);
and I_34053 (I581432,I581415,I160366);
or I_34054 (I581449,I581432,I160354);
DFFARX1 I_34055 (I581449,I2507,I581042,I581475,);
nor I_34056 (I581483,I581475,I581226);
DFFARX1 I_34057 (I581483,I2507,I581042,I581010,);
DFFARX1 I_34058 (I581475,I2507,I581042,I581034,);
not I_34059 (I581528,I581475);
nor I_34060 (I581545,I581528,I581102);
nor I_34061 (I581562,I581367,I581545);
DFFARX1 I_34062 (I581562,I2507,I581042,I581031,);
not I_34063 (I581620,I2514);
DFFARX1 I_34064 (I1371952,I2507,I581620,I581646,);
not I_34065 (I581654,I581646);
DFFARX1 I_34066 (I1371952,I2507,I581620,I581680,);
not I_34067 (I581688,I1371976);
nand I_34068 (I581705,I581688,I1371958);
not I_34069 (I581722,I581705);
nor I_34070 (I581739,I581722,I1371973);
nor I_34071 (I581756,I581654,I581739);
DFFARX1 I_34072 (I581756,I2507,I581620,I581606,);
not I_34073 (I581787,I1371973);
nand I_34074 (I581804,I581787,I581722);
and I_34075 (I581821,I581787,I1371955);
nand I_34076 (I581838,I581821,I1371964);
nor I_34077 (I581603,I581838,I581787);
and I_34078 (I581594,I581680,I581838);
not I_34079 (I581883,I581838);
nand I_34080 (I581597,I581680,I581883);
nor I_34081 (I581591,I581646,I581838);
not I_34082 (I581928,I1371961);
nor I_34083 (I581945,I581928,I1371955);
nand I_34084 (I581962,I581945,I581787);
nor I_34085 (I581600,I581705,I581962);
nor I_34086 (I581993,I581928,I1371970);
and I_34087 (I582010,I581993,I1371979);
or I_34088 (I582027,I582010,I1371967);
DFFARX1 I_34089 (I582027,I2507,I581620,I582053,);
nor I_34090 (I582061,I582053,I581804);
DFFARX1 I_34091 (I582061,I2507,I581620,I581588,);
DFFARX1 I_34092 (I582053,I2507,I581620,I581612,);
not I_34093 (I582106,I582053);
nor I_34094 (I582123,I582106,I581680);
nor I_34095 (I582140,I581945,I582123);
DFFARX1 I_34096 (I582140,I2507,I581620,I581609,);
not I_34097 (I582198,I2514);
DFFARX1 I_34098 (I242470,I2507,I582198,I582224,);
not I_34099 (I582232,I582224);
DFFARX1 I_34100 (I242455,I2507,I582198,I582258,);
not I_34101 (I582266,I242473);
nand I_34102 (I582283,I582266,I242458);
not I_34103 (I582300,I582283);
nor I_34104 (I582317,I582300,I242455);
nor I_34105 (I582334,I582232,I582317);
DFFARX1 I_34106 (I582334,I2507,I582198,I582184,);
not I_34107 (I582365,I242455);
nand I_34108 (I582382,I582365,I582300);
and I_34109 (I582399,I582365,I242458);
nand I_34110 (I582416,I582399,I242479);
nor I_34111 (I582181,I582416,I582365);
and I_34112 (I582172,I582258,I582416);
not I_34113 (I582461,I582416);
nand I_34114 (I582175,I582258,I582461);
nor I_34115 (I582169,I582224,I582416);
not I_34116 (I582506,I242467);
nor I_34117 (I582523,I582506,I242458);
nand I_34118 (I582540,I582523,I582365);
nor I_34119 (I582178,I582283,I582540);
nor I_34120 (I582571,I582506,I242461);
and I_34121 (I582588,I582571,I242476);
or I_34122 (I582605,I582588,I242464);
DFFARX1 I_34123 (I582605,I2507,I582198,I582631,);
nor I_34124 (I582639,I582631,I582382);
DFFARX1 I_34125 (I582639,I2507,I582198,I582166,);
DFFARX1 I_34126 (I582631,I2507,I582198,I582190,);
not I_34127 (I582684,I582631);
nor I_34128 (I582701,I582684,I582258);
nor I_34129 (I582718,I582523,I582701);
DFFARX1 I_34130 (I582718,I2507,I582198,I582187,);
not I_34131 (I582776,I2514);
DFFARX1 I_34132 (I694876,I2507,I582776,I582802,);
not I_34133 (I582810,I582802);
DFFARX1 I_34134 (I694888,I2507,I582776,I582836,);
not I_34135 (I582844,I694879);
nand I_34136 (I582861,I582844,I694882);
not I_34137 (I582878,I582861);
nor I_34138 (I582895,I582878,I694885);
nor I_34139 (I582912,I582810,I582895);
DFFARX1 I_34140 (I582912,I2507,I582776,I582762,);
not I_34141 (I582943,I694885);
nand I_34142 (I582960,I582943,I582878);
and I_34143 (I582977,I582943,I694879);
nand I_34144 (I582994,I582977,I694891);
nor I_34145 (I582759,I582994,I582943);
and I_34146 (I582750,I582836,I582994);
not I_34147 (I583039,I582994);
nand I_34148 (I582753,I582836,I583039);
nor I_34149 (I582747,I582802,I582994);
not I_34150 (I583084,I694897);
nor I_34151 (I583101,I583084,I694879);
nand I_34152 (I583118,I583101,I582943);
nor I_34153 (I582756,I582861,I583118);
nor I_34154 (I583149,I583084,I694876);
and I_34155 (I583166,I583149,I694894);
or I_34156 (I583183,I583166,I694900);
DFFARX1 I_34157 (I583183,I2507,I582776,I583209,);
nor I_34158 (I583217,I583209,I582960);
DFFARX1 I_34159 (I583217,I2507,I582776,I582744,);
DFFARX1 I_34160 (I583209,I2507,I582776,I582768,);
not I_34161 (I583262,I583209);
nor I_34162 (I583279,I583262,I582836);
nor I_34163 (I583296,I583101,I583279);
DFFARX1 I_34164 (I583296,I2507,I582776,I582765,);
not I_34165 (I583354,I2514);
DFFARX1 I_34166 (I492027,I2507,I583354,I583380,);
not I_34167 (I583388,I583380);
DFFARX1 I_34168 (I492039,I2507,I583354,I583414,);
not I_34169 (I583422,I492015);
nand I_34170 (I583439,I583422,I492042);
not I_34171 (I583456,I583439);
nor I_34172 (I583473,I583456,I492030);
nor I_34173 (I583490,I583388,I583473);
DFFARX1 I_34174 (I583490,I2507,I583354,I583340,);
not I_34175 (I583521,I492030);
nand I_34176 (I583538,I583521,I583456);
and I_34177 (I583555,I583521,I492015);
nand I_34178 (I583572,I583555,I492018);
nor I_34179 (I583337,I583572,I583521);
and I_34180 (I583328,I583414,I583572);
not I_34181 (I583617,I583572);
nand I_34182 (I583331,I583414,I583617);
nor I_34183 (I583325,I583380,I583572);
not I_34184 (I583662,I492024);
nor I_34185 (I583679,I583662,I492015);
nand I_34186 (I583696,I583679,I583521);
nor I_34187 (I583334,I583439,I583696);
nor I_34188 (I583727,I583662,I492033);
and I_34189 (I583744,I583727,I492021);
or I_34190 (I583761,I583744,I492036);
DFFARX1 I_34191 (I583761,I2507,I583354,I583787,);
nor I_34192 (I583795,I583787,I583538);
DFFARX1 I_34193 (I583795,I2507,I583354,I583322,);
DFFARX1 I_34194 (I583787,I2507,I583354,I583346,);
not I_34195 (I583840,I583787);
nor I_34196 (I583857,I583840,I583414);
nor I_34197 (I583874,I583679,I583857);
DFFARX1 I_34198 (I583874,I2507,I583354,I583343,);
not I_34199 (I583932,I2514);
DFFARX1 I_34200 (I984477,I2507,I583932,I583958,);
not I_34201 (I583966,I583958);
DFFARX1 I_34202 (I984474,I2507,I583932,I583992,);
not I_34203 (I584000,I984471);
nand I_34204 (I584017,I584000,I984498);
not I_34205 (I584034,I584017);
nor I_34206 (I584051,I584034,I984486);
nor I_34207 (I584068,I583966,I584051);
DFFARX1 I_34208 (I584068,I2507,I583932,I583918,);
not I_34209 (I584099,I984486);
nand I_34210 (I584116,I584099,I584034);
and I_34211 (I584133,I584099,I984492);
nand I_34212 (I584150,I584133,I984483);
nor I_34213 (I583915,I584150,I584099);
and I_34214 (I583906,I583992,I584150);
not I_34215 (I584195,I584150);
nand I_34216 (I583909,I583992,I584195);
nor I_34217 (I583903,I583958,I584150);
not I_34218 (I584240,I984480);
nor I_34219 (I584257,I584240,I984492);
nand I_34220 (I584274,I584257,I584099);
nor I_34221 (I583912,I584017,I584274);
nor I_34222 (I584305,I584240,I984495);
and I_34223 (I584322,I584305,I984489);
or I_34224 (I584339,I584322,I984471);
DFFARX1 I_34225 (I584339,I2507,I583932,I584365,);
nor I_34226 (I584373,I584365,I584116);
DFFARX1 I_34227 (I584373,I2507,I583932,I583900,);
DFFARX1 I_34228 (I584365,I2507,I583932,I583924,);
not I_34229 (I584418,I584365);
nor I_34230 (I584435,I584418,I583992);
nor I_34231 (I584452,I584257,I584435);
DFFARX1 I_34232 (I584452,I2507,I583932,I583921,);
not I_34233 (I584510,I2514);
DFFARX1 I_34234 (I397371,I2507,I584510,I584536,);
not I_34235 (I584544,I584536);
DFFARX1 I_34236 (I397383,I2507,I584510,I584570,);
not I_34237 (I584578,I397359);
nand I_34238 (I584595,I584578,I397386);
not I_34239 (I584612,I584595);
nor I_34240 (I584629,I584612,I397374);
nor I_34241 (I584646,I584544,I584629);
DFFARX1 I_34242 (I584646,I2507,I584510,I584496,);
not I_34243 (I584677,I397374);
nand I_34244 (I584694,I584677,I584612);
and I_34245 (I584711,I584677,I397359);
nand I_34246 (I584728,I584711,I397362);
nor I_34247 (I584493,I584728,I584677);
and I_34248 (I584484,I584570,I584728);
not I_34249 (I584773,I584728);
nand I_34250 (I584487,I584570,I584773);
nor I_34251 (I584481,I584536,I584728);
not I_34252 (I584818,I397368);
nor I_34253 (I584835,I584818,I397359);
nand I_34254 (I584852,I584835,I584677);
nor I_34255 (I584490,I584595,I584852);
nor I_34256 (I584883,I584818,I397377);
and I_34257 (I584900,I584883,I397365);
or I_34258 (I584917,I584900,I397380);
DFFARX1 I_34259 (I584917,I2507,I584510,I584943,);
nor I_34260 (I584951,I584943,I584694);
DFFARX1 I_34261 (I584951,I2507,I584510,I584478,);
DFFARX1 I_34262 (I584943,I2507,I584510,I584502,);
not I_34263 (I584996,I584943);
nor I_34264 (I585013,I584996,I584570);
nor I_34265 (I585030,I584835,I585013);
DFFARX1 I_34266 (I585030,I2507,I584510,I584499,);
not I_34267 (I585088,I2514);
DFFARX1 I_34268 (I166310,I2507,I585088,I585114,);
not I_34269 (I585122,I585114);
DFFARX1 I_34270 (I166295,I2507,I585088,I585148,);
not I_34271 (I585156,I166313);
nand I_34272 (I585173,I585156,I166298);
not I_34273 (I585190,I585173);
nor I_34274 (I585207,I585190,I166295);
nor I_34275 (I585224,I585122,I585207);
DFFARX1 I_34276 (I585224,I2507,I585088,I585074,);
not I_34277 (I585255,I166295);
nand I_34278 (I585272,I585255,I585190);
and I_34279 (I585289,I585255,I166298);
nand I_34280 (I585306,I585289,I166319);
nor I_34281 (I585071,I585306,I585255);
and I_34282 (I585062,I585148,I585306);
not I_34283 (I585351,I585306);
nand I_34284 (I585065,I585148,I585351);
nor I_34285 (I585059,I585114,I585306);
not I_34286 (I585396,I166307);
nor I_34287 (I585413,I585396,I166298);
nand I_34288 (I585430,I585413,I585255);
nor I_34289 (I585068,I585173,I585430);
nor I_34290 (I585461,I585396,I166301);
and I_34291 (I585478,I585461,I166316);
or I_34292 (I585495,I585478,I166304);
DFFARX1 I_34293 (I585495,I2507,I585088,I585521,);
nor I_34294 (I585529,I585521,I585272);
DFFARX1 I_34295 (I585529,I2507,I585088,I585056,);
DFFARX1 I_34296 (I585521,I2507,I585088,I585080,);
not I_34297 (I585574,I585521);
nor I_34298 (I585591,I585574,I585148);
nor I_34299 (I585608,I585413,I585591);
DFFARX1 I_34300 (I585608,I2507,I585088,I585077,);
not I_34301 (I585666,I2514);
DFFARX1 I_34302 (I811213,I2507,I585666,I585692,);
not I_34303 (I585700,I585692);
DFFARX1 I_34304 (I811213,I2507,I585666,I585726,);
not I_34305 (I585734,I811210);
nand I_34306 (I585751,I585734,I811225);
not I_34307 (I585768,I585751);
nor I_34308 (I585785,I585768,I811219);
nor I_34309 (I585802,I585700,I585785);
DFFARX1 I_34310 (I585802,I2507,I585666,I585652,);
not I_34311 (I585833,I811219);
nand I_34312 (I585850,I585833,I585768);
and I_34313 (I585867,I585833,I811216);
nand I_34314 (I585884,I585867,I811207);
nor I_34315 (I585649,I585884,I585833);
and I_34316 (I585640,I585726,I585884);
not I_34317 (I585929,I585884);
nand I_34318 (I585643,I585726,I585929);
nor I_34319 (I585637,I585692,I585884);
not I_34320 (I585974,I811228);
nor I_34321 (I585991,I585974,I811216);
nand I_34322 (I586008,I585991,I585833);
nor I_34323 (I585646,I585751,I586008);
nor I_34324 (I586039,I585974,I811207);
and I_34325 (I586056,I586039,I811210);
or I_34326 (I586073,I586056,I811222);
DFFARX1 I_34327 (I586073,I2507,I585666,I586099,);
nor I_34328 (I586107,I586099,I585850);
DFFARX1 I_34329 (I586107,I2507,I585666,I585634,);
DFFARX1 I_34330 (I586099,I2507,I585666,I585658,);
not I_34331 (I586152,I586099);
nor I_34332 (I586169,I586152,I585726);
nor I_34333 (I586186,I585991,I586169);
DFFARX1 I_34334 (I586186,I2507,I585666,I585655,);
not I_34335 (I586244,I2514);
DFFARX1 I_34336 (I783809,I2507,I586244,I586270,);
not I_34337 (I586278,I586270);
DFFARX1 I_34338 (I783809,I2507,I586244,I586304,);
not I_34339 (I586312,I783806);
nand I_34340 (I586329,I586312,I783821);
not I_34341 (I586346,I586329);
nor I_34342 (I586363,I586346,I783815);
nor I_34343 (I586380,I586278,I586363);
DFFARX1 I_34344 (I586380,I2507,I586244,I586230,);
not I_34345 (I586411,I783815);
nand I_34346 (I586428,I586411,I586346);
and I_34347 (I586445,I586411,I783812);
nand I_34348 (I586462,I586445,I783803);
nor I_34349 (I586227,I586462,I586411);
and I_34350 (I586218,I586304,I586462);
not I_34351 (I586507,I586462);
nand I_34352 (I586221,I586304,I586507);
nor I_34353 (I586215,I586270,I586462);
not I_34354 (I586552,I783824);
nor I_34355 (I586569,I586552,I783812);
nand I_34356 (I586586,I586569,I586411);
nor I_34357 (I586224,I586329,I586586);
nor I_34358 (I586617,I586552,I783803);
and I_34359 (I586634,I586617,I783806);
or I_34360 (I586651,I586634,I783818);
DFFARX1 I_34361 (I586651,I2507,I586244,I586677,);
nor I_34362 (I586685,I586677,I586428);
DFFARX1 I_34363 (I586685,I2507,I586244,I586212,);
DFFARX1 I_34364 (I586677,I2507,I586244,I586236,);
not I_34365 (I586730,I586677);
nor I_34366 (I586747,I586730,I586304);
nor I_34367 (I586764,I586569,I586747);
DFFARX1 I_34368 (I586764,I2507,I586244,I586233,);
not I_34369 (I586822,I2514);
DFFARX1 I_34370 (I1255922,I2507,I586822,I586848,);
not I_34371 (I586856,I586848);
DFFARX1 I_34372 (I1255934,I2507,I586822,I586882,);
not I_34373 (I586890,I1255925);
nand I_34374 (I586907,I586890,I1255913);
not I_34375 (I586924,I586907);
nor I_34376 (I586941,I586924,I1255910);
nor I_34377 (I586958,I586856,I586941);
DFFARX1 I_34378 (I586958,I2507,I586822,I586808,);
not I_34379 (I586989,I1255910);
nand I_34380 (I587006,I586989,I586924);
and I_34381 (I587023,I586989,I1255916);
nand I_34382 (I587040,I587023,I1255913);
nor I_34383 (I586805,I587040,I586989);
and I_34384 (I586796,I586882,I587040);
not I_34385 (I587085,I587040);
nand I_34386 (I586799,I586882,I587085);
nor I_34387 (I586793,I586848,I587040);
not I_34388 (I587130,I1255931);
nor I_34389 (I587147,I587130,I1255916);
nand I_34390 (I587164,I587147,I586989);
nor I_34391 (I586802,I586907,I587164);
nor I_34392 (I587195,I587130,I1255919);
and I_34393 (I587212,I587195,I1255910);
or I_34394 (I587229,I587212,I1255928);
DFFARX1 I_34395 (I587229,I2507,I586822,I587255,);
nor I_34396 (I587263,I587255,I587006);
DFFARX1 I_34397 (I587263,I2507,I586822,I586790,);
DFFARX1 I_34398 (I587255,I2507,I586822,I586814,);
not I_34399 (I587308,I587255);
nor I_34400 (I587325,I587308,I586882);
nor I_34401 (I587342,I587147,I587325);
DFFARX1 I_34402 (I587342,I2507,I586822,I586811,);
not I_34403 (I587400,I2514);
DFFARX1 I_34404 (I743428,I2507,I587400,I587426,);
not I_34405 (I587434,I587426);
DFFARX1 I_34406 (I743440,I2507,I587400,I587460,);
not I_34407 (I587468,I743431);
nand I_34408 (I587485,I587468,I743434);
not I_34409 (I587502,I587485);
nor I_34410 (I587519,I587502,I743437);
nor I_34411 (I587536,I587434,I587519);
DFFARX1 I_34412 (I587536,I2507,I587400,I587386,);
not I_34413 (I587567,I743437);
nand I_34414 (I587584,I587567,I587502);
and I_34415 (I587601,I587567,I743431);
nand I_34416 (I587618,I587601,I743443);
nor I_34417 (I587383,I587618,I587567);
and I_34418 (I587374,I587460,I587618);
not I_34419 (I587663,I587618);
nand I_34420 (I587377,I587460,I587663);
nor I_34421 (I587371,I587426,I587618);
not I_34422 (I587708,I743449);
nor I_34423 (I587725,I587708,I743431);
nand I_34424 (I587742,I587725,I587567);
nor I_34425 (I587380,I587485,I587742);
nor I_34426 (I587773,I587708,I743428);
and I_34427 (I587790,I587773,I743446);
or I_34428 (I587807,I587790,I743452);
DFFARX1 I_34429 (I587807,I2507,I587400,I587833,);
nor I_34430 (I587841,I587833,I587584);
DFFARX1 I_34431 (I587841,I2507,I587400,I587368,);
DFFARX1 I_34432 (I587833,I2507,I587400,I587392,);
not I_34433 (I587886,I587833);
nor I_34434 (I587903,I587886,I587460);
nor I_34435 (I587920,I587725,I587903);
DFFARX1 I_34436 (I587920,I2507,I587400,I587389,);
not I_34437 (I587978,I2514);
DFFARX1 I_34438 (I79126,I2507,I587978,I588004,);
not I_34439 (I588012,I588004);
DFFARX1 I_34440 (I79105,I2507,I587978,I588038,);
not I_34441 (I588046,I79102);
nand I_34442 (I588063,I588046,I79117);
not I_34443 (I588080,I588063);
nor I_34444 (I588097,I588080,I79105);
nor I_34445 (I588114,I588012,I588097);
DFFARX1 I_34446 (I588114,I2507,I587978,I587964,);
not I_34447 (I588145,I79105);
nand I_34448 (I588162,I588145,I588080);
and I_34449 (I588179,I588145,I79108);
nand I_34450 (I588196,I588179,I79123);
nor I_34451 (I587961,I588196,I588145);
and I_34452 (I587952,I588038,I588196);
not I_34453 (I588241,I588196);
nand I_34454 (I587955,I588038,I588241);
nor I_34455 (I587949,I588004,I588196);
not I_34456 (I588286,I79114);
nor I_34457 (I588303,I588286,I79108);
nand I_34458 (I588320,I588303,I588145);
nor I_34459 (I587958,I588063,I588320);
nor I_34460 (I588351,I588286,I79102);
and I_34461 (I588368,I588351,I79111);
or I_34462 (I588385,I588368,I79120);
DFFARX1 I_34463 (I588385,I2507,I587978,I588411,);
nor I_34464 (I588419,I588411,I588162);
DFFARX1 I_34465 (I588419,I2507,I587978,I587946,);
DFFARX1 I_34466 (I588411,I2507,I587978,I587970,);
not I_34467 (I588464,I588411);
nor I_34468 (I588481,I588464,I588038);
nor I_34469 (I588498,I588303,I588481);
DFFARX1 I_34470 (I588498,I2507,I587978,I587967,);
not I_34471 (I588556,I2514);
DFFARX1 I_34472 (I1128886,I2507,I588556,I588582,);
not I_34473 (I588590,I588582);
DFFARX1 I_34474 (I1128892,I2507,I588556,I588616,);
not I_34475 (I588624,I1128886);
nand I_34476 (I588641,I588624,I1128889);
not I_34477 (I588658,I588641);
nor I_34478 (I588675,I588658,I1128907);
nor I_34479 (I588692,I588590,I588675);
DFFARX1 I_34480 (I588692,I2507,I588556,I588542,);
not I_34481 (I588723,I1128907);
nand I_34482 (I588740,I588723,I588658);
and I_34483 (I588757,I588723,I1128910);
nand I_34484 (I588774,I588757,I1128889);
nor I_34485 (I588539,I588774,I588723);
and I_34486 (I588530,I588616,I588774);
not I_34487 (I588819,I588774);
nand I_34488 (I588533,I588616,I588819);
nor I_34489 (I588527,I588582,I588774);
not I_34490 (I588864,I1128895);
nor I_34491 (I588881,I588864,I1128910);
nand I_34492 (I588898,I588881,I588723);
nor I_34493 (I588536,I588641,I588898);
nor I_34494 (I588929,I588864,I1128901);
and I_34495 (I588946,I588929,I1128898);
or I_34496 (I588963,I588946,I1128904);
DFFARX1 I_34497 (I588963,I2507,I588556,I588989,);
nor I_34498 (I588997,I588989,I588740);
DFFARX1 I_34499 (I588997,I2507,I588556,I588524,);
DFFARX1 I_34500 (I588989,I2507,I588556,I588548,);
not I_34501 (I589042,I588989);
nor I_34502 (I589059,I589042,I588616);
nor I_34503 (I589076,I588881,I589059);
DFFARX1 I_34504 (I589076,I2507,I588556,I588545,);
not I_34505 (I589134,I2514);
DFFARX1 I_34506 (I101787,I2507,I589134,I589160,);
not I_34507 (I589168,I589160);
DFFARX1 I_34508 (I101766,I2507,I589134,I589194,);
not I_34509 (I589202,I101763);
nand I_34510 (I589219,I589202,I101778);
not I_34511 (I589236,I589219);
nor I_34512 (I589253,I589236,I101766);
nor I_34513 (I589270,I589168,I589253);
DFFARX1 I_34514 (I589270,I2507,I589134,I589120,);
not I_34515 (I589301,I101766);
nand I_34516 (I589318,I589301,I589236);
and I_34517 (I589335,I589301,I101769);
nand I_34518 (I589352,I589335,I101784);
nor I_34519 (I589117,I589352,I589301);
and I_34520 (I589108,I589194,I589352);
not I_34521 (I589397,I589352);
nand I_34522 (I589111,I589194,I589397);
nor I_34523 (I589105,I589160,I589352);
not I_34524 (I589442,I101775);
nor I_34525 (I589459,I589442,I101769);
nand I_34526 (I589476,I589459,I589301);
nor I_34527 (I589114,I589219,I589476);
nor I_34528 (I589507,I589442,I101763);
and I_34529 (I589524,I589507,I101772);
or I_34530 (I589541,I589524,I101781);
DFFARX1 I_34531 (I589541,I2507,I589134,I589567,);
nor I_34532 (I589575,I589567,I589318);
DFFARX1 I_34533 (I589575,I2507,I589134,I589102,);
DFFARX1 I_34534 (I589567,I2507,I589134,I589126,);
not I_34535 (I589620,I589567);
nor I_34536 (I589637,I589620,I589194);
nor I_34537 (I589654,I589459,I589637);
DFFARX1 I_34538 (I589654,I2507,I589134,I589123,);
not I_34539 (I589712,I2514);
DFFARX1 I_34540 (I1378497,I2507,I589712,I589738,);
not I_34541 (I589746,I589738);
DFFARX1 I_34542 (I1378497,I2507,I589712,I589772,);
not I_34543 (I589780,I1378521);
nand I_34544 (I589797,I589780,I1378503);
not I_34545 (I589814,I589797);
nor I_34546 (I589831,I589814,I1378518);
nor I_34547 (I589848,I589746,I589831);
DFFARX1 I_34548 (I589848,I2507,I589712,I589698,);
not I_34549 (I589879,I1378518);
nand I_34550 (I589896,I589879,I589814);
and I_34551 (I589913,I589879,I1378500);
nand I_34552 (I589930,I589913,I1378509);
nor I_34553 (I589695,I589930,I589879);
and I_34554 (I589686,I589772,I589930);
not I_34555 (I589975,I589930);
nand I_34556 (I589689,I589772,I589975);
nor I_34557 (I589683,I589738,I589930);
not I_34558 (I590020,I1378506);
nor I_34559 (I590037,I590020,I1378500);
nand I_34560 (I590054,I590037,I589879);
nor I_34561 (I589692,I589797,I590054);
nor I_34562 (I590085,I590020,I1378515);
and I_34563 (I590102,I590085,I1378524);
or I_34564 (I590119,I590102,I1378512);
DFFARX1 I_34565 (I590119,I2507,I589712,I590145,);
nor I_34566 (I590153,I590145,I589896);
DFFARX1 I_34567 (I590153,I2507,I589712,I589680,);
DFFARX1 I_34568 (I590145,I2507,I589712,I589704,);
not I_34569 (I590198,I590145);
nor I_34570 (I590215,I590198,I589772);
nor I_34571 (I590232,I590037,I590215);
DFFARX1 I_34572 (I590232,I2507,I589712,I589701,);
not I_34573 (I590290,I2514);
DFFARX1 I_34574 (I1330897,I2507,I590290,I590316,);
not I_34575 (I590324,I590316);
DFFARX1 I_34576 (I1330897,I2507,I590290,I590350,);
not I_34577 (I590358,I1330921);
nand I_34578 (I590375,I590358,I1330903);
not I_34579 (I590392,I590375);
nor I_34580 (I590409,I590392,I1330918);
nor I_34581 (I590426,I590324,I590409);
DFFARX1 I_34582 (I590426,I2507,I590290,I590276,);
not I_34583 (I590457,I1330918);
nand I_34584 (I590474,I590457,I590392);
and I_34585 (I590491,I590457,I1330900);
nand I_34586 (I590508,I590491,I1330909);
nor I_34587 (I590273,I590508,I590457);
and I_34588 (I590264,I590350,I590508);
not I_34589 (I590553,I590508);
nand I_34590 (I590267,I590350,I590553);
nor I_34591 (I590261,I590316,I590508);
not I_34592 (I590598,I1330906);
nor I_34593 (I590615,I590598,I1330900);
nand I_34594 (I590632,I590615,I590457);
nor I_34595 (I590270,I590375,I590632);
nor I_34596 (I590663,I590598,I1330915);
and I_34597 (I590680,I590663,I1330924);
or I_34598 (I590697,I590680,I1330912);
DFFARX1 I_34599 (I590697,I2507,I590290,I590723,);
nor I_34600 (I590731,I590723,I590474);
DFFARX1 I_34601 (I590731,I2507,I590290,I590258,);
DFFARX1 I_34602 (I590723,I2507,I590290,I590282,);
not I_34603 (I590776,I590723);
nor I_34604 (I590793,I590776,I590350);
nor I_34605 (I590810,I590615,I590793);
DFFARX1 I_34606 (I590810,I2507,I590290,I590279,);
not I_34607 (I590868,I2514);
DFFARX1 I_34608 (I244850,I2507,I590868,I590894,);
not I_34609 (I590902,I590894);
DFFARX1 I_34610 (I244835,I2507,I590868,I590928,);
not I_34611 (I590936,I244853);
nand I_34612 (I590953,I590936,I244838);
not I_34613 (I590970,I590953);
nor I_34614 (I590987,I590970,I244835);
nor I_34615 (I591004,I590902,I590987);
DFFARX1 I_34616 (I591004,I2507,I590868,I590854,);
not I_34617 (I591035,I244835);
nand I_34618 (I591052,I591035,I590970);
and I_34619 (I591069,I591035,I244838);
nand I_34620 (I591086,I591069,I244859);
nor I_34621 (I590851,I591086,I591035);
and I_34622 (I590842,I590928,I591086);
not I_34623 (I591131,I591086);
nand I_34624 (I590845,I590928,I591131);
nor I_34625 (I590839,I590894,I591086);
not I_34626 (I591176,I244847);
nor I_34627 (I591193,I591176,I244838);
nand I_34628 (I591210,I591193,I591035);
nor I_34629 (I590848,I590953,I591210);
nor I_34630 (I591241,I591176,I244841);
and I_34631 (I591258,I591241,I244856);
or I_34632 (I591275,I591258,I244844);
DFFARX1 I_34633 (I591275,I2507,I590868,I591301,);
nor I_34634 (I591309,I591301,I591052);
DFFARX1 I_34635 (I591309,I2507,I590868,I590836,);
DFFARX1 I_34636 (I591301,I2507,I590868,I590860,);
not I_34637 (I591354,I591301);
nor I_34638 (I591371,I591354,I590928);
nor I_34639 (I591388,I591193,I591371);
DFFARX1 I_34640 (I591388,I2507,I590868,I590857,);
not I_34641 (I591446,I2514);
DFFARX1 I_34642 (I486043,I2507,I591446,I591472,);
not I_34643 (I591480,I591472);
DFFARX1 I_34644 (I486055,I2507,I591446,I591506,);
not I_34645 (I591514,I486031);
nand I_34646 (I591531,I591514,I486058);
not I_34647 (I591548,I591531);
nor I_34648 (I591565,I591548,I486046);
nor I_34649 (I591582,I591480,I591565);
DFFARX1 I_34650 (I591582,I2507,I591446,I591432,);
not I_34651 (I591613,I486046);
nand I_34652 (I591630,I591613,I591548);
and I_34653 (I591647,I591613,I486031);
nand I_34654 (I591664,I591647,I486034);
nor I_34655 (I591429,I591664,I591613);
and I_34656 (I591420,I591506,I591664);
not I_34657 (I591709,I591664);
nand I_34658 (I591423,I591506,I591709);
nor I_34659 (I591417,I591472,I591664);
not I_34660 (I591754,I486040);
nor I_34661 (I591771,I591754,I486031);
nand I_34662 (I591788,I591771,I591613);
nor I_34663 (I591426,I591531,I591788);
nor I_34664 (I591819,I591754,I486049);
and I_34665 (I591836,I591819,I486037);
or I_34666 (I591853,I591836,I486052);
DFFARX1 I_34667 (I591853,I2507,I591446,I591879,);
nor I_34668 (I591887,I591879,I591630);
DFFARX1 I_34669 (I591887,I2507,I591446,I591414,);
DFFARX1 I_34670 (I591879,I2507,I591446,I591438,);
not I_34671 (I591932,I591879);
nor I_34672 (I591949,I591932,I591506);
nor I_34673 (I591966,I591771,I591949);
DFFARX1 I_34674 (I591966,I2507,I591446,I591435,);
not I_34675 (I592024,I2514);
DFFARX1 I_34676 (I416411,I2507,I592024,I592050,);
not I_34677 (I592058,I592050);
DFFARX1 I_34678 (I416423,I2507,I592024,I592084,);
not I_34679 (I592092,I416399);
nand I_34680 (I592109,I592092,I416426);
not I_34681 (I592126,I592109);
nor I_34682 (I592143,I592126,I416414);
nor I_34683 (I592160,I592058,I592143);
DFFARX1 I_34684 (I592160,I2507,I592024,I592010,);
not I_34685 (I592191,I416414);
nand I_34686 (I592208,I592191,I592126);
and I_34687 (I592225,I592191,I416399);
nand I_34688 (I592242,I592225,I416402);
nor I_34689 (I592007,I592242,I592191);
and I_34690 (I591998,I592084,I592242);
not I_34691 (I592287,I592242);
nand I_34692 (I592001,I592084,I592287);
nor I_34693 (I591995,I592050,I592242);
not I_34694 (I592332,I416408);
nor I_34695 (I592349,I592332,I416399);
nand I_34696 (I592366,I592349,I592191);
nor I_34697 (I592004,I592109,I592366);
nor I_34698 (I592397,I592332,I416417);
and I_34699 (I592414,I592397,I416405);
or I_34700 (I592431,I592414,I416420);
DFFARX1 I_34701 (I592431,I2507,I592024,I592457,);
nor I_34702 (I592465,I592457,I592208);
DFFARX1 I_34703 (I592465,I2507,I592024,I591992,);
DFFARX1 I_34704 (I592457,I2507,I592024,I592016,);
not I_34705 (I592510,I592457);
nor I_34706 (I592527,I592510,I592084);
nor I_34707 (I592544,I592349,I592527);
DFFARX1 I_34708 (I592544,I2507,I592024,I592013,);
not I_34709 (I592602,I2514);
DFFARX1 I_34710 (I628984,I2507,I592602,I592628,);
not I_34711 (I592636,I592628);
DFFARX1 I_34712 (I628996,I2507,I592602,I592662,);
not I_34713 (I592670,I628987);
nand I_34714 (I592687,I592670,I628990);
not I_34715 (I592704,I592687);
nor I_34716 (I592721,I592704,I628993);
nor I_34717 (I592738,I592636,I592721);
DFFARX1 I_34718 (I592738,I2507,I592602,I592588,);
not I_34719 (I592769,I628993);
nand I_34720 (I592786,I592769,I592704);
and I_34721 (I592803,I592769,I628987);
nand I_34722 (I592820,I592803,I628999);
nor I_34723 (I592585,I592820,I592769);
and I_34724 (I592576,I592662,I592820);
not I_34725 (I592865,I592820);
nand I_34726 (I592579,I592662,I592865);
nor I_34727 (I592573,I592628,I592820);
not I_34728 (I592910,I629005);
nor I_34729 (I592927,I592910,I628987);
nand I_34730 (I592944,I592927,I592769);
nor I_34731 (I592582,I592687,I592944);
nor I_34732 (I592975,I592910,I628984);
and I_34733 (I592992,I592975,I629002);
or I_34734 (I593009,I592992,I629008);
DFFARX1 I_34735 (I593009,I2507,I592602,I593035,);
nor I_34736 (I593043,I593035,I592786);
DFFARX1 I_34737 (I593043,I2507,I592602,I592570,);
DFFARX1 I_34738 (I593035,I2507,I592602,I592594,);
not I_34739 (I593088,I593035);
nor I_34740 (I593105,I593088,I592662);
nor I_34741 (I593122,I592927,I593105);
DFFARX1 I_34742 (I593122,I2507,I592602,I592591,);
not I_34743 (I593180,I2514);
DFFARX1 I_34744 (I1281354,I2507,I593180,I593206,);
not I_34745 (I593214,I593206);
DFFARX1 I_34746 (I1281366,I2507,I593180,I593240,);
not I_34747 (I593248,I1281357);
nand I_34748 (I593265,I593248,I1281345);
not I_34749 (I593282,I593265);
nor I_34750 (I593299,I593282,I1281342);
nor I_34751 (I593316,I593214,I593299);
DFFARX1 I_34752 (I593316,I2507,I593180,I593166,);
not I_34753 (I593347,I1281342);
nand I_34754 (I593364,I593347,I593282);
and I_34755 (I593381,I593347,I1281348);
nand I_34756 (I593398,I593381,I1281345);
nor I_34757 (I593163,I593398,I593347);
and I_34758 (I593154,I593240,I593398);
not I_34759 (I593443,I593398);
nand I_34760 (I593157,I593240,I593443);
nor I_34761 (I593151,I593206,I593398);
not I_34762 (I593488,I1281363);
nor I_34763 (I593505,I593488,I1281348);
nand I_34764 (I593522,I593505,I593347);
nor I_34765 (I593160,I593265,I593522);
nor I_34766 (I593553,I593488,I1281351);
and I_34767 (I593570,I593553,I1281342);
or I_34768 (I593587,I593570,I1281360);
DFFARX1 I_34769 (I593587,I2507,I593180,I593613,);
nor I_34770 (I593621,I593613,I593364);
DFFARX1 I_34771 (I593621,I2507,I593180,I593148,);
DFFARX1 I_34772 (I593613,I2507,I593180,I593172,);
not I_34773 (I593666,I593613);
nor I_34774 (I593683,I593666,I593240);
nor I_34775 (I593700,I593505,I593683);
DFFARX1 I_34776 (I593700,I2507,I593180,I593169,);
not I_34777 (I593758,I2514);
DFFARX1 I_34778 (I884466,I2507,I593758,I593784,);
not I_34779 (I593792,I593784);
DFFARX1 I_34780 (I884466,I2507,I593758,I593818,);
not I_34781 (I593826,I884463);
nand I_34782 (I593843,I593826,I884478);
not I_34783 (I593860,I593843);
nor I_34784 (I593877,I593860,I884472);
nor I_34785 (I593894,I593792,I593877);
DFFARX1 I_34786 (I593894,I2507,I593758,I593744,);
not I_34787 (I593925,I884472);
nand I_34788 (I593942,I593925,I593860);
and I_34789 (I593959,I593925,I884469);
nand I_34790 (I593976,I593959,I884460);
nor I_34791 (I593741,I593976,I593925);
and I_34792 (I593732,I593818,I593976);
not I_34793 (I594021,I593976);
nand I_34794 (I593735,I593818,I594021);
nor I_34795 (I593729,I593784,I593976);
not I_34796 (I594066,I884481);
nor I_34797 (I594083,I594066,I884469);
nand I_34798 (I594100,I594083,I593925);
nor I_34799 (I593738,I593843,I594100);
nor I_34800 (I594131,I594066,I884460);
and I_34801 (I594148,I594131,I884463);
or I_34802 (I594165,I594148,I884475);
DFFARX1 I_34803 (I594165,I2507,I593758,I594191,);
nor I_34804 (I594199,I594191,I593942);
DFFARX1 I_34805 (I594199,I2507,I593758,I593726,);
DFFARX1 I_34806 (I594191,I2507,I593758,I593750,);
not I_34807 (I594244,I594191);
nor I_34808 (I594261,I594244,I593818);
nor I_34809 (I594278,I594083,I594261);
DFFARX1 I_34810 (I594278,I2507,I593758,I593747,);
not I_34811 (I594336,I2514);
DFFARX1 I_34812 (I663664,I2507,I594336,I594362,);
not I_34813 (I594370,I594362);
DFFARX1 I_34814 (I663676,I2507,I594336,I594396,);
not I_34815 (I594404,I663667);
nand I_34816 (I594421,I594404,I663670);
not I_34817 (I594438,I594421);
nor I_34818 (I594455,I594438,I663673);
nor I_34819 (I594472,I594370,I594455);
DFFARX1 I_34820 (I594472,I2507,I594336,I594322,);
not I_34821 (I594503,I663673);
nand I_34822 (I594520,I594503,I594438);
and I_34823 (I594537,I594503,I663667);
nand I_34824 (I594554,I594537,I663679);
nor I_34825 (I594319,I594554,I594503);
and I_34826 (I594310,I594396,I594554);
not I_34827 (I594599,I594554);
nand I_34828 (I594313,I594396,I594599);
nor I_34829 (I594307,I594362,I594554);
not I_34830 (I594644,I663685);
nor I_34831 (I594661,I594644,I663667);
nand I_34832 (I594678,I594661,I594503);
nor I_34833 (I594316,I594421,I594678);
nor I_34834 (I594709,I594644,I663664);
and I_34835 (I594726,I594709,I663682);
or I_34836 (I594743,I594726,I663688);
DFFARX1 I_34837 (I594743,I2507,I594336,I594769,);
nor I_34838 (I594777,I594769,I594520);
DFFARX1 I_34839 (I594777,I2507,I594336,I594304,);
DFFARX1 I_34840 (I594769,I2507,I594336,I594328,);
not I_34841 (I594822,I594769);
nor I_34842 (I594839,I594822,I594396);
nor I_34843 (I594856,I594661,I594839);
DFFARX1 I_34844 (I594856,I2507,I594336,I594325,);
not I_34845 (I594914,I2514);
DFFARX1 I_34846 (I1379092,I2507,I594914,I594940,);
not I_34847 (I594948,I594940);
DFFARX1 I_34848 (I1379092,I2507,I594914,I594974,);
not I_34849 (I594982,I1379116);
nand I_34850 (I594999,I594982,I1379098);
not I_34851 (I595016,I594999);
nor I_34852 (I595033,I595016,I1379113);
nor I_34853 (I595050,I594948,I595033);
DFFARX1 I_34854 (I595050,I2507,I594914,I594900,);
not I_34855 (I595081,I1379113);
nand I_34856 (I595098,I595081,I595016);
and I_34857 (I595115,I595081,I1379095);
nand I_34858 (I595132,I595115,I1379104);
nor I_34859 (I594897,I595132,I595081);
and I_34860 (I594888,I594974,I595132);
not I_34861 (I595177,I595132);
nand I_34862 (I594891,I594974,I595177);
nor I_34863 (I594885,I594940,I595132);
not I_34864 (I595222,I1379101);
nor I_34865 (I595239,I595222,I1379095);
nand I_34866 (I595256,I595239,I595081);
nor I_34867 (I594894,I594999,I595256);
nor I_34868 (I595287,I595222,I1379110);
and I_34869 (I595304,I595287,I1379119);
or I_34870 (I595321,I595304,I1379107);
DFFARX1 I_34871 (I595321,I2507,I594914,I595347,);
nor I_34872 (I595355,I595347,I595098);
DFFARX1 I_34873 (I595355,I2507,I594914,I594882,);
DFFARX1 I_34874 (I595347,I2507,I594914,I594906,);
not I_34875 (I595400,I595347);
nor I_34876 (I595417,I595400,I594974);
nor I_34877 (I595434,I595239,I595417);
DFFARX1 I_34878 (I595434,I2507,I594914,I594903,);
not I_34879 (I595492,I2514);
DFFARX1 I_34880 (I305531,I2507,I595492,I595518,);
not I_34881 (I595526,I595518);
DFFARX1 I_34882 (I305546,I2507,I595492,I595552,);
not I_34883 (I595560,I305549);
nand I_34884 (I595577,I595560,I305528);
not I_34885 (I595594,I595577);
nor I_34886 (I595611,I595594,I305552);
nor I_34887 (I595628,I595526,I595611);
DFFARX1 I_34888 (I595628,I2507,I595492,I595478,);
not I_34889 (I595659,I305552);
nand I_34890 (I595676,I595659,I595594);
and I_34891 (I595693,I595659,I305534);
nand I_34892 (I595710,I595693,I305525);
nor I_34893 (I595475,I595710,I595659);
and I_34894 (I595466,I595552,I595710);
not I_34895 (I595755,I595710);
nand I_34896 (I595469,I595552,I595755);
nor I_34897 (I595463,I595518,I595710);
not I_34898 (I595800,I305525);
nor I_34899 (I595817,I595800,I305534);
nand I_34900 (I595834,I595817,I595659);
nor I_34901 (I595472,I595577,I595834);
nor I_34902 (I595865,I595800,I305540);
and I_34903 (I595882,I595865,I305543);
or I_34904 (I595899,I595882,I305537);
DFFARX1 I_34905 (I595899,I2507,I595492,I595925,);
nor I_34906 (I595933,I595925,I595676);
DFFARX1 I_34907 (I595933,I2507,I595492,I595460,);
DFFARX1 I_34908 (I595925,I2507,I595492,I595484,);
not I_34909 (I595978,I595925);
nor I_34910 (I595995,I595978,I595552);
nor I_34911 (I596012,I595817,I595995);
DFFARX1 I_34912 (I596012,I2507,I595492,I595481,);
not I_34913 (I596070,I2514);
DFFARX1 I_34914 (I271276,I2507,I596070,I596096,);
not I_34915 (I596104,I596096);
DFFARX1 I_34916 (I271291,I2507,I596070,I596130,);
not I_34917 (I596138,I271294);
nand I_34918 (I596155,I596138,I271273);
not I_34919 (I596172,I596155);
nor I_34920 (I596189,I596172,I271297);
nor I_34921 (I596206,I596104,I596189);
DFFARX1 I_34922 (I596206,I2507,I596070,I596056,);
not I_34923 (I596237,I271297);
nand I_34924 (I596254,I596237,I596172);
and I_34925 (I596271,I596237,I271279);
nand I_34926 (I596288,I596271,I271270);
nor I_34927 (I596053,I596288,I596237);
and I_34928 (I596044,I596130,I596288);
not I_34929 (I596333,I596288);
nand I_34930 (I596047,I596130,I596333);
nor I_34931 (I596041,I596096,I596288);
not I_34932 (I596378,I271270);
nor I_34933 (I596395,I596378,I271279);
nand I_34934 (I596412,I596395,I596237);
nor I_34935 (I596050,I596155,I596412);
nor I_34936 (I596443,I596378,I271285);
and I_34937 (I596460,I596443,I271288);
or I_34938 (I596477,I596460,I271282);
DFFARX1 I_34939 (I596477,I2507,I596070,I596503,);
nor I_34940 (I596511,I596503,I596254);
DFFARX1 I_34941 (I596511,I2507,I596070,I596038,);
DFFARX1 I_34942 (I596503,I2507,I596070,I596062,);
not I_34943 (I596556,I596503);
nor I_34944 (I596573,I596556,I596130);
nor I_34945 (I596590,I596395,I596573);
DFFARX1 I_34946 (I596590,I2507,I596070,I596059,);
not I_34947 (I596648,I2514);
DFFARX1 I_34948 (I1014089,I2507,I596648,I596674,);
not I_34949 (I596682,I596674);
DFFARX1 I_34950 (I1014080,I2507,I596648,I596708,);
not I_34951 (I596716,I1014074);
nand I_34952 (I596733,I596716,I1014086);
not I_34953 (I596750,I596733);
nor I_34954 (I596767,I596750,I1014077);
nor I_34955 (I596784,I596682,I596767);
DFFARX1 I_34956 (I596784,I2507,I596648,I596634,);
not I_34957 (I596815,I1014077);
nand I_34958 (I596832,I596815,I596750);
and I_34959 (I596849,I596815,I1014083);
nand I_34960 (I596866,I596849,I1014068);
nor I_34961 (I596631,I596866,I596815);
and I_34962 (I596622,I596708,I596866);
not I_34963 (I596911,I596866);
nand I_34964 (I596625,I596708,I596911);
nor I_34965 (I596619,I596674,I596866);
not I_34966 (I596956,I1014068);
nor I_34967 (I596973,I596956,I1014083);
nand I_34968 (I596990,I596973,I596815);
nor I_34969 (I596628,I596733,I596990);
nor I_34970 (I597021,I596956,I1014071);
and I_34971 (I597038,I597021,I1014074);
or I_34972 (I597055,I597038,I1014071);
DFFARX1 I_34973 (I597055,I2507,I596648,I597081,);
nor I_34974 (I597089,I597081,I596832);
DFFARX1 I_34975 (I597089,I2507,I596648,I596616,);
DFFARX1 I_34976 (I597081,I2507,I596648,I596640,);
not I_34977 (I597134,I597081);
nor I_34978 (I597151,I597134,I596708);
nor I_34979 (I597168,I596973,I597151);
DFFARX1 I_34980 (I597168,I2507,I596648,I596637,);
not I_34981 (I597226,I2514);
DFFARX1 I_34982 (I806997,I2507,I597226,I597252,);
not I_34983 (I597260,I597252);
DFFARX1 I_34984 (I806997,I2507,I597226,I597286,);
not I_34985 (I597294,I806994);
nand I_34986 (I597311,I597294,I807009);
not I_34987 (I597328,I597311);
nor I_34988 (I597345,I597328,I807003);
nor I_34989 (I597362,I597260,I597345);
DFFARX1 I_34990 (I597362,I2507,I597226,I597212,);
not I_34991 (I597393,I807003);
nand I_34992 (I597410,I597393,I597328);
and I_34993 (I597427,I597393,I807000);
nand I_34994 (I597444,I597427,I806991);
nor I_34995 (I597209,I597444,I597393);
and I_34996 (I597200,I597286,I597444);
not I_34997 (I597489,I597444);
nand I_34998 (I597203,I597286,I597489);
nor I_34999 (I597197,I597252,I597444);
not I_35000 (I597534,I807012);
nor I_35001 (I597551,I597534,I807000);
nand I_35002 (I597568,I597551,I597393);
nor I_35003 (I597206,I597311,I597568);
nor I_35004 (I597599,I597534,I806991);
and I_35005 (I597616,I597599,I806994);
or I_35006 (I597633,I597616,I807006);
DFFARX1 I_35007 (I597633,I2507,I597226,I597659,);
nor I_35008 (I597667,I597659,I597410);
DFFARX1 I_35009 (I597667,I2507,I597226,I597194,);
DFFARX1 I_35010 (I597659,I2507,I597226,I597218,);
not I_35011 (I597712,I597659);
nor I_35012 (I597729,I597712,I597286);
nor I_35013 (I597746,I597551,I597729);
DFFARX1 I_35014 (I597746,I2507,I597226,I597215,);
not I_35015 (I597804,I2514);
DFFARX1 I_35016 (I1206900,I2507,I597804,I597830,);
not I_35017 (I597838,I597830);
DFFARX1 I_35018 (I1206894,I2507,I597804,I597864,);
not I_35019 (I597872,I1206903);
nand I_35020 (I597889,I597872,I1206882);
not I_35021 (I597906,I597889);
nor I_35022 (I597923,I597906,I1206891);
nor I_35023 (I597940,I597838,I597923);
DFFARX1 I_35024 (I597940,I2507,I597804,I597790,);
not I_35025 (I597971,I1206891);
nand I_35026 (I597988,I597971,I597906);
and I_35027 (I598005,I597971,I1206906);
nand I_35028 (I598022,I598005,I1206885);
nor I_35029 (I597787,I598022,I597971);
and I_35030 (I597778,I597864,I598022);
not I_35031 (I598067,I598022);
nand I_35032 (I597781,I597864,I598067);
nor I_35033 (I597775,I597830,I598022);
not I_35034 (I598112,I1206888);
nor I_35035 (I598129,I598112,I1206906);
nand I_35036 (I598146,I598129,I597971);
nor I_35037 (I597784,I597889,I598146);
nor I_35038 (I598177,I598112,I1206897);
and I_35039 (I598194,I598177,I1206885);
or I_35040 (I598211,I598194,I1206882);
DFFARX1 I_35041 (I598211,I2507,I597804,I598237,);
nor I_35042 (I598245,I598237,I597988);
DFFARX1 I_35043 (I598245,I2507,I597804,I597772,);
DFFARX1 I_35044 (I598237,I2507,I597804,I597796,);
not I_35045 (I598290,I598237);
nor I_35046 (I598307,I598290,I597864);
nor I_35047 (I598324,I598129,I598307);
DFFARX1 I_35048 (I598324,I2507,I597804,I597793,);
not I_35049 (I598382,I2514);
DFFARX1 I_35050 (I852846,I2507,I598382,I598408,);
not I_35051 (I598416,I598408);
DFFARX1 I_35052 (I852846,I2507,I598382,I598442,);
not I_35053 (I598450,I852843);
nand I_35054 (I598467,I598450,I852858);
not I_35055 (I598484,I598467);
nor I_35056 (I598501,I598484,I852852);
nor I_35057 (I598518,I598416,I598501);
DFFARX1 I_35058 (I598518,I2507,I598382,I598368,);
not I_35059 (I598549,I852852);
nand I_35060 (I598566,I598549,I598484);
and I_35061 (I598583,I598549,I852849);
nand I_35062 (I598600,I598583,I852840);
nor I_35063 (I598365,I598600,I598549);
and I_35064 (I598356,I598442,I598600);
not I_35065 (I598645,I598600);
nand I_35066 (I598359,I598442,I598645);
nor I_35067 (I598353,I598408,I598600);
not I_35068 (I598690,I852861);
nor I_35069 (I598707,I598690,I852849);
nand I_35070 (I598724,I598707,I598549);
nor I_35071 (I598362,I598467,I598724);
nor I_35072 (I598755,I598690,I852840);
and I_35073 (I598772,I598755,I852843);
or I_35074 (I598789,I598772,I852855);
DFFARX1 I_35075 (I598789,I2507,I598382,I598815,);
nor I_35076 (I598823,I598815,I598566);
DFFARX1 I_35077 (I598823,I2507,I598382,I598350,);
DFFARX1 I_35078 (I598815,I2507,I598382,I598374,);
not I_35079 (I598868,I598815);
nor I_35080 (I598885,I598868,I598442);
nor I_35081 (I598902,I598707,I598885);
DFFARX1 I_35082 (I598902,I2507,I598382,I598371,);
not I_35083 (I598960,I2514);
DFFARX1 I_35084 (I1385637,I2507,I598960,I598986,);
not I_35085 (I598994,I598986);
DFFARX1 I_35086 (I1385637,I2507,I598960,I599020,);
not I_35087 (I599028,I1385661);
nand I_35088 (I599045,I599028,I1385643);
not I_35089 (I599062,I599045);
nor I_35090 (I599079,I599062,I1385658);
nor I_35091 (I599096,I598994,I599079);
DFFARX1 I_35092 (I599096,I2507,I598960,I598946,);
not I_35093 (I599127,I1385658);
nand I_35094 (I599144,I599127,I599062);
and I_35095 (I599161,I599127,I1385640);
nand I_35096 (I599178,I599161,I1385649);
nor I_35097 (I598943,I599178,I599127);
and I_35098 (I598934,I599020,I599178);
not I_35099 (I599223,I599178);
nand I_35100 (I598937,I599020,I599223);
nor I_35101 (I598931,I598986,I599178);
not I_35102 (I599268,I1385646);
nor I_35103 (I599285,I599268,I1385640);
nand I_35104 (I599302,I599285,I599127);
nor I_35105 (I598940,I599045,I599302);
nor I_35106 (I599333,I599268,I1385655);
and I_35107 (I599350,I599333,I1385664);
or I_35108 (I599367,I599350,I1385652);
DFFARX1 I_35109 (I599367,I2507,I598960,I599393,);
nor I_35110 (I599401,I599393,I599144);
DFFARX1 I_35111 (I599401,I2507,I598960,I598928,);
DFFARX1 I_35112 (I599393,I2507,I598960,I598952,);
not I_35113 (I599446,I599393);
nor I_35114 (I599463,I599446,I599020);
nor I_35115 (I599480,I599285,I599463);
DFFARX1 I_35116 (I599480,I2507,I598960,I598949,);
not I_35117 (I599538,I2514);
DFFARX1 I_35118 (I1296931,I2507,I599538,I599564,);
not I_35119 (I599572,I599564);
DFFARX1 I_35120 (I1296949,I2507,I599538,I599598,);
not I_35121 (I599606,I1296946);
nand I_35122 (I599623,I599606,I1296937);
not I_35123 (I599640,I599623);
nor I_35124 (I599657,I599640,I1296934);
nor I_35125 (I599674,I599572,I599657);
DFFARX1 I_35126 (I599674,I2507,I599538,I599524,);
not I_35127 (I599705,I1296934);
nand I_35128 (I599722,I599705,I599640);
and I_35129 (I599739,I599705,I1296940);
nand I_35130 (I599756,I599739,I1296955);
nor I_35131 (I599521,I599756,I599705);
and I_35132 (I599512,I599598,I599756);
not I_35133 (I599801,I599756);
nand I_35134 (I599515,I599598,I599801);
nor I_35135 (I599509,I599564,I599756);
not I_35136 (I599846,I1296931);
nor I_35137 (I599863,I599846,I1296940);
nand I_35138 (I599880,I599863,I599705);
nor I_35139 (I599518,I599623,I599880);
nor I_35140 (I599911,I599846,I1296952);
and I_35141 (I599928,I599911,I1296943);
or I_35142 (I599945,I599928,I1296958);
DFFARX1 I_35143 (I599945,I2507,I599538,I599971,);
nor I_35144 (I599979,I599971,I599722);
DFFARX1 I_35145 (I599979,I2507,I599538,I599506,);
DFFARX1 I_35146 (I599971,I2507,I599538,I599530,);
not I_35147 (I600024,I599971);
nor I_35148 (I600041,I600024,I599598);
nor I_35149 (I600058,I599863,I600041);
DFFARX1 I_35150 (I600058,I2507,I599538,I599527,);
not I_35151 (I600116,I2514);
DFFARX1 I_35152 (I973495,I2507,I600116,I600142,);
not I_35153 (I600150,I600142);
DFFARX1 I_35154 (I973492,I2507,I600116,I600176,);
not I_35155 (I600184,I973489);
nand I_35156 (I600201,I600184,I973516);
not I_35157 (I600218,I600201);
nor I_35158 (I600235,I600218,I973504);
nor I_35159 (I600252,I600150,I600235);
DFFARX1 I_35160 (I600252,I2507,I600116,I600102,);
not I_35161 (I600283,I973504);
nand I_35162 (I600300,I600283,I600218);
and I_35163 (I600317,I600283,I973510);
nand I_35164 (I600334,I600317,I973501);
nor I_35165 (I600099,I600334,I600283);
and I_35166 (I600090,I600176,I600334);
not I_35167 (I600379,I600334);
nand I_35168 (I600093,I600176,I600379);
nor I_35169 (I600087,I600142,I600334);
not I_35170 (I600424,I973498);
nor I_35171 (I600441,I600424,I973510);
nand I_35172 (I600458,I600441,I600283);
nor I_35173 (I600096,I600201,I600458);
nor I_35174 (I600489,I600424,I973513);
and I_35175 (I600506,I600489,I973507);
or I_35176 (I600523,I600506,I973489);
DFFARX1 I_35177 (I600523,I2507,I600116,I600549,);
nor I_35178 (I600557,I600549,I600300);
DFFARX1 I_35179 (I600557,I2507,I600116,I600084,);
DFFARX1 I_35180 (I600549,I2507,I600116,I600108,);
not I_35181 (I600602,I600549);
nor I_35182 (I600619,I600602,I600176);
nor I_35183 (I600636,I600441,I600619);
DFFARX1 I_35184 (I600636,I2507,I600116,I600105,);
not I_35185 (I600694,I2514);
DFFARX1 I_35186 (I794349,I2507,I600694,I600720,);
not I_35187 (I600728,I600720);
DFFARX1 I_35188 (I794349,I2507,I600694,I600754,);
not I_35189 (I600762,I794346);
nand I_35190 (I600779,I600762,I794361);
not I_35191 (I600796,I600779);
nor I_35192 (I600813,I600796,I794355);
nor I_35193 (I600830,I600728,I600813);
DFFARX1 I_35194 (I600830,I2507,I600694,I600680,);
not I_35195 (I600861,I794355);
nand I_35196 (I600878,I600861,I600796);
and I_35197 (I600895,I600861,I794352);
nand I_35198 (I600912,I600895,I794343);
nor I_35199 (I600677,I600912,I600861);
and I_35200 (I600668,I600754,I600912);
not I_35201 (I600957,I600912);
nand I_35202 (I600671,I600754,I600957);
nor I_35203 (I600665,I600720,I600912);
not I_35204 (I601002,I794364);
nor I_35205 (I601019,I601002,I794352);
nand I_35206 (I601036,I601019,I600861);
nor I_35207 (I600674,I600779,I601036);
nor I_35208 (I601067,I601002,I794343);
and I_35209 (I601084,I601067,I794346);
or I_35210 (I601101,I601084,I794358);
DFFARX1 I_35211 (I601101,I2507,I600694,I601127,);
nor I_35212 (I601135,I601127,I600878);
DFFARX1 I_35213 (I601135,I2507,I600694,I600662,);
DFFARX1 I_35214 (I601127,I2507,I600694,I600686,);
not I_35215 (I601180,I601127);
nor I_35216 (I601197,I601180,I600754);
nor I_35217 (I601214,I601019,I601197);
DFFARX1 I_35218 (I601214,I2507,I600694,I600683,);
not I_35219 (I601272,I2514);
DFFARX1 I_35220 (I858643,I2507,I601272,I601298,);
not I_35221 (I601306,I601298);
DFFARX1 I_35222 (I858643,I2507,I601272,I601332,);
not I_35223 (I601340,I858640);
nand I_35224 (I601357,I601340,I858655);
not I_35225 (I601374,I601357);
nor I_35226 (I601391,I601374,I858649);
nor I_35227 (I601408,I601306,I601391);
DFFARX1 I_35228 (I601408,I2507,I601272,I601258,);
not I_35229 (I601439,I858649);
nand I_35230 (I601456,I601439,I601374);
and I_35231 (I601473,I601439,I858646);
nand I_35232 (I601490,I601473,I858637);
nor I_35233 (I601255,I601490,I601439);
and I_35234 (I601246,I601332,I601490);
not I_35235 (I601535,I601490);
nand I_35236 (I601249,I601332,I601535);
nor I_35237 (I601243,I601298,I601490);
not I_35238 (I601580,I858658);
nor I_35239 (I601597,I601580,I858646);
nand I_35240 (I601614,I601597,I601439);
nor I_35241 (I601252,I601357,I601614);
nor I_35242 (I601645,I601580,I858637);
and I_35243 (I601662,I601645,I858640);
or I_35244 (I601679,I601662,I858652);
DFFARX1 I_35245 (I601679,I2507,I601272,I601705,);
nor I_35246 (I601713,I601705,I601456);
DFFARX1 I_35247 (I601713,I2507,I601272,I601240,);
DFFARX1 I_35248 (I601705,I2507,I601272,I601264,);
not I_35249 (I601758,I601705);
nor I_35250 (I601775,I601758,I601332);
nor I_35251 (I601792,I601597,I601775);
DFFARX1 I_35252 (I601792,I2507,I601272,I601261,);
not I_35253 (I601850,I2514);
DFFARX1 I_35254 (I266006,I2507,I601850,I601876,);
not I_35255 (I601884,I601876);
DFFARX1 I_35256 (I266021,I2507,I601850,I601910,);
not I_35257 (I601918,I266024);
nand I_35258 (I601935,I601918,I266003);
not I_35259 (I601952,I601935);
nor I_35260 (I601969,I601952,I266027);
nor I_35261 (I601986,I601884,I601969);
DFFARX1 I_35262 (I601986,I2507,I601850,I601836,);
not I_35263 (I602017,I266027);
nand I_35264 (I602034,I602017,I601952);
and I_35265 (I602051,I602017,I266009);
nand I_35266 (I602068,I602051,I266000);
nor I_35267 (I601833,I602068,I602017);
and I_35268 (I601824,I601910,I602068);
not I_35269 (I602113,I602068);
nand I_35270 (I601827,I601910,I602113);
nor I_35271 (I601821,I601876,I602068);
not I_35272 (I602158,I266000);
nor I_35273 (I602175,I602158,I266009);
nand I_35274 (I602192,I602175,I602017);
nor I_35275 (I601830,I601935,I602192);
nor I_35276 (I602223,I602158,I266015);
and I_35277 (I602240,I602223,I266018);
or I_35278 (I602257,I602240,I266012);
DFFARX1 I_35279 (I602257,I2507,I601850,I602283,);
nor I_35280 (I602291,I602283,I602034);
DFFARX1 I_35281 (I602291,I2507,I601850,I601818,);
DFFARX1 I_35282 (I602283,I2507,I601850,I601842,);
not I_35283 (I602336,I602283);
nor I_35284 (I602353,I602336,I601910);
nor I_35285 (I602370,I602175,I602353);
DFFARX1 I_35286 (I602370,I2507,I601850,I601839,);
not I_35287 (I602428,I2514);
DFFARX1 I_35288 (I1227572,I2507,I602428,I602454,);
not I_35289 (I602462,I602454);
DFFARX1 I_35290 (I1227566,I2507,I602428,I602488,);
not I_35291 (I602496,I1227575);
nand I_35292 (I602513,I602496,I1227554);
not I_35293 (I602530,I602513);
nor I_35294 (I602547,I602530,I1227563);
nor I_35295 (I602564,I602462,I602547);
DFFARX1 I_35296 (I602564,I2507,I602428,I602414,);
not I_35297 (I602595,I1227563);
nand I_35298 (I602612,I602595,I602530);
and I_35299 (I602629,I602595,I1227578);
nand I_35300 (I602646,I602629,I1227557);
nor I_35301 (I602411,I602646,I602595);
and I_35302 (I602402,I602488,I602646);
not I_35303 (I602691,I602646);
nand I_35304 (I602405,I602488,I602691);
nor I_35305 (I602399,I602454,I602646);
not I_35306 (I602736,I1227560);
nor I_35307 (I602753,I602736,I1227578);
nand I_35308 (I602770,I602753,I602595);
nor I_35309 (I602408,I602513,I602770);
nor I_35310 (I602801,I602736,I1227569);
and I_35311 (I602818,I602801,I1227557);
or I_35312 (I602835,I602818,I1227554);
DFFARX1 I_35313 (I602835,I2507,I602428,I602861,);
nor I_35314 (I602869,I602861,I602612);
DFFARX1 I_35315 (I602869,I2507,I602428,I602396,);
DFFARX1 I_35316 (I602861,I2507,I602428,I602420,);
not I_35317 (I602914,I602861);
nor I_35318 (I602931,I602914,I602488);
nor I_35319 (I602948,I602753,I602931);
DFFARX1 I_35320 (I602948,I2507,I602428,I602417,);
not I_35321 (I603006,I2514);
DFFARX1 I_35322 (I926337,I2507,I603006,I603032,);
not I_35323 (I603040,I603032);
DFFARX1 I_35324 (I926334,I2507,I603006,I603066,);
not I_35325 (I603074,I926331);
nand I_35326 (I603091,I603074,I926358);
not I_35327 (I603108,I603091);
nor I_35328 (I603125,I603108,I926346);
nor I_35329 (I603142,I603040,I603125);
DFFARX1 I_35330 (I603142,I2507,I603006,I602992,);
not I_35331 (I603173,I926346);
nand I_35332 (I603190,I603173,I603108);
and I_35333 (I603207,I603173,I926352);
nand I_35334 (I603224,I603207,I926343);
nor I_35335 (I602989,I603224,I603173);
and I_35336 (I602980,I603066,I603224);
not I_35337 (I603269,I603224);
nand I_35338 (I602983,I603066,I603269);
nor I_35339 (I602977,I603032,I603224);
not I_35340 (I603314,I926340);
nor I_35341 (I603331,I603314,I926352);
nand I_35342 (I603348,I603331,I603173);
nor I_35343 (I602986,I603091,I603348);
nor I_35344 (I603379,I603314,I926355);
and I_35345 (I603396,I603379,I926349);
or I_35346 (I603413,I603396,I926331);
DFFARX1 I_35347 (I603413,I2507,I603006,I603439,);
nor I_35348 (I603447,I603439,I603190);
DFFARX1 I_35349 (I603447,I2507,I603006,I602974,);
DFFARX1 I_35350 (I603439,I2507,I603006,I602998,);
not I_35351 (I603492,I603439);
nor I_35352 (I603509,I603492,I603066);
nor I_35353 (I603526,I603331,I603509);
DFFARX1 I_35354 (I603526,I2507,I603006,I602995,);
not I_35355 (I603584,I2514);
DFFARX1 I_35356 (I1852,I2507,I603584,I603610,);
not I_35357 (I603618,I603610);
DFFARX1 I_35358 (I2412,I2507,I603584,I603644,);
not I_35359 (I603652,I2180);
nand I_35360 (I603669,I603652,I2092);
not I_35361 (I603686,I603669);
nor I_35362 (I603703,I603686,I1556);
nor I_35363 (I603720,I603618,I603703);
DFFARX1 I_35364 (I603720,I2507,I603584,I603570,);
not I_35365 (I603751,I1556);
nand I_35366 (I603768,I603751,I603686);
and I_35367 (I603785,I603751,I2396);
nand I_35368 (I603802,I603785,I1708);
nor I_35369 (I603567,I603802,I603751);
and I_35370 (I603558,I603644,I603802);
not I_35371 (I603847,I603802);
nand I_35372 (I603561,I603644,I603847);
nor I_35373 (I603555,I603610,I603802);
not I_35374 (I603892,I1644);
nor I_35375 (I603909,I603892,I2396);
nand I_35376 (I603926,I603909,I603751);
nor I_35377 (I603564,I603669,I603926);
nor I_35378 (I603957,I603892,I2028);
and I_35379 (I603974,I603957,I1900);
or I_35380 (I603991,I603974,I2436);
DFFARX1 I_35381 (I603991,I2507,I603584,I604017,);
nor I_35382 (I604025,I604017,I603768);
DFFARX1 I_35383 (I604025,I2507,I603584,I603552,);
DFFARX1 I_35384 (I604017,I2507,I603584,I603576,);
not I_35385 (I604070,I604017);
nor I_35386 (I604087,I604070,I603644);
nor I_35387 (I604104,I603909,I604087);
DFFARX1 I_35388 (I604104,I2507,I603584,I603573,);
not I_35389 (I604162,I2514);
DFFARX1 I_35390 (I1280198,I2507,I604162,I604188,);
not I_35391 (I604196,I604188);
DFFARX1 I_35392 (I1280210,I2507,I604162,I604222,);
not I_35393 (I604230,I1280201);
nand I_35394 (I604247,I604230,I1280189);
not I_35395 (I604264,I604247);
nor I_35396 (I604281,I604264,I1280186);
nor I_35397 (I604298,I604196,I604281);
DFFARX1 I_35398 (I604298,I2507,I604162,I604148,);
not I_35399 (I604329,I1280186);
nand I_35400 (I604346,I604329,I604264);
and I_35401 (I604363,I604329,I1280192);
nand I_35402 (I604380,I604363,I1280189);
nor I_35403 (I604145,I604380,I604329);
and I_35404 (I604136,I604222,I604380);
not I_35405 (I604425,I604380);
nand I_35406 (I604139,I604222,I604425);
nor I_35407 (I604133,I604188,I604380);
not I_35408 (I604470,I1280207);
nor I_35409 (I604487,I604470,I1280192);
nand I_35410 (I604504,I604487,I604329);
nor I_35411 (I604142,I604247,I604504);
nor I_35412 (I604535,I604470,I1280195);
and I_35413 (I604552,I604535,I1280186);
or I_35414 (I604569,I604552,I1280204);
DFFARX1 I_35415 (I604569,I2507,I604162,I604595,);
nor I_35416 (I604603,I604595,I604346);
DFFARX1 I_35417 (I604603,I2507,I604162,I604130,);
DFFARX1 I_35418 (I604595,I2507,I604162,I604154,);
not I_35419 (I604648,I604595);
nor I_35420 (I604665,I604648,I604222);
nor I_35421 (I604682,I604487,I604665);
DFFARX1 I_35422 (I604682,I2507,I604162,I604151,);
not I_35423 (I604740,I2514);
DFFARX1 I_35424 (I1383852,I2507,I604740,I604766,);
not I_35425 (I604774,I604766);
DFFARX1 I_35426 (I1383852,I2507,I604740,I604800,);
not I_35427 (I604808,I1383876);
nand I_35428 (I604825,I604808,I1383858);
not I_35429 (I604842,I604825);
nor I_35430 (I604859,I604842,I1383873);
nor I_35431 (I604876,I604774,I604859);
DFFARX1 I_35432 (I604876,I2507,I604740,I604726,);
not I_35433 (I604907,I1383873);
nand I_35434 (I604924,I604907,I604842);
and I_35435 (I604941,I604907,I1383855);
nand I_35436 (I604958,I604941,I1383864);
nor I_35437 (I604723,I604958,I604907);
and I_35438 (I604714,I604800,I604958);
not I_35439 (I605003,I604958);
nand I_35440 (I604717,I604800,I605003);
nor I_35441 (I604711,I604766,I604958);
not I_35442 (I605048,I1383861);
nor I_35443 (I605065,I605048,I1383855);
nand I_35444 (I605082,I605065,I604907);
nor I_35445 (I604720,I604825,I605082);
nor I_35446 (I605113,I605048,I1383870);
and I_35447 (I605130,I605113,I1383879);
or I_35448 (I605147,I605130,I1383867);
DFFARX1 I_35449 (I605147,I2507,I604740,I605173,);
nor I_35450 (I605181,I605173,I604924);
DFFARX1 I_35451 (I605181,I2507,I604740,I604708,);
DFFARX1 I_35452 (I605173,I2507,I604740,I604732,);
not I_35453 (I605226,I605173);
nor I_35454 (I605243,I605226,I604800);
nor I_35455 (I605260,I605065,I605243);
DFFARX1 I_35456 (I605260,I2507,I604740,I604729,);
not I_35457 (I605318,I2514);
DFFARX1 I_35458 (I689096,I2507,I605318,I605344,);
not I_35459 (I605352,I605344);
DFFARX1 I_35460 (I689108,I2507,I605318,I605378,);
not I_35461 (I605386,I689099);
nand I_35462 (I605403,I605386,I689102);
not I_35463 (I605420,I605403);
nor I_35464 (I605437,I605420,I689105);
nor I_35465 (I605454,I605352,I605437);
DFFARX1 I_35466 (I605454,I2507,I605318,I605304,);
not I_35467 (I605485,I689105);
nand I_35468 (I605502,I605485,I605420);
and I_35469 (I605519,I605485,I689099);
nand I_35470 (I605536,I605519,I689111);
nor I_35471 (I605301,I605536,I605485);
and I_35472 (I605292,I605378,I605536);
not I_35473 (I605581,I605536);
nand I_35474 (I605295,I605378,I605581);
nor I_35475 (I605289,I605344,I605536);
not I_35476 (I605626,I689117);
nor I_35477 (I605643,I605626,I689099);
nand I_35478 (I605660,I605643,I605485);
nor I_35479 (I605298,I605403,I605660);
nor I_35480 (I605691,I605626,I689096);
and I_35481 (I605708,I605691,I689114);
or I_35482 (I605725,I605708,I689120);
DFFARX1 I_35483 (I605725,I2507,I605318,I605751,);
nor I_35484 (I605759,I605751,I605502);
DFFARX1 I_35485 (I605759,I2507,I605318,I605286,);
DFFARX1 I_35486 (I605751,I2507,I605318,I605310,);
not I_35487 (I605804,I605751);
nor I_35488 (I605821,I605804,I605378);
nor I_35489 (I605838,I605643,I605821);
DFFARX1 I_35490 (I605838,I2507,I605318,I605307,);
not I_35491 (I605896,I2514);
DFFARX1 I_35492 (I304477,I2507,I605896,I605922,);
not I_35493 (I605930,I605922);
DFFARX1 I_35494 (I304492,I2507,I605896,I605956,);
not I_35495 (I605964,I304495);
nand I_35496 (I605981,I605964,I304474);
not I_35497 (I605998,I605981);
nor I_35498 (I606015,I605998,I304498);
nor I_35499 (I606032,I605930,I606015);
DFFARX1 I_35500 (I606032,I2507,I605896,I605882,);
not I_35501 (I606063,I304498);
nand I_35502 (I606080,I606063,I605998);
and I_35503 (I606097,I606063,I304480);
nand I_35504 (I606114,I606097,I304471);
nor I_35505 (I605879,I606114,I606063);
and I_35506 (I605870,I605956,I606114);
not I_35507 (I606159,I606114);
nand I_35508 (I605873,I605956,I606159);
nor I_35509 (I605867,I605922,I606114);
not I_35510 (I606204,I304471);
nor I_35511 (I606221,I606204,I304480);
nand I_35512 (I606238,I606221,I606063);
nor I_35513 (I605876,I605981,I606238);
nor I_35514 (I606269,I606204,I304486);
and I_35515 (I606286,I606269,I304489);
or I_35516 (I606303,I606286,I304483);
DFFARX1 I_35517 (I606303,I2507,I605896,I606329,);
nor I_35518 (I606337,I606329,I606080);
DFFARX1 I_35519 (I606337,I2507,I605896,I605864,);
DFFARX1 I_35520 (I606329,I2507,I605896,I605888,);
not I_35521 (I606382,I606329);
nor I_35522 (I606399,I606382,I605956);
nor I_35523 (I606416,I606221,I606399);
DFFARX1 I_35524 (I606416,I2507,I605896,I605885,);
not I_35525 (I606474,I2514);
DFFARX1 I_35526 (I476795,I2507,I606474,I606500,);
not I_35527 (I606508,I606500);
DFFARX1 I_35528 (I476807,I2507,I606474,I606534,);
not I_35529 (I606542,I476783);
nand I_35530 (I606559,I606542,I476810);
not I_35531 (I606576,I606559);
nor I_35532 (I606593,I606576,I476798);
nor I_35533 (I606610,I606508,I606593);
DFFARX1 I_35534 (I606610,I2507,I606474,I606460,);
not I_35535 (I606641,I476798);
nand I_35536 (I606658,I606641,I606576);
and I_35537 (I606675,I606641,I476783);
nand I_35538 (I606692,I606675,I476786);
nor I_35539 (I606457,I606692,I606641);
and I_35540 (I606448,I606534,I606692);
not I_35541 (I606737,I606692);
nand I_35542 (I606451,I606534,I606737);
nor I_35543 (I606445,I606500,I606692);
not I_35544 (I606782,I476792);
nor I_35545 (I606799,I606782,I476783);
nand I_35546 (I606816,I606799,I606641);
nor I_35547 (I606454,I606559,I606816);
nor I_35548 (I606847,I606782,I476801);
and I_35549 (I606864,I606847,I476789);
or I_35550 (I606881,I606864,I476804);
DFFARX1 I_35551 (I606881,I2507,I606474,I606907,);
nor I_35552 (I606915,I606907,I606658);
DFFARX1 I_35553 (I606915,I2507,I606474,I606442,);
DFFARX1 I_35554 (I606907,I2507,I606474,I606466,);
not I_35555 (I606960,I606907);
nor I_35556 (I606977,I606960,I606534);
nor I_35557 (I606994,I606799,I606977);
DFFARX1 I_35558 (I606994,I2507,I606474,I606463,);
not I_35559 (I607052,I2514);
DFFARX1 I_35560 (I417499,I2507,I607052,I607078,);
not I_35561 (I607086,I607078);
DFFARX1 I_35562 (I417511,I2507,I607052,I607112,);
not I_35563 (I607120,I417487);
nand I_35564 (I607137,I607120,I417514);
not I_35565 (I607154,I607137);
nor I_35566 (I607171,I607154,I417502);
nor I_35567 (I607188,I607086,I607171);
DFFARX1 I_35568 (I607188,I2507,I607052,I607038,);
not I_35569 (I607219,I417502);
nand I_35570 (I607236,I607219,I607154);
and I_35571 (I607253,I607219,I417487);
nand I_35572 (I607270,I607253,I417490);
nor I_35573 (I607035,I607270,I607219);
and I_35574 (I607026,I607112,I607270);
not I_35575 (I607315,I607270);
nand I_35576 (I607029,I607112,I607315);
nor I_35577 (I607023,I607078,I607270);
not I_35578 (I607360,I417496);
nor I_35579 (I607377,I607360,I417487);
nand I_35580 (I607394,I607377,I607219);
nor I_35581 (I607032,I607137,I607394);
nor I_35582 (I607425,I607360,I417505);
and I_35583 (I607442,I607425,I417493);
or I_35584 (I607459,I607442,I417508);
DFFARX1 I_35585 (I607459,I2507,I607052,I607485,);
nor I_35586 (I607493,I607485,I607236);
DFFARX1 I_35587 (I607493,I2507,I607052,I607020,);
DFFARX1 I_35588 (I607485,I2507,I607052,I607044,);
not I_35589 (I607538,I607485);
nor I_35590 (I607555,I607538,I607112);
nor I_35591 (I607572,I607377,I607555);
DFFARX1 I_35592 (I607572,I2507,I607052,I607041,);
not I_35593 (I607630,I2514);
DFFARX1 I_35594 (I1204026,I2507,I607630,I607656,);
not I_35595 (I607664,I607656);
DFFARX1 I_35596 (I1204032,I2507,I607630,I607690,);
not I_35597 (I607698,I1204026);
nand I_35598 (I607715,I607698,I1204029);
not I_35599 (I607732,I607715);
nor I_35600 (I607749,I607732,I1204047);
nor I_35601 (I607766,I607664,I607749);
DFFARX1 I_35602 (I607766,I2507,I607630,I607616,);
not I_35603 (I607797,I1204047);
nand I_35604 (I607814,I607797,I607732);
and I_35605 (I607831,I607797,I1204050);
nand I_35606 (I607848,I607831,I1204029);
nor I_35607 (I607613,I607848,I607797);
and I_35608 (I607604,I607690,I607848);
not I_35609 (I607893,I607848);
nand I_35610 (I607607,I607690,I607893);
nor I_35611 (I607601,I607656,I607848);
not I_35612 (I607938,I1204035);
nor I_35613 (I607955,I607938,I1204050);
nand I_35614 (I607972,I607955,I607797);
nor I_35615 (I607610,I607715,I607972);
nor I_35616 (I608003,I607938,I1204041);
and I_35617 (I608020,I608003,I1204038);
or I_35618 (I608037,I608020,I1204044);
DFFARX1 I_35619 (I608037,I2507,I607630,I608063,);
nor I_35620 (I608071,I608063,I607814);
DFFARX1 I_35621 (I608071,I2507,I607630,I607598,);
DFFARX1 I_35622 (I608063,I2507,I607630,I607622,);
not I_35623 (I608116,I608063);
nor I_35624 (I608133,I608116,I607690);
nor I_35625 (I608150,I607955,I608133);
DFFARX1 I_35626 (I608150,I2507,I607630,I607619,);
not I_35627 (I608208,I2514);
DFFARX1 I_35628 (I842306,I2507,I608208,I608234,);
not I_35629 (I608242,I608234);
DFFARX1 I_35630 (I842306,I2507,I608208,I608268,);
not I_35631 (I608276,I842303);
nand I_35632 (I608293,I608276,I842318);
not I_35633 (I608310,I608293);
nor I_35634 (I608327,I608310,I842312);
nor I_35635 (I608344,I608242,I608327);
DFFARX1 I_35636 (I608344,I2507,I608208,I608194,);
not I_35637 (I608375,I842312);
nand I_35638 (I608392,I608375,I608310);
and I_35639 (I608409,I608375,I842309);
nand I_35640 (I608426,I608409,I842300);
nor I_35641 (I608191,I608426,I608375);
and I_35642 (I608182,I608268,I608426);
not I_35643 (I608471,I608426);
nand I_35644 (I608185,I608268,I608471);
nor I_35645 (I608179,I608234,I608426);
not I_35646 (I608516,I842321);
nor I_35647 (I608533,I608516,I842309);
nand I_35648 (I608550,I608533,I608375);
nor I_35649 (I608188,I608293,I608550);
nor I_35650 (I608581,I608516,I842300);
and I_35651 (I608598,I608581,I842303);
or I_35652 (I608615,I608598,I842315);
DFFARX1 I_35653 (I608615,I2507,I608208,I608641,);
nor I_35654 (I608649,I608641,I608392);
DFFARX1 I_35655 (I608649,I2507,I608208,I608176,);
DFFARX1 I_35656 (I608641,I2507,I608208,I608200,);
not I_35657 (I608694,I608641);
nor I_35658 (I608711,I608694,I608268);
nor I_35659 (I608728,I608533,I608711);
DFFARX1 I_35660 (I608728,I2507,I608208,I608197,);
not I_35661 (I608786,I2514);
DFFARX1 I_35662 (I1078022,I2507,I608786,I608812,);
not I_35663 (I608820,I608812);
DFFARX1 I_35664 (I1078028,I2507,I608786,I608846,);
not I_35665 (I608854,I1078022);
nand I_35666 (I608871,I608854,I1078025);
not I_35667 (I608888,I608871);
nor I_35668 (I608905,I608888,I1078043);
nor I_35669 (I608922,I608820,I608905);
DFFARX1 I_35670 (I608922,I2507,I608786,I608772,);
not I_35671 (I608953,I1078043);
nand I_35672 (I608970,I608953,I608888);
and I_35673 (I608987,I608953,I1078046);
nand I_35674 (I609004,I608987,I1078025);
nor I_35675 (I608769,I609004,I608953);
and I_35676 (I608760,I608846,I609004);
not I_35677 (I609049,I609004);
nand I_35678 (I608763,I608846,I609049);
nor I_35679 (I608757,I608812,I609004);
not I_35680 (I609094,I1078031);
nor I_35681 (I609111,I609094,I1078046);
nand I_35682 (I609128,I609111,I608953);
nor I_35683 (I608766,I608871,I609128);
nor I_35684 (I609159,I609094,I1078037);
and I_35685 (I609176,I609159,I1078034);
or I_35686 (I609193,I609176,I1078040);
DFFARX1 I_35687 (I609193,I2507,I608786,I609219,);
nor I_35688 (I609227,I609219,I608970);
DFFARX1 I_35689 (I609227,I2507,I608786,I608754,);
DFFARX1 I_35690 (I609219,I2507,I608786,I608778,);
not I_35691 (I609272,I609219);
nor I_35692 (I609289,I609272,I608846);
nor I_35693 (I609306,I609111,I609289);
DFFARX1 I_35694 (I609306,I2507,I608786,I608775,);
not I_35695 (I609364,I2514);
DFFARX1 I_35696 (I51195,I2507,I609364,I609390,);
not I_35697 (I609398,I609390);
DFFARX1 I_35698 (I51174,I2507,I609364,I609424,);
not I_35699 (I609432,I51171);
nand I_35700 (I609449,I609432,I51186);
not I_35701 (I609466,I609449);
nor I_35702 (I609483,I609466,I51174);
nor I_35703 (I609500,I609398,I609483);
DFFARX1 I_35704 (I609500,I2507,I609364,I609350,);
not I_35705 (I609531,I51174);
nand I_35706 (I609548,I609531,I609466);
and I_35707 (I609565,I609531,I51177);
nand I_35708 (I609582,I609565,I51192);
nor I_35709 (I609347,I609582,I609531);
and I_35710 (I609338,I609424,I609582);
not I_35711 (I609627,I609582);
nand I_35712 (I609341,I609424,I609627);
nor I_35713 (I609335,I609390,I609582);
not I_35714 (I609672,I51183);
nor I_35715 (I609689,I609672,I51177);
nand I_35716 (I609706,I609689,I609531);
nor I_35717 (I609344,I609449,I609706);
nor I_35718 (I609737,I609672,I51171);
and I_35719 (I609754,I609737,I51180);
or I_35720 (I609771,I609754,I51189);
DFFARX1 I_35721 (I609771,I2507,I609364,I609797,);
nor I_35722 (I609805,I609797,I609548);
DFFARX1 I_35723 (I609805,I2507,I609364,I609332,);
DFFARX1 I_35724 (I609797,I2507,I609364,I609356,);
not I_35725 (I609850,I609797);
nor I_35726 (I609867,I609850,I609424);
nor I_35727 (I609884,I609689,I609867);
DFFARX1 I_35728 (I609884,I2507,I609364,I609353,);
not I_35729 (I609942,I2514);
DFFARX1 I_35730 (I110219,I2507,I609942,I609968,);
not I_35731 (I609976,I609968);
DFFARX1 I_35732 (I110198,I2507,I609942,I610002,);
not I_35733 (I610010,I110195);
nand I_35734 (I610027,I610010,I110210);
not I_35735 (I610044,I610027);
nor I_35736 (I610061,I610044,I110198);
nor I_35737 (I610078,I609976,I610061);
DFFARX1 I_35738 (I610078,I2507,I609942,I609928,);
not I_35739 (I610109,I110198);
nand I_35740 (I610126,I610109,I610044);
and I_35741 (I610143,I610109,I110201);
nand I_35742 (I610160,I610143,I110216);
nor I_35743 (I609925,I610160,I610109);
and I_35744 (I609916,I610002,I610160);
not I_35745 (I610205,I610160);
nand I_35746 (I609919,I610002,I610205);
nor I_35747 (I609913,I609968,I610160);
not I_35748 (I610250,I110207);
nor I_35749 (I610267,I610250,I110201);
nand I_35750 (I610284,I610267,I610109);
nor I_35751 (I609922,I610027,I610284);
nor I_35752 (I610315,I610250,I110195);
and I_35753 (I610332,I610315,I110204);
or I_35754 (I610349,I610332,I110213);
DFFARX1 I_35755 (I610349,I2507,I609942,I610375,);
nor I_35756 (I610383,I610375,I610126);
DFFARX1 I_35757 (I610383,I2507,I609942,I609910,);
DFFARX1 I_35758 (I610375,I2507,I609942,I609934,);
not I_35759 (I610428,I610375);
nor I_35760 (I610445,I610428,I610002);
nor I_35761 (I610462,I610267,I610445);
DFFARX1 I_35762 (I610462,I2507,I609942,I609931,);
not I_35763 (I610520,I2514);
DFFARX1 I_35764 (I295518,I2507,I610520,I610546,);
not I_35765 (I610554,I610546);
DFFARX1 I_35766 (I295533,I2507,I610520,I610580,);
not I_35767 (I610588,I295536);
nand I_35768 (I610605,I610588,I295515);
not I_35769 (I610622,I610605);
nor I_35770 (I610639,I610622,I295539);
nor I_35771 (I610656,I610554,I610639);
DFFARX1 I_35772 (I610656,I2507,I610520,I610506,);
not I_35773 (I610687,I295539);
nand I_35774 (I610704,I610687,I610622);
and I_35775 (I610721,I610687,I295521);
nand I_35776 (I610738,I610721,I295512);
nor I_35777 (I610503,I610738,I610687);
and I_35778 (I610494,I610580,I610738);
not I_35779 (I610783,I610738);
nand I_35780 (I610497,I610580,I610783);
nor I_35781 (I610491,I610546,I610738);
not I_35782 (I610828,I295512);
nor I_35783 (I610845,I610828,I295521);
nand I_35784 (I610862,I610845,I610687);
nor I_35785 (I610500,I610605,I610862);
nor I_35786 (I610893,I610828,I295527);
and I_35787 (I610910,I610893,I295530);
or I_35788 (I610927,I610910,I295524);
DFFARX1 I_35789 (I610927,I2507,I610520,I610953,);
nor I_35790 (I610961,I610953,I610704);
DFFARX1 I_35791 (I610961,I2507,I610520,I610488,);
DFFARX1 I_35792 (I610953,I2507,I610520,I610512,);
not I_35793 (I611006,I610953);
nor I_35794 (I611023,I611006,I610580);
nor I_35795 (I611040,I610845,I611023);
DFFARX1 I_35796 (I611040,I2507,I610520,I610509,);
not I_35797 (I611098,I2514);
DFFARX1 I_35798 (I630718,I2507,I611098,I611124,);
not I_35799 (I611132,I611124);
DFFARX1 I_35800 (I630730,I2507,I611098,I611158,);
not I_35801 (I611166,I630721);
nand I_35802 (I611183,I611166,I630724);
not I_35803 (I611200,I611183);
nor I_35804 (I611217,I611200,I630727);
nor I_35805 (I611234,I611132,I611217);
DFFARX1 I_35806 (I611234,I2507,I611098,I611084,);
not I_35807 (I611265,I630727);
nand I_35808 (I611282,I611265,I611200);
and I_35809 (I611299,I611265,I630721);
nand I_35810 (I611316,I611299,I630733);
nor I_35811 (I611081,I611316,I611265);
and I_35812 (I611072,I611158,I611316);
not I_35813 (I611361,I611316);
nand I_35814 (I611075,I611158,I611361);
nor I_35815 (I611069,I611124,I611316);
not I_35816 (I611406,I630739);
nor I_35817 (I611423,I611406,I630721);
nand I_35818 (I611440,I611423,I611265);
nor I_35819 (I611078,I611183,I611440);
nor I_35820 (I611471,I611406,I630718);
and I_35821 (I611488,I611471,I630736);
or I_35822 (I611505,I611488,I630742);
DFFARX1 I_35823 (I611505,I2507,I611098,I611531,);
nor I_35824 (I611539,I611531,I611282);
DFFARX1 I_35825 (I611539,I2507,I611098,I611066,);
DFFARX1 I_35826 (I611531,I2507,I611098,I611090,);
not I_35827 (I611584,I611531);
nor I_35828 (I611601,I611584,I611158);
nor I_35829 (I611618,I611423,I611601);
DFFARX1 I_35830 (I611618,I2507,I611098,I611087,);
not I_35831 (I611676,I2514);
DFFARX1 I_35832 (I1283666,I2507,I611676,I611702,);
not I_35833 (I611710,I611702);
DFFARX1 I_35834 (I1283678,I2507,I611676,I611736,);
not I_35835 (I611744,I1283669);
nand I_35836 (I611761,I611744,I1283657);
not I_35837 (I611778,I611761);
nor I_35838 (I611795,I611778,I1283654);
nor I_35839 (I611812,I611710,I611795);
DFFARX1 I_35840 (I611812,I2507,I611676,I611662,);
not I_35841 (I611843,I1283654);
nand I_35842 (I611860,I611843,I611778);
and I_35843 (I611877,I611843,I1283660);
nand I_35844 (I611894,I611877,I1283657);
nor I_35845 (I611659,I611894,I611843);
and I_35846 (I611650,I611736,I611894);
not I_35847 (I611939,I611894);
nand I_35848 (I611653,I611736,I611939);
nor I_35849 (I611647,I611702,I611894);
not I_35850 (I611984,I1283675);
nor I_35851 (I612001,I611984,I1283660);
nand I_35852 (I612018,I612001,I611843);
nor I_35853 (I611656,I611761,I612018);
nor I_35854 (I612049,I611984,I1283663);
and I_35855 (I612066,I612049,I1283654);
or I_35856 (I612083,I612066,I1283672);
DFFARX1 I_35857 (I612083,I2507,I611676,I612109,);
nor I_35858 (I612117,I612109,I611860);
DFFARX1 I_35859 (I612117,I2507,I611676,I611644,);
DFFARX1 I_35860 (I612109,I2507,I611676,I611668,);
not I_35861 (I612162,I612109);
nor I_35862 (I612179,I612162,I611736);
nor I_35863 (I612196,I612001,I612179);
DFFARX1 I_35864 (I612196,I2507,I611676,I611665,);
not I_35865 (I612254,I2514);
DFFARX1 I_35866 (I1370167,I2507,I612254,I612280,);
not I_35867 (I612288,I612280);
DFFARX1 I_35868 (I1370167,I2507,I612254,I612314,);
not I_35869 (I612322,I1370191);
nand I_35870 (I612339,I612322,I1370173);
not I_35871 (I612356,I612339);
nor I_35872 (I612373,I612356,I1370188);
nor I_35873 (I612390,I612288,I612373);
DFFARX1 I_35874 (I612390,I2507,I612254,I612240,);
not I_35875 (I612421,I1370188);
nand I_35876 (I612438,I612421,I612356);
and I_35877 (I612455,I612421,I1370170);
nand I_35878 (I612472,I612455,I1370179);
nor I_35879 (I612237,I612472,I612421);
and I_35880 (I612228,I612314,I612472);
not I_35881 (I612517,I612472);
nand I_35882 (I612231,I612314,I612517);
nor I_35883 (I612225,I612280,I612472);
not I_35884 (I612562,I1370176);
nor I_35885 (I612579,I612562,I1370170);
nand I_35886 (I612596,I612579,I612421);
nor I_35887 (I612234,I612339,I612596);
nor I_35888 (I612627,I612562,I1370185);
and I_35889 (I612644,I612627,I1370194);
or I_35890 (I612661,I612644,I1370182);
DFFARX1 I_35891 (I612661,I2507,I612254,I612687,);
nor I_35892 (I612695,I612687,I612438);
DFFARX1 I_35893 (I612695,I2507,I612254,I612222,);
DFFARX1 I_35894 (I612687,I2507,I612254,I612246,);
not I_35895 (I612740,I612687);
nor I_35896 (I612757,I612740,I612314);
nor I_35897 (I612774,I612579,I612757);
DFFARX1 I_35898 (I612774,I2507,I612254,I612243,);
not I_35899 (I612832,I2514);
DFFARX1 I_35900 (I1048310,I2507,I612832,I612858,);
not I_35901 (I612866,I612858);
DFFARX1 I_35902 (I1048301,I2507,I612832,I612892,);
not I_35903 (I612900,I1048295);
nand I_35904 (I612917,I612900,I1048307);
not I_35905 (I612934,I612917);
nor I_35906 (I612951,I612934,I1048298);
nor I_35907 (I612968,I612866,I612951);
DFFARX1 I_35908 (I612968,I2507,I612832,I612818,);
not I_35909 (I612999,I1048298);
nand I_35910 (I613016,I612999,I612934);
and I_35911 (I613033,I612999,I1048304);
nand I_35912 (I613050,I613033,I1048289);
nor I_35913 (I612815,I613050,I612999);
and I_35914 (I612806,I612892,I613050);
not I_35915 (I613095,I613050);
nand I_35916 (I612809,I612892,I613095);
nor I_35917 (I612803,I612858,I613050);
not I_35918 (I613140,I1048289);
nor I_35919 (I613157,I613140,I1048304);
nand I_35920 (I613174,I613157,I612999);
nor I_35921 (I612812,I612917,I613174);
nor I_35922 (I613205,I613140,I1048292);
and I_35923 (I613222,I613205,I1048295);
or I_35924 (I613239,I613222,I1048292);
DFFARX1 I_35925 (I613239,I2507,I612832,I613265,);
nor I_35926 (I613273,I613265,I613016);
DFFARX1 I_35927 (I613273,I2507,I612832,I612800,);
DFFARX1 I_35928 (I613265,I2507,I612832,I612824,);
not I_35929 (I613318,I613265);
nor I_35930 (I613335,I613318,I612892);
nor I_35931 (I613352,I613157,I613335);
DFFARX1 I_35932 (I613352,I2507,I612832,I612821,);
not I_35933 (I613410,I2514);
DFFARX1 I_35934 (I1169924,I2507,I613410,I613436,);
not I_35935 (I613444,I613436);
DFFARX1 I_35936 (I1169930,I2507,I613410,I613470,);
not I_35937 (I613478,I1169924);
nand I_35938 (I613495,I613478,I1169927);
not I_35939 (I613512,I613495);
nor I_35940 (I613529,I613512,I1169945);
nor I_35941 (I613546,I613444,I613529);
DFFARX1 I_35942 (I613546,I2507,I613410,I613396,);
not I_35943 (I613577,I1169945);
nand I_35944 (I613594,I613577,I613512);
and I_35945 (I613611,I613577,I1169948);
nand I_35946 (I613628,I613611,I1169927);
nor I_35947 (I613393,I613628,I613577);
and I_35948 (I613384,I613470,I613628);
not I_35949 (I613673,I613628);
nand I_35950 (I613387,I613470,I613673);
nor I_35951 (I613381,I613436,I613628);
not I_35952 (I613718,I1169933);
nor I_35953 (I613735,I613718,I1169948);
nand I_35954 (I613752,I613735,I613577);
nor I_35955 (I613390,I613495,I613752);
nor I_35956 (I613783,I613718,I1169939);
and I_35957 (I613800,I613783,I1169936);
or I_35958 (I613817,I613800,I1169942);
DFFARX1 I_35959 (I613817,I2507,I613410,I613843,);
nor I_35960 (I613851,I613843,I613594);
DFFARX1 I_35961 (I613851,I2507,I613410,I613378,);
DFFARX1 I_35962 (I613843,I2507,I613410,I613402,);
not I_35963 (I613896,I613843);
nor I_35964 (I613913,I613896,I613470);
nor I_35965 (I613930,I613735,I613913);
DFFARX1 I_35966 (I613930,I2507,I613410,I613399,);
not I_35967 (I613988,I2514);
DFFARX1 I_35968 (I488763,I2507,I613988,I614014,);
not I_35969 (I614022,I614014);
DFFARX1 I_35970 (I488775,I2507,I613988,I614048,);
not I_35971 (I614056,I488751);
nand I_35972 (I614073,I614056,I488778);
not I_35973 (I614090,I614073);
nor I_35974 (I614107,I614090,I488766);
nor I_35975 (I614124,I614022,I614107);
DFFARX1 I_35976 (I614124,I2507,I613988,I613974,);
not I_35977 (I614155,I488766);
nand I_35978 (I614172,I614155,I614090);
and I_35979 (I614189,I614155,I488751);
nand I_35980 (I614206,I614189,I488754);
nor I_35981 (I613971,I614206,I614155);
and I_35982 (I613962,I614048,I614206);
not I_35983 (I614251,I614206);
nand I_35984 (I613965,I614048,I614251);
nor I_35985 (I613959,I614014,I614206);
not I_35986 (I614296,I488760);
nor I_35987 (I614313,I614296,I488751);
nand I_35988 (I614330,I614313,I614155);
nor I_35989 (I613968,I614073,I614330);
nor I_35990 (I614361,I614296,I488769);
and I_35991 (I614378,I614361,I488757);
or I_35992 (I614395,I614378,I488772);
DFFARX1 I_35993 (I614395,I2507,I613988,I614421,);
nor I_35994 (I614429,I614421,I614172);
DFFARX1 I_35995 (I614429,I2507,I613988,I613956,);
DFFARX1 I_35996 (I614421,I2507,I613988,I613980,);
not I_35997 (I614474,I614421);
nor I_35998 (I614491,I614474,I614048);
nor I_35999 (I614508,I614313,I614491);
DFFARX1 I_36000 (I614508,I2507,I613988,I613977,);
not I_36001 (I614566,I2514);
DFFARX1 I_36002 (I307639,I2507,I614566,I614592,);
not I_36003 (I614600,I614592);
DFFARX1 I_36004 (I307654,I2507,I614566,I614626,);
not I_36005 (I614634,I307657);
nand I_36006 (I614651,I614634,I307636);
not I_36007 (I614668,I614651);
nor I_36008 (I614685,I614668,I307660);
nor I_36009 (I614702,I614600,I614685);
DFFARX1 I_36010 (I614702,I2507,I614566,I614552,);
not I_36011 (I614733,I307660);
nand I_36012 (I614750,I614733,I614668);
and I_36013 (I614767,I614733,I307642);
nand I_36014 (I614784,I614767,I307633);
nor I_36015 (I614549,I614784,I614733);
and I_36016 (I614540,I614626,I614784);
not I_36017 (I614829,I614784);
nand I_36018 (I614543,I614626,I614829);
nor I_36019 (I614537,I614592,I614784);
not I_36020 (I614874,I307633);
nor I_36021 (I614891,I614874,I307642);
nand I_36022 (I614908,I614891,I614733);
nor I_36023 (I614546,I614651,I614908);
nor I_36024 (I614939,I614874,I307648);
and I_36025 (I614956,I614939,I307651);
or I_36026 (I614973,I614956,I307645);
DFFARX1 I_36027 (I614973,I2507,I614566,I614999,);
nor I_36028 (I615007,I614999,I614750);
DFFARX1 I_36029 (I615007,I2507,I614566,I614534,);
DFFARX1 I_36030 (I614999,I2507,I614566,I614558,);
not I_36031 (I615052,I614999);
nor I_36032 (I615069,I615052,I614626);
nor I_36033 (I615086,I614891,I615069);
DFFARX1 I_36034 (I615086,I2507,I614566,I614555,);
not I_36035 (I615144,I2514);
DFFARX1 I_36036 (I954761,I2507,I615144,I615170,);
not I_36037 (I615178,I615170);
DFFARX1 I_36038 (I954758,I2507,I615144,I615204,);
not I_36039 (I615212,I954755);
nand I_36040 (I615229,I615212,I954782);
not I_36041 (I615246,I615229);
nor I_36042 (I615263,I615246,I954770);
nor I_36043 (I615280,I615178,I615263);
DFFARX1 I_36044 (I615280,I2507,I615144,I615130,);
not I_36045 (I615311,I954770);
nand I_36046 (I615328,I615311,I615246);
and I_36047 (I615345,I615311,I954776);
nand I_36048 (I615362,I615345,I954767);
nor I_36049 (I615127,I615362,I615311);
and I_36050 (I615118,I615204,I615362);
not I_36051 (I615407,I615362);
nand I_36052 (I615121,I615204,I615407);
nor I_36053 (I615115,I615170,I615362);
not I_36054 (I615452,I954764);
nor I_36055 (I615469,I615452,I954776);
nand I_36056 (I615486,I615469,I615311);
nor I_36057 (I615124,I615229,I615486);
nor I_36058 (I615517,I615452,I954779);
and I_36059 (I615534,I615517,I954773);
or I_36060 (I615551,I615534,I954755);
DFFARX1 I_36061 (I615551,I2507,I615144,I615577,);
nor I_36062 (I615585,I615577,I615328);
DFFARX1 I_36063 (I615585,I2507,I615144,I615112,);
DFFARX1 I_36064 (I615577,I2507,I615144,I615136,);
not I_36065 (I615630,I615577);
nor I_36066 (I615647,I615630,I615204);
nor I_36067 (I615664,I615469,I615647);
DFFARX1 I_36068 (I615664,I2507,I615144,I615133,);
not I_36069 (I615722,I2514);
DFFARX1 I_36070 (I1389207,I2507,I615722,I615748,);
not I_36071 (I615756,I615748);
DFFARX1 I_36072 (I1389207,I2507,I615722,I615782,);
not I_36073 (I615790,I1389231);
nand I_36074 (I615807,I615790,I1389213);
not I_36075 (I615824,I615807);
nor I_36076 (I615841,I615824,I1389228);
nor I_36077 (I615858,I615756,I615841);
DFFARX1 I_36078 (I615858,I2507,I615722,I615708,);
not I_36079 (I615889,I1389228);
nand I_36080 (I615906,I615889,I615824);
and I_36081 (I615923,I615889,I1389210);
nand I_36082 (I615940,I615923,I1389219);
nor I_36083 (I615705,I615940,I615889);
and I_36084 (I615696,I615782,I615940);
not I_36085 (I615985,I615940);
nand I_36086 (I615699,I615782,I615985);
nor I_36087 (I615693,I615748,I615940);
not I_36088 (I616030,I1389216);
nor I_36089 (I616047,I616030,I1389210);
nand I_36090 (I616064,I616047,I615889);
nor I_36091 (I615702,I615807,I616064);
nor I_36092 (I616095,I616030,I1389225);
and I_36093 (I616112,I616095,I1389234);
or I_36094 (I616129,I616112,I1389222);
DFFARX1 I_36095 (I616129,I2507,I615722,I616155,);
nor I_36096 (I616163,I616155,I615906);
DFFARX1 I_36097 (I616163,I2507,I615722,I615690,);
DFFARX1 I_36098 (I616155,I2507,I615722,I615714,);
not I_36099 (I616208,I616155);
nor I_36100 (I616225,I616208,I615782);
nor I_36101 (I616242,I616047,I616225);
DFFARX1 I_36102 (I616242,I2507,I615722,I615711,);
not I_36103 (I616300,I2514);
DFFARX1 I_36104 (I433819,I2507,I616300,I616326,);
not I_36105 (I616334,I616326);
DFFARX1 I_36106 (I433831,I2507,I616300,I616360,);
not I_36107 (I616368,I433807);
nand I_36108 (I616385,I616368,I433834);
not I_36109 (I616402,I616385);
nor I_36110 (I616419,I616402,I433822);
nor I_36111 (I616436,I616334,I616419);
DFFARX1 I_36112 (I616436,I2507,I616300,I616286,);
not I_36113 (I616467,I433822);
nand I_36114 (I616484,I616467,I616402);
and I_36115 (I616501,I616467,I433807);
nand I_36116 (I616518,I616501,I433810);
nor I_36117 (I616283,I616518,I616467);
and I_36118 (I616274,I616360,I616518);
not I_36119 (I616563,I616518);
nand I_36120 (I616277,I616360,I616563);
nor I_36121 (I616271,I616326,I616518);
not I_36122 (I616608,I433816);
nor I_36123 (I616625,I616608,I433807);
nand I_36124 (I616642,I616625,I616467);
nor I_36125 (I616280,I616385,I616642);
nor I_36126 (I616673,I616608,I433825);
and I_36127 (I616690,I616673,I433813);
or I_36128 (I616707,I616690,I433828);
DFFARX1 I_36129 (I616707,I2507,I616300,I616733,);
nor I_36130 (I616741,I616733,I616484);
DFFARX1 I_36131 (I616741,I2507,I616300,I616268,);
DFFARX1 I_36132 (I616733,I2507,I616300,I616292,);
not I_36133 (I616786,I616733);
nor I_36134 (I616803,I616786,I616360);
nor I_36135 (I616820,I616625,I616803);
DFFARX1 I_36136 (I616820,I2507,I616300,I616289,);
not I_36137 (I616878,I2514);
DFFARX1 I_36138 (I1041578,I2507,I616878,I616904,);
not I_36139 (I616912,I616904);
DFFARX1 I_36140 (I1041569,I2507,I616878,I616938,);
not I_36141 (I616946,I1041563);
nand I_36142 (I616963,I616946,I1041575);
not I_36143 (I616980,I616963);
nor I_36144 (I616997,I616980,I1041566);
nor I_36145 (I617014,I616912,I616997);
DFFARX1 I_36146 (I617014,I2507,I616878,I616864,);
not I_36147 (I617045,I1041566);
nand I_36148 (I617062,I617045,I616980);
and I_36149 (I617079,I617045,I1041572);
nand I_36150 (I617096,I617079,I1041557);
nor I_36151 (I616861,I617096,I617045);
and I_36152 (I616852,I616938,I617096);
not I_36153 (I617141,I617096);
nand I_36154 (I616855,I616938,I617141);
nor I_36155 (I616849,I616904,I617096);
not I_36156 (I617186,I1041557);
nor I_36157 (I617203,I617186,I1041572);
nand I_36158 (I617220,I617203,I617045);
nor I_36159 (I616858,I616963,I617220);
nor I_36160 (I617251,I617186,I1041560);
and I_36161 (I617268,I617251,I1041563);
or I_36162 (I617285,I617268,I1041560);
DFFARX1 I_36163 (I617285,I2507,I616878,I617311,);
nor I_36164 (I617319,I617311,I617062);
DFFARX1 I_36165 (I617319,I2507,I616878,I616846,);
DFFARX1 I_36166 (I617311,I2507,I616878,I616870,);
not I_36167 (I617364,I617311);
nor I_36168 (I617381,I617364,I616938);
nor I_36169 (I617398,I617203,I617381);
DFFARX1 I_36170 (I617398,I2507,I616878,I616867,);
not I_36171 (I617456,I2514);
DFFARX1 I_36172 (I647480,I2507,I617456,I617482,);
not I_36173 (I617490,I617482);
DFFARX1 I_36174 (I647492,I2507,I617456,I617516,);
not I_36175 (I617524,I647483);
nand I_36176 (I617541,I617524,I647486);
not I_36177 (I617558,I617541);
nor I_36178 (I617575,I617558,I647489);
nor I_36179 (I617592,I617490,I617575);
DFFARX1 I_36180 (I617592,I2507,I617456,I617442,);
not I_36181 (I617623,I647489);
nand I_36182 (I617640,I617623,I617558);
and I_36183 (I617657,I617623,I647483);
nand I_36184 (I617674,I617657,I647495);
nor I_36185 (I617439,I617674,I617623);
and I_36186 (I617430,I617516,I617674);
not I_36187 (I617719,I617674);
nand I_36188 (I617433,I617516,I617719);
nor I_36189 (I617427,I617482,I617674);
not I_36190 (I617764,I647501);
nor I_36191 (I617781,I617764,I647483);
nand I_36192 (I617798,I617781,I617623);
nor I_36193 (I617436,I617541,I617798);
nor I_36194 (I617829,I617764,I647480);
and I_36195 (I617846,I617829,I647498);
or I_36196 (I617863,I617846,I647504);
DFFARX1 I_36197 (I617863,I2507,I617456,I617889,);
nor I_36198 (I617897,I617889,I617640);
DFFARX1 I_36199 (I617897,I2507,I617456,I617424,);
DFFARX1 I_36200 (I617889,I2507,I617456,I617448,);
not I_36201 (I617942,I617889);
nor I_36202 (I617959,I617942,I617516);
nor I_36203 (I617976,I617781,I617959);
DFFARX1 I_36204 (I617976,I2507,I617456,I617445,);
not I_36205 (I618034,I2514);
DFFARX1 I_36206 (I732446,I2507,I618034,I618060,);
not I_36207 (I618068,I618060);
DFFARX1 I_36208 (I732458,I2507,I618034,I618094,);
not I_36209 (I618102,I732449);
nand I_36210 (I618119,I618102,I732452);
not I_36211 (I618136,I618119);
nor I_36212 (I618153,I618136,I732455);
nor I_36213 (I618170,I618068,I618153);
DFFARX1 I_36214 (I618170,I2507,I618034,I618020,);
not I_36215 (I618201,I732455);
nand I_36216 (I618218,I618201,I618136);
and I_36217 (I618235,I618201,I732449);
nand I_36218 (I618252,I618235,I732461);
nor I_36219 (I618017,I618252,I618201);
and I_36220 (I618008,I618094,I618252);
not I_36221 (I618297,I618252);
nand I_36222 (I618011,I618094,I618297);
nor I_36223 (I618005,I618060,I618252);
not I_36224 (I618342,I732467);
nor I_36225 (I618359,I618342,I732449);
nand I_36226 (I618376,I618359,I618201);
nor I_36227 (I618014,I618119,I618376);
nor I_36228 (I618407,I618342,I732446);
and I_36229 (I618424,I618407,I732464);
or I_36230 (I618441,I618424,I732470);
DFFARX1 I_36231 (I618441,I2507,I618034,I618467,);
nor I_36232 (I618475,I618467,I618218);
DFFARX1 I_36233 (I618475,I2507,I618034,I618002,);
DFFARX1 I_36234 (I618467,I2507,I618034,I618026,);
not I_36235 (I618520,I618467);
nor I_36236 (I618537,I618520,I618094);
nor I_36237 (I618554,I618359,I618537);
DFFARX1 I_36238 (I618554,I2507,I618034,I618023,);
not I_36239 (I618612,I2514);
DFFARX1 I_36240 (I199035,I2507,I618612,I618638,);
not I_36241 (I618646,I618638);
DFFARX1 I_36242 (I199020,I2507,I618612,I618672,);
not I_36243 (I618680,I199038);
nand I_36244 (I618697,I618680,I199023);
not I_36245 (I618714,I618697);
nor I_36246 (I618731,I618714,I199020);
nor I_36247 (I618748,I618646,I618731);
DFFARX1 I_36248 (I618748,I2507,I618612,I618598,);
not I_36249 (I618779,I199020);
nand I_36250 (I618796,I618779,I618714);
and I_36251 (I618813,I618779,I199023);
nand I_36252 (I618830,I618813,I199044);
nor I_36253 (I618595,I618830,I618779);
and I_36254 (I618586,I618672,I618830);
not I_36255 (I618875,I618830);
nand I_36256 (I618589,I618672,I618875);
nor I_36257 (I618583,I618638,I618830);
not I_36258 (I618920,I199032);
nor I_36259 (I618937,I618920,I199023);
nand I_36260 (I618954,I618937,I618779);
nor I_36261 (I618592,I618697,I618954);
nor I_36262 (I618985,I618920,I199026);
and I_36263 (I619002,I618985,I199041);
or I_36264 (I619019,I619002,I199029);
DFFARX1 I_36265 (I619019,I2507,I618612,I619045,);
nor I_36266 (I619053,I619045,I618796);
DFFARX1 I_36267 (I619053,I2507,I618612,I618580,);
DFFARX1 I_36268 (I619045,I2507,I618612,I618604,);
not I_36269 (I619098,I619045);
nor I_36270 (I619115,I619098,I618672);
nor I_36271 (I619132,I618937,I619115);
DFFARX1 I_36272 (I619132,I2507,I618612,I618601,);
not I_36273 (I619190,I2514);
DFFARX1 I_36274 (I427291,I2507,I619190,I619216,);
not I_36275 (I619224,I619216);
DFFARX1 I_36276 (I427303,I2507,I619190,I619250,);
not I_36277 (I619258,I427279);
nand I_36278 (I619275,I619258,I427306);
not I_36279 (I619292,I619275);
nor I_36280 (I619309,I619292,I427294);
nor I_36281 (I619326,I619224,I619309);
DFFARX1 I_36282 (I619326,I2507,I619190,I619176,);
not I_36283 (I619357,I427294);
nand I_36284 (I619374,I619357,I619292);
and I_36285 (I619391,I619357,I427279);
nand I_36286 (I619408,I619391,I427282);
nor I_36287 (I619173,I619408,I619357);
and I_36288 (I619164,I619250,I619408);
not I_36289 (I619453,I619408);
nand I_36290 (I619167,I619250,I619453);
nor I_36291 (I619161,I619216,I619408);
not I_36292 (I619498,I427288);
nor I_36293 (I619515,I619498,I427279);
nand I_36294 (I619532,I619515,I619357);
nor I_36295 (I619170,I619275,I619532);
nor I_36296 (I619563,I619498,I427297);
and I_36297 (I619580,I619563,I427285);
or I_36298 (I619597,I619580,I427300);
DFFARX1 I_36299 (I619597,I2507,I619190,I619623,);
nor I_36300 (I619631,I619623,I619374);
DFFARX1 I_36301 (I619631,I2507,I619190,I619158,);
DFFARX1 I_36302 (I619623,I2507,I619190,I619182,);
not I_36303 (I619676,I619623);
nor I_36304 (I619693,I619676,I619250);
nor I_36305 (I619710,I619515,I619693);
DFFARX1 I_36306 (I619710,I2507,I619190,I619179,);
not I_36307 (I619768,I2514);
DFFARX1 I_36308 (I753832,I2507,I619768,I619794,);
not I_36309 (I619802,I619794);
DFFARX1 I_36310 (I753844,I2507,I619768,I619828,);
not I_36311 (I619836,I753835);
nand I_36312 (I619853,I619836,I753838);
not I_36313 (I619870,I619853);
nor I_36314 (I619887,I619870,I753841);
nor I_36315 (I619904,I619802,I619887);
DFFARX1 I_36316 (I619904,I2507,I619768,I619754,);
not I_36317 (I619935,I753841);
nand I_36318 (I619952,I619935,I619870);
and I_36319 (I619969,I619935,I753835);
nand I_36320 (I619986,I619969,I753847);
nor I_36321 (I619751,I619986,I619935);
and I_36322 (I619742,I619828,I619986);
not I_36323 (I620031,I619986);
nand I_36324 (I619745,I619828,I620031);
nor I_36325 (I619739,I619794,I619986);
not I_36326 (I620076,I753853);
nor I_36327 (I620093,I620076,I753835);
nand I_36328 (I620110,I620093,I619935);
nor I_36329 (I619748,I619853,I620110);
nor I_36330 (I620141,I620076,I753832);
and I_36331 (I620158,I620141,I753850);
or I_36332 (I620175,I620158,I753856);
DFFARX1 I_36333 (I620175,I2507,I619768,I620201,);
nor I_36334 (I620209,I620201,I619952);
DFFARX1 I_36335 (I620209,I2507,I619768,I619736,);
DFFARX1 I_36336 (I620201,I2507,I619768,I619760,);
not I_36337 (I620254,I620201);
nor I_36338 (I620271,I620254,I619828);
nor I_36339 (I620288,I620093,I620271);
DFFARX1 I_36340 (I620288,I2507,I619768,I619757,);
not I_36341 (I620346,I2514);
DFFARX1 I_36342 (I1150272,I2507,I620346,I620372,);
not I_36343 (I620380,I620372);
DFFARX1 I_36344 (I1150278,I2507,I620346,I620406,);
not I_36345 (I620414,I1150272);
nand I_36346 (I620431,I620414,I1150275);
not I_36347 (I620448,I620431);
nor I_36348 (I620465,I620448,I1150293);
nor I_36349 (I620482,I620380,I620465);
DFFARX1 I_36350 (I620482,I2507,I620346,I620332,);
not I_36351 (I620513,I1150293);
nand I_36352 (I620530,I620513,I620448);
and I_36353 (I620547,I620513,I1150296);
nand I_36354 (I620564,I620547,I1150275);
nor I_36355 (I620329,I620564,I620513);
and I_36356 (I620320,I620406,I620564);
not I_36357 (I620609,I620564);
nand I_36358 (I620323,I620406,I620609);
nor I_36359 (I620317,I620372,I620564);
not I_36360 (I620654,I1150281);
nor I_36361 (I620671,I620654,I1150296);
nand I_36362 (I620688,I620671,I620513);
nor I_36363 (I620326,I620431,I620688);
nor I_36364 (I620719,I620654,I1150287);
and I_36365 (I620736,I620719,I1150284);
or I_36366 (I620753,I620736,I1150290);
DFFARX1 I_36367 (I620753,I2507,I620346,I620779,);
nor I_36368 (I620787,I620779,I620530);
DFFARX1 I_36369 (I620787,I2507,I620346,I620314,);
DFFARX1 I_36370 (I620779,I2507,I620346,I620338,);
not I_36371 (I620832,I620779);
nor I_36372 (I620849,I620832,I620406);
nor I_36373 (I620866,I620671,I620849);
DFFARX1 I_36374 (I620866,I2507,I620346,I620335,);
not I_36375 (I620924,I2514);
DFFARX1 I_36376 (I1362432,I2507,I620924,I620950,);
not I_36377 (I620958,I620950);
DFFARX1 I_36378 (I1362432,I2507,I620924,I620984,);
not I_36379 (I620992,I1362456);
nand I_36380 (I621009,I620992,I1362438);
not I_36381 (I621026,I621009);
nor I_36382 (I621043,I621026,I1362453);
nor I_36383 (I621060,I620958,I621043);
DFFARX1 I_36384 (I621060,I2507,I620924,I620910,);
not I_36385 (I621091,I1362453);
nand I_36386 (I621108,I621091,I621026);
and I_36387 (I621125,I621091,I1362435);
nand I_36388 (I621142,I621125,I1362444);
nor I_36389 (I620907,I621142,I621091);
and I_36390 (I620898,I620984,I621142);
not I_36391 (I621187,I621142);
nand I_36392 (I620901,I620984,I621187);
nor I_36393 (I620895,I620950,I621142);
not I_36394 (I621232,I1362441);
nor I_36395 (I621249,I621232,I1362435);
nand I_36396 (I621266,I621249,I621091);
nor I_36397 (I620904,I621009,I621266);
nor I_36398 (I621297,I621232,I1362450);
and I_36399 (I621314,I621297,I1362459);
or I_36400 (I621331,I621314,I1362447);
DFFARX1 I_36401 (I621331,I2507,I620924,I621357,);
nor I_36402 (I621365,I621357,I621108);
DFFARX1 I_36403 (I621365,I2507,I620924,I620892,);
DFFARX1 I_36404 (I621357,I2507,I620924,I620916,);
not I_36405 (I621410,I621357);
nor I_36406 (I621427,I621410,I620984);
nor I_36407 (I621444,I621249,I621427);
DFFARX1 I_36408 (I621444,I2507,I620924,I620913,);
not I_36409 (I621502,I2514);
DFFARX1 I_36410 (I1231924,I2507,I621502,I621528,);
not I_36411 (I621536,I621528);
DFFARX1 I_36412 (I1231918,I2507,I621502,I621562,);
not I_36413 (I621570,I1231927);
nand I_36414 (I621587,I621570,I1231906);
not I_36415 (I621604,I621587);
nor I_36416 (I621621,I621604,I1231915);
nor I_36417 (I621638,I621536,I621621);
DFFARX1 I_36418 (I621638,I2507,I621502,I621488,);
not I_36419 (I621669,I1231915);
nand I_36420 (I621686,I621669,I621604);
and I_36421 (I621703,I621669,I1231930);
nand I_36422 (I621720,I621703,I1231909);
nor I_36423 (I621485,I621720,I621669);
and I_36424 (I621476,I621562,I621720);
not I_36425 (I621765,I621720);
nand I_36426 (I621479,I621562,I621765);
nor I_36427 (I621473,I621528,I621720);
not I_36428 (I621810,I1231912);
nor I_36429 (I621827,I621810,I1231930);
nand I_36430 (I621844,I621827,I621669);
nor I_36431 (I621482,I621587,I621844);
nor I_36432 (I621875,I621810,I1231921);
and I_36433 (I621892,I621875,I1231909);
or I_36434 (I621909,I621892,I1231906);
DFFARX1 I_36435 (I621909,I2507,I621502,I621935,);
nor I_36436 (I621943,I621935,I621686);
DFFARX1 I_36437 (I621943,I2507,I621502,I621470,);
DFFARX1 I_36438 (I621935,I2507,I621502,I621494,);
not I_36439 (I621988,I621935);
nor I_36440 (I622005,I621988,I621562);
nor I_36441 (I622022,I621827,I622005);
DFFARX1 I_36442 (I622022,I2507,I621502,I621491,);
not I_36443 (I622080,I2514);
DFFARX1 I_36444 (I447963,I2507,I622080,I622106,);
not I_36445 (I622114,I622106);
DFFARX1 I_36446 (I447975,I2507,I622080,I622140,);
not I_36447 (I622148,I447951);
nand I_36448 (I622165,I622148,I447978);
not I_36449 (I622182,I622165);
nor I_36450 (I622199,I622182,I447966);
nor I_36451 (I622216,I622114,I622199);
DFFARX1 I_36452 (I622216,I2507,I622080,I622066,);
not I_36453 (I622247,I447966);
nand I_36454 (I622264,I622247,I622182);
and I_36455 (I622281,I622247,I447951);
nand I_36456 (I622298,I622281,I447954);
nor I_36457 (I622063,I622298,I622247);
and I_36458 (I622054,I622140,I622298);
not I_36459 (I622343,I622298);
nand I_36460 (I622057,I622140,I622343);
nor I_36461 (I622051,I622106,I622298);
not I_36462 (I622388,I447960);
nor I_36463 (I622405,I622388,I447951);
nand I_36464 (I622422,I622405,I622247);
nor I_36465 (I622060,I622165,I622422);
nor I_36466 (I622453,I622388,I447969);
and I_36467 (I622470,I622453,I447957);
or I_36468 (I622487,I622470,I447972);
DFFARX1 I_36469 (I622487,I2507,I622080,I622513,);
nor I_36470 (I622521,I622513,I622264);
DFFARX1 I_36471 (I622521,I2507,I622080,I622048,);
DFFARX1 I_36472 (I622513,I2507,I622080,I622072,);
not I_36473 (I622566,I622513);
nor I_36474 (I622583,I622566,I622140);
nor I_36475 (I622600,I622405,I622583);
DFFARX1 I_36476 (I622600,I2507,I622080,I622069,);
not I_36477 (I622658,I2514);
DFFARX1 I_36478 (I1167612,I2507,I622658,I622684,);
not I_36479 (I622692,I622684);
DFFARX1 I_36480 (I1167618,I2507,I622658,I622718,);
not I_36481 (I622726,I1167612);
nand I_36482 (I622743,I622726,I1167615);
not I_36483 (I622760,I622743);
nor I_36484 (I622777,I622760,I1167633);
nor I_36485 (I622794,I622692,I622777);
DFFARX1 I_36486 (I622794,I2507,I622658,I622644,);
not I_36487 (I622825,I1167633);
nand I_36488 (I622842,I622825,I622760);
and I_36489 (I622859,I622825,I1167636);
nand I_36490 (I622876,I622859,I1167615);
nor I_36491 (I622641,I622876,I622825);
and I_36492 (I622632,I622718,I622876);
not I_36493 (I622921,I622876);
nand I_36494 (I622635,I622718,I622921);
nor I_36495 (I622629,I622684,I622876);
not I_36496 (I622966,I1167621);
nor I_36497 (I622983,I622966,I1167636);
nand I_36498 (I623000,I622983,I622825);
nor I_36499 (I622638,I622743,I623000);
nor I_36500 (I623031,I622966,I1167627);
and I_36501 (I623048,I623031,I1167624);
or I_36502 (I623065,I623048,I1167630);
DFFARX1 I_36503 (I623065,I2507,I622658,I623091,);
nor I_36504 (I623099,I623091,I622842);
DFFARX1 I_36505 (I623099,I2507,I622658,I622626,);
DFFARX1 I_36506 (I623091,I2507,I622658,I622650,);
not I_36507 (I623144,I623091);
nor I_36508 (I623161,I623144,I622718);
nor I_36509 (I623178,I622983,I623161);
DFFARX1 I_36510 (I623178,I2507,I622658,I622647,);
not I_36511 (I623236,I2514);
DFFARX1 I_36512 (I1370762,I2507,I623236,I623262,);
not I_36513 (I623270,I623262);
DFFARX1 I_36514 (I1370762,I2507,I623236,I623296,);
not I_36515 (I623304,I1370786);
nand I_36516 (I623321,I623304,I1370768);
not I_36517 (I623338,I623321);
nor I_36518 (I623355,I623338,I1370783);
nor I_36519 (I623372,I623270,I623355);
DFFARX1 I_36520 (I623372,I2507,I623236,I623222,);
not I_36521 (I623403,I1370783);
nand I_36522 (I623420,I623403,I623338);
and I_36523 (I623437,I623403,I1370765);
nand I_36524 (I623454,I623437,I1370774);
nor I_36525 (I623219,I623454,I623403);
and I_36526 (I623210,I623296,I623454);
not I_36527 (I623499,I623454);
nand I_36528 (I623213,I623296,I623499);
nor I_36529 (I623207,I623262,I623454);
not I_36530 (I623544,I1370771);
nor I_36531 (I623561,I623544,I1370765);
nand I_36532 (I623578,I623561,I623403);
nor I_36533 (I623216,I623321,I623578);
nor I_36534 (I623609,I623544,I1370780);
and I_36535 (I623626,I623609,I1370789);
or I_36536 (I623643,I623626,I1370777);
DFFARX1 I_36537 (I623643,I2507,I623236,I623669,);
nor I_36538 (I623677,I623669,I623420);
DFFARX1 I_36539 (I623677,I2507,I623236,I623204,);
DFFARX1 I_36540 (I623669,I2507,I623236,I623228,);
not I_36541 (I623722,I623669);
nor I_36542 (I623739,I623722,I623296);
nor I_36543 (I623756,I623561,I623739);
DFFARX1 I_36544 (I623756,I2507,I623236,I623225,);
not I_36545 (I623814,I2514);
DFFARX1 I_36546 (I682738,I2507,I623814,I623840,);
not I_36547 (I623848,I623840);
DFFARX1 I_36548 (I682750,I2507,I623814,I623874,);
not I_36549 (I623882,I682741);
nand I_36550 (I623899,I623882,I682744);
not I_36551 (I623916,I623899);
nor I_36552 (I623933,I623916,I682747);
nor I_36553 (I623950,I623848,I623933);
DFFARX1 I_36554 (I623950,I2507,I623814,I623800,);
not I_36555 (I623981,I682747);
nand I_36556 (I623998,I623981,I623916);
and I_36557 (I624015,I623981,I682741);
nand I_36558 (I624032,I624015,I682753);
nor I_36559 (I623797,I624032,I623981);
and I_36560 (I623788,I623874,I624032);
not I_36561 (I624077,I624032);
nand I_36562 (I623791,I623874,I624077);
nor I_36563 (I623785,I623840,I624032);
not I_36564 (I624122,I682759);
nor I_36565 (I624139,I624122,I682741);
nand I_36566 (I624156,I624139,I623981);
nor I_36567 (I623794,I623899,I624156);
nor I_36568 (I624187,I624122,I682738);
and I_36569 (I624204,I624187,I682756);
or I_36570 (I624221,I624204,I682762);
DFFARX1 I_36571 (I624221,I2507,I623814,I624247,);
nor I_36572 (I624255,I624247,I623998);
DFFARX1 I_36573 (I624255,I2507,I623814,I623782,);
DFFARX1 I_36574 (I624247,I2507,I623814,I623806,);
not I_36575 (I624300,I624247);
nor I_36576 (I624317,I624300,I623874);
nor I_36577 (I624334,I624139,I624317);
DFFARX1 I_36578 (I624334,I2507,I623814,I623803,);
not I_36579 (I624392,I2514);
DFFARX1 I_36580 (I838617,I2507,I624392,I624418,);
not I_36581 (I624426,I624418);
DFFARX1 I_36582 (I838617,I2507,I624392,I624452,);
not I_36583 (I624460,I838614);
nand I_36584 (I624477,I624460,I838629);
not I_36585 (I624494,I624477);
nor I_36586 (I624511,I624494,I838623);
nor I_36587 (I624528,I624426,I624511);
DFFARX1 I_36588 (I624528,I2507,I624392,I624378,);
not I_36589 (I624559,I838623);
nand I_36590 (I624576,I624559,I624494);
and I_36591 (I624593,I624559,I838620);
nand I_36592 (I624610,I624593,I838611);
nor I_36593 (I624375,I624610,I624559);
and I_36594 (I624366,I624452,I624610);
not I_36595 (I624655,I624610);
nand I_36596 (I624369,I624452,I624655);
nor I_36597 (I624363,I624418,I624610);
not I_36598 (I624700,I838632);
nor I_36599 (I624717,I624700,I838620);
nand I_36600 (I624734,I624717,I624559);
nor I_36601 (I624372,I624477,I624734);
nor I_36602 (I624765,I624700,I838611);
and I_36603 (I624782,I624765,I838614);
or I_36604 (I624799,I624782,I838626);
DFFARX1 I_36605 (I624799,I2507,I624392,I624825,);
nor I_36606 (I624833,I624825,I624576);
DFFARX1 I_36607 (I624833,I2507,I624392,I624360,);
DFFARX1 I_36608 (I624825,I2507,I624392,I624384,);
not I_36609 (I624878,I624825);
nor I_36610 (I624895,I624878,I624452);
nor I_36611 (I624912,I624717,I624895);
DFFARX1 I_36612 (I624912,I2507,I624392,I624381,);
not I_36613 (I624970,I2514);
DFFARX1 I_36614 (I1365407,I2507,I624970,I624996,);
not I_36615 (I625004,I624996);
DFFARX1 I_36616 (I1365407,I2507,I624970,I625030,);
not I_36617 (I625038,I1365431);
nand I_36618 (I625055,I625038,I1365413);
not I_36619 (I625072,I625055);
nor I_36620 (I625089,I625072,I1365428);
nor I_36621 (I625106,I625004,I625089);
DFFARX1 I_36622 (I625106,I2507,I624970,I624956,);
not I_36623 (I625137,I1365428);
nand I_36624 (I625154,I625137,I625072);
and I_36625 (I625171,I625137,I1365410);
nand I_36626 (I625188,I625171,I1365419);
nor I_36627 (I624953,I625188,I625137);
and I_36628 (I624944,I625030,I625188);
not I_36629 (I625233,I625188);
nand I_36630 (I624947,I625030,I625233);
nor I_36631 (I624941,I624996,I625188);
not I_36632 (I625278,I1365416);
nor I_36633 (I625295,I625278,I1365410);
nand I_36634 (I625312,I625295,I625137);
nor I_36635 (I624950,I625055,I625312);
nor I_36636 (I625343,I625278,I1365425);
and I_36637 (I625360,I625343,I1365434);
or I_36638 (I625377,I625360,I1365422);
DFFARX1 I_36639 (I625377,I2507,I624970,I625403,);
nor I_36640 (I625411,I625403,I625154);
DFFARX1 I_36641 (I625411,I2507,I624970,I624938,);
DFFARX1 I_36642 (I625403,I2507,I624970,I624962,);
not I_36643 (I625456,I625403);
nor I_36644 (I625473,I625456,I625030);
nor I_36645 (I625490,I625295,I625473);
DFFARX1 I_36646 (I625490,I2507,I624970,I624959,);
not I_36647 (I625548,I2514);
DFFARX1 I_36648 (I977371,I2507,I625548,I625574,);
not I_36649 (I625582,I625574);
DFFARX1 I_36650 (I977368,I2507,I625548,I625608,);
not I_36651 (I625616,I977365);
nand I_36652 (I625633,I625616,I977392);
not I_36653 (I625650,I625633);
nor I_36654 (I625667,I625650,I977380);
nor I_36655 (I625684,I625582,I625667);
DFFARX1 I_36656 (I625684,I2507,I625548,I625534,);
not I_36657 (I625715,I977380);
nand I_36658 (I625732,I625715,I625650);
and I_36659 (I625749,I625715,I977386);
nand I_36660 (I625766,I625749,I977377);
nor I_36661 (I625531,I625766,I625715);
and I_36662 (I625522,I625608,I625766);
not I_36663 (I625811,I625766);
nand I_36664 (I625525,I625608,I625811);
nor I_36665 (I625519,I625574,I625766);
not I_36666 (I625856,I977374);
nor I_36667 (I625873,I625856,I977386);
nand I_36668 (I625890,I625873,I625715);
nor I_36669 (I625528,I625633,I625890);
nor I_36670 (I625921,I625856,I977389);
and I_36671 (I625938,I625921,I977383);
or I_36672 (I625955,I625938,I977365);
DFFARX1 I_36673 (I625955,I2507,I625548,I625981,);
nor I_36674 (I625989,I625981,I625732);
DFFARX1 I_36675 (I625989,I2507,I625548,I625516,);
DFFARX1 I_36676 (I625981,I2507,I625548,I625540,);
not I_36677 (I626034,I625981);
nor I_36678 (I626051,I626034,I625608);
nor I_36679 (I626068,I625873,I626051);
DFFARX1 I_36680 (I626068,I2507,I625548,I625537,);
not I_36681 (I626126,I2514);
DFFARX1 I_36682 (I1201714,I2507,I626126,I626152,);
not I_36683 (I626160,I626152);
DFFARX1 I_36684 (I1201720,I2507,I626126,I626186,);
not I_36685 (I626194,I1201714);
nand I_36686 (I626211,I626194,I1201717);
not I_36687 (I626228,I626211);
nor I_36688 (I626245,I626228,I1201735);
nor I_36689 (I626262,I626160,I626245);
DFFARX1 I_36690 (I626262,I2507,I626126,I626112,);
not I_36691 (I626293,I1201735);
nand I_36692 (I626310,I626293,I626228);
and I_36693 (I626327,I626293,I1201738);
nand I_36694 (I626344,I626327,I1201717);
nor I_36695 (I626109,I626344,I626293);
and I_36696 (I626100,I626186,I626344);
not I_36697 (I626389,I626344);
nand I_36698 (I626103,I626186,I626389);
nor I_36699 (I626097,I626152,I626344);
not I_36700 (I626434,I1201723);
nor I_36701 (I626451,I626434,I1201738);
nand I_36702 (I626468,I626451,I626293);
nor I_36703 (I626106,I626211,I626468);
nor I_36704 (I626499,I626434,I1201729);
and I_36705 (I626516,I626499,I1201726);
or I_36706 (I626533,I626516,I1201732);
DFFARX1 I_36707 (I626533,I2507,I626126,I626559,);
nor I_36708 (I626567,I626559,I626310);
DFFARX1 I_36709 (I626567,I2507,I626126,I626094,);
DFFARX1 I_36710 (I626559,I2507,I626126,I626118,);
not I_36711 (I626612,I626559);
nor I_36712 (I626629,I626612,I626186);
nor I_36713 (I626646,I626451,I626629);
DFFARX1 I_36714 (I626646,I2507,I626126,I626115,);
not I_36715 (I626704,I2514);
DFFARX1 I_36716 (I261790,I2507,I626704,I626730,);
not I_36717 (I626738,I626730);
DFFARX1 I_36718 (I261805,I2507,I626704,I626764,);
not I_36719 (I626772,I261808);
nand I_36720 (I626789,I626772,I261787);
not I_36721 (I626806,I626789);
nor I_36722 (I626823,I626806,I261811);
nor I_36723 (I626840,I626738,I626823);
DFFARX1 I_36724 (I626840,I2507,I626704,I626690,);
not I_36725 (I626871,I261811);
nand I_36726 (I626888,I626871,I626806);
and I_36727 (I626905,I626871,I261793);
nand I_36728 (I626922,I626905,I261784);
nor I_36729 (I626687,I626922,I626871);
and I_36730 (I626678,I626764,I626922);
not I_36731 (I626967,I626922);
nand I_36732 (I626681,I626764,I626967);
nor I_36733 (I626675,I626730,I626922);
not I_36734 (I627012,I261784);
nor I_36735 (I627029,I627012,I261793);
nand I_36736 (I627046,I627029,I626871);
nor I_36737 (I626684,I626789,I627046);
nor I_36738 (I627077,I627012,I261799);
and I_36739 (I627094,I627077,I261802);
or I_36740 (I627111,I627094,I261796);
DFFARX1 I_36741 (I627111,I2507,I626704,I627137,);
nor I_36742 (I627145,I627137,I626888);
DFFARX1 I_36743 (I627145,I2507,I626704,I626672,);
DFFARX1 I_36744 (I627137,I2507,I626704,I626696,);
not I_36745 (I627190,I627137);
nor I_36746 (I627207,I627190,I626764);
nor I_36747 (I627224,I627029,I627207);
DFFARX1 I_36748 (I627224,I2507,I626704,I626693,);
not I_36749 (I627282,I2514);
DFFARX1 I_36750 (I434904,I2507,I627282,I627308,);
not I_36751 (I627316,I627308);
nand I_36752 (I627333,I434895,I434913);
and I_36753 (I627350,I627333,I434916);
DFFARX1 I_36754 (I627350,I2507,I627282,I627376,);
not I_36755 (I627384,I434910);
DFFARX1 I_36756 (I434898,I2507,I627282,I627410,);
not I_36757 (I627418,I627410);
nor I_36758 (I627435,I627418,I627316);
and I_36759 (I627452,I627435,I434910);
nor I_36760 (I627469,I627418,I627384);
nor I_36761 (I627265,I627376,I627469);
DFFARX1 I_36762 (I434907,I2507,I627282,I627509,);
nor I_36763 (I627517,I627509,I627376);
not I_36764 (I627534,I627517);
not I_36765 (I627551,I627509);
nor I_36766 (I627568,I627551,I627452);
DFFARX1 I_36767 (I627568,I2507,I627282,I627268,);
nand I_36768 (I627599,I434922,I434919);
and I_36769 (I627616,I627599,I434901);
DFFARX1 I_36770 (I627616,I2507,I627282,I627642,);
nor I_36771 (I627650,I627642,I627509);
DFFARX1 I_36772 (I627650,I2507,I627282,I627250,);
nand I_36773 (I627681,I627642,I627551);
nand I_36774 (I627259,I627534,I627681);
not I_36775 (I627712,I627642);
nor I_36776 (I627729,I627712,I627452);
DFFARX1 I_36777 (I627729,I2507,I627282,I627271,);
nor I_36778 (I627760,I434895,I434919);
or I_36779 (I627262,I627509,I627760);
nor I_36780 (I627253,I627642,I627760);
or I_36781 (I627256,I627376,I627760);
DFFARX1 I_36782 (I627760,I2507,I627282,I627274,);
not I_36783 (I627860,I2514);
DFFARX1 I_36784 (I617424,I2507,I627860,I627886,);
not I_36785 (I627894,I627886);
nand I_36786 (I627911,I617433,I617442);
and I_36787 (I627928,I627911,I617448);
DFFARX1 I_36788 (I627928,I2507,I627860,I627954,);
not I_36789 (I627962,I617445);
DFFARX1 I_36790 (I617430,I2507,I627860,I627988,);
not I_36791 (I627996,I627988);
nor I_36792 (I628013,I627996,I627894);
and I_36793 (I628030,I628013,I617445);
nor I_36794 (I628047,I627996,I627962);
nor I_36795 (I627843,I627954,I628047);
DFFARX1 I_36796 (I617439,I2507,I627860,I628087,);
nor I_36797 (I628095,I628087,I627954);
not I_36798 (I628112,I628095);
not I_36799 (I628129,I628087);
nor I_36800 (I628146,I628129,I628030);
DFFARX1 I_36801 (I628146,I2507,I627860,I627846,);
nand I_36802 (I628177,I617436,I617427);
and I_36803 (I628194,I628177,I617424);
DFFARX1 I_36804 (I628194,I2507,I627860,I628220,);
nor I_36805 (I628228,I628220,I628087);
DFFARX1 I_36806 (I628228,I2507,I627860,I627828,);
nand I_36807 (I628259,I628220,I628129);
nand I_36808 (I627837,I628112,I628259);
not I_36809 (I628290,I628220);
nor I_36810 (I628307,I628290,I628030);
DFFARX1 I_36811 (I628307,I2507,I627860,I627849,);
nor I_36812 (I628338,I617427,I617427);
or I_36813 (I627840,I628087,I628338);
nor I_36814 (I627831,I628220,I628338);
or I_36815 (I627834,I627954,I628338);
DFFARX1 I_36816 (I628338,I2507,I627860,I627852,);
not I_36817 (I628438,I2514);
DFFARX1 I_36818 (I181170,I2507,I628438,I628464,);
not I_36819 (I628472,I628464);
nand I_36820 (I628489,I181173,I181194);
and I_36821 (I628506,I628489,I181182);
DFFARX1 I_36822 (I628506,I2507,I628438,I628532,);
not I_36823 (I628540,I181179);
DFFARX1 I_36824 (I181170,I2507,I628438,I628566,);
not I_36825 (I628574,I628566);
nor I_36826 (I628591,I628574,I628472);
and I_36827 (I628608,I628591,I181179);
nor I_36828 (I628625,I628574,I628540);
nor I_36829 (I628421,I628532,I628625);
DFFARX1 I_36830 (I181188,I2507,I628438,I628665,);
nor I_36831 (I628673,I628665,I628532);
not I_36832 (I628690,I628673);
not I_36833 (I628707,I628665);
nor I_36834 (I628724,I628707,I628608);
DFFARX1 I_36835 (I628724,I2507,I628438,I628424,);
nand I_36836 (I628755,I181173,I181176);
and I_36837 (I628772,I628755,I181185);
DFFARX1 I_36838 (I628772,I2507,I628438,I628798,);
nor I_36839 (I628806,I628798,I628665);
DFFARX1 I_36840 (I628806,I2507,I628438,I628406,);
nand I_36841 (I628837,I628798,I628707);
nand I_36842 (I628415,I628690,I628837);
not I_36843 (I628868,I628798);
nor I_36844 (I628885,I628868,I628608);
DFFARX1 I_36845 (I628885,I2507,I628438,I628427,);
nor I_36846 (I628916,I181191,I181176);
or I_36847 (I628418,I628665,I628916);
nor I_36848 (I628409,I628798,I628916);
or I_36849 (I628412,I628532,I628916);
DFFARX1 I_36850 (I628916,I2507,I628438,I628430,);
not I_36851 (I629016,I2514);
DFFARX1 I_36852 (I958009,I2507,I629016,I629042,);
not I_36853 (I629050,I629042);
nand I_36854 (I629067,I957985,I958000);
and I_36855 (I629084,I629067,I958012);
DFFARX1 I_36856 (I629084,I2507,I629016,I629110,);
not I_36857 (I629118,I957997);
DFFARX1 I_36858 (I957988,I2507,I629016,I629144,);
not I_36859 (I629152,I629144);
nor I_36860 (I629169,I629152,I629050);
and I_36861 (I629186,I629169,I957997);
nor I_36862 (I629203,I629152,I629118);
nor I_36863 (I628999,I629110,I629203);
DFFARX1 I_36864 (I957985,I2507,I629016,I629243,);
nor I_36865 (I629251,I629243,I629110);
not I_36866 (I629268,I629251);
not I_36867 (I629285,I629243);
nor I_36868 (I629302,I629285,I629186);
DFFARX1 I_36869 (I629302,I2507,I629016,I629002,);
nand I_36870 (I629333,I958003,I957994);
and I_36871 (I629350,I629333,I958006);
DFFARX1 I_36872 (I629350,I2507,I629016,I629376,);
nor I_36873 (I629384,I629376,I629243);
DFFARX1 I_36874 (I629384,I2507,I629016,I628984,);
nand I_36875 (I629415,I629376,I629285);
nand I_36876 (I628993,I629268,I629415);
not I_36877 (I629446,I629376);
nor I_36878 (I629463,I629446,I629186);
DFFARX1 I_36879 (I629463,I2507,I629016,I629005,);
nor I_36880 (I629494,I957991,I957994);
or I_36881 (I628996,I629243,I629494);
nor I_36882 (I628987,I629376,I629494);
or I_36883 (I628990,I629110,I629494);
DFFARX1 I_36884 (I629494,I2507,I629016,I629008,);
not I_36885 (I629594,I2514);
DFFARX1 I_36886 (I1218306,I2507,I629594,I629620,);
not I_36887 (I629628,I629620);
nand I_36888 (I629645,I1218309,I1218318);
and I_36889 (I629662,I629645,I1218321);
DFFARX1 I_36890 (I629662,I2507,I629594,I629688,);
not I_36891 (I629696,I1218330);
DFFARX1 I_36892 (I1218312,I2507,I629594,I629722,);
not I_36893 (I629730,I629722);
nor I_36894 (I629747,I629730,I629628);
and I_36895 (I629764,I629747,I1218330);
nor I_36896 (I629781,I629730,I629696);
nor I_36897 (I629577,I629688,I629781);
DFFARX1 I_36898 (I1218309,I2507,I629594,I629821,);
nor I_36899 (I629829,I629821,I629688);
not I_36900 (I629846,I629829);
not I_36901 (I629863,I629821);
nor I_36902 (I629880,I629863,I629764);
DFFARX1 I_36903 (I629880,I2507,I629594,I629580,);
nand I_36904 (I629911,I1218327,I1218306);
and I_36905 (I629928,I629911,I1218324);
DFFARX1 I_36906 (I629928,I2507,I629594,I629954,);
nor I_36907 (I629962,I629954,I629821);
DFFARX1 I_36908 (I629962,I2507,I629594,I629562,);
nand I_36909 (I629993,I629954,I629863);
nand I_36910 (I629571,I629846,I629993);
not I_36911 (I630024,I629954);
nor I_36912 (I630041,I630024,I629764);
DFFARX1 I_36913 (I630041,I2507,I629594,I629583,);
nor I_36914 (I630072,I1218315,I1218306);
or I_36915 (I629574,I629821,I630072);
nor I_36916 (I629565,I629954,I630072);
or I_36917 (I629568,I629688,I630072);
DFFARX1 I_36918 (I630072,I2507,I629594,I629586,);
not I_36919 (I630172,I2514);
DFFARX1 I_36920 (I1285388,I2507,I630172,I630198,);
not I_36921 (I630206,I630198);
nand I_36922 (I630223,I1285412,I1285394);
and I_36923 (I630240,I630223,I1285400);
DFFARX1 I_36924 (I630240,I2507,I630172,I630266,);
not I_36925 (I630274,I1285406);
DFFARX1 I_36926 (I1285391,I2507,I630172,I630300,);
not I_36927 (I630308,I630300);
nor I_36928 (I630325,I630308,I630206);
and I_36929 (I630342,I630325,I1285406);
nor I_36930 (I630359,I630308,I630274);
nor I_36931 (I630155,I630266,I630359);
DFFARX1 I_36932 (I1285403,I2507,I630172,I630399,);
nor I_36933 (I630407,I630399,I630266);
not I_36934 (I630424,I630407);
not I_36935 (I630441,I630399);
nor I_36936 (I630458,I630441,I630342);
DFFARX1 I_36937 (I630458,I2507,I630172,I630158,);
nand I_36938 (I630489,I1285409,I1285397);
and I_36939 (I630506,I630489,I1285391);
DFFARX1 I_36940 (I630506,I2507,I630172,I630532,);
nor I_36941 (I630540,I630532,I630399);
DFFARX1 I_36942 (I630540,I2507,I630172,I630140,);
nand I_36943 (I630571,I630532,I630441);
nand I_36944 (I630149,I630424,I630571);
not I_36945 (I630602,I630532);
nor I_36946 (I630619,I630602,I630342);
DFFARX1 I_36947 (I630619,I2507,I630172,I630161,);
nor I_36948 (I630650,I1285388,I1285397);
or I_36949 (I630152,I630399,I630650);
nor I_36950 (I630143,I630532,I630650);
or I_36951 (I630146,I630266,I630650);
DFFARX1 I_36952 (I630650,I2507,I630172,I630164,);
not I_36953 (I630750,I2514);
DFFARX1 I_36954 (I1215586,I2507,I630750,I630776,);
not I_36955 (I630784,I630776);
nand I_36956 (I630801,I1215589,I1215598);
and I_36957 (I630818,I630801,I1215601);
DFFARX1 I_36958 (I630818,I2507,I630750,I630844,);
not I_36959 (I630852,I1215610);
DFFARX1 I_36960 (I1215592,I2507,I630750,I630878,);
not I_36961 (I630886,I630878);
nor I_36962 (I630903,I630886,I630784);
and I_36963 (I630920,I630903,I1215610);
nor I_36964 (I630937,I630886,I630852);
nor I_36965 (I630733,I630844,I630937);
DFFARX1 I_36966 (I1215589,I2507,I630750,I630977,);
nor I_36967 (I630985,I630977,I630844);
not I_36968 (I631002,I630985);
not I_36969 (I631019,I630977);
nor I_36970 (I631036,I631019,I630920);
DFFARX1 I_36971 (I631036,I2507,I630750,I630736,);
nand I_36972 (I631067,I1215607,I1215586);
and I_36973 (I631084,I631067,I1215604);
DFFARX1 I_36974 (I631084,I2507,I630750,I631110,);
nor I_36975 (I631118,I631110,I630977);
DFFARX1 I_36976 (I631118,I2507,I630750,I630718,);
nand I_36977 (I631149,I631110,I631019);
nand I_36978 (I630727,I631002,I631149);
not I_36979 (I631180,I631110);
nor I_36980 (I631197,I631180,I630920);
DFFARX1 I_36981 (I631197,I2507,I630750,I630739,);
nor I_36982 (I631228,I1215595,I1215586);
or I_36983 (I630730,I630977,I631228);
nor I_36984 (I630721,I631110,I631228);
or I_36985 (I630724,I630844,I631228);
DFFARX1 I_36986 (I631228,I2507,I630750,I630742,);
not I_36987 (I631328,I2514);
DFFARX1 I_36988 (I1163006,I2507,I631328,I631354,);
not I_36989 (I631362,I631354);
nand I_36990 (I631379,I1162988,I1163000);
and I_36991 (I631396,I631379,I1163003);
DFFARX1 I_36992 (I631396,I2507,I631328,I631422,);
not I_36993 (I631430,I1162997);
DFFARX1 I_36994 (I1162994,I2507,I631328,I631456,);
not I_36995 (I631464,I631456);
nor I_36996 (I631481,I631464,I631362);
and I_36997 (I631498,I631481,I1162997);
nor I_36998 (I631515,I631464,I631430);
nor I_36999 (I631311,I631422,I631515);
DFFARX1 I_37000 (I1163012,I2507,I631328,I631555,);
nor I_37001 (I631563,I631555,I631422);
not I_37002 (I631580,I631563);
not I_37003 (I631597,I631555);
nor I_37004 (I631614,I631597,I631498);
DFFARX1 I_37005 (I631614,I2507,I631328,I631314,);
nand I_37006 (I631645,I1162991,I1162991);
and I_37007 (I631662,I631645,I1162988);
DFFARX1 I_37008 (I631662,I2507,I631328,I631688,);
nor I_37009 (I631696,I631688,I631555);
DFFARX1 I_37010 (I631696,I2507,I631328,I631296,);
nand I_37011 (I631727,I631688,I631597);
nand I_37012 (I631305,I631580,I631727);
not I_37013 (I631758,I631688);
nor I_37014 (I631775,I631758,I631498);
DFFARX1 I_37015 (I631775,I2507,I631328,I631317,);
nor I_37016 (I631806,I1163009,I1162991);
or I_37017 (I631308,I631555,I631806);
nor I_37018 (I631299,I631688,I631806);
or I_37019 (I631302,I631422,I631806);
DFFARX1 I_37020 (I631806,I2507,I631328,I631320,);
not I_37021 (I631906,I2514);
DFFARX1 I_37022 (I194855,I2507,I631906,I631932,);
not I_37023 (I631940,I631932);
nand I_37024 (I631957,I194858,I194879);
and I_37025 (I631974,I631957,I194867);
DFFARX1 I_37026 (I631974,I2507,I631906,I632000,);
not I_37027 (I632008,I194864);
DFFARX1 I_37028 (I194855,I2507,I631906,I632034,);
not I_37029 (I632042,I632034);
nor I_37030 (I632059,I632042,I631940);
and I_37031 (I632076,I632059,I194864);
nor I_37032 (I632093,I632042,I632008);
nor I_37033 (I631889,I632000,I632093);
DFFARX1 I_37034 (I194873,I2507,I631906,I632133,);
nor I_37035 (I632141,I632133,I632000);
not I_37036 (I632158,I632141);
not I_37037 (I632175,I632133);
nor I_37038 (I632192,I632175,I632076);
DFFARX1 I_37039 (I632192,I2507,I631906,I631892,);
nand I_37040 (I632223,I194858,I194861);
and I_37041 (I632240,I632223,I194870);
DFFARX1 I_37042 (I632240,I2507,I631906,I632266,);
nor I_37043 (I632274,I632266,I632133);
DFFARX1 I_37044 (I632274,I2507,I631906,I631874,);
nand I_37045 (I632305,I632266,I632175);
nand I_37046 (I631883,I632158,I632305);
not I_37047 (I632336,I632266);
nor I_37048 (I632353,I632336,I632076);
DFFARX1 I_37049 (I632353,I2507,I631906,I631895,);
nor I_37050 (I632384,I194876,I194861);
or I_37051 (I631886,I632133,I632384);
nor I_37052 (I631877,I632266,I632384);
or I_37053 (I631880,I632000,I632384);
DFFARX1 I_37054 (I632384,I2507,I631906,I631898,);
not I_37055 (I632484,I2514);
DFFARX1 I_37056 (I389752,I2507,I632484,I632510,);
not I_37057 (I632518,I632510);
nand I_37058 (I632535,I389743,I389761);
and I_37059 (I632552,I632535,I389764);
DFFARX1 I_37060 (I632552,I2507,I632484,I632578,);
not I_37061 (I632586,I389758);
DFFARX1 I_37062 (I389746,I2507,I632484,I632612,);
not I_37063 (I632620,I632612);
nor I_37064 (I632637,I632620,I632518);
and I_37065 (I632654,I632637,I389758);
nor I_37066 (I632671,I632620,I632586);
nor I_37067 (I632467,I632578,I632671);
DFFARX1 I_37068 (I389755,I2507,I632484,I632711,);
nor I_37069 (I632719,I632711,I632578);
not I_37070 (I632736,I632719);
not I_37071 (I632753,I632711);
nor I_37072 (I632770,I632753,I632654);
DFFARX1 I_37073 (I632770,I2507,I632484,I632470,);
nand I_37074 (I632801,I389770,I389767);
and I_37075 (I632818,I632801,I389749);
DFFARX1 I_37076 (I632818,I2507,I632484,I632844,);
nor I_37077 (I632852,I632844,I632711);
DFFARX1 I_37078 (I632852,I2507,I632484,I632452,);
nand I_37079 (I632883,I632844,I632753);
nand I_37080 (I632461,I632736,I632883);
not I_37081 (I632914,I632844);
nor I_37082 (I632931,I632914,I632654);
DFFARX1 I_37083 (I632931,I2507,I632484,I632473,);
nor I_37084 (I632962,I389743,I389767);
or I_37085 (I632464,I632711,I632962);
nor I_37086 (I632455,I632844,I632962);
or I_37087 (I632458,I632578,I632962);
DFFARX1 I_37088 (I632962,I2507,I632484,I632476,);
not I_37089 (I633062,I2514);
DFFARX1 I_37090 (I272348,I2507,I633062,I633088,);
not I_37091 (I633096,I633088);
nand I_37092 (I633113,I272351,I272327);
and I_37093 (I633130,I633113,I272324);
DFFARX1 I_37094 (I633130,I2507,I633062,I633156,);
not I_37095 (I633164,I272330);
DFFARX1 I_37096 (I272324,I2507,I633062,I633190,);
not I_37097 (I633198,I633190);
nor I_37098 (I633215,I633198,I633096);
and I_37099 (I633232,I633215,I272330);
nor I_37100 (I633249,I633198,I633164);
nor I_37101 (I633045,I633156,I633249);
DFFARX1 I_37102 (I272333,I2507,I633062,I633289,);
nor I_37103 (I633297,I633289,I633156);
not I_37104 (I633314,I633297);
not I_37105 (I633331,I633289);
nor I_37106 (I633348,I633331,I633232);
DFFARX1 I_37107 (I633348,I2507,I633062,I633048,);
nand I_37108 (I633379,I272336,I272345);
and I_37109 (I633396,I633379,I272342);
DFFARX1 I_37110 (I633396,I2507,I633062,I633422,);
nor I_37111 (I633430,I633422,I633289);
DFFARX1 I_37112 (I633430,I2507,I633062,I633030,);
nand I_37113 (I633461,I633422,I633331);
nand I_37114 (I633039,I633314,I633461);
not I_37115 (I633492,I633422);
nor I_37116 (I633509,I633492,I633232);
DFFARX1 I_37117 (I633509,I2507,I633062,I633051,);
nor I_37118 (I633540,I272339,I272345);
or I_37119 (I633042,I633289,I633540);
nor I_37120 (I633033,I633422,I633540);
or I_37121 (I633036,I633156,I633540);
DFFARX1 I_37122 (I633540,I2507,I633062,I633054,);
not I_37123 (I633640,I2514);
DFFARX1 I_37124 (I947027,I2507,I633640,I633666,);
not I_37125 (I633674,I633666);
nand I_37126 (I633691,I947003,I947018);
and I_37127 (I633708,I633691,I947030);
DFFARX1 I_37128 (I633708,I2507,I633640,I633734,);
not I_37129 (I633742,I947015);
DFFARX1 I_37130 (I947006,I2507,I633640,I633768,);
not I_37131 (I633776,I633768);
nor I_37132 (I633793,I633776,I633674);
and I_37133 (I633810,I633793,I947015);
nor I_37134 (I633827,I633776,I633742);
nor I_37135 (I633623,I633734,I633827);
DFFARX1 I_37136 (I947003,I2507,I633640,I633867,);
nor I_37137 (I633875,I633867,I633734);
not I_37138 (I633892,I633875);
not I_37139 (I633909,I633867);
nor I_37140 (I633926,I633909,I633810);
DFFARX1 I_37141 (I633926,I2507,I633640,I633626,);
nand I_37142 (I633957,I947021,I947012);
and I_37143 (I633974,I633957,I947024);
DFFARX1 I_37144 (I633974,I2507,I633640,I634000,);
nor I_37145 (I634008,I634000,I633867);
DFFARX1 I_37146 (I634008,I2507,I633640,I633608,);
nand I_37147 (I634039,I634000,I633909);
nand I_37148 (I633617,I633892,I634039);
not I_37149 (I634070,I634000);
nor I_37150 (I634087,I634070,I633810);
DFFARX1 I_37151 (I634087,I2507,I633640,I633629,);
nor I_37152 (I634118,I947009,I947012);
or I_37153 (I633620,I633867,I634118);
nor I_37154 (I633611,I634000,I634118);
or I_37155 (I633614,I633734,I634118);
DFFARX1 I_37156 (I634118,I2507,I633640,I633632,);
not I_37157 (I634218,I2514);
DFFARX1 I_37158 (I1059544,I2507,I634218,I634244,);
not I_37159 (I634252,I634244);
nand I_37160 (I634269,I1059526,I1059538);
and I_37161 (I634286,I634269,I1059541);
DFFARX1 I_37162 (I634286,I2507,I634218,I634312,);
not I_37163 (I634320,I1059535);
DFFARX1 I_37164 (I1059532,I2507,I634218,I634346,);
not I_37165 (I634354,I634346);
nor I_37166 (I634371,I634354,I634252);
and I_37167 (I634388,I634371,I1059535);
nor I_37168 (I634405,I634354,I634320);
nor I_37169 (I634201,I634312,I634405);
DFFARX1 I_37170 (I1059550,I2507,I634218,I634445,);
nor I_37171 (I634453,I634445,I634312);
not I_37172 (I634470,I634453);
not I_37173 (I634487,I634445);
nor I_37174 (I634504,I634487,I634388);
DFFARX1 I_37175 (I634504,I2507,I634218,I634204,);
nand I_37176 (I634535,I1059529,I1059529);
and I_37177 (I634552,I634535,I1059526);
DFFARX1 I_37178 (I634552,I2507,I634218,I634578,);
nor I_37179 (I634586,I634578,I634445);
DFFARX1 I_37180 (I634586,I2507,I634218,I634186,);
nand I_37181 (I634617,I634578,I634487);
nand I_37182 (I634195,I634470,I634617);
not I_37183 (I634648,I634578);
nor I_37184 (I634665,I634648,I634388);
DFFARX1 I_37185 (I634665,I2507,I634218,I634207,);
nor I_37186 (I634696,I1059547,I1059529);
or I_37187 (I634198,I634445,I634696);
nor I_37188 (I634189,I634578,I634696);
or I_37189 (I634192,I634312,I634696);
DFFARX1 I_37190 (I634696,I2507,I634218,I634210,);
not I_37191 (I634796,I2514);
DFFARX1 I_37192 (I291320,I2507,I634796,I634822,);
not I_37193 (I634830,I634822);
nand I_37194 (I634847,I291323,I291299);
and I_37195 (I634864,I634847,I291296);
DFFARX1 I_37196 (I634864,I2507,I634796,I634890,);
not I_37197 (I634898,I291302);
DFFARX1 I_37198 (I291296,I2507,I634796,I634924,);
not I_37199 (I634932,I634924);
nor I_37200 (I634949,I634932,I634830);
and I_37201 (I634966,I634949,I291302);
nor I_37202 (I634983,I634932,I634898);
nor I_37203 (I634779,I634890,I634983);
DFFARX1 I_37204 (I291305,I2507,I634796,I635023,);
nor I_37205 (I635031,I635023,I634890);
not I_37206 (I635048,I635031);
not I_37207 (I635065,I635023);
nor I_37208 (I635082,I635065,I634966);
DFFARX1 I_37209 (I635082,I2507,I634796,I634782,);
nand I_37210 (I635113,I291308,I291317);
and I_37211 (I635130,I635113,I291314);
DFFARX1 I_37212 (I635130,I2507,I634796,I635156,);
nor I_37213 (I635164,I635156,I635023);
DFFARX1 I_37214 (I635164,I2507,I634796,I634764,);
nand I_37215 (I635195,I635156,I635065);
nand I_37216 (I634773,I635048,I635195);
not I_37217 (I635226,I635156);
nor I_37218 (I635243,I635226,I634966);
DFFARX1 I_37219 (I635243,I2507,I634796,I634785,);
nor I_37220 (I635274,I291311,I291317);
or I_37221 (I634776,I635023,I635274);
nor I_37222 (I634767,I635156,I635274);
or I_37223 (I634770,I634890,I635274);
DFFARX1 I_37224 (I635274,I2507,I634796,I634788,);
not I_37225 (I635374,I2514);
DFFARX1 I_37226 (I812803,I2507,I635374,I635400,);
not I_37227 (I635408,I635400);
nand I_37228 (I635425,I812791,I812809);
and I_37229 (I635442,I635425,I812806);
DFFARX1 I_37230 (I635442,I2507,I635374,I635468,);
not I_37231 (I635476,I812797);
DFFARX1 I_37232 (I812794,I2507,I635374,I635502,);
not I_37233 (I635510,I635502);
nor I_37234 (I635527,I635510,I635408);
and I_37235 (I635544,I635527,I812797);
nor I_37236 (I635561,I635510,I635476);
nor I_37237 (I635357,I635468,I635561);
DFFARX1 I_37238 (I812788,I2507,I635374,I635601,);
nor I_37239 (I635609,I635601,I635468);
not I_37240 (I635626,I635609);
not I_37241 (I635643,I635601);
nor I_37242 (I635660,I635643,I635544);
DFFARX1 I_37243 (I635660,I2507,I635374,I635360,);
nand I_37244 (I635691,I812788,I812791);
and I_37245 (I635708,I635691,I812794);
DFFARX1 I_37246 (I635708,I2507,I635374,I635734,);
nor I_37247 (I635742,I635734,I635601);
DFFARX1 I_37248 (I635742,I2507,I635374,I635342,);
nand I_37249 (I635773,I635734,I635643);
nand I_37250 (I635351,I635626,I635773);
not I_37251 (I635804,I635734);
nor I_37252 (I635821,I635804,I635544);
DFFARX1 I_37253 (I635821,I2507,I635374,I635363,);
nor I_37254 (I635852,I812800,I812791);
or I_37255 (I635354,I635601,I635852);
nor I_37256 (I635345,I635734,I635852);
or I_37257 (I635348,I635468,I635852);
DFFARX1 I_37258 (I635852,I2507,I635374,I635366,);
not I_37259 (I635952,I2514);
DFFARX1 I_37260 (I799628,I2507,I635952,I635978,);
not I_37261 (I635986,I635978);
nand I_37262 (I636003,I799616,I799634);
and I_37263 (I636020,I636003,I799631);
DFFARX1 I_37264 (I636020,I2507,I635952,I636046,);
not I_37265 (I636054,I799622);
DFFARX1 I_37266 (I799619,I2507,I635952,I636080,);
not I_37267 (I636088,I636080);
nor I_37268 (I636105,I636088,I635986);
and I_37269 (I636122,I636105,I799622);
nor I_37270 (I636139,I636088,I636054);
nor I_37271 (I635935,I636046,I636139);
DFFARX1 I_37272 (I799613,I2507,I635952,I636179,);
nor I_37273 (I636187,I636179,I636046);
not I_37274 (I636204,I636187);
not I_37275 (I636221,I636179);
nor I_37276 (I636238,I636221,I636122);
DFFARX1 I_37277 (I636238,I2507,I635952,I635938,);
nand I_37278 (I636269,I799613,I799616);
and I_37279 (I636286,I636269,I799619);
DFFARX1 I_37280 (I636286,I2507,I635952,I636312,);
nor I_37281 (I636320,I636312,I636179);
DFFARX1 I_37282 (I636320,I2507,I635952,I635920,);
nand I_37283 (I636351,I636312,I636221);
nand I_37284 (I635929,I636204,I636351);
not I_37285 (I636382,I636312);
nor I_37286 (I636399,I636382,I636122);
DFFARX1 I_37287 (I636399,I2507,I635952,I635941,);
nor I_37288 (I636430,I799625,I799616);
or I_37289 (I635932,I636179,I636430);
nor I_37290 (I635923,I636312,I636430);
or I_37291 (I635926,I636046,I636430);
DFFARX1 I_37292 (I636430,I2507,I635952,I635944,);
not I_37293 (I636530,I2514);
DFFARX1 I_37294 (I1107518,I2507,I636530,I636556,);
not I_37295 (I636564,I636556);
nand I_37296 (I636581,I1107500,I1107512);
and I_37297 (I636598,I636581,I1107515);
DFFARX1 I_37298 (I636598,I2507,I636530,I636624,);
not I_37299 (I636632,I1107509);
DFFARX1 I_37300 (I1107506,I2507,I636530,I636658,);
not I_37301 (I636666,I636658);
nor I_37302 (I636683,I636666,I636564);
and I_37303 (I636700,I636683,I1107509);
nor I_37304 (I636717,I636666,I636632);
nor I_37305 (I636513,I636624,I636717);
DFFARX1 I_37306 (I1107524,I2507,I636530,I636757,);
nor I_37307 (I636765,I636757,I636624);
not I_37308 (I636782,I636765);
not I_37309 (I636799,I636757);
nor I_37310 (I636816,I636799,I636700);
DFFARX1 I_37311 (I636816,I2507,I636530,I636516,);
nand I_37312 (I636847,I1107503,I1107503);
and I_37313 (I636864,I636847,I1107500);
DFFARX1 I_37314 (I636864,I2507,I636530,I636890,);
nor I_37315 (I636898,I636890,I636757);
DFFARX1 I_37316 (I636898,I2507,I636530,I636498,);
nand I_37317 (I636929,I636890,I636799);
nand I_37318 (I636507,I636782,I636929);
not I_37319 (I636960,I636890);
nor I_37320 (I636977,I636960,I636700);
DFFARX1 I_37321 (I636977,I2507,I636530,I636519,);
nor I_37322 (I637008,I1107521,I1107503);
or I_37323 (I636510,I636757,I637008);
nor I_37324 (I636501,I636890,I637008);
or I_37325 (I636504,I636624,I637008);
DFFARX1 I_37326 (I637008,I2507,I636530,I636522,);
not I_37327 (I637108,I2514);
DFFARX1 I_37328 (I1284810,I2507,I637108,I637134,);
not I_37329 (I637142,I637134);
nand I_37330 (I637159,I1284834,I1284816);
and I_37331 (I637176,I637159,I1284822);
DFFARX1 I_37332 (I637176,I2507,I637108,I637202,);
not I_37333 (I637210,I1284828);
DFFARX1 I_37334 (I1284813,I2507,I637108,I637236,);
not I_37335 (I637244,I637236);
nor I_37336 (I637261,I637244,I637142);
and I_37337 (I637278,I637261,I1284828);
nor I_37338 (I637295,I637244,I637210);
nor I_37339 (I637091,I637202,I637295);
DFFARX1 I_37340 (I1284825,I2507,I637108,I637335,);
nor I_37341 (I637343,I637335,I637202);
not I_37342 (I637360,I637343);
not I_37343 (I637377,I637335);
nor I_37344 (I637394,I637377,I637278);
DFFARX1 I_37345 (I637394,I2507,I637108,I637094,);
nand I_37346 (I637425,I1284831,I1284819);
and I_37347 (I637442,I637425,I1284813);
DFFARX1 I_37348 (I637442,I2507,I637108,I637468,);
nor I_37349 (I637476,I637468,I637335);
DFFARX1 I_37350 (I637476,I2507,I637108,I637076,);
nand I_37351 (I637507,I637468,I637377);
nand I_37352 (I637085,I637360,I637507);
not I_37353 (I637538,I637468);
nor I_37354 (I637555,I637538,I637278);
DFFARX1 I_37355 (I637555,I2507,I637108,I637097,);
nor I_37356 (I637586,I1284810,I1284819);
or I_37357 (I637088,I637335,I637586);
nor I_37358 (I637079,I637468,I637586);
or I_37359 (I637082,I637202,I637586);
DFFARX1 I_37360 (I637586,I2507,I637108,I637100,);
not I_37361 (I637686,I2514);
DFFARX1 I_37362 (I975451,I2507,I637686,I637712,);
not I_37363 (I637720,I637712);
nand I_37364 (I637737,I975427,I975442);
and I_37365 (I637754,I637737,I975454);
DFFARX1 I_37366 (I637754,I2507,I637686,I637780,);
not I_37367 (I637788,I975439);
DFFARX1 I_37368 (I975430,I2507,I637686,I637814,);
not I_37369 (I637822,I637814);
nor I_37370 (I637839,I637822,I637720);
and I_37371 (I637856,I637839,I975439);
nor I_37372 (I637873,I637822,I637788);
nor I_37373 (I637669,I637780,I637873);
DFFARX1 I_37374 (I975427,I2507,I637686,I637913,);
nor I_37375 (I637921,I637913,I637780);
not I_37376 (I637938,I637921);
not I_37377 (I637955,I637913);
nor I_37378 (I637972,I637955,I637856);
DFFARX1 I_37379 (I637972,I2507,I637686,I637672,);
nand I_37380 (I638003,I975445,I975436);
and I_37381 (I638020,I638003,I975448);
DFFARX1 I_37382 (I638020,I2507,I637686,I638046,);
nor I_37383 (I638054,I638046,I637913);
DFFARX1 I_37384 (I638054,I2507,I637686,I637654,);
nand I_37385 (I638085,I638046,I637955);
nand I_37386 (I637663,I637938,I638085);
not I_37387 (I638116,I638046);
nor I_37388 (I638133,I638116,I637856);
DFFARX1 I_37389 (I638133,I2507,I637686,I637675,);
nor I_37390 (I638164,I975433,I975436);
or I_37391 (I637666,I637913,I638164);
nor I_37392 (I637657,I638046,I638164);
or I_37393 (I637660,I637780,I638164);
DFFARX1 I_37394 (I638164,I2507,I637686,I637678,);
not I_37395 (I638264,I2514);
DFFARX1 I_37396 (I1153758,I2507,I638264,I638290,);
not I_37397 (I638298,I638290);
nand I_37398 (I638315,I1153740,I1153752);
and I_37399 (I638332,I638315,I1153755);
DFFARX1 I_37400 (I638332,I2507,I638264,I638358,);
not I_37401 (I638366,I1153749);
DFFARX1 I_37402 (I1153746,I2507,I638264,I638392,);
not I_37403 (I638400,I638392);
nor I_37404 (I638417,I638400,I638298);
and I_37405 (I638434,I638417,I1153749);
nor I_37406 (I638451,I638400,I638366);
nor I_37407 (I638247,I638358,I638451);
DFFARX1 I_37408 (I1153764,I2507,I638264,I638491,);
nor I_37409 (I638499,I638491,I638358);
not I_37410 (I638516,I638499);
not I_37411 (I638533,I638491);
nor I_37412 (I638550,I638533,I638434);
DFFARX1 I_37413 (I638550,I2507,I638264,I638250,);
nand I_37414 (I638581,I1153743,I1153743);
and I_37415 (I638598,I638581,I1153740);
DFFARX1 I_37416 (I638598,I2507,I638264,I638624,);
nor I_37417 (I638632,I638624,I638491);
DFFARX1 I_37418 (I638632,I2507,I638264,I638232,);
nand I_37419 (I638663,I638624,I638533);
nand I_37420 (I638241,I638516,I638663);
not I_37421 (I638694,I638624);
nor I_37422 (I638711,I638694,I638434);
DFFARX1 I_37423 (I638711,I2507,I638264,I638253,);
nor I_37424 (I638742,I1153761,I1153743);
or I_37425 (I638244,I638491,I638742);
nor I_37426 (I638235,I638624,I638742);
or I_37427 (I638238,I638358,I638742);
DFFARX1 I_37428 (I638742,I2507,I638264,I638256,);
not I_37429 (I638842,I2514);
DFFARX1 I_37430 (I376152,I2507,I638842,I638868,);
not I_37431 (I638876,I638868);
nand I_37432 (I638893,I376143,I376161);
and I_37433 (I638910,I638893,I376164);
DFFARX1 I_37434 (I638910,I2507,I638842,I638936,);
not I_37435 (I638944,I376158);
DFFARX1 I_37436 (I376146,I2507,I638842,I638970,);
not I_37437 (I638978,I638970);
nor I_37438 (I638995,I638978,I638876);
and I_37439 (I639012,I638995,I376158);
nor I_37440 (I639029,I638978,I638944);
nor I_37441 (I638825,I638936,I639029);
DFFARX1 I_37442 (I376155,I2507,I638842,I639069,);
nor I_37443 (I639077,I639069,I638936);
not I_37444 (I639094,I639077);
not I_37445 (I639111,I639069);
nor I_37446 (I639128,I639111,I639012);
DFFARX1 I_37447 (I639128,I2507,I638842,I638828,);
nand I_37448 (I639159,I376170,I376167);
and I_37449 (I639176,I639159,I376149);
DFFARX1 I_37450 (I639176,I2507,I638842,I639202,);
nor I_37451 (I639210,I639202,I639069);
DFFARX1 I_37452 (I639210,I2507,I638842,I638810,);
nand I_37453 (I639241,I639202,I639111);
nand I_37454 (I638819,I639094,I639241);
not I_37455 (I639272,I639202);
nor I_37456 (I639289,I639272,I639012);
DFFARX1 I_37457 (I639289,I2507,I638842,I638831,);
nor I_37458 (I639320,I376143,I376167);
or I_37459 (I638822,I639069,I639320);
nor I_37460 (I638813,I639202,I639320);
or I_37461 (I638816,I638936,I639320);
DFFARX1 I_37462 (I639320,I2507,I638842,I638834,);
not I_37463 (I639420,I2514);
DFFARX1 I_37464 (I794885,I2507,I639420,I639446,);
not I_37465 (I639454,I639446);
nand I_37466 (I639471,I794873,I794891);
and I_37467 (I639488,I639471,I794888);
DFFARX1 I_37468 (I639488,I2507,I639420,I639514,);
not I_37469 (I639522,I794879);
DFFARX1 I_37470 (I794876,I2507,I639420,I639548,);
not I_37471 (I639556,I639548);
nor I_37472 (I639573,I639556,I639454);
and I_37473 (I639590,I639573,I794879);
nor I_37474 (I639607,I639556,I639522);
nor I_37475 (I639403,I639514,I639607);
DFFARX1 I_37476 (I794870,I2507,I639420,I639647,);
nor I_37477 (I639655,I639647,I639514);
not I_37478 (I639672,I639655);
not I_37479 (I639689,I639647);
nor I_37480 (I639706,I639689,I639590);
DFFARX1 I_37481 (I639706,I2507,I639420,I639406,);
nand I_37482 (I639737,I794870,I794873);
and I_37483 (I639754,I639737,I794876);
DFFARX1 I_37484 (I639754,I2507,I639420,I639780,);
nor I_37485 (I639788,I639780,I639647);
DFFARX1 I_37486 (I639788,I2507,I639420,I639388,);
nand I_37487 (I639819,I639780,I639689);
nand I_37488 (I639397,I639672,I639819);
not I_37489 (I639850,I639780);
nor I_37490 (I639867,I639850,I639590);
DFFARX1 I_37491 (I639867,I2507,I639420,I639409,);
nor I_37492 (I639898,I794882,I794873);
or I_37493 (I639400,I639647,I639898);
nor I_37494 (I639391,I639780,I639898);
or I_37495 (I639394,I639514,I639898);
DFFARX1 I_37496 (I639898,I2507,I639420,I639412,);
not I_37497 (I639998,I2514);
DFFARX1 I_37498 (I14293,I2507,I639998,I640024,);
not I_37499 (I640032,I640024);
nand I_37500 (I640049,I14290,I14281);
and I_37501 (I640066,I640049,I14281);
DFFARX1 I_37502 (I640066,I2507,I639998,I640092,);
not I_37503 (I640100,I14284);
DFFARX1 I_37504 (I14299,I2507,I639998,I640126,);
not I_37505 (I640134,I640126);
nor I_37506 (I640151,I640134,I640032);
and I_37507 (I640168,I640151,I14284);
nor I_37508 (I640185,I640134,I640100);
nor I_37509 (I639981,I640092,I640185);
DFFARX1 I_37510 (I14284,I2507,I639998,I640225,);
nor I_37511 (I640233,I640225,I640092);
not I_37512 (I640250,I640233);
not I_37513 (I640267,I640225);
nor I_37514 (I640284,I640267,I640168);
DFFARX1 I_37515 (I640284,I2507,I639998,I639984,);
nand I_37516 (I640315,I14302,I14287);
and I_37517 (I640332,I640315,I14305);
DFFARX1 I_37518 (I640332,I2507,I639998,I640358,);
nor I_37519 (I640366,I640358,I640225);
DFFARX1 I_37520 (I640366,I2507,I639998,I639966,);
nand I_37521 (I640397,I640358,I640267);
nand I_37522 (I639975,I640250,I640397);
not I_37523 (I640428,I640358);
nor I_37524 (I640445,I640428,I640168);
DFFARX1 I_37525 (I640445,I2507,I639998,I639987,);
nor I_37526 (I640476,I14296,I14287);
or I_37527 (I639978,I640225,I640476);
nor I_37528 (I639969,I640358,I640476);
or I_37529 (I639972,I640092,I640476);
DFFARX1 I_37530 (I640476,I2507,I639998,I639990,);
not I_37531 (I640576,I2514);
DFFARX1 I_37532 (I1326164,I2507,I640576,I640602,);
not I_37533 (I640610,I640602);
nand I_37534 (I640627,I1326149,I1326137);
and I_37535 (I640644,I640627,I1326152);
DFFARX1 I_37536 (I640644,I2507,I640576,I640670,);
not I_37537 (I640678,I1326137);
DFFARX1 I_37538 (I1326155,I2507,I640576,I640704,);
not I_37539 (I640712,I640704);
nor I_37540 (I640729,I640712,I640610);
and I_37541 (I640746,I640729,I1326137);
nor I_37542 (I640763,I640712,I640678);
nor I_37543 (I640559,I640670,I640763);
DFFARX1 I_37544 (I1326143,I2507,I640576,I640803,);
nor I_37545 (I640811,I640803,I640670);
not I_37546 (I640828,I640811);
not I_37547 (I640845,I640803);
nor I_37548 (I640862,I640845,I640746);
DFFARX1 I_37549 (I640862,I2507,I640576,I640562,);
nand I_37550 (I640893,I1326140,I1326146);
and I_37551 (I640910,I640893,I1326161);
DFFARX1 I_37552 (I640910,I2507,I640576,I640936,);
nor I_37553 (I640944,I640936,I640803);
DFFARX1 I_37554 (I640944,I2507,I640576,I640544,);
nand I_37555 (I640975,I640936,I640845);
nand I_37556 (I640553,I640828,I640975);
not I_37557 (I641006,I640936);
nor I_37558 (I641023,I641006,I640746);
DFFARX1 I_37559 (I641023,I2507,I640576,I640565,);
nor I_37560 (I641054,I1326158,I1326146);
or I_37561 (I640556,I640803,I641054);
nor I_37562 (I640547,I640936,I641054);
or I_37563 (I640550,I640670,I641054);
DFFARX1 I_37564 (I641054,I2507,I640576,I640568,);
not I_37565 (I641154,I2514);
DFFARX1 I_37566 (I1018001,I2507,I641154,I641180,);
not I_37567 (I641188,I641180);
nand I_37568 (I641205,I1017998,I1018016);
and I_37569 (I641222,I641205,I1018013);
DFFARX1 I_37570 (I641222,I2507,I641154,I641248,);
not I_37571 (I641256,I1017995);
DFFARX1 I_37572 (I1017998,I2507,I641154,I641282,);
not I_37573 (I641290,I641282);
nor I_37574 (I641307,I641290,I641188);
and I_37575 (I641324,I641307,I1017995);
nor I_37576 (I641341,I641290,I641256);
nor I_37577 (I641137,I641248,I641341);
DFFARX1 I_37578 (I1018007,I2507,I641154,I641381,);
nor I_37579 (I641389,I641381,I641248);
not I_37580 (I641406,I641389);
not I_37581 (I641423,I641381);
nor I_37582 (I641440,I641423,I641324);
DFFARX1 I_37583 (I641440,I2507,I641154,I641140,);
nand I_37584 (I641471,I1018010,I1017995);
and I_37585 (I641488,I641471,I1018001);
DFFARX1 I_37586 (I641488,I2507,I641154,I641514,);
nor I_37587 (I641522,I641514,I641381);
DFFARX1 I_37588 (I641522,I2507,I641154,I641122,);
nand I_37589 (I641553,I641514,I641423);
nand I_37590 (I641131,I641406,I641553);
not I_37591 (I641584,I641514);
nor I_37592 (I641601,I641584,I641324);
DFFARX1 I_37593 (I641601,I2507,I641154,I641143,);
nor I_37594 (I641632,I1018004,I1017995);
or I_37595 (I641134,I641381,I641632);
nor I_37596 (I641125,I641514,I641632);
or I_37597 (I641128,I641248,I641632);
DFFARX1 I_37598 (I641632,I2507,I641154,I641146,);
not I_37599 (I641732,I2514);
DFFARX1 I_37600 (I452856,I2507,I641732,I641758,);
not I_37601 (I641766,I641758);
nand I_37602 (I641783,I452847,I452865);
and I_37603 (I641800,I641783,I452868);
DFFARX1 I_37604 (I641800,I2507,I641732,I641826,);
not I_37605 (I641834,I452862);
DFFARX1 I_37606 (I452850,I2507,I641732,I641860,);
not I_37607 (I641868,I641860);
nor I_37608 (I641885,I641868,I641766);
and I_37609 (I641902,I641885,I452862);
nor I_37610 (I641919,I641868,I641834);
nor I_37611 (I641715,I641826,I641919);
DFFARX1 I_37612 (I452859,I2507,I641732,I641959,);
nor I_37613 (I641967,I641959,I641826);
not I_37614 (I641984,I641967);
not I_37615 (I642001,I641959);
nor I_37616 (I642018,I642001,I641902);
DFFARX1 I_37617 (I642018,I2507,I641732,I641718,);
nand I_37618 (I642049,I452874,I452871);
and I_37619 (I642066,I642049,I452853);
DFFARX1 I_37620 (I642066,I2507,I641732,I642092,);
nor I_37621 (I642100,I642092,I641959);
DFFARX1 I_37622 (I642100,I2507,I641732,I641700,);
nand I_37623 (I642131,I642092,I642001);
nand I_37624 (I641709,I641984,I642131);
not I_37625 (I642162,I642092);
nor I_37626 (I642179,I642162,I641902);
DFFARX1 I_37627 (I642179,I2507,I641732,I641721,);
nor I_37628 (I642210,I452847,I452871);
or I_37629 (I641712,I641959,I642210);
nor I_37630 (I641703,I642092,I642210);
or I_37631 (I641706,I641826,I642210);
DFFARX1 I_37632 (I642210,I2507,I641732,I641724,);
not I_37633 (I642310,I2514);
DFFARX1 I_37634 (I167485,I2507,I642310,I642336,);
not I_37635 (I642344,I642336);
nand I_37636 (I642361,I167488,I167509);
and I_37637 (I642378,I642361,I167497);
DFFARX1 I_37638 (I642378,I2507,I642310,I642404,);
not I_37639 (I642412,I167494);
DFFARX1 I_37640 (I167485,I2507,I642310,I642438,);
not I_37641 (I642446,I642438);
nor I_37642 (I642463,I642446,I642344);
and I_37643 (I642480,I642463,I167494);
nor I_37644 (I642497,I642446,I642412);
nor I_37645 (I642293,I642404,I642497);
DFFARX1 I_37646 (I167503,I2507,I642310,I642537,);
nor I_37647 (I642545,I642537,I642404);
not I_37648 (I642562,I642545);
not I_37649 (I642579,I642537);
nor I_37650 (I642596,I642579,I642480);
DFFARX1 I_37651 (I642596,I2507,I642310,I642296,);
nand I_37652 (I642627,I167488,I167491);
and I_37653 (I642644,I642627,I167500);
DFFARX1 I_37654 (I642644,I2507,I642310,I642670,);
nor I_37655 (I642678,I642670,I642537);
DFFARX1 I_37656 (I642678,I2507,I642310,I642278,);
nand I_37657 (I642709,I642670,I642579);
nand I_37658 (I642287,I642562,I642709);
not I_37659 (I642740,I642670);
nor I_37660 (I642757,I642740,I642480);
DFFARX1 I_37661 (I642757,I2507,I642310,I642299,);
nor I_37662 (I642788,I167506,I167491);
or I_37663 (I642290,I642537,I642788);
nor I_37664 (I642281,I642670,I642788);
or I_37665 (I642284,I642404,I642788);
DFFARX1 I_37666 (I642788,I2507,I642310,I642302,);
not I_37667 (I642888,I2514);
DFFARX1 I_37668 (I385400,I2507,I642888,I642914,);
not I_37669 (I642922,I642914);
nand I_37670 (I642939,I385391,I385409);
and I_37671 (I642956,I642939,I385412);
DFFARX1 I_37672 (I642956,I2507,I642888,I642982,);
not I_37673 (I642990,I385406);
DFFARX1 I_37674 (I385394,I2507,I642888,I643016,);
not I_37675 (I643024,I643016);
nor I_37676 (I643041,I643024,I642922);
and I_37677 (I643058,I643041,I385406);
nor I_37678 (I643075,I643024,I642990);
nor I_37679 (I642871,I642982,I643075);
DFFARX1 I_37680 (I385403,I2507,I642888,I643115,);
nor I_37681 (I643123,I643115,I642982);
not I_37682 (I643140,I643123);
not I_37683 (I643157,I643115);
nor I_37684 (I643174,I643157,I643058);
DFFARX1 I_37685 (I643174,I2507,I642888,I642874,);
nand I_37686 (I643205,I385418,I385415);
and I_37687 (I643222,I643205,I385397);
DFFARX1 I_37688 (I643222,I2507,I642888,I643248,);
nor I_37689 (I643256,I643248,I643115);
DFFARX1 I_37690 (I643256,I2507,I642888,I642856,);
nand I_37691 (I643287,I643248,I643157);
nand I_37692 (I642865,I643140,I643287);
not I_37693 (I643318,I643248);
nor I_37694 (I643335,I643318,I643058);
DFFARX1 I_37695 (I643335,I2507,I642888,I642877,);
nor I_37696 (I643366,I385391,I385415);
or I_37697 (I642868,I643115,I643366);
nor I_37698 (I642859,I643248,I643366);
or I_37699 (I642862,I642982,I643366);
DFFARX1 I_37700 (I643366,I2507,I642888,I642880,);
not I_37701 (I643466,I2514);
DFFARX1 I_37702 (I29576,I2507,I643466,I643492,);
not I_37703 (I643500,I643492);
nand I_37704 (I643517,I29573,I29564);
and I_37705 (I643534,I643517,I29564);
DFFARX1 I_37706 (I643534,I2507,I643466,I643560,);
not I_37707 (I643568,I29567);
DFFARX1 I_37708 (I29582,I2507,I643466,I643594,);
not I_37709 (I643602,I643594);
nor I_37710 (I643619,I643602,I643500);
and I_37711 (I643636,I643619,I29567);
nor I_37712 (I643653,I643602,I643568);
nor I_37713 (I643449,I643560,I643653);
DFFARX1 I_37714 (I29567,I2507,I643466,I643693,);
nor I_37715 (I643701,I643693,I643560);
not I_37716 (I643718,I643701);
not I_37717 (I643735,I643693);
nor I_37718 (I643752,I643735,I643636);
DFFARX1 I_37719 (I643752,I2507,I643466,I643452,);
nand I_37720 (I643783,I29585,I29570);
and I_37721 (I643800,I643783,I29588);
DFFARX1 I_37722 (I643800,I2507,I643466,I643826,);
nor I_37723 (I643834,I643826,I643693);
DFFARX1 I_37724 (I643834,I2507,I643466,I643434,);
nand I_37725 (I643865,I643826,I643735);
nand I_37726 (I643443,I643718,I643865);
not I_37727 (I643896,I643826);
nor I_37728 (I643913,I643896,I643636);
DFFARX1 I_37729 (I643913,I2507,I643466,I643455,);
nor I_37730 (I643944,I29579,I29570);
or I_37731 (I643446,I643693,I643944);
nor I_37732 (I643437,I643826,I643944);
or I_37733 (I643440,I643560,I643944);
DFFARX1 I_37734 (I643944,I2507,I643466,I643458,);
not I_37735 (I644044,I2514);
DFFARX1 I_37736 (I1251490,I2507,I644044,I644070,);
not I_37737 (I644078,I644070);
nand I_37738 (I644095,I1251493,I1251502);
and I_37739 (I644112,I644095,I1251505);
DFFARX1 I_37740 (I644112,I2507,I644044,I644138,);
not I_37741 (I644146,I1251514);
DFFARX1 I_37742 (I1251496,I2507,I644044,I644172,);
not I_37743 (I644180,I644172);
nor I_37744 (I644197,I644180,I644078);
and I_37745 (I644214,I644197,I1251514);
nor I_37746 (I644231,I644180,I644146);
nor I_37747 (I644027,I644138,I644231);
DFFARX1 I_37748 (I1251493,I2507,I644044,I644271,);
nor I_37749 (I644279,I644271,I644138);
not I_37750 (I644296,I644279);
not I_37751 (I644313,I644271);
nor I_37752 (I644330,I644313,I644214);
DFFARX1 I_37753 (I644330,I2507,I644044,I644030,);
nand I_37754 (I644361,I1251511,I1251490);
and I_37755 (I644378,I644361,I1251508);
DFFARX1 I_37756 (I644378,I2507,I644044,I644404,);
nor I_37757 (I644412,I644404,I644271);
DFFARX1 I_37758 (I644412,I2507,I644044,I644012,);
nand I_37759 (I644443,I644404,I644313);
nand I_37760 (I644021,I644296,I644443);
not I_37761 (I644474,I644404);
nor I_37762 (I644491,I644474,I644214);
DFFARX1 I_37763 (I644491,I2507,I644044,I644033,);
nor I_37764 (I644522,I1251499,I1251490);
or I_37765 (I644024,I644271,I644522);
nor I_37766 (I644015,I644404,I644522);
or I_37767 (I644018,I644138,I644522);
DFFARX1 I_37768 (I644522,I2507,I644044,I644036,);
not I_37769 (I644622,I2514);
DFFARX1 I_37770 (I461016,I2507,I644622,I644648,);
not I_37771 (I644656,I644648);
nand I_37772 (I644673,I461007,I461025);
and I_37773 (I644690,I644673,I461028);
DFFARX1 I_37774 (I644690,I2507,I644622,I644716,);
not I_37775 (I644724,I461022);
DFFARX1 I_37776 (I461010,I2507,I644622,I644750,);
not I_37777 (I644758,I644750);
nor I_37778 (I644775,I644758,I644656);
and I_37779 (I644792,I644775,I461022);
nor I_37780 (I644809,I644758,I644724);
nor I_37781 (I644605,I644716,I644809);
DFFARX1 I_37782 (I461019,I2507,I644622,I644849,);
nor I_37783 (I644857,I644849,I644716);
not I_37784 (I644874,I644857);
not I_37785 (I644891,I644849);
nor I_37786 (I644908,I644891,I644792);
DFFARX1 I_37787 (I644908,I2507,I644622,I644608,);
nand I_37788 (I644939,I461034,I461031);
and I_37789 (I644956,I644939,I461013);
DFFARX1 I_37790 (I644956,I2507,I644622,I644982,);
nor I_37791 (I644990,I644982,I644849);
DFFARX1 I_37792 (I644990,I2507,I644622,I644590,);
nand I_37793 (I645021,I644982,I644891);
nand I_37794 (I644599,I644874,I645021);
not I_37795 (I645052,I644982);
nor I_37796 (I645069,I645052,I644792);
DFFARX1 I_37797 (I645069,I2507,I644622,I644611,);
nor I_37798 (I645100,I461007,I461031);
or I_37799 (I644602,I644849,I645100);
nor I_37800 (I644593,I644982,I645100);
or I_37801 (I644596,I644716,I645100);
DFFARX1 I_37802 (I645100,I2507,I644622,I644614,);
not I_37803 (I645200,I2514);
DFFARX1 I_37804 (I1337469,I2507,I645200,I645226,);
not I_37805 (I645234,I645226);
nand I_37806 (I645251,I1337454,I1337442);
and I_37807 (I645268,I645251,I1337457);
DFFARX1 I_37808 (I645268,I2507,I645200,I645294,);
not I_37809 (I645302,I1337442);
DFFARX1 I_37810 (I1337460,I2507,I645200,I645328,);
not I_37811 (I645336,I645328);
nor I_37812 (I645353,I645336,I645234);
and I_37813 (I645370,I645353,I1337442);
nor I_37814 (I645387,I645336,I645302);
nor I_37815 (I645183,I645294,I645387);
DFFARX1 I_37816 (I1337448,I2507,I645200,I645427,);
nor I_37817 (I645435,I645427,I645294);
not I_37818 (I645452,I645435);
not I_37819 (I645469,I645427);
nor I_37820 (I645486,I645469,I645370);
DFFARX1 I_37821 (I645486,I2507,I645200,I645186,);
nand I_37822 (I645517,I1337445,I1337451);
and I_37823 (I645534,I645517,I1337466);
DFFARX1 I_37824 (I645534,I2507,I645200,I645560,);
nor I_37825 (I645568,I645560,I645427);
DFFARX1 I_37826 (I645568,I2507,I645200,I645168,);
nand I_37827 (I645599,I645560,I645469);
nand I_37828 (I645177,I645452,I645599);
not I_37829 (I645630,I645560);
nor I_37830 (I645647,I645630,I645370);
DFFARX1 I_37831 (I645647,I2507,I645200,I645189,);
nor I_37832 (I645678,I1337463,I1337451);
or I_37833 (I645180,I645427,I645678);
nor I_37834 (I645171,I645560,I645678);
or I_37835 (I645174,I645294,I645678);
DFFARX1 I_37836 (I645678,I2507,I645200,I645192,);
not I_37837 (I645778,I2514);
DFFARX1 I_37838 (I1348774,I2507,I645778,I645804,);
not I_37839 (I645812,I645804);
nand I_37840 (I645829,I1348759,I1348747);
and I_37841 (I645846,I645829,I1348762);
DFFARX1 I_37842 (I645846,I2507,I645778,I645872,);
not I_37843 (I645880,I1348747);
DFFARX1 I_37844 (I1348765,I2507,I645778,I645906,);
not I_37845 (I645914,I645906);
nor I_37846 (I645931,I645914,I645812);
and I_37847 (I645948,I645931,I1348747);
nor I_37848 (I645965,I645914,I645880);
nor I_37849 (I645761,I645872,I645965);
DFFARX1 I_37850 (I1348753,I2507,I645778,I646005,);
nor I_37851 (I646013,I646005,I645872);
not I_37852 (I646030,I646013);
not I_37853 (I646047,I646005);
nor I_37854 (I646064,I646047,I645948);
DFFARX1 I_37855 (I646064,I2507,I645778,I645764,);
nand I_37856 (I646095,I1348750,I1348756);
and I_37857 (I646112,I646095,I1348771);
DFFARX1 I_37858 (I646112,I2507,I645778,I646138,);
nor I_37859 (I646146,I646138,I646005);
DFFARX1 I_37860 (I646146,I2507,I645778,I645746,);
nand I_37861 (I646177,I646138,I646047);
nand I_37862 (I645755,I646030,I646177);
not I_37863 (I646208,I646138);
nor I_37864 (I646225,I646208,I645948);
DFFARX1 I_37865 (I646225,I2507,I645778,I645767,);
nor I_37866 (I646256,I1348768,I1348756);
or I_37867 (I645758,I646005,I646256);
nor I_37868 (I645749,I646138,I646256);
or I_37869 (I645752,I645872,I646256);
DFFARX1 I_37870 (I646256,I2507,I645778,I645770,);
not I_37871 (I646356,I2514);
DFFARX1 I_37872 (I1269204,I2507,I646356,I646382,);
not I_37873 (I646390,I646382);
nand I_37874 (I646407,I1269228,I1269210);
and I_37875 (I646424,I646407,I1269216);
DFFARX1 I_37876 (I646424,I2507,I646356,I646450,);
not I_37877 (I646458,I1269222);
DFFARX1 I_37878 (I1269207,I2507,I646356,I646484,);
not I_37879 (I646492,I646484);
nor I_37880 (I646509,I646492,I646390);
and I_37881 (I646526,I646509,I1269222);
nor I_37882 (I646543,I646492,I646458);
nor I_37883 (I646339,I646450,I646543);
DFFARX1 I_37884 (I1269219,I2507,I646356,I646583,);
nor I_37885 (I646591,I646583,I646450);
not I_37886 (I646608,I646591);
not I_37887 (I646625,I646583);
nor I_37888 (I646642,I646625,I646526);
DFFARX1 I_37889 (I646642,I2507,I646356,I646342,);
nand I_37890 (I646673,I1269225,I1269213);
and I_37891 (I646690,I646673,I1269207);
DFFARX1 I_37892 (I646690,I2507,I646356,I646716,);
nor I_37893 (I646724,I646716,I646583);
DFFARX1 I_37894 (I646724,I2507,I646356,I646324,);
nand I_37895 (I646755,I646716,I646625);
nand I_37896 (I646333,I646608,I646755);
not I_37897 (I646786,I646716);
nor I_37898 (I646803,I646786,I646526);
DFFARX1 I_37899 (I646803,I2507,I646356,I646345,);
nor I_37900 (I646834,I1269204,I1269213);
or I_37901 (I646336,I646583,I646834);
nor I_37902 (I646327,I646716,I646834);
or I_37903 (I646330,I646450,I646834);
DFFARX1 I_37904 (I646834,I2507,I646356,I646348,);
not I_37905 (I646934,I2514);
DFFARX1 I_37906 (I373532,I2507,I646934,I646960,);
not I_37907 (I646968,I646960);
nand I_37908 (I646985,I373535,I373511);
and I_37909 (I647002,I646985,I373508);
DFFARX1 I_37910 (I647002,I2507,I646934,I647028,);
not I_37911 (I647036,I373514);
DFFARX1 I_37912 (I373508,I2507,I646934,I647062,);
not I_37913 (I647070,I647062);
nor I_37914 (I647087,I647070,I646968);
and I_37915 (I647104,I647087,I373514);
nor I_37916 (I647121,I647070,I647036);
nor I_37917 (I646917,I647028,I647121);
DFFARX1 I_37918 (I373517,I2507,I646934,I647161,);
nor I_37919 (I647169,I647161,I647028);
not I_37920 (I647186,I647169);
not I_37921 (I647203,I647161);
nor I_37922 (I647220,I647203,I647104);
DFFARX1 I_37923 (I647220,I2507,I646934,I646920,);
nand I_37924 (I647251,I373520,I373529);
and I_37925 (I647268,I647251,I373526);
DFFARX1 I_37926 (I647268,I2507,I646934,I647294,);
nor I_37927 (I647302,I647294,I647161);
DFFARX1 I_37928 (I647302,I2507,I646934,I646902,);
nand I_37929 (I647333,I647294,I647203);
nand I_37930 (I646911,I647186,I647333);
not I_37931 (I647364,I647294);
nor I_37932 (I647381,I647364,I647104);
DFFARX1 I_37933 (I647381,I2507,I646934,I646923,);
nor I_37934 (I647412,I373523,I373529);
or I_37935 (I646914,I647161,I647412);
nor I_37936 (I646905,I647294,I647412);
or I_37937 (I646908,I647028,I647412);
DFFARX1 I_37938 (I647412,I2507,I646934,I646926,);
not I_37939 (I647512,I2514);
DFFARX1 I_37940 (I626672,I2507,I647512,I647538,);
not I_37941 (I647546,I647538);
nand I_37942 (I647563,I626681,I626690);
and I_37943 (I647580,I647563,I626696);
DFFARX1 I_37944 (I647580,I2507,I647512,I647606,);
not I_37945 (I647614,I626693);
DFFARX1 I_37946 (I626678,I2507,I647512,I647640,);
not I_37947 (I647648,I647640);
nor I_37948 (I647665,I647648,I647546);
and I_37949 (I647682,I647665,I626693);
nor I_37950 (I647699,I647648,I647614);
nor I_37951 (I647495,I647606,I647699);
DFFARX1 I_37952 (I626687,I2507,I647512,I647739,);
nor I_37953 (I647747,I647739,I647606);
not I_37954 (I647764,I647747);
not I_37955 (I647781,I647739);
nor I_37956 (I647798,I647781,I647682);
DFFARX1 I_37957 (I647798,I2507,I647512,I647498,);
nand I_37958 (I647829,I626684,I626675);
and I_37959 (I647846,I647829,I626672);
DFFARX1 I_37960 (I647846,I2507,I647512,I647872,);
nor I_37961 (I647880,I647872,I647739);
DFFARX1 I_37962 (I647880,I2507,I647512,I647480,);
nand I_37963 (I647911,I647872,I647781);
nand I_37964 (I647489,I647764,I647911);
not I_37965 (I647942,I647872);
nor I_37966 (I647959,I647942,I647682);
DFFARX1 I_37967 (I647959,I2507,I647512,I647501,);
nor I_37968 (I647990,I626675,I626675);
or I_37969 (I647492,I647739,I647990);
nor I_37970 (I647483,I647872,I647990);
or I_37971 (I647486,I647606,I647990);
DFFARX1 I_37972 (I647990,I2507,I647512,I647504,);
not I_37973 (I648090,I2514);
DFFARX1 I_37974 (I1367814,I2507,I648090,I648116,);
not I_37975 (I648124,I648116);
nand I_37976 (I648141,I1367799,I1367787);
and I_37977 (I648158,I648141,I1367802);
DFFARX1 I_37978 (I648158,I2507,I648090,I648184,);
not I_37979 (I648192,I1367787);
DFFARX1 I_37980 (I1367805,I2507,I648090,I648218,);
not I_37981 (I648226,I648218);
nor I_37982 (I648243,I648226,I648124);
and I_37983 (I648260,I648243,I1367787);
nor I_37984 (I648277,I648226,I648192);
nor I_37985 (I648073,I648184,I648277);
DFFARX1 I_37986 (I1367793,I2507,I648090,I648317,);
nor I_37987 (I648325,I648317,I648184);
not I_37988 (I648342,I648325);
not I_37989 (I648359,I648317);
nor I_37990 (I648376,I648359,I648260);
DFFARX1 I_37991 (I648376,I2507,I648090,I648076,);
nand I_37992 (I648407,I1367790,I1367796);
and I_37993 (I648424,I648407,I1367811);
DFFARX1 I_37994 (I648424,I2507,I648090,I648450,);
nor I_37995 (I648458,I648450,I648317);
DFFARX1 I_37996 (I648458,I2507,I648090,I648058,);
nand I_37997 (I648489,I648450,I648359);
nand I_37998 (I648067,I648342,I648489);
not I_37999 (I648520,I648450);
nor I_38000 (I648537,I648520,I648260);
DFFARX1 I_38001 (I648537,I2507,I648090,I648079,);
nor I_38002 (I648568,I1367808,I1367796);
or I_38003 (I648070,I648317,I648568);
nor I_38004 (I648061,I648450,I648568);
or I_38005 (I648064,I648184,I648568);
DFFARX1 I_38006 (I648568,I2507,I648090,I648082,);
not I_38007 (I648668,I2514);
DFFARX1 I_38008 (I89118,I2507,I648668,I648694,);
not I_38009 (I648702,I648694);
nand I_38010 (I648719,I89127,I89136);
and I_38011 (I648736,I648719,I89115);
DFFARX1 I_38012 (I648736,I2507,I648668,I648762,);
not I_38013 (I648770,I89118);
DFFARX1 I_38014 (I89133,I2507,I648668,I648796,);
not I_38015 (I648804,I648796);
nor I_38016 (I648821,I648804,I648702);
and I_38017 (I648838,I648821,I89118);
nor I_38018 (I648855,I648804,I648770);
nor I_38019 (I648651,I648762,I648855);
DFFARX1 I_38020 (I89124,I2507,I648668,I648895,);
nor I_38021 (I648903,I648895,I648762);
not I_38022 (I648920,I648903);
not I_38023 (I648937,I648895);
nor I_38024 (I648954,I648937,I648838);
DFFARX1 I_38025 (I648954,I2507,I648668,I648654,);
nand I_38026 (I648985,I89139,I89115);
and I_38027 (I649002,I648985,I89121);
DFFARX1 I_38028 (I649002,I2507,I648668,I649028,);
nor I_38029 (I649036,I649028,I648895);
DFFARX1 I_38030 (I649036,I2507,I648668,I648636,);
nand I_38031 (I649067,I649028,I648937);
nand I_38032 (I648645,I648920,I649067);
not I_38033 (I649098,I649028);
nor I_38034 (I649115,I649098,I648838);
DFFARX1 I_38035 (I649115,I2507,I648668,I648657,);
nor I_38036 (I649146,I89130,I89115);
or I_38037 (I648648,I648895,I649146);
nor I_38038 (I648639,I649028,I649146);
or I_38039 (I648642,I648762,I649146);
DFFARX1 I_38040 (I649146,I2507,I648668,I648660,);
not I_38041 (I649246,I2514);
DFFARX1 I_38042 (I269186,I2507,I649246,I649272,);
not I_38043 (I649280,I649272);
nand I_38044 (I649297,I269189,I269165);
and I_38045 (I649314,I649297,I269162);
DFFARX1 I_38046 (I649314,I2507,I649246,I649340,);
not I_38047 (I649348,I269168);
DFFARX1 I_38048 (I269162,I2507,I649246,I649374,);
not I_38049 (I649382,I649374);
nor I_38050 (I649399,I649382,I649280);
and I_38051 (I649416,I649399,I269168);
nor I_38052 (I649433,I649382,I649348);
nor I_38053 (I649229,I649340,I649433);
DFFARX1 I_38054 (I269171,I2507,I649246,I649473,);
nor I_38055 (I649481,I649473,I649340);
not I_38056 (I649498,I649481);
not I_38057 (I649515,I649473);
nor I_38058 (I649532,I649515,I649416);
DFFARX1 I_38059 (I649532,I2507,I649246,I649232,);
nand I_38060 (I649563,I269174,I269183);
and I_38061 (I649580,I649563,I269180);
DFFARX1 I_38062 (I649580,I2507,I649246,I649606,);
nor I_38063 (I649614,I649606,I649473);
DFFARX1 I_38064 (I649614,I2507,I649246,I649214,);
nand I_38065 (I649645,I649606,I649515);
nand I_38066 (I649223,I649498,I649645);
not I_38067 (I649676,I649606);
nor I_38068 (I649693,I649676,I649416);
DFFARX1 I_38069 (I649693,I2507,I649246,I649235,);
nor I_38070 (I649724,I269177,I269183);
or I_38071 (I649226,I649473,I649724);
nor I_38072 (I649217,I649606,I649724);
or I_38073 (I649220,I649340,I649724);
DFFARX1 I_38074 (I649724,I2507,I649246,I649238,);
not I_38075 (I649824,I2514);
DFFARX1 I_38076 (I919895,I2507,I649824,I649850,);
not I_38077 (I649858,I649850);
nand I_38078 (I649875,I919871,I919886);
and I_38079 (I649892,I649875,I919898);
DFFARX1 I_38080 (I649892,I2507,I649824,I649918,);
not I_38081 (I649926,I919883);
DFFARX1 I_38082 (I919874,I2507,I649824,I649952,);
not I_38083 (I649960,I649952);
nor I_38084 (I649977,I649960,I649858);
and I_38085 (I649994,I649977,I919883);
nor I_38086 (I650011,I649960,I649926);
nor I_38087 (I649807,I649918,I650011);
DFFARX1 I_38088 (I919871,I2507,I649824,I650051,);
nor I_38089 (I650059,I650051,I649918);
not I_38090 (I650076,I650059);
not I_38091 (I650093,I650051);
nor I_38092 (I650110,I650093,I649994);
DFFARX1 I_38093 (I650110,I2507,I649824,I649810,);
nand I_38094 (I650141,I919889,I919880);
and I_38095 (I650158,I650141,I919892);
DFFARX1 I_38096 (I650158,I2507,I649824,I650184,);
nor I_38097 (I650192,I650184,I650051);
DFFARX1 I_38098 (I650192,I2507,I649824,I649792,);
nand I_38099 (I650223,I650184,I650093);
nand I_38100 (I649801,I650076,I650223);
not I_38101 (I650254,I650184);
nor I_38102 (I650271,I650254,I649994);
DFFARX1 I_38103 (I650271,I2507,I649824,I649813,);
nor I_38104 (I650302,I919877,I919880);
or I_38105 (I649804,I650051,I650302);
nor I_38106 (I649795,I650184,I650302);
or I_38107 (I649798,I649918,I650302);
DFFARX1 I_38108 (I650302,I2507,I649824,I649816,);
not I_38109 (I650402,I2514);
DFFARX1 I_38110 (I1079196,I2507,I650402,I650428,);
not I_38111 (I650436,I650428);
nand I_38112 (I650453,I1079178,I1079190);
and I_38113 (I650470,I650453,I1079193);
DFFARX1 I_38114 (I650470,I2507,I650402,I650496,);
not I_38115 (I650504,I1079187);
DFFARX1 I_38116 (I1079184,I2507,I650402,I650530,);
not I_38117 (I650538,I650530);
nor I_38118 (I650555,I650538,I650436);
and I_38119 (I650572,I650555,I1079187);
nor I_38120 (I650589,I650538,I650504);
nor I_38121 (I650385,I650496,I650589);
DFFARX1 I_38122 (I1079202,I2507,I650402,I650629,);
nor I_38123 (I650637,I650629,I650496);
not I_38124 (I650654,I650637);
not I_38125 (I650671,I650629);
nor I_38126 (I650688,I650671,I650572);
DFFARX1 I_38127 (I650688,I2507,I650402,I650388,);
nand I_38128 (I650719,I1079181,I1079181);
and I_38129 (I650736,I650719,I1079178);
DFFARX1 I_38130 (I650736,I2507,I650402,I650762,);
nor I_38131 (I650770,I650762,I650629);
DFFARX1 I_38132 (I650770,I2507,I650402,I650370,);
nand I_38133 (I650801,I650762,I650671);
nand I_38134 (I650379,I650654,I650801);
not I_38135 (I650832,I650762);
nor I_38136 (I650849,I650832,I650572);
DFFARX1 I_38137 (I650849,I2507,I650402,I650391,);
nor I_38138 (I650880,I1079199,I1079181);
or I_38139 (I650382,I650629,I650880);
nor I_38140 (I650373,I650762,I650880);
or I_38141 (I650376,I650496,I650880);
DFFARX1 I_38142 (I650880,I2507,I650402,I650394,);
not I_38143 (I650980,I2514);
DFFARX1 I_38144 (I301860,I2507,I650980,I651006,);
not I_38145 (I651014,I651006);
nand I_38146 (I651031,I301863,I301839);
and I_38147 (I651048,I651031,I301836);
DFFARX1 I_38148 (I651048,I2507,I650980,I651074,);
not I_38149 (I651082,I301842);
DFFARX1 I_38150 (I301836,I2507,I650980,I651108,);
not I_38151 (I651116,I651108);
nor I_38152 (I651133,I651116,I651014);
and I_38153 (I651150,I651133,I301842);
nor I_38154 (I651167,I651116,I651082);
nor I_38155 (I650963,I651074,I651167);
DFFARX1 I_38156 (I301845,I2507,I650980,I651207,);
nor I_38157 (I651215,I651207,I651074);
not I_38158 (I651232,I651215);
not I_38159 (I651249,I651207);
nor I_38160 (I651266,I651249,I651150);
DFFARX1 I_38161 (I651266,I2507,I650980,I650966,);
nand I_38162 (I651297,I301848,I301857);
and I_38163 (I651314,I651297,I301854);
DFFARX1 I_38164 (I651314,I2507,I650980,I651340,);
nor I_38165 (I651348,I651340,I651207);
DFFARX1 I_38166 (I651348,I2507,I650980,I650948,);
nand I_38167 (I651379,I651340,I651249);
nand I_38168 (I650957,I651232,I651379);
not I_38169 (I651410,I651340);
nor I_38170 (I651427,I651410,I651150);
DFFARX1 I_38171 (I651427,I2507,I650980,I650969,);
nor I_38172 (I651458,I301851,I301857);
or I_38173 (I650960,I651207,I651458);
nor I_38174 (I650951,I651340,I651458);
or I_38175 (I650954,I651074,I651458);
DFFARX1 I_38176 (I651458,I2507,I650980,I650972,);
not I_38177 (I651558,I2514);
DFFARX1 I_38178 (I407160,I2507,I651558,I651584,);
not I_38179 (I651592,I651584);
nand I_38180 (I651609,I407151,I407169);
and I_38181 (I651626,I651609,I407172);
DFFARX1 I_38182 (I651626,I2507,I651558,I651652,);
not I_38183 (I651660,I407166);
DFFARX1 I_38184 (I407154,I2507,I651558,I651686,);
not I_38185 (I651694,I651686);
nor I_38186 (I651711,I651694,I651592);
and I_38187 (I651728,I651711,I407166);
nor I_38188 (I651745,I651694,I651660);
nor I_38189 (I651541,I651652,I651745);
DFFARX1 I_38190 (I407163,I2507,I651558,I651785,);
nor I_38191 (I651793,I651785,I651652);
not I_38192 (I651810,I651793);
not I_38193 (I651827,I651785);
nor I_38194 (I651844,I651827,I651728);
DFFARX1 I_38195 (I651844,I2507,I651558,I651544,);
nand I_38196 (I651875,I407178,I407175);
and I_38197 (I651892,I651875,I407157);
DFFARX1 I_38198 (I651892,I2507,I651558,I651918,);
nor I_38199 (I651926,I651918,I651785);
DFFARX1 I_38200 (I651926,I2507,I651558,I651526,);
nand I_38201 (I651957,I651918,I651827);
nand I_38202 (I651535,I651810,I651957);
not I_38203 (I651988,I651918);
nor I_38204 (I652005,I651988,I651728);
DFFARX1 I_38205 (I652005,I2507,I651558,I651547,);
nor I_38206 (I652036,I407151,I407175);
or I_38207 (I651538,I651785,I652036);
nor I_38208 (I651529,I651918,I652036);
or I_38209 (I651532,I651652,I652036);
DFFARX1 I_38210 (I652036,I2507,I651558,I651550,);
not I_38211 (I652136,I2514);
DFFARX1 I_38212 (I62768,I2507,I652136,I652162,);
not I_38213 (I652170,I652162);
nand I_38214 (I652187,I62777,I62786);
and I_38215 (I652204,I652187,I62765);
DFFARX1 I_38216 (I652204,I2507,I652136,I652230,);
not I_38217 (I652238,I62768);
DFFARX1 I_38218 (I62783,I2507,I652136,I652264,);
not I_38219 (I652272,I652264);
nor I_38220 (I652289,I652272,I652170);
and I_38221 (I652306,I652289,I62768);
nor I_38222 (I652323,I652272,I652238);
nor I_38223 (I652119,I652230,I652323);
DFFARX1 I_38224 (I62774,I2507,I652136,I652363,);
nor I_38225 (I652371,I652363,I652230);
not I_38226 (I652388,I652371);
not I_38227 (I652405,I652363);
nor I_38228 (I652422,I652405,I652306);
DFFARX1 I_38229 (I652422,I2507,I652136,I652122,);
nand I_38230 (I652453,I62789,I62765);
and I_38231 (I652470,I652453,I62771);
DFFARX1 I_38232 (I652470,I2507,I652136,I652496,);
nor I_38233 (I652504,I652496,I652363);
DFFARX1 I_38234 (I652504,I2507,I652136,I652104,);
nand I_38235 (I652535,I652496,I652405);
nand I_38236 (I652113,I652388,I652535);
not I_38237 (I652566,I652496);
nor I_38238 (I652583,I652566,I652306);
DFFARX1 I_38239 (I652583,I2507,I652136,I652125,);
nor I_38240 (I652614,I62780,I62765);
or I_38241 (I652116,I652363,I652614);
nor I_38242 (I652107,I652496,I652614);
or I_38243 (I652110,I652230,I652614);
DFFARX1 I_38244 (I652614,I2507,I652136,I652128,);
not I_38245 (I652714,I2514);
DFFARX1 I_38246 (I438168,I2507,I652714,I652740,);
not I_38247 (I652748,I652740);
nand I_38248 (I652765,I438159,I438177);
and I_38249 (I652782,I652765,I438180);
DFFARX1 I_38250 (I652782,I2507,I652714,I652808,);
not I_38251 (I652816,I438174);
DFFARX1 I_38252 (I438162,I2507,I652714,I652842,);
not I_38253 (I652850,I652842);
nor I_38254 (I652867,I652850,I652748);
and I_38255 (I652884,I652867,I438174);
nor I_38256 (I652901,I652850,I652816);
nor I_38257 (I652697,I652808,I652901);
DFFARX1 I_38258 (I438171,I2507,I652714,I652941,);
nor I_38259 (I652949,I652941,I652808);
not I_38260 (I652966,I652949);
not I_38261 (I652983,I652941);
nor I_38262 (I653000,I652983,I652884);
DFFARX1 I_38263 (I653000,I2507,I652714,I652700,);
nand I_38264 (I653031,I438186,I438183);
and I_38265 (I653048,I653031,I438165);
DFFARX1 I_38266 (I653048,I2507,I652714,I653074,);
nor I_38267 (I653082,I653074,I652941);
DFFARX1 I_38268 (I653082,I2507,I652714,I652682,);
nand I_38269 (I653113,I653074,I652983);
nand I_38270 (I652691,I652966,I653113);
not I_38271 (I653144,I653074);
nor I_38272 (I653161,I653144,I652884);
DFFARX1 I_38273 (I653161,I2507,I652714,I652703,);
nor I_38274 (I653192,I438159,I438183);
or I_38275 (I652694,I652941,I653192);
nor I_38276 (I652685,I653074,I653192);
or I_38277 (I652688,I652808,I653192);
DFFARX1 I_38278 (I653192,I2507,I652714,I652706,);
not I_38279 (I653292,I2514);
DFFARX1 I_38280 (I430552,I2507,I653292,I653318,);
not I_38281 (I653326,I653318);
nand I_38282 (I653343,I430543,I430561);
and I_38283 (I653360,I653343,I430564);
DFFARX1 I_38284 (I653360,I2507,I653292,I653386,);
not I_38285 (I653394,I430558);
DFFARX1 I_38286 (I430546,I2507,I653292,I653420,);
not I_38287 (I653428,I653420);
nor I_38288 (I653445,I653428,I653326);
and I_38289 (I653462,I653445,I430558);
nor I_38290 (I653479,I653428,I653394);
nor I_38291 (I653275,I653386,I653479);
DFFARX1 I_38292 (I430555,I2507,I653292,I653519,);
nor I_38293 (I653527,I653519,I653386);
not I_38294 (I653544,I653527);
not I_38295 (I653561,I653519);
nor I_38296 (I653578,I653561,I653462);
DFFARX1 I_38297 (I653578,I2507,I653292,I653278,);
nand I_38298 (I653609,I430570,I430567);
and I_38299 (I653626,I653609,I430549);
DFFARX1 I_38300 (I653626,I2507,I653292,I653652,);
nor I_38301 (I653660,I653652,I653519);
DFFARX1 I_38302 (I653660,I2507,I653292,I653260,);
nand I_38303 (I653691,I653652,I653561);
nand I_38304 (I653269,I653544,I653691);
not I_38305 (I653722,I653652);
nor I_38306 (I653739,I653722,I653462);
DFFARX1 I_38307 (I653739,I2507,I653292,I653281,);
nor I_38308 (I653770,I430543,I430567);
or I_38309 (I653272,I653519,I653770);
nor I_38310 (I653263,I653652,I653770);
or I_38311 (I653266,I653386,I653770);
DFFARX1 I_38312 (I653770,I2507,I653292,I653284,);
not I_38313 (I653870,I2514);
DFFARX1 I_38314 (I833883,I2507,I653870,I653896,);
not I_38315 (I653904,I653896);
nand I_38316 (I653921,I833871,I833889);
and I_38317 (I653938,I653921,I833886);
DFFARX1 I_38318 (I653938,I2507,I653870,I653964,);
not I_38319 (I653972,I833877);
DFFARX1 I_38320 (I833874,I2507,I653870,I653998,);
not I_38321 (I654006,I653998);
nor I_38322 (I654023,I654006,I653904);
and I_38323 (I654040,I654023,I833877);
nor I_38324 (I654057,I654006,I653972);
nor I_38325 (I653853,I653964,I654057);
DFFARX1 I_38326 (I833868,I2507,I653870,I654097,);
nor I_38327 (I654105,I654097,I653964);
not I_38328 (I654122,I654105);
not I_38329 (I654139,I654097);
nor I_38330 (I654156,I654139,I654040);
DFFARX1 I_38331 (I654156,I2507,I653870,I653856,);
nand I_38332 (I654187,I833868,I833871);
and I_38333 (I654204,I654187,I833874);
DFFARX1 I_38334 (I654204,I2507,I653870,I654230,);
nor I_38335 (I654238,I654230,I654097);
DFFARX1 I_38336 (I654238,I2507,I653870,I653838,);
nand I_38337 (I654269,I654230,I654139);
nand I_38338 (I653847,I654122,I654269);
not I_38339 (I654300,I654230);
nor I_38340 (I654317,I654300,I654040);
DFFARX1 I_38341 (I654317,I2507,I653870,I653859,);
nor I_38342 (I654348,I833880,I833871);
or I_38343 (I653850,I654097,I654348);
nor I_38344 (I653841,I654230,I654348);
or I_38345 (I653844,I653964,I654348);
DFFARX1 I_38346 (I654348,I2507,I653870,I653862,);
not I_38347 (I654448,I2514);
DFFARX1 I_38348 (I2523,I2507,I654448,I654474,);
not I_38349 (I654482,I654474);
nand I_38350 (I654499,I2526,I2538);
and I_38351 (I654516,I654499,I2517);
DFFARX1 I_38352 (I654516,I2507,I654448,I654542,);
not I_38353 (I654550,I2517);
DFFARX1 I_38354 (I2520,I2507,I654448,I654576,);
not I_38355 (I654584,I654576);
nor I_38356 (I654601,I654584,I654482);
and I_38357 (I654618,I654601,I2517);
nor I_38358 (I654635,I654584,I654550);
nor I_38359 (I654431,I654542,I654635);
DFFARX1 I_38360 (I2532,I2507,I654448,I654675,);
nor I_38361 (I654683,I654675,I654542);
not I_38362 (I654700,I654683);
not I_38363 (I654717,I654675);
nor I_38364 (I654734,I654717,I654618);
DFFARX1 I_38365 (I654734,I2507,I654448,I654434,);
nand I_38366 (I654765,I2535,I2520);
and I_38367 (I654782,I654765,I2529);
DFFARX1 I_38368 (I654782,I2507,I654448,I654808,);
nor I_38369 (I654816,I654808,I654675);
DFFARX1 I_38370 (I654816,I2507,I654448,I654416,);
nand I_38371 (I654847,I654808,I654717);
nand I_38372 (I654425,I654700,I654847);
not I_38373 (I654878,I654808);
nor I_38374 (I654895,I654878,I654618);
DFFARX1 I_38375 (I654895,I2507,I654448,I654437,);
nor I_38376 (I654926,I2523,I2520);
or I_38377 (I654428,I654675,I654926);
nor I_38378 (I654419,I654808,I654926);
or I_38379 (I654422,I654542,I654926);
DFFARX1 I_38380 (I654926,I2507,I654448,I654440,);
not I_38381 (I655026,I2514);
DFFARX1 I_38382 (I579854,I2507,I655026,I655052,);
not I_38383 (I655060,I655052);
nand I_38384 (I655077,I579863,I579872);
and I_38385 (I655094,I655077,I579878);
DFFARX1 I_38386 (I655094,I2507,I655026,I655120,);
not I_38387 (I655128,I579875);
DFFARX1 I_38388 (I579860,I2507,I655026,I655154,);
not I_38389 (I655162,I655154);
nor I_38390 (I655179,I655162,I655060);
and I_38391 (I655196,I655179,I579875);
nor I_38392 (I655213,I655162,I655128);
nor I_38393 (I655009,I655120,I655213);
DFFARX1 I_38394 (I579869,I2507,I655026,I655253,);
nor I_38395 (I655261,I655253,I655120);
not I_38396 (I655278,I655261);
not I_38397 (I655295,I655253);
nor I_38398 (I655312,I655295,I655196);
DFFARX1 I_38399 (I655312,I2507,I655026,I655012,);
nand I_38400 (I655343,I579866,I579857);
and I_38401 (I655360,I655343,I579854);
DFFARX1 I_38402 (I655360,I2507,I655026,I655386,);
nor I_38403 (I655394,I655386,I655253);
DFFARX1 I_38404 (I655394,I2507,I655026,I654994,);
nand I_38405 (I655425,I655386,I655295);
nand I_38406 (I655003,I655278,I655425);
not I_38407 (I655456,I655386);
nor I_38408 (I655473,I655456,I655196);
DFFARX1 I_38409 (I655473,I2507,I655026,I655015,);
nor I_38410 (I655504,I579857,I579857);
or I_38411 (I655006,I655253,I655504);
nor I_38412 (I654997,I655386,I655504);
or I_38413 (I655000,I655120,I655504);
DFFARX1 I_38414 (I655504,I2507,I655026,I655018,);
not I_38415 (I655604,I2514);
DFFARX1 I_38416 (I458840,I2507,I655604,I655630,);
not I_38417 (I655638,I655630);
nand I_38418 (I655655,I458831,I458849);
and I_38419 (I655672,I655655,I458852);
DFFARX1 I_38420 (I655672,I2507,I655604,I655698,);
not I_38421 (I655706,I458846);
DFFARX1 I_38422 (I458834,I2507,I655604,I655732,);
not I_38423 (I655740,I655732);
nor I_38424 (I655757,I655740,I655638);
and I_38425 (I655774,I655757,I458846);
nor I_38426 (I655791,I655740,I655706);
nor I_38427 (I655587,I655698,I655791);
DFFARX1 I_38428 (I458843,I2507,I655604,I655831,);
nor I_38429 (I655839,I655831,I655698);
not I_38430 (I655856,I655839);
not I_38431 (I655873,I655831);
nor I_38432 (I655890,I655873,I655774);
DFFARX1 I_38433 (I655890,I2507,I655604,I655590,);
nand I_38434 (I655921,I458858,I458855);
and I_38435 (I655938,I655921,I458837);
DFFARX1 I_38436 (I655938,I2507,I655604,I655964,);
nor I_38437 (I655972,I655964,I655831);
DFFARX1 I_38438 (I655972,I2507,I655604,I655572,);
nand I_38439 (I656003,I655964,I655873);
nand I_38440 (I655581,I655856,I656003);
not I_38441 (I656034,I655964);
nor I_38442 (I656051,I656034,I655774);
DFFARX1 I_38443 (I656051,I2507,I655604,I655593,);
nor I_38444 (I656082,I458831,I458855);
or I_38445 (I655584,I655831,I656082);
nor I_38446 (I655575,I655964,I656082);
or I_38447 (I655578,I655698,I656082);
DFFARX1 I_38448 (I656082,I2507,I655604,I655596,);
not I_38449 (I656182,I2514);
DFFARX1 I_38450 (I1311289,I2507,I656182,I656208,);
not I_38451 (I656216,I656208);
nand I_38452 (I656233,I1311274,I1311262);
and I_38453 (I656250,I656233,I1311277);
DFFARX1 I_38454 (I656250,I2507,I656182,I656276,);
not I_38455 (I656284,I1311262);
DFFARX1 I_38456 (I1311280,I2507,I656182,I656310,);
not I_38457 (I656318,I656310);
nor I_38458 (I656335,I656318,I656216);
and I_38459 (I656352,I656335,I1311262);
nor I_38460 (I656369,I656318,I656284);
nor I_38461 (I656165,I656276,I656369);
DFFARX1 I_38462 (I1311268,I2507,I656182,I656409,);
nor I_38463 (I656417,I656409,I656276);
not I_38464 (I656434,I656417);
not I_38465 (I656451,I656409);
nor I_38466 (I656468,I656451,I656352);
DFFARX1 I_38467 (I656468,I2507,I656182,I656168,);
nand I_38468 (I656499,I1311265,I1311271);
and I_38469 (I656516,I656499,I1311286);
DFFARX1 I_38470 (I656516,I2507,I656182,I656542,);
nor I_38471 (I656550,I656542,I656409);
DFFARX1 I_38472 (I656550,I2507,I656182,I656150,);
nand I_38473 (I656581,I656542,I656451);
nand I_38474 (I656159,I656434,I656581);
not I_38475 (I656612,I656542);
nor I_38476 (I656629,I656612,I656352);
DFFARX1 I_38477 (I656629,I2507,I656182,I656171,);
nor I_38478 (I656660,I1311283,I1311271);
or I_38479 (I656162,I656409,I656660);
nor I_38480 (I656153,I656542,I656660);
or I_38481 (I656156,I656276,I656660);
DFFARX1 I_38482 (I656660,I2507,I656182,I656174,);
not I_38483 (I656760,I2514);
DFFARX1 I_38484 (I261281,I2507,I656760,I656786,);
not I_38485 (I656794,I656786);
nand I_38486 (I656811,I261284,I261260);
and I_38487 (I656828,I656811,I261257);
DFFARX1 I_38488 (I656828,I2507,I656760,I656854,);
not I_38489 (I656862,I261263);
DFFARX1 I_38490 (I261257,I2507,I656760,I656888,);
not I_38491 (I656896,I656888);
nor I_38492 (I656913,I656896,I656794);
and I_38493 (I656930,I656913,I261263);
nor I_38494 (I656947,I656896,I656862);
nor I_38495 (I656743,I656854,I656947);
DFFARX1 I_38496 (I261266,I2507,I656760,I656987,);
nor I_38497 (I656995,I656987,I656854);
not I_38498 (I657012,I656995);
not I_38499 (I657029,I656987);
nor I_38500 (I657046,I657029,I656930);
DFFARX1 I_38501 (I657046,I2507,I656760,I656746,);
nand I_38502 (I657077,I261269,I261278);
and I_38503 (I657094,I657077,I261275);
DFFARX1 I_38504 (I657094,I2507,I656760,I657120,);
nor I_38505 (I657128,I657120,I656987);
DFFARX1 I_38506 (I657128,I2507,I656760,I656728,);
nand I_38507 (I657159,I657120,I657029);
nand I_38508 (I656737,I657012,I657159);
not I_38509 (I657190,I657120);
nor I_38510 (I657207,I657190,I656930);
DFFARX1 I_38511 (I657207,I2507,I656760,I656749,);
nor I_38512 (I657238,I261272,I261278);
or I_38513 (I656740,I656987,I657238);
nor I_38514 (I656731,I657120,I657238);
or I_38515 (I656734,I656854,I657238);
DFFARX1 I_38516 (I657238,I2507,I656760,I656752,);
not I_38517 (I657338,I2514);
DFFARX1 I_38518 (I293428,I2507,I657338,I657364,);
not I_38519 (I657372,I657364);
nand I_38520 (I657389,I293431,I293407);
and I_38521 (I657406,I657389,I293404);
DFFARX1 I_38522 (I657406,I2507,I657338,I657432,);
not I_38523 (I657440,I293410);
DFFARX1 I_38524 (I293404,I2507,I657338,I657466,);
not I_38525 (I657474,I657466);
nor I_38526 (I657491,I657474,I657372);
and I_38527 (I657508,I657491,I293410);
nor I_38528 (I657525,I657474,I657440);
nor I_38529 (I657321,I657432,I657525);
DFFARX1 I_38530 (I293413,I2507,I657338,I657565,);
nor I_38531 (I657573,I657565,I657432);
not I_38532 (I657590,I657573);
not I_38533 (I657607,I657565);
nor I_38534 (I657624,I657607,I657508);
DFFARX1 I_38535 (I657624,I2507,I657338,I657324,);
nand I_38536 (I657655,I293416,I293425);
and I_38537 (I657672,I657655,I293422);
DFFARX1 I_38538 (I657672,I2507,I657338,I657698,);
nor I_38539 (I657706,I657698,I657565);
DFFARX1 I_38540 (I657706,I2507,I657338,I657306,);
nand I_38541 (I657737,I657698,I657607);
nand I_38542 (I657315,I657590,I657737);
not I_38543 (I657768,I657698);
nor I_38544 (I657785,I657768,I657508);
DFFARX1 I_38545 (I657785,I2507,I657338,I657327,);
nor I_38546 (I657816,I293419,I293425);
or I_38547 (I657318,I657565,I657816);
nor I_38548 (I657309,I657698,I657816);
or I_38549 (I657312,I657432,I657816);
DFFARX1 I_38550 (I657816,I2507,I657338,I657330,);
not I_38551 (I657916,I2514);
DFFARX1 I_38552 (I931523,I2507,I657916,I657942,);
not I_38553 (I657950,I657942);
nand I_38554 (I657967,I931499,I931514);
and I_38555 (I657984,I657967,I931526);
DFFARX1 I_38556 (I657984,I2507,I657916,I658010,);
not I_38557 (I658018,I931511);
DFFARX1 I_38558 (I931502,I2507,I657916,I658044,);
not I_38559 (I658052,I658044);
nor I_38560 (I658069,I658052,I657950);
and I_38561 (I658086,I658069,I931511);
nor I_38562 (I658103,I658052,I658018);
nor I_38563 (I657899,I658010,I658103);
DFFARX1 I_38564 (I931499,I2507,I657916,I658143,);
nor I_38565 (I658151,I658143,I658010);
not I_38566 (I658168,I658151);
not I_38567 (I658185,I658143);
nor I_38568 (I658202,I658185,I658086);
DFFARX1 I_38569 (I658202,I2507,I657916,I657902,);
nand I_38570 (I658233,I931517,I931508);
and I_38571 (I658250,I658233,I931520);
DFFARX1 I_38572 (I658250,I2507,I657916,I658276,);
nor I_38573 (I658284,I658276,I658143);
DFFARX1 I_38574 (I658284,I2507,I657916,I657884,);
nand I_38575 (I658315,I658276,I658185);
nand I_38576 (I657893,I658168,I658315);
not I_38577 (I658346,I658276);
nor I_38578 (I658363,I658346,I658086);
DFFARX1 I_38579 (I658363,I2507,I657916,I657905,);
nor I_38580 (I658394,I931505,I931508);
or I_38581 (I657896,I658143,I658394);
nor I_38582 (I657887,I658276,I658394);
or I_38583 (I657890,I658010,I658394);
DFFARX1 I_38584 (I658394,I2507,I657916,I657908,);
not I_38585 (I658494,I2514);
DFFARX1 I_38586 (I856544,I2507,I658494,I658520,);
not I_38587 (I658528,I658520);
nand I_38588 (I658545,I856532,I856550);
and I_38589 (I658562,I658545,I856547);
DFFARX1 I_38590 (I658562,I2507,I658494,I658588,);
not I_38591 (I658596,I856538);
DFFARX1 I_38592 (I856535,I2507,I658494,I658622,);
not I_38593 (I658630,I658622);
nor I_38594 (I658647,I658630,I658528);
and I_38595 (I658664,I658647,I856538);
nor I_38596 (I658681,I658630,I658596);
nor I_38597 (I658477,I658588,I658681);
DFFARX1 I_38598 (I856529,I2507,I658494,I658721,);
nor I_38599 (I658729,I658721,I658588);
not I_38600 (I658746,I658729);
not I_38601 (I658763,I658721);
nor I_38602 (I658780,I658763,I658664);
DFFARX1 I_38603 (I658780,I2507,I658494,I658480,);
nand I_38604 (I658811,I856529,I856532);
and I_38605 (I658828,I658811,I856535);
DFFARX1 I_38606 (I658828,I2507,I658494,I658854,);
nor I_38607 (I658862,I658854,I658721);
DFFARX1 I_38608 (I658862,I2507,I658494,I658462,);
nand I_38609 (I658893,I658854,I658763);
nand I_38610 (I658471,I658746,I658893);
not I_38611 (I658924,I658854);
nor I_38612 (I658941,I658924,I658664);
DFFARX1 I_38613 (I658941,I2507,I658494,I658483,);
nor I_38614 (I658972,I856541,I856532);
or I_38615 (I658474,I658721,I658972);
nor I_38616 (I658465,I658854,I658972);
or I_38617 (I658468,I658588,I658972);
DFFARX1 I_38618 (I658972,I2507,I658494,I658486,);
not I_38619 (I659072,I2514);
DFFARX1 I_38620 (I498849,I2507,I659072,I659098,);
not I_38621 (I659106,I659098);
nand I_38622 (I659123,I498864,I498849);
and I_38623 (I659140,I659123,I498852);
DFFARX1 I_38624 (I659140,I2507,I659072,I659166,);
not I_38625 (I659174,I498852);
DFFARX1 I_38626 (I498861,I2507,I659072,I659200,);
not I_38627 (I659208,I659200);
nor I_38628 (I659225,I659208,I659106);
and I_38629 (I659242,I659225,I498852);
nor I_38630 (I659259,I659208,I659174);
nor I_38631 (I659055,I659166,I659259);
DFFARX1 I_38632 (I498855,I2507,I659072,I659299,);
nor I_38633 (I659307,I659299,I659166);
not I_38634 (I659324,I659307);
not I_38635 (I659341,I659299);
nor I_38636 (I659358,I659341,I659242);
DFFARX1 I_38637 (I659358,I2507,I659072,I659058,);
nand I_38638 (I659389,I498858,I498867);
and I_38639 (I659406,I659389,I498873);
DFFARX1 I_38640 (I659406,I2507,I659072,I659432,);
nor I_38641 (I659440,I659432,I659299);
DFFARX1 I_38642 (I659440,I2507,I659072,I659040,);
nand I_38643 (I659471,I659432,I659341);
nand I_38644 (I659049,I659324,I659471);
not I_38645 (I659502,I659432);
nor I_38646 (I659519,I659502,I659242);
DFFARX1 I_38647 (I659519,I2507,I659072,I659061,);
nor I_38648 (I659550,I498870,I498867);
or I_38649 (I659052,I659299,I659550);
nor I_38650 (I659043,I659432,I659550);
or I_38651 (I659046,I659166,I659550);
DFFARX1 I_38652 (I659550,I2507,I659072,I659064,);
not I_38653 (I659650,I2514);
DFFARX1 I_38654 (I325048,I2507,I659650,I659676,);
not I_38655 (I659684,I659676);
nand I_38656 (I659701,I325051,I325027);
and I_38657 (I659718,I659701,I325024);
DFFARX1 I_38658 (I659718,I2507,I659650,I659744,);
not I_38659 (I659752,I325030);
DFFARX1 I_38660 (I325024,I2507,I659650,I659778,);
not I_38661 (I659786,I659778);
nor I_38662 (I659803,I659786,I659684);
and I_38663 (I659820,I659803,I325030);
nor I_38664 (I659837,I659786,I659752);
nor I_38665 (I659633,I659744,I659837);
DFFARX1 I_38666 (I325033,I2507,I659650,I659877,);
nor I_38667 (I659885,I659877,I659744);
not I_38668 (I659902,I659885);
not I_38669 (I659919,I659877);
nor I_38670 (I659936,I659919,I659820);
DFFARX1 I_38671 (I659936,I2507,I659650,I659636,);
nand I_38672 (I659967,I325036,I325045);
and I_38673 (I659984,I659967,I325042);
DFFARX1 I_38674 (I659984,I2507,I659650,I660010,);
nor I_38675 (I660018,I660010,I659877);
DFFARX1 I_38676 (I660018,I2507,I659650,I659618,);
nand I_38677 (I660049,I660010,I659919);
nand I_38678 (I659627,I659902,I660049);
not I_38679 (I660080,I660010);
nor I_38680 (I660097,I660080,I659820);
DFFARX1 I_38681 (I660097,I2507,I659650,I659639,);
nor I_38682 (I660128,I325039,I325045);
or I_38683 (I659630,I659877,I660128);
nor I_38684 (I659621,I660010,I660128);
or I_38685 (I659624,I659744,I660128);
DFFARX1 I_38686 (I660128,I2507,I659650,I659642,);
not I_38687 (I660228,I2514);
DFFARX1 I_38688 (I994831,I2507,I660228,I660254,);
not I_38689 (I660262,I660254);
nand I_38690 (I660279,I994807,I994822);
and I_38691 (I660296,I660279,I994834);
DFFARX1 I_38692 (I660296,I2507,I660228,I660322,);
not I_38693 (I660330,I994819);
DFFARX1 I_38694 (I994810,I2507,I660228,I660356,);
not I_38695 (I660364,I660356);
nor I_38696 (I660381,I660364,I660262);
and I_38697 (I660398,I660381,I994819);
nor I_38698 (I660415,I660364,I660330);
nor I_38699 (I660211,I660322,I660415);
DFFARX1 I_38700 (I994807,I2507,I660228,I660455,);
nor I_38701 (I660463,I660455,I660322);
not I_38702 (I660480,I660463);
not I_38703 (I660497,I660455);
nor I_38704 (I660514,I660497,I660398);
DFFARX1 I_38705 (I660514,I2507,I660228,I660214,);
nand I_38706 (I660545,I994825,I994816);
and I_38707 (I660562,I660545,I994828);
DFFARX1 I_38708 (I660562,I2507,I660228,I660588,);
nor I_38709 (I660596,I660588,I660455);
DFFARX1 I_38710 (I660596,I2507,I660228,I660196,);
nand I_38711 (I660627,I660588,I660497);
nand I_38712 (I660205,I660480,I660627);
not I_38713 (I660658,I660588);
nor I_38714 (I660675,I660658,I660398);
DFFARX1 I_38715 (I660675,I2507,I660228,I660217,);
nor I_38716 (I660706,I994813,I994816);
or I_38717 (I660208,I660455,I660706);
nor I_38718 (I660199,I660588,I660706);
or I_38719 (I660202,I660322,I660706);
DFFARX1 I_38720 (I660706,I2507,I660228,I660220,);
not I_38721 (I660806,I2514);
DFFARX1 I_38722 (I537524,I2507,I660806,I660832,);
not I_38723 (I660840,I660832);
nand I_38724 (I660857,I537539,I537524);
and I_38725 (I660874,I660857,I537527);
DFFARX1 I_38726 (I660874,I2507,I660806,I660900,);
not I_38727 (I660908,I537527);
DFFARX1 I_38728 (I537536,I2507,I660806,I660934,);
not I_38729 (I660942,I660934);
nor I_38730 (I660959,I660942,I660840);
and I_38731 (I660976,I660959,I537527);
nor I_38732 (I660993,I660942,I660908);
nor I_38733 (I660789,I660900,I660993);
DFFARX1 I_38734 (I537530,I2507,I660806,I661033,);
nor I_38735 (I661041,I661033,I660900);
not I_38736 (I661058,I661041);
not I_38737 (I661075,I661033);
nor I_38738 (I661092,I661075,I660976);
DFFARX1 I_38739 (I661092,I2507,I660806,I660792,);
nand I_38740 (I661123,I537533,I537542);
and I_38741 (I661140,I661123,I537548);
DFFARX1 I_38742 (I661140,I2507,I660806,I661166,);
nor I_38743 (I661174,I661166,I661033);
DFFARX1 I_38744 (I661174,I2507,I660806,I660774,);
nand I_38745 (I661205,I661166,I661075);
nand I_38746 (I660783,I661058,I661205);
not I_38747 (I661236,I661166);
nor I_38748 (I661253,I661236,I660976);
DFFARX1 I_38749 (I661253,I2507,I660806,I660795,);
nor I_38750 (I661284,I537545,I537542);
or I_38751 (I660786,I661033,I661284);
nor I_38752 (I660777,I661166,I661284);
or I_38753 (I660780,I660900,I661284);
DFFARX1 I_38754 (I661284,I2507,I660806,I660798,);
not I_38755 (I661384,I2514);
DFFARX1 I_38756 (I495279,I2507,I661384,I661410,);
not I_38757 (I661418,I661410);
nand I_38758 (I661435,I495294,I495279);
and I_38759 (I661452,I661435,I495282);
DFFARX1 I_38760 (I661452,I2507,I661384,I661478,);
not I_38761 (I661486,I495282);
DFFARX1 I_38762 (I495291,I2507,I661384,I661512,);
not I_38763 (I661520,I661512);
nor I_38764 (I661537,I661520,I661418);
and I_38765 (I661554,I661537,I495282);
nor I_38766 (I661571,I661520,I661486);
nor I_38767 (I661367,I661478,I661571);
DFFARX1 I_38768 (I495285,I2507,I661384,I661611,);
nor I_38769 (I661619,I661611,I661478);
not I_38770 (I661636,I661619);
not I_38771 (I661653,I661611);
nor I_38772 (I661670,I661653,I661554);
DFFARX1 I_38773 (I661670,I2507,I661384,I661370,);
nand I_38774 (I661701,I495288,I495297);
and I_38775 (I661718,I661701,I495303);
DFFARX1 I_38776 (I661718,I2507,I661384,I661744,);
nor I_38777 (I661752,I661744,I661611);
DFFARX1 I_38778 (I661752,I2507,I661384,I661352,);
nand I_38779 (I661783,I661744,I661653);
nand I_38780 (I661361,I661636,I661783);
not I_38781 (I661814,I661744);
nor I_38782 (I661831,I661814,I661554);
DFFARX1 I_38783 (I661831,I2507,I661384,I661373,);
nor I_38784 (I661862,I495300,I495297);
or I_38785 (I661364,I661611,I661862);
nor I_38786 (I661355,I661744,I661862);
or I_38787 (I661358,I661478,I661862);
DFFARX1 I_38788 (I661862,I2507,I661384,I661376,);
not I_38789 (I661962,I2514);
DFFARX1 I_38790 (I834937,I2507,I661962,I661988,);
not I_38791 (I661996,I661988);
nand I_38792 (I662013,I834925,I834943);
and I_38793 (I662030,I662013,I834940);
DFFARX1 I_38794 (I662030,I2507,I661962,I662056,);
not I_38795 (I662064,I834931);
DFFARX1 I_38796 (I834928,I2507,I661962,I662090,);
not I_38797 (I662098,I662090);
nor I_38798 (I662115,I662098,I661996);
and I_38799 (I662132,I662115,I834931);
nor I_38800 (I662149,I662098,I662064);
nor I_38801 (I661945,I662056,I662149);
DFFARX1 I_38802 (I834922,I2507,I661962,I662189,);
nor I_38803 (I662197,I662189,I662056);
not I_38804 (I662214,I662197);
not I_38805 (I662231,I662189);
nor I_38806 (I662248,I662231,I662132);
DFFARX1 I_38807 (I662248,I2507,I661962,I661948,);
nand I_38808 (I662279,I834922,I834925);
and I_38809 (I662296,I662279,I834928);
DFFARX1 I_38810 (I662296,I2507,I661962,I662322,);
nor I_38811 (I662330,I662322,I662189);
DFFARX1 I_38812 (I662330,I2507,I661962,I661930,);
nand I_38813 (I662361,I662322,I662231);
nand I_38814 (I661939,I662214,I662361);
not I_38815 (I662392,I662322);
nor I_38816 (I662409,I662392,I662132);
DFFARX1 I_38817 (I662409,I2507,I661962,I661951,);
nor I_38818 (I662440,I834934,I834925);
or I_38819 (I661942,I662189,I662440);
nor I_38820 (I661933,I662322,I662440);
or I_38821 (I661936,I662056,I662440);
DFFARX1 I_38822 (I662440,I2507,I661962,I661954,);
not I_38823 (I662540,I2514);
DFFARX1 I_38824 (I1173410,I2507,I662540,I662566,);
not I_38825 (I662574,I662566);
nand I_38826 (I662591,I1173392,I1173404);
and I_38827 (I662608,I662591,I1173407);
DFFARX1 I_38828 (I662608,I2507,I662540,I662634,);
not I_38829 (I662642,I1173401);
DFFARX1 I_38830 (I1173398,I2507,I662540,I662668,);
not I_38831 (I662676,I662668);
nor I_38832 (I662693,I662676,I662574);
and I_38833 (I662710,I662693,I1173401);
nor I_38834 (I662727,I662676,I662642);
nor I_38835 (I662523,I662634,I662727);
DFFARX1 I_38836 (I1173416,I2507,I662540,I662767,);
nor I_38837 (I662775,I662767,I662634);
not I_38838 (I662792,I662775);
not I_38839 (I662809,I662767);
nor I_38840 (I662826,I662809,I662710);
DFFARX1 I_38841 (I662826,I2507,I662540,I662526,);
nand I_38842 (I662857,I1173395,I1173395);
and I_38843 (I662874,I662857,I1173392);
DFFARX1 I_38844 (I662874,I2507,I662540,I662900,);
nor I_38845 (I662908,I662900,I662767);
DFFARX1 I_38846 (I662908,I2507,I662540,I662508,);
nand I_38847 (I662939,I662900,I662809);
nand I_38848 (I662517,I662792,I662939);
not I_38849 (I662970,I662900);
nor I_38850 (I662987,I662970,I662710);
DFFARX1 I_38851 (I662987,I2507,I662540,I662529,);
nor I_38852 (I663018,I1173413,I1173395);
or I_38853 (I662520,I662767,I663018);
nor I_38854 (I662511,I662900,I663018);
or I_38855 (I662514,I662634,I663018);
DFFARX1 I_38856 (I663018,I2507,I662540,I662532,);
not I_38857 (I663118,I2514);
DFFARX1 I_38858 (I790669,I2507,I663118,I663144,);
not I_38859 (I663152,I663144);
nand I_38860 (I663169,I790657,I790675);
and I_38861 (I663186,I663169,I790672);
DFFARX1 I_38862 (I663186,I2507,I663118,I663212,);
not I_38863 (I663220,I790663);
DFFARX1 I_38864 (I790660,I2507,I663118,I663246,);
not I_38865 (I663254,I663246);
nor I_38866 (I663271,I663254,I663152);
and I_38867 (I663288,I663271,I790663);
nor I_38868 (I663305,I663254,I663220);
nor I_38869 (I663101,I663212,I663305);
DFFARX1 I_38870 (I790654,I2507,I663118,I663345,);
nor I_38871 (I663353,I663345,I663212);
not I_38872 (I663370,I663353);
not I_38873 (I663387,I663345);
nor I_38874 (I663404,I663387,I663288);
DFFARX1 I_38875 (I663404,I2507,I663118,I663104,);
nand I_38876 (I663435,I790654,I790657);
and I_38877 (I663452,I663435,I790660);
DFFARX1 I_38878 (I663452,I2507,I663118,I663478,);
nor I_38879 (I663486,I663478,I663345);
DFFARX1 I_38880 (I663486,I2507,I663118,I663086,);
nand I_38881 (I663517,I663478,I663387);
nand I_38882 (I663095,I663370,I663517);
not I_38883 (I663548,I663478);
nor I_38884 (I663565,I663548,I663288);
DFFARX1 I_38885 (I663565,I2507,I663118,I663107,);
nor I_38886 (I663596,I790666,I790657);
or I_38887 (I663098,I663345,I663596);
nor I_38888 (I663089,I663478,I663596);
or I_38889 (I663092,I663212,I663596);
DFFARX1 I_38890 (I663596,I2507,I663118,I663110,);
not I_38891 (I663696,I2514);
DFFARX1 I_38892 (I1242242,I2507,I663696,I663722,);
not I_38893 (I663730,I663722);
nand I_38894 (I663747,I1242245,I1242254);
and I_38895 (I663764,I663747,I1242257);
DFFARX1 I_38896 (I663764,I2507,I663696,I663790,);
not I_38897 (I663798,I1242266);
DFFARX1 I_38898 (I1242248,I2507,I663696,I663824,);
not I_38899 (I663832,I663824);
nor I_38900 (I663849,I663832,I663730);
and I_38901 (I663866,I663849,I1242266);
nor I_38902 (I663883,I663832,I663798);
nor I_38903 (I663679,I663790,I663883);
DFFARX1 I_38904 (I1242245,I2507,I663696,I663923,);
nor I_38905 (I663931,I663923,I663790);
not I_38906 (I663948,I663931);
not I_38907 (I663965,I663923);
nor I_38908 (I663982,I663965,I663866);
DFFARX1 I_38909 (I663982,I2507,I663696,I663682,);
nand I_38910 (I664013,I1242263,I1242242);
and I_38911 (I664030,I664013,I1242260);
DFFARX1 I_38912 (I664030,I2507,I663696,I664056,);
nor I_38913 (I664064,I664056,I663923);
DFFARX1 I_38914 (I664064,I2507,I663696,I663664,);
nand I_38915 (I664095,I664056,I663965);
nand I_38916 (I663673,I663948,I664095);
not I_38917 (I664126,I664056);
nor I_38918 (I664143,I664126,I663866);
DFFARX1 I_38919 (I664143,I2507,I663696,I663685,);
nor I_38920 (I664174,I1242251,I1242242);
or I_38921 (I663676,I663923,I664174);
nor I_38922 (I663667,I664056,I664174);
or I_38923 (I663670,I663790,I664174);
DFFARX1 I_38924 (I664174,I2507,I663696,I663688,);
not I_38925 (I664274,I2514);
DFFARX1 I_38926 (I1202888,I2507,I664274,I664300,);
not I_38927 (I664308,I664300);
nand I_38928 (I664325,I1202870,I1202882);
and I_38929 (I664342,I664325,I1202885);
DFFARX1 I_38930 (I664342,I2507,I664274,I664368,);
not I_38931 (I664376,I1202879);
DFFARX1 I_38932 (I1202876,I2507,I664274,I664402,);
not I_38933 (I664410,I664402);
nor I_38934 (I664427,I664410,I664308);
and I_38935 (I664444,I664427,I1202879);
nor I_38936 (I664461,I664410,I664376);
nor I_38937 (I664257,I664368,I664461);
DFFARX1 I_38938 (I1202894,I2507,I664274,I664501,);
nor I_38939 (I664509,I664501,I664368);
not I_38940 (I664526,I664509);
not I_38941 (I664543,I664501);
nor I_38942 (I664560,I664543,I664444);
DFFARX1 I_38943 (I664560,I2507,I664274,I664260,);
nand I_38944 (I664591,I1202873,I1202873);
and I_38945 (I664608,I664591,I1202870);
DFFARX1 I_38946 (I664608,I2507,I664274,I664634,);
nor I_38947 (I664642,I664634,I664501);
DFFARX1 I_38948 (I664642,I2507,I664274,I664242,);
nand I_38949 (I664673,I664634,I664543);
nand I_38950 (I664251,I664526,I664673);
not I_38951 (I664704,I664634);
nor I_38952 (I664721,I664704,I664444);
DFFARX1 I_38953 (I664721,I2507,I664274,I664263,);
nor I_38954 (I664752,I1202891,I1202873);
or I_38955 (I664254,I664501,I664752);
nor I_38956 (I664245,I664634,I664752);
or I_38957 (I664248,I664368,I664752);
DFFARX1 I_38958 (I664752,I2507,I664274,I664266,);
not I_38959 (I664852,I2514);
DFFARX1 I_38960 (I340331,I2507,I664852,I664878,);
not I_38961 (I664886,I664878);
nand I_38962 (I664903,I340334,I340310);
and I_38963 (I664920,I664903,I340307);
DFFARX1 I_38964 (I664920,I2507,I664852,I664946,);
not I_38965 (I664954,I340313);
DFFARX1 I_38966 (I340307,I2507,I664852,I664980,);
not I_38967 (I664988,I664980);
nor I_38968 (I665005,I664988,I664886);
and I_38969 (I665022,I665005,I340313);
nor I_38970 (I665039,I664988,I664954);
nor I_38971 (I664835,I664946,I665039);
DFFARX1 I_38972 (I340316,I2507,I664852,I665079,);
nor I_38973 (I665087,I665079,I664946);
not I_38974 (I665104,I665087);
not I_38975 (I665121,I665079);
nor I_38976 (I665138,I665121,I665022);
DFFARX1 I_38977 (I665138,I2507,I664852,I664838,);
nand I_38978 (I665169,I340319,I340328);
and I_38979 (I665186,I665169,I340325);
DFFARX1 I_38980 (I665186,I2507,I664852,I665212,);
nor I_38981 (I665220,I665212,I665079);
DFFARX1 I_38982 (I665220,I2507,I664852,I664820,);
nand I_38983 (I665251,I665212,I665121);
nand I_38984 (I664829,I665104,I665251);
not I_38985 (I665282,I665212);
nor I_38986 (I665299,I665282,I665022);
DFFARX1 I_38987 (I665299,I2507,I664852,I664841,);
nor I_38988 (I665330,I340322,I340328);
or I_38989 (I664832,I665079,I665330);
nor I_38990 (I664823,I665212,I665330);
or I_38991 (I664826,I664946,I665330);
DFFARX1 I_38992 (I665330,I2507,I664852,I664844,);
not I_38993 (I665430,I2514);
DFFARX1 I_38994 (I1053905,I2507,I665430,I665456,);
not I_38995 (I665464,I665456);
nand I_38996 (I665481,I1053902,I1053920);
and I_38997 (I665498,I665481,I1053917);
DFFARX1 I_38998 (I665498,I2507,I665430,I665524,);
not I_38999 (I665532,I1053899);
DFFARX1 I_39000 (I1053902,I2507,I665430,I665558,);
not I_39001 (I665566,I665558);
nor I_39002 (I665583,I665566,I665464);
and I_39003 (I665600,I665583,I1053899);
nor I_39004 (I665617,I665566,I665532);
nor I_39005 (I665413,I665524,I665617);
DFFARX1 I_39006 (I1053911,I2507,I665430,I665657,);
nor I_39007 (I665665,I665657,I665524);
not I_39008 (I665682,I665665);
not I_39009 (I665699,I665657);
nor I_39010 (I665716,I665699,I665600);
DFFARX1 I_39011 (I665716,I2507,I665430,I665416,);
nand I_39012 (I665747,I1053914,I1053899);
and I_39013 (I665764,I665747,I1053905);
DFFARX1 I_39014 (I665764,I2507,I665430,I665790,);
nor I_39015 (I665798,I665790,I665657);
DFFARX1 I_39016 (I665798,I2507,I665430,I665398,);
nand I_39017 (I665829,I665790,I665699);
nand I_39018 (I665407,I665682,I665829);
not I_39019 (I665860,I665790);
nor I_39020 (I665877,I665860,I665600);
DFFARX1 I_39021 (I665877,I2507,I665430,I665419,);
nor I_39022 (I665908,I1053908,I1053899);
or I_39023 (I665410,I665657,I665908);
nor I_39024 (I665401,I665790,I665908);
or I_39025 (I665404,I665524,I665908);
DFFARX1 I_39026 (I665908,I2507,I665430,I665422,);
not I_39027 (I666008,I2514);
DFFARX1 I_39028 (I1289434,I2507,I666008,I666034,);
not I_39029 (I666042,I666034);
nand I_39030 (I666059,I1289458,I1289440);
and I_39031 (I666076,I666059,I1289446);
DFFARX1 I_39032 (I666076,I2507,I666008,I666102,);
not I_39033 (I666110,I1289452);
DFFARX1 I_39034 (I1289437,I2507,I666008,I666136,);
not I_39035 (I666144,I666136);
nor I_39036 (I666161,I666144,I666042);
and I_39037 (I666178,I666161,I1289452);
nor I_39038 (I666195,I666144,I666110);
nor I_39039 (I665991,I666102,I666195);
DFFARX1 I_39040 (I1289449,I2507,I666008,I666235,);
nor I_39041 (I666243,I666235,I666102);
not I_39042 (I666260,I666243);
not I_39043 (I666277,I666235);
nor I_39044 (I666294,I666277,I666178);
DFFARX1 I_39045 (I666294,I2507,I666008,I665994,);
nand I_39046 (I666325,I1289455,I1289443);
and I_39047 (I666342,I666325,I1289437);
DFFARX1 I_39048 (I666342,I2507,I666008,I666368,);
nor I_39049 (I666376,I666368,I666235);
DFFARX1 I_39050 (I666376,I2507,I666008,I665976,);
nand I_39051 (I666407,I666368,I666277);
nand I_39052 (I665985,I666260,I666407);
not I_39053 (I666438,I666368);
nor I_39054 (I666455,I666438,I666178);
DFFARX1 I_39055 (I666455,I2507,I666008,I665997,);
nor I_39056 (I666486,I1289434,I1289443);
or I_39057 (I665988,I666235,I666486);
nor I_39058 (I665979,I666368,I666486);
or I_39059 (I665982,I666102,I666486);
DFFARX1 I_39060 (I666486,I2507,I666008,I666000,);
not I_39061 (I666586,I2514);
DFFARX1 I_39062 (I463192,I2507,I666586,I666612,);
not I_39063 (I666620,I666612);
nand I_39064 (I666637,I463183,I463201);
and I_39065 (I666654,I666637,I463204);
DFFARX1 I_39066 (I666654,I2507,I666586,I666680,);
not I_39067 (I666688,I463198);
DFFARX1 I_39068 (I463186,I2507,I666586,I666714,);
not I_39069 (I666722,I666714);
nor I_39070 (I666739,I666722,I666620);
and I_39071 (I666756,I666739,I463198);
nor I_39072 (I666773,I666722,I666688);
nor I_39073 (I666569,I666680,I666773);
DFFARX1 I_39074 (I463195,I2507,I666586,I666813,);
nor I_39075 (I666821,I666813,I666680);
not I_39076 (I666838,I666821);
not I_39077 (I666855,I666813);
nor I_39078 (I666872,I666855,I666756);
DFFARX1 I_39079 (I666872,I2507,I666586,I666572,);
nand I_39080 (I666903,I463210,I463207);
and I_39081 (I666920,I666903,I463189);
DFFARX1 I_39082 (I666920,I2507,I666586,I666946,);
nor I_39083 (I666954,I666946,I666813);
DFFARX1 I_39084 (I666954,I2507,I666586,I666554,);
nand I_39085 (I666985,I666946,I666855);
nand I_39086 (I666563,I666838,I666985);
not I_39087 (I667016,I666946);
nor I_39088 (I667033,I667016,I666756);
DFFARX1 I_39089 (I667033,I2507,I666586,I666575,);
nor I_39090 (I667064,I463183,I463207);
or I_39091 (I666566,I666813,I667064);
nor I_39092 (I666557,I666946,I667064);
or I_39093 (I666560,I666680,I667064);
DFFARX1 I_39094 (I667064,I2507,I666586,I666578,);
not I_39095 (I667164,I2514);
DFFARX1 I_39096 (I40116,I2507,I667164,I667190,);
not I_39097 (I667198,I667190);
nand I_39098 (I667215,I40113,I40104);
and I_39099 (I667232,I667215,I40104);
DFFARX1 I_39100 (I667232,I2507,I667164,I667258,);
not I_39101 (I667266,I40107);
DFFARX1 I_39102 (I40122,I2507,I667164,I667292,);
not I_39103 (I667300,I667292);
nor I_39104 (I667317,I667300,I667198);
and I_39105 (I667334,I667317,I40107);
nor I_39106 (I667351,I667300,I667266);
nor I_39107 (I667147,I667258,I667351);
DFFARX1 I_39108 (I40107,I2507,I667164,I667391,);
nor I_39109 (I667399,I667391,I667258);
not I_39110 (I667416,I667399);
not I_39111 (I667433,I667391);
nor I_39112 (I667450,I667433,I667334);
DFFARX1 I_39113 (I667450,I2507,I667164,I667150,);
nand I_39114 (I667481,I40125,I40110);
and I_39115 (I667498,I667481,I40128);
DFFARX1 I_39116 (I667498,I2507,I667164,I667524,);
nor I_39117 (I667532,I667524,I667391);
DFFARX1 I_39118 (I667532,I2507,I667164,I667132,);
nand I_39119 (I667563,I667524,I667433);
nand I_39120 (I667141,I667416,I667563);
not I_39121 (I667594,I667524);
nor I_39122 (I667611,I667594,I667334);
DFFARX1 I_39123 (I667611,I2507,I667164,I667153,);
nor I_39124 (I667642,I40119,I40110);
or I_39125 (I667144,I667391,I667642);
nor I_39126 (I667135,I667524,I667642);
or I_39127 (I667138,I667258,I667642);
DFFARX1 I_39128 (I667642,I2507,I667164,I667156,);
not I_39129 (I667742,I2514);
DFFARX1 I_39130 (I1162428,I2507,I667742,I667768,);
not I_39131 (I667776,I667768);
nand I_39132 (I667793,I1162410,I1162422);
and I_39133 (I667810,I667793,I1162425);
DFFARX1 I_39134 (I667810,I2507,I667742,I667836,);
not I_39135 (I667844,I1162419);
DFFARX1 I_39136 (I1162416,I2507,I667742,I667870,);
not I_39137 (I667878,I667870);
nor I_39138 (I667895,I667878,I667776);
and I_39139 (I667912,I667895,I1162419);
nor I_39140 (I667929,I667878,I667844);
nor I_39141 (I667725,I667836,I667929);
DFFARX1 I_39142 (I1162434,I2507,I667742,I667969,);
nor I_39143 (I667977,I667969,I667836);
not I_39144 (I667994,I667977);
not I_39145 (I668011,I667969);
nor I_39146 (I668028,I668011,I667912);
DFFARX1 I_39147 (I668028,I2507,I667742,I667728,);
nand I_39148 (I668059,I1162413,I1162413);
and I_39149 (I668076,I668059,I1162410);
DFFARX1 I_39150 (I668076,I2507,I667742,I668102,);
nor I_39151 (I668110,I668102,I667969);
DFFARX1 I_39152 (I668110,I2507,I667742,I667710,);
nand I_39153 (I668141,I668102,I668011);
nand I_39154 (I667719,I667994,I668141);
not I_39155 (I668172,I668102);
nor I_39156 (I668189,I668172,I667912);
DFFARX1 I_39157 (I668189,I2507,I667742,I667731,);
nor I_39158 (I668220,I1162431,I1162413);
or I_39159 (I667722,I667969,I668220);
nor I_39160 (I667713,I668102,I668220);
or I_39161 (I667716,I667836,I668220);
DFFARX1 I_39162 (I668220,I2507,I667742,I667734,);
not I_39163 (I668320,I2514);
DFFARX1 I_39164 (I929585,I2507,I668320,I668346,);
not I_39165 (I668354,I668346);
nand I_39166 (I668371,I929561,I929576);
and I_39167 (I668388,I668371,I929588);
DFFARX1 I_39168 (I668388,I2507,I668320,I668414,);
not I_39169 (I668422,I929573);
DFFARX1 I_39170 (I929564,I2507,I668320,I668448,);
not I_39171 (I668456,I668448);
nor I_39172 (I668473,I668456,I668354);
and I_39173 (I668490,I668473,I929573);
nor I_39174 (I668507,I668456,I668422);
nor I_39175 (I668303,I668414,I668507);
DFFARX1 I_39176 (I929561,I2507,I668320,I668547,);
nor I_39177 (I668555,I668547,I668414);
not I_39178 (I668572,I668555);
not I_39179 (I668589,I668547);
nor I_39180 (I668606,I668589,I668490);
DFFARX1 I_39181 (I668606,I2507,I668320,I668306,);
nand I_39182 (I668637,I929579,I929570);
and I_39183 (I668654,I668637,I929582);
DFFARX1 I_39184 (I668654,I2507,I668320,I668680,);
nor I_39185 (I668688,I668680,I668547);
DFFARX1 I_39186 (I668688,I2507,I668320,I668288,);
nand I_39187 (I668719,I668680,I668589);
nand I_39188 (I668297,I668572,I668719);
not I_39189 (I668750,I668680);
nor I_39190 (I668767,I668750,I668490);
DFFARX1 I_39191 (I668767,I2507,I668320,I668309,);
nor I_39192 (I668798,I929567,I929570);
or I_39193 (I668300,I668547,I668798);
nor I_39194 (I668291,I668680,I668798);
or I_39195 (I668294,I668414,I668798);
DFFARX1 I_39196 (I668798,I2507,I668320,I668312,);
not I_39197 (I668898,I2514);
DFFARX1 I_39198 (I605286,I2507,I668898,I668924,);
not I_39199 (I668932,I668924);
nand I_39200 (I668949,I605295,I605304);
and I_39201 (I668966,I668949,I605310);
DFFARX1 I_39202 (I668966,I2507,I668898,I668992,);
not I_39203 (I669000,I605307);
DFFARX1 I_39204 (I605292,I2507,I668898,I669026,);
not I_39205 (I669034,I669026);
nor I_39206 (I669051,I669034,I668932);
and I_39207 (I669068,I669051,I605307);
nor I_39208 (I669085,I669034,I669000);
nor I_39209 (I668881,I668992,I669085);
DFFARX1 I_39210 (I605301,I2507,I668898,I669125,);
nor I_39211 (I669133,I669125,I668992);
not I_39212 (I669150,I669133);
not I_39213 (I669167,I669125);
nor I_39214 (I669184,I669167,I669068);
DFFARX1 I_39215 (I669184,I2507,I668898,I668884,);
nand I_39216 (I669215,I605298,I605289);
and I_39217 (I669232,I669215,I605286);
DFFARX1 I_39218 (I669232,I2507,I668898,I669258,);
nor I_39219 (I669266,I669258,I669125);
DFFARX1 I_39220 (I669266,I2507,I668898,I668866,);
nand I_39221 (I669297,I669258,I669167);
nand I_39222 (I668875,I669150,I669297);
not I_39223 (I669328,I669258);
nor I_39224 (I669345,I669328,I669068);
DFFARX1 I_39225 (I669345,I2507,I668898,I668887,);
nor I_39226 (I669376,I605289,I605289);
or I_39227 (I668878,I669125,I669376);
nor I_39228 (I668869,I669258,I669376);
or I_39229 (I668872,I668992,I669376);
DFFARX1 I_39230 (I669376,I2507,I668898,I668890,);
not I_39231 (I669476,I2514);
DFFARX1 I_39232 (I824924,I2507,I669476,I669502,);
not I_39233 (I669510,I669502);
nand I_39234 (I669527,I824912,I824930);
and I_39235 (I669544,I669527,I824927);
DFFARX1 I_39236 (I669544,I2507,I669476,I669570,);
not I_39237 (I669578,I824918);
DFFARX1 I_39238 (I824915,I2507,I669476,I669604,);
not I_39239 (I669612,I669604);
nor I_39240 (I669629,I669612,I669510);
and I_39241 (I669646,I669629,I824918);
nor I_39242 (I669663,I669612,I669578);
nor I_39243 (I669459,I669570,I669663);
DFFARX1 I_39244 (I824909,I2507,I669476,I669703,);
nor I_39245 (I669711,I669703,I669570);
not I_39246 (I669728,I669711);
not I_39247 (I669745,I669703);
nor I_39248 (I669762,I669745,I669646);
DFFARX1 I_39249 (I669762,I2507,I669476,I669462,);
nand I_39250 (I669793,I824909,I824912);
and I_39251 (I669810,I669793,I824915);
DFFARX1 I_39252 (I669810,I2507,I669476,I669836,);
nor I_39253 (I669844,I669836,I669703);
DFFARX1 I_39254 (I669844,I2507,I669476,I669444,);
nand I_39255 (I669875,I669836,I669745);
nand I_39256 (I669453,I669728,I669875);
not I_39257 (I669906,I669836);
nor I_39258 (I669923,I669906,I669646);
DFFARX1 I_39259 (I669923,I2507,I669476,I669465,);
nor I_39260 (I669954,I824921,I824912);
or I_39261 (I669456,I669703,I669954);
nor I_39262 (I669447,I669836,I669954);
or I_39263 (I669450,I669570,I669954);
DFFARX1 I_39264 (I669954,I2507,I669476,I669468,);
not I_39265 (I670054,I2514);
DFFARX1 I_39266 (I45913,I2507,I670054,I670080,);
not I_39267 (I670088,I670080);
nand I_39268 (I670105,I45910,I45901);
and I_39269 (I670122,I670105,I45901);
DFFARX1 I_39270 (I670122,I2507,I670054,I670148,);
not I_39271 (I670156,I45904);
DFFARX1 I_39272 (I45919,I2507,I670054,I670182,);
not I_39273 (I670190,I670182);
nor I_39274 (I670207,I670190,I670088);
and I_39275 (I670224,I670207,I45904);
nor I_39276 (I670241,I670190,I670156);
nor I_39277 (I670037,I670148,I670241);
DFFARX1 I_39278 (I45904,I2507,I670054,I670281,);
nor I_39279 (I670289,I670281,I670148);
not I_39280 (I670306,I670289);
not I_39281 (I670323,I670281);
nor I_39282 (I670340,I670323,I670224);
DFFARX1 I_39283 (I670340,I2507,I670054,I670040,);
nand I_39284 (I670371,I45922,I45907);
and I_39285 (I670388,I670371,I45925);
DFFARX1 I_39286 (I670388,I2507,I670054,I670414,);
nor I_39287 (I670422,I670414,I670281);
DFFARX1 I_39288 (I670422,I2507,I670054,I670022,);
nand I_39289 (I670453,I670414,I670323);
nand I_39290 (I670031,I670306,I670453);
not I_39291 (I670484,I670414);
nor I_39292 (I670501,I670484,I670224);
DFFARX1 I_39293 (I670501,I2507,I670054,I670043,);
nor I_39294 (I670532,I45916,I45907);
or I_39295 (I670034,I670281,I670532);
nor I_39296 (I670025,I670414,I670532);
or I_39297 (I670028,I670148,I670532);
DFFARX1 I_39298 (I670532,I2507,I670054,I670046,);
not I_39299 (I670632,I2514);
DFFARX1 I_39300 (I579276,I2507,I670632,I670658,);
not I_39301 (I670666,I670658);
nand I_39302 (I670683,I579285,I579294);
and I_39303 (I670700,I670683,I579300);
DFFARX1 I_39304 (I670700,I2507,I670632,I670726,);
not I_39305 (I670734,I579297);
DFFARX1 I_39306 (I579282,I2507,I670632,I670760,);
not I_39307 (I670768,I670760);
nor I_39308 (I670785,I670768,I670666);
and I_39309 (I670802,I670785,I579297);
nor I_39310 (I670819,I670768,I670734);
nor I_39311 (I670615,I670726,I670819);
DFFARX1 I_39312 (I579291,I2507,I670632,I670859,);
nor I_39313 (I670867,I670859,I670726);
not I_39314 (I670884,I670867);
not I_39315 (I670901,I670859);
nor I_39316 (I670918,I670901,I670802);
DFFARX1 I_39317 (I670918,I2507,I670632,I670618,);
nand I_39318 (I670949,I579288,I579279);
and I_39319 (I670966,I670949,I579276);
DFFARX1 I_39320 (I670966,I2507,I670632,I670992,);
nor I_39321 (I671000,I670992,I670859);
DFFARX1 I_39322 (I671000,I2507,I670632,I670600,);
nand I_39323 (I671031,I670992,I670901);
nand I_39324 (I670609,I670884,I671031);
not I_39325 (I671062,I670992);
nor I_39326 (I671079,I671062,I670802);
DFFARX1 I_39327 (I671079,I2507,I670632,I670621,);
nor I_39328 (I671110,I579279,I579279);
or I_39329 (I670612,I670859,I671110);
nor I_39330 (I670603,I670992,I671110);
or I_39331 (I670606,I670726,I671110);
DFFARX1 I_39332 (I671110,I2507,I670632,I670624,);
not I_39333 (I671210,I2514);
DFFARX1 I_39334 (I1150868,I2507,I671210,I671236,);
not I_39335 (I671244,I671236);
nand I_39336 (I671261,I1150850,I1150862);
and I_39337 (I671278,I671261,I1150865);
DFFARX1 I_39338 (I671278,I2507,I671210,I671304,);
not I_39339 (I671312,I1150859);
DFFARX1 I_39340 (I1150856,I2507,I671210,I671338,);
not I_39341 (I671346,I671338);
nor I_39342 (I671363,I671346,I671244);
and I_39343 (I671380,I671363,I1150859);
nor I_39344 (I671397,I671346,I671312);
nor I_39345 (I671193,I671304,I671397);
DFFARX1 I_39346 (I1150874,I2507,I671210,I671437,);
nor I_39347 (I671445,I671437,I671304);
not I_39348 (I671462,I671445);
not I_39349 (I671479,I671437);
nor I_39350 (I671496,I671479,I671380);
DFFARX1 I_39351 (I671496,I2507,I671210,I671196,);
nand I_39352 (I671527,I1150853,I1150853);
and I_39353 (I671544,I671527,I1150850);
DFFARX1 I_39354 (I671544,I2507,I671210,I671570,);
nor I_39355 (I671578,I671570,I671437);
DFFARX1 I_39356 (I671578,I2507,I671210,I671178,);
nand I_39357 (I671609,I671570,I671479);
nand I_39358 (I671187,I671462,I671609);
not I_39359 (I671640,I671570);
nor I_39360 (I671657,I671640,I671380);
DFFARX1 I_39361 (I671657,I2507,I671210,I671199,);
nor I_39362 (I671688,I1150871,I1150853);
or I_39363 (I671190,I671437,I671688);
nor I_39364 (I671181,I671570,I671688);
or I_39365 (I671184,I671304,I671688);
DFFARX1 I_39366 (I671688,I2507,I671210,I671202,);
not I_39367 (I671788,I2514);
DFFARX1 I_39368 (I949611,I2507,I671788,I671814,);
not I_39369 (I671822,I671814);
nand I_39370 (I671839,I949587,I949602);
and I_39371 (I671856,I671839,I949614);
DFFARX1 I_39372 (I671856,I2507,I671788,I671882,);
not I_39373 (I671890,I949599);
DFFARX1 I_39374 (I949590,I2507,I671788,I671916,);
not I_39375 (I671924,I671916);
nor I_39376 (I671941,I671924,I671822);
and I_39377 (I671958,I671941,I949599);
nor I_39378 (I671975,I671924,I671890);
nor I_39379 (I671771,I671882,I671975);
DFFARX1 I_39380 (I949587,I2507,I671788,I672015,);
nor I_39381 (I672023,I672015,I671882);
not I_39382 (I672040,I672023);
not I_39383 (I672057,I672015);
nor I_39384 (I672074,I672057,I671958);
DFFARX1 I_39385 (I672074,I2507,I671788,I671774,);
nand I_39386 (I672105,I949605,I949596);
and I_39387 (I672122,I672105,I949608);
DFFARX1 I_39388 (I672122,I2507,I671788,I672148,);
nor I_39389 (I672156,I672148,I672015);
DFFARX1 I_39390 (I672156,I2507,I671788,I671756,);
nand I_39391 (I672187,I672148,I672057);
nand I_39392 (I671765,I672040,I672187);
not I_39393 (I672218,I672148);
nor I_39394 (I672235,I672218,I671958);
DFFARX1 I_39395 (I672235,I2507,I671788,I671777,);
nor I_39396 (I672266,I949593,I949596);
or I_39397 (I671768,I672015,I672266);
nor I_39398 (I671759,I672148,I672266);
or I_39399 (I671762,I671882,I672266);
DFFARX1 I_39400 (I672266,I2507,I671788,I671780,);
not I_39401 (I672366,I2514);
DFFARX1 I_39402 (I944443,I2507,I672366,I672392,);
not I_39403 (I672400,I672392);
nand I_39404 (I672417,I944419,I944434);
and I_39405 (I672434,I672417,I944446);
DFFARX1 I_39406 (I672434,I2507,I672366,I672460,);
not I_39407 (I672468,I944431);
DFFARX1 I_39408 (I944422,I2507,I672366,I672494,);
not I_39409 (I672502,I672494);
nor I_39410 (I672519,I672502,I672400);
and I_39411 (I672536,I672519,I944431);
nor I_39412 (I672553,I672502,I672468);
nor I_39413 (I672349,I672460,I672553);
DFFARX1 I_39414 (I944419,I2507,I672366,I672593,);
nor I_39415 (I672601,I672593,I672460);
not I_39416 (I672618,I672601);
not I_39417 (I672635,I672593);
nor I_39418 (I672652,I672635,I672536);
DFFARX1 I_39419 (I672652,I2507,I672366,I672352,);
nand I_39420 (I672683,I944437,I944428);
and I_39421 (I672700,I672683,I944440);
DFFARX1 I_39422 (I672700,I2507,I672366,I672726,);
nor I_39423 (I672734,I672726,I672593);
DFFARX1 I_39424 (I672734,I2507,I672366,I672334,);
nand I_39425 (I672765,I672726,I672635);
nand I_39426 (I672343,I672618,I672765);
not I_39427 (I672796,I672726);
nor I_39428 (I672813,I672796,I672536);
DFFARX1 I_39429 (I672813,I2507,I672366,I672355,);
nor I_39430 (I672844,I944425,I944428);
or I_39431 (I672346,I672593,I672844);
nor I_39432 (I672337,I672726,I672844);
or I_39433 (I672340,I672460,I672844);
DFFARX1 I_39434 (I672844,I2507,I672366,I672358,);
not I_39435 (I672944,I2514);
DFFARX1 I_39436 (I233530,I2507,I672944,I672970,);
not I_39437 (I672978,I672970);
nand I_39438 (I672995,I233533,I233554);
and I_39439 (I673012,I672995,I233542);
DFFARX1 I_39440 (I673012,I2507,I672944,I673038,);
not I_39441 (I673046,I233539);
DFFARX1 I_39442 (I233530,I2507,I672944,I673072,);
not I_39443 (I673080,I673072);
nor I_39444 (I673097,I673080,I672978);
and I_39445 (I673114,I673097,I233539);
nor I_39446 (I673131,I673080,I673046);
nor I_39447 (I672927,I673038,I673131);
DFFARX1 I_39448 (I233548,I2507,I672944,I673171,);
nor I_39449 (I673179,I673171,I673038);
not I_39450 (I673196,I673179);
not I_39451 (I673213,I673171);
nor I_39452 (I673230,I673213,I673114);
DFFARX1 I_39453 (I673230,I2507,I672944,I672930,);
nand I_39454 (I673261,I233533,I233536);
and I_39455 (I673278,I673261,I233545);
DFFARX1 I_39456 (I673278,I2507,I672944,I673304,);
nor I_39457 (I673312,I673304,I673171);
DFFARX1 I_39458 (I673312,I2507,I672944,I672912,);
nand I_39459 (I673343,I673304,I673213);
nand I_39460 (I672921,I673196,I673343);
not I_39461 (I673374,I673304);
nor I_39462 (I673391,I673374,I673114);
DFFARX1 I_39463 (I673391,I2507,I672944,I672933,);
nor I_39464 (I673422,I233551,I233536);
or I_39465 (I672924,I673171,I673422);
nor I_39466 (I672915,I673304,I673422);
or I_39467 (I672918,I673038,I673422);
DFFARX1 I_39468 (I673422,I2507,I672944,I672936,);
not I_39469 (I673522,I2514);
DFFARX1 I_39470 (I1000645,I2507,I673522,I673548,);
not I_39471 (I673556,I673548);
nand I_39472 (I673573,I1000621,I1000636);
and I_39473 (I673590,I673573,I1000648);
DFFARX1 I_39474 (I673590,I2507,I673522,I673616,);
not I_39475 (I673624,I1000633);
DFFARX1 I_39476 (I1000624,I2507,I673522,I673650,);
not I_39477 (I673658,I673650);
nor I_39478 (I673675,I673658,I673556);
and I_39479 (I673692,I673675,I1000633);
nor I_39480 (I673709,I673658,I673624);
nor I_39481 (I673505,I673616,I673709);
DFFARX1 I_39482 (I1000621,I2507,I673522,I673749,);
nor I_39483 (I673757,I673749,I673616);
not I_39484 (I673774,I673757);
not I_39485 (I673791,I673749);
nor I_39486 (I673808,I673791,I673692);
DFFARX1 I_39487 (I673808,I2507,I673522,I673508,);
nand I_39488 (I673839,I1000639,I1000630);
and I_39489 (I673856,I673839,I1000642);
DFFARX1 I_39490 (I673856,I2507,I673522,I673882,);
nor I_39491 (I673890,I673882,I673749);
DFFARX1 I_39492 (I673890,I2507,I673522,I673490,);
nand I_39493 (I673921,I673882,I673791);
nand I_39494 (I673499,I673774,I673921);
not I_39495 (I673952,I673882);
nor I_39496 (I673969,I673952,I673692);
DFFARX1 I_39497 (I673969,I2507,I673522,I673511,);
nor I_39498 (I674000,I1000627,I1000630);
or I_39499 (I673502,I673749,I674000);
nor I_39500 (I673493,I673882,I674000);
or I_39501 (I673496,I673616,I674000);
DFFARX1 I_39502 (I674000,I2507,I673522,I673514,);
not I_39503 (I674100,I2514);
DFFARX1 I_39504 (I1314264,I2507,I674100,I674126,);
not I_39505 (I674134,I674126);
nand I_39506 (I674151,I1314249,I1314237);
and I_39507 (I674168,I674151,I1314252);
DFFARX1 I_39508 (I674168,I2507,I674100,I674194,);
not I_39509 (I674202,I1314237);
DFFARX1 I_39510 (I1314255,I2507,I674100,I674228,);
not I_39511 (I674236,I674228);
nor I_39512 (I674253,I674236,I674134);
and I_39513 (I674270,I674253,I1314237);
nor I_39514 (I674287,I674236,I674202);
nor I_39515 (I674083,I674194,I674287);
DFFARX1 I_39516 (I1314243,I2507,I674100,I674327,);
nor I_39517 (I674335,I674327,I674194);
not I_39518 (I674352,I674335);
not I_39519 (I674369,I674327);
nor I_39520 (I674386,I674369,I674270);
DFFARX1 I_39521 (I674386,I2507,I674100,I674086,);
nand I_39522 (I674417,I1314240,I1314246);
and I_39523 (I674434,I674417,I1314261);
DFFARX1 I_39524 (I674434,I2507,I674100,I674460,);
nor I_39525 (I674468,I674460,I674327);
DFFARX1 I_39526 (I674468,I2507,I674100,I674068,);
nand I_39527 (I674499,I674460,I674369);
nand I_39528 (I674077,I674352,I674499);
not I_39529 (I674530,I674460);
nor I_39530 (I674547,I674530,I674270);
DFFARX1 I_39531 (I674547,I2507,I674100,I674089,);
nor I_39532 (I674578,I1314258,I1314246);
or I_39533 (I674080,I674327,I674578);
nor I_39534 (I674071,I674460,I674578);
or I_39535 (I674074,I674194,I674578);
DFFARX1 I_39536 (I674578,I2507,I674100,I674092,);
not I_39537 (I674678,I2514);
DFFARX1 I_39538 (I137152,I2507,I674678,I674704,);
not I_39539 (I674712,I674704);
nand I_39540 (I674729,I137167,I137140);
and I_39541 (I674746,I674729,I137155);
DFFARX1 I_39542 (I674746,I2507,I674678,I674772,);
not I_39543 (I674780,I137158);
DFFARX1 I_39544 (I137143,I2507,I674678,I674806,);
not I_39545 (I674814,I674806);
nor I_39546 (I674831,I674814,I674712);
and I_39547 (I674848,I674831,I137158);
nor I_39548 (I674865,I674814,I674780);
nor I_39549 (I674661,I674772,I674865);
DFFARX1 I_39550 (I137149,I2507,I674678,I674905,);
nor I_39551 (I674913,I674905,I674772);
not I_39552 (I674930,I674913);
not I_39553 (I674947,I674905);
nor I_39554 (I674964,I674947,I674848);
DFFARX1 I_39555 (I674964,I2507,I674678,I674664,);
nand I_39556 (I674995,I137164,I137146);
and I_39557 (I675012,I674995,I137161);
DFFARX1 I_39558 (I675012,I2507,I674678,I675038,);
nor I_39559 (I675046,I675038,I674905);
DFFARX1 I_39560 (I675046,I2507,I674678,I674646,);
nand I_39561 (I675077,I675038,I674947);
nand I_39562 (I674655,I674930,I675077);
not I_39563 (I675108,I675038);
nor I_39564 (I675125,I675108,I674848);
DFFARX1 I_39565 (I675125,I2507,I674678,I674667,);
nor I_39566 (I675156,I137140,I137146);
or I_39567 (I674658,I674905,I675156);
nor I_39568 (I674649,I675038,I675156);
or I_39569 (I674652,I674772,I675156);
DFFARX1 I_39570 (I675156,I2507,I674678,I674670,);
not I_39571 (I675256,I2514);
DFFARX1 I_39572 (I1135262,I2507,I675256,I675282,);
not I_39573 (I675290,I675282);
nand I_39574 (I675307,I1135244,I1135256);
and I_39575 (I675324,I675307,I1135259);
DFFARX1 I_39576 (I675324,I2507,I675256,I675350,);
not I_39577 (I675358,I1135253);
DFFARX1 I_39578 (I1135250,I2507,I675256,I675384,);
not I_39579 (I675392,I675384);
nor I_39580 (I675409,I675392,I675290);
and I_39581 (I675426,I675409,I1135253);
nor I_39582 (I675443,I675392,I675358);
nor I_39583 (I675239,I675350,I675443);
DFFARX1 I_39584 (I1135268,I2507,I675256,I675483,);
nor I_39585 (I675491,I675483,I675350);
not I_39586 (I675508,I675491);
not I_39587 (I675525,I675483);
nor I_39588 (I675542,I675525,I675426);
DFFARX1 I_39589 (I675542,I2507,I675256,I675242,);
nand I_39590 (I675573,I1135247,I1135247);
and I_39591 (I675590,I675573,I1135244);
DFFARX1 I_39592 (I675590,I2507,I675256,I675616,);
nor I_39593 (I675624,I675616,I675483);
DFFARX1 I_39594 (I675624,I2507,I675256,I675224,);
nand I_39595 (I675655,I675616,I675525);
nand I_39596 (I675233,I675508,I675655);
not I_39597 (I675686,I675616);
nor I_39598 (I675703,I675686,I675426);
DFFARX1 I_39599 (I675703,I2507,I675256,I675245,);
nor I_39600 (I675734,I1135265,I1135247);
or I_39601 (I675236,I675483,I675734);
nor I_39602 (I675227,I675616,I675734);
or I_39603 (I675230,I675350,I675734);
DFFARX1 I_39604 (I675734,I2507,I675256,I675248,);
not I_39605 (I675834,I2514);
DFFARX1 I_39606 (I981265,I2507,I675834,I675860,);
not I_39607 (I675868,I675860);
nand I_39608 (I675885,I981241,I981256);
and I_39609 (I675902,I675885,I981268);
DFFARX1 I_39610 (I675902,I2507,I675834,I675928,);
not I_39611 (I675936,I981253);
DFFARX1 I_39612 (I981244,I2507,I675834,I675962,);
not I_39613 (I675970,I675962);
nor I_39614 (I675987,I675970,I675868);
and I_39615 (I676004,I675987,I981253);
nor I_39616 (I676021,I675970,I675936);
nor I_39617 (I675817,I675928,I676021);
DFFARX1 I_39618 (I981241,I2507,I675834,I676061,);
nor I_39619 (I676069,I676061,I675928);
not I_39620 (I676086,I676069);
not I_39621 (I676103,I676061);
nor I_39622 (I676120,I676103,I676004);
DFFARX1 I_39623 (I676120,I2507,I675834,I675820,);
nand I_39624 (I676151,I981259,I981250);
and I_39625 (I676168,I676151,I981262);
DFFARX1 I_39626 (I676168,I2507,I675834,I676194,);
nor I_39627 (I676202,I676194,I676061);
DFFARX1 I_39628 (I676202,I2507,I675834,I675802,);
nand I_39629 (I676233,I676194,I676103);
nand I_39630 (I675811,I676086,I676233);
not I_39631 (I676264,I676194);
nor I_39632 (I676281,I676264,I676004);
DFFARX1 I_39633 (I676281,I2507,I675834,I675823,);
nor I_39634 (I676312,I981247,I981250);
or I_39635 (I675814,I676061,I676312);
nor I_39636 (I675805,I676194,I676312);
or I_39637 (I675808,I675928,I676312);
DFFARX1 I_39638 (I676312,I2507,I675834,I675826,);
not I_39639 (I676412,I2514);
DFFARX1 I_39640 (I151420,I2507,I676412,I676438,);
not I_39641 (I676446,I676438);
nand I_39642 (I676463,I151423,I151444);
and I_39643 (I676480,I676463,I151432);
DFFARX1 I_39644 (I676480,I2507,I676412,I676506,);
not I_39645 (I676514,I151429);
DFFARX1 I_39646 (I151420,I2507,I676412,I676540,);
not I_39647 (I676548,I676540);
nor I_39648 (I676565,I676548,I676446);
and I_39649 (I676582,I676565,I151429);
nor I_39650 (I676599,I676548,I676514);
nor I_39651 (I676395,I676506,I676599);
DFFARX1 I_39652 (I151438,I2507,I676412,I676639,);
nor I_39653 (I676647,I676639,I676506);
not I_39654 (I676664,I676647);
not I_39655 (I676681,I676639);
nor I_39656 (I676698,I676681,I676582);
DFFARX1 I_39657 (I676698,I2507,I676412,I676398,);
nand I_39658 (I676729,I151423,I151426);
and I_39659 (I676746,I676729,I151435);
DFFARX1 I_39660 (I676746,I2507,I676412,I676772,);
nor I_39661 (I676780,I676772,I676639);
DFFARX1 I_39662 (I676780,I2507,I676412,I676380,);
nand I_39663 (I676811,I676772,I676681);
nand I_39664 (I676389,I676664,I676811);
not I_39665 (I676842,I676772);
nor I_39666 (I676859,I676842,I676582);
DFFARX1 I_39667 (I676859,I2507,I676412,I676401,);
nor I_39668 (I676890,I151441,I151426);
or I_39669 (I676392,I676639,I676890);
nor I_39670 (I676383,I676772,I676890);
or I_39671 (I676386,I676506,I676890);
DFFARX1 I_39672 (I676890,I2507,I676412,I676404,);
not I_39673 (I676990,I2514);
DFFARX1 I_39674 (I1335089,I2507,I676990,I677016,);
not I_39675 (I677024,I677016);
nand I_39676 (I677041,I1335074,I1335062);
and I_39677 (I677058,I677041,I1335077);
DFFARX1 I_39678 (I677058,I2507,I676990,I677084,);
not I_39679 (I677092,I1335062);
DFFARX1 I_39680 (I1335080,I2507,I676990,I677118,);
not I_39681 (I677126,I677118);
nor I_39682 (I677143,I677126,I677024);
and I_39683 (I677160,I677143,I1335062);
nor I_39684 (I677177,I677126,I677092);
nor I_39685 (I676973,I677084,I677177);
DFFARX1 I_39686 (I1335068,I2507,I676990,I677217,);
nor I_39687 (I677225,I677217,I677084);
not I_39688 (I677242,I677225);
not I_39689 (I677259,I677217);
nor I_39690 (I677276,I677259,I677160);
DFFARX1 I_39691 (I677276,I2507,I676990,I676976,);
nand I_39692 (I677307,I1335065,I1335071);
and I_39693 (I677324,I677307,I1335086);
DFFARX1 I_39694 (I677324,I2507,I676990,I677350,);
nor I_39695 (I677358,I677350,I677217);
DFFARX1 I_39696 (I677358,I2507,I676990,I676958,);
nand I_39697 (I677389,I677350,I677259);
nand I_39698 (I676967,I677242,I677389);
not I_39699 (I677420,I677350);
nor I_39700 (I677437,I677420,I677160);
DFFARX1 I_39701 (I677437,I2507,I676990,I676979,);
nor I_39702 (I677468,I1335083,I1335071);
or I_39703 (I676970,I677217,I677468);
nor I_39704 (I676961,I677350,I677468);
or I_39705 (I676964,I677084,I677468);
DFFARX1 I_39706 (I677468,I2507,I676990,I676982,);
not I_39707 (I677568,I2514);
DFFARX1 I_39708 (I853382,I2507,I677568,I677594,);
not I_39709 (I677602,I677594);
nand I_39710 (I677619,I853370,I853388);
and I_39711 (I677636,I677619,I853385);
DFFARX1 I_39712 (I677636,I2507,I677568,I677662,);
not I_39713 (I677670,I853376);
DFFARX1 I_39714 (I853373,I2507,I677568,I677696,);
not I_39715 (I677704,I677696);
nor I_39716 (I677721,I677704,I677602);
and I_39717 (I677738,I677721,I853376);
nor I_39718 (I677755,I677704,I677670);
nor I_39719 (I677551,I677662,I677755);
DFFARX1 I_39720 (I853367,I2507,I677568,I677795,);
nor I_39721 (I677803,I677795,I677662);
not I_39722 (I677820,I677803);
not I_39723 (I677837,I677795);
nor I_39724 (I677854,I677837,I677738);
DFFARX1 I_39725 (I677854,I2507,I677568,I677554,);
nand I_39726 (I677885,I853367,I853370);
and I_39727 (I677902,I677885,I853373);
DFFARX1 I_39728 (I677902,I2507,I677568,I677928,);
nor I_39729 (I677936,I677928,I677795);
DFFARX1 I_39730 (I677936,I2507,I677568,I677536,);
nand I_39731 (I677967,I677928,I677837);
nand I_39732 (I677545,I677820,I677967);
not I_39733 (I677998,I677928);
nor I_39734 (I678015,I677998,I677738);
DFFARX1 I_39735 (I678015,I2507,I677568,I677557,);
nor I_39736 (I678046,I853379,I853370);
or I_39737 (I677548,I677795,I678046);
nor I_39738 (I677539,I677928,I678046);
or I_39739 (I677542,I677662,I678046);
DFFARX1 I_39740 (I678046,I2507,I677568,I677560,);
not I_39741 (I678146,I2514);
DFFARX1 I_39742 (I1182080,I2507,I678146,I678172,);
not I_39743 (I678180,I678172);
nand I_39744 (I678197,I1182062,I1182074);
and I_39745 (I678214,I678197,I1182077);
DFFARX1 I_39746 (I678214,I2507,I678146,I678240,);
not I_39747 (I678248,I1182071);
DFFARX1 I_39748 (I1182068,I2507,I678146,I678274,);
not I_39749 (I678282,I678274);
nor I_39750 (I678299,I678282,I678180);
and I_39751 (I678316,I678299,I1182071);
nor I_39752 (I678333,I678282,I678248);
nor I_39753 (I678129,I678240,I678333);
DFFARX1 I_39754 (I1182086,I2507,I678146,I678373,);
nor I_39755 (I678381,I678373,I678240);
not I_39756 (I678398,I678381);
not I_39757 (I678415,I678373);
nor I_39758 (I678432,I678415,I678316);
DFFARX1 I_39759 (I678432,I2507,I678146,I678132,);
nand I_39760 (I678463,I1182065,I1182065);
and I_39761 (I678480,I678463,I1182062);
DFFARX1 I_39762 (I678480,I2507,I678146,I678506,);
nor I_39763 (I678514,I678506,I678373);
DFFARX1 I_39764 (I678514,I2507,I678146,I678114,);
nand I_39765 (I678545,I678506,I678415);
nand I_39766 (I678123,I678398,I678545);
not I_39767 (I678576,I678506);
nor I_39768 (I678593,I678576,I678316);
DFFARX1 I_39769 (I678593,I2507,I678146,I678135,);
nor I_39770 (I678624,I1182083,I1182065);
or I_39771 (I678126,I678373,I678624);
nor I_39772 (I678117,I678506,I678624);
or I_39773 (I678120,I678240,I678624);
DFFARX1 I_39774 (I678624,I2507,I678146,I678138,);
not I_39775 (I678724,I2514);
DFFARX1 I_39776 (I1153180,I2507,I678724,I678750,);
not I_39777 (I678758,I678750);
nand I_39778 (I678775,I1153162,I1153174);
and I_39779 (I678792,I678775,I1153177);
DFFARX1 I_39780 (I678792,I2507,I678724,I678818,);
not I_39781 (I678826,I1153171);
DFFARX1 I_39782 (I1153168,I2507,I678724,I678852,);
not I_39783 (I678860,I678852);
nor I_39784 (I678877,I678860,I678758);
and I_39785 (I678894,I678877,I1153171);
nor I_39786 (I678911,I678860,I678826);
nor I_39787 (I678707,I678818,I678911);
DFFARX1 I_39788 (I1153186,I2507,I678724,I678951,);
nor I_39789 (I678959,I678951,I678818);
not I_39790 (I678976,I678959);
not I_39791 (I678993,I678951);
nor I_39792 (I679010,I678993,I678894);
DFFARX1 I_39793 (I679010,I2507,I678724,I678710,);
nand I_39794 (I679041,I1153165,I1153165);
and I_39795 (I679058,I679041,I1153162);
DFFARX1 I_39796 (I679058,I2507,I678724,I679084,);
nor I_39797 (I679092,I679084,I678951);
DFFARX1 I_39798 (I679092,I2507,I678724,I678692,);
nand I_39799 (I679123,I679084,I678993);
nand I_39800 (I678701,I678976,I679123);
not I_39801 (I679154,I679084);
nor I_39802 (I679171,I679154,I678894);
DFFARX1 I_39803 (I679171,I2507,I678724,I678713,);
nor I_39804 (I679202,I1153183,I1153165);
or I_39805 (I678704,I678951,I679202);
nor I_39806 (I678695,I679084,I679202);
or I_39807 (I678698,I678818,I679202);
DFFARX1 I_39808 (I679202,I2507,I678724,I678716,);
not I_39809 (I679302,I2514);
DFFARX1 I_39810 (I531574,I2507,I679302,I679328,);
not I_39811 (I679336,I679328);
nand I_39812 (I679353,I531589,I531574);
and I_39813 (I679370,I679353,I531577);
DFFARX1 I_39814 (I679370,I2507,I679302,I679396,);
not I_39815 (I679404,I531577);
DFFARX1 I_39816 (I531586,I2507,I679302,I679430,);
not I_39817 (I679438,I679430);
nor I_39818 (I679455,I679438,I679336);
and I_39819 (I679472,I679455,I531577);
nor I_39820 (I679489,I679438,I679404);
nor I_39821 (I679285,I679396,I679489);
DFFARX1 I_39822 (I531580,I2507,I679302,I679529,);
nor I_39823 (I679537,I679529,I679396);
not I_39824 (I679554,I679537);
not I_39825 (I679571,I679529);
nor I_39826 (I679588,I679571,I679472);
DFFARX1 I_39827 (I679588,I2507,I679302,I679288,);
nand I_39828 (I679619,I531583,I531592);
and I_39829 (I679636,I679619,I531598);
DFFARX1 I_39830 (I679636,I2507,I679302,I679662,);
nor I_39831 (I679670,I679662,I679529);
DFFARX1 I_39832 (I679670,I2507,I679302,I679270,);
nand I_39833 (I679701,I679662,I679571);
nand I_39834 (I679279,I679554,I679701);
not I_39835 (I679732,I679662);
nor I_39836 (I679749,I679732,I679472);
DFFARX1 I_39837 (I679749,I2507,I679302,I679291,);
nor I_39838 (I679780,I531595,I531592);
or I_39839 (I679282,I679529,I679780);
nor I_39840 (I679273,I679662,I679780);
or I_39841 (I679276,I679396,I679780);
DFFARX1 I_39842 (I679780,I2507,I679302,I679294,);
not I_39843 (I679880,I2514);
DFFARX1 I_39844 (I105982,I2507,I679880,I679906,);
not I_39845 (I679914,I679906);
nand I_39846 (I679931,I105991,I106000);
and I_39847 (I679948,I679931,I105979);
DFFARX1 I_39848 (I679948,I2507,I679880,I679974,);
not I_39849 (I679982,I105982);
DFFARX1 I_39850 (I105997,I2507,I679880,I680008,);
not I_39851 (I680016,I680008);
nor I_39852 (I680033,I680016,I679914);
and I_39853 (I680050,I680033,I105982);
nor I_39854 (I680067,I680016,I679982);
nor I_39855 (I679863,I679974,I680067);
DFFARX1 I_39856 (I105988,I2507,I679880,I680107,);
nor I_39857 (I680115,I680107,I679974);
not I_39858 (I680132,I680115);
not I_39859 (I680149,I680107);
nor I_39860 (I680166,I680149,I680050);
DFFARX1 I_39861 (I680166,I2507,I679880,I679866,);
nand I_39862 (I680197,I106003,I105979);
and I_39863 (I680214,I680197,I105985);
DFFARX1 I_39864 (I680214,I2507,I679880,I680240,);
nor I_39865 (I680248,I680240,I680107);
DFFARX1 I_39866 (I680248,I2507,I679880,I679848,);
nand I_39867 (I680279,I680240,I680149);
nand I_39868 (I679857,I680132,I680279);
not I_39869 (I680310,I680240);
nor I_39870 (I680327,I680310,I680050);
DFFARX1 I_39871 (I680327,I2507,I679880,I679869,);
nor I_39872 (I680358,I105994,I105979);
or I_39873 (I679860,I680107,I680358);
nor I_39874 (I679851,I680240,I680358);
or I_39875 (I679854,I679974,I680358);
DFFARX1 I_39876 (I680358,I2507,I679880,I679872,);
not I_39877 (I680458,I2514);
DFFARX1 I_39878 (I515509,I2507,I680458,I680484,);
not I_39879 (I680492,I680484);
nand I_39880 (I680509,I515524,I515509);
and I_39881 (I680526,I680509,I515512);
DFFARX1 I_39882 (I680526,I2507,I680458,I680552,);
not I_39883 (I680560,I515512);
DFFARX1 I_39884 (I515521,I2507,I680458,I680586,);
not I_39885 (I680594,I680586);
nor I_39886 (I680611,I680594,I680492);
and I_39887 (I680628,I680611,I515512);
nor I_39888 (I680645,I680594,I680560);
nor I_39889 (I680441,I680552,I680645);
DFFARX1 I_39890 (I515515,I2507,I680458,I680685,);
nor I_39891 (I680693,I680685,I680552);
not I_39892 (I680710,I680693);
not I_39893 (I680727,I680685);
nor I_39894 (I680744,I680727,I680628);
DFFARX1 I_39895 (I680744,I2507,I680458,I680444,);
nand I_39896 (I680775,I515518,I515527);
and I_39897 (I680792,I680775,I515533);
DFFARX1 I_39898 (I680792,I2507,I680458,I680818,);
nor I_39899 (I680826,I680818,I680685);
DFFARX1 I_39900 (I680826,I2507,I680458,I680426,);
nand I_39901 (I680857,I680818,I680727);
nand I_39902 (I680435,I680710,I680857);
not I_39903 (I680888,I680818);
nor I_39904 (I680905,I680888,I680628);
DFFARX1 I_39905 (I680905,I2507,I680458,I680447,);
nor I_39906 (I680936,I515530,I515527);
or I_39907 (I680438,I680685,I680936);
nor I_39908 (I680429,I680818,I680936);
or I_39909 (I680432,I680552,I680936);
DFFARX1 I_39910 (I680936,I2507,I680458,I680450,);
not I_39911 (I681036,I2514);
DFFARX1 I_39912 (I496469,I2507,I681036,I681062,);
not I_39913 (I681070,I681062);
nand I_39914 (I681087,I496484,I496469);
and I_39915 (I681104,I681087,I496472);
DFFARX1 I_39916 (I681104,I2507,I681036,I681130,);
not I_39917 (I681138,I496472);
DFFARX1 I_39918 (I496481,I2507,I681036,I681164,);
not I_39919 (I681172,I681164);
nor I_39920 (I681189,I681172,I681070);
and I_39921 (I681206,I681189,I496472);
nor I_39922 (I681223,I681172,I681138);
nor I_39923 (I681019,I681130,I681223);
DFFARX1 I_39924 (I496475,I2507,I681036,I681263,);
nor I_39925 (I681271,I681263,I681130);
not I_39926 (I681288,I681271);
not I_39927 (I681305,I681263);
nor I_39928 (I681322,I681305,I681206);
DFFARX1 I_39929 (I681322,I2507,I681036,I681022,);
nand I_39930 (I681353,I496478,I496487);
and I_39931 (I681370,I681353,I496493);
DFFARX1 I_39932 (I681370,I2507,I681036,I681396,);
nor I_39933 (I681404,I681396,I681263);
DFFARX1 I_39934 (I681404,I2507,I681036,I681004,);
nand I_39935 (I681435,I681396,I681305);
nand I_39936 (I681013,I681288,I681435);
not I_39937 (I681466,I681396);
nor I_39938 (I681483,I681466,I681206);
DFFARX1 I_39939 (I681483,I2507,I681036,I681025,);
nor I_39940 (I681514,I496490,I496487);
or I_39941 (I681016,I681263,I681514);
nor I_39942 (I681007,I681396,I681514);
or I_39943 (I681010,I681130,I681514);
DFFARX1 I_39944 (I681514,I2507,I681036,I681028,);
not I_39945 (I681614,I2514);
DFFARX1 I_39946 (I228175,I2507,I681614,I681640,);
not I_39947 (I681648,I681640);
nand I_39948 (I681665,I228178,I228199);
and I_39949 (I681682,I681665,I228187);
DFFARX1 I_39950 (I681682,I2507,I681614,I681708,);
not I_39951 (I681716,I228184);
DFFARX1 I_39952 (I228175,I2507,I681614,I681742,);
not I_39953 (I681750,I681742);
nor I_39954 (I681767,I681750,I681648);
and I_39955 (I681784,I681767,I228184);
nor I_39956 (I681801,I681750,I681716);
nor I_39957 (I681597,I681708,I681801);
DFFARX1 I_39958 (I228193,I2507,I681614,I681841,);
nor I_39959 (I681849,I681841,I681708);
not I_39960 (I681866,I681849);
not I_39961 (I681883,I681841);
nor I_39962 (I681900,I681883,I681784);
DFFARX1 I_39963 (I681900,I2507,I681614,I681600,);
nand I_39964 (I681931,I228178,I228181);
and I_39965 (I681948,I681931,I228190);
DFFARX1 I_39966 (I681948,I2507,I681614,I681974,);
nor I_39967 (I681982,I681974,I681841);
DFFARX1 I_39968 (I681982,I2507,I681614,I681582,);
nand I_39969 (I682013,I681974,I681883);
nand I_39970 (I681591,I681866,I682013);
not I_39971 (I682044,I681974);
nor I_39972 (I682061,I682044,I681784);
DFFARX1 I_39973 (I682061,I2507,I681614,I681603,);
nor I_39974 (I682092,I228196,I228181);
or I_39975 (I681594,I681841,I682092);
nor I_39976 (I681585,I681974,I682092);
or I_39977 (I681588,I681708,I682092);
DFFARX1 I_39978 (I682092,I2507,I681614,I681606,);
not I_39979 (I682192,I2514);
DFFARX1 I_39980 (I615690,I2507,I682192,I682218,);
not I_39981 (I682226,I682218);
nand I_39982 (I682243,I615699,I615708);
and I_39983 (I682260,I682243,I615714);
DFFARX1 I_39984 (I682260,I2507,I682192,I682286,);
not I_39985 (I682294,I615711);
DFFARX1 I_39986 (I615696,I2507,I682192,I682320,);
not I_39987 (I682328,I682320);
nor I_39988 (I682345,I682328,I682226);
and I_39989 (I682362,I682345,I615711);
nor I_39990 (I682379,I682328,I682294);
nor I_39991 (I682175,I682286,I682379);
DFFARX1 I_39992 (I615705,I2507,I682192,I682419,);
nor I_39993 (I682427,I682419,I682286);
not I_39994 (I682444,I682427);
not I_39995 (I682461,I682419);
nor I_39996 (I682478,I682461,I682362);
DFFARX1 I_39997 (I682478,I2507,I682192,I682178,);
nand I_39998 (I682509,I615702,I615693);
and I_39999 (I682526,I682509,I615690);
DFFARX1 I_40000 (I682526,I2507,I682192,I682552,);
nor I_40001 (I682560,I682552,I682419);
DFFARX1 I_40002 (I682560,I2507,I682192,I682160,);
nand I_40003 (I682591,I682552,I682461);
nand I_40004 (I682169,I682444,I682591);
not I_40005 (I682622,I682552);
nor I_40006 (I682639,I682622,I682362);
DFFARX1 I_40007 (I682639,I2507,I682192,I682181,);
nor I_40008 (I682670,I615693,I615693);
or I_40009 (I682172,I682419,I682670);
nor I_40010 (I682163,I682552,I682670);
or I_40011 (I682166,I682286,I682670);
DFFARX1 I_40012 (I682670,I2507,I682192,I682184,);
not I_40013 (I682770,I2514);
DFFARX1 I_40014 (I1268048,I2507,I682770,I682796,);
not I_40015 (I682804,I682796);
nand I_40016 (I682821,I1268072,I1268054);
and I_40017 (I682838,I682821,I1268060);
DFFARX1 I_40018 (I682838,I2507,I682770,I682864,);
not I_40019 (I682872,I1268066);
DFFARX1 I_40020 (I1268051,I2507,I682770,I682898,);
not I_40021 (I682906,I682898);
nor I_40022 (I682923,I682906,I682804);
and I_40023 (I682940,I682923,I1268066);
nor I_40024 (I682957,I682906,I682872);
nor I_40025 (I682753,I682864,I682957);
DFFARX1 I_40026 (I1268063,I2507,I682770,I682997,);
nor I_40027 (I683005,I682997,I682864);
not I_40028 (I683022,I683005);
not I_40029 (I683039,I682997);
nor I_40030 (I683056,I683039,I682940);
DFFARX1 I_40031 (I683056,I2507,I682770,I682756,);
nand I_40032 (I683087,I1268069,I1268057);
and I_40033 (I683104,I683087,I1268051);
DFFARX1 I_40034 (I683104,I2507,I682770,I683130,);
nor I_40035 (I683138,I683130,I682997);
DFFARX1 I_40036 (I683138,I2507,I682770,I682738,);
nand I_40037 (I683169,I683130,I683039);
nand I_40038 (I682747,I683022,I683169);
not I_40039 (I683200,I683130);
nor I_40040 (I683217,I683200,I682940);
DFFARX1 I_40041 (I683217,I2507,I682770,I682759,);
nor I_40042 (I683248,I1268048,I1268057);
or I_40043 (I682750,I682997,I683248);
nor I_40044 (I682741,I683130,I683248);
or I_40045 (I682744,I682864,I683248);
DFFARX1 I_40046 (I683248,I2507,I682770,I682762,);
not I_40047 (I683348,I2514);
DFFARX1 I_40048 (I203185,I2507,I683348,I683374,);
not I_40049 (I683382,I683374);
nand I_40050 (I683399,I203188,I203209);
and I_40051 (I683416,I683399,I203197);
DFFARX1 I_40052 (I683416,I2507,I683348,I683442,);
not I_40053 (I683450,I203194);
DFFARX1 I_40054 (I203185,I2507,I683348,I683476,);
not I_40055 (I683484,I683476);
nor I_40056 (I683501,I683484,I683382);
and I_40057 (I683518,I683501,I203194);
nor I_40058 (I683535,I683484,I683450);
nor I_40059 (I683331,I683442,I683535);
DFFARX1 I_40060 (I203203,I2507,I683348,I683575,);
nor I_40061 (I683583,I683575,I683442);
not I_40062 (I683600,I683583);
not I_40063 (I683617,I683575);
nor I_40064 (I683634,I683617,I683518);
DFFARX1 I_40065 (I683634,I2507,I683348,I683334,);
nand I_40066 (I683665,I203188,I203191);
and I_40067 (I683682,I683665,I203200);
DFFARX1 I_40068 (I683682,I2507,I683348,I683708,);
nor I_40069 (I683716,I683708,I683575);
DFFARX1 I_40070 (I683716,I2507,I683348,I683316,);
nand I_40071 (I683747,I683708,I683617);
nand I_40072 (I683325,I683600,I683747);
not I_40073 (I683778,I683708);
nor I_40074 (I683795,I683778,I683518);
DFFARX1 I_40075 (I683795,I2507,I683348,I683337,);
nor I_40076 (I683826,I203206,I203191);
or I_40077 (I683328,I683575,I683826);
nor I_40078 (I683319,I683708,I683826);
or I_40079 (I683322,I683442,I683826);
DFFARX1 I_40080 (I683826,I2507,I683348,I683340,);
not I_40081 (I683926,I2514);
DFFARX1 I_40082 (I1095380,I2507,I683926,I683952,);
not I_40083 (I683960,I683952);
nand I_40084 (I683977,I1095362,I1095374);
and I_40085 (I683994,I683977,I1095377);
DFFARX1 I_40086 (I683994,I2507,I683926,I684020,);
not I_40087 (I684028,I1095371);
DFFARX1 I_40088 (I1095368,I2507,I683926,I684054,);
not I_40089 (I684062,I684054);
nor I_40090 (I684079,I684062,I683960);
and I_40091 (I684096,I684079,I1095371);
nor I_40092 (I684113,I684062,I684028);
nor I_40093 (I683909,I684020,I684113);
DFFARX1 I_40094 (I1095386,I2507,I683926,I684153,);
nor I_40095 (I684161,I684153,I684020);
not I_40096 (I684178,I684161);
not I_40097 (I684195,I684153);
nor I_40098 (I684212,I684195,I684096);
DFFARX1 I_40099 (I684212,I2507,I683926,I683912,);
nand I_40100 (I684243,I1095365,I1095365);
and I_40101 (I684260,I684243,I1095362);
DFFARX1 I_40102 (I684260,I2507,I683926,I684286,);
nor I_40103 (I684294,I684286,I684153);
DFFARX1 I_40104 (I684294,I2507,I683926,I683894,);
nand I_40105 (I684325,I684286,I684195);
nand I_40106 (I683903,I684178,I684325);
not I_40107 (I684356,I684286);
nor I_40108 (I684373,I684356,I684096);
DFFARX1 I_40109 (I684373,I2507,I683926,I683915,);
nor I_40110 (I684404,I1095383,I1095365);
or I_40111 (I683906,I684153,I684404);
nor I_40112 (I683897,I684286,I684404);
or I_40113 (I683900,I684020,I684404);
DFFARX1 I_40114 (I684404,I2507,I683926,I683918,);
not I_40115 (I684504,I2514);
DFFARX1 I_40116 (I225795,I2507,I684504,I684530,);
not I_40117 (I684538,I684530);
nand I_40118 (I684555,I225798,I225819);
and I_40119 (I684572,I684555,I225807);
DFFARX1 I_40120 (I684572,I2507,I684504,I684598,);
not I_40121 (I684606,I225804);
DFFARX1 I_40122 (I225795,I2507,I684504,I684632,);
not I_40123 (I684640,I684632);
nor I_40124 (I684657,I684640,I684538);
and I_40125 (I684674,I684657,I225804);
nor I_40126 (I684691,I684640,I684606);
nor I_40127 (I684487,I684598,I684691);
DFFARX1 I_40128 (I225813,I2507,I684504,I684731,);
nor I_40129 (I684739,I684731,I684598);
not I_40130 (I684756,I684739);
not I_40131 (I684773,I684731);
nor I_40132 (I684790,I684773,I684674);
DFFARX1 I_40133 (I684790,I2507,I684504,I684490,);
nand I_40134 (I684821,I225798,I225801);
and I_40135 (I684838,I684821,I225810);
DFFARX1 I_40136 (I684838,I2507,I684504,I684864,);
nor I_40137 (I684872,I684864,I684731);
DFFARX1 I_40138 (I684872,I2507,I684504,I684472,);
nand I_40139 (I684903,I684864,I684773);
nand I_40140 (I684481,I684756,I684903);
not I_40141 (I684934,I684864);
nor I_40142 (I684951,I684934,I684674);
DFFARX1 I_40143 (I684951,I2507,I684504,I684493,);
nor I_40144 (I684982,I225816,I225801);
or I_40145 (I684484,I684731,I684982);
nor I_40146 (I684475,I684864,I684982);
or I_40147 (I684478,I684598,I684982);
DFFARX1 I_40148 (I684982,I2507,I684504,I684496,);
not I_40149 (I685082,I2514);
DFFARX1 I_40150 (I958655,I2507,I685082,I685108,);
not I_40151 (I685116,I685108);
nand I_40152 (I685133,I958631,I958646);
and I_40153 (I685150,I685133,I958658);
DFFARX1 I_40154 (I685150,I2507,I685082,I685176,);
not I_40155 (I685184,I958643);
DFFARX1 I_40156 (I958634,I2507,I685082,I685210,);
not I_40157 (I685218,I685210);
nor I_40158 (I685235,I685218,I685116);
and I_40159 (I685252,I685235,I958643);
nor I_40160 (I685269,I685218,I685184);
nor I_40161 (I685065,I685176,I685269);
DFFARX1 I_40162 (I958631,I2507,I685082,I685309,);
nor I_40163 (I685317,I685309,I685176);
not I_40164 (I685334,I685317);
not I_40165 (I685351,I685309);
nor I_40166 (I685368,I685351,I685252);
DFFARX1 I_40167 (I685368,I2507,I685082,I685068,);
nand I_40168 (I685399,I958649,I958640);
and I_40169 (I685416,I685399,I958652);
DFFARX1 I_40170 (I685416,I2507,I685082,I685442,);
nor I_40171 (I685450,I685442,I685309);
DFFARX1 I_40172 (I685450,I2507,I685082,I685050,);
nand I_40173 (I685481,I685442,I685351);
nand I_40174 (I685059,I685334,I685481);
not I_40175 (I685512,I685442);
nor I_40176 (I685529,I685512,I685252);
DFFARX1 I_40177 (I685529,I2507,I685082,I685071,);
nor I_40178 (I685560,I958637,I958640);
or I_40179 (I685062,I685309,I685560);
nor I_40180 (I685053,I685442,I685560);
or I_40181 (I685056,I685176,I685560);
DFFARX1 I_40182 (I685560,I2507,I685082,I685074,);
not I_40183 (I685660,I2514);
DFFARX1 I_40184 (I39589,I2507,I685660,I685686,);
not I_40185 (I685694,I685686);
nand I_40186 (I685711,I39586,I39577);
and I_40187 (I685728,I685711,I39577);
DFFARX1 I_40188 (I685728,I2507,I685660,I685754,);
not I_40189 (I685762,I39580);
DFFARX1 I_40190 (I39595,I2507,I685660,I685788,);
not I_40191 (I685796,I685788);
nor I_40192 (I685813,I685796,I685694);
and I_40193 (I685830,I685813,I39580);
nor I_40194 (I685847,I685796,I685762);
nor I_40195 (I685643,I685754,I685847);
DFFARX1 I_40196 (I39580,I2507,I685660,I685887,);
nor I_40197 (I685895,I685887,I685754);
not I_40198 (I685912,I685895);
not I_40199 (I685929,I685887);
nor I_40200 (I685946,I685929,I685830);
DFFARX1 I_40201 (I685946,I2507,I685660,I685646,);
nand I_40202 (I685977,I39598,I39583);
and I_40203 (I685994,I685977,I39601);
DFFARX1 I_40204 (I685994,I2507,I685660,I686020,);
nor I_40205 (I686028,I686020,I685887);
DFFARX1 I_40206 (I686028,I2507,I685660,I685628,);
nand I_40207 (I686059,I686020,I685929);
nand I_40208 (I685637,I685912,I686059);
not I_40209 (I686090,I686020);
nor I_40210 (I686107,I686090,I685830);
DFFARX1 I_40211 (I686107,I2507,I685660,I685649,);
nor I_40212 (I686138,I39592,I39583);
or I_40213 (I685640,I685887,I686138);
nor I_40214 (I685631,I686020,I686138);
or I_40215 (I685634,I685754,I686138);
DFFARX1 I_40216 (I686138,I2507,I685660,I685652,);
not I_40217 (I686238,I2514);
DFFARX1 I_40218 (I1212866,I2507,I686238,I686264,);
not I_40219 (I686272,I686264);
nand I_40220 (I686289,I1212869,I1212878);
and I_40221 (I686306,I686289,I1212881);
DFFARX1 I_40222 (I686306,I2507,I686238,I686332,);
not I_40223 (I686340,I1212890);
DFFARX1 I_40224 (I1212872,I2507,I686238,I686366,);
not I_40225 (I686374,I686366);
nor I_40226 (I686391,I686374,I686272);
and I_40227 (I686408,I686391,I1212890);
nor I_40228 (I686425,I686374,I686340);
nor I_40229 (I686221,I686332,I686425);
DFFARX1 I_40230 (I1212869,I2507,I686238,I686465,);
nor I_40231 (I686473,I686465,I686332);
not I_40232 (I686490,I686473);
not I_40233 (I686507,I686465);
nor I_40234 (I686524,I686507,I686408);
DFFARX1 I_40235 (I686524,I2507,I686238,I686224,);
nand I_40236 (I686555,I1212887,I1212866);
and I_40237 (I686572,I686555,I1212884);
DFFARX1 I_40238 (I686572,I2507,I686238,I686598,);
nor I_40239 (I686606,I686598,I686465);
DFFARX1 I_40240 (I686606,I2507,I686238,I686206,);
nand I_40241 (I686637,I686598,I686507);
nand I_40242 (I686215,I686490,I686637);
not I_40243 (I686668,I686598);
nor I_40244 (I686685,I686668,I686408);
DFFARX1 I_40245 (I686685,I2507,I686238,I686227,);
nor I_40246 (I686716,I1212875,I1212866);
or I_40247 (I686218,I686465,I686716);
nor I_40248 (I686209,I686598,I686716);
or I_40249 (I686212,I686332,I686716);
DFFARX1 I_40250 (I686716,I2507,I686238,I686230,);
not I_40251 (I686816,I2514);
DFFARX1 I_40252 (I15347,I2507,I686816,I686842,);
not I_40253 (I686850,I686842);
nand I_40254 (I686867,I15344,I15335);
and I_40255 (I686884,I686867,I15335);
DFFARX1 I_40256 (I686884,I2507,I686816,I686910,);
not I_40257 (I686918,I15338);
DFFARX1 I_40258 (I15353,I2507,I686816,I686944,);
not I_40259 (I686952,I686944);
nor I_40260 (I686969,I686952,I686850);
and I_40261 (I686986,I686969,I15338);
nor I_40262 (I687003,I686952,I686918);
nor I_40263 (I686799,I686910,I687003);
DFFARX1 I_40264 (I15338,I2507,I686816,I687043,);
nor I_40265 (I687051,I687043,I686910);
not I_40266 (I687068,I687051);
not I_40267 (I687085,I687043);
nor I_40268 (I687102,I687085,I686986);
DFFARX1 I_40269 (I687102,I2507,I686816,I686802,);
nand I_40270 (I687133,I15356,I15341);
and I_40271 (I687150,I687133,I15359);
DFFARX1 I_40272 (I687150,I2507,I686816,I687176,);
nor I_40273 (I687184,I687176,I687043);
DFFARX1 I_40274 (I687184,I2507,I686816,I686784,);
nand I_40275 (I687215,I687176,I687085);
nand I_40276 (I686793,I687068,I687215);
not I_40277 (I687246,I687176);
nor I_40278 (I687263,I687246,I686986);
DFFARX1 I_40279 (I687263,I2507,I686816,I686805,);
nor I_40280 (I687294,I15350,I15341);
or I_40281 (I686796,I687043,I687294);
nor I_40282 (I686787,I687176,I687294);
or I_40283 (I686790,I686910,I687294);
DFFARX1 I_40284 (I687294,I2507,I686816,I686808,);
not I_40285 (I687394,I2514);
DFFARX1 I_40286 (I326629,I2507,I687394,I687420,);
not I_40287 (I687428,I687420);
nand I_40288 (I687445,I326632,I326608);
and I_40289 (I687462,I687445,I326605);
DFFARX1 I_40290 (I687462,I2507,I687394,I687488,);
not I_40291 (I687496,I326611);
DFFARX1 I_40292 (I326605,I2507,I687394,I687522,);
not I_40293 (I687530,I687522);
nor I_40294 (I687547,I687530,I687428);
and I_40295 (I687564,I687547,I326611);
nor I_40296 (I687581,I687530,I687496);
nor I_40297 (I687377,I687488,I687581);
DFFARX1 I_40298 (I326614,I2507,I687394,I687621,);
nor I_40299 (I687629,I687621,I687488);
not I_40300 (I687646,I687629);
not I_40301 (I687663,I687621);
nor I_40302 (I687680,I687663,I687564);
DFFARX1 I_40303 (I687680,I2507,I687394,I687380,);
nand I_40304 (I687711,I326617,I326626);
and I_40305 (I687728,I687711,I326623);
DFFARX1 I_40306 (I687728,I2507,I687394,I687754,);
nor I_40307 (I687762,I687754,I687621);
DFFARX1 I_40308 (I687762,I2507,I687394,I687362,);
nand I_40309 (I687793,I687754,I687663);
nand I_40310 (I687371,I687646,I687793);
not I_40311 (I687824,I687754);
nor I_40312 (I687841,I687824,I687564);
DFFARX1 I_40313 (I687841,I2507,I687394,I687383,);
nor I_40314 (I687872,I326620,I326626);
or I_40315 (I687374,I687621,I687872);
nor I_40316 (I687365,I687754,I687872);
or I_40317 (I687368,I687488,I687872);
DFFARX1 I_40318 (I687872,I2507,I687394,I687386,);
not I_40319 (I687972,I2514);
DFFARX1 I_40320 (I355614,I2507,I687972,I687998,);
not I_40321 (I688006,I687998);
nand I_40322 (I688023,I355617,I355593);
and I_40323 (I688040,I688023,I355590);
DFFARX1 I_40324 (I688040,I2507,I687972,I688066,);
not I_40325 (I688074,I355596);
DFFARX1 I_40326 (I355590,I2507,I687972,I688100,);
not I_40327 (I688108,I688100);
nor I_40328 (I688125,I688108,I688006);
and I_40329 (I688142,I688125,I355596);
nor I_40330 (I688159,I688108,I688074);
nor I_40331 (I687955,I688066,I688159);
DFFARX1 I_40332 (I355599,I2507,I687972,I688199,);
nor I_40333 (I688207,I688199,I688066);
not I_40334 (I688224,I688207);
not I_40335 (I688241,I688199);
nor I_40336 (I688258,I688241,I688142);
DFFARX1 I_40337 (I688258,I2507,I687972,I687958,);
nand I_40338 (I688289,I355602,I355611);
and I_40339 (I688306,I688289,I355608);
DFFARX1 I_40340 (I688306,I2507,I687972,I688332,);
nor I_40341 (I688340,I688332,I688199);
DFFARX1 I_40342 (I688340,I2507,I687972,I687940,);
nand I_40343 (I688371,I688332,I688241);
nand I_40344 (I687949,I688224,I688371);
not I_40345 (I688402,I688332);
nor I_40346 (I688419,I688402,I688142);
DFFARX1 I_40347 (I688419,I2507,I687972,I687961,);
nor I_40348 (I688450,I355605,I355611);
or I_40349 (I687952,I688199,I688450);
nor I_40350 (I687943,I688332,I688450);
or I_40351 (I687946,I688066,I688450);
DFFARX1 I_40352 (I688450,I2507,I687972,I687964,);
not I_40353 (I688550,I2514);
DFFARX1 I_40354 (I408792,I2507,I688550,I688576,);
not I_40355 (I688584,I688576);
nand I_40356 (I688601,I408783,I408801);
and I_40357 (I688618,I688601,I408804);
DFFARX1 I_40358 (I688618,I2507,I688550,I688644,);
not I_40359 (I688652,I408798);
DFFARX1 I_40360 (I408786,I2507,I688550,I688678,);
not I_40361 (I688686,I688678);
nor I_40362 (I688703,I688686,I688584);
and I_40363 (I688720,I688703,I408798);
nor I_40364 (I688737,I688686,I688652);
nor I_40365 (I688533,I688644,I688737);
DFFARX1 I_40366 (I408795,I2507,I688550,I688777,);
nor I_40367 (I688785,I688777,I688644);
not I_40368 (I688802,I688785);
not I_40369 (I688819,I688777);
nor I_40370 (I688836,I688819,I688720);
DFFARX1 I_40371 (I688836,I2507,I688550,I688536,);
nand I_40372 (I688867,I408810,I408807);
and I_40373 (I688884,I688867,I408789);
DFFARX1 I_40374 (I688884,I2507,I688550,I688910,);
nor I_40375 (I688918,I688910,I688777);
DFFARX1 I_40376 (I688918,I2507,I688550,I688518,);
nand I_40377 (I688949,I688910,I688819);
nand I_40378 (I688527,I688802,I688949);
not I_40379 (I688980,I688910);
nor I_40380 (I688997,I688980,I688720);
DFFARX1 I_40381 (I688997,I2507,I688550,I688539,);
nor I_40382 (I689028,I408783,I408807);
or I_40383 (I688530,I688777,I689028);
nor I_40384 (I688521,I688910,I689028);
or I_40385 (I688524,I688644,I689028);
DFFARX1 I_40386 (I689028,I2507,I688550,I688542,);
not I_40387 (I689128,I2514);
DFFARX1 I_40388 (I99131,I2507,I689128,I689154,);
not I_40389 (I689162,I689154);
nand I_40390 (I689179,I99140,I99149);
and I_40391 (I689196,I689179,I99128);
DFFARX1 I_40392 (I689196,I2507,I689128,I689222,);
not I_40393 (I689230,I99131);
DFFARX1 I_40394 (I99146,I2507,I689128,I689256,);
not I_40395 (I689264,I689256);
nor I_40396 (I689281,I689264,I689162);
and I_40397 (I689298,I689281,I99131);
nor I_40398 (I689315,I689264,I689230);
nor I_40399 (I689111,I689222,I689315);
DFFARX1 I_40400 (I99137,I2507,I689128,I689355,);
nor I_40401 (I689363,I689355,I689222);
not I_40402 (I689380,I689363);
not I_40403 (I689397,I689355);
nor I_40404 (I689414,I689397,I689298);
DFFARX1 I_40405 (I689414,I2507,I689128,I689114,);
nand I_40406 (I689445,I99152,I99128);
and I_40407 (I689462,I689445,I99134);
DFFARX1 I_40408 (I689462,I2507,I689128,I689488,);
nor I_40409 (I689496,I689488,I689355);
DFFARX1 I_40410 (I689496,I2507,I689128,I689096,);
nand I_40411 (I689527,I689488,I689397);
nand I_40412 (I689105,I689380,I689527);
not I_40413 (I689558,I689488);
nor I_40414 (I689575,I689558,I689298);
DFFARX1 I_40415 (I689575,I2507,I689128,I689117,);
nor I_40416 (I689606,I99143,I99128);
or I_40417 (I689108,I689355,I689606);
nor I_40418 (I689099,I689488,I689606);
or I_40419 (I689102,I689222,I689606);
DFFARX1 I_40420 (I689606,I2507,I689128,I689120,);
not I_40421 (I689706,I2514);
DFFARX1 I_40422 (I1226466,I2507,I689706,I689732,);
not I_40423 (I689740,I689732);
nand I_40424 (I689757,I1226469,I1226478);
and I_40425 (I689774,I689757,I1226481);
DFFARX1 I_40426 (I689774,I2507,I689706,I689800,);
not I_40427 (I689808,I1226490);
DFFARX1 I_40428 (I1226472,I2507,I689706,I689834,);
not I_40429 (I689842,I689834);
nor I_40430 (I689859,I689842,I689740);
and I_40431 (I689876,I689859,I1226490);
nor I_40432 (I689893,I689842,I689808);
nor I_40433 (I689689,I689800,I689893);
DFFARX1 I_40434 (I1226469,I2507,I689706,I689933,);
nor I_40435 (I689941,I689933,I689800);
not I_40436 (I689958,I689941);
not I_40437 (I689975,I689933);
nor I_40438 (I689992,I689975,I689876);
DFFARX1 I_40439 (I689992,I2507,I689706,I689692,);
nand I_40440 (I690023,I1226487,I1226466);
and I_40441 (I690040,I690023,I1226484);
DFFARX1 I_40442 (I690040,I2507,I689706,I690066,);
nor I_40443 (I690074,I690066,I689933);
DFFARX1 I_40444 (I690074,I2507,I689706,I689674,);
nand I_40445 (I690105,I690066,I689975);
nand I_40446 (I689683,I689958,I690105);
not I_40447 (I690136,I690066);
nor I_40448 (I690153,I690136,I689876);
DFFARX1 I_40449 (I690153,I2507,I689706,I689695,);
nor I_40450 (I690184,I1226475,I1226466);
or I_40451 (I689686,I689933,I690184);
nor I_40452 (I689677,I690066,I690184);
or I_40453 (I689680,I689800,I690184);
DFFARX1 I_40454 (I690184,I2507,I689706,I689698,);
not I_40455 (I690284,I2514);
DFFARX1 I_40456 (I1035953,I2507,I690284,I690310,);
not I_40457 (I690318,I690310);
nand I_40458 (I690335,I1035950,I1035968);
and I_40459 (I690352,I690335,I1035965);
DFFARX1 I_40460 (I690352,I2507,I690284,I690378,);
not I_40461 (I690386,I1035947);
DFFARX1 I_40462 (I1035950,I2507,I690284,I690412,);
not I_40463 (I690420,I690412);
nor I_40464 (I690437,I690420,I690318);
and I_40465 (I690454,I690437,I1035947);
nor I_40466 (I690471,I690420,I690386);
nor I_40467 (I690267,I690378,I690471);
DFFARX1 I_40468 (I1035959,I2507,I690284,I690511,);
nor I_40469 (I690519,I690511,I690378);
not I_40470 (I690536,I690519);
not I_40471 (I690553,I690511);
nor I_40472 (I690570,I690553,I690454);
DFFARX1 I_40473 (I690570,I2507,I690284,I690270,);
nand I_40474 (I690601,I1035962,I1035947);
and I_40475 (I690618,I690601,I1035953);
DFFARX1 I_40476 (I690618,I2507,I690284,I690644,);
nor I_40477 (I690652,I690644,I690511);
DFFARX1 I_40478 (I690652,I2507,I690284,I690252,);
nand I_40479 (I690683,I690644,I690553);
nand I_40480 (I690261,I690536,I690683);
not I_40481 (I690714,I690644);
nor I_40482 (I690731,I690714,I690454);
DFFARX1 I_40483 (I690731,I2507,I690284,I690273,);
nor I_40484 (I690762,I1035956,I1035947);
or I_40485 (I690264,I690511,I690762);
nor I_40486 (I690255,I690644,I690762);
or I_40487 (I690258,I690378,I690762);
DFFARX1 I_40488 (I690762,I2507,I690284,I690276,);
not I_40489 (I690862,I2514);
DFFARX1 I_40490 (I941859,I2507,I690862,I690888,);
not I_40491 (I690896,I690888);
nand I_40492 (I690913,I941835,I941850);
and I_40493 (I690930,I690913,I941862);
DFFARX1 I_40494 (I690930,I2507,I690862,I690956,);
not I_40495 (I690964,I941847);
DFFARX1 I_40496 (I941838,I2507,I690862,I690990,);
not I_40497 (I690998,I690990);
nor I_40498 (I691015,I690998,I690896);
and I_40499 (I691032,I691015,I941847);
nor I_40500 (I691049,I690998,I690964);
nor I_40501 (I690845,I690956,I691049);
DFFARX1 I_40502 (I941835,I2507,I690862,I691089,);
nor I_40503 (I691097,I691089,I690956);
not I_40504 (I691114,I691097);
not I_40505 (I691131,I691089);
nor I_40506 (I691148,I691131,I691032);
DFFARX1 I_40507 (I691148,I2507,I690862,I690848,);
nand I_40508 (I691179,I941853,I941844);
and I_40509 (I691196,I691179,I941856);
DFFARX1 I_40510 (I691196,I2507,I690862,I691222,);
nor I_40511 (I691230,I691222,I691089);
DFFARX1 I_40512 (I691230,I2507,I690862,I690830,);
nand I_40513 (I691261,I691222,I691131);
nand I_40514 (I690839,I691114,I691261);
not I_40515 (I691292,I691222);
nor I_40516 (I691309,I691292,I691032);
DFFARX1 I_40517 (I691309,I2507,I690862,I690851,);
nor I_40518 (I691340,I941841,I941844);
or I_40519 (I690842,I691089,I691340);
nor I_40520 (I690833,I691222,I691340);
or I_40521 (I690836,I690956,I691340);
DFFARX1 I_40522 (I691340,I2507,I690862,I690854,);
not I_40523 (I691440,I2514);
DFFARX1 I_40524 (I576964,I2507,I691440,I691466,);
not I_40525 (I691474,I691466);
nand I_40526 (I691491,I576973,I576982);
and I_40527 (I691508,I691491,I576988);
DFFARX1 I_40528 (I691508,I2507,I691440,I691534,);
not I_40529 (I691542,I576985);
DFFARX1 I_40530 (I576970,I2507,I691440,I691568,);
not I_40531 (I691576,I691568);
nor I_40532 (I691593,I691576,I691474);
and I_40533 (I691610,I691593,I576985);
nor I_40534 (I691627,I691576,I691542);
nor I_40535 (I691423,I691534,I691627);
DFFARX1 I_40536 (I576979,I2507,I691440,I691667,);
nor I_40537 (I691675,I691667,I691534);
not I_40538 (I691692,I691675);
not I_40539 (I691709,I691667);
nor I_40540 (I691726,I691709,I691610);
DFFARX1 I_40541 (I691726,I2507,I691440,I691426,);
nand I_40542 (I691757,I576976,I576967);
and I_40543 (I691774,I691757,I576964);
DFFARX1 I_40544 (I691774,I2507,I691440,I691800,);
nor I_40545 (I691808,I691800,I691667);
DFFARX1 I_40546 (I691808,I2507,I691440,I691408,);
nand I_40547 (I691839,I691800,I691709);
nand I_40548 (I691417,I691692,I691839);
not I_40549 (I691870,I691800);
nor I_40550 (I691887,I691870,I691610);
DFFARX1 I_40551 (I691887,I2507,I691440,I691429,);
nor I_40552 (I691918,I576967,I576967);
or I_40553 (I691420,I691667,I691918);
nor I_40554 (I691411,I691800,I691918);
or I_40555 (I691414,I691534,I691918);
DFFARX1 I_40556 (I691918,I2507,I691440,I691432,);
not I_40557 (I692018,I2514);
DFFARX1 I_40558 (I111252,I2507,I692018,I692044,);
not I_40559 (I692052,I692044);
nand I_40560 (I692069,I111261,I111270);
and I_40561 (I692086,I692069,I111249);
DFFARX1 I_40562 (I692086,I2507,I692018,I692112,);
not I_40563 (I692120,I111252);
DFFARX1 I_40564 (I111267,I2507,I692018,I692146,);
not I_40565 (I692154,I692146);
nor I_40566 (I692171,I692154,I692052);
and I_40567 (I692188,I692171,I111252);
nor I_40568 (I692205,I692154,I692120);
nor I_40569 (I692001,I692112,I692205);
DFFARX1 I_40570 (I111258,I2507,I692018,I692245,);
nor I_40571 (I692253,I692245,I692112);
not I_40572 (I692270,I692253);
not I_40573 (I692287,I692245);
nor I_40574 (I692304,I692287,I692188);
DFFARX1 I_40575 (I692304,I2507,I692018,I692004,);
nand I_40576 (I692335,I111273,I111249);
and I_40577 (I692352,I692335,I111255);
DFFARX1 I_40578 (I692352,I2507,I692018,I692378,);
nor I_40579 (I692386,I692378,I692245);
DFFARX1 I_40580 (I692386,I2507,I692018,I691986,);
nand I_40581 (I692417,I692378,I692287);
nand I_40582 (I691995,I692270,I692417);
not I_40583 (I692448,I692378);
nor I_40584 (I692465,I692448,I692188);
DFFARX1 I_40585 (I692465,I2507,I692018,I692007,);
nor I_40586 (I692496,I111264,I111249);
or I_40587 (I691998,I692245,I692496);
nor I_40588 (I691989,I692378,I692496);
or I_40589 (I691992,I692112,I692496);
DFFARX1 I_40590 (I692496,I2507,I692018,I692010,);
not I_40591 (I692596,I2514);
DFFARX1 I_40592 (I1332114,I2507,I692596,I692622,);
not I_40593 (I692630,I692622);
nand I_40594 (I692647,I1332099,I1332087);
and I_40595 (I692664,I692647,I1332102);
DFFARX1 I_40596 (I692664,I2507,I692596,I692690,);
not I_40597 (I692698,I1332087);
DFFARX1 I_40598 (I1332105,I2507,I692596,I692724,);
not I_40599 (I692732,I692724);
nor I_40600 (I692749,I692732,I692630);
and I_40601 (I692766,I692749,I1332087);
nor I_40602 (I692783,I692732,I692698);
nor I_40603 (I692579,I692690,I692783);
DFFARX1 I_40604 (I1332093,I2507,I692596,I692823,);
nor I_40605 (I692831,I692823,I692690);
not I_40606 (I692848,I692831);
not I_40607 (I692865,I692823);
nor I_40608 (I692882,I692865,I692766);
DFFARX1 I_40609 (I692882,I2507,I692596,I692582,);
nand I_40610 (I692913,I1332090,I1332096);
and I_40611 (I692930,I692913,I1332111);
DFFARX1 I_40612 (I692930,I2507,I692596,I692956,);
nor I_40613 (I692964,I692956,I692823);
DFFARX1 I_40614 (I692964,I2507,I692596,I692564,);
nand I_40615 (I692995,I692956,I692865);
nand I_40616 (I692573,I692848,I692995);
not I_40617 (I693026,I692956);
nor I_40618 (I693043,I693026,I692766);
DFFARX1 I_40619 (I693043,I2507,I692596,I692585,);
nor I_40620 (I693074,I1332108,I1332096);
or I_40621 (I692576,I692823,I693074);
nor I_40622 (I692567,I692956,I693074);
or I_40623 (I692570,I692690,I693074);
DFFARX1 I_40624 (I693074,I2507,I692596,I692588,);
not I_40625 (I693174,I2514);
DFFARX1 I_40626 (I1058393,I2507,I693174,I693200,);
not I_40627 (I693208,I693200);
nand I_40628 (I693225,I1058390,I1058408);
and I_40629 (I693242,I693225,I1058405);
DFFARX1 I_40630 (I693242,I2507,I693174,I693268,);
not I_40631 (I693276,I1058387);
DFFARX1 I_40632 (I1058390,I2507,I693174,I693302,);
not I_40633 (I693310,I693302);
nor I_40634 (I693327,I693310,I693208);
and I_40635 (I693344,I693327,I1058387);
nor I_40636 (I693361,I693310,I693276);
nor I_40637 (I693157,I693268,I693361);
DFFARX1 I_40638 (I1058399,I2507,I693174,I693401,);
nor I_40639 (I693409,I693401,I693268);
not I_40640 (I693426,I693409);
not I_40641 (I693443,I693401);
nor I_40642 (I693460,I693443,I693344);
DFFARX1 I_40643 (I693460,I2507,I693174,I693160,);
nand I_40644 (I693491,I1058402,I1058387);
and I_40645 (I693508,I693491,I1058393);
DFFARX1 I_40646 (I693508,I2507,I693174,I693534,);
nor I_40647 (I693542,I693534,I693401);
DFFARX1 I_40648 (I693542,I2507,I693174,I693142,);
nand I_40649 (I693573,I693534,I693443);
nand I_40650 (I693151,I693426,I693573);
not I_40651 (I693604,I693534);
nor I_40652 (I693621,I693604,I693344);
DFFARX1 I_40653 (I693621,I2507,I693174,I693163,);
nor I_40654 (I693652,I1058396,I1058387);
or I_40655 (I693154,I693401,I693652);
nor I_40656 (I693145,I693534,I693652);
or I_40657 (I693148,I693268,I693652);
DFFARX1 I_40658 (I693652,I2507,I693174,I693166,);
not I_40659 (I693752,I2514);
DFFARX1 I_40660 (I215085,I2507,I693752,I693778,);
not I_40661 (I693786,I693778);
nand I_40662 (I693803,I215088,I215109);
and I_40663 (I693820,I693803,I215097);
DFFARX1 I_40664 (I693820,I2507,I693752,I693846,);
not I_40665 (I693854,I215094);
DFFARX1 I_40666 (I215085,I2507,I693752,I693880,);
not I_40667 (I693888,I693880);
nor I_40668 (I693905,I693888,I693786);
and I_40669 (I693922,I693905,I215094);
nor I_40670 (I693939,I693888,I693854);
nor I_40671 (I693735,I693846,I693939);
DFFARX1 I_40672 (I215103,I2507,I693752,I693979,);
nor I_40673 (I693987,I693979,I693846);
not I_40674 (I694004,I693987);
not I_40675 (I694021,I693979);
nor I_40676 (I694038,I694021,I693922);
DFFARX1 I_40677 (I694038,I2507,I693752,I693738,);
nand I_40678 (I694069,I215088,I215091);
and I_40679 (I694086,I694069,I215100);
DFFARX1 I_40680 (I694086,I2507,I693752,I694112,);
nor I_40681 (I694120,I694112,I693979);
DFFARX1 I_40682 (I694120,I2507,I693752,I693720,);
nand I_40683 (I694151,I694112,I694021);
nand I_40684 (I693729,I694004,I694151);
not I_40685 (I694182,I694112);
nor I_40686 (I694199,I694182,I693922);
DFFARX1 I_40687 (I694199,I2507,I693752,I693741,);
nor I_40688 (I694230,I215106,I215091);
or I_40689 (I693732,I693979,I694230);
nor I_40690 (I693723,I694112,I694230);
or I_40691 (I693726,I693846,I694230);
DFFARX1 I_40692 (I694230,I2507,I693752,I693744,);
not I_40693 (I694330,I2514);
DFFARX1 I_40694 (I826505,I2507,I694330,I694356,);
not I_40695 (I694364,I694356);
nand I_40696 (I694381,I826493,I826511);
and I_40697 (I694398,I694381,I826508);
DFFARX1 I_40698 (I694398,I2507,I694330,I694424,);
not I_40699 (I694432,I826499);
DFFARX1 I_40700 (I826496,I2507,I694330,I694458,);
not I_40701 (I694466,I694458);
nor I_40702 (I694483,I694466,I694364);
and I_40703 (I694500,I694483,I826499);
nor I_40704 (I694517,I694466,I694432);
nor I_40705 (I694313,I694424,I694517);
DFFARX1 I_40706 (I826490,I2507,I694330,I694557,);
nor I_40707 (I694565,I694557,I694424);
not I_40708 (I694582,I694565);
not I_40709 (I694599,I694557);
nor I_40710 (I694616,I694599,I694500);
DFFARX1 I_40711 (I694616,I2507,I694330,I694316,);
nand I_40712 (I694647,I826490,I826493);
and I_40713 (I694664,I694647,I826496);
DFFARX1 I_40714 (I694664,I2507,I694330,I694690,);
nor I_40715 (I694698,I694690,I694557);
DFFARX1 I_40716 (I694698,I2507,I694330,I694298,);
nand I_40717 (I694729,I694690,I694599);
nand I_40718 (I694307,I694582,I694729);
not I_40719 (I694760,I694690);
nor I_40720 (I694777,I694760,I694500);
DFFARX1 I_40721 (I694777,I2507,I694330,I694319,);
nor I_40722 (I694808,I826502,I826493);
or I_40723 (I694310,I694557,I694808);
nor I_40724 (I694301,I694690,I694808);
or I_40725 (I694304,I694424,I694808);
DFFARX1 I_40726 (I694808,I2507,I694330,I694322,);
not I_40727 (I694908,I2514);
DFFARX1 I_40728 (I224605,I2507,I694908,I694934,);
not I_40729 (I694942,I694934);
nand I_40730 (I694959,I224608,I224629);
and I_40731 (I694976,I694959,I224617);
DFFARX1 I_40732 (I694976,I2507,I694908,I695002,);
not I_40733 (I695010,I224614);
DFFARX1 I_40734 (I224605,I2507,I694908,I695036,);
not I_40735 (I695044,I695036);
nor I_40736 (I695061,I695044,I694942);
and I_40737 (I695078,I695061,I224614);
nor I_40738 (I695095,I695044,I695010);
nor I_40739 (I694891,I695002,I695095);
DFFARX1 I_40740 (I224623,I2507,I694908,I695135,);
nor I_40741 (I695143,I695135,I695002);
not I_40742 (I695160,I695143);
not I_40743 (I695177,I695135);
nor I_40744 (I695194,I695177,I695078);
DFFARX1 I_40745 (I695194,I2507,I694908,I694894,);
nand I_40746 (I695225,I224608,I224611);
and I_40747 (I695242,I695225,I224620);
DFFARX1 I_40748 (I695242,I2507,I694908,I695268,);
nor I_40749 (I695276,I695268,I695135);
DFFARX1 I_40750 (I695276,I2507,I694908,I694876,);
nand I_40751 (I695307,I695268,I695177);
nand I_40752 (I694885,I695160,I695307);
not I_40753 (I695338,I695268);
nor I_40754 (I695355,I695338,I695078);
DFFARX1 I_40755 (I695355,I2507,I694908,I694897,);
nor I_40756 (I695386,I224626,I224611);
or I_40757 (I694888,I695135,I695386);
nor I_40758 (I694879,I695268,I695386);
or I_40759 (I694882,I695002,I695386);
DFFARX1 I_40760 (I695386,I2507,I694908,I694900,);
not I_40761 (I695486,I2514);
DFFARX1 I_40762 (I936691,I2507,I695486,I695512,);
not I_40763 (I695520,I695512);
nand I_40764 (I695537,I936667,I936682);
and I_40765 (I695554,I695537,I936694);
DFFARX1 I_40766 (I695554,I2507,I695486,I695580,);
not I_40767 (I695588,I936679);
DFFARX1 I_40768 (I936670,I2507,I695486,I695614,);
not I_40769 (I695622,I695614);
nor I_40770 (I695639,I695622,I695520);
and I_40771 (I695656,I695639,I936679);
nor I_40772 (I695673,I695622,I695588);
nor I_40773 (I695469,I695580,I695673);
DFFARX1 I_40774 (I936667,I2507,I695486,I695713,);
nor I_40775 (I695721,I695713,I695580);
not I_40776 (I695738,I695721);
not I_40777 (I695755,I695713);
nor I_40778 (I695772,I695755,I695656);
DFFARX1 I_40779 (I695772,I2507,I695486,I695472,);
nand I_40780 (I695803,I936685,I936676);
and I_40781 (I695820,I695803,I936688);
DFFARX1 I_40782 (I695820,I2507,I695486,I695846,);
nor I_40783 (I695854,I695846,I695713);
DFFARX1 I_40784 (I695854,I2507,I695486,I695454,);
nand I_40785 (I695885,I695846,I695755);
nand I_40786 (I695463,I695738,I695885);
not I_40787 (I695916,I695846);
nor I_40788 (I695933,I695916,I695656);
DFFARX1 I_40789 (I695933,I2507,I695486,I695475,);
nor I_40790 (I695964,I936673,I936676);
or I_40791 (I695466,I695713,I695964);
nor I_40792 (I695457,I695846,I695964);
or I_40793 (I695460,I695580,I695964);
DFFARX1 I_40794 (I695964,I2507,I695486,I695478,);
not I_40795 (I696064,I2514);
DFFARX1 I_40796 (I1197108,I2507,I696064,I696090,);
not I_40797 (I696098,I696090);
nand I_40798 (I696115,I1197090,I1197102);
and I_40799 (I696132,I696115,I1197105);
DFFARX1 I_40800 (I696132,I2507,I696064,I696158,);
not I_40801 (I696166,I1197099);
DFFARX1 I_40802 (I1197096,I2507,I696064,I696192,);
not I_40803 (I696200,I696192);
nor I_40804 (I696217,I696200,I696098);
and I_40805 (I696234,I696217,I1197099);
nor I_40806 (I696251,I696200,I696166);
nor I_40807 (I696047,I696158,I696251);
DFFARX1 I_40808 (I1197114,I2507,I696064,I696291,);
nor I_40809 (I696299,I696291,I696158);
not I_40810 (I696316,I696299);
not I_40811 (I696333,I696291);
nor I_40812 (I696350,I696333,I696234);
DFFARX1 I_40813 (I696350,I2507,I696064,I696050,);
nand I_40814 (I696381,I1197093,I1197093);
and I_40815 (I696398,I696381,I1197090);
DFFARX1 I_40816 (I696398,I2507,I696064,I696424,);
nor I_40817 (I696432,I696424,I696291);
DFFARX1 I_40818 (I696432,I2507,I696064,I696032,);
nand I_40819 (I696463,I696424,I696333);
nand I_40820 (I696041,I696316,I696463);
not I_40821 (I696494,I696424);
nor I_40822 (I696511,I696494,I696234);
DFFARX1 I_40823 (I696511,I2507,I696064,I696053,);
nor I_40824 (I696542,I1197111,I1197093);
or I_40825 (I696044,I696291,I696542);
nor I_40826 (I696035,I696424,I696542);
or I_40827 (I696038,I696158,I696542);
DFFARX1 I_40828 (I696542,I2507,I696064,I696056,);
not I_40829 (I696642,I2514);
DFFARX1 I_40830 (I1105784,I2507,I696642,I696668,);
not I_40831 (I696676,I696668);
nand I_40832 (I696693,I1105766,I1105778);
and I_40833 (I696710,I696693,I1105781);
DFFARX1 I_40834 (I696710,I2507,I696642,I696736,);
not I_40835 (I696744,I1105775);
DFFARX1 I_40836 (I1105772,I2507,I696642,I696770,);
not I_40837 (I696778,I696770);
nor I_40838 (I696795,I696778,I696676);
and I_40839 (I696812,I696795,I1105775);
nor I_40840 (I696829,I696778,I696744);
nor I_40841 (I696625,I696736,I696829);
DFFARX1 I_40842 (I1105790,I2507,I696642,I696869,);
nor I_40843 (I696877,I696869,I696736);
not I_40844 (I696894,I696877);
not I_40845 (I696911,I696869);
nor I_40846 (I696928,I696911,I696812);
DFFARX1 I_40847 (I696928,I2507,I696642,I696628,);
nand I_40848 (I696959,I1105769,I1105769);
and I_40849 (I696976,I696959,I1105766);
DFFARX1 I_40850 (I696976,I2507,I696642,I697002,);
nor I_40851 (I697010,I697002,I696869);
DFFARX1 I_40852 (I697010,I2507,I696642,I696610,);
nand I_40853 (I697041,I697002,I696911);
nand I_40854 (I696619,I696894,I697041);
not I_40855 (I697072,I697002);
nor I_40856 (I697089,I697072,I696812);
DFFARX1 I_40857 (I697089,I2507,I696642,I696631,);
nor I_40858 (I697120,I1105787,I1105769);
or I_40859 (I696622,I696869,I697120);
nor I_40860 (I696613,I697002,I697120);
or I_40861 (I696616,I696736,I697120);
DFFARX1 I_40862 (I697120,I2507,I696642,I696634,);
not I_40863 (I697220,I2514);
DFFARX1 I_40864 (I24833,I2507,I697220,I697246,);
not I_40865 (I697254,I697246);
nand I_40866 (I697271,I24830,I24821);
and I_40867 (I697288,I697271,I24821);
DFFARX1 I_40868 (I697288,I2507,I697220,I697314,);
not I_40869 (I697322,I24824);
DFFARX1 I_40870 (I24839,I2507,I697220,I697348,);
not I_40871 (I697356,I697348);
nor I_40872 (I697373,I697356,I697254);
and I_40873 (I697390,I697373,I24824);
nor I_40874 (I697407,I697356,I697322);
nor I_40875 (I697203,I697314,I697407);
DFFARX1 I_40876 (I24824,I2507,I697220,I697447,);
nor I_40877 (I697455,I697447,I697314);
not I_40878 (I697472,I697455);
not I_40879 (I697489,I697447);
nor I_40880 (I697506,I697489,I697390);
DFFARX1 I_40881 (I697506,I2507,I697220,I697206,);
nand I_40882 (I697537,I24842,I24827);
and I_40883 (I697554,I697537,I24845);
DFFARX1 I_40884 (I697554,I2507,I697220,I697580,);
nor I_40885 (I697588,I697580,I697447);
DFFARX1 I_40886 (I697588,I2507,I697220,I697188,);
nand I_40887 (I697619,I697580,I697489);
nand I_40888 (I697197,I697472,I697619);
not I_40889 (I697650,I697580);
nor I_40890 (I697667,I697650,I697390);
DFFARX1 I_40891 (I697667,I2507,I697220,I697209,);
nor I_40892 (I697698,I24836,I24827);
or I_40893 (I697200,I697447,I697698);
nor I_40894 (I697191,I697580,I697698);
or I_40895 (I697194,I697314,I697698);
DFFARX1 I_40896 (I697698,I2507,I697220,I697212,);
not I_40897 (I697798,I2514);
DFFARX1 I_40898 (I1207426,I2507,I697798,I697824,);
not I_40899 (I697832,I697824);
nand I_40900 (I697849,I1207429,I1207438);
and I_40901 (I697866,I697849,I1207441);
DFFARX1 I_40902 (I697866,I2507,I697798,I697892,);
not I_40903 (I697900,I1207450);
DFFARX1 I_40904 (I1207432,I2507,I697798,I697926,);
not I_40905 (I697934,I697926);
nor I_40906 (I697951,I697934,I697832);
and I_40907 (I697968,I697951,I1207450);
nor I_40908 (I697985,I697934,I697900);
nor I_40909 (I697781,I697892,I697985);
DFFARX1 I_40910 (I1207429,I2507,I697798,I698025,);
nor I_40911 (I698033,I698025,I697892);
not I_40912 (I698050,I698033);
not I_40913 (I698067,I698025);
nor I_40914 (I698084,I698067,I697968);
DFFARX1 I_40915 (I698084,I2507,I697798,I697784,);
nand I_40916 (I698115,I1207447,I1207426);
and I_40917 (I698132,I698115,I1207444);
DFFARX1 I_40918 (I698132,I2507,I697798,I698158,);
nor I_40919 (I698166,I698158,I698025);
DFFARX1 I_40920 (I698166,I2507,I697798,I697766,);
nand I_40921 (I698197,I698158,I698067);
nand I_40922 (I697775,I698050,I698197);
not I_40923 (I698228,I698158);
nor I_40924 (I698245,I698228,I697968);
DFFARX1 I_40925 (I698245,I2507,I697798,I697787,);
nor I_40926 (I698276,I1207435,I1207426);
or I_40927 (I697778,I698025,I698276);
nor I_40928 (I697769,I698158,I698276);
or I_40929 (I697772,I697892,I698276);
DFFARX1 I_40930 (I698276,I2507,I697798,I697790,);
not I_40931 (I698376,I2514);
DFFARX1 I_40932 (I1041002,I2507,I698376,I698402,);
not I_40933 (I698410,I698402);
nand I_40934 (I698427,I1040999,I1041017);
and I_40935 (I698444,I698427,I1041014);
DFFARX1 I_40936 (I698444,I2507,I698376,I698470,);
not I_40937 (I698478,I1040996);
DFFARX1 I_40938 (I1040999,I2507,I698376,I698504,);
not I_40939 (I698512,I698504);
nor I_40940 (I698529,I698512,I698410);
and I_40941 (I698546,I698529,I1040996);
nor I_40942 (I698563,I698512,I698478);
nor I_40943 (I698359,I698470,I698563);
DFFARX1 I_40944 (I1041008,I2507,I698376,I698603,);
nor I_40945 (I698611,I698603,I698470);
not I_40946 (I698628,I698611);
not I_40947 (I698645,I698603);
nor I_40948 (I698662,I698645,I698546);
DFFARX1 I_40949 (I698662,I2507,I698376,I698362,);
nand I_40950 (I698693,I1041011,I1040996);
and I_40951 (I698710,I698693,I1041002);
DFFARX1 I_40952 (I698710,I2507,I698376,I698736,);
nor I_40953 (I698744,I698736,I698603);
DFFARX1 I_40954 (I698744,I2507,I698376,I698344,);
nand I_40955 (I698775,I698736,I698645);
nand I_40956 (I698353,I698628,I698775);
not I_40957 (I698806,I698736);
nor I_40958 (I698823,I698806,I698546);
DFFARX1 I_40959 (I698823,I2507,I698376,I698365,);
nor I_40960 (I698854,I1041005,I1040996);
or I_40961 (I698356,I698603,I698854);
nor I_40962 (I698347,I698736,I698854);
or I_40963 (I698350,I698470,I698854);
DFFARX1 I_40964 (I698854,I2507,I698376,I698368,);
not I_40965 (I698954,I2514);
DFFARX1 I_40966 (I334007,I2507,I698954,I698980,);
not I_40967 (I698988,I698980);
nand I_40968 (I699005,I334010,I333986);
and I_40969 (I699022,I699005,I333983);
DFFARX1 I_40970 (I699022,I2507,I698954,I699048,);
not I_40971 (I699056,I333989);
DFFARX1 I_40972 (I333983,I2507,I698954,I699082,);
not I_40973 (I699090,I699082);
nor I_40974 (I699107,I699090,I698988);
and I_40975 (I699124,I699107,I333989);
nor I_40976 (I699141,I699090,I699056);
nor I_40977 (I698937,I699048,I699141);
DFFARX1 I_40978 (I333992,I2507,I698954,I699181,);
nor I_40979 (I699189,I699181,I699048);
not I_40980 (I699206,I699189);
not I_40981 (I699223,I699181);
nor I_40982 (I699240,I699223,I699124);
DFFARX1 I_40983 (I699240,I2507,I698954,I698940,);
nand I_40984 (I699271,I333995,I334004);
and I_40985 (I699288,I699271,I334001);
DFFARX1 I_40986 (I699288,I2507,I698954,I699314,);
nor I_40987 (I699322,I699314,I699181);
DFFARX1 I_40988 (I699322,I2507,I698954,I698922,);
nand I_40989 (I699353,I699314,I699223);
nand I_40990 (I698931,I699206,I699353);
not I_40991 (I699384,I699314);
nor I_40992 (I699401,I699384,I699124);
DFFARX1 I_40993 (I699401,I2507,I698954,I698943,);
nor I_40994 (I699432,I333998,I334004);
or I_40995 (I698934,I699181,I699432);
nor I_40996 (I698925,I699314,I699432);
or I_40997 (I698928,I699048,I699432);
DFFARX1 I_40998 (I699432,I2507,I698954,I698946,);
not I_40999 (I699532,I2514);
DFFARX1 I_41000 (I999353,I2507,I699532,I699558,);
not I_41001 (I699566,I699558);
nand I_41002 (I699583,I999329,I999344);
and I_41003 (I699600,I699583,I999356);
DFFARX1 I_41004 (I699600,I2507,I699532,I699626,);
not I_41005 (I699634,I999341);
DFFARX1 I_41006 (I999332,I2507,I699532,I699660,);
not I_41007 (I699668,I699660);
nor I_41008 (I699685,I699668,I699566);
and I_41009 (I699702,I699685,I999341);
nor I_41010 (I699719,I699668,I699634);
nor I_41011 (I699515,I699626,I699719);
DFFARX1 I_41012 (I999329,I2507,I699532,I699759,);
nor I_41013 (I699767,I699759,I699626);
not I_41014 (I699784,I699767);
not I_41015 (I699801,I699759);
nor I_41016 (I699818,I699801,I699702);
DFFARX1 I_41017 (I699818,I2507,I699532,I699518,);
nand I_41018 (I699849,I999347,I999338);
and I_41019 (I699866,I699849,I999350);
DFFARX1 I_41020 (I699866,I2507,I699532,I699892,);
nor I_41021 (I699900,I699892,I699759);
DFFARX1 I_41022 (I699900,I2507,I699532,I699500,);
nand I_41023 (I699931,I699892,I699801);
nand I_41024 (I699509,I699784,I699931);
not I_41025 (I699962,I699892);
nor I_41026 (I699979,I699962,I699702);
DFFARX1 I_41027 (I699979,I2507,I699532,I699521,);
nor I_41028 (I700010,I999335,I999338);
or I_41029 (I699512,I699759,I700010);
nor I_41030 (I699503,I699892,I700010);
or I_41031 (I699506,I699626,I700010);
DFFARX1 I_41032 (I700010,I2507,I699532,I699524,);
not I_41033 (I700110,I2514);
DFFARX1 I_41034 (I492568,I2507,I700110,I700136,);
not I_41035 (I700144,I700136);
nand I_41036 (I700161,I492559,I492577);
and I_41037 (I700178,I700161,I492580);
DFFARX1 I_41038 (I700178,I2507,I700110,I700204,);
not I_41039 (I700212,I492574);
DFFARX1 I_41040 (I492562,I2507,I700110,I700238,);
not I_41041 (I700246,I700238);
nor I_41042 (I700263,I700246,I700144);
and I_41043 (I700280,I700263,I492574);
nor I_41044 (I700297,I700246,I700212);
nor I_41045 (I700093,I700204,I700297);
DFFARX1 I_41046 (I492571,I2507,I700110,I700337,);
nor I_41047 (I700345,I700337,I700204);
not I_41048 (I700362,I700345);
not I_41049 (I700379,I700337);
nor I_41050 (I700396,I700379,I700280);
DFFARX1 I_41051 (I700396,I2507,I700110,I700096,);
nand I_41052 (I700427,I492586,I492583);
and I_41053 (I700444,I700427,I492565);
DFFARX1 I_41054 (I700444,I2507,I700110,I700470,);
nor I_41055 (I700478,I700470,I700337);
DFFARX1 I_41056 (I700478,I2507,I700110,I700078,);
nand I_41057 (I700509,I700470,I700379);
nand I_41058 (I700087,I700362,I700509);
not I_41059 (I700540,I700470);
nor I_41060 (I700557,I700540,I700280);
DFFARX1 I_41061 (I700557,I2507,I700110,I700099,);
nor I_41062 (I700588,I492559,I492583);
or I_41063 (I700090,I700337,I700588);
nor I_41064 (I700081,I700470,I700588);
or I_41065 (I700084,I700204,I700588);
DFFARX1 I_41066 (I700588,I2507,I700110,I700102,);
not I_41067 (I700688,I2514);
DFFARX1 I_41068 (I511939,I2507,I700688,I700714,);
not I_41069 (I700722,I700714);
nand I_41070 (I700739,I511954,I511939);
and I_41071 (I700756,I700739,I511942);
DFFARX1 I_41072 (I700756,I2507,I700688,I700782,);
not I_41073 (I700790,I511942);
DFFARX1 I_41074 (I511951,I2507,I700688,I700816,);
not I_41075 (I700824,I700816);
nor I_41076 (I700841,I700824,I700722);
and I_41077 (I700858,I700841,I511942);
nor I_41078 (I700875,I700824,I700790);
nor I_41079 (I700671,I700782,I700875);
DFFARX1 I_41080 (I511945,I2507,I700688,I700915,);
nor I_41081 (I700923,I700915,I700782);
not I_41082 (I700940,I700923);
not I_41083 (I700957,I700915);
nor I_41084 (I700974,I700957,I700858);
DFFARX1 I_41085 (I700974,I2507,I700688,I700674,);
nand I_41086 (I701005,I511948,I511957);
and I_41087 (I701022,I701005,I511963);
DFFARX1 I_41088 (I701022,I2507,I700688,I701048,);
nor I_41089 (I701056,I701048,I700915);
DFFARX1 I_41090 (I701056,I2507,I700688,I700656,);
nand I_41091 (I701087,I701048,I700957);
nand I_41092 (I700665,I700940,I701087);
not I_41093 (I701118,I701048);
nor I_41094 (I701135,I701118,I700858);
DFFARX1 I_41095 (I701135,I2507,I700688,I700677,);
nor I_41096 (I701166,I511960,I511957);
or I_41097 (I700668,I700915,I701166);
nor I_41098 (I700659,I701048,I701166);
or I_41099 (I700662,I700782,I701166);
DFFARX1 I_41100 (I701166,I2507,I700688,I700680,);
not I_41101 (I701266,I2514);
DFFARX1 I_41102 (I1358889,I2507,I701266,I701292,);
not I_41103 (I701300,I701292);
nand I_41104 (I701317,I1358874,I1358862);
and I_41105 (I701334,I701317,I1358877);
DFFARX1 I_41106 (I701334,I2507,I701266,I701360,);
not I_41107 (I701368,I1358862);
DFFARX1 I_41108 (I1358880,I2507,I701266,I701394,);
not I_41109 (I701402,I701394);
nor I_41110 (I701419,I701402,I701300);
and I_41111 (I701436,I701419,I1358862);
nor I_41112 (I701453,I701402,I701368);
nor I_41113 (I701249,I701360,I701453);
DFFARX1 I_41114 (I1358868,I2507,I701266,I701493,);
nor I_41115 (I701501,I701493,I701360);
not I_41116 (I701518,I701501);
not I_41117 (I701535,I701493);
nor I_41118 (I701552,I701535,I701436);
DFFARX1 I_41119 (I701552,I2507,I701266,I701252,);
nand I_41120 (I701583,I1358865,I1358871);
and I_41121 (I701600,I701583,I1358886);
DFFARX1 I_41122 (I701600,I2507,I701266,I701626,);
nor I_41123 (I701634,I701626,I701493);
DFFARX1 I_41124 (I701634,I2507,I701266,I701234,);
nand I_41125 (I701665,I701626,I701535);
nand I_41126 (I701243,I701518,I701665);
not I_41127 (I701696,I701626);
nor I_41128 (I701713,I701696,I701436);
DFFARX1 I_41129 (I701713,I2507,I701266,I701255,);
nor I_41130 (I701744,I1358883,I1358871);
or I_41131 (I701246,I701493,I701744);
nor I_41132 (I701237,I701626,I701744);
or I_41133 (I701240,I701360,I701744);
DFFARX1 I_41134 (I701744,I2507,I701266,I701258,);
not I_41135 (I701844,I2514);
DFFARX1 I_41136 (I406072,I2507,I701844,I701870,);
not I_41137 (I701878,I701870);
nand I_41138 (I701895,I406063,I406081);
and I_41139 (I701912,I701895,I406084);
DFFARX1 I_41140 (I701912,I2507,I701844,I701938,);
not I_41141 (I701946,I406078);
DFFARX1 I_41142 (I406066,I2507,I701844,I701972,);
not I_41143 (I701980,I701972);
nor I_41144 (I701997,I701980,I701878);
and I_41145 (I702014,I701997,I406078);
nor I_41146 (I702031,I701980,I701946);
nor I_41147 (I701827,I701938,I702031);
DFFARX1 I_41148 (I406075,I2507,I701844,I702071,);
nor I_41149 (I702079,I702071,I701938);
not I_41150 (I702096,I702079);
not I_41151 (I702113,I702071);
nor I_41152 (I702130,I702113,I702014);
DFFARX1 I_41153 (I702130,I2507,I701844,I701830,);
nand I_41154 (I702161,I406090,I406087);
and I_41155 (I702178,I702161,I406069);
DFFARX1 I_41156 (I702178,I2507,I701844,I702204,);
nor I_41157 (I702212,I702204,I702071);
DFFARX1 I_41158 (I702212,I2507,I701844,I701812,);
nand I_41159 (I702243,I702204,I702113);
nand I_41160 (I701821,I702096,I702243);
not I_41161 (I702274,I702204);
nor I_41162 (I702291,I702274,I702014);
DFFARX1 I_41163 (I702291,I2507,I701844,I701833,);
nor I_41164 (I702322,I406063,I406087);
or I_41165 (I701824,I702071,I702322);
nor I_41166 (I701815,I702204,I702322);
or I_41167 (I701818,I701938,I702322);
DFFARX1 I_41168 (I702322,I2507,I701844,I701836,);
not I_41169 (I702422,I2514);
DFFARX1 I_41170 (I781183,I2507,I702422,I702448,);
not I_41171 (I702456,I702448);
nand I_41172 (I702473,I781171,I781189);
and I_41173 (I702490,I702473,I781186);
DFFARX1 I_41174 (I702490,I2507,I702422,I702516,);
not I_41175 (I702524,I781177);
DFFARX1 I_41176 (I781174,I2507,I702422,I702550,);
not I_41177 (I702558,I702550);
nor I_41178 (I702575,I702558,I702456);
and I_41179 (I702592,I702575,I781177);
nor I_41180 (I702609,I702558,I702524);
nor I_41181 (I702405,I702516,I702609);
DFFARX1 I_41182 (I781168,I2507,I702422,I702649,);
nor I_41183 (I702657,I702649,I702516);
not I_41184 (I702674,I702657);
not I_41185 (I702691,I702649);
nor I_41186 (I702708,I702691,I702592);
DFFARX1 I_41187 (I702708,I2507,I702422,I702408,);
nand I_41188 (I702739,I781168,I781171);
and I_41189 (I702756,I702739,I781174);
DFFARX1 I_41190 (I702756,I2507,I702422,I702782,);
nor I_41191 (I702790,I702782,I702649);
DFFARX1 I_41192 (I702790,I2507,I702422,I702390,);
nand I_41193 (I702821,I702782,I702691);
nand I_41194 (I702399,I702674,I702821);
not I_41195 (I702852,I702782);
nor I_41196 (I702869,I702852,I702592);
DFFARX1 I_41197 (I702869,I2507,I702422,I702411,);
nor I_41198 (I702900,I781180,I781171);
or I_41199 (I702402,I702649,I702900);
nor I_41200 (I702393,I702782,I702900);
or I_41201 (I702396,I702516,I702900);
DFFARX1 I_41202 (I702900,I2507,I702422,I702414,);
not I_41203 (I703000,I2514);
DFFARX1 I_41204 (I618002,I2507,I703000,I703026,);
not I_41205 (I703034,I703026);
nand I_41206 (I703051,I618011,I618020);
and I_41207 (I703068,I703051,I618026);
DFFARX1 I_41208 (I703068,I2507,I703000,I703094,);
not I_41209 (I703102,I618023);
DFFARX1 I_41210 (I618008,I2507,I703000,I703128,);
not I_41211 (I703136,I703128);
nor I_41212 (I703153,I703136,I703034);
and I_41213 (I703170,I703153,I618023);
nor I_41214 (I703187,I703136,I703102);
nor I_41215 (I702983,I703094,I703187);
DFFARX1 I_41216 (I618017,I2507,I703000,I703227,);
nor I_41217 (I703235,I703227,I703094);
not I_41218 (I703252,I703235);
not I_41219 (I703269,I703227);
nor I_41220 (I703286,I703269,I703170);
DFFARX1 I_41221 (I703286,I2507,I703000,I702986,);
nand I_41222 (I703317,I618014,I618005);
and I_41223 (I703334,I703317,I618002);
DFFARX1 I_41224 (I703334,I2507,I703000,I703360,);
nor I_41225 (I703368,I703360,I703227);
DFFARX1 I_41226 (I703368,I2507,I703000,I702968,);
nand I_41227 (I703399,I703360,I703269);
nand I_41228 (I702977,I703252,I703399);
not I_41229 (I703430,I703360);
nor I_41230 (I703447,I703430,I703170);
DFFARX1 I_41231 (I703447,I2507,I703000,I702989,);
nor I_41232 (I703478,I618005,I618005);
or I_41233 (I702980,I703227,I703478);
nor I_41234 (I702971,I703360,I703478);
or I_41235 (I702974,I703094,I703478);
DFFARX1 I_41236 (I703478,I2507,I703000,I702992,);
not I_41237 (I703578,I2514);
DFFARX1 I_41238 (I786980,I2507,I703578,I703604,);
not I_41239 (I703612,I703604);
nand I_41240 (I703629,I786968,I786986);
and I_41241 (I703646,I703629,I786983);
DFFARX1 I_41242 (I703646,I2507,I703578,I703672,);
not I_41243 (I703680,I786974);
DFFARX1 I_41244 (I786971,I2507,I703578,I703706,);
not I_41245 (I703714,I703706);
nor I_41246 (I703731,I703714,I703612);
and I_41247 (I703748,I703731,I786974);
nor I_41248 (I703765,I703714,I703680);
nor I_41249 (I703561,I703672,I703765);
DFFARX1 I_41250 (I786965,I2507,I703578,I703805,);
nor I_41251 (I703813,I703805,I703672);
not I_41252 (I703830,I703813);
not I_41253 (I703847,I703805);
nor I_41254 (I703864,I703847,I703748);
DFFARX1 I_41255 (I703864,I2507,I703578,I703564,);
nand I_41256 (I703895,I786965,I786968);
and I_41257 (I703912,I703895,I786971);
DFFARX1 I_41258 (I703912,I2507,I703578,I703938,);
nor I_41259 (I703946,I703938,I703805);
DFFARX1 I_41260 (I703946,I2507,I703578,I703546,);
nand I_41261 (I703977,I703938,I703847);
nand I_41262 (I703555,I703830,I703977);
not I_41263 (I704008,I703938);
nor I_41264 (I704025,I704008,I703748);
DFFARX1 I_41265 (I704025,I2507,I703578,I703567,);
nor I_41266 (I704056,I786977,I786968);
or I_41267 (I703558,I703805,I704056);
nor I_41268 (I703549,I703938,I704056);
or I_41269 (I703552,I703672,I704056);
DFFARX1 I_41270 (I704056,I2507,I703578,I703570,);
not I_41271 (I704156,I2514);
DFFARX1 I_41272 (I412600,I2507,I704156,I704182,);
not I_41273 (I704190,I704182);
nand I_41274 (I704207,I412591,I412609);
and I_41275 (I704224,I704207,I412612);
DFFARX1 I_41276 (I704224,I2507,I704156,I704250,);
not I_41277 (I704258,I412606);
DFFARX1 I_41278 (I412594,I2507,I704156,I704284,);
not I_41279 (I704292,I704284);
nor I_41280 (I704309,I704292,I704190);
and I_41281 (I704326,I704309,I412606);
nor I_41282 (I704343,I704292,I704258);
nor I_41283 (I704139,I704250,I704343);
DFFARX1 I_41284 (I412603,I2507,I704156,I704383,);
nor I_41285 (I704391,I704383,I704250);
not I_41286 (I704408,I704391);
not I_41287 (I704425,I704383);
nor I_41288 (I704442,I704425,I704326);
DFFARX1 I_41289 (I704442,I2507,I704156,I704142,);
nand I_41290 (I704473,I412618,I412615);
and I_41291 (I704490,I704473,I412597);
DFFARX1 I_41292 (I704490,I2507,I704156,I704516,);
nor I_41293 (I704524,I704516,I704383);
DFFARX1 I_41294 (I704524,I2507,I704156,I704124,);
nand I_41295 (I704555,I704516,I704425);
nand I_41296 (I704133,I704408,I704555);
not I_41297 (I704586,I704516);
nor I_41298 (I704603,I704586,I704326);
DFFARX1 I_41299 (I704603,I2507,I704156,I704145,);
nor I_41300 (I704634,I412591,I412615);
or I_41301 (I704136,I704383,I704634);
nor I_41302 (I704127,I704516,I704634);
or I_41303 (I704130,I704250,I704634);
DFFARX1 I_41304 (I704634,I2507,I704156,I704148,);
not I_41305 (I704734,I2514);
DFFARX1 I_41306 (I80159,I2507,I704734,I704760,);
not I_41307 (I704768,I704760);
nand I_41308 (I704785,I80168,I80177);
and I_41309 (I704802,I704785,I80156);
DFFARX1 I_41310 (I704802,I2507,I704734,I704828,);
not I_41311 (I704836,I80159);
DFFARX1 I_41312 (I80174,I2507,I704734,I704862,);
not I_41313 (I704870,I704862);
nor I_41314 (I704887,I704870,I704768);
and I_41315 (I704904,I704887,I80159);
nor I_41316 (I704921,I704870,I704836);
nor I_41317 (I704717,I704828,I704921);
DFFARX1 I_41318 (I80165,I2507,I704734,I704961,);
nor I_41319 (I704969,I704961,I704828);
not I_41320 (I704986,I704969);
not I_41321 (I705003,I704961);
nor I_41322 (I705020,I705003,I704904);
DFFARX1 I_41323 (I705020,I2507,I704734,I704720,);
nand I_41324 (I705051,I80180,I80156);
and I_41325 (I705068,I705051,I80162);
DFFARX1 I_41326 (I705068,I2507,I704734,I705094,);
nor I_41327 (I705102,I705094,I704961);
DFFARX1 I_41328 (I705102,I2507,I704734,I704702,);
nand I_41329 (I705133,I705094,I705003);
nand I_41330 (I704711,I704986,I705133);
not I_41331 (I705164,I705094);
nor I_41332 (I705181,I705164,I704904);
DFFARX1 I_41333 (I705181,I2507,I704734,I704723,);
nor I_41334 (I705212,I80171,I80156);
or I_41335 (I704714,I704961,I705212);
nor I_41336 (I704705,I705094,I705212);
or I_41337 (I704708,I704828,I705212);
DFFARX1 I_41338 (I705212,I2507,I704734,I704726,);
not I_41339 (I705312,I2514);
DFFARX1 I_41340 (I1320809,I2507,I705312,I705338,);
not I_41341 (I705346,I705338);
nand I_41342 (I705363,I1320794,I1320782);
and I_41343 (I705380,I705363,I1320797);
DFFARX1 I_41344 (I705380,I2507,I705312,I705406,);
not I_41345 (I705414,I1320782);
DFFARX1 I_41346 (I1320800,I2507,I705312,I705440,);
not I_41347 (I705448,I705440);
nor I_41348 (I705465,I705448,I705346);
and I_41349 (I705482,I705465,I1320782);
nor I_41350 (I705499,I705448,I705414);
nor I_41351 (I705295,I705406,I705499);
DFFARX1 I_41352 (I1320788,I2507,I705312,I705539,);
nor I_41353 (I705547,I705539,I705406);
not I_41354 (I705564,I705547);
not I_41355 (I705581,I705539);
nor I_41356 (I705598,I705581,I705482);
DFFARX1 I_41357 (I705598,I2507,I705312,I705298,);
nand I_41358 (I705629,I1320785,I1320791);
and I_41359 (I705646,I705629,I1320806);
DFFARX1 I_41360 (I705646,I2507,I705312,I705672,);
nor I_41361 (I705680,I705672,I705539);
DFFARX1 I_41362 (I705680,I2507,I705312,I705280,);
nand I_41363 (I705711,I705672,I705581);
nand I_41364 (I705289,I705564,I705711);
not I_41365 (I705742,I705672);
nor I_41366 (I705759,I705742,I705482);
DFFARX1 I_41367 (I705759,I2507,I705312,I705301,);
nor I_41368 (I705790,I1320803,I1320791);
or I_41369 (I705292,I705539,I705790);
nor I_41370 (I705283,I705672,I705790);
or I_41371 (I705286,I705406,I705790);
DFFARX1 I_41372 (I705790,I2507,I705312,I705304,);
not I_41373 (I705890,I2514);
DFFARX1 I_41374 (I25887,I2507,I705890,I705916,);
not I_41375 (I705924,I705916);
nand I_41376 (I705941,I25884,I25875);
and I_41377 (I705958,I705941,I25875);
DFFARX1 I_41378 (I705958,I2507,I705890,I705984,);
not I_41379 (I705992,I25878);
DFFARX1 I_41380 (I25893,I2507,I705890,I706018,);
not I_41381 (I706026,I706018);
nor I_41382 (I706043,I706026,I705924);
and I_41383 (I706060,I706043,I25878);
nor I_41384 (I706077,I706026,I705992);
nor I_41385 (I705873,I705984,I706077);
DFFARX1 I_41386 (I25878,I2507,I705890,I706117,);
nor I_41387 (I706125,I706117,I705984);
not I_41388 (I706142,I706125);
not I_41389 (I706159,I706117);
nor I_41390 (I706176,I706159,I706060);
DFFARX1 I_41391 (I706176,I2507,I705890,I705876,);
nand I_41392 (I706207,I25896,I25881);
and I_41393 (I706224,I706207,I25899);
DFFARX1 I_41394 (I706224,I2507,I705890,I706250,);
nor I_41395 (I706258,I706250,I706117);
DFFARX1 I_41396 (I706258,I2507,I705890,I705858,);
nand I_41397 (I706289,I706250,I706159);
nand I_41398 (I705867,I706142,I706289);
not I_41399 (I706320,I706250);
nor I_41400 (I706337,I706320,I706060);
DFFARX1 I_41401 (I706337,I2507,I705890,I705879,);
nor I_41402 (I706368,I25890,I25881);
or I_41403 (I705870,I706117,I706368);
nor I_41404 (I705861,I706250,I706368);
or I_41405 (I705864,I705984,I706368);
DFFARX1 I_41406 (I706368,I2507,I705890,I705882,);
not I_41407 (I706468,I2514);
DFFARX1 I_41408 (I319778,I2507,I706468,I706494,);
not I_41409 (I706502,I706494);
nand I_41410 (I706519,I319781,I319757);
and I_41411 (I706536,I706519,I319754);
DFFARX1 I_41412 (I706536,I2507,I706468,I706562,);
not I_41413 (I706570,I319760);
DFFARX1 I_41414 (I319754,I2507,I706468,I706596,);
not I_41415 (I706604,I706596);
nor I_41416 (I706621,I706604,I706502);
and I_41417 (I706638,I706621,I319760);
nor I_41418 (I706655,I706604,I706570);
nor I_41419 (I706451,I706562,I706655);
DFFARX1 I_41420 (I319763,I2507,I706468,I706695,);
nor I_41421 (I706703,I706695,I706562);
not I_41422 (I706720,I706703);
not I_41423 (I706737,I706695);
nor I_41424 (I706754,I706737,I706638);
DFFARX1 I_41425 (I706754,I2507,I706468,I706454,);
nand I_41426 (I706785,I319766,I319775);
and I_41427 (I706802,I706785,I319772);
DFFARX1 I_41428 (I706802,I2507,I706468,I706828,);
nor I_41429 (I706836,I706828,I706695);
DFFARX1 I_41430 (I706836,I2507,I706468,I706436,);
nand I_41431 (I706867,I706828,I706737);
nand I_41432 (I706445,I706720,I706867);
not I_41433 (I706898,I706828);
nor I_41434 (I706915,I706898,I706638);
DFFARX1 I_41435 (I706915,I2507,I706468,I706457,);
nor I_41436 (I706946,I319769,I319775);
or I_41437 (I706448,I706695,I706946);
nor I_41438 (I706439,I706828,I706946);
or I_41439 (I706442,I706562,I706946);
DFFARX1 I_41440 (I706946,I2507,I706468,I706460,);
not I_41441 (I707046,I2514);
DFFARX1 I_41442 (I1188438,I2507,I707046,I707072,);
not I_41443 (I707080,I707072);
nand I_41444 (I707097,I1188420,I1188432);
and I_41445 (I707114,I707097,I1188435);
DFFARX1 I_41446 (I707114,I2507,I707046,I707140,);
not I_41447 (I707148,I1188429);
DFFARX1 I_41448 (I1188426,I2507,I707046,I707174,);
not I_41449 (I707182,I707174);
nor I_41450 (I707199,I707182,I707080);
and I_41451 (I707216,I707199,I1188429);
nor I_41452 (I707233,I707182,I707148);
nor I_41453 (I707029,I707140,I707233);
DFFARX1 I_41454 (I1188444,I2507,I707046,I707273,);
nor I_41455 (I707281,I707273,I707140);
not I_41456 (I707298,I707281);
not I_41457 (I707315,I707273);
nor I_41458 (I707332,I707315,I707216);
DFFARX1 I_41459 (I707332,I2507,I707046,I707032,);
nand I_41460 (I707363,I1188423,I1188423);
and I_41461 (I707380,I707363,I1188420);
DFFARX1 I_41462 (I707380,I2507,I707046,I707406,);
nor I_41463 (I707414,I707406,I707273);
DFFARX1 I_41464 (I707414,I2507,I707046,I707014,);
nand I_41465 (I707445,I707406,I707315);
nand I_41466 (I707023,I707298,I707445);
not I_41467 (I707476,I707406);
nor I_41468 (I707493,I707476,I707216);
DFFARX1 I_41469 (I707493,I2507,I707046,I707035,);
nor I_41470 (I707524,I1188441,I1188423);
or I_41471 (I707026,I707273,I707524);
nor I_41472 (I707017,I707406,I707524);
or I_41473 (I707020,I707140,I707524);
DFFARX1 I_41474 (I707524,I2507,I707046,I707038,);
not I_41475 (I707624,I2514);
DFFARX1 I_41476 (I228770,I2507,I707624,I707650,);
not I_41477 (I707658,I707650);
nand I_41478 (I707675,I228773,I228794);
and I_41479 (I707692,I707675,I228782);
DFFARX1 I_41480 (I707692,I2507,I707624,I707718,);
not I_41481 (I707726,I228779);
DFFARX1 I_41482 (I228770,I2507,I707624,I707752,);
not I_41483 (I707760,I707752);
nor I_41484 (I707777,I707760,I707658);
and I_41485 (I707794,I707777,I228779);
nor I_41486 (I707811,I707760,I707726);
nor I_41487 (I707607,I707718,I707811);
DFFARX1 I_41488 (I228788,I2507,I707624,I707851,);
nor I_41489 (I707859,I707851,I707718);
not I_41490 (I707876,I707859);
not I_41491 (I707893,I707851);
nor I_41492 (I707910,I707893,I707794);
DFFARX1 I_41493 (I707910,I2507,I707624,I707610,);
nand I_41494 (I707941,I228773,I228776);
and I_41495 (I707958,I707941,I228785);
DFFARX1 I_41496 (I707958,I2507,I707624,I707984,);
nor I_41497 (I707992,I707984,I707851);
DFFARX1 I_41498 (I707992,I2507,I707624,I707592,);
nand I_41499 (I708023,I707984,I707893);
nand I_41500 (I707601,I707876,I708023);
not I_41501 (I708054,I707984);
nor I_41502 (I708071,I708054,I707794);
DFFARX1 I_41503 (I708071,I2507,I707624,I707613,);
nor I_41504 (I708102,I228791,I228776);
or I_41505 (I707604,I707851,I708102);
nor I_41506 (I707595,I707984,I708102);
or I_41507 (I707598,I707718,I708102);
DFFARX1 I_41508 (I708102,I2507,I707624,I707616,);
not I_41509 (I708202,I2514);
DFFARX1 I_41510 (I1056710,I2507,I708202,I708228,);
not I_41511 (I708236,I708228);
nand I_41512 (I708253,I1056707,I1056725);
and I_41513 (I708270,I708253,I1056722);
DFFARX1 I_41514 (I708270,I2507,I708202,I708296,);
not I_41515 (I708304,I1056704);
DFFARX1 I_41516 (I1056707,I2507,I708202,I708330,);
not I_41517 (I708338,I708330);
nor I_41518 (I708355,I708338,I708236);
and I_41519 (I708372,I708355,I1056704);
nor I_41520 (I708389,I708338,I708304);
nor I_41521 (I708185,I708296,I708389);
DFFARX1 I_41522 (I1056716,I2507,I708202,I708429,);
nor I_41523 (I708437,I708429,I708296);
not I_41524 (I708454,I708437);
not I_41525 (I708471,I708429);
nor I_41526 (I708488,I708471,I708372);
DFFARX1 I_41527 (I708488,I2507,I708202,I708188,);
nand I_41528 (I708519,I1056719,I1056704);
and I_41529 (I708536,I708519,I1056710);
DFFARX1 I_41530 (I708536,I2507,I708202,I708562,);
nor I_41531 (I708570,I708562,I708429);
DFFARX1 I_41532 (I708570,I2507,I708202,I708170,);
nand I_41533 (I708601,I708562,I708471);
nand I_41534 (I708179,I708454,I708601);
not I_41535 (I708632,I708562);
nor I_41536 (I708649,I708632,I708372);
DFFARX1 I_41537 (I708649,I2507,I708202,I708191,);
nor I_41538 (I708680,I1056713,I1056704);
or I_41539 (I708182,I708429,I708680);
nor I_41540 (I708173,I708562,I708680);
or I_41541 (I708176,I708296,I708680);
DFFARX1 I_41542 (I708680,I2507,I708202,I708194,);
not I_41543 (I708780,I2514);
DFFARX1 I_41544 (I779602,I2507,I708780,I708806,);
not I_41545 (I708814,I708806);
nand I_41546 (I708831,I779590,I779608);
and I_41547 (I708848,I708831,I779605);
DFFARX1 I_41548 (I708848,I2507,I708780,I708874,);
not I_41549 (I708882,I779596);
DFFARX1 I_41550 (I779593,I2507,I708780,I708908,);
not I_41551 (I708916,I708908);
nor I_41552 (I708933,I708916,I708814);
and I_41553 (I708950,I708933,I779596);
nor I_41554 (I708967,I708916,I708882);
nor I_41555 (I708763,I708874,I708967);
DFFARX1 I_41556 (I779587,I2507,I708780,I709007,);
nor I_41557 (I709015,I709007,I708874);
not I_41558 (I709032,I709015);
not I_41559 (I709049,I709007);
nor I_41560 (I709066,I709049,I708950);
DFFARX1 I_41561 (I709066,I2507,I708780,I708766,);
nand I_41562 (I709097,I779587,I779590);
and I_41563 (I709114,I709097,I779593);
DFFARX1 I_41564 (I709114,I2507,I708780,I709140,);
nor I_41565 (I709148,I709140,I709007);
DFFARX1 I_41566 (I709148,I2507,I708780,I708748,);
nand I_41567 (I709179,I709140,I709049);
nand I_41568 (I708757,I709032,I709179);
not I_41569 (I709210,I709140);
nor I_41570 (I709227,I709210,I708950);
DFFARX1 I_41571 (I709227,I2507,I708780,I708769,);
nor I_41572 (I709258,I779599,I779590);
or I_41573 (I708760,I709007,I709258);
nor I_41574 (I708751,I709140,I709258);
or I_41575 (I708754,I708874,I709258);
DFFARX1 I_41576 (I709258,I2507,I708780,I708772,);
not I_41577 (I709358,I2514);
DFFARX1 I_41578 (I1057832,I2507,I709358,I709384,);
not I_41579 (I709392,I709384);
nand I_41580 (I709409,I1057829,I1057847);
and I_41581 (I709426,I709409,I1057844);
DFFARX1 I_41582 (I709426,I2507,I709358,I709452,);
not I_41583 (I709460,I1057826);
DFFARX1 I_41584 (I1057829,I2507,I709358,I709486,);
not I_41585 (I709494,I709486);
nor I_41586 (I709511,I709494,I709392);
and I_41587 (I709528,I709511,I1057826);
nor I_41588 (I709545,I709494,I709460);
nor I_41589 (I709341,I709452,I709545);
DFFARX1 I_41590 (I1057838,I2507,I709358,I709585,);
nor I_41591 (I709593,I709585,I709452);
not I_41592 (I709610,I709593);
not I_41593 (I709627,I709585);
nor I_41594 (I709644,I709627,I709528);
DFFARX1 I_41595 (I709644,I2507,I709358,I709344,);
nand I_41596 (I709675,I1057841,I1057826);
and I_41597 (I709692,I709675,I1057832);
DFFARX1 I_41598 (I709692,I2507,I709358,I709718,);
nor I_41599 (I709726,I709718,I709585);
DFFARX1 I_41600 (I709726,I2507,I709358,I709326,);
nand I_41601 (I709757,I709718,I709627);
nand I_41602 (I709335,I709610,I709757);
not I_41603 (I709788,I709718);
nor I_41604 (I709805,I709788,I709528);
DFFARX1 I_41605 (I709805,I2507,I709358,I709347,);
nor I_41606 (I709836,I1057835,I1057826);
or I_41607 (I709338,I709585,I709836);
nor I_41608 (I709329,I709718,I709836);
or I_41609 (I709332,I709452,I709836);
DFFARX1 I_41610 (I709836,I2507,I709358,I709350,);
not I_41611 (I709936,I2514);
DFFARX1 I_41612 (I807533,I2507,I709936,I709962,);
not I_41613 (I709970,I709962);
nand I_41614 (I709987,I807521,I807539);
and I_41615 (I710004,I709987,I807536);
DFFARX1 I_41616 (I710004,I2507,I709936,I710030,);
not I_41617 (I710038,I807527);
DFFARX1 I_41618 (I807524,I2507,I709936,I710064,);
not I_41619 (I710072,I710064);
nor I_41620 (I710089,I710072,I709970);
and I_41621 (I710106,I710089,I807527);
nor I_41622 (I710123,I710072,I710038);
nor I_41623 (I709919,I710030,I710123);
DFFARX1 I_41624 (I807518,I2507,I709936,I710163,);
nor I_41625 (I710171,I710163,I710030);
not I_41626 (I710188,I710171);
not I_41627 (I710205,I710163);
nor I_41628 (I710222,I710205,I710106);
DFFARX1 I_41629 (I710222,I2507,I709936,I709922,);
nand I_41630 (I710253,I807518,I807521);
and I_41631 (I710270,I710253,I807524);
DFFARX1 I_41632 (I710270,I2507,I709936,I710296,);
nor I_41633 (I710304,I710296,I710163);
DFFARX1 I_41634 (I710304,I2507,I709936,I709904,);
nand I_41635 (I710335,I710296,I710205);
nand I_41636 (I709913,I710188,I710335);
not I_41637 (I710366,I710296);
nor I_41638 (I710383,I710366,I710106);
DFFARX1 I_41639 (I710383,I2507,I709936,I709925,);
nor I_41640 (I710414,I807530,I807521);
or I_41641 (I709916,I710163,I710414);
nor I_41642 (I709907,I710296,I710414);
or I_41643 (I709910,I710030,I710414);
DFFARX1 I_41644 (I710414,I2507,I709936,I709928,);
not I_41645 (I710514,I2514);
DFFARX1 I_41646 (I964469,I2507,I710514,I710540,);
not I_41647 (I710548,I710540);
nand I_41648 (I710565,I964445,I964460);
and I_41649 (I710582,I710565,I964472);
DFFARX1 I_41650 (I710582,I2507,I710514,I710608,);
not I_41651 (I710616,I964457);
DFFARX1 I_41652 (I964448,I2507,I710514,I710642,);
not I_41653 (I710650,I710642);
nor I_41654 (I710667,I710650,I710548);
and I_41655 (I710684,I710667,I964457);
nor I_41656 (I710701,I710650,I710616);
nor I_41657 (I710497,I710608,I710701);
DFFARX1 I_41658 (I964445,I2507,I710514,I710741,);
nor I_41659 (I710749,I710741,I710608);
not I_41660 (I710766,I710749);
not I_41661 (I710783,I710741);
nor I_41662 (I710800,I710783,I710684);
DFFARX1 I_41663 (I710800,I2507,I710514,I710500,);
nand I_41664 (I710831,I964463,I964454);
and I_41665 (I710848,I710831,I964466);
DFFARX1 I_41666 (I710848,I2507,I710514,I710874,);
nor I_41667 (I710882,I710874,I710741);
DFFARX1 I_41668 (I710882,I2507,I710514,I710482,);
nand I_41669 (I710913,I710874,I710783);
nand I_41670 (I710491,I710766,I710913);
not I_41671 (I710944,I710874);
nor I_41672 (I710961,I710944,I710684);
DFFARX1 I_41673 (I710961,I2507,I710514,I710503,);
nor I_41674 (I710992,I964451,I964454);
or I_41675 (I710494,I710741,I710992);
nor I_41676 (I710485,I710874,I710992);
or I_41677 (I710488,I710608,I710992);
DFFARX1 I_41678 (I710992,I2507,I710514,I710506,);
not I_41679 (I711092,I2514);
DFFARX1 I_41680 (I569450,I2507,I711092,I711118,);
not I_41681 (I711126,I711118);
nand I_41682 (I711143,I569459,I569468);
and I_41683 (I711160,I711143,I569474);
DFFARX1 I_41684 (I711160,I2507,I711092,I711186,);
not I_41685 (I711194,I569471);
DFFARX1 I_41686 (I569456,I2507,I711092,I711220,);
not I_41687 (I711228,I711220);
nor I_41688 (I711245,I711228,I711126);
and I_41689 (I711262,I711245,I569471);
nor I_41690 (I711279,I711228,I711194);
nor I_41691 (I711075,I711186,I711279);
DFFARX1 I_41692 (I569465,I2507,I711092,I711319,);
nor I_41693 (I711327,I711319,I711186);
not I_41694 (I711344,I711327);
not I_41695 (I711361,I711319);
nor I_41696 (I711378,I711361,I711262);
DFFARX1 I_41697 (I711378,I2507,I711092,I711078,);
nand I_41698 (I711409,I569462,I569453);
and I_41699 (I711426,I711409,I569450);
DFFARX1 I_41700 (I711426,I2507,I711092,I711452,);
nor I_41701 (I711460,I711452,I711319);
DFFARX1 I_41702 (I711460,I2507,I711092,I711060,);
nand I_41703 (I711491,I711452,I711361);
nand I_41704 (I711069,I711344,I711491);
not I_41705 (I711522,I711452);
nor I_41706 (I711539,I711522,I711262);
DFFARX1 I_41707 (I711539,I2507,I711092,I711081,);
nor I_41708 (I711570,I569453,I569453);
or I_41709 (I711072,I711319,I711570);
nor I_41710 (I711063,I711452,I711570);
or I_41711 (I711066,I711186,I711570);
DFFARX1 I_41712 (I711570,I2507,I711092,I711084,);
not I_41713 (I711670,I2514);
DFFARX1 I_41714 (I434360,I2507,I711670,I711696,);
not I_41715 (I711704,I711696);
nand I_41716 (I711721,I434351,I434369);
and I_41717 (I711738,I711721,I434372);
DFFARX1 I_41718 (I711738,I2507,I711670,I711764,);
not I_41719 (I711772,I434366);
DFFARX1 I_41720 (I434354,I2507,I711670,I711798,);
not I_41721 (I711806,I711798);
nor I_41722 (I711823,I711806,I711704);
and I_41723 (I711840,I711823,I434366);
nor I_41724 (I711857,I711806,I711772);
nor I_41725 (I711653,I711764,I711857);
DFFARX1 I_41726 (I434363,I2507,I711670,I711897,);
nor I_41727 (I711905,I711897,I711764);
not I_41728 (I711922,I711905);
not I_41729 (I711939,I711897);
nor I_41730 (I711956,I711939,I711840);
DFFARX1 I_41731 (I711956,I2507,I711670,I711656,);
nand I_41732 (I711987,I434378,I434375);
and I_41733 (I712004,I711987,I434357);
DFFARX1 I_41734 (I712004,I2507,I711670,I712030,);
nor I_41735 (I712038,I712030,I711897);
DFFARX1 I_41736 (I712038,I2507,I711670,I711638,);
nand I_41737 (I712069,I712030,I711939);
nand I_41738 (I711647,I711922,I712069);
not I_41739 (I712100,I712030);
nor I_41740 (I712117,I712100,I711840);
DFFARX1 I_41741 (I712117,I2507,I711670,I711659,);
nor I_41742 (I712148,I434351,I434375);
or I_41743 (I711650,I711897,I712148);
nor I_41744 (I711641,I712030,I712148);
or I_41745 (I711644,I711764,I712148);
DFFARX1 I_41746 (I712148,I2507,I711670,I711662,);
not I_41747 (I712248,I2514);
DFFARX1 I_41748 (I1368409,I2507,I712248,I712274,);
not I_41749 (I712282,I712274);
nand I_41750 (I712299,I1368394,I1368382);
and I_41751 (I712316,I712299,I1368397);
DFFARX1 I_41752 (I712316,I2507,I712248,I712342,);
not I_41753 (I712350,I1368382);
DFFARX1 I_41754 (I1368400,I2507,I712248,I712376,);
not I_41755 (I712384,I712376);
nor I_41756 (I712401,I712384,I712282);
and I_41757 (I712418,I712401,I1368382);
nor I_41758 (I712435,I712384,I712350);
nor I_41759 (I712231,I712342,I712435);
DFFARX1 I_41760 (I1368388,I2507,I712248,I712475,);
nor I_41761 (I712483,I712475,I712342);
not I_41762 (I712500,I712483);
not I_41763 (I712517,I712475);
nor I_41764 (I712534,I712517,I712418);
DFFARX1 I_41765 (I712534,I2507,I712248,I712234,);
nand I_41766 (I712565,I1368385,I1368391);
and I_41767 (I712582,I712565,I1368406);
DFFARX1 I_41768 (I712582,I2507,I712248,I712608,);
nor I_41769 (I712616,I712608,I712475);
DFFARX1 I_41770 (I712616,I2507,I712248,I712216,);
nand I_41771 (I712647,I712608,I712517);
nand I_41772 (I712225,I712500,I712647);
not I_41773 (I712678,I712608);
nor I_41774 (I712695,I712678,I712418);
DFFARX1 I_41775 (I712695,I2507,I712248,I712237,);
nor I_41776 (I712726,I1368403,I1368391);
or I_41777 (I712228,I712475,I712726);
nor I_41778 (I712219,I712608,I712726);
or I_41779 (I712222,I712342,I712726);
DFFARX1 I_41780 (I712726,I2507,I712248,I712240,);
not I_41781 (I712826,I2514);
DFFARX1 I_41782 (I35373,I2507,I712826,I712852,);
not I_41783 (I712860,I712852);
nand I_41784 (I712877,I35370,I35361);
and I_41785 (I712894,I712877,I35361);
DFFARX1 I_41786 (I712894,I2507,I712826,I712920,);
not I_41787 (I712928,I35364);
DFFARX1 I_41788 (I35379,I2507,I712826,I712954,);
not I_41789 (I712962,I712954);
nor I_41790 (I712979,I712962,I712860);
and I_41791 (I712996,I712979,I35364);
nor I_41792 (I713013,I712962,I712928);
nor I_41793 (I712809,I712920,I713013);
DFFARX1 I_41794 (I35364,I2507,I712826,I713053,);
nor I_41795 (I713061,I713053,I712920);
not I_41796 (I713078,I713061);
not I_41797 (I713095,I713053);
nor I_41798 (I713112,I713095,I712996);
DFFARX1 I_41799 (I713112,I2507,I712826,I712812,);
nand I_41800 (I713143,I35382,I35367);
and I_41801 (I713160,I713143,I35385);
DFFARX1 I_41802 (I713160,I2507,I712826,I713186,);
nor I_41803 (I713194,I713186,I713053);
DFFARX1 I_41804 (I713194,I2507,I712826,I712794,);
nand I_41805 (I713225,I713186,I713095);
nand I_41806 (I712803,I713078,I713225);
not I_41807 (I713256,I713186);
nor I_41808 (I713273,I713256,I712996);
DFFARX1 I_41809 (I713273,I2507,I712826,I712815,);
nor I_41810 (I713304,I35376,I35367);
or I_41811 (I712806,I713053,I713304);
nor I_41812 (I712797,I713186,I713304);
or I_41813 (I712800,I712920,I713304);
DFFARX1 I_41814 (I713304,I2507,I712826,I712818,);
not I_41815 (I713404,I2514);
DFFARX1 I_41816 (I1304239,I2507,I713404,I713430,);
not I_41817 (I713438,I713430);
nand I_41818 (I713455,I1304227,I1304245);
and I_41819 (I713472,I713455,I1304236);
DFFARX1 I_41820 (I713472,I2507,I713404,I713498,);
not I_41821 (I713506,I1304251);
DFFARX1 I_41822 (I1304248,I2507,I713404,I713532,);
not I_41823 (I713540,I713532);
nor I_41824 (I713557,I713540,I713438);
and I_41825 (I713574,I713557,I1304251);
nor I_41826 (I713591,I713540,I713506);
nor I_41827 (I713387,I713498,I713591);
DFFARX1 I_41828 (I1304230,I2507,I713404,I713631,);
nor I_41829 (I713639,I713631,I713498);
not I_41830 (I713656,I713639);
not I_41831 (I713673,I713631);
nor I_41832 (I713690,I713673,I713574);
DFFARX1 I_41833 (I713690,I2507,I713404,I713390,);
nand I_41834 (I713721,I1304224,I1304224);
and I_41835 (I713738,I713721,I1304233);
DFFARX1 I_41836 (I713738,I2507,I713404,I713764,);
nor I_41837 (I713772,I713764,I713631);
DFFARX1 I_41838 (I713772,I2507,I713404,I713372,);
nand I_41839 (I713803,I713764,I713673);
nand I_41840 (I713381,I713656,I713803);
not I_41841 (I713834,I713764);
nor I_41842 (I713851,I713834,I713574);
DFFARX1 I_41843 (I713851,I2507,I713404,I713393,);
nor I_41844 (I713882,I1304242,I1304224);
or I_41845 (I713384,I713631,I713882);
nor I_41846 (I713375,I713764,I713882);
or I_41847 (I713378,I713498,I713882);
DFFARX1 I_41848 (I713882,I2507,I713404,I713396,);
not I_41849 (I713982,I2514);
DFFARX1 I_41850 (I831248,I2507,I713982,I714008,);
not I_41851 (I714016,I714008);
nand I_41852 (I714033,I831236,I831254);
and I_41853 (I714050,I714033,I831251);
DFFARX1 I_41854 (I714050,I2507,I713982,I714076,);
not I_41855 (I714084,I831242);
DFFARX1 I_41856 (I831239,I2507,I713982,I714110,);
not I_41857 (I714118,I714110);
nor I_41858 (I714135,I714118,I714016);
and I_41859 (I714152,I714135,I831242);
nor I_41860 (I714169,I714118,I714084);
nor I_41861 (I713965,I714076,I714169);
DFFARX1 I_41862 (I831233,I2507,I713982,I714209,);
nor I_41863 (I714217,I714209,I714076);
not I_41864 (I714234,I714217);
not I_41865 (I714251,I714209);
nor I_41866 (I714268,I714251,I714152);
DFFARX1 I_41867 (I714268,I2507,I713982,I713968,);
nand I_41868 (I714299,I831233,I831236);
and I_41869 (I714316,I714299,I831239);
DFFARX1 I_41870 (I714316,I2507,I713982,I714342,);
nor I_41871 (I714350,I714342,I714209);
DFFARX1 I_41872 (I714350,I2507,I713982,I713950,);
nand I_41873 (I714381,I714342,I714251);
nand I_41874 (I713959,I714234,I714381);
not I_41875 (I714412,I714342);
nor I_41876 (I714429,I714412,I714152);
DFFARX1 I_41877 (I714429,I2507,I713982,I713971,);
nor I_41878 (I714460,I831245,I831236);
or I_41879 (I713962,I714209,I714460);
nor I_41880 (I713953,I714342,I714460);
or I_41881 (I713956,I714076,I714460);
DFFARX1 I_41882 (I714460,I2507,I713982,I713974,);
not I_41883 (I714560,I2514);
DFFARX1 I_41884 (I1010147,I2507,I714560,I714586,);
not I_41885 (I714594,I714586);
nand I_41886 (I714611,I1010144,I1010162);
and I_41887 (I714628,I714611,I1010159);
DFFARX1 I_41888 (I714628,I2507,I714560,I714654,);
not I_41889 (I714662,I1010141);
DFFARX1 I_41890 (I1010144,I2507,I714560,I714688,);
not I_41891 (I714696,I714688);
nor I_41892 (I714713,I714696,I714594);
and I_41893 (I714730,I714713,I1010141);
nor I_41894 (I714747,I714696,I714662);
nor I_41895 (I714543,I714654,I714747);
DFFARX1 I_41896 (I1010153,I2507,I714560,I714787,);
nor I_41897 (I714795,I714787,I714654);
not I_41898 (I714812,I714795);
not I_41899 (I714829,I714787);
nor I_41900 (I714846,I714829,I714730);
DFFARX1 I_41901 (I714846,I2507,I714560,I714546,);
nand I_41902 (I714877,I1010156,I1010141);
and I_41903 (I714894,I714877,I1010147);
DFFARX1 I_41904 (I714894,I2507,I714560,I714920,);
nor I_41905 (I714928,I714920,I714787);
DFFARX1 I_41906 (I714928,I2507,I714560,I714528,);
nand I_41907 (I714959,I714920,I714829);
nand I_41908 (I714537,I714812,I714959);
not I_41909 (I714990,I714920);
nor I_41910 (I715007,I714990,I714730);
DFFARX1 I_41911 (I715007,I2507,I714560,I714549,);
nor I_41912 (I715038,I1010150,I1010141);
or I_41913 (I714540,I714787,I715038);
nor I_41914 (I714531,I714920,I715038);
or I_41915 (I714534,I714654,I715038);
DFFARX1 I_41916 (I715038,I2507,I714560,I714552,);
not I_41917 (I715138,I2514);
DFFARX1 I_41918 (I1245506,I2507,I715138,I715164,);
not I_41919 (I715172,I715164);
nand I_41920 (I715189,I1245509,I1245518);
and I_41921 (I715206,I715189,I1245521);
DFFARX1 I_41922 (I715206,I2507,I715138,I715232,);
not I_41923 (I715240,I1245530);
DFFARX1 I_41924 (I1245512,I2507,I715138,I715266,);
not I_41925 (I715274,I715266);
nor I_41926 (I715291,I715274,I715172);
and I_41927 (I715308,I715291,I1245530);
nor I_41928 (I715325,I715274,I715240);
nor I_41929 (I715121,I715232,I715325);
DFFARX1 I_41930 (I1245509,I2507,I715138,I715365,);
nor I_41931 (I715373,I715365,I715232);
not I_41932 (I715390,I715373);
not I_41933 (I715407,I715365);
nor I_41934 (I715424,I715407,I715308);
DFFARX1 I_41935 (I715424,I2507,I715138,I715124,);
nand I_41936 (I715455,I1245527,I1245506);
and I_41937 (I715472,I715455,I1245524);
DFFARX1 I_41938 (I715472,I2507,I715138,I715498,);
nor I_41939 (I715506,I715498,I715365);
DFFARX1 I_41940 (I715506,I2507,I715138,I715106,);
nand I_41941 (I715537,I715498,I715407);
nand I_41942 (I715115,I715390,I715537);
not I_41943 (I715568,I715498);
nor I_41944 (I715585,I715568,I715308);
DFFARX1 I_41945 (I715585,I2507,I715138,I715127,);
nor I_41946 (I715616,I1245515,I1245506);
or I_41947 (I715118,I715365,I715616);
nor I_41948 (I715109,I715498,I715616);
or I_41949 (I715112,I715232,I715616);
DFFARX1 I_41950 (I715616,I2507,I715138,I715130,);
not I_41951 (I715716,I2514);
DFFARX1 I_41952 (I1029782,I2507,I715716,I715742,);
not I_41953 (I715750,I715742);
nand I_41954 (I715767,I1029779,I1029797);
and I_41955 (I715784,I715767,I1029794);
DFFARX1 I_41956 (I715784,I2507,I715716,I715810,);
not I_41957 (I715818,I1029776);
DFFARX1 I_41958 (I1029779,I2507,I715716,I715844,);
not I_41959 (I715852,I715844);
nor I_41960 (I715869,I715852,I715750);
and I_41961 (I715886,I715869,I1029776);
nor I_41962 (I715903,I715852,I715818);
nor I_41963 (I715699,I715810,I715903);
DFFARX1 I_41964 (I1029788,I2507,I715716,I715943,);
nor I_41965 (I715951,I715943,I715810);
not I_41966 (I715968,I715951);
not I_41967 (I715985,I715943);
nor I_41968 (I716002,I715985,I715886);
DFFARX1 I_41969 (I716002,I2507,I715716,I715702,);
nand I_41970 (I716033,I1029791,I1029776);
and I_41971 (I716050,I716033,I1029782);
DFFARX1 I_41972 (I716050,I2507,I715716,I716076,);
nor I_41973 (I716084,I716076,I715943);
DFFARX1 I_41974 (I716084,I2507,I715716,I715684,);
nand I_41975 (I716115,I716076,I715985);
nand I_41976 (I715693,I715968,I716115);
not I_41977 (I716146,I716076);
nor I_41978 (I716163,I716146,I715886);
DFFARX1 I_41979 (I716163,I2507,I715716,I715705,);
nor I_41980 (I716194,I1029785,I1029776);
or I_41981 (I715696,I715943,I716194);
nor I_41982 (I715687,I716076,I716194);
or I_41983 (I715690,I715810,I716194);
DFFARX1 I_41984 (I716194,I2507,I715716,I715708,);
not I_41985 (I716294,I2514);
DFFARX1 I_41986 (I1071682,I2507,I716294,I716320,);
not I_41987 (I716328,I716320);
nand I_41988 (I716345,I1071664,I1071676);
and I_41989 (I716362,I716345,I1071679);
DFFARX1 I_41990 (I716362,I2507,I716294,I716388,);
not I_41991 (I716396,I1071673);
DFFARX1 I_41992 (I1071670,I2507,I716294,I716422,);
not I_41993 (I716430,I716422);
nor I_41994 (I716447,I716430,I716328);
and I_41995 (I716464,I716447,I1071673);
nor I_41996 (I716481,I716430,I716396);
nor I_41997 (I716277,I716388,I716481);
DFFARX1 I_41998 (I1071688,I2507,I716294,I716521,);
nor I_41999 (I716529,I716521,I716388);
not I_42000 (I716546,I716529);
not I_42001 (I716563,I716521);
nor I_42002 (I716580,I716563,I716464);
DFFARX1 I_42003 (I716580,I2507,I716294,I716280,);
nand I_42004 (I716611,I1071667,I1071667);
and I_42005 (I716628,I716611,I1071664);
DFFARX1 I_42006 (I716628,I2507,I716294,I716654,);
nor I_42007 (I716662,I716654,I716521);
DFFARX1 I_42008 (I716662,I2507,I716294,I716262,);
nand I_42009 (I716693,I716654,I716563);
nand I_42010 (I716271,I716546,I716693);
not I_42011 (I716724,I716654);
nor I_42012 (I716741,I716724,I716464);
DFFARX1 I_42013 (I716741,I2507,I716294,I716283,);
nor I_42014 (I716772,I1071685,I1071667);
or I_42015 (I716274,I716521,I716772);
nor I_42016 (I716265,I716654,I716772);
or I_42017 (I716268,I716388,I716772);
DFFARX1 I_42018 (I716772,I2507,I716294,I716286,);
not I_42019 (I716872,I2514);
DFFARX1 I_42020 (I1372574,I2507,I716872,I716898,);
not I_42021 (I716906,I716898);
nand I_42022 (I716923,I1372559,I1372547);
and I_42023 (I716940,I716923,I1372562);
DFFARX1 I_42024 (I716940,I2507,I716872,I716966,);
not I_42025 (I716974,I1372547);
DFFARX1 I_42026 (I1372565,I2507,I716872,I717000,);
not I_42027 (I717008,I717000);
nor I_42028 (I717025,I717008,I716906);
and I_42029 (I717042,I717025,I1372547);
nor I_42030 (I717059,I717008,I716974);
nor I_42031 (I716855,I716966,I717059);
DFFARX1 I_42032 (I1372553,I2507,I716872,I717099,);
nor I_42033 (I717107,I717099,I716966);
not I_42034 (I717124,I717107);
not I_42035 (I717141,I717099);
nor I_42036 (I717158,I717141,I717042);
DFFARX1 I_42037 (I717158,I2507,I716872,I716858,);
nand I_42038 (I717189,I1372550,I1372556);
and I_42039 (I717206,I717189,I1372571);
DFFARX1 I_42040 (I717206,I2507,I716872,I717232,);
nor I_42041 (I717240,I717232,I717099);
DFFARX1 I_42042 (I717240,I2507,I716872,I716840,);
nand I_42043 (I717271,I717232,I717141);
nand I_42044 (I716849,I717124,I717271);
not I_42045 (I717302,I717232);
nor I_42046 (I717319,I717302,I717042);
DFFARX1 I_42047 (I717319,I2507,I716872,I716861,);
nor I_42048 (I717350,I1372568,I1372556);
or I_42049 (I716852,I717099,I717350);
nor I_42050 (I716843,I717232,I717350);
or I_42051 (I716846,I716966,I717350);
DFFARX1 I_42052 (I717350,I2507,I716872,I716864,);
not I_42053 (I717450,I2514);
DFFARX1 I_42054 (I249595,I2507,I717450,I717476,);
not I_42055 (I717484,I717476);
nand I_42056 (I717501,I249598,I249619);
and I_42057 (I717518,I717501,I249607);
DFFARX1 I_42058 (I717518,I2507,I717450,I717544,);
not I_42059 (I717552,I249604);
DFFARX1 I_42060 (I249595,I2507,I717450,I717578,);
not I_42061 (I717586,I717578);
nor I_42062 (I717603,I717586,I717484);
and I_42063 (I717620,I717603,I249604);
nor I_42064 (I717637,I717586,I717552);
nor I_42065 (I717433,I717544,I717637);
DFFARX1 I_42066 (I249613,I2507,I717450,I717677,);
nor I_42067 (I717685,I717677,I717544);
not I_42068 (I717702,I717685);
not I_42069 (I717719,I717677);
nor I_42070 (I717736,I717719,I717620);
DFFARX1 I_42071 (I717736,I2507,I717450,I717436,);
nand I_42072 (I717767,I249598,I249601);
and I_42073 (I717784,I717767,I249610);
DFFARX1 I_42074 (I717784,I2507,I717450,I717810,);
nor I_42075 (I717818,I717810,I717677);
DFFARX1 I_42076 (I717818,I2507,I717450,I717418,);
nand I_42077 (I717849,I717810,I717719);
nand I_42078 (I717427,I717702,I717849);
not I_42079 (I717880,I717810);
nor I_42080 (I717897,I717880,I717620);
DFFARX1 I_42081 (I717897,I2507,I717450,I717439,);
nor I_42082 (I717928,I249616,I249601);
or I_42083 (I717430,I717677,I717928);
nor I_42084 (I717421,I717810,I717928);
or I_42085 (I717424,I717544,I717928);
DFFARX1 I_42086 (I717928,I2507,I717450,I717442,);
not I_42087 (I718028,I2514);
DFFARX1 I_42088 (I985787,I2507,I718028,I718054,);
not I_42089 (I718062,I718054);
nand I_42090 (I718079,I985763,I985778);
and I_42091 (I718096,I718079,I985790);
DFFARX1 I_42092 (I718096,I2507,I718028,I718122,);
not I_42093 (I718130,I985775);
DFFARX1 I_42094 (I985766,I2507,I718028,I718156,);
not I_42095 (I718164,I718156);
nor I_42096 (I718181,I718164,I718062);
and I_42097 (I718198,I718181,I985775);
nor I_42098 (I718215,I718164,I718130);
nor I_42099 (I718011,I718122,I718215);
DFFARX1 I_42100 (I985763,I2507,I718028,I718255,);
nor I_42101 (I718263,I718255,I718122);
not I_42102 (I718280,I718263);
not I_42103 (I718297,I718255);
nor I_42104 (I718314,I718297,I718198);
DFFARX1 I_42105 (I718314,I2507,I718028,I718014,);
nand I_42106 (I718345,I985781,I985772);
and I_42107 (I718362,I718345,I985784);
DFFARX1 I_42108 (I718362,I2507,I718028,I718388,);
nor I_42109 (I718396,I718388,I718255);
DFFARX1 I_42110 (I718396,I2507,I718028,I717996,);
nand I_42111 (I718427,I718388,I718297);
nand I_42112 (I718005,I718280,I718427);
not I_42113 (I718458,I718388);
nor I_42114 (I718475,I718458,I718198);
DFFARX1 I_42115 (I718475,I2507,I718028,I718017,);
nor I_42116 (I718506,I985769,I985772);
or I_42117 (I718008,I718255,I718506);
nor I_42118 (I717999,I718388,I718506);
or I_42119 (I718002,I718122,I718506);
DFFARX1 I_42120 (I718506,I2507,I718028,I718020,);
not I_42121 (I718606,I2514);
DFFARX1 I_42122 (I369843,I2507,I718606,I718632,);
not I_42123 (I718640,I718632);
nand I_42124 (I718657,I369846,I369822);
and I_42125 (I718674,I718657,I369819);
DFFARX1 I_42126 (I718674,I2507,I718606,I718700,);
not I_42127 (I718708,I369825);
DFFARX1 I_42128 (I369819,I2507,I718606,I718734,);
not I_42129 (I718742,I718734);
nor I_42130 (I718759,I718742,I718640);
and I_42131 (I718776,I718759,I369825);
nor I_42132 (I718793,I718742,I718708);
nor I_42133 (I718589,I718700,I718793);
DFFARX1 I_42134 (I369828,I2507,I718606,I718833,);
nor I_42135 (I718841,I718833,I718700);
not I_42136 (I718858,I718841);
not I_42137 (I718875,I718833);
nor I_42138 (I718892,I718875,I718776);
DFFARX1 I_42139 (I718892,I2507,I718606,I718592,);
nand I_42140 (I718923,I369831,I369840);
and I_42141 (I718940,I718923,I369837);
DFFARX1 I_42142 (I718940,I2507,I718606,I718966,);
nor I_42143 (I718974,I718966,I718833);
DFFARX1 I_42144 (I718974,I2507,I718606,I718574,);
nand I_42145 (I719005,I718966,I718875);
nand I_42146 (I718583,I718858,I719005);
not I_42147 (I719036,I718966);
nor I_42148 (I719053,I719036,I718776);
DFFARX1 I_42149 (I719053,I2507,I718606,I718595,);
nor I_42150 (I719084,I369834,I369840);
or I_42151 (I718586,I718833,I719084);
nor I_42152 (I718577,I718966,I719084);
or I_42153 (I718580,I718700,I719084);
DFFARX1 I_42154 (I719084,I2507,I718606,I718598,);
not I_42155 (I719184,I2514);
DFFARX1 I_42156 (I1764,I2507,I719184,I719210,);
not I_42157 (I719218,I719210);
nand I_42158 (I719235,I1372,I1868);
and I_42159 (I719252,I719235,I1748);
DFFARX1 I_42160 (I719252,I2507,I719184,I719278,);
not I_42161 (I719286,I1564);
DFFARX1 I_42162 (I2044,I2507,I719184,I719312,);
not I_42163 (I719320,I719312);
nor I_42164 (I719337,I719320,I719218);
and I_42165 (I719354,I719337,I1564);
nor I_42166 (I719371,I719320,I719286);
nor I_42167 (I719167,I719278,I719371);
DFFARX1 I_42168 (I2244,I2507,I719184,I719411,);
nor I_42169 (I719419,I719411,I719278);
not I_42170 (I719436,I719419);
not I_42171 (I719453,I719411);
nor I_42172 (I719470,I719453,I719354);
DFFARX1 I_42173 (I719470,I2507,I719184,I719170,);
nand I_42174 (I719501,I2156,I1724);
and I_42175 (I719518,I719501,I2340);
DFFARX1 I_42176 (I719518,I2507,I719184,I719544,);
nor I_42177 (I719552,I719544,I719411);
DFFARX1 I_42178 (I719552,I2507,I719184,I719152,);
nand I_42179 (I719583,I719544,I719453);
nand I_42180 (I719161,I719436,I719583);
not I_42181 (I719614,I719544);
nor I_42182 (I719631,I719614,I719354);
DFFARX1 I_42183 (I719631,I2507,I719184,I719173,);
nor I_42184 (I719662,I2324,I1724);
or I_42185 (I719164,I719411,I719662);
nor I_42186 (I719155,I719544,I719662);
or I_42187 (I719158,I719278,I719662);
DFFARX1 I_42188 (I719662,I2507,I719184,I719176,);
not I_42189 (I719762,I2514);
DFFARX1 I_42190 (I450680,I2507,I719762,I719788,);
not I_42191 (I719796,I719788);
nand I_42192 (I719813,I450671,I450689);
and I_42193 (I719830,I719813,I450692);
DFFARX1 I_42194 (I719830,I2507,I719762,I719856,);
not I_42195 (I719864,I450686);
DFFARX1 I_42196 (I450674,I2507,I719762,I719890,);
not I_42197 (I719898,I719890);
nor I_42198 (I719915,I719898,I719796);
and I_42199 (I719932,I719915,I450686);
nor I_42200 (I719949,I719898,I719864);
nor I_42201 (I719745,I719856,I719949);
DFFARX1 I_42202 (I450683,I2507,I719762,I719989,);
nor I_42203 (I719997,I719989,I719856);
not I_42204 (I720014,I719997);
not I_42205 (I720031,I719989);
nor I_42206 (I720048,I720031,I719932);
DFFARX1 I_42207 (I720048,I2507,I719762,I719748,);
nand I_42208 (I720079,I450698,I450695);
and I_42209 (I720096,I720079,I450677);
DFFARX1 I_42210 (I720096,I2507,I719762,I720122,);
nor I_42211 (I720130,I720122,I719989);
DFFARX1 I_42212 (I720130,I2507,I719762,I719730,);
nand I_42213 (I720161,I720122,I720031);
nand I_42214 (I719739,I720014,I720161);
not I_42215 (I720192,I720122);
nor I_42216 (I720209,I720192,I719932);
DFFARX1 I_42217 (I720209,I2507,I719762,I719751,);
nor I_42218 (I720240,I450671,I450695);
or I_42219 (I719742,I719989,I720240);
nor I_42220 (I719733,I720122,I720240);
or I_42221 (I719736,I719856,I720240);
DFFARX1 I_42222 (I720240,I2507,I719762,I719754,);
not I_42223 (I720340,I2514);
DFFARX1 I_42224 (I159750,I2507,I720340,I720366,);
not I_42225 (I720374,I720366);
nand I_42226 (I720391,I159753,I159774);
and I_42227 (I720408,I720391,I159762);
DFFARX1 I_42228 (I720408,I2507,I720340,I720434,);
not I_42229 (I720442,I159759);
DFFARX1 I_42230 (I159750,I2507,I720340,I720468,);
not I_42231 (I720476,I720468);
nor I_42232 (I720493,I720476,I720374);
and I_42233 (I720510,I720493,I159759);
nor I_42234 (I720527,I720476,I720442);
nor I_42235 (I720323,I720434,I720527);
DFFARX1 I_42236 (I159768,I2507,I720340,I720567,);
nor I_42237 (I720575,I720567,I720434);
not I_42238 (I720592,I720575);
not I_42239 (I720609,I720567);
nor I_42240 (I720626,I720609,I720510);
DFFARX1 I_42241 (I720626,I2507,I720340,I720326,);
nand I_42242 (I720657,I159753,I159756);
and I_42243 (I720674,I720657,I159765);
DFFARX1 I_42244 (I720674,I2507,I720340,I720700,);
nor I_42245 (I720708,I720700,I720567);
DFFARX1 I_42246 (I720708,I2507,I720340,I720308,);
nand I_42247 (I720739,I720700,I720609);
nand I_42248 (I720317,I720592,I720739);
not I_42249 (I720770,I720700);
nor I_42250 (I720787,I720770,I720510);
DFFARX1 I_42251 (I720787,I2507,I720340,I720329,);
nor I_42252 (I720818,I159771,I159756);
or I_42253 (I720320,I720567,I720818);
nor I_42254 (I720311,I720700,I720818);
or I_42255 (I720314,I720434,I720818);
DFFARX1 I_42256 (I720818,I2507,I720340,I720332,);
not I_42257 (I720918,I2514);
DFFARX1 I_42258 (I98604,I2507,I720918,I720944,);
not I_42259 (I720952,I720944);
nand I_42260 (I720969,I98613,I98622);
and I_42261 (I720986,I720969,I98601);
DFFARX1 I_42262 (I720986,I2507,I720918,I721012,);
not I_42263 (I721020,I98604);
DFFARX1 I_42264 (I98619,I2507,I720918,I721046,);
not I_42265 (I721054,I721046);
nor I_42266 (I721071,I721054,I720952);
and I_42267 (I721088,I721071,I98604);
nor I_42268 (I721105,I721054,I721020);
nor I_42269 (I720901,I721012,I721105);
DFFARX1 I_42270 (I98610,I2507,I720918,I721145,);
nor I_42271 (I721153,I721145,I721012);
not I_42272 (I721170,I721153);
not I_42273 (I721187,I721145);
nor I_42274 (I721204,I721187,I721088);
DFFARX1 I_42275 (I721204,I2507,I720918,I720904,);
nand I_42276 (I721235,I98625,I98601);
and I_42277 (I721252,I721235,I98607);
DFFARX1 I_42278 (I721252,I2507,I720918,I721278,);
nor I_42279 (I721286,I721278,I721145);
DFFARX1 I_42280 (I721286,I2507,I720918,I720886,);
nand I_42281 (I721317,I721278,I721187);
nand I_42282 (I720895,I721170,I721317);
not I_42283 (I721348,I721278);
nor I_42284 (I721365,I721348,I721088);
DFFARX1 I_42285 (I721365,I2507,I720918,I720907,);
nor I_42286 (I721396,I98616,I98601);
or I_42287 (I720898,I721145,I721396);
nor I_42288 (I720889,I721278,I721396);
or I_42289 (I720892,I721012,I721396);
DFFARX1 I_42290 (I721396,I2507,I720918,I720910,);
not I_42291 (I721496,I2514);
DFFARX1 I_42292 (I1265736,I2507,I721496,I721522,);
not I_42293 (I721530,I721522);
nand I_42294 (I721547,I1265760,I1265742);
and I_42295 (I721564,I721547,I1265748);
DFFARX1 I_42296 (I721564,I2507,I721496,I721590,);
not I_42297 (I721598,I1265754);
DFFARX1 I_42298 (I1265739,I2507,I721496,I721624,);
not I_42299 (I721632,I721624);
nor I_42300 (I721649,I721632,I721530);
and I_42301 (I721666,I721649,I1265754);
nor I_42302 (I721683,I721632,I721598);
nor I_42303 (I721479,I721590,I721683);
DFFARX1 I_42304 (I1265751,I2507,I721496,I721723,);
nor I_42305 (I721731,I721723,I721590);
not I_42306 (I721748,I721731);
not I_42307 (I721765,I721723);
nor I_42308 (I721782,I721765,I721666);
DFFARX1 I_42309 (I721782,I2507,I721496,I721482,);
nand I_42310 (I721813,I1265757,I1265745);
and I_42311 (I721830,I721813,I1265739);
DFFARX1 I_42312 (I721830,I2507,I721496,I721856,);
nor I_42313 (I721864,I721856,I721723);
DFFARX1 I_42314 (I721864,I2507,I721496,I721464,);
nand I_42315 (I721895,I721856,I721765);
nand I_42316 (I721473,I721748,I721895);
not I_42317 (I721926,I721856);
nor I_42318 (I721943,I721926,I721666);
DFFARX1 I_42319 (I721943,I2507,I721496,I721485,);
nor I_42320 (I721974,I1265736,I1265745);
or I_42321 (I721476,I721723,I721974);
nor I_42322 (I721467,I721856,I721974);
or I_42323 (I721470,I721590,I721974);
DFFARX1 I_42324 (I721974,I2507,I721496,I721488,);
not I_42325 (I722074,I2514);
DFFARX1 I_42326 (I310819,I2507,I722074,I722100,);
not I_42327 (I722108,I722100);
nand I_42328 (I722125,I310822,I310798);
and I_42329 (I722142,I722125,I310795);
DFFARX1 I_42330 (I722142,I2507,I722074,I722168,);
not I_42331 (I722176,I310801);
DFFARX1 I_42332 (I310795,I2507,I722074,I722202,);
not I_42333 (I722210,I722202);
nor I_42334 (I722227,I722210,I722108);
and I_42335 (I722244,I722227,I310801);
nor I_42336 (I722261,I722210,I722176);
nor I_42337 (I722057,I722168,I722261);
DFFARX1 I_42338 (I310804,I2507,I722074,I722301,);
nor I_42339 (I722309,I722301,I722168);
not I_42340 (I722326,I722309);
not I_42341 (I722343,I722301);
nor I_42342 (I722360,I722343,I722244);
DFFARX1 I_42343 (I722360,I2507,I722074,I722060,);
nand I_42344 (I722391,I310807,I310816);
and I_42345 (I722408,I722391,I310813);
DFFARX1 I_42346 (I722408,I2507,I722074,I722434,);
nor I_42347 (I722442,I722434,I722301);
DFFARX1 I_42348 (I722442,I2507,I722074,I722042,);
nand I_42349 (I722473,I722434,I722343);
nand I_42350 (I722051,I722326,I722473);
not I_42351 (I722504,I722434);
nor I_42352 (I722521,I722504,I722244);
DFFARX1 I_42353 (I722521,I2507,I722074,I722063,);
nor I_42354 (I722552,I310810,I310816);
or I_42355 (I722054,I722301,I722552);
nor I_42356 (I722045,I722434,I722552);
or I_42357 (I722048,I722168,I722552);
DFFARX1 I_42358 (I722552,I2507,I722074,I722066,);
not I_42359 (I722652,I2514);
DFFARX1 I_42360 (I396280,I2507,I722652,I722678,);
not I_42361 (I722686,I722678);
nand I_42362 (I722703,I396271,I396289);
and I_42363 (I722720,I722703,I396292);
DFFARX1 I_42364 (I722720,I2507,I722652,I722746,);
not I_42365 (I722754,I396286);
DFFARX1 I_42366 (I396274,I2507,I722652,I722780,);
not I_42367 (I722788,I722780);
nor I_42368 (I722805,I722788,I722686);
and I_42369 (I722822,I722805,I396286);
nor I_42370 (I722839,I722788,I722754);
nor I_42371 (I722635,I722746,I722839);
DFFARX1 I_42372 (I396283,I2507,I722652,I722879,);
nor I_42373 (I722887,I722879,I722746);
not I_42374 (I722904,I722887);
not I_42375 (I722921,I722879);
nor I_42376 (I722938,I722921,I722822);
DFFARX1 I_42377 (I722938,I2507,I722652,I722638,);
nand I_42378 (I722969,I396298,I396295);
and I_42379 (I722986,I722969,I396277);
DFFARX1 I_42380 (I722986,I2507,I722652,I723012,);
nor I_42381 (I723020,I723012,I722879);
DFFARX1 I_42382 (I723020,I2507,I722652,I722620,);
nand I_42383 (I723051,I723012,I722921);
nand I_42384 (I722629,I722904,I723051);
not I_42385 (I723082,I723012);
nor I_42386 (I723099,I723082,I722822);
DFFARX1 I_42387 (I723099,I2507,I722652,I722641,);
nor I_42388 (I723130,I396271,I396295);
or I_42389 (I722632,I722879,I723130);
nor I_42390 (I722623,I723012,I723130);
or I_42391 (I722626,I722746,I723130);
DFFARX1 I_42392 (I723130,I2507,I722652,I722644,);
not I_42393 (I723230,I2514);
DFFARX1 I_42394 (I1092490,I2507,I723230,I723256,);
not I_42395 (I723264,I723256);
nand I_42396 (I723281,I1092472,I1092484);
and I_42397 (I723298,I723281,I1092487);
DFFARX1 I_42398 (I723298,I2507,I723230,I723324,);
not I_42399 (I723332,I1092481);
DFFARX1 I_42400 (I1092478,I2507,I723230,I723358,);
not I_42401 (I723366,I723358);
nor I_42402 (I723383,I723366,I723264);
and I_42403 (I723400,I723383,I1092481);
nor I_42404 (I723417,I723366,I723332);
nor I_42405 (I723213,I723324,I723417);
DFFARX1 I_42406 (I1092496,I2507,I723230,I723457,);
nor I_42407 (I723465,I723457,I723324);
not I_42408 (I723482,I723465);
not I_42409 (I723499,I723457);
nor I_42410 (I723516,I723499,I723400);
DFFARX1 I_42411 (I723516,I2507,I723230,I723216,);
nand I_42412 (I723547,I1092475,I1092475);
and I_42413 (I723564,I723547,I1092472);
DFFARX1 I_42414 (I723564,I2507,I723230,I723590,);
nor I_42415 (I723598,I723590,I723457);
DFFARX1 I_42416 (I723598,I2507,I723230,I723198,);
nand I_42417 (I723629,I723590,I723499);
nand I_42418 (I723207,I723482,I723629);
not I_42419 (I723660,I723590);
nor I_42420 (I723677,I723660,I723400);
DFFARX1 I_42421 (I723677,I2507,I723230,I723219,);
nor I_42422 (I723708,I1092493,I1092475);
or I_42423 (I723210,I723457,I723708);
nor I_42424 (I723201,I723590,I723708);
or I_42425 (I723204,I723324,I723708);
DFFARX1 I_42426 (I723708,I2507,I723230,I723222,);
not I_42427 (I723808,I2514);
DFFARX1 I_42428 (I501229,I2507,I723808,I723834,);
not I_42429 (I723842,I723834);
nand I_42430 (I723859,I501244,I501229);
and I_42431 (I723876,I723859,I501232);
DFFARX1 I_42432 (I723876,I2507,I723808,I723902,);
not I_42433 (I723910,I501232);
DFFARX1 I_42434 (I501241,I2507,I723808,I723936,);
not I_42435 (I723944,I723936);
nor I_42436 (I723961,I723944,I723842);
and I_42437 (I723978,I723961,I501232);
nor I_42438 (I723995,I723944,I723910);
nor I_42439 (I723791,I723902,I723995);
DFFARX1 I_42440 (I501235,I2507,I723808,I724035,);
nor I_42441 (I724043,I724035,I723902);
not I_42442 (I724060,I724043);
not I_42443 (I724077,I724035);
nor I_42444 (I724094,I724077,I723978);
DFFARX1 I_42445 (I724094,I2507,I723808,I723794,);
nand I_42446 (I724125,I501238,I501247);
and I_42447 (I724142,I724125,I501253);
DFFARX1 I_42448 (I724142,I2507,I723808,I724168,);
nor I_42449 (I724176,I724168,I724035);
DFFARX1 I_42450 (I724176,I2507,I723808,I723776,);
nand I_42451 (I724207,I724168,I724077);
nand I_42452 (I723785,I724060,I724207);
not I_42453 (I724238,I724168);
nor I_42454 (I724255,I724238,I723978);
DFFARX1 I_42455 (I724255,I2507,I723808,I723797,);
nor I_42456 (I724286,I501250,I501247);
or I_42457 (I723788,I724035,I724286);
nor I_42458 (I723779,I724168,I724286);
or I_42459 (I723782,I723902,I724286);
DFFARX1 I_42460 (I724286,I2507,I723808,I723800,);
not I_42461 (I724386,I2514);
DFFARX1 I_42462 (I1268626,I2507,I724386,I724412,);
not I_42463 (I724420,I724412);
nand I_42464 (I724437,I1268650,I1268632);
and I_42465 (I724454,I724437,I1268638);
DFFARX1 I_42466 (I724454,I2507,I724386,I724480,);
not I_42467 (I724488,I1268644);
DFFARX1 I_42468 (I1268629,I2507,I724386,I724514,);
not I_42469 (I724522,I724514);
nor I_42470 (I724539,I724522,I724420);
and I_42471 (I724556,I724539,I1268644);
nor I_42472 (I724573,I724522,I724488);
nor I_42473 (I724369,I724480,I724573);
DFFARX1 I_42474 (I1268641,I2507,I724386,I724613,);
nor I_42475 (I724621,I724613,I724480);
not I_42476 (I724638,I724621);
not I_42477 (I724655,I724613);
nor I_42478 (I724672,I724655,I724556);
DFFARX1 I_42479 (I724672,I2507,I724386,I724372,);
nand I_42480 (I724703,I1268647,I1268635);
and I_42481 (I724720,I724703,I1268629);
DFFARX1 I_42482 (I724720,I2507,I724386,I724746,);
nor I_42483 (I724754,I724746,I724613);
DFFARX1 I_42484 (I724754,I2507,I724386,I724354,);
nand I_42485 (I724785,I724746,I724655);
nand I_42486 (I724363,I724638,I724785);
not I_42487 (I724816,I724746);
nor I_42488 (I724833,I724816,I724556);
DFFARX1 I_42489 (I724833,I2507,I724386,I724375,);
nor I_42490 (I724864,I1268626,I1268635);
or I_42491 (I724366,I724613,I724864);
nor I_42492 (I724357,I724746,I724864);
or I_42493 (I724360,I724480,I724864);
DFFARX1 I_42494 (I724864,I2507,I724386,I724378,);
not I_42495 (I724964,I2514);
DFFARX1 I_42496 (I409336,I2507,I724964,I724990,);
not I_42497 (I724998,I724990);
nand I_42498 (I725015,I409327,I409345);
and I_42499 (I725032,I725015,I409348);
DFFARX1 I_42500 (I725032,I2507,I724964,I725058,);
not I_42501 (I725066,I409342);
DFFARX1 I_42502 (I409330,I2507,I724964,I725092,);
not I_42503 (I725100,I725092);
nor I_42504 (I725117,I725100,I724998);
and I_42505 (I725134,I725117,I409342);
nor I_42506 (I725151,I725100,I725066);
nor I_42507 (I724947,I725058,I725151);
DFFARX1 I_42508 (I409339,I2507,I724964,I725191,);
nor I_42509 (I725199,I725191,I725058);
not I_42510 (I725216,I725199);
not I_42511 (I725233,I725191);
nor I_42512 (I725250,I725233,I725134);
DFFARX1 I_42513 (I725250,I2507,I724964,I724950,);
nand I_42514 (I725281,I409354,I409351);
and I_42515 (I725298,I725281,I409333);
DFFARX1 I_42516 (I725298,I2507,I724964,I725324,);
nor I_42517 (I725332,I725324,I725191);
DFFARX1 I_42518 (I725332,I2507,I724964,I724932,);
nand I_42519 (I725363,I725324,I725233);
nand I_42520 (I724941,I725216,I725363);
not I_42521 (I725394,I725324);
nor I_42522 (I725411,I725394,I725134);
DFFARX1 I_42523 (I725411,I2507,I724964,I724953,);
nor I_42524 (I725442,I409327,I409351);
or I_42525 (I724944,I725191,I725442);
nor I_42526 (I724935,I725324,I725442);
or I_42527 (I724938,I725058,I725442);
DFFARX1 I_42528 (I725442,I2507,I724964,I724956,);
not I_42529 (I725542,I2514);
DFFARX1 I_42530 (I546330,I2507,I725542,I725568,);
not I_42531 (I725576,I725568);
nand I_42532 (I725593,I546339,I546348);
and I_42533 (I725610,I725593,I546354);
DFFARX1 I_42534 (I725610,I2507,I725542,I725636,);
not I_42535 (I725644,I546351);
DFFARX1 I_42536 (I546336,I2507,I725542,I725670,);
not I_42537 (I725678,I725670);
nor I_42538 (I725695,I725678,I725576);
and I_42539 (I725712,I725695,I546351);
nor I_42540 (I725729,I725678,I725644);
nor I_42541 (I725525,I725636,I725729);
DFFARX1 I_42542 (I546345,I2507,I725542,I725769,);
nor I_42543 (I725777,I725769,I725636);
not I_42544 (I725794,I725777);
not I_42545 (I725811,I725769);
nor I_42546 (I725828,I725811,I725712);
DFFARX1 I_42547 (I725828,I2507,I725542,I725528,);
nand I_42548 (I725859,I546342,I546333);
and I_42549 (I725876,I725859,I546330);
DFFARX1 I_42550 (I725876,I2507,I725542,I725902,);
nor I_42551 (I725910,I725902,I725769);
DFFARX1 I_42552 (I725910,I2507,I725542,I725510,);
nand I_42553 (I725941,I725902,I725811);
nand I_42554 (I725519,I725794,I725941);
not I_42555 (I725972,I725902);
nor I_42556 (I725989,I725972,I725712);
DFFARX1 I_42557 (I725989,I2507,I725542,I725531,);
nor I_42558 (I726020,I546333,I546333);
or I_42559 (I725522,I725769,I726020);
nor I_42560 (I725513,I725902,I726020);
or I_42561 (I725516,I725636,I726020);
DFFARX1 I_42562 (I726020,I2507,I725542,I725534,);
not I_42563 (I726120,I2514);
DFFARX1 I_42564 (I241265,I2507,I726120,I726146,);
not I_42565 (I726154,I726146);
nand I_42566 (I726171,I241268,I241289);
and I_42567 (I726188,I726171,I241277);
DFFARX1 I_42568 (I726188,I2507,I726120,I726214,);
not I_42569 (I726222,I241274);
DFFARX1 I_42570 (I241265,I2507,I726120,I726248,);
not I_42571 (I726256,I726248);
nor I_42572 (I726273,I726256,I726154);
and I_42573 (I726290,I726273,I241274);
nor I_42574 (I726307,I726256,I726222);
nor I_42575 (I726103,I726214,I726307);
DFFARX1 I_42576 (I241283,I2507,I726120,I726347,);
nor I_42577 (I726355,I726347,I726214);
not I_42578 (I726372,I726355);
not I_42579 (I726389,I726347);
nor I_42580 (I726406,I726389,I726290);
DFFARX1 I_42581 (I726406,I2507,I726120,I726106,);
nand I_42582 (I726437,I241268,I241271);
and I_42583 (I726454,I726437,I241280);
DFFARX1 I_42584 (I726454,I2507,I726120,I726480,);
nor I_42585 (I726488,I726480,I726347);
DFFARX1 I_42586 (I726488,I2507,I726120,I726088,);
nand I_42587 (I726519,I726480,I726389);
nand I_42588 (I726097,I726372,I726519);
not I_42589 (I726550,I726480);
nor I_42590 (I726567,I726550,I726290);
DFFARX1 I_42591 (I726567,I2507,I726120,I726109,);
nor I_42592 (I726598,I241286,I241271);
or I_42593 (I726100,I726347,I726598);
nor I_42594 (I726091,I726480,I726598);
or I_42595 (I726094,I726214,I726598);
DFFARX1 I_42596 (I726598,I2507,I726120,I726112,);
not I_42597 (I726698,I2514);
DFFARX1 I_42598 (I957363,I2507,I726698,I726724,);
not I_42599 (I726732,I726724);
nand I_42600 (I726749,I957339,I957354);
and I_42601 (I726766,I726749,I957366);
DFFARX1 I_42602 (I726766,I2507,I726698,I726792,);
not I_42603 (I726800,I957351);
DFFARX1 I_42604 (I957342,I2507,I726698,I726826,);
not I_42605 (I726834,I726826);
nor I_42606 (I726851,I726834,I726732);
and I_42607 (I726868,I726851,I957351);
nor I_42608 (I726885,I726834,I726800);
nor I_42609 (I726681,I726792,I726885);
DFFARX1 I_42610 (I957339,I2507,I726698,I726925,);
nor I_42611 (I726933,I726925,I726792);
not I_42612 (I726950,I726933);
not I_42613 (I726967,I726925);
nor I_42614 (I726984,I726967,I726868);
DFFARX1 I_42615 (I726984,I2507,I726698,I726684,);
nand I_42616 (I727015,I957357,I957348);
and I_42617 (I727032,I727015,I957360);
DFFARX1 I_42618 (I727032,I2507,I726698,I727058,);
nor I_42619 (I727066,I727058,I726925);
DFFARX1 I_42620 (I727066,I2507,I726698,I726666,);
nand I_42621 (I727097,I727058,I726967);
nand I_42622 (I726675,I726950,I727097);
not I_42623 (I727128,I727058);
nor I_42624 (I727145,I727128,I726868);
DFFARX1 I_42625 (I727145,I2507,I726698,I726687,);
nor I_42626 (I727176,I957345,I957348);
or I_42627 (I726678,I726925,I727176);
nor I_42628 (I726669,I727058,I727176);
or I_42629 (I726672,I726792,I727176);
DFFARX1 I_42630 (I727176,I2507,I726698,I726690,);
not I_42631 (I727276,I2514);
DFFARX1 I_42632 (I249000,I2507,I727276,I727302,);
not I_42633 (I727310,I727302);
nand I_42634 (I727327,I249003,I249024);
and I_42635 (I727344,I727327,I249012);
DFFARX1 I_42636 (I727344,I2507,I727276,I727370,);
not I_42637 (I727378,I249009);
DFFARX1 I_42638 (I249000,I2507,I727276,I727404,);
not I_42639 (I727412,I727404);
nor I_42640 (I727429,I727412,I727310);
and I_42641 (I727446,I727429,I249009);
nor I_42642 (I727463,I727412,I727378);
nor I_42643 (I727259,I727370,I727463);
DFFARX1 I_42644 (I249018,I2507,I727276,I727503,);
nor I_42645 (I727511,I727503,I727370);
not I_42646 (I727528,I727511);
not I_42647 (I727545,I727503);
nor I_42648 (I727562,I727545,I727446);
DFFARX1 I_42649 (I727562,I2507,I727276,I727262,);
nand I_42650 (I727593,I249003,I249006);
and I_42651 (I727610,I727593,I249015);
DFFARX1 I_42652 (I727610,I2507,I727276,I727636,);
nor I_42653 (I727644,I727636,I727503);
DFFARX1 I_42654 (I727644,I2507,I727276,I727244,);
nand I_42655 (I727675,I727636,I727545);
nand I_42656 (I727253,I727528,I727675);
not I_42657 (I727706,I727636);
nor I_42658 (I727723,I727706,I727446);
DFFARX1 I_42659 (I727723,I2507,I727276,I727265,);
nor I_42660 (I727754,I249021,I249006);
or I_42661 (I727256,I727503,I727754);
nor I_42662 (I727247,I727636,I727754);
or I_42663 (I727250,I727370,I727754);
DFFARX1 I_42664 (I727754,I2507,I727276,I727268,);
not I_42665 (I727854,I2514);
DFFARX1 I_42666 (I885657,I2507,I727854,I727880,);
not I_42667 (I727888,I727880);
nand I_42668 (I727905,I885633,I885648);
and I_42669 (I727922,I727905,I885660);
DFFARX1 I_42670 (I727922,I2507,I727854,I727948,);
not I_42671 (I727956,I885645);
DFFARX1 I_42672 (I885636,I2507,I727854,I727982,);
not I_42673 (I727990,I727982);
nor I_42674 (I728007,I727990,I727888);
and I_42675 (I728024,I728007,I885645);
nor I_42676 (I728041,I727990,I727956);
nor I_42677 (I727837,I727948,I728041);
DFFARX1 I_42678 (I885633,I2507,I727854,I728081,);
nor I_42679 (I728089,I728081,I727948);
not I_42680 (I728106,I728089);
not I_42681 (I728123,I728081);
nor I_42682 (I728140,I728123,I728024);
DFFARX1 I_42683 (I728140,I2507,I727854,I727840,);
nand I_42684 (I728171,I885651,I885642);
and I_42685 (I728188,I728171,I885654);
DFFARX1 I_42686 (I728188,I2507,I727854,I728214,);
nor I_42687 (I728222,I728214,I728081);
DFFARX1 I_42688 (I728222,I2507,I727854,I727822,);
nand I_42689 (I728253,I728214,I728123);
nand I_42690 (I727831,I728106,I728253);
not I_42691 (I728284,I728214);
nor I_42692 (I728301,I728284,I728024);
DFFARX1 I_42693 (I728301,I2507,I727854,I727843,);
nor I_42694 (I728332,I885639,I885642);
or I_42695 (I727834,I728081,I728332);
nor I_42696 (I727825,I728214,I728332);
or I_42697 (I727828,I727948,I728332);
DFFARX1 I_42698 (I728332,I2507,I727854,I727846,);
not I_42699 (I728432,I2514);
DFFARX1 I_42700 (I450136,I2507,I728432,I728458,);
not I_42701 (I728466,I728458);
nand I_42702 (I728483,I450127,I450145);
and I_42703 (I728500,I728483,I450148);
DFFARX1 I_42704 (I728500,I2507,I728432,I728526,);
not I_42705 (I728534,I450142);
DFFARX1 I_42706 (I450130,I2507,I728432,I728560,);
not I_42707 (I728568,I728560);
nor I_42708 (I728585,I728568,I728466);
and I_42709 (I728602,I728585,I450142);
nor I_42710 (I728619,I728568,I728534);
nor I_42711 (I728415,I728526,I728619);
DFFARX1 I_42712 (I450139,I2507,I728432,I728659,);
nor I_42713 (I728667,I728659,I728526);
not I_42714 (I728684,I728667);
not I_42715 (I728701,I728659);
nor I_42716 (I728718,I728701,I728602);
DFFARX1 I_42717 (I728718,I2507,I728432,I728418,);
nand I_42718 (I728749,I450154,I450151);
and I_42719 (I728766,I728749,I450133);
DFFARX1 I_42720 (I728766,I2507,I728432,I728792,);
nor I_42721 (I728800,I728792,I728659);
DFFARX1 I_42722 (I728800,I2507,I728432,I728400,);
nand I_42723 (I728831,I728792,I728701);
nand I_42724 (I728409,I728684,I728831);
not I_42725 (I728862,I728792);
nor I_42726 (I728879,I728862,I728602);
DFFARX1 I_42727 (I728879,I2507,I728432,I728421,);
nor I_42728 (I728910,I450127,I450151);
or I_42729 (I728412,I728659,I728910);
nor I_42730 (I728403,I728792,I728910);
or I_42731 (I728406,I728526,I728910);
DFFARX1 I_42732 (I728910,I2507,I728432,I728424,);
not I_42733 (I729010,I2514);
DFFARX1 I_42734 (I482776,I2507,I729010,I729036,);
not I_42735 (I729044,I729036);
nand I_42736 (I729061,I482767,I482785);
and I_42737 (I729078,I729061,I482788);
DFFARX1 I_42738 (I729078,I2507,I729010,I729104,);
not I_42739 (I729112,I482782);
DFFARX1 I_42740 (I482770,I2507,I729010,I729138,);
not I_42741 (I729146,I729138);
nor I_42742 (I729163,I729146,I729044);
and I_42743 (I729180,I729163,I482782);
nor I_42744 (I729197,I729146,I729112);
nor I_42745 (I728993,I729104,I729197);
DFFARX1 I_42746 (I482779,I2507,I729010,I729237,);
nor I_42747 (I729245,I729237,I729104);
not I_42748 (I729262,I729245);
not I_42749 (I729279,I729237);
nor I_42750 (I729296,I729279,I729180);
DFFARX1 I_42751 (I729296,I2507,I729010,I728996,);
nand I_42752 (I729327,I482794,I482791);
and I_42753 (I729344,I729327,I482773);
DFFARX1 I_42754 (I729344,I2507,I729010,I729370,);
nor I_42755 (I729378,I729370,I729237);
DFFARX1 I_42756 (I729378,I2507,I729010,I728978,);
nand I_42757 (I729409,I729370,I729279);
nand I_42758 (I728987,I729262,I729409);
not I_42759 (I729440,I729370);
nor I_42760 (I729457,I729440,I729180);
DFFARX1 I_42761 (I729457,I2507,I729010,I728999,);
nor I_42762 (I729488,I482767,I482791);
or I_42763 (I728990,I729237,I729488);
nor I_42764 (I728981,I729370,I729488);
or I_42765 (I728984,I729104,I729488);
DFFARX1 I_42766 (I729488,I2507,I729010,I729002,);
not I_42767 (I729588,I2514);
DFFARX1 I_42768 (I1225378,I2507,I729588,I729614,);
not I_42769 (I729622,I729614);
nand I_42770 (I729639,I1225381,I1225390);
and I_42771 (I729656,I729639,I1225393);
DFFARX1 I_42772 (I729656,I2507,I729588,I729682,);
not I_42773 (I729690,I1225402);
DFFARX1 I_42774 (I1225384,I2507,I729588,I729716,);
not I_42775 (I729724,I729716);
nor I_42776 (I729741,I729724,I729622);
and I_42777 (I729758,I729741,I1225402);
nor I_42778 (I729775,I729724,I729690);
nor I_42779 (I729571,I729682,I729775);
DFFARX1 I_42780 (I1225381,I2507,I729588,I729815,);
nor I_42781 (I729823,I729815,I729682);
not I_42782 (I729840,I729823);
not I_42783 (I729857,I729815);
nor I_42784 (I729874,I729857,I729758);
DFFARX1 I_42785 (I729874,I2507,I729588,I729574,);
nand I_42786 (I729905,I1225399,I1225378);
and I_42787 (I729922,I729905,I1225396);
DFFARX1 I_42788 (I729922,I2507,I729588,I729948,);
nor I_42789 (I729956,I729948,I729815);
DFFARX1 I_42790 (I729956,I2507,I729588,I729556,);
nand I_42791 (I729987,I729948,I729857);
nand I_42792 (I729565,I729840,I729987);
not I_42793 (I730018,I729948);
nor I_42794 (I730035,I730018,I729758);
DFFARX1 I_42795 (I730035,I2507,I729588,I729577,);
nor I_42796 (I730066,I1225387,I1225378);
or I_42797 (I729568,I729815,I730066);
nor I_42798 (I729559,I729948,I730066);
or I_42799 (I729562,I729682,I730066);
DFFARX1 I_42800 (I730066,I2507,I729588,I729580,);
not I_42801 (I730166,I2514);
DFFARX1 I_42802 (I1146822,I2507,I730166,I730192,);
not I_42803 (I730200,I730192);
nand I_42804 (I730217,I1146804,I1146816);
and I_42805 (I730234,I730217,I1146819);
DFFARX1 I_42806 (I730234,I2507,I730166,I730260,);
not I_42807 (I730268,I1146813);
DFFARX1 I_42808 (I1146810,I2507,I730166,I730294,);
not I_42809 (I730302,I730294);
nor I_42810 (I730319,I730302,I730200);
and I_42811 (I730336,I730319,I1146813);
nor I_42812 (I730353,I730302,I730268);
nor I_42813 (I730149,I730260,I730353);
DFFARX1 I_42814 (I1146828,I2507,I730166,I730393,);
nor I_42815 (I730401,I730393,I730260);
not I_42816 (I730418,I730401);
not I_42817 (I730435,I730393);
nor I_42818 (I730452,I730435,I730336);
DFFARX1 I_42819 (I730452,I2507,I730166,I730152,);
nand I_42820 (I730483,I1146807,I1146807);
and I_42821 (I730500,I730483,I1146804);
DFFARX1 I_42822 (I730500,I2507,I730166,I730526,);
nor I_42823 (I730534,I730526,I730393);
DFFARX1 I_42824 (I730534,I2507,I730166,I730134,);
nand I_42825 (I730565,I730526,I730435);
nand I_42826 (I730143,I730418,I730565);
not I_42827 (I730596,I730526);
nor I_42828 (I730613,I730596,I730336);
DFFARX1 I_42829 (I730613,I2507,I730166,I730155,);
nor I_42830 (I730644,I1146825,I1146807);
or I_42831 (I730146,I730393,I730644);
nor I_42832 (I730137,I730526,I730644);
or I_42833 (I730140,I730260,I730644);
DFFARX1 I_42834 (I730644,I2507,I730166,I730158,);
not I_42835 (I730744,I2514);
DFFARX1 I_42836 (I1172832,I2507,I730744,I730770,);
not I_42837 (I730778,I730770);
nand I_42838 (I730795,I1172814,I1172826);
and I_42839 (I730812,I730795,I1172829);
DFFARX1 I_42840 (I730812,I2507,I730744,I730838,);
not I_42841 (I730846,I1172823);
DFFARX1 I_42842 (I1172820,I2507,I730744,I730872,);
not I_42843 (I730880,I730872);
nor I_42844 (I730897,I730880,I730778);
and I_42845 (I730914,I730897,I1172823);
nor I_42846 (I730931,I730880,I730846);
nor I_42847 (I730727,I730838,I730931);
DFFARX1 I_42848 (I1172838,I2507,I730744,I730971,);
nor I_42849 (I730979,I730971,I730838);
not I_42850 (I730996,I730979);
not I_42851 (I731013,I730971);
nor I_42852 (I731030,I731013,I730914);
DFFARX1 I_42853 (I731030,I2507,I730744,I730730,);
nand I_42854 (I731061,I1172817,I1172817);
and I_42855 (I731078,I731061,I1172814);
DFFARX1 I_42856 (I731078,I2507,I730744,I731104,);
nor I_42857 (I731112,I731104,I730971);
DFFARX1 I_42858 (I731112,I2507,I730744,I730712,);
nand I_42859 (I731143,I731104,I731013);
nand I_42860 (I730721,I730996,I731143);
not I_42861 (I731174,I731104);
nor I_42862 (I731191,I731174,I730914);
DFFARX1 I_42863 (I731191,I2507,I730744,I730733,);
nor I_42864 (I731222,I1172835,I1172817);
or I_42865 (I730724,I730971,I731222);
nor I_42866 (I730715,I731104,I731222);
or I_42867 (I730718,I730838,I731222);
DFFARX1 I_42868 (I731222,I2507,I730744,I730736,);
not I_42869 (I731322,I2514);
DFFARX1 I_42870 (I337696,I2507,I731322,I731348,);
not I_42871 (I731356,I731348);
nand I_42872 (I731373,I337699,I337675);
and I_42873 (I731390,I731373,I337672);
DFFARX1 I_42874 (I731390,I2507,I731322,I731416,);
not I_42875 (I731424,I337678);
DFFARX1 I_42876 (I337672,I2507,I731322,I731450,);
not I_42877 (I731458,I731450);
nor I_42878 (I731475,I731458,I731356);
and I_42879 (I731492,I731475,I337678);
nor I_42880 (I731509,I731458,I731424);
nor I_42881 (I731305,I731416,I731509);
DFFARX1 I_42882 (I337681,I2507,I731322,I731549,);
nor I_42883 (I731557,I731549,I731416);
not I_42884 (I731574,I731557);
not I_42885 (I731591,I731549);
nor I_42886 (I731608,I731591,I731492);
DFFARX1 I_42887 (I731608,I2507,I731322,I731308,);
nand I_42888 (I731639,I337684,I337693);
and I_42889 (I731656,I731639,I337690);
DFFARX1 I_42890 (I731656,I2507,I731322,I731682,);
nor I_42891 (I731690,I731682,I731549);
DFFARX1 I_42892 (I731690,I2507,I731322,I731290,);
nand I_42893 (I731721,I731682,I731591);
nand I_42894 (I731299,I731574,I731721);
not I_42895 (I731752,I731682);
nor I_42896 (I731769,I731752,I731492);
DFFARX1 I_42897 (I731769,I2507,I731322,I731311,);
nor I_42898 (I731800,I337687,I337693);
or I_42899 (I731302,I731549,I731800);
nor I_42900 (I731293,I731682,I731800);
or I_42901 (I731296,I731416,I731800);
DFFARX1 I_42902 (I731800,I2507,I731322,I731314,);
not I_42903 (I731900,I2514);
DFFARX1 I_42904 (I1024733,I2507,I731900,I731926,);
not I_42905 (I731934,I731926);
nand I_42906 (I731951,I1024730,I1024748);
and I_42907 (I731968,I731951,I1024745);
DFFARX1 I_42908 (I731968,I2507,I731900,I731994,);
not I_42909 (I732002,I1024727);
DFFARX1 I_42910 (I1024730,I2507,I731900,I732028,);
not I_42911 (I732036,I732028);
nor I_42912 (I732053,I732036,I731934);
and I_42913 (I732070,I732053,I1024727);
nor I_42914 (I732087,I732036,I732002);
nor I_42915 (I731883,I731994,I732087);
DFFARX1 I_42916 (I1024739,I2507,I731900,I732127,);
nor I_42917 (I732135,I732127,I731994);
not I_42918 (I732152,I732135);
not I_42919 (I732169,I732127);
nor I_42920 (I732186,I732169,I732070);
DFFARX1 I_42921 (I732186,I2507,I731900,I731886,);
nand I_42922 (I732217,I1024742,I1024727);
and I_42923 (I732234,I732217,I1024733);
DFFARX1 I_42924 (I732234,I2507,I731900,I732260,);
nor I_42925 (I732268,I732260,I732127);
DFFARX1 I_42926 (I732268,I2507,I731900,I731868,);
nand I_42927 (I732299,I732260,I732169);
nand I_42928 (I731877,I732152,I732299);
not I_42929 (I732330,I732260);
nor I_42930 (I732347,I732330,I732070);
DFFARX1 I_42931 (I732347,I2507,I731900,I731889,);
nor I_42932 (I732378,I1024736,I1024727);
or I_42933 (I731880,I732127,I732378);
nor I_42934 (I731871,I732260,I732378);
or I_42935 (I731874,I731994,I732378);
DFFARX1 I_42936 (I732378,I2507,I731900,I731892,);
not I_42937 (I732478,I2514);
DFFARX1 I_42938 (I845477,I2507,I732478,I732504,);
not I_42939 (I732512,I732504);
nand I_42940 (I732529,I845465,I845483);
and I_42941 (I732546,I732529,I845480);
DFFARX1 I_42942 (I732546,I2507,I732478,I732572,);
not I_42943 (I732580,I845471);
DFFARX1 I_42944 (I845468,I2507,I732478,I732606,);
not I_42945 (I732614,I732606);
nor I_42946 (I732631,I732614,I732512);
and I_42947 (I732648,I732631,I845471);
nor I_42948 (I732665,I732614,I732580);
nor I_42949 (I732461,I732572,I732665);
DFFARX1 I_42950 (I845462,I2507,I732478,I732705,);
nor I_42951 (I732713,I732705,I732572);
not I_42952 (I732730,I732713);
not I_42953 (I732747,I732705);
nor I_42954 (I732764,I732747,I732648);
DFFARX1 I_42955 (I732764,I2507,I732478,I732464,);
nand I_42956 (I732795,I845462,I845465);
and I_42957 (I732812,I732795,I845468);
DFFARX1 I_42958 (I732812,I2507,I732478,I732838,);
nor I_42959 (I732846,I732838,I732705);
DFFARX1 I_42960 (I732846,I2507,I732478,I732446,);
nand I_42961 (I732877,I732838,I732747);
nand I_42962 (I732455,I732730,I732877);
not I_42963 (I732908,I732838);
nor I_42964 (I732925,I732908,I732648);
DFFARX1 I_42965 (I732925,I2507,I732478,I732467,);
nor I_42966 (I732956,I845474,I845465);
or I_42967 (I732458,I732705,I732956);
nor I_42968 (I732449,I732838,I732956);
or I_42969 (I732452,I732572,I732956);
DFFARX1 I_42970 (I732956,I2507,I732478,I732470,);
not I_42971 (I733056,I2514);
DFFARX1 I_42972 (I1142198,I2507,I733056,I733082,);
not I_42973 (I733090,I733082);
nand I_42974 (I733107,I1142180,I1142192);
and I_42975 (I733124,I733107,I1142195);
DFFARX1 I_42976 (I733124,I2507,I733056,I733150,);
not I_42977 (I733158,I1142189);
DFFARX1 I_42978 (I1142186,I2507,I733056,I733184,);
not I_42979 (I733192,I733184);
nor I_42980 (I733209,I733192,I733090);
and I_42981 (I733226,I733209,I1142189);
nor I_42982 (I733243,I733192,I733158);
nor I_42983 (I733039,I733150,I733243);
DFFARX1 I_42984 (I1142204,I2507,I733056,I733283,);
nor I_42985 (I733291,I733283,I733150);
not I_42986 (I733308,I733291);
not I_42987 (I733325,I733283);
nor I_42988 (I733342,I733325,I733226);
DFFARX1 I_42989 (I733342,I2507,I733056,I733042,);
nand I_42990 (I733373,I1142183,I1142183);
and I_42991 (I733390,I733373,I1142180);
DFFARX1 I_42992 (I733390,I2507,I733056,I733416,);
nor I_42993 (I733424,I733416,I733283);
DFFARX1 I_42994 (I733424,I2507,I733056,I733024,);
nand I_42995 (I733455,I733416,I733325);
nand I_42996 (I733033,I733308,I733455);
not I_42997 (I733486,I733416);
nor I_42998 (I733503,I733486,I733226);
DFFARX1 I_42999 (I733503,I2507,I733056,I733045,);
nor I_43000 (I733534,I1142201,I1142183);
or I_43001 (I733036,I733283,I733534);
nor I_43002 (I733027,I733416,I733534);
or I_43003 (I733030,I733150,I733534);
DFFARX1 I_43004 (I733534,I2507,I733056,I733048,);
not I_43005 (I733634,I2514);
DFFARX1 I_43006 (I1309504,I2507,I733634,I733660,);
not I_43007 (I733668,I733660);
nand I_43008 (I733685,I1309489,I1309477);
and I_43009 (I733702,I733685,I1309492);
DFFARX1 I_43010 (I733702,I2507,I733634,I733728,);
not I_43011 (I733736,I1309477);
DFFARX1 I_43012 (I1309495,I2507,I733634,I733762,);
not I_43013 (I733770,I733762);
nor I_43014 (I733787,I733770,I733668);
and I_43015 (I733804,I733787,I1309477);
nor I_43016 (I733821,I733770,I733736);
nor I_43017 (I733617,I733728,I733821);
DFFARX1 I_43018 (I1309483,I2507,I733634,I733861,);
nor I_43019 (I733869,I733861,I733728);
not I_43020 (I733886,I733869);
not I_43021 (I733903,I733861);
nor I_43022 (I733920,I733903,I733804);
DFFARX1 I_43023 (I733920,I2507,I733634,I733620,);
nand I_43024 (I733951,I1309480,I1309486);
and I_43025 (I733968,I733951,I1309501);
DFFARX1 I_43026 (I733968,I2507,I733634,I733994,);
nor I_43027 (I734002,I733994,I733861);
DFFARX1 I_43028 (I734002,I2507,I733634,I733602,);
nand I_43029 (I734033,I733994,I733903);
nand I_43030 (I733611,I733886,I734033);
not I_43031 (I734064,I733994);
nor I_43032 (I734081,I734064,I733804);
DFFARX1 I_43033 (I734081,I2507,I733634,I733623,);
nor I_43034 (I734112,I1309498,I1309486);
or I_43035 (I733614,I733861,I734112);
nor I_43036 (I733605,I733994,I734112);
or I_43037 (I733608,I733728,I734112);
DFFARX1 I_43038 (I734112,I2507,I733634,I733626,);
not I_43039 (I734212,I2514);
DFFARX1 I_43040 (I287104,I2507,I734212,I734238,);
not I_43041 (I734246,I734238);
nand I_43042 (I734263,I287107,I287083);
and I_43043 (I734280,I734263,I287080);
DFFARX1 I_43044 (I734280,I2507,I734212,I734306,);
not I_43045 (I734314,I287086);
DFFARX1 I_43046 (I287080,I2507,I734212,I734340,);
not I_43047 (I734348,I734340);
nor I_43048 (I734365,I734348,I734246);
and I_43049 (I734382,I734365,I287086);
nor I_43050 (I734399,I734348,I734314);
nor I_43051 (I734195,I734306,I734399);
DFFARX1 I_43052 (I287089,I2507,I734212,I734439,);
nor I_43053 (I734447,I734439,I734306);
not I_43054 (I734464,I734447);
not I_43055 (I734481,I734439);
nor I_43056 (I734498,I734481,I734382);
DFFARX1 I_43057 (I734498,I2507,I734212,I734198,);
nand I_43058 (I734529,I287092,I287101);
and I_43059 (I734546,I734529,I287098);
DFFARX1 I_43060 (I734546,I2507,I734212,I734572,);
nor I_43061 (I734580,I734572,I734439);
DFFARX1 I_43062 (I734580,I2507,I734212,I734180,);
nand I_43063 (I734611,I734572,I734481);
nand I_43064 (I734189,I734464,I734611);
not I_43065 (I734642,I734572);
nor I_43066 (I734659,I734642,I734382);
DFFARX1 I_43067 (I734659,I2507,I734212,I734201,);
nor I_43068 (I734690,I287095,I287101);
or I_43069 (I734192,I734439,I734690);
nor I_43070 (I734183,I734572,I734690);
or I_43071 (I734186,I734306,I734690);
DFFARX1 I_43072 (I734690,I2507,I734212,I734204,);
not I_43073 (I734790,I2514);
DFFARX1 I_43074 (I247215,I2507,I734790,I734816,);
not I_43075 (I734824,I734816);
nand I_43076 (I734841,I247218,I247239);
and I_43077 (I734858,I734841,I247227);
DFFARX1 I_43078 (I734858,I2507,I734790,I734884,);
not I_43079 (I734892,I247224);
DFFARX1 I_43080 (I247215,I2507,I734790,I734918,);
not I_43081 (I734926,I734918);
nor I_43082 (I734943,I734926,I734824);
and I_43083 (I734960,I734943,I247224);
nor I_43084 (I734977,I734926,I734892);
nor I_43085 (I734773,I734884,I734977);
DFFARX1 I_43086 (I247233,I2507,I734790,I735017,);
nor I_43087 (I735025,I735017,I734884);
not I_43088 (I735042,I735025);
not I_43089 (I735059,I735017);
nor I_43090 (I735076,I735059,I734960);
DFFARX1 I_43091 (I735076,I2507,I734790,I734776,);
nand I_43092 (I735107,I247218,I247221);
and I_43093 (I735124,I735107,I247230);
DFFARX1 I_43094 (I735124,I2507,I734790,I735150,);
nor I_43095 (I735158,I735150,I735017);
DFFARX1 I_43096 (I735158,I2507,I734790,I734758,);
nand I_43097 (I735189,I735150,I735059);
nand I_43098 (I734767,I735042,I735189);
not I_43099 (I735220,I735150);
nor I_43100 (I735237,I735220,I734960);
DFFARX1 I_43101 (I735237,I2507,I734790,I734779,);
nor I_43102 (I735268,I247236,I247221);
or I_43103 (I734770,I735017,I735268);
nor I_43104 (I734761,I735150,I735268);
or I_43105 (I734764,I734884,I735268);
DFFARX1 I_43106 (I735268,I2507,I734790,I734782,);
not I_43107 (I735368,I2514);
DFFARX1 I_43108 (I1229186,I2507,I735368,I735394,);
not I_43109 (I735402,I735394);
nand I_43110 (I735419,I1229189,I1229198);
and I_43111 (I735436,I735419,I1229201);
DFFARX1 I_43112 (I735436,I2507,I735368,I735462,);
not I_43113 (I735470,I1229210);
DFFARX1 I_43114 (I1229192,I2507,I735368,I735496,);
not I_43115 (I735504,I735496);
nor I_43116 (I735521,I735504,I735402);
and I_43117 (I735538,I735521,I1229210);
nor I_43118 (I735555,I735504,I735470);
nor I_43119 (I735351,I735462,I735555);
DFFARX1 I_43120 (I1229189,I2507,I735368,I735595,);
nor I_43121 (I735603,I735595,I735462);
not I_43122 (I735620,I735603);
not I_43123 (I735637,I735595);
nor I_43124 (I735654,I735637,I735538);
DFFARX1 I_43125 (I735654,I2507,I735368,I735354,);
nand I_43126 (I735685,I1229207,I1229186);
and I_43127 (I735702,I735685,I1229204);
DFFARX1 I_43128 (I735702,I2507,I735368,I735728,);
nor I_43129 (I735736,I735728,I735595);
DFFARX1 I_43130 (I735736,I2507,I735368,I735336,);
nand I_43131 (I735767,I735728,I735637);
nand I_43132 (I735345,I735620,I735767);
not I_43133 (I735798,I735728);
nor I_43134 (I735815,I735798,I735538);
DFFARX1 I_43135 (I735815,I2507,I735368,I735357,);
nor I_43136 (I735846,I1229195,I1229186);
or I_43137 (I735348,I735595,I735846);
nor I_43138 (I735339,I735728,I735846);
or I_43139 (I735342,I735462,I735846);
DFFARX1 I_43140 (I735846,I2507,I735368,I735360,);
not I_43141 (I735946,I2514);
DFFARX1 I_43142 (I424568,I2507,I735946,I735972,);
not I_43143 (I735980,I735972);
nand I_43144 (I735997,I424559,I424577);
and I_43145 (I736014,I735997,I424580);
DFFARX1 I_43146 (I736014,I2507,I735946,I736040,);
not I_43147 (I736048,I424574);
DFFARX1 I_43148 (I424562,I2507,I735946,I736074,);
not I_43149 (I736082,I736074);
nor I_43150 (I736099,I736082,I735980);
and I_43151 (I736116,I736099,I424574);
nor I_43152 (I736133,I736082,I736048);
nor I_43153 (I735929,I736040,I736133);
DFFARX1 I_43154 (I424571,I2507,I735946,I736173,);
nor I_43155 (I736181,I736173,I736040);
not I_43156 (I736198,I736181);
not I_43157 (I736215,I736173);
nor I_43158 (I736232,I736215,I736116);
DFFARX1 I_43159 (I736232,I2507,I735946,I735932,);
nand I_43160 (I736263,I424586,I424583);
and I_43161 (I736280,I736263,I424565);
DFFARX1 I_43162 (I736280,I2507,I735946,I736306,);
nor I_43163 (I736314,I736306,I736173);
DFFARX1 I_43164 (I736314,I2507,I735946,I735914,);
nand I_43165 (I736345,I736306,I736215);
nand I_43166 (I735923,I736198,I736345);
not I_43167 (I736376,I736306);
nor I_43168 (I736393,I736376,I736116);
DFFARX1 I_43169 (I736393,I2507,I735946,I735935,);
nor I_43170 (I736424,I424559,I424583);
or I_43171 (I735926,I736173,I736424);
nor I_43172 (I735917,I736306,I736424);
or I_43173 (I735920,I736040,I736424);
DFFARX1 I_43174 (I736424,I2507,I735946,I735938,);
not I_43175 (I736524,I2514);
DFFARX1 I_43176 (I472984,I2507,I736524,I736550,);
not I_43177 (I736558,I736550);
nand I_43178 (I736575,I472975,I472993);
and I_43179 (I736592,I736575,I472996);
DFFARX1 I_43180 (I736592,I2507,I736524,I736618,);
not I_43181 (I736626,I472990);
DFFARX1 I_43182 (I472978,I2507,I736524,I736652,);
not I_43183 (I736660,I736652);
nor I_43184 (I736677,I736660,I736558);
and I_43185 (I736694,I736677,I472990);
nor I_43186 (I736711,I736660,I736626);
nor I_43187 (I736507,I736618,I736711);
DFFARX1 I_43188 (I472987,I2507,I736524,I736751,);
nor I_43189 (I736759,I736751,I736618);
not I_43190 (I736776,I736759);
not I_43191 (I736793,I736751);
nor I_43192 (I736810,I736793,I736694);
DFFARX1 I_43193 (I736810,I2507,I736524,I736510,);
nand I_43194 (I736841,I473002,I472999);
and I_43195 (I736858,I736841,I472981);
DFFARX1 I_43196 (I736858,I2507,I736524,I736884,);
nor I_43197 (I736892,I736884,I736751);
DFFARX1 I_43198 (I736892,I2507,I736524,I736492,);
nand I_43199 (I736923,I736884,I736793);
nand I_43200 (I736501,I736776,I736923);
not I_43201 (I736954,I736884);
nor I_43202 (I736971,I736954,I736694);
DFFARX1 I_43203 (I736971,I2507,I736524,I736513,);
nor I_43204 (I737002,I472975,I472999);
or I_43205 (I736504,I736751,I737002);
nor I_43206 (I736495,I736884,I737002);
or I_43207 (I736498,I736618,I737002);
DFFARX1 I_43208 (I737002,I2507,I736524,I736516,);
not I_43209 (I737102,I2514);
DFFARX1 I_43210 (I940567,I2507,I737102,I737128,);
not I_43211 (I737136,I737128);
nand I_43212 (I737153,I940543,I940558);
and I_43213 (I737170,I737153,I940570);
DFFARX1 I_43214 (I737170,I2507,I737102,I737196,);
not I_43215 (I737204,I940555);
DFFARX1 I_43216 (I940546,I2507,I737102,I737230,);
not I_43217 (I737238,I737230);
nor I_43218 (I737255,I737238,I737136);
and I_43219 (I737272,I737255,I940555);
nor I_43220 (I737289,I737238,I737204);
nor I_43221 (I737085,I737196,I737289);
DFFARX1 I_43222 (I940543,I2507,I737102,I737329,);
nor I_43223 (I737337,I737329,I737196);
not I_43224 (I737354,I737337);
not I_43225 (I737371,I737329);
nor I_43226 (I737388,I737371,I737272);
DFFARX1 I_43227 (I737388,I2507,I737102,I737088,);
nand I_43228 (I737419,I940561,I940552);
and I_43229 (I737436,I737419,I940564);
DFFARX1 I_43230 (I737436,I2507,I737102,I737462,);
nor I_43231 (I737470,I737462,I737329);
DFFARX1 I_43232 (I737470,I2507,I737102,I737070,);
nand I_43233 (I737501,I737462,I737371);
nand I_43234 (I737079,I737354,I737501);
not I_43235 (I737532,I737462);
nor I_43236 (I737549,I737532,I737272);
DFFARX1 I_43237 (I737549,I2507,I737102,I737091,);
nor I_43238 (I737580,I940549,I940552);
or I_43239 (I737082,I737329,I737580);
nor I_43240 (I737073,I737462,I737580);
or I_43241 (I737076,I737196,I737580);
DFFARX1 I_43242 (I737580,I2507,I737102,I737094,);
not I_43243 (I737680,I2514);
DFFARX1 I_43244 (I4903,I2507,I737680,I737706,);
not I_43245 (I737714,I737706);
nand I_43246 (I737731,I4906,I4918);
and I_43247 (I737748,I737731,I4897);
DFFARX1 I_43248 (I737748,I2507,I737680,I737774,);
not I_43249 (I737782,I4897);
DFFARX1 I_43250 (I4900,I2507,I737680,I737808,);
not I_43251 (I737816,I737808);
nor I_43252 (I737833,I737816,I737714);
and I_43253 (I737850,I737833,I4897);
nor I_43254 (I737867,I737816,I737782);
nor I_43255 (I737663,I737774,I737867);
DFFARX1 I_43256 (I4912,I2507,I737680,I737907,);
nor I_43257 (I737915,I737907,I737774);
not I_43258 (I737932,I737915);
not I_43259 (I737949,I737907);
nor I_43260 (I737966,I737949,I737850);
DFFARX1 I_43261 (I737966,I2507,I737680,I737666,);
nand I_43262 (I737997,I4915,I4900);
and I_43263 (I738014,I737997,I4909);
DFFARX1 I_43264 (I738014,I2507,I737680,I738040,);
nor I_43265 (I738048,I738040,I737907);
DFFARX1 I_43266 (I738048,I2507,I737680,I737648,);
nand I_43267 (I738079,I738040,I737949);
nand I_43268 (I737657,I737932,I738079);
not I_43269 (I738110,I738040);
nor I_43270 (I738127,I738110,I737850);
DFFARX1 I_43271 (I738127,I2507,I737680,I737669,);
nor I_43272 (I738158,I4903,I4900);
or I_43273 (I737660,I737907,I738158);
nor I_43274 (I737651,I738040,I738158);
or I_43275 (I737654,I737774,I738158);
DFFARX1 I_43276 (I738158,I2507,I737680,I737672,);
not I_43277 (I738258,I2514);
DFFARX1 I_43278 (I404440,I2507,I738258,I738284,);
not I_43279 (I738292,I738284);
nand I_43280 (I738309,I404431,I404449);
and I_43281 (I738326,I738309,I404452);
DFFARX1 I_43282 (I738326,I2507,I738258,I738352,);
not I_43283 (I738360,I404446);
DFFARX1 I_43284 (I404434,I2507,I738258,I738386,);
not I_43285 (I738394,I738386);
nor I_43286 (I738411,I738394,I738292);
and I_43287 (I738428,I738411,I404446);
nor I_43288 (I738445,I738394,I738360);
nor I_43289 (I738241,I738352,I738445);
DFFARX1 I_43290 (I404443,I2507,I738258,I738485,);
nor I_43291 (I738493,I738485,I738352);
not I_43292 (I738510,I738493);
not I_43293 (I738527,I738485);
nor I_43294 (I738544,I738527,I738428);
DFFARX1 I_43295 (I738544,I2507,I738258,I738244,);
nand I_43296 (I738575,I404458,I404455);
and I_43297 (I738592,I738575,I404437);
DFFARX1 I_43298 (I738592,I2507,I738258,I738618,);
nor I_43299 (I738626,I738618,I738485);
DFFARX1 I_43300 (I738626,I2507,I738258,I738226,);
nand I_43301 (I738657,I738618,I738527);
nand I_43302 (I738235,I738510,I738657);
not I_43303 (I738688,I738618);
nor I_43304 (I738705,I738688,I738428);
DFFARX1 I_43305 (I738705,I2507,I738258,I738247,);
nor I_43306 (I738736,I404431,I404455);
or I_43307 (I738238,I738485,I738736);
nor I_43308 (I738229,I738618,I738736);
or I_43309 (I738232,I738352,I738736);
DFFARX1 I_43310 (I738736,I2507,I738258,I738250,);
not I_43311 (I738836,I2514);
DFFARX1 I_43312 (I841788,I2507,I738836,I738862,);
not I_43313 (I738870,I738862);
nand I_43314 (I738887,I841776,I841794);
and I_43315 (I738904,I738887,I841791);
DFFARX1 I_43316 (I738904,I2507,I738836,I738930,);
not I_43317 (I738938,I841782);
DFFARX1 I_43318 (I841779,I2507,I738836,I738964,);
not I_43319 (I738972,I738964);
nor I_43320 (I738989,I738972,I738870);
and I_43321 (I739006,I738989,I841782);
nor I_43322 (I739023,I738972,I738938);
nor I_43323 (I738819,I738930,I739023);
DFFARX1 I_43324 (I841773,I2507,I738836,I739063,);
nor I_43325 (I739071,I739063,I738930);
not I_43326 (I739088,I739071);
not I_43327 (I739105,I739063);
nor I_43328 (I739122,I739105,I739006);
DFFARX1 I_43329 (I739122,I2507,I738836,I738822,);
nand I_43330 (I739153,I841773,I841776);
and I_43331 (I739170,I739153,I841779);
DFFARX1 I_43332 (I739170,I2507,I738836,I739196,);
nor I_43333 (I739204,I739196,I739063);
DFFARX1 I_43334 (I739204,I2507,I738836,I738804,);
nand I_43335 (I739235,I739196,I739105);
nand I_43336 (I738813,I739088,I739235);
not I_43337 (I739266,I739196);
nor I_43338 (I739283,I739266,I739006);
DFFARX1 I_43339 (I739283,I2507,I738836,I738825,);
nor I_43340 (I739314,I841785,I841776);
or I_43341 (I738816,I739063,I739314);
nor I_43342 (I738807,I739196,I739314);
or I_43343 (I738810,I738930,I739314);
DFFARX1 I_43344 (I739314,I2507,I738836,I738828,);
not I_43345 (I739414,I2514);
DFFARX1 I_43346 (I183550,I2507,I739414,I739440,);
not I_43347 (I739448,I739440);
nand I_43348 (I739465,I183553,I183574);
and I_43349 (I739482,I739465,I183562);
DFFARX1 I_43350 (I739482,I2507,I739414,I739508,);
not I_43351 (I739516,I183559);
DFFARX1 I_43352 (I183550,I2507,I739414,I739542,);
not I_43353 (I739550,I739542);
nor I_43354 (I739567,I739550,I739448);
and I_43355 (I739584,I739567,I183559);
nor I_43356 (I739601,I739550,I739516);
nor I_43357 (I739397,I739508,I739601);
DFFARX1 I_43358 (I183568,I2507,I739414,I739641,);
nor I_43359 (I739649,I739641,I739508);
not I_43360 (I739666,I739649);
not I_43361 (I739683,I739641);
nor I_43362 (I739700,I739683,I739584);
DFFARX1 I_43363 (I739700,I2507,I739414,I739400,);
nand I_43364 (I739731,I183553,I183556);
and I_43365 (I739748,I739731,I183565);
DFFARX1 I_43366 (I739748,I2507,I739414,I739774,);
nor I_43367 (I739782,I739774,I739641);
DFFARX1 I_43368 (I739782,I2507,I739414,I739382,);
nand I_43369 (I739813,I739774,I739683);
nand I_43370 (I739391,I739666,I739813);
not I_43371 (I739844,I739774);
nor I_43372 (I739861,I739844,I739584);
DFFARX1 I_43373 (I739861,I2507,I739414,I739403,);
nor I_43374 (I739892,I183571,I183556);
or I_43375 (I739394,I739641,I739892);
nor I_43376 (I739385,I739774,I739892);
or I_43377 (I739388,I739508,I739892);
DFFARX1 I_43378 (I739892,I2507,I739414,I739406,);
not I_43379 (I739992,I2514);
DFFARX1 I_43380 (I587946,I2507,I739992,I740018,);
not I_43381 (I740026,I740018);
nand I_43382 (I740043,I587955,I587964);
and I_43383 (I740060,I740043,I587970);
DFFARX1 I_43384 (I740060,I2507,I739992,I740086,);
not I_43385 (I740094,I587967);
DFFARX1 I_43386 (I587952,I2507,I739992,I740120,);
not I_43387 (I740128,I740120);
nor I_43388 (I740145,I740128,I740026);
and I_43389 (I740162,I740145,I587967);
nor I_43390 (I740179,I740128,I740094);
nor I_43391 (I739975,I740086,I740179);
DFFARX1 I_43392 (I587961,I2507,I739992,I740219,);
nor I_43393 (I740227,I740219,I740086);
not I_43394 (I740244,I740227);
not I_43395 (I740261,I740219);
nor I_43396 (I740278,I740261,I740162);
DFFARX1 I_43397 (I740278,I2507,I739992,I739978,);
nand I_43398 (I740309,I587958,I587949);
and I_43399 (I740326,I740309,I587946);
DFFARX1 I_43400 (I740326,I2507,I739992,I740352,);
nor I_43401 (I740360,I740352,I740219);
DFFARX1 I_43402 (I740360,I2507,I739992,I739960,);
nand I_43403 (I740391,I740352,I740261);
nand I_43404 (I739969,I740244,I740391);
not I_43405 (I740422,I740352);
nor I_43406 (I740439,I740422,I740162);
DFFARX1 I_43407 (I740439,I2507,I739992,I739981,);
nor I_43408 (I740470,I587949,I587949);
or I_43409 (I739972,I740219,I740470);
nor I_43410 (I739963,I740352,I740470);
or I_43411 (I739966,I740086,I740470);
DFFARX1 I_43412 (I740470,I2507,I739992,I739984,);
not I_43413 (I740570,I2514);
DFFARX1 I_43414 (I1382689,I2507,I740570,I740596,);
not I_43415 (I740604,I740596);
nand I_43416 (I740621,I1382674,I1382662);
and I_43417 (I740638,I740621,I1382677);
DFFARX1 I_43418 (I740638,I2507,I740570,I740664,);
not I_43419 (I740672,I1382662);
DFFARX1 I_43420 (I1382680,I2507,I740570,I740698,);
not I_43421 (I740706,I740698);
nor I_43422 (I740723,I740706,I740604);
and I_43423 (I740740,I740723,I1382662);
nor I_43424 (I740757,I740706,I740672);
nor I_43425 (I740553,I740664,I740757);
DFFARX1 I_43426 (I1382668,I2507,I740570,I740797,);
nor I_43427 (I740805,I740797,I740664);
not I_43428 (I740822,I740805);
not I_43429 (I740839,I740797);
nor I_43430 (I740856,I740839,I740740);
DFFARX1 I_43431 (I740856,I2507,I740570,I740556,);
nand I_43432 (I740887,I1382665,I1382671);
and I_43433 (I740904,I740887,I1382686);
DFFARX1 I_43434 (I740904,I2507,I740570,I740930,);
nor I_43435 (I740938,I740930,I740797);
DFFARX1 I_43436 (I740938,I2507,I740570,I740538,);
nand I_43437 (I740969,I740930,I740839);
nand I_43438 (I740547,I740822,I740969);
not I_43439 (I741000,I740930);
nor I_43440 (I741017,I741000,I740740);
DFFARX1 I_43441 (I741017,I2507,I740570,I740559,);
nor I_43442 (I741048,I1382683,I1382671);
or I_43443 (I740550,I740797,I741048);
nor I_43444 (I740541,I740930,I741048);
or I_43445 (I740544,I740664,I741048);
DFFARX1 I_43446 (I741048,I2507,I740570,I740562,);
not I_43447 (I741148,I2514);
DFFARX1 I_43448 (I933461,I2507,I741148,I741174,);
not I_43449 (I741182,I741174);
nand I_43450 (I741199,I933437,I933452);
and I_43451 (I741216,I741199,I933464);
DFFARX1 I_43452 (I741216,I2507,I741148,I741242,);
not I_43453 (I741250,I933449);
DFFARX1 I_43454 (I933440,I2507,I741148,I741276,);
not I_43455 (I741284,I741276);
nor I_43456 (I741301,I741284,I741182);
and I_43457 (I741318,I741301,I933449);
nor I_43458 (I741335,I741284,I741250);
nor I_43459 (I741131,I741242,I741335);
DFFARX1 I_43460 (I933437,I2507,I741148,I741375,);
nor I_43461 (I741383,I741375,I741242);
not I_43462 (I741400,I741383);
not I_43463 (I741417,I741375);
nor I_43464 (I741434,I741417,I741318);
DFFARX1 I_43465 (I741434,I2507,I741148,I741134,);
nand I_43466 (I741465,I933455,I933446);
and I_43467 (I741482,I741465,I933458);
DFFARX1 I_43468 (I741482,I2507,I741148,I741508,);
nor I_43469 (I741516,I741508,I741375);
DFFARX1 I_43470 (I741516,I2507,I741148,I741116,);
nand I_43471 (I741547,I741508,I741417);
nand I_43472 (I741125,I741400,I741547);
not I_43473 (I741578,I741508);
nor I_43474 (I741595,I741578,I741318);
DFFARX1 I_43475 (I741595,I2507,I741148,I741137,);
nor I_43476 (I741626,I933443,I933446);
or I_43477 (I741128,I741375,I741626);
nor I_43478 (I741119,I741508,I741626);
or I_43479 (I741122,I741242,I741626);
DFFARX1 I_43480 (I741626,I2507,I741148,I741140,);
not I_43481 (I741726,I2514);
DFFARX1 I_43482 (I486584,I2507,I741726,I741752,);
not I_43483 (I741760,I741752);
nand I_43484 (I741777,I486575,I486593);
and I_43485 (I741794,I741777,I486596);
DFFARX1 I_43486 (I741794,I2507,I741726,I741820,);
not I_43487 (I741828,I486590);
DFFARX1 I_43488 (I486578,I2507,I741726,I741854,);
not I_43489 (I741862,I741854);
nor I_43490 (I741879,I741862,I741760);
and I_43491 (I741896,I741879,I486590);
nor I_43492 (I741913,I741862,I741828);
nor I_43493 (I741709,I741820,I741913);
DFFARX1 I_43494 (I486587,I2507,I741726,I741953,);
nor I_43495 (I741961,I741953,I741820);
not I_43496 (I741978,I741961);
not I_43497 (I741995,I741953);
nor I_43498 (I742012,I741995,I741896);
DFFARX1 I_43499 (I742012,I2507,I741726,I741712,);
nand I_43500 (I742043,I486602,I486599);
and I_43501 (I742060,I742043,I486581);
DFFARX1 I_43502 (I742060,I2507,I741726,I742086,);
nor I_43503 (I742094,I742086,I741953);
DFFARX1 I_43504 (I742094,I2507,I741726,I741694,);
nand I_43505 (I742125,I742086,I741995);
nand I_43506 (I741703,I741978,I742125);
not I_43507 (I742156,I742086);
nor I_43508 (I742173,I742156,I741896);
DFFARX1 I_43509 (I742173,I2507,I741726,I741715,);
nor I_43510 (I742204,I486575,I486599);
or I_43511 (I741706,I741953,I742204);
nor I_43512 (I741697,I742086,I742204);
or I_43513 (I741700,I741820,I742204);
DFFARX1 I_43514 (I742204,I2507,I741726,I741718,);
not I_43515 (I742304,I2514);
DFFARX1 I_43516 (I298698,I2507,I742304,I742330,);
not I_43517 (I742338,I742330);
nand I_43518 (I742355,I298701,I298677);
and I_43519 (I742372,I742355,I298674);
DFFARX1 I_43520 (I742372,I2507,I742304,I742398,);
not I_43521 (I742406,I298680);
DFFARX1 I_43522 (I298674,I2507,I742304,I742432,);
not I_43523 (I742440,I742432);
nor I_43524 (I742457,I742440,I742338);
and I_43525 (I742474,I742457,I298680);
nor I_43526 (I742491,I742440,I742406);
nor I_43527 (I742287,I742398,I742491);
DFFARX1 I_43528 (I298683,I2507,I742304,I742531,);
nor I_43529 (I742539,I742531,I742398);
not I_43530 (I742556,I742539);
not I_43531 (I742573,I742531);
nor I_43532 (I742590,I742573,I742474);
DFFARX1 I_43533 (I742590,I2507,I742304,I742290,);
nand I_43534 (I742621,I298686,I298695);
and I_43535 (I742638,I742621,I298692);
DFFARX1 I_43536 (I742638,I2507,I742304,I742664,);
nor I_43537 (I742672,I742664,I742531);
DFFARX1 I_43538 (I742672,I2507,I742304,I742272,);
nand I_43539 (I742703,I742664,I742573);
nand I_43540 (I742281,I742556,I742703);
not I_43541 (I742734,I742664);
nor I_43542 (I742751,I742734,I742474);
DFFARX1 I_43543 (I742751,I2507,I742304,I742293,);
nor I_43544 (I742782,I298689,I298695);
or I_43545 (I742284,I742531,I742782);
nor I_43546 (I742275,I742664,I742782);
or I_43547 (I742278,I742398,I742782);
DFFARX1 I_43548 (I742782,I2507,I742304,I742296,);
not I_43549 (I742882,I2514);
DFFARX1 I_43550 (I1156070,I2507,I742882,I742908,);
not I_43551 (I742916,I742908);
nand I_43552 (I742933,I1156052,I1156064);
and I_43553 (I742950,I742933,I1156067);
DFFARX1 I_43554 (I742950,I2507,I742882,I742976,);
not I_43555 (I742984,I1156061);
DFFARX1 I_43556 (I1156058,I2507,I742882,I743010,);
not I_43557 (I743018,I743010);
nor I_43558 (I743035,I743018,I742916);
and I_43559 (I743052,I743035,I1156061);
nor I_43560 (I743069,I743018,I742984);
nor I_43561 (I742865,I742976,I743069);
DFFARX1 I_43562 (I1156076,I2507,I742882,I743109,);
nor I_43563 (I743117,I743109,I742976);
not I_43564 (I743134,I743117);
not I_43565 (I743151,I743109);
nor I_43566 (I743168,I743151,I743052);
DFFARX1 I_43567 (I743168,I2507,I742882,I742868,);
nand I_43568 (I743199,I1156055,I1156055);
and I_43569 (I743216,I743199,I1156052);
DFFARX1 I_43570 (I743216,I2507,I742882,I743242,);
nor I_43571 (I743250,I743242,I743109);
DFFARX1 I_43572 (I743250,I2507,I742882,I742850,);
nand I_43573 (I743281,I743242,I743151);
nand I_43574 (I742859,I743134,I743281);
not I_43575 (I743312,I743242);
nor I_43576 (I743329,I743312,I743052);
DFFARX1 I_43577 (I743329,I2507,I742882,I742871,);
nor I_43578 (I743360,I1156073,I1156055);
or I_43579 (I742862,I743109,I743360);
nor I_43580 (I742853,I743242,I743360);
or I_43581 (I742856,I742976,I743360);
DFFARX1 I_43582 (I743360,I2507,I742882,I742874,);
not I_43583 (I743460,I2514);
DFFARX1 I_43584 (I428920,I2507,I743460,I743486,);
not I_43585 (I743494,I743486);
nand I_43586 (I743511,I428911,I428929);
and I_43587 (I743528,I743511,I428932);
DFFARX1 I_43588 (I743528,I2507,I743460,I743554,);
not I_43589 (I743562,I428926);
DFFARX1 I_43590 (I428914,I2507,I743460,I743588,);
not I_43591 (I743596,I743588);
nor I_43592 (I743613,I743596,I743494);
and I_43593 (I743630,I743613,I428926);
nor I_43594 (I743647,I743596,I743562);
nor I_43595 (I743443,I743554,I743647);
DFFARX1 I_43596 (I428923,I2507,I743460,I743687,);
nor I_43597 (I743695,I743687,I743554);
not I_43598 (I743712,I743695);
not I_43599 (I743729,I743687);
nor I_43600 (I743746,I743729,I743630);
DFFARX1 I_43601 (I743746,I2507,I743460,I743446,);
nand I_43602 (I743777,I428938,I428935);
and I_43603 (I743794,I743777,I428917);
DFFARX1 I_43604 (I743794,I2507,I743460,I743820,);
nor I_43605 (I743828,I743820,I743687);
DFFARX1 I_43606 (I743828,I2507,I743460,I743428,);
nand I_43607 (I743859,I743820,I743729);
nand I_43608 (I743437,I743712,I743859);
not I_43609 (I743890,I743820);
nor I_43610 (I743907,I743890,I743630);
DFFARX1 I_43611 (I743907,I2507,I743460,I743449,);
nor I_43612 (I743938,I428911,I428935);
or I_43613 (I743440,I743687,I743938);
nor I_43614 (I743431,I743820,I743938);
or I_43615 (I743434,I743554,I743938);
DFFARX1 I_43616 (I743938,I2507,I743460,I743452,);
not I_43617 (I744038,I2514);
DFFARX1 I_43618 (I58025,I2507,I744038,I744064,);
not I_43619 (I744072,I744064);
nand I_43620 (I744089,I58034,I58043);
and I_43621 (I744106,I744089,I58022);
DFFARX1 I_43622 (I744106,I2507,I744038,I744132,);
not I_43623 (I744140,I58025);
DFFARX1 I_43624 (I58040,I2507,I744038,I744166,);
not I_43625 (I744174,I744166);
nor I_43626 (I744191,I744174,I744072);
and I_43627 (I744208,I744191,I58025);
nor I_43628 (I744225,I744174,I744140);
nor I_43629 (I744021,I744132,I744225);
DFFARX1 I_43630 (I58031,I2507,I744038,I744265,);
nor I_43631 (I744273,I744265,I744132);
not I_43632 (I744290,I744273);
not I_43633 (I744307,I744265);
nor I_43634 (I744324,I744307,I744208);
DFFARX1 I_43635 (I744324,I2507,I744038,I744024,);
nand I_43636 (I744355,I58046,I58022);
and I_43637 (I744372,I744355,I58028);
DFFARX1 I_43638 (I744372,I2507,I744038,I744398,);
nor I_43639 (I744406,I744398,I744265);
DFFARX1 I_43640 (I744406,I2507,I744038,I744006,);
nand I_43641 (I744437,I744398,I744307);
nand I_43642 (I744015,I744290,I744437);
not I_43643 (I744468,I744398);
nor I_43644 (I744485,I744468,I744208);
DFFARX1 I_43645 (I744485,I2507,I744038,I744027,);
nor I_43646 (I744516,I58037,I58022);
or I_43647 (I744018,I744265,I744516);
nor I_43648 (I744009,I744398,I744516);
or I_43649 (I744012,I744132,I744516);
DFFARX1 I_43650 (I744516,I2507,I744038,I744030,);
not I_43651 (I744616,I2514);
DFFARX1 I_43652 (I1351749,I2507,I744616,I744642,);
not I_43653 (I744650,I744642);
nand I_43654 (I744667,I1351734,I1351722);
and I_43655 (I744684,I744667,I1351737);
DFFARX1 I_43656 (I744684,I2507,I744616,I744710,);
not I_43657 (I744718,I1351722);
DFFARX1 I_43658 (I1351740,I2507,I744616,I744744,);
not I_43659 (I744752,I744744);
nor I_43660 (I744769,I744752,I744650);
and I_43661 (I744786,I744769,I1351722);
nor I_43662 (I744803,I744752,I744718);
nor I_43663 (I744599,I744710,I744803);
DFFARX1 I_43664 (I1351728,I2507,I744616,I744843,);
nor I_43665 (I744851,I744843,I744710);
not I_43666 (I744868,I744851);
not I_43667 (I744885,I744843);
nor I_43668 (I744902,I744885,I744786);
DFFARX1 I_43669 (I744902,I2507,I744616,I744602,);
nand I_43670 (I744933,I1351725,I1351731);
and I_43671 (I744950,I744933,I1351746);
DFFARX1 I_43672 (I744950,I2507,I744616,I744976,);
nor I_43673 (I744984,I744976,I744843);
DFFARX1 I_43674 (I744984,I2507,I744616,I744584,);
nand I_43675 (I745015,I744976,I744885);
nand I_43676 (I744593,I744868,I745015);
not I_43677 (I745046,I744976);
nor I_43678 (I745063,I745046,I744786);
DFFARX1 I_43679 (I745063,I2507,I744616,I744605,);
nor I_43680 (I745094,I1351743,I1351731);
or I_43681 (I744596,I744843,I745094);
nor I_43682 (I744587,I744976,I745094);
or I_43683 (I744590,I744710,I745094);
DFFARX1 I_43684 (I745094,I2507,I744616,I744608,);
not I_43685 (I745194,I2514);
DFFARX1 I_43686 (I256538,I2507,I745194,I745220,);
not I_43687 (I745228,I745220);
nand I_43688 (I745245,I256541,I256517);
and I_43689 (I745262,I745245,I256514);
DFFARX1 I_43690 (I745262,I2507,I745194,I745288,);
not I_43691 (I745296,I256520);
DFFARX1 I_43692 (I256514,I2507,I745194,I745322,);
not I_43693 (I745330,I745322);
nor I_43694 (I745347,I745330,I745228);
and I_43695 (I745364,I745347,I256520);
nor I_43696 (I745381,I745330,I745296);
nor I_43697 (I745177,I745288,I745381);
DFFARX1 I_43698 (I256523,I2507,I745194,I745421,);
nor I_43699 (I745429,I745421,I745288);
not I_43700 (I745446,I745429);
not I_43701 (I745463,I745421);
nor I_43702 (I745480,I745463,I745364);
DFFARX1 I_43703 (I745480,I2507,I745194,I745180,);
nand I_43704 (I745511,I256526,I256535);
and I_43705 (I745528,I745511,I256532);
DFFARX1 I_43706 (I745528,I2507,I745194,I745554,);
nor I_43707 (I745562,I745554,I745421);
DFFARX1 I_43708 (I745562,I2507,I745194,I745162,);
nand I_43709 (I745593,I745554,I745463);
nand I_43710 (I745171,I745446,I745593);
not I_43711 (I745624,I745554);
nor I_43712 (I745641,I745624,I745364);
DFFARX1 I_43713 (I745641,I2507,I745194,I745183,);
nor I_43714 (I745672,I256529,I256535);
or I_43715 (I745174,I745421,I745672);
nor I_43716 (I745165,I745554,I745672);
or I_43717 (I745168,I745288,I745672);
DFFARX1 I_43718 (I745672,I2507,I745194,I745186,);
not I_43719 (I745772,I2514);
DFFARX1 I_43720 (I601818,I2507,I745772,I745798,);
not I_43721 (I745806,I745798);
nand I_43722 (I745823,I601827,I601836);
and I_43723 (I745840,I745823,I601842);
DFFARX1 I_43724 (I745840,I2507,I745772,I745866,);
not I_43725 (I745874,I601839);
DFFARX1 I_43726 (I601824,I2507,I745772,I745900,);
not I_43727 (I745908,I745900);
nor I_43728 (I745925,I745908,I745806);
and I_43729 (I745942,I745925,I601839);
nor I_43730 (I745959,I745908,I745874);
nor I_43731 (I745755,I745866,I745959);
DFFARX1 I_43732 (I601833,I2507,I745772,I745999,);
nor I_43733 (I746007,I745999,I745866);
not I_43734 (I746024,I746007);
not I_43735 (I746041,I745999);
nor I_43736 (I746058,I746041,I745942);
DFFARX1 I_43737 (I746058,I2507,I745772,I745758,);
nand I_43738 (I746089,I601830,I601821);
and I_43739 (I746106,I746089,I601818);
DFFARX1 I_43740 (I746106,I2507,I745772,I746132,);
nor I_43741 (I746140,I746132,I745999);
DFFARX1 I_43742 (I746140,I2507,I745772,I745740,);
nand I_43743 (I746171,I746132,I746041);
nand I_43744 (I745749,I746024,I746171);
not I_43745 (I746202,I746132);
nor I_43746 (I746219,I746202,I745942);
DFFARX1 I_43747 (I746219,I2507,I745772,I745761,);
nor I_43748 (I746250,I601821,I601821);
or I_43749 (I745752,I745999,I746250);
nor I_43750 (I745743,I746132,I746250);
or I_43751 (I745746,I745866,I746250);
DFFARX1 I_43752 (I746250,I2507,I745772,I745764,);
not I_43753 (I746350,I2514);
DFFARX1 I_43754 (I1189594,I2507,I746350,I746376,);
not I_43755 (I746384,I746376);
nand I_43756 (I746401,I1189576,I1189588);
and I_43757 (I746418,I746401,I1189591);
DFFARX1 I_43758 (I746418,I2507,I746350,I746444,);
not I_43759 (I746452,I1189585);
DFFARX1 I_43760 (I1189582,I2507,I746350,I746478,);
not I_43761 (I746486,I746478);
nor I_43762 (I746503,I746486,I746384);
and I_43763 (I746520,I746503,I1189585);
nor I_43764 (I746537,I746486,I746452);
nor I_43765 (I746333,I746444,I746537);
DFFARX1 I_43766 (I1189600,I2507,I746350,I746577,);
nor I_43767 (I746585,I746577,I746444);
not I_43768 (I746602,I746585);
not I_43769 (I746619,I746577);
nor I_43770 (I746636,I746619,I746520);
DFFARX1 I_43771 (I746636,I2507,I746350,I746336,);
nand I_43772 (I746667,I1189579,I1189579);
and I_43773 (I746684,I746667,I1189576);
DFFARX1 I_43774 (I746684,I2507,I746350,I746710,);
nor I_43775 (I746718,I746710,I746577);
DFFARX1 I_43776 (I746718,I2507,I746350,I746318,);
nand I_43777 (I746749,I746710,I746619);
nand I_43778 (I746327,I746602,I746749);
not I_43779 (I746780,I746710);
nor I_43780 (I746797,I746780,I746520);
DFFARX1 I_43781 (I746797,I2507,I746350,I746339,);
nor I_43782 (I746828,I1189597,I1189579);
or I_43783 (I746330,I746577,I746828);
nor I_43784 (I746321,I746710,I746828);
or I_43785 (I746324,I746444,I746828);
DFFARX1 I_43786 (I746828,I2507,I746350,I746342,);
not I_43787 (I746928,I2514);
DFFARX1 I_43788 (I1069370,I2507,I746928,I746954,);
not I_43789 (I746962,I746954);
nand I_43790 (I746979,I1069352,I1069364);
and I_43791 (I746996,I746979,I1069367);
DFFARX1 I_43792 (I746996,I2507,I746928,I747022,);
not I_43793 (I747030,I1069361);
DFFARX1 I_43794 (I1069358,I2507,I746928,I747056,);
not I_43795 (I747064,I747056);
nor I_43796 (I747081,I747064,I746962);
and I_43797 (I747098,I747081,I1069361);
nor I_43798 (I747115,I747064,I747030);
nor I_43799 (I746911,I747022,I747115);
DFFARX1 I_43800 (I1069376,I2507,I746928,I747155,);
nor I_43801 (I747163,I747155,I747022);
not I_43802 (I747180,I747163);
not I_43803 (I747197,I747155);
nor I_43804 (I747214,I747197,I747098);
DFFARX1 I_43805 (I747214,I2507,I746928,I746914,);
nand I_43806 (I747245,I1069355,I1069355);
and I_43807 (I747262,I747245,I1069352);
DFFARX1 I_43808 (I747262,I2507,I746928,I747288,);
nor I_43809 (I747296,I747288,I747155);
DFFARX1 I_43810 (I747296,I2507,I746928,I746896,);
nand I_43811 (I747327,I747288,I747197);
nand I_43812 (I746905,I747180,I747327);
not I_43813 (I747358,I747288);
nor I_43814 (I747375,I747358,I747098);
DFFARX1 I_43815 (I747375,I2507,I746928,I746917,);
nor I_43816 (I747406,I1069373,I1069355);
or I_43817 (I746908,I747155,I747406);
nor I_43818 (I746899,I747288,I747406);
or I_43819 (I746902,I747022,I747406);
DFFARX1 I_43820 (I747406,I2507,I746928,I746920,);
not I_43821 (I747506,I2514);
DFFARX1 I_43822 (I795939,I2507,I747506,I747532,);
not I_43823 (I747540,I747532);
nand I_43824 (I747557,I795927,I795945);
and I_43825 (I747574,I747557,I795942);
DFFARX1 I_43826 (I747574,I2507,I747506,I747600,);
not I_43827 (I747608,I795933);
DFFARX1 I_43828 (I795930,I2507,I747506,I747634,);
not I_43829 (I747642,I747634);
nor I_43830 (I747659,I747642,I747540);
and I_43831 (I747676,I747659,I795933);
nor I_43832 (I747693,I747642,I747608);
nor I_43833 (I747489,I747600,I747693);
DFFARX1 I_43834 (I795924,I2507,I747506,I747733,);
nor I_43835 (I747741,I747733,I747600);
not I_43836 (I747758,I747741);
not I_43837 (I747775,I747733);
nor I_43838 (I747792,I747775,I747676);
DFFARX1 I_43839 (I747792,I2507,I747506,I747492,);
nand I_43840 (I747823,I795924,I795927);
and I_43841 (I747840,I747823,I795930);
DFFARX1 I_43842 (I747840,I2507,I747506,I747866,);
nor I_43843 (I747874,I747866,I747733);
DFFARX1 I_43844 (I747874,I2507,I747506,I747474,);
nand I_43845 (I747905,I747866,I747775);
nand I_43846 (I747483,I747758,I747905);
not I_43847 (I747936,I747866);
nor I_43848 (I747953,I747936,I747676);
DFFARX1 I_43849 (I747953,I2507,I747506,I747495,);
nor I_43850 (I747984,I795936,I795927);
or I_43851 (I747486,I747733,I747984);
nor I_43852 (I747477,I747866,I747984);
or I_43853 (I747480,I747600,I747984);
DFFARX1 I_43854 (I747984,I2507,I747506,I747498,);
not I_43855 (I748084,I2514);
DFFARX1 I_43856 (I1102894,I2507,I748084,I748110,);
not I_43857 (I748118,I748110);
nand I_43858 (I748135,I1102876,I1102888);
and I_43859 (I748152,I748135,I1102891);
DFFARX1 I_43860 (I748152,I2507,I748084,I748178,);
not I_43861 (I748186,I1102885);
DFFARX1 I_43862 (I1102882,I2507,I748084,I748212,);
not I_43863 (I748220,I748212);
nor I_43864 (I748237,I748220,I748118);
and I_43865 (I748254,I748237,I1102885);
nor I_43866 (I748271,I748220,I748186);
nor I_43867 (I748067,I748178,I748271);
DFFARX1 I_43868 (I1102900,I2507,I748084,I748311,);
nor I_43869 (I748319,I748311,I748178);
not I_43870 (I748336,I748319);
not I_43871 (I748353,I748311);
nor I_43872 (I748370,I748353,I748254);
DFFARX1 I_43873 (I748370,I2507,I748084,I748070,);
nand I_43874 (I748401,I1102879,I1102879);
and I_43875 (I748418,I748401,I1102876);
DFFARX1 I_43876 (I748418,I2507,I748084,I748444,);
nor I_43877 (I748452,I748444,I748311);
DFFARX1 I_43878 (I748452,I2507,I748084,I748052,);
nand I_43879 (I748483,I748444,I748353);
nand I_43880 (I748061,I748336,I748483);
not I_43881 (I748514,I748444);
nor I_43882 (I748531,I748514,I748254);
DFFARX1 I_43883 (I748531,I2507,I748084,I748073,);
nor I_43884 (I748562,I1102897,I1102879);
or I_43885 (I748064,I748311,I748562);
nor I_43886 (I748055,I748444,I748562);
or I_43887 (I748058,I748178,I748562);
DFFARX1 I_43888 (I748562,I2507,I748084,I748076,);
not I_43889 (I748662,I2514);
DFFARX1 I_43890 (I614534,I2507,I748662,I748688,);
not I_43891 (I748696,I748688);
nand I_43892 (I748713,I614543,I614552);
and I_43893 (I748730,I748713,I614558);
DFFARX1 I_43894 (I748730,I2507,I748662,I748756,);
not I_43895 (I748764,I614555);
DFFARX1 I_43896 (I614540,I2507,I748662,I748790,);
not I_43897 (I748798,I748790);
nor I_43898 (I748815,I748798,I748696);
and I_43899 (I748832,I748815,I614555);
nor I_43900 (I748849,I748798,I748764);
nor I_43901 (I748645,I748756,I748849);
DFFARX1 I_43902 (I614549,I2507,I748662,I748889,);
nor I_43903 (I748897,I748889,I748756);
not I_43904 (I748914,I748897);
not I_43905 (I748931,I748889);
nor I_43906 (I748948,I748931,I748832);
DFFARX1 I_43907 (I748948,I2507,I748662,I748648,);
nand I_43908 (I748979,I614546,I614537);
and I_43909 (I748996,I748979,I614534);
DFFARX1 I_43910 (I748996,I2507,I748662,I749022,);
nor I_43911 (I749030,I749022,I748889);
DFFARX1 I_43912 (I749030,I2507,I748662,I748630,);
nand I_43913 (I749061,I749022,I748931);
nand I_43914 (I748639,I748914,I749061);
not I_43915 (I749092,I749022);
nor I_43916 (I749109,I749092,I748832);
DFFARX1 I_43917 (I749109,I2507,I748662,I748651,);
nor I_43918 (I749140,I614537,I614537);
or I_43919 (I748642,I748889,I749140);
nor I_43920 (I748633,I749022,I749140);
or I_43921 (I748636,I748756,I749140);
DFFARX1 I_43922 (I749140,I2507,I748662,I748654,);
not I_43923 (I749240,I2514);
DFFARX1 I_43924 (I1110986,I2507,I749240,I749266,);
not I_43925 (I749274,I749266);
nand I_43926 (I749291,I1110968,I1110980);
and I_43927 (I749308,I749291,I1110983);
DFFARX1 I_43928 (I749308,I2507,I749240,I749334,);
not I_43929 (I749342,I1110977);
DFFARX1 I_43930 (I1110974,I2507,I749240,I749368,);
not I_43931 (I749376,I749368);
nor I_43932 (I749393,I749376,I749274);
and I_43933 (I749410,I749393,I1110977);
nor I_43934 (I749427,I749376,I749342);
nor I_43935 (I749223,I749334,I749427);
DFFARX1 I_43936 (I1110992,I2507,I749240,I749467,);
nor I_43937 (I749475,I749467,I749334);
not I_43938 (I749492,I749475);
not I_43939 (I749509,I749467);
nor I_43940 (I749526,I749509,I749410);
DFFARX1 I_43941 (I749526,I2507,I749240,I749226,);
nand I_43942 (I749557,I1110971,I1110971);
and I_43943 (I749574,I749557,I1110968);
DFFARX1 I_43944 (I749574,I2507,I749240,I749600,);
nor I_43945 (I749608,I749600,I749467);
DFFARX1 I_43946 (I749608,I2507,I749240,I749208,);
nand I_43947 (I749639,I749600,I749509);
nand I_43948 (I749217,I749492,I749639);
not I_43949 (I749670,I749600);
nor I_43950 (I749687,I749670,I749410);
DFFARX1 I_43951 (I749687,I2507,I749240,I749229,);
nor I_43952 (I749718,I1110989,I1110971);
or I_43953 (I749220,I749467,I749718);
nor I_43954 (I749211,I749600,I749718);
or I_43955 (I749214,I749334,I749718);
DFFARX1 I_43956 (I749718,I2507,I749240,I749232,);
not I_43957 (I749818,I2514);
DFFARX1 I_43958 (I321886,I2507,I749818,I749844,);
not I_43959 (I749852,I749844);
nand I_43960 (I749869,I321889,I321865);
and I_43961 (I749886,I749869,I321862);
DFFARX1 I_43962 (I749886,I2507,I749818,I749912,);
not I_43963 (I749920,I321868);
DFFARX1 I_43964 (I321862,I2507,I749818,I749946,);
not I_43965 (I749954,I749946);
nor I_43966 (I749971,I749954,I749852);
and I_43967 (I749988,I749971,I321868);
nor I_43968 (I750005,I749954,I749920);
nor I_43969 (I749801,I749912,I750005);
DFFARX1 I_43970 (I321871,I2507,I749818,I750045,);
nor I_43971 (I750053,I750045,I749912);
not I_43972 (I750070,I750053);
not I_43973 (I750087,I750045);
nor I_43974 (I750104,I750087,I749988);
DFFARX1 I_43975 (I750104,I2507,I749818,I749804,);
nand I_43976 (I750135,I321874,I321883);
and I_43977 (I750152,I750135,I321880);
DFFARX1 I_43978 (I750152,I2507,I749818,I750178,);
nor I_43979 (I750186,I750178,I750045);
DFFARX1 I_43980 (I750186,I2507,I749818,I749786,);
nand I_43981 (I750217,I750178,I750087);
nand I_43982 (I749795,I750070,I750217);
not I_43983 (I750248,I750178);
nor I_43984 (I750265,I750248,I749988);
DFFARX1 I_43985 (I750265,I2507,I749818,I749807,);
nor I_43986 (I750296,I321877,I321883);
or I_43987 (I749798,I750045,I750296);
nor I_43988 (I749789,I750178,I750296);
or I_43989 (I749792,I749912,I750296);
DFFARX1 I_43990 (I750296,I2507,I749818,I749810,);
not I_43991 (I750396,I2514);
DFFARX1 I_43992 (I69619,I2507,I750396,I750422,);
not I_43993 (I750430,I750422);
nand I_43994 (I750447,I69628,I69637);
and I_43995 (I750464,I750447,I69616);
DFFARX1 I_43996 (I750464,I2507,I750396,I750490,);
not I_43997 (I750498,I69619);
DFFARX1 I_43998 (I69634,I2507,I750396,I750524,);
not I_43999 (I750532,I750524);
nor I_44000 (I750549,I750532,I750430);
and I_44001 (I750566,I750549,I69619);
nor I_44002 (I750583,I750532,I750498);
nor I_44003 (I750379,I750490,I750583);
DFFARX1 I_44004 (I69625,I2507,I750396,I750623,);
nor I_44005 (I750631,I750623,I750490);
not I_44006 (I750648,I750631);
not I_44007 (I750665,I750623);
nor I_44008 (I750682,I750665,I750566);
DFFARX1 I_44009 (I750682,I2507,I750396,I750382,);
nand I_44010 (I750713,I69640,I69616);
and I_44011 (I750730,I750713,I69622);
DFFARX1 I_44012 (I750730,I2507,I750396,I750756,);
nor I_44013 (I750764,I750756,I750623);
DFFARX1 I_44014 (I750764,I2507,I750396,I750364,);
nand I_44015 (I750795,I750756,I750665);
nand I_44016 (I750373,I750648,I750795);
not I_44017 (I750826,I750756);
nor I_44018 (I750843,I750826,I750566);
DFFARX1 I_44019 (I750843,I2507,I750396,I750385,);
nor I_44020 (I750874,I69631,I69616);
or I_44021 (I750376,I750623,I750874);
nor I_44022 (I750367,I750756,I750874);
or I_44023 (I750370,I750490,I750874);
DFFARX1 I_44024 (I750874,I2507,I750396,I750388,);
not I_44025 (I750974,I2514);
DFFARX1 I_44026 (I259173,I2507,I750974,I751000,);
not I_44027 (I751008,I751000);
nand I_44028 (I751025,I259176,I259152);
and I_44029 (I751042,I751025,I259149);
DFFARX1 I_44030 (I751042,I2507,I750974,I751068,);
not I_44031 (I751076,I259155);
DFFARX1 I_44032 (I259149,I2507,I750974,I751102,);
not I_44033 (I751110,I751102);
nor I_44034 (I751127,I751110,I751008);
and I_44035 (I751144,I751127,I259155);
nor I_44036 (I751161,I751110,I751076);
nor I_44037 (I750957,I751068,I751161);
DFFARX1 I_44038 (I259158,I2507,I750974,I751201,);
nor I_44039 (I751209,I751201,I751068);
not I_44040 (I751226,I751209);
not I_44041 (I751243,I751201);
nor I_44042 (I751260,I751243,I751144);
DFFARX1 I_44043 (I751260,I2507,I750974,I750960,);
nand I_44044 (I751291,I259161,I259170);
and I_44045 (I751308,I751291,I259167);
DFFARX1 I_44046 (I751308,I2507,I750974,I751334,);
nor I_44047 (I751342,I751334,I751201);
DFFARX1 I_44048 (I751342,I2507,I750974,I750942,);
nand I_44049 (I751373,I751334,I751243);
nand I_44050 (I750951,I751226,I751373);
not I_44051 (I751404,I751334);
nor I_44052 (I751421,I751404,I751144);
DFFARX1 I_44053 (I751421,I2507,I750974,I750963,);
nor I_44054 (I751452,I259164,I259170);
or I_44055 (I750954,I751201,I751452);
nor I_44056 (I750945,I751334,I751452);
or I_44057 (I750948,I751068,I751452);
DFFARX1 I_44058 (I751452,I2507,I750974,I750966,);
not I_44059 (I751552,I2514);
DFFARX1 I_44060 (I258646,I2507,I751552,I751578,);
not I_44061 (I751586,I751578);
nand I_44062 (I751603,I258649,I258625);
and I_44063 (I751620,I751603,I258622);
DFFARX1 I_44064 (I751620,I2507,I751552,I751646,);
not I_44065 (I751654,I258628);
DFFARX1 I_44066 (I258622,I2507,I751552,I751680,);
not I_44067 (I751688,I751680);
nor I_44068 (I751705,I751688,I751586);
and I_44069 (I751722,I751705,I258628);
nor I_44070 (I751739,I751688,I751654);
nor I_44071 (I751535,I751646,I751739);
DFFARX1 I_44072 (I258631,I2507,I751552,I751779,);
nor I_44073 (I751787,I751779,I751646);
not I_44074 (I751804,I751787);
not I_44075 (I751821,I751779);
nor I_44076 (I751838,I751821,I751722);
DFFARX1 I_44077 (I751838,I2507,I751552,I751538,);
nand I_44078 (I751869,I258634,I258643);
and I_44079 (I751886,I751869,I258640);
DFFARX1 I_44080 (I751886,I2507,I751552,I751912,);
nor I_44081 (I751920,I751912,I751779);
DFFARX1 I_44082 (I751920,I2507,I751552,I751520,);
nand I_44083 (I751951,I751912,I751821);
nand I_44084 (I751529,I751804,I751951);
not I_44085 (I751982,I751912);
nor I_44086 (I751999,I751982,I751722);
DFFARX1 I_44087 (I751999,I2507,I751552,I751541,);
nor I_44088 (I752030,I258637,I258643);
or I_44089 (I751532,I751779,I752030);
nor I_44090 (I751523,I751912,I752030);
or I_44091 (I751526,I751646,I752030);
DFFARX1 I_44092 (I752030,I2507,I751552,I751544,);
not I_44093 (I752130,I2514);
DFFARX1 I_44094 (I118103,I2507,I752130,I752156,);
not I_44095 (I752164,I752156);
nand I_44096 (I752181,I118112,I118121);
and I_44097 (I752198,I752181,I118100);
DFFARX1 I_44098 (I752198,I2507,I752130,I752224,);
not I_44099 (I752232,I118103);
DFFARX1 I_44100 (I118118,I2507,I752130,I752258,);
not I_44101 (I752266,I752258);
nor I_44102 (I752283,I752266,I752164);
and I_44103 (I752300,I752283,I118103);
nor I_44104 (I752317,I752266,I752232);
nor I_44105 (I752113,I752224,I752317);
DFFARX1 I_44106 (I118109,I2507,I752130,I752357,);
nor I_44107 (I752365,I752357,I752224);
not I_44108 (I752382,I752365);
not I_44109 (I752399,I752357);
nor I_44110 (I752416,I752399,I752300);
DFFARX1 I_44111 (I752416,I2507,I752130,I752116,);
nand I_44112 (I752447,I118124,I118100);
and I_44113 (I752464,I752447,I118106);
DFFARX1 I_44114 (I752464,I2507,I752130,I752490,);
nor I_44115 (I752498,I752490,I752357);
DFFARX1 I_44116 (I752498,I2507,I752130,I752098,);
nand I_44117 (I752529,I752490,I752399);
nand I_44118 (I752107,I752382,I752529);
not I_44119 (I752560,I752490);
nor I_44120 (I752577,I752560,I752300);
DFFARX1 I_44121 (I752577,I2507,I752130,I752119,);
nor I_44122 (I752608,I118115,I118100);
or I_44123 (I752110,I752357,I752608);
nor I_44124 (I752101,I752490,I752608);
or I_44125 (I752104,I752224,I752608);
DFFARX1 I_44126 (I752608,I2507,I752130,I752122,);
not I_44127 (I752708,I2514);
DFFARX1 I_44128 (I200805,I2507,I752708,I752734,);
not I_44129 (I752742,I752734);
nand I_44130 (I752759,I200808,I200829);
and I_44131 (I752776,I752759,I200817);
DFFARX1 I_44132 (I752776,I2507,I752708,I752802,);
not I_44133 (I752810,I200814);
DFFARX1 I_44134 (I200805,I2507,I752708,I752836,);
not I_44135 (I752844,I752836);
nor I_44136 (I752861,I752844,I752742);
and I_44137 (I752878,I752861,I200814);
nor I_44138 (I752895,I752844,I752810);
nor I_44139 (I752691,I752802,I752895);
DFFARX1 I_44140 (I200823,I2507,I752708,I752935,);
nor I_44141 (I752943,I752935,I752802);
not I_44142 (I752960,I752943);
not I_44143 (I752977,I752935);
nor I_44144 (I752994,I752977,I752878);
DFFARX1 I_44145 (I752994,I2507,I752708,I752694,);
nand I_44146 (I753025,I200808,I200811);
and I_44147 (I753042,I753025,I200820);
DFFARX1 I_44148 (I753042,I2507,I752708,I753068,);
nor I_44149 (I753076,I753068,I752935);
DFFARX1 I_44150 (I753076,I2507,I752708,I752676,);
nand I_44151 (I753107,I753068,I752977);
nand I_44152 (I752685,I752960,I753107);
not I_44153 (I753138,I753068);
nor I_44154 (I753155,I753138,I752878);
DFFARX1 I_44155 (I753155,I2507,I752708,I752697,);
nor I_44156 (I753186,I200826,I200811);
or I_44157 (I752688,I752935,I753186);
nor I_44158 (I752679,I753068,I753186);
or I_44159 (I752682,I752802,I753186);
DFFARX1 I_44160 (I753186,I2507,I752708,I752700,);
not I_44161 (I753286,I2514);
DFFARX1 I_44162 (I1193062,I2507,I753286,I753312,);
not I_44163 (I753320,I753312);
nand I_44164 (I753337,I1193044,I1193056);
and I_44165 (I753354,I753337,I1193059);
DFFARX1 I_44166 (I753354,I2507,I753286,I753380,);
not I_44167 (I753388,I1193053);
DFFARX1 I_44168 (I1193050,I2507,I753286,I753414,);
not I_44169 (I753422,I753414);
nor I_44170 (I753439,I753422,I753320);
and I_44171 (I753456,I753439,I1193053);
nor I_44172 (I753473,I753422,I753388);
nor I_44173 (I753269,I753380,I753473);
DFFARX1 I_44174 (I1193068,I2507,I753286,I753513,);
nor I_44175 (I753521,I753513,I753380);
not I_44176 (I753538,I753521);
not I_44177 (I753555,I753513);
nor I_44178 (I753572,I753555,I753456);
DFFARX1 I_44179 (I753572,I2507,I753286,I753272,);
nand I_44180 (I753603,I1193047,I1193047);
and I_44181 (I753620,I753603,I1193044);
DFFARX1 I_44182 (I753620,I2507,I753286,I753646,);
nor I_44183 (I753654,I753646,I753513);
DFFARX1 I_44184 (I753654,I2507,I753286,I753254,);
nand I_44185 (I753685,I753646,I753555);
nand I_44186 (I753263,I753538,I753685);
not I_44187 (I753716,I753646);
nor I_44188 (I753733,I753716,I753456);
DFFARX1 I_44189 (I753733,I2507,I753286,I753275,);
nor I_44190 (I753764,I1193065,I1193047);
or I_44191 (I753266,I753513,I753764);
nor I_44192 (I753257,I753646,I753764);
or I_44193 (I753260,I753380,I753764);
DFFARX1 I_44194 (I753764,I2507,I753286,I753278,);
not I_44195 (I753864,I2514);
DFFARX1 I_44196 (I623204,I2507,I753864,I753890,);
not I_44197 (I753898,I753890);
nand I_44198 (I753915,I623213,I623222);
and I_44199 (I753932,I753915,I623228);
DFFARX1 I_44200 (I753932,I2507,I753864,I753958,);
not I_44201 (I753966,I623225);
DFFARX1 I_44202 (I623210,I2507,I753864,I753992,);
not I_44203 (I754000,I753992);
nor I_44204 (I754017,I754000,I753898);
and I_44205 (I754034,I754017,I623225);
nor I_44206 (I754051,I754000,I753966);
nor I_44207 (I753847,I753958,I754051);
DFFARX1 I_44208 (I623219,I2507,I753864,I754091,);
nor I_44209 (I754099,I754091,I753958);
not I_44210 (I754116,I754099);
not I_44211 (I754133,I754091);
nor I_44212 (I754150,I754133,I754034);
DFFARX1 I_44213 (I754150,I2507,I753864,I753850,);
nand I_44214 (I754181,I623216,I623207);
and I_44215 (I754198,I754181,I623204);
DFFARX1 I_44216 (I754198,I2507,I753864,I754224,);
nor I_44217 (I754232,I754224,I754091);
DFFARX1 I_44218 (I754232,I2507,I753864,I753832,);
nand I_44219 (I754263,I754224,I754133);
nand I_44220 (I753841,I754116,I754263);
not I_44221 (I754294,I754224);
nor I_44222 (I754311,I754294,I754034);
DFFARX1 I_44223 (I754311,I2507,I753864,I753853,);
nor I_44224 (I754342,I623207,I623207);
or I_44225 (I753844,I754091,I754342);
nor I_44226 (I753835,I754224,I754342);
or I_44227 (I753838,I753958,I754342);
DFFARX1 I_44228 (I754342,I2507,I753864,I753856,);
not I_44229 (I754442,I2514);
DFFARX1 I_44230 (I410424,I2507,I754442,I754468,);
not I_44231 (I754476,I754468);
nand I_44232 (I754493,I410415,I410433);
and I_44233 (I754510,I754493,I410436);
DFFARX1 I_44234 (I754510,I2507,I754442,I754536,);
not I_44235 (I754544,I410430);
DFFARX1 I_44236 (I410418,I2507,I754442,I754570,);
not I_44237 (I754578,I754570);
nor I_44238 (I754595,I754578,I754476);
and I_44239 (I754612,I754595,I410430);
nor I_44240 (I754629,I754578,I754544);
nor I_44241 (I754425,I754536,I754629);
DFFARX1 I_44242 (I410427,I2507,I754442,I754669,);
nor I_44243 (I754677,I754669,I754536);
not I_44244 (I754694,I754677);
not I_44245 (I754711,I754669);
nor I_44246 (I754728,I754711,I754612);
DFFARX1 I_44247 (I754728,I2507,I754442,I754428,);
nand I_44248 (I754759,I410442,I410439);
and I_44249 (I754776,I754759,I410421);
DFFARX1 I_44250 (I754776,I2507,I754442,I754802,);
nor I_44251 (I754810,I754802,I754669);
DFFARX1 I_44252 (I754810,I2507,I754442,I754410,);
nand I_44253 (I754841,I754802,I754711);
nand I_44254 (I754419,I754694,I754841);
not I_44255 (I754872,I754802);
nor I_44256 (I754889,I754872,I754612);
DFFARX1 I_44257 (I754889,I2507,I754442,I754431,);
nor I_44258 (I754920,I410415,I410439);
or I_44259 (I754422,I754669,I754920);
nor I_44260 (I754413,I754802,I754920);
or I_44261 (I754416,I754536,I754920);
DFFARX1 I_44262 (I754920,I2507,I754442,I754434,);
not I_44263 (I755020,I2514);
DFFARX1 I_44264 (I1090178,I2507,I755020,I755046,);
not I_44265 (I755054,I755046);
nand I_44266 (I755071,I1090160,I1090172);
and I_44267 (I755088,I755071,I1090175);
DFFARX1 I_44268 (I755088,I2507,I755020,I755114,);
not I_44269 (I755122,I1090169);
DFFARX1 I_44270 (I1090166,I2507,I755020,I755148,);
not I_44271 (I755156,I755148);
nor I_44272 (I755173,I755156,I755054);
and I_44273 (I755190,I755173,I1090169);
nor I_44274 (I755207,I755156,I755122);
nor I_44275 (I755003,I755114,I755207);
DFFARX1 I_44276 (I1090184,I2507,I755020,I755247,);
nor I_44277 (I755255,I755247,I755114);
not I_44278 (I755272,I755255);
not I_44279 (I755289,I755247);
nor I_44280 (I755306,I755289,I755190);
DFFARX1 I_44281 (I755306,I2507,I755020,I755006,);
nand I_44282 (I755337,I1090163,I1090163);
and I_44283 (I755354,I755337,I1090160);
DFFARX1 I_44284 (I755354,I2507,I755020,I755380,);
nor I_44285 (I755388,I755380,I755247);
DFFARX1 I_44286 (I755388,I2507,I755020,I754988,);
nand I_44287 (I755419,I755380,I755289);
nand I_44288 (I754997,I755272,I755419);
not I_44289 (I755450,I755380);
nor I_44290 (I755467,I755450,I755190);
DFFARX1 I_44291 (I755467,I2507,I755020,I755009,);
nor I_44292 (I755498,I1090181,I1090163);
or I_44293 (I755000,I755247,I755498);
nor I_44294 (I754991,I755380,I755498);
or I_44295 (I754994,I755114,I755498);
DFFARX1 I_44296 (I755498,I2507,I755020,I755012,);
not I_44297 (I755598,I2514);
DFFARX1 I_44298 (I23779,I2507,I755598,I755624,);
not I_44299 (I755632,I755624);
nand I_44300 (I755649,I23776,I23767);
and I_44301 (I755666,I755649,I23767);
DFFARX1 I_44302 (I755666,I2507,I755598,I755692,);
not I_44303 (I755700,I23770);
DFFARX1 I_44304 (I23785,I2507,I755598,I755726,);
not I_44305 (I755734,I755726);
nor I_44306 (I755751,I755734,I755632);
and I_44307 (I755768,I755751,I23770);
nor I_44308 (I755785,I755734,I755700);
nor I_44309 (I755581,I755692,I755785);
DFFARX1 I_44310 (I23770,I2507,I755598,I755825,);
nor I_44311 (I755833,I755825,I755692);
not I_44312 (I755850,I755833);
not I_44313 (I755867,I755825);
nor I_44314 (I755884,I755867,I755768);
DFFARX1 I_44315 (I755884,I2507,I755598,I755584,);
nand I_44316 (I755915,I23788,I23773);
and I_44317 (I755932,I755915,I23791);
DFFARX1 I_44318 (I755932,I2507,I755598,I755958,);
nor I_44319 (I755966,I755958,I755825);
DFFARX1 I_44320 (I755966,I2507,I755598,I755566,);
nand I_44321 (I755997,I755958,I755867);
nand I_44322 (I755575,I755850,I755997);
not I_44323 (I756028,I755958);
nor I_44324 (I756045,I756028,I755768);
DFFARX1 I_44325 (I756045,I2507,I755598,I755587,);
nor I_44326 (I756076,I23782,I23773);
or I_44327 (I755578,I755825,I756076);
nor I_44328 (I755569,I755958,I756076);
or I_44329 (I755572,I755692,I756076);
DFFARX1 I_44330 (I756076,I2507,I755598,I755590,);
not I_44331 (I756176,I2514);
DFFARX1 I_44332 (I1388639,I2507,I756176,I756202,);
not I_44333 (I756210,I756202);
nand I_44334 (I756227,I1388624,I1388612);
and I_44335 (I756244,I756227,I1388627);
DFFARX1 I_44336 (I756244,I2507,I756176,I756270,);
not I_44337 (I756278,I1388612);
DFFARX1 I_44338 (I1388630,I2507,I756176,I756304,);
not I_44339 (I756312,I756304);
nor I_44340 (I756329,I756312,I756210);
and I_44341 (I756346,I756329,I1388612);
nor I_44342 (I756363,I756312,I756278);
nor I_44343 (I756159,I756270,I756363);
DFFARX1 I_44344 (I1388618,I2507,I756176,I756403,);
nor I_44345 (I756411,I756403,I756270);
not I_44346 (I756428,I756411);
not I_44347 (I756445,I756403);
nor I_44348 (I756462,I756445,I756346);
DFFARX1 I_44349 (I756462,I2507,I756176,I756162,);
nand I_44350 (I756493,I1388615,I1388621);
and I_44351 (I756510,I756493,I1388636);
DFFARX1 I_44352 (I756510,I2507,I756176,I756536,);
nor I_44353 (I756544,I756536,I756403);
DFFARX1 I_44354 (I756544,I2507,I756176,I756144,);
nand I_44355 (I756575,I756536,I756445);
nand I_44356 (I756153,I756428,I756575);
not I_44357 (I756606,I756536);
nor I_44358 (I756623,I756606,I756346);
DFFARX1 I_44359 (I756623,I2507,I756176,I756165,);
nor I_44360 (I756654,I1388633,I1388621);
or I_44361 (I756156,I756403,I756654);
nor I_44362 (I756147,I756536,I756654);
or I_44363 (I756150,I756270,I756654);
DFFARX1 I_44364 (I756654,I2507,I756176,I756168,);
not I_44365 (I756754,I2514);
DFFARX1 I_44366 (I1065902,I2507,I756754,I756780,);
not I_44367 (I756788,I756780);
nand I_44368 (I756805,I1065884,I1065896);
and I_44369 (I756822,I756805,I1065899);
DFFARX1 I_44370 (I756822,I2507,I756754,I756848,);
not I_44371 (I756856,I1065893);
DFFARX1 I_44372 (I1065890,I2507,I756754,I756882,);
not I_44373 (I756890,I756882);
nor I_44374 (I756907,I756890,I756788);
and I_44375 (I756924,I756907,I1065893);
nor I_44376 (I756941,I756890,I756856);
nor I_44377 (I756737,I756848,I756941);
DFFARX1 I_44378 (I1065908,I2507,I756754,I756981,);
nor I_44379 (I756989,I756981,I756848);
not I_44380 (I757006,I756989);
not I_44381 (I757023,I756981);
nor I_44382 (I757040,I757023,I756924);
DFFARX1 I_44383 (I757040,I2507,I756754,I756740,);
nand I_44384 (I757071,I1065887,I1065887);
and I_44385 (I757088,I757071,I1065884);
DFFARX1 I_44386 (I757088,I2507,I756754,I757114,);
nor I_44387 (I757122,I757114,I756981);
DFFARX1 I_44388 (I757122,I2507,I756754,I756722,);
nand I_44389 (I757153,I757114,I757023);
nand I_44390 (I756731,I757006,I757153);
not I_44391 (I757184,I757114);
nor I_44392 (I757201,I757184,I756924);
DFFARX1 I_44393 (I757201,I2507,I756754,I756743,);
nor I_44394 (I757232,I1065905,I1065887);
or I_44395 (I756734,I756981,I757232);
nor I_44396 (I756725,I757114,I757232);
or I_44397 (I756728,I756848,I757232);
DFFARX1 I_44398 (I757232,I2507,I756754,I756746,);
not I_44399 (I757332,I2514);
DFFARX1 I_44400 (I561358,I2507,I757332,I757358,);
not I_44401 (I757366,I757358);
nand I_44402 (I757383,I561367,I561376);
and I_44403 (I757400,I757383,I561382);
DFFARX1 I_44404 (I757400,I2507,I757332,I757426,);
not I_44405 (I757434,I561379);
DFFARX1 I_44406 (I561364,I2507,I757332,I757460,);
not I_44407 (I757468,I757460);
nor I_44408 (I757485,I757468,I757366);
and I_44409 (I757502,I757485,I561379);
nor I_44410 (I757519,I757468,I757434);
nor I_44411 (I757315,I757426,I757519);
DFFARX1 I_44412 (I561373,I2507,I757332,I757559,);
nor I_44413 (I757567,I757559,I757426);
not I_44414 (I757584,I757567);
not I_44415 (I757601,I757559);
nor I_44416 (I757618,I757601,I757502);
DFFARX1 I_44417 (I757618,I2507,I757332,I757318,);
nand I_44418 (I757649,I561370,I561361);
and I_44419 (I757666,I757649,I561358);
DFFARX1 I_44420 (I757666,I2507,I757332,I757692,);
nor I_44421 (I757700,I757692,I757559);
DFFARX1 I_44422 (I757700,I2507,I757332,I757300,);
nand I_44423 (I757731,I757692,I757601);
nand I_44424 (I757309,I757584,I757731);
not I_44425 (I757762,I757692);
nor I_44426 (I757779,I757762,I757502);
DFFARX1 I_44427 (I757779,I2507,I757332,I757321,);
nor I_44428 (I757810,I561361,I561361);
or I_44429 (I757312,I757559,I757810);
nor I_44430 (I757303,I757692,I757810);
or I_44431 (I757306,I757426,I757810);
DFFARX1 I_44432 (I757810,I2507,I757332,I757324,);
not I_44433 (I757910,I2514);
DFFARX1 I_44434 (I402264,I2507,I757910,I757936,);
not I_44435 (I757944,I757936);
nand I_44436 (I757961,I402255,I402273);
and I_44437 (I757978,I757961,I402276);
DFFARX1 I_44438 (I757978,I2507,I757910,I758004,);
not I_44439 (I758012,I402270);
DFFARX1 I_44440 (I402258,I2507,I757910,I758038,);
not I_44441 (I758046,I758038);
nor I_44442 (I758063,I758046,I757944);
and I_44443 (I758080,I758063,I402270);
nor I_44444 (I758097,I758046,I758012);
nor I_44445 (I757893,I758004,I758097);
DFFARX1 I_44446 (I402267,I2507,I757910,I758137,);
nor I_44447 (I758145,I758137,I758004);
not I_44448 (I758162,I758145);
not I_44449 (I758179,I758137);
nor I_44450 (I758196,I758179,I758080);
DFFARX1 I_44451 (I758196,I2507,I757910,I757896,);
nand I_44452 (I758227,I402282,I402279);
and I_44453 (I758244,I758227,I402261);
DFFARX1 I_44454 (I758244,I2507,I757910,I758270,);
nor I_44455 (I758278,I758270,I758137);
DFFARX1 I_44456 (I758278,I2507,I757910,I757878,);
nand I_44457 (I758309,I758270,I758179);
nand I_44458 (I757887,I758162,I758309);
not I_44459 (I758340,I758270);
nor I_44460 (I758357,I758340,I758080);
DFFARX1 I_44461 (I758357,I2507,I757910,I757899,);
nor I_44462 (I758388,I402255,I402279);
or I_44463 (I757890,I758137,I758388);
nor I_44464 (I757881,I758270,I758388);
or I_44465 (I757884,I758004,I758388);
DFFARX1 I_44466 (I758388,I2507,I757910,I757902,);
not I_44467 (I758488,I2514);
DFFARX1 I_44468 (I1335684,I2507,I758488,I758514,);
not I_44469 (I758522,I758514);
nand I_44470 (I758539,I1335669,I1335657);
and I_44471 (I758556,I758539,I1335672);
DFFARX1 I_44472 (I758556,I2507,I758488,I758582,);
not I_44473 (I758590,I1335657);
DFFARX1 I_44474 (I1335675,I2507,I758488,I758616,);
not I_44475 (I758624,I758616);
nor I_44476 (I758641,I758624,I758522);
and I_44477 (I758658,I758641,I1335657);
nor I_44478 (I758675,I758624,I758590);
nor I_44479 (I758471,I758582,I758675);
DFFARX1 I_44480 (I1335663,I2507,I758488,I758715,);
nor I_44481 (I758723,I758715,I758582);
not I_44482 (I758740,I758723);
not I_44483 (I758757,I758715);
nor I_44484 (I758774,I758757,I758658);
DFFARX1 I_44485 (I758774,I2507,I758488,I758474,);
nand I_44486 (I758805,I1335660,I1335666);
and I_44487 (I758822,I758805,I1335681);
DFFARX1 I_44488 (I758822,I2507,I758488,I758848,);
nor I_44489 (I758856,I758848,I758715);
DFFARX1 I_44490 (I758856,I2507,I758488,I758456,);
nand I_44491 (I758887,I758848,I758757);
nand I_44492 (I758465,I758740,I758887);
not I_44493 (I758918,I758848);
nor I_44494 (I758935,I758918,I758658);
DFFARX1 I_44495 (I758935,I2507,I758488,I758477,);
nor I_44496 (I758966,I1335678,I1335666);
or I_44497 (I758468,I758715,I758966);
nor I_44498 (I758459,I758848,I758966);
or I_44499 (I758462,I758582,I758966);
DFFARX1 I_44500 (I758966,I2507,I758488,I758480,);
not I_44501 (I759066,I2514);
DFFARX1 I_44502 (I1021367,I2507,I759066,I759092,);
not I_44503 (I759100,I759092);
nand I_44504 (I759117,I1021364,I1021382);
and I_44505 (I759134,I759117,I1021379);
DFFARX1 I_44506 (I759134,I2507,I759066,I759160,);
not I_44507 (I759168,I1021361);
DFFARX1 I_44508 (I1021364,I2507,I759066,I759194,);
not I_44509 (I759202,I759194);
nor I_44510 (I759219,I759202,I759100);
and I_44511 (I759236,I759219,I1021361);
nor I_44512 (I759253,I759202,I759168);
nor I_44513 (I759049,I759160,I759253);
DFFARX1 I_44514 (I1021373,I2507,I759066,I759293,);
nor I_44515 (I759301,I759293,I759160);
not I_44516 (I759318,I759301);
not I_44517 (I759335,I759293);
nor I_44518 (I759352,I759335,I759236);
DFFARX1 I_44519 (I759352,I2507,I759066,I759052,);
nand I_44520 (I759383,I1021376,I1021361);
and I_44521 (I759400,I759383,I1021367);
DFFARX1 I_44522 (I759400,I2507,I759066,I759426,);
nor I_44523 (I759434,I759426,I759293);
DFFARX1 I_44524 (I759434,I2507,I759066,I759034,);
nand I_44525 (I759465,I759426,I759335);
nand I_44526 (I759043,I759318,I759465);
not I_44527 (I759496,I759426);
nor I_44528 (I759513,I759496,I759236);
DFFARX1 I_44529 (I759513,I2507,I759066,I759055,);
nor I_44530 (I759544,I1021370,I1021361);
or I_44531 (I759046,I759293,I759544);
nor I_44532 (I759037,I759426,I759544);
or I_44533 (I759040,I759160,I759544);
DFFARX1 I_44534 (I759544,I2507,I759066,I759058,);
not I_44535 (I759644,I2514);
DFFARX1 I_44536 (I1271516,I2507,I759644,I759670,);
not I_44537 (I759678,I759670);
nand I_44538 (I759695,I1271540,I1271522);
and I_44539 (I759712,I759695,I1271528);
DFFARX1 I_44540 (I759712,I2507,I759644,I759738,);
not I_44541 (I759746,I1271534);
DFFARX1 I_44542 (I1271519,I2507,I759644,I759772,);
not I_44543 (I759780,I759772);
nor I_44544 (I759797,I759780,I759678);
and I_44545 (I759814,I759797,I1271534);
nor I_44546 (I759831,I759780,I759746);
nor I_44547 (I759627,I759738,I759831);
DFFARX1 I_44548 (I1271531,I2507,I759644,I759871,);
nor I_44549 (I759879,I759871,I759738);
not I_44550 (I759896,I759879);
not I_44551 (I759913,I759871);
nor I_44552 (I759930,I759913,I759814);
DFFARX1 I_44553 (I759930,I2507,I759644,I759630,);
nand I_44554 (I759961,I1271537,I1271525);
and I_44555 (I759978,I759961,I1271519);
DFFARX1 I_44556 (I759978,I2507,I759644,I760004,);
nor I_44557 (I760012,I760004,I759871);
DFFARX1 I_44558 (I760012,I2507,I759644,I759612,);
nand I_44559 (I760043,I760004,I759913);
nand I_44560 (I759621,I759896,I760043);
not I_44561 (I760074,I760004);
nor I_44562 (I760091,I760074,I759814);
DFFARX1 I_44563 (I760091,I2507,I759644,I759633,);
nor I_44564 (I760122,I1271516,I1271525);
or I_44565 (I759624,I759871,I760122);
nor I_44566 (I759615,I760004,I760122);
or I_44567 (I759618,I759738,I760122);
DFFARX1 I_44568 (I760122,I2507,I759644,I759636,);
not I_44569 (I760222,I2514);
DFFARX1 I_44570 (I1145088,I2507,I760222,I760248,);
not I_44571 (I760256,I760248);
nand I_44572 (I760273,I1145070,I1145082);
and I_44573 (I760290,I760273,I1145085);
DFFARX1 I_44574 (I760290,I2507,I760222,I760316,);
not I_44575 (I760324,I1145079);
DFFARX1 I_44576 (I1145076,I2507,I760222,I760350,);
not I_44577 (I760358,I760350);
nor I_44578 (I760375,I760358,I760256);
and I_44579 (I760392,I760375,I1145079);
nor I_44580 (I760409,I760358,I760324);
nor I_44581 (I760205,I760316,I760409);
DFFARX1 I_44582 (I1145094,I2507,I760222,I760449,);
nor I_44583 (I760457,I760449,I760316);
not I_44584 (I760474,I760457);
not I_44585 (I760491,I760449);
nor I_44586 (I760508,I760491,I760392);
DFFARX1 I_44587 (I760508,I2507,I760222,I760208,);
nand I_44588 (I760539,I1145073,I1145073);
and I_44589 (I760556,I760539,I1145070);
DFFARX1 I_44590 (I760556,I2507,I760222,I760582,);
nor I_44591 (I760590,I760582,I760449);
DFFARX1 I_44592 (I760590,I2507,I760222,I760190,);
nand I_44593 (I760621,I760582,I760491);
nand I_44594 (I760199,I760474,I760621);
not I_44595 (I760652,I760582);
nor I_44596 (I760669,I760652,I760392);
DFFARX1 I_44597 (I760669,I2507,I760222,I760211,);
nor I_44598 (I760700,I1145091,I1145073);
or I_44599 (I760202,I760449,I760700);
nor I_44600 (I760193,I760582,I760700);
or I_44601 (I760196,I760316,I760700);
DFFARX1 I_44602 (I760700,I2507,I760222,I760214,);
not I_44603 (I760800,I2514);
DFFARX1 I_44604 (I435448,I2507,I760800,I760826,);
not I_44605 (I760834,I760826);
nand I_44606 (I760851,I435439,I435457);
and I_44607 (I760868,I760851,I435460);
DFFARX1 I_44608 (I760868,I2507,I760800,I760894,);
not I_44609 (I760902,I435454);
DFFARX1 I_44610 (I435442,I2507,I760800,I760928,);
not I_44611 (I760936,I760928);
nor I_44612 (I760953,I760936,I760834);
and I_44613 (I760970,I760953,I435454);
nor I_44614 (I760987,I760936,I760902);
nor I_44615 (I760783,I760894,I760987);
DFFARX1 I_44616 (I435451,I2507,I760800,I761027,);
nor I_44617 (I761035,I761027,I760894);
not I_44618 (I761052,I761035);
not I_44619 (I761069,I761027);
nor I_44620 (I761086,I761069,I760970);
DFFARX1 I_44621 (I761086,I2507,I760800,I760786,);
nand I_44622 (I761117,I435466,I435463);
and I_44623 (I761134,I761117,I435445);
DFFARX1 I_44624 (I761134,I2507,I760800,I761160,);
nor I_44625 (I761168,I761160,I761027);
DFFARX1 I_44626 (I761168,I2507,I760800,I760768,);
nand I_44627 (I761199,I761160,I761069);
nand I_44628 (I760777,I761052,I761199);
not I_44629 (I761230,I761160);
nor I_44630 (I761247,I761230,I760970);
DFFARX1 I_44631 (I761247,I2507,I760800,I760789,);
nor I_44632 (I761278,I435439,I435463);
or I_44633 (I760780,I761027,I761278);
nor I_44634 (I760771,I761160,I761278);
or I_44635 (I760774,I760894,I761278);
DFFARX1 I_44636 (I761278,I2507,I760800,I760792,);
not I_44637 (I761378,I2514);
DFFARX1 I_44638 (I1716,I2507,I761378,I761404,);
not I_44639 (I761412,I761404);
nand I_44640 (I761429,I2476,I2036);
and I_44641 (I761446,I761429,I1388);
DFFARX1 I_44642 (I761446,I2507,I761378,I761472,);
not I_44643 (I761480,I1404);
DFFARX1 I_44644 (I2212,I2507,I761378,I761506,);
not I_44645 (I761514,I761506);
nor I_44646 (I761531,I761514,I761412);
and I_44647 (I761548,I761531,I1404);
nor I_44648 (I761565,I761514,I761480);
nor I_44649 (I761361,I761472,I761565);
DFFARX1 I_44650 (I1772,I2507,I761378,I761605,);
nor I_44651 (I761613,I761605,I761472);
not I_44652 (I761630,I761613);
not I_44653 (I761647,I761605);
nor I_44654 (I761664,I761647,I761548);
DFFARX1 I_44655 (I761664,I2507,I761378,I761364,);
nand I_44656 (I761695,I2004,I1604);
and I_44657 (I761712,I761695,I2188);
DFFARX1 I_44658 (I761712,I2507,I761378,I761738,);
nor I_44659 (I761746,I761738,I761605);
DFFARX1 I_44660 (I761746,I2507,I761378,I761346,);
nand I_44661 (I761777,I761738,I761647);
nand I_44662 (I761355,I761630,I761777);
not I_44663 (I761808,I761738);
nor I_44664 (I761825,I761808,I761548);
DFFARX1 I_44665 (I761825,I2507,I761378,I761367,);
nor I_44666 (I761856,I1940,I1604);
or I_44667 (I761358,I761605,I761856);
nor I_44668 (I761349,I761738,I761856);
or I_44669 (I761352,I761472,I761856);
DFFARX1 I_44670 (I761856,I2507,I761378,I761370,);
not I_44671 (I761956,I2514);
DFFARX1 I_44672 (I800155,I2507,I761956,I761982,);
not I_44673 (I761990,I761982);
nand I_44674 (I762007,I800143,I800161);
and I_44675 (I762024,I762007,I800158);
DFFARX1 I_44676 (I762024,I2507,I761956,I762050,);
not I_44677 (I762058,I800149);
DFFARX1 I_44678 (I800146,I2507,I761956,I762084,);
not I_44679 (I762092,I762084);
nor I_44680 (I762109,I762092,I761990);
and I_44681 (I762126,I762109,I800149);
nor I_44682 (I762143,I762092,I762058);
nor I_44683 (I761939,I762050,I762143);
DFFARX1 I_44684 (I800140,I2507,I761956,I762183,);
nor I_44685 (I762191,I762183,I762050);
not I_44686 (I762208,I762191);
not I_44687 (I762225,I762183);
nor I_44688 (I762242,I762225,I762126);
DFFARX1 I_44689 (I762242,I2507,I761956,I761942,);
nand I_44690 (I762273,I800140,I800143);
and I_44691 (I762290,I762273,I800146);
DFFARX1 I_44692 (I762290,I2507,I761956,I762316,);
nor I_44693 (I762324,I762316,I762183);
DFFARX1 I_44694 (I762324,I2507,I761956,I761924,);
nand I_44695 (I762355,I762316,I762225);
nand I_44696 (I761933,I762208,I762355);
not I_44697 (I762386,I762316);
nor I_44698 (I762403,I762386,I762126);
DFFARX1 I_44699 (I762403,I2507,I761956,I761945,);
nor I_44700 (I762434,I800152,I800143);
or I_44701 (I761936,I762183,I762434);
nor I_44702 (I761927,I762316,I762434);
or I_44703 (I761930,I762050,I762434);
DFFARX1 I_44704 (I762434,I2507,I761956,I761948,);
not I_44705 (I762534,I2514);
DFFARX1 I_44706 (I836518,I2507,I762534,I762560,);
not I_44707 (I762568,I762560);
nand I_44708 (I762585,I836506,I836524);
and I_44709 (I762602,I762585,I836521);
DFFARX1 I_44710 (I762602,I2507,I762534,I762628,);
not I_44711 (I762636,I836512);
DFFARX1 I_44712 (I836509,I2507,I762534,I762662,);
not I_44713 (I762670,I762662);
nor I_44714 (I762687,I762670,I762568);
and I_44715 (I762704,I762687,I836512);
nor I_44716 (I762721,I762670,I762636);
nor I_44717 (I762517,I762628,I762721);
DFFARX1 I_44718 (I836503,I2507,I762534,I762761,);
nor I_44719 (I762769,I762761,I762628);
not I_44720 (I762786,I762769);
not I_44721 (I762803,I762761);
nor I_44722 (I762820,I762803,I762704);
DFFARX1 I_44723 (I762820,I2507,I762534,I762520,);
nand I_44724 (I762851,I836503,I836506);
and I_44725 (I762868,I762851,I836509);
DFFARX1 I_44726 (I762868,I2507,I762534,I762894,);
nor I_44727 (I762902,I762894,I762761);
DFFARX1 I_44728 (I762902,I2507,I762534,I762502,);
nand I_44729 (I762933,I762894,I762803);
nand I_44730 (I762511,I762786,I762933);
not I_44731 (I762964,I762894);
nor I_44732 (I762981,I762964,I762704);
DFFARX1 I_44733 (I762981,I2507,I762534,I762523,);
nor I_44734 (I763012,I836515,I836506);
or I_44735 (I762514,I762761,I763012);
nor I_44736 (I762505,I762894,I763012);
or I_44737 (I762508,I762628,I763012);
DFFARX1 I_44738 (I763012,I2507,I762534,I762526,);
not I_44739 (I763112,I2514);
DFFARX1 I_44740 (I107563,I2507,I763112,I763138,);
not I_44741 (I763146,I763138);
nand I_44742 (I763163,I107572,I107581);
and I_44743 (I763180,I763163,I107560);
DFFARX1 I_44744 (I763180,I2507,I763112,I763206,);
not I_44745 (I763214,I107563);
DFFARX1 I_44746 (I107578,I2507,I763112,I763240,);
not I_44747 (I763248,I763240);
nor I_44748 (I763265,I763248,I763146);
and I_44749 (I763282,I763265,I107563);
nor I_44750 (I763299,I763248,I763214);
nor I_44751 (I763095,I763206,I763299);
DFFARX1 I_44752 (I107569,I2507,I763112,I763339,);
nor I_44753 (I763347,I763339,I763206);
not I_44754 (I763364,I763347);
not I_44755 (I763381,I763339);
nor I_44756 (I763398,I763381,I763282);
DFFARX1 I_44757 (I763398,I2507,I763112,I763098,);
nand I_44758 (I763429,I107584,I107560);
and I_44759 (I763446,I763429,I107566);
DFFARX1 I_44760 (I763446,I2507,I763112,I763472,);
nor I_44761 (I763480,I763472,I763339);
DFFARX1 I_44762 (I763480,I2507,I763112,I763080,);
nand I_44763 (I763511,I763472,I763381);
nand I_44764 (I763089,I763364,I763511);
not I_44765 (I763542,I763472);
nor I_44766 (I763559,I763542,I763282);
DFFARX1 I_44767 (I763559,I2507,I763112,I763101,);
nor I_44768 (I763590,I107575,I107560);
or I_44769 (I763092,I763339,I763590);
nor I_44770 (I763083,I763472,I763590);
or I_44771 (I763086,I763206,I763590);
DFFARX1 I_44772 (I763590,I2507,I763112,I763104,);
not I_44773 (I763690,I2514);
DFFARX1 I_44774 (I160940,I2507,I763690,I763716,);
not I_44775 (I763724,I763716);
nand I_44776 (I763741,I160943,I160964);
and I_44777 (I763758,I763741,I160952);
DFFARX1 I_44778 (I763758,I2507,I763690,I763784,);
not I_44779 (I763792,I160949);
DFFARX1 I_44780 (I160940,I2507,I763690,I763818,);
not I_44781 (I763826,I763818);
nor I_44782 (I763843,I763826,I763724);
and I_44783 (I763860,I763843,I160949);
nor I_44784 (I763877,I763826,I763792);
nor I_44785 (I763673,I763784,I763877);
DFFARX1 I_44786 (I160958,I2507,I763690,I763917,);
nor I_44787 (I763925,I763917,I763784);
not I_44788 (I763942,I763925);
not I_44789 (I763959,I763917);
nor I_44790 (I763976,I763959,I763860);
DFFARX1 I_44791 (I763976,I2507,I763690,I763676,);
nand I_44792 (I764007,I160943,I160946);
and I_44793 (I764024,I764007,I160955);
DFFARX1 I_44794 (I764024,I2507,I763690,I764050,);
nor I_44795 (I764058,I764050,I763917);
DFFARX1 I_44796 (I764058,I2507,I763690,I763658,);
nand I_44797 (I764089,I764050,I763959);
nand I_44798 (I763667,I763942,I764089);
not I_44799 (I764120,I764050);
nor I_44800 (I764137,I764120,I763860);
DFFARX1 I_44801 (I764137,I2507,I763690,I763679,);
nor I_44802 (I764168,I160961,I160946);
or I_44803 (I763670,I763917,I764168);
nor I_44804 (I763661,I764050,I764168);
or I_44805 (I763664,I763784,I764168);
DFFARX1 I_44806 (I764168,I2507,I763690,I763682,);
not I_44807 (I764268,I2514);
DFFARX1 I_44808 (I94388,I2507,I764268,I764294,);
not I_44809 (I764302,I764294);
nand I_44810 (I764319,I94397,I94406);
and I_44811 (I764336,I764319,I94385);
DFFARX1 I_44812 (I764336,I2507,I764268,I764362,);
not I_44813 (I764370,I94388);
DFFARX1 I_44814 (I94403,I2507,I764268,I764396,);
not I_44815 (I764404,I764396);
nor I_44816 (I764421,I764404,I764302);
and I_44817 (I764438,I764421,I94388);
nor I_44818 (I764455,I764404,I764370);
nor I_44819 (I764251,I764362,I764455);
DFFARX1 I_44820 (I94394,I2507,I764268,I764495,);
nor I_44821 (I764503,I764495,I764362);
not I_44822 (I764520,I764503);
not I_44823 (I764537,I764495);
nor I_44824 (I764554,I764537,I764438);
DFFARX1 I_44825 (I764554,I2507,I764268,I764254,);
nand I_44826 (I764585,I94409,I94385);
and I_44827 (I764602,I764585,I94391);
DFFARX1 I_44828 (I764602,I2507,I764268,I764628,);
nor I_44829 (I764636,I764628,I764495);
DFFARX1 I_44830 (I764636,I2507,I764268,I764236,);
nand I_44831 (I764667,I764628,I764537);
nand I_44832 (I764245,I764520,I764667);
not I_44833 (I764698,I764628);
nor I_44834 (I764715,I764698,I764438);
DFFARX1 I_44835 (I764715,I2507,I764268,I764257,);
nor I_44836 (I764746,I94400,I94385);
or I_44837 (I764248,I764495,I764746);
nor I_44838 (I764239,I764628,I764746);
or I_44839 (I764242,I764362,I764746);
DFFARX1 I_44840 (I764746,I2507,I764268,I764260,);
not I_44841 (I764846,I2514);
DFFARX1 I_44842 (I986433,I2507,I764846,I764872,);
not I_44843 (I764880,I764872);
nand I_44844 (I764897,I986409,I986424);
and I_44845 (I764914,I764897,I986436);
DFFARX1 I_44846 (I764914,I2507,I764846,I764940,);
not I_44847 (I764948,I986421);
DFFARX1 I_44848 (I986412,I2507,I764846,I764974,);
not I_44849 (I764982,I764974);
nor I_44850 (I764999,I764982,I764880);
and I_44851 (I765016,I764999,I986421);
nor I_44852 (I765033,I764982,I764948);
nor I_44853 (I764829,I764940,I765033);
DFFARX1 I_44854 (I986409,I2507,I764846,I765073,);
nor I_44855 (I765081,I765073,I764940);
not I_44856 (I765098,I765081);
not I_44857 (I765115,I765073);
nor I_44858 (I765132,I765115,I765016);
DFFARX1 I_44859 (I765132,I2507,I764846,I764832,);
nand I_44860 (I765163,I986427,I986418);
and I_44861 (I765180,I765163,I986430);
DFFARX1 I_44862 (I765180,I2507,I764846,I765206,);
nor I_44863 (I765214,I765206,I765073);
DFFARX1 I_44864 (I765214,I2507,I764846,I764814,);
nand I_44865 (I765245,I765206,I765115);
nand I_44866 (I764823,I765098,I765245);
not I_44867 (I765276,I765206);
nor I_44868 (I765293,I765276,I765016);
DFFARX1 I_44869 (I765293,I2507,I764846,I764835,);
nor I_44870 (I765324,I986415,I986418);
or I_44871 (I764826,I765073,I765324);
nor I_44872 (I764817,I765206,I765324);
or I_44873 (I764820,I764940,I765324);
DFFARX1 I_44874 (I765324,I2507,I764846,I764838,);
not I_44875 (I765424,I2514);
DFFARX1 I_44876 (I422936,I2507,I765424,I765450,);
not I_44877 (I765458,I765450);
nand I_44878 (I765475,I422927,I422945);
and I_44879 (I765492,I765475,I422948);
DFFARX1 I_44880 (I765492,I2507,I765424,I765518,);
not I_44881 (I765526,I422942);
DFFARX1 I_44882 (I422930,I2507,I765424,I765552,);
not I_44883 (I765560,I765552);
nor I_44884 (I765577,I765560,I765458);
and I_44885 (I765594,I765577,I422942);
nor I_44886 (I765611,I765560,I765526);
nor I_44887 (I765407,I765518,I765611);
DFFARX1 I_44888 (I422939,I2507,I765424,I765651,);
nor I_44889 (I765659,I765651,I765518);
not I_44890 (I765676,I765659);
not I_44891 (I765693,I765651);
nor I_44892 (I765710,I765693,I765594);
DFFARX1 I_44893 (I765710,I2507,I765424,I765410,);
nand I_44894 (I765741,I422954,I422951);
and I_44895 (I765758,I765741,I422933);
DFFARX1 I_44896 (I765758,I2507,I765424,I765784,);
nor I_44897 (I765792,I765784,I765651);
DFFARX1 I_44898 (I765792,I2507,I765424,I765392,);
nand I_44899 (I765823,I765784,I765693);
nand I_44900 (I765401,I765676,I765823);
not I_44901 (I765854,I765784);
nor I_44902 (I765871,I765854,I765594);
DFFARX1 I_44903 (I765871,I2507,I765424,I765413,);
nor I_44904 (I765902,I422927,I422951);
or I_44905 (I765404,I765651,I765902);
nor I_44906 (I765395,I765784,I765902);
or I_44907 (I765398,I765518,I765902);
DFFARX1 I_44908 (I765902,I2507,I765424,I765416,);
not I_44909 (I766002,I2514);
DFFARX1 I_44910 (I878678,I2507,I766002,I766028,);
not I_44911 (I766036,I766028);
nand I_44912 (I766053,I878666,I878684);
and I_44913 (I766070,I766053,I878681);
DFFARX1 I_44914 (I766070,I2507,I766002,I766096,);
not I_44915 (I766104,I878672);
DFFARX1 I_44916 (I878669,I2507,I766002,I766130,);
not I_44917 (I766138,I766130);
nor I_44918 (I766155,I766138,I766036);
and I_44919 (I766172,I766155,I878672);
nor I_44920 (I766189,I766138,I766104);
nor I_44921 (I765985,I766096,I766189);
DFFARX1 I_44922 (I878663,I2507,I766002,I766229,);
nor I_44923 (I766237,I766229,I766096);
not I_44924 (I766254,I766237);
not I_44925 (I766271,I766229);
nor I_44926 (I766288,I766271,I766172);
DFFARX1 I_44927 (I766288,I2507,I766002,I765988,);
nand I_44928 (I766319,I878663,I878666);
and I_44929 (I766336,I766319,I878669);
DFFARX1 I_44930 (I766336,I2507,I766002,I766362,);
nor I_44931 (I766370,I766362,I766229);
DFFARX1 I_44932 (I766370,I2507,I766002,I765970,);
nand I_44933 (I766401,I766362,I766271);
nand I_44934 (I765979,I766254,I766401);
not I_44935 (I766432,I766362);
nor I_44936 (I766449,I766432,I766172);
DFFARX1 I_44937 (I766449,I2507,I766002,I765991,);
nor I_44938 (I766480,I878675,I878666);
or I_44939 (I765982,I766229,I766480);
nor I_44940 (I765973,I766362,I766480);
or I_44941 (I765976,I766096,I766480);
DFFARX1 I_44942 (I766480,I2507,I766002,I765994,);
not I_44943 (I766580,I2514);
DFFARX1 I_44944 (I1007105,I2507,I766580,I766606,);
not I_44945 (I766614,I766606);
nand I_44946 (I766631,I1007081,I1007096);
and I_44947 (I766648,I766631,I1007108);
DFFARX1 I_44948 (I766648,I2507,I766580,I766674,);
not I_44949 (I766682,I1007093);
DFFARX1 I_44950 (I1007084,I2507,I766580,I766708,);
not I_44951 (I766716,I766708);
nor I_44952 (I766733,I766716,I766614);
and I_44953 (I766750,I766733,I1007093);
nor I_44954 (I766767,I766716,I766682);
nor I_44955 (I766563,I766674,I766767);
DFFARX1 I_44956 (I1007081,I2507,I766580,I766807,);
nor I_44957 (I766815,I766807,I766674);
not I_44958 (I766832,I766815);
not I_44959 (I766849,I766807);
nor I_44960 (I766866,I766849,I766750);
DFFARX1 I_44961 (I766866,I2507,I766580,I766566,);
nand I_44962 (I766897,I1007099,I1007090);
and I_44963 (I766914,I766897,I1007102);
DFFARX1 I_44964 (I766914,I2507,I766580,I766940,);
nor I_44965 (I766948,I766940,I766807);
DFFARX1 I_44966 (I766948,I2507,I766580,I766548,);
nand I_44967 (I766979,I766940,I766849);
nand I_44968 (I766557,I766832,I766979);
not I_44969 (I767010,I766940);
nor I_44970 (I767027,I767010,I766750);
DFFARX1 I_44971 (I767027,I2507,I766580,I766569,);
nor I_44972 (I767058,I1007087,I1007090);
or I_44973 (I766560,I766807,I767058);
nor I_44974 (I766551,I766940,I767058);
or I_44975 (I766554,I766674,I767058);
DFFARX1 I_44976 (I767058,I2507,I766580,I766572,);
not I_44977 (I767158,I2514);
DFFARX1 I_44978 (I241860,I2507,I767158,I767184,);
not I_44979 (I767192,I767184);
nand I_44980 (I767209,I241863,I241884);
and I_44981 (I767226,I767209,I241872);
DFFARX1 I_44982 (I767226,I2507,I767158,I767252,);
not I_44983 (I767260,I241869);
DFFARX1 I_44984 (I241860,I2507,I767158,I767286,);
not I_44985 (I767294,I767286);
nor I_44986 (I767311,I767294,I767192);
and I_44987 (I767328,I767311,I241869);
nor I_44988 (I767345,I767294,I767260);
nor I_44989 (I767141,I767252,I767345);
DFFARX1 I_44990 (I241878,I2507,I767158,I767385,);
nor I_44991 (I767393,I767385,I767252);
not I_44992 (I767410,I767393);
not I_44993 (I767427,I767385);
nor I_44994 (I767444,I767427,I767328);
DFFARX1 I_44995 (I767444,I2507,I767158,I767144,);
nand I_44996 (I767475,I241863,I241866);
and I_44997 (I767492,I767475,I241875);
DFFARX1 I_44998 (I767492,I2507,I767158,I767518,);
nor I_44999 (I767526,I767518,I767385);
DFFARX1 I_45000 (I767526,I2507,I767158,I767126,);
nand I_45001 (I767557,I767518,I767427);
nand I_45002 (I767135,I767410,I767557);
not I_45003 (I767588,I767518);
nor I_45004 (I767605,I767588,I767328);
DFFARX1 I_45005 (I767605,I2507,I767158,I767147,);
nor I_45006 (I767636,I241881,I241866);
or I_45007 (I767138,I767385,I767636);
nor I_45008 (I767129,I767518,I767636);
or I_45009 (I767132,I767252,I767636);
DFFARX1 I_45010 (I767636,I2507,I767158,I767150,);
not I_45011 (I767736,I2514);
DFFARX1 I_45012 (I439256,I2507,I767736,I767762,);
not I_45013 (I767770,I767762);
nand I_45014 (I767787,I439247,I439265);
and I_45015 (I767804,I767787,I439268);
DFFARX1 I_45016 (I767804,I2507,I767736,I767830,);
not I_45017 (I767838,I439262);
DFFARX1 I_45018 (I439250,I2507,I767736,I767864,);
not I_45019 (I767872,I767864);
nor I_45020 (I767889,I767872,I767770);
and I_45021 (I767906,I767889,I439262);
nor I_45022 (I767923,I767872,I767838);
nor I_45023 (I767719,I767830,I767923);
DFFARX1 I_45024 (I439259,I2507,I767736,I767963,);
nor I_45025 (I767971,I767963,I767830);
not I_45026 (I767988,I767971);
not I_45027 (I768005,I767963);
nor I_45028 (I768022,I768005,I767906);
DFFARX1 I_45029 (I768022,I2507,I767736,I767722,);
nand I_45030 (I768053,I439274,I439271);
and I_45031 (I768070,I768053,I439253);
DFFARX1 I_45032 (I768070,I2507,I767736,I768096,);
nor I_45033 (I768104,I768096,I767963);
DFFARX1 I_45034 (I768104,I2507,I767736,I767704,);
nand I_45035 (I768135,I768096,I768005);
nand I_45036 (I767713,I767988,I768135);
not I_45037 (I768166,I768096);
nor I_45038 (I768183,I768166,I767906);
DFFARX1 I_45039 (I768183,I2507,I767736,I767725,);
nor I_45040 (I768214,I439247,I439271);
or I_45041 (I767716,I767963,I768214);
nor I_45042 (I767707,I768096,I768214);
or I_45043 (I767710,I767830,I768214);
DFFARX1 I_45044 (I768214,I2507,I767736,I767728,);
not I_45045 (I768314,I2514);
DFFARX1 I_45046 (I1068214,I2507,I768314,I768340,);
not I_45047 (I768348,I768340);
nand I_45048 (I768365,I1068196,I1068208);
and I_45049 (I768382,I768365,I1068211);
DFFARX1 I_45050 (I768382,I2507,I768314,I768408,);
not I_45051 (I768416,I1068205);
DFFARX1 I_45052 (I1068202,I2507,I768314,I768442,);
not I_45053 (I768450,I768442);
nor I_45054 (I768467,I768450,I768348);
and I_45055 (I768484,I768467,I1068205);
nor I_45056 (I768501,I768450,I768416);
nor I_45057 (I768297,I768408,I768501);
DFFARX1 I_45058 (I1068220,I2507,I768314,I768541,);
nor I_45059 (I768549,I768541,I768408);
not I_45060 (I768566,I768549);
not I_45061 (I768583,I768541);
nor I_45062 (I768600,I768583,I768484);
DFFARX1 I_45063 (I768600,I2507,I768314,I768300,);
nand I_45064 (I768631,I1068199,I1068199);
and I_45065 (I768648,I768631,I1068196);
DFFARX1 I_45066 (I768648,I2507,I768314,I768674,);
nor I_45067 (I768682,I768674,I768541);
DFFARX1 I_45068 (I768682,I2507,I768314,I768282,);
nand I_45069 (I768713,I768674,I768583);
nand I_45070 (I768291,I768566,I768713);
not I_45071 (I768744,I768674);
nor I_45072 (I768761,I768744,I768484);
DFFARX1 I_45073 (I768761,I2507,I768314,I768303,);
nor I_45074 (I768792,I1068217,I1068199);
or I_45075 (I768294,I768541,I768792);
nor I_45076 (I768285,I768674,I768792);
or I_45077 (I768288,I768408,I768792);
DFFARX1 I_45078 (I768792,I2507,I768314,I768306,);
not I_45079 (I768892,I2514);
DFFARX1 I_45080 (I1049978,I2507,I768892,I768918,);
not I_45081 (I768926,I768918);
nand I_45082 (I768943,I1049975,I1049993);
and I_45083 (I768960,I768943,I1049990);
DFFARX1 I_45084 (I768960,I2507,I768892,I768986,);
not I_45085 (I768994,I1049972);
DFFARX1 I_45086 (I1049975,I2507,I768892,I769020,);
not I_45087 (I769028,I769020);
nor I_45088 (I769045,I769028,I768926);
and I_45089 (I769062,I769045,I1049972);
nor I_45090 (I769079,I769028,I768994);
nor I_45091 (I768875,I768986,I769079);
DFFARX1 I_45092 (I1049984,I2507,I768892,I769119,);
nor I_45093 (I769127,I769119,I768986);
not I_45094 (I769144,I769127);
not I_45095 (I769161,I769119);
nor I_45096 (I769178,I769161,I769062);
DFFARX1 I_45097 (I769178,I2507,I768892,I768878,);
nand I_45098 (I769209,I1049987,I1049972);
and I_45099 (I769226,I769209,I1049978);
DFFARX1 I_45100 (I769226,I2507,I768892,I769252,);
nor I_45101 (I769260,I769252,I769119);
DFFARX1 I_45102 (I769260,I2507,I768892,I768860,);
nand I_45103 (I769291,I769252,I769161);
nand I_45104 (I768869,I769144,I769291);
not I_45105 (I769322,I769252);
nor I_45106 (I769339,I769322,I769062);
DFFARX1 I_45107 (I769339,I2507,I768892,I768881,);
nor I_45108 (I769370,I1049981,I1049972);
or I_45109 (I768872,I769119,I769370);
nor I_45110 (I768863,I769252,I769370);
or I_45111 (I768866,I768986,I769370);
DFFARX1 I_45112 (I769370,I2507,I768892,I768884,);
not I_45113 (I769470,I2514);
DFFARX1 I_45114 (I544018,I2507,I769470,I769496,);
not I_45115 (I769504,I769496);
nand I_45116 (I769521,I544027,I544036);
and I_45117 (I769538,I769521,I544042);
DFFARX1 I_45118 (I769538,I2507,I769470,I769564,);
not I_45119 (I769572,I544039);
DFFARX1 I_45120 (I544024,I2507,I769470,I769598,);
not I_45121 (I769606,I769598);
nor I_45122 (I769623,I769606,I769504);
and I_45123 (I769640,I769623,I544039);
nor I_45124 (I769657,I769606,I769572);
nor I_45125 (I769453,I769564,I769657);
DFFARX1 I_45126 (I544033,I2507,I769470,I769697,);
nor I_45127 (I769705,I769697,I769564);
not I_45128 (I769722,I769705);
not I_45129 (I769739,I769697);
nor I_45130 (I769756,I769739,I769640);
DFFARX1 I_45131 (I769756,I2507,I769470,I769456,);
nand I_45132 (I769787,I544030,I544021);
and I_45133 (I769804,I769787,I544018);
DFFARX1 I_45134 (I769804,I2507,I769470,I769830,);
nor I_45135 (I769838,I769830,I769697);
DFFARX1 I_45136 (I769838,I2507,I769470,I769438,);
nand I_45137 (I769869,I769830,I769739);
nand I_45138 (I769447,I769722,I769869);
not I_45139 (I769900,I769830);
nor I_45140 (I769917,I769900,I769640);
DFFARX1 I_45141 (I769917,I2507,I769470,I769459,);
nor I_45142 (I769948,I544021,I544021);
or I_45143 (I769450,I769697,I769948);
nor I_45144 (I769441,I769830,I769948);
or I_45145 (I769444,I769564,I769948);
DFFARX1 I_45146 (I769948,I2507,I769470,I769462,);
not I_45147 (I770048,I2514);
DFFARX1 I_45148 (I872354,I2507,I770048,I770074,);
not I_45149 (I770082,I770074);
nand I_45150 (I770099,I872342,I872360);
and I_45151 (I770116,I770099,I872357);
DFFARX1 I_45152 (I770116,I2507,I770048,I770142,);
not I_45153 (I770150,I872348);
DFFARX1 I_45154 (I872345,I2507,I770048,I770176,);
not I_45155 (I770184,I770176);
nor I_45156 (I770201,I770184,I770082);
and I_45157 (I770218,I770201,I872348);
nor I_45158 (I770235,I770184,I770150);
nor I_45159 (I770031,I770142,I770235);
DFFARX1 I_45160 (I872339,I2507,I770048,I770275,);
nor I_45161 (I770283,I770275,I770142);
not I_45162 (I770300,I770283);
not I_45163 (I770317,I770275);
nor I_45164 (I770334,I770317,I770218);
DFFARX1 I_45165 (I770334,I2507,I770048,I770034,);
nand I_45166 (I770365,I872339,I872342);
and I_45167 (I770382,I770365,I872345);
DFFARX1 I_45168 (I770382,I2507,I770048,I770408,);
nor I_45169 (I770416,I770408,I770275);
DFFARX1 I_45170 (I770416,I2507,I770048,I770016,);
nand I_45171 (I770447,I770408,I770317);
nand I_45172 (I770025,I770300,I770447);
not I_45173 (I770478,I770408);
nor I_45174 (I770495,I770478,I770218);
DFFARX1 I_45175 (I770495,I2507,I770048,I770037,);
nor I_45176 (I770526,I872351,I872342);
or I_45177 (I770028,I770275,I770526);
nor I_45178 (I770019,I770408,I770526);
or I_45179 (I770022,I770142,I770526);
DFFARX1 I_45180 (I770526,I2507,I770048,I770040,);
not I_45181 (I770626,I2514);
DFFARX1 I_45182 (I510749,I2507,I770626,I770652,);
not I_45183 (I770660,I770652);
nand I_45184 (I770677,I510764,I510749);
and I_45185 (I770694,I770677,I510752);
DFFARX1 I_45186 (I770694,I2507,I770626,I770720,);
not I_45187 (I770728,I510752);
DFFARX1 I_45188 (I510761,I2507,I770626,I770754,);
not I_45189 (I770762,I770754);
nor I_45190 (I770779,I770762,I770660);
and I_45191 (I770796,I770779,I510752);
nor I_45192 (I770813,I770762,I770728);
nor I_45193 (I770609,I770720,I770813);
DFFARX1 I_45194 (I510755,I2507,I770626,I770853,);
nor I_45195 (I770861,I770853,I770720);
not I_45196 (I770878,I770861);
not I_45197 (I770895,I770853);
nor I_45198 (I770912,I770895,I770796);
DFFARX1 I_45199 (I770912,I2507,I770626,I770612,);
nand I_45200 (I770943,I510758,I510767);
and I_45201 (I770960,I770943,I510773);
DFFARX1 I_45202 (I770960,I2507,I770626,I770986,);
nor I_45203 (I770994,I770986,I770853);
DFFARX1 I_45204 (I770994,I2507,I770626,I770594,);
nand I_45205 (I771025,I770986,I770895);
nand I_45206 (I770603,I770878,I771025);
not I_45207 (I771056,I770986);
nor I_45208 (I771073,I771056,I770796);
DFFARX1 I_45209 (I771073,I2507,I770626,I770615,);
nor I_45210 (I771104,I510770,I510767);
or I_45211 (I770606,I770853,I771104);
nor I_45212 (I770597,I770986,I771104);
or I_45213 (I770600,I770720,I771104);
DFFARX1 I_45214 (I771104,I2507,I770626,I770618,);
not I_45215 (I771204,I2514);
DFFARX1 I_45216 (I501824,I2507,I771204,I771230,);
not I_45217 (I771238,I771230);
nand I_45218 (I771255,I501839,I501824);
and I_45219 (I771272,I771255,I501827);
DFFARX1 I_45220 (I771272,I2507,I771204,I771298,);
not I_45221 (I771306,I501827);
DFFARX1 I_45222 (I501836,I2507,I771204,I771332,);
not I_45223 (I771340,I771332);
nor I_45224 (I771357,I771340,I771238);
and I_45225 (I771374,I771357,I501827);
nor I_45226 (I771391,I771340,I771306);
nor I_45227 (I771187,I771298,I771391);
DFFARX1 I_45228 (I501830,I2507,I771204,I771431,);
nor I_45229 (I771439,I771431,I771298);
not I_45230 (I771456,I771439);
not I_45231 (I771473,I771431);
nor I_45232 (I771490,I771473,I771374);
DFFARX1 I_45233 (I771490,I2507,I771204,I771190,);
nand I_45234 (I771521,I501833,I501842);
and I_45235 (I771538,I771521,I501848);
DFFARX1 I_45236 (I771538,I2507,I771204,I771564,);
nor I_45237 (I771572,I771564,I771431);
DFFARX1 I_45238 (I771572,I2507,I771204,I771172,);
nand I_45239 (I771603,I771564,I771473);
nand I_45240 (I771181,I771456,I771603);
not I_45241 (I771634,I771564);
nor I_45242 (I771651,I771634,I771374);
DFFARX1 I_45243 (I771651,I2507,I771204,I771193,);
nor I_45244 (I771682,I501845,I501842);
or I_45245 (I771184,I771431,I771682);
nor I_45246 (I771175,I771564,I771682);
or I_45247 (I771178,I771298,I771682);
DFFARX1 I_45248 (I771682,I2507,I771204,I771196,);
not I_45249 (I771782,I2514);
DFFARX1 I_45250 (I251795,I2507,I771782,I771808,);
not I_45251 (I771816,I771808);
nand I_45252 (I771833,I251798,I251774);
and I_45253 (I771850,I771833,I251771);
DFFARX1 I_45254 (I771850,I2507,I771782,I771876,);
not I_45255 (I771884,I251777);
DFFARX1 I_45256 (I251771,I2507,I771782,I771910,);
not I_45257 (I771918,I771910);
nor I_45258 (I771935,I771918,I771816);
and I_45259 (I771952,I771935,I251777);
nor I_45260 (I771969,I771918,I771884);
nor I_45261 (I771765,I771876,I771969);
DFFARX1 I_45262 (I251780,I2507,I771782,I772009,);
nor I_45263 (I772017,I772009,I771876);
not I_45264 (I772034,I772017);
not I_45265 (I772051,I772009);
nor I_45266 (I772068,I772051,I771952);
DFFARX1 I_45267 (I772068,I2507,I771782,I771768,);
nand I_45268 (I772099,I251783,I251792);
and I_45269 (I772116,I772099,I251789);
DFFARX1 I_45270 (I772116,I2507,I771782,I772142,);
nor I_45271 (I772150,I772142,I772009);
DFFARX1 I_45272 (I772150,I2507,I771782,I771750,);
nand I_45273 (I772181,I772142,I772051);
nand I_45274 (I771759,I772034,I772181);
not I_45275 (I772212,I772142);
nor I_45276 (I772229,I772212,I771952);
DFFARX1 I_45277 (I772229,I2507,I771782,I771771,);
nor I_45278 (I772260,I251786,I251792);
or I_45279 (I771762,I772009,I772260);
nor I_45280 (I771753,I772142,I772260);
or I_45281 (I771756,I771876,I772260);
DFFARX1 I_45282 (I772260,I2507,I771782,I771774,);
not I_45283 (I772360,I2514);
DFFARX1 I_45284 (I879732,I2507,I772360,I772386,);
not I_45285 (I772394,I772386);
nand I_45286 (I772411,I879720,I879738);
and I_45287 (I772428,I772411,I879735);
DFFARX1 I_45288 (I772428,I2507,I772360,I772454,);
not I_45289 (I772462,I879726);
DFFARX1 I_45290 (I879723,I2507,I772360,I772488,);
not I_45291 (I772496,I772488);
nor I_45292 (I772513,I772496,I772394);
and I_45293 (I772530,I772513,I879726);
nor I_45294 (I772547,I772496,I772462);
nor I_45295 (I772343,I772454,I772547);
DFFARX1 I_45296 (I879717,I2507,I772360,I772587,);
nor I_45297 (I772595,I772587,I772454);
not I_45298 (I772612,I772595);
not I_45299 (I772629,I772587);
nor I_45300 (I772646,I772629,I772530);
DFFARX1 I_45301 (I772646,I2507,I772360,I772346,);
nand I_45302 (I772677,I879717,I879720);
and I_45303 (I772694,I772677,I879723);
DFFARX1 I_45304 (I772694,I2507,I772360,I772720,);
nor I_45305 (I772728,I772720,I772587);
DFFARX1 I_45306 (I772728,I2507,I772360,I772328,);
nand I_45307 (I772759,I772720,I772629);
nand I_45308 (I772337,I772612,I772759);
not I_45309 (I772790,I772720);
nor I_45310 (I772807,I772790,I772530);
DFFARX1 I_45311 (I772807,I2507,I772360,I772349,);
nor I_45312 (I772838,I879729,I879720);
or I_45313 (I772340,I772587,I772838);
nor I_45314 (I772331,I772720,I772838);
or I_45315 (I772334,I772454,I772838);
DFFARX1 I_45316 (I772838,I2507,I772360,I772352,);
not I_45317 (I772938,I2514);
DFFARX1 I_45318 (I813330,I2507,I772938,I772964,);
not I_45319 (I772972,I772964);
nand I_45320 (I772989,I813318,I813336);
and I_45321 (I773006,I772989,I813333);
DFFARX1 I_45322 (I773006,I2507,I772938,I773032,);
not I_45323 (I773040,I813324);
DFFARX1 I_45324 (I813321,I2507,I772938,I773066,);
not I_45325 (I773074,I773066);
nor I_45326 (I773091,I773074,I772972);
and I_45327 (I773108,I773091,I813324);
nor I_45328 (I773125,I773074,I773040);
nor I_45329 (I772921,I773032,I773125);
DFFARX1 I_45330 (I813315,I2507,I772938,I773165,);
nor I_45331 (I773173,I773165,I773032);
not I_45332 (I773190,I773173);
not I_45333 (I773207,I773165);
nor I_45334 (I773224,I773207,I773108);
DFFARX1 I_45335 (I773224,I2507,I772938,I772924,);
nand I_45336 (I773255,I813315,I813318);
and I_45337 (I773272,I773255,I813321);
DFFARX1 I_45338 (I773272,I2507,I772938,I773298,);
nor I_45339 (I773306,I773298,I773165);
DFFARX1 I_45340 (I773306,I2507,I772938,I772906,);
nand I_45341 (I773337,I773298,I773207);
nand I_45342 (I772915,I773190,I773337);
not I_45343 (I773368,I773298);
nor I_45344 (I773385,I773368,I773108);
DFFARX1 I_45345 (I773385,I2507,I772938,I772927,);
nor I_45346 (I773416,I813327,I813318);
or I_45347 (I772918,I773165,I773416);
nor I_45348 (I772909,I773298,I773416);
or I_45349 (I772912,I773032,I773416);
DFFARX1 I_45350 (I773416,I2507,I772938,I772930,);
not I_45351 (I773516,I2514);
DFFARX1 I_45352 (I1288856,I2507,I773516,I773542,);
not I_45353 (I773550,I773542);
nand I_45354 (I773567,I1288880,I1288862);
and I_45355 (I773584,I773567,I1288868);
DFFARX1 I_45356 (I773584,I2507,I773516,I773610,);
not I_45357 (I773618,I1288874);
DFFARX1 I_45358 (I1288859,I2507,I773516,I773644,);
not I_45359 (I773652,I773644);
nor I_45360 (I773669,I773652,I773550);
and I_45361 (I773686,I773669,I1288874);
nor I_45362 (I773703,I773652,I773618);
nor I_45363 (I773499,I773610,I773703);
DFFARX1 I_45364 (I1288871,I2507,I773516,I773743,);
nor I_45365 (I773751,I773743,I773610);
not I_45366 (I773768,I773751);
not I_45367 (I773785,I773743);
nor I_45368 (I773802,I773785,I773686);
DFFARX1 I_45369 (I773802,I2507,I773516,I773502,);
nand I_45370 (I773833,I1288877,I1288865);
and I_45371 (I773850,I773833,I1288859);
DFFARX1 I_45372 (I773850,I2507,I773516,I773876,);
nor I_45373 (I773884,I773876,I773743);
DFFARX1 I_45374 (I773884,I2507,I773516,I773484,);
nand I_45375 (I773915,I773876,I773785);
nand I_45376 (I773493,I773768,I773915);
not I_45377 (I773946,I773876);
nor I_45378 (I773963,I773946,I773686);
DFFARX1 I_45379 (I773963,I2507,I773516,I773505,);
nor I_45380 (I773994,I1288856,I1288865);
or I_45381 (I773496,I773743,I773994);
nor I_45382 (I773487,I773876,I773994);
or I_45383 (I773490,I773610,I773994);
DFFARX1 I_45384 (I773994,I2507,I773516,I773508,);
not I_45385 (I774094,I2514);
DFFARX1 I_45386 (I219845,I2507,I774094,I774120,);
not I_45387 (I774128,I774120);
nand I_45388 (I774145,I219848,I219869);
and I_45389 (I774162,I774145,I219857);
DFFARX1 I_45390 (I774162,I2507,I774094,I774188,);
not I_45391 (I774196,I219854);
DFFARX1 I_45392 (I219845,I2507,I774094,I774222,);
not I_45393 (I774230,I774222);
nor I_45394 (I774247,I774230,I774128);
and I_45395 (I774264,I774247,I219854);
nor I_45396 (I774281,I774230,I774196);
nor I_45397 (I774077,I774188,I774281);
DFFARX1 I_45398 (I219863,I2507,I774094,I774321,);
nor I_45399 (I774329,I774321,I774188);
not I_45400 (I774346,I774329);
not I_45401 (I774363,I774321);
nor I_45402 (I774380,I774363,I774264);
DFFARX1 I_45403 (I774380,I2507,I774094,I774080,);
nand I_45404 (I774411,I219848,I219851);
and I_45405 (I774428,I774411,I219860);
DFFARX1 I_45406 (I774428,I2507,I774094,I774454,);
nor I_45407 (I774462,I774454,I774321);
DFFARX1 I_45408 (I774462,I2507,I774094,I774062,);
nand I_45409 (I774493,I774454,I774363);
nand I_45410 (I774071,I774346,I774493);
not I_45411 (I774524,I774454);
nor I_45412 (I774541,I774524,I774264);
DFFARX1 I_45413 (I774541,I2507,I774094,I774083,);
nor I_45414 (I774572,I219866,I219851);
or I_45415 (I774074,I774321,I774572);
nor I_45416 (I774065,I774454,I774572);
or I_45417 (I774068,I774188,I774572);
DFFARX1 I_45418 (I774572,I2507,I774094,I774086,);
not I_45419 (I774672,I2514);
DFFARX1 I_45420 (I1037636,I2507,I774672,I774698,);
not I_45421 (I774706,I774698);
nand I_45422 (I774723,I1037633,I1037651);
and I_45423 (I774740,I774723,I1037648);
DFFARX1 I_45424 (I774740,I2507,I774672,I774766,);
not I_45425 (I774774,I1037630);
DFFARX1 I_45426 (I1037633,I2507,I774672,I774800,);
not I_45427 (I774808,I774800);
nor I_45428 (I774825,I774808,I774706);
and I_45429 (I774842,I774825,I1037630);
nor I_45430 (I774859,I774808,I774774);
nor I_45431 (I774655,I774766,I774859);
DFFARX1 I_45432 (I1037642,I2507,I774672,I774899,);
nor I_45433 (I774907,I774899,I774766);
not I_45434 (I774924,I774907);
not I_45435 (I774941,I774899);
nor I_45436 (I774958,I774941,I774842);
DFFARX1 I_45437 (I774958,I2507,I774672,I774658,);
nand I_45438 (I774989,I1037645,I1037630);
and I_45439 (I775006,I774989,I1037636);
DFFARX1 I_45440 (I775006,I2507,I774672,I775032,);
nor I_45441 (I775040,I775032,I774899);
DFFARX1 I_45442 (I775040,I2507,I774672,I774640,);
nand I_45443 (I775071,I775032,I774941);
nand I_45444 (I774649,I774924,I775071);
not I_45445 (I775102,I775032);
nor I_45446 (I775119,I775102,I774842);
DFFARX1 I_45447 (I775119,I2507,I774672,I774661,);
nor I_45448 (I775150,I1037639,I1037630);
or I_45449 (I774652,I774899,I775150);
nor I_45450 (I774643,I775032,I775150);
or I_45451 (I774646,I774766,I775150);
DFFARX1 I_45452 (I775150,I2507,I774672,I774664,);
not I_45453 (I775250,I2514);
DFFARX1 I_45454 (I72781,I2507,I775250,I775276,);
not I_45455 (I775284,I775276);
nand I_45456 (I775301,I72790,I72799);
and I_45457 (I775318,I775301,I72778);
DFFARX1 I_45458 (I775318,I2507,I775250,I775344,);
not I_45459 (I775352,I72781);
DFFARX1 I_45460 (I72796,I2507,I775250,I775378,);
not I_45461 (I775386,I775378);
nor I_45462 (I775403,I775386,I775284);
and I_45463 (I775420,I775403,I72781);
nor I_45464 (I775437,I775386,I775352);
nor I_45465 (I775233,I775344,I775437);
DFFARX1 I_45466 (I72787,I2507,I775250,I775477,);
nor I_45467 (I775485,I775477,I775344);
not I_45468 (I775502,I775485);
not I_45469 (I775519,I775477);
nor I_45470 (I775536,I775519,I775420);
DFFARX1 I_45471 (I775536,I2507,I775250,I775236,);
nand I_45472 (I775567,I72802,I72778);
and I_45473 (I775584,I775567,I72784);
DFFARX1 I_45474 (I775584,I2507,I775250,I775610,);
nor I_45475 (I775618,I775610,I775477);
DFFARX1 I_45476 (I775618,I2507,I775250,I775218,);
nand I_45477 (I775649,I775610,I775519);
nand I_45478 (I775227,I775502,I775649);
not I_45479 (I775680,I775610);
nor I_45480 (I775697,I775680,I775420);
DFFARX1 I_45481 (I775697,I2507,I775250,I775239,);
nor I_45482 (I775728,I72793,I72778);
or I_45483 (I775230,I775477,I775728);
nor I_45484 (I775221,I775610,I775728);
or I_45485 (I775224,I775344,I775728);
DFFARX1 I_45486 (I775728,I2507,I775250,I775242,);
not I_45487 (I775828,I2514);
DFFARX1 I_45488 (I1014635,I2507,I775828,I775854,);
not I_45489 (I775862,I775854);
nand I_45490 (I775879,I1014632,I1014650);
and I_45491 (I775896,I775879,I1014647);
DFFARX1 I_45492 (I775896,I2507,I775828,I775922,);
not I_45493 (I775930,I1014629);
DFFARX1 I_45494 (I1014632,I2507,I775828,I775956,);
not I_45495 (I775964,I775956);
nor I_45496 (I775981,I775964,I775862);
and I_45497 (I775998,I775981,I1014629);
nor I_45498 (I776015,I775964,I775930);
nor I_45499 (I775811,I775922,I776015);
DFFARX1 I_45500 (I1014641,I2507,I775828,I776055,);
nor I_45501 (I776063,I776055,I775922);
not I_45502 (I776080,I776063);
not I_45503 (I776097,I776055);
nor I_45504 (I776114,I776097,I775998);
DFFARX1 I_45505 (I776114,I2507,I775828,I775814,);
nand I_45506 (I776145,I1014644,I1014629);
and I_45507 (I776162,I776145,I1014635);
DFFARX1 I_45508 (I776162,I2507,I775828,I776188,);
nor I_45509 (I776196,I776188,I776055);
DFFARX1 I_45510 (I776196,I2507,I775828,I775796,);
nand I_45511 (I776227,I776188,I776097);
nand I_45512 (I775805,I776080,I776227);
not I_45513 (I776258,I776188);
nor I_45514 (I776275,I776258,I775998);
DFFARX1 I_45515 (I776275,I2507,I775828,I775817,);
nor I_45516 (I776306,I1014638,I1014629);
or I_45517 (I775808,I776055,I776306);
nor I_45518 (I775799,I776188,I776306);
or I_45519 (I775802,I775922,I776306);
DFFARX1 I_45520 (I776306,I2507,I775828,I775820,);
not I_45521 (I776406,I2514);
DFFARX1 I_45522 (I396824,I2507,I776406,I776432,);
not I_45523 (I776440,I776432);
nand I_45524 (I776457,I396815,I396833);
and I_45525 (I776474,I776457,I396836);
DFFARX1 I_45526 (I776474,I2507,I776406,I776500,);
not I_45527 (I776508,I396830);
DFFARX1 I_45528 (I396818,I2507,I776406,I776534,);
not I_45529 (I776542,I776534);
nor I_45530 (I776559,I776542,I776440);
and I_45531 (I776576,I776559,I396830);
nor I_45532 (I776593,I776542,I776508);
nor I_45533 (I776389,I776500,I776593);
DFFARX1 I_45534 (I396827,I2507,I776406,I776633,);
nor I_45535 (I776641,I776633,I776500);
not I_45536 (I776658,I776641);
not I_45537 (I776675,I776633);
nor I_45538 (I776692,I776675,I776576);
DFFARX1 I_45539 (I776692,I2507,I776406,I776392,);
nand I_45540 (I776723,I396842,I396839);
and I_45541 (I776740,I776723,I396821);
DFFARX1 I_45542 (I776740,I2507,I776406,I776766,);
nor I_45543 (I776774,I776766,I776633);
DFFARX1 I_45544 (I776774,I2507,I776406,I776374,);
nand I_45545 (I776805,I776766,I776675);
nand I_45546 (I776383,I776658,I776805);
not I_45547 (I776836,I776766);
nor I_45548 (I776853,I776836,I776576);
DFFARX1 I_45549 (I776853,I2507,I776406,I776395,);
nor I_45550 (I776884,I396815,I396839);
or I_45551 (I776386,I776633,I776884);
nor I_45552 (I776377,I776766,I776884);
or I_45553 (I776380,I776500,I776884);
DFFARX1 I_45554 (I776884,I2507,I776406,I776398,);
not I_45555 (I776981,I2514);
DFFARX1 I_45556 (I1042127,I2507,I776981,I777007,);
not I_45557 (I777015,I777007);
nand I_45558 (I777032,I1042136,I1042124);
and I_45559 (I777049,I777032,I1042121);
DFFARX1 I_45560 (I777049,I2507,I776981,I777075,);
DFFARX1 I_45561 (I777075,I2507,I776981,I776970,);
DFFARX1 I_45562 (I1042121,I2507,I776981,I777106,);
nand I_45563 (I777114,I777106,I1042118);
not I_45564 (I777131,I777114);
DFFARX1 I_45565 (I777131,I2507,I776981,I777157,);
not I_45566 (I777165,I777157);
nor I_45567 (I776973,I777015,I777165);
DFFARX1 I_45568 (I1042124,I2507,I776981,I777205,);
nor I_45569 (I776964,I777205,I777075);
nor I_45570 (I776955,I777205,I777131);
nand I_45571 (I777241,I1042139,I1042130);
and I_45572 (I777258,I777241,I1042133);
DFFARX1 I_45573 (I777258,I2507,I776981,I777284,);
not I_45574 (I777292,I777284);
nand I_45575 (I777309,I777292,I777205);
nand I_45576 (I776958,I777292,I777114);
nor I_45577 (I777340,I1042118,I1042130);
and I_45578 (I777357,I777205,I777340);
nor I_45579 (I777374,I777292,I777357);
DFFARX1 I_45580 (I777374,I2507,I776981,I776967,);
nor I_45581 (I777405,I777007,I777340);
DFFARX1 I_45582 (I777405,I2507,I776981,I776952,);
nor I_45583 (I777436,I777284,I777340);
not I_45584 (I777453,I777436);
nand I_45585 (I776961,I777453,I777309);
not I_45586 (I777508,I2514);
DFFARX1 I_45587 (I71748,I2507,I777508,I777534,);
not I_45588 (I777542,I777534);
nand I_45589 (I777559,I71724,I71733);
and I_45590 (I777576,I777559,I71727);
DFFARX1 I_45591 (I777576,I2507,I777508,I777602,);
DFFARX1 I_45592 (I777602,I2507,I777508,I777497,);
DFFARX1 I_45593 (I71745,I2507,I777508,I777633,);
nand I_45594 (I777641,I777633,I71736);
not I_45595 (I777658,I777641);
DFFARX1 I_45596 (I777658,I2507,I777508,I777684,);
not I_45597 (I777692,I777684);
nor I_45598 (I777500,I777542,I777692);
DFFARX1 I_45599 (I71730,I2507,I777508,I777732,);
nor I_45600 (I777491,I777732,I777602);
nor I_45601 (I777482,I777732,I777658);
nand I_45602 (I777768,I71742,I71739);
and I_45603 (I777785,I777768,I71727);
DFFARX1 I_45604 (I777785,I2507,I777508,I777811,);
not I_45605 (I777819,I777811);
nand I_45606 (I777836,I777819,I777732);
nand I_45607 (I777485,I777819,I777641);
nor I_45608 (I777867,I71724,I71739);
and I_45609 (I777884,I777732,I777867);
nor I_45610 (I777901,I777819,I777884);
DFFARX1 I_45611 (I777901,I2507,I777508,I777494,);
nor I_45612 (I777932,I777534,I777867);
DFFARX1 I_45613 (I777932,I2507,I777508,I777479,);
nor I_45614 (I777963,I777811,I777867);
not I_45615 (I777980,I777963);
nand I_45616 (I777488,I777980,I777836);
not I_45617 (I778035,I2514);
DFFARX1 I_45618 (I522655,I2507,I778035,I778061,);
not I_45619 (I778069,I778061);
nand I_45620 (I778086,I522673,I522664);
and I_45621 (I778103,I778086,I522667);
DFFARX1 I_45622 (I778103,I2507,I778035,I778129,);
DFFARX1 I_45623 (I778129,I2507,I778035,I778024,);
DFFARX1 I_45624 (I522661,I2507,I778035,I778160,);
nand I_45625 (I778168,I778160,I522652);
not I_45626 (I778185,I778168);
DFFARX1 I_45627 (I778185,I2507,I778035,I778211,);
not I_45628 (I778219,I778211);
nor I_45629 (I778027,I778069,I778219);
DFFARX1 I_45630 (I522658,I2507,I778035,I778259,);
nor I_45631 (I778018,I778259,I778129);
nor I_45632 (I778009,I778259,I778185);
nand I_45633 (I778295,I522652,I522649);
and I_45634 (I778312,I778295,I522670);
DFFARX1 I_45635 (I778312,I2507,I778035,I778338,);
not I_45636 (I778346,I778338);
nand I_45637 (I778363,I778346,I778259);
nand I_45638 (I778012,I778346,I778168);
nor I_45639 (I778394,I522649,I522649);
and I_45640 (I778411,I778259,I778394);
nor I_45641 (I778428,I778346,I778411);
DFFARX1 I_45642 (I778428,I2507,I778035,I778021,);
nor I_45643 (I778459,I778061,I778394);
DFFARX1 I_45644 (I778459,I2507,I778035,I778006,);
nor I_45645 (I778490,I778338,I778394);
not I_45646 (I778507,I778490);
nand I_45647 (I778015,I778507,I778363);
not I_45648 (I778562,I2514);
DFFARX1 I_45649 (I321344,I2507,I778562,I778588,);
not I_45650 (I778596,I778588);
nand I_45651 (I778613,I321335,I321335);
and I_45652 (I778630,I778613,I321353);
DFFARX1 I_45653 (I778630,I2507,I778562,I778656,);
DFFARX1 I_45654 (I778656,I2507,I778562,I778551,);
DFFARX1 I_45655 (I321356,I2507,I778562,I778687,);
nand I_45656 (I778695,I778687,I321338);
not I_45657 (I778712,I778695);
DFFARX1 I_45658 (I778712,I2507,I778562,I778738,);
not I_45659 (I778746,I778738);
nor I_45660 (I778554,I778596,I778746);
DFFARX1 I_45661 (I321350,I2507,I778562,I778786,);
nor I_45662 (I778545,I778786,I778656);
nor I_45663 (I778536,I778786,I778712);
nand I_45664 (I778822,I321362,I321341);
and I_45665 (I778839,I778822,I321347);
DFFARX1 I_45666 (I778839,I2507,I778562,I778865,);
not I_45667 (I778873,I778865);
nand I_45668 (I778890,I778873,I778786);
nand I_45669 (I778539,I778873,I778695);
nor I_45670 (I778921,I321359,I321341);
and I_45671 (I778938,I778786,I778921);
nor I_45672 (I778955,I778873,I778938);
DFFARX1 I_45673 (I778955,I2507,I778562,I778548,);
nor I_45674 (I778986,I778588,I778921);
DFFARX1 I_45675 (I778986,I2507,I778562,I778533,);
nor I_45676 (I779017,I778865,I778921);
not I_45677 (I779034,I779017);
nand I_45678 (I778542,I779034,I778890);
not I_45679 (I779089,I2514);
DFFARX1 I_45680 (I170466,I2507,I779089,I779115,);
not I_45681 (I779123,I779115);
nand I_45682 (I779140,I170463,I170481);
and I_45683 (I779157,I779140,I170472);
DFFARX1 I_45684 (I779157,I2507,I779089,I779183,);
DFFARX1 I_45685 (I779183,I2507,I779089,I779078,);
DFFARX1 I_45686 (I170478,I2507,I779089,I779214,);
nand I_45687 (I779222,I779214,I170475);
not I_45688 (I779239,I779222);
DFFARX1 I_45689 (I779239,I2507,I779089,I779265,);
not I_45690 (I779273,I779265);
nor I_45691 (I779081,I779123,I779273);
DFFARX1 I_45692 (I170469,I2507,I779089,I779313,);
nor I_45693 (I779072,I779313,I779183);
nor I_45694 (I779063,I779313,I779239);
nand I_45695 (I779349,I170460,I170484);
and I_45696 (I779366,I779349,I170463);
DFFARX1 I_45697 (I779366,I2507,I779089,I779392,);
not I_45698 (I779400,I779392);
nand I_45699 (I779417,I779400,I779313);
nand I_45700 (I779066,I779400,I779222);
nor I_45701 (I779448,I170460,I170484);
and I_45702 (I779465,I779313,I779448);
nor I_45703 (I779482,I779400,I779465);
DFFARX1 I_45704 (I779482,I2507,I779089,I779075,);
nor I_45705 (I779513,I779115,I779448);
DFFARX1 I_45706 (I779513,I2507,I779089,I779060,);
nor I_45707 (I779544,I779392,I779448);
not I_45708 (I779561,I779544);
nand I_45709 (I779069,I779561,I779417);
not I_45710 (I779616,I2514);
DFFARX1 I_45711 (I115489,I2507,I779616,I779642,);
not I_45712 (I779650,I779642);
nand I_45713 (I779667,I115465,I115474);
and I_45714 (I779684,I779667,I115468);
DFFARX1 I_45715 (I779684,I2507,I779616,I779710,);
DFFARX1 I_45716 (I779710,I2507,I779616,I779605,);
DFFARX1 I_45717 (I115486,I2507,I779616,I779741,);
nand I_45718 (I779749,I779741,I115477);
not I_45719 (I779766,I779749);
DFFARX1 I_45720 (I779766,I2507,I779616,I779792,);
not I_45721 (I779800,I779792);
nor I_45722 (I779608,I779650,I779800);
DFFARX1 I_45723 (I115471,I2507,I779616,I779840,);
nor I_45724 (I779599,I779840,I779710);
nor I_45725 (I779590,I779840,I779766);
nand I_45726 (I779876,I115483,I115480);
and I_45727 (I779893,I779876,I115468);
DFFARX1 I_45728 (I779893,I2507,I779616,I779919,);
not I_45729 (I779927,I779919);
nand I_45730 (I779944,I779927,I779840);
nand I_45731 (I779593,I779927,I779749);
nor I_45732 (I779975,I115465,I115480);
and I_45733 (I779992,I779840,I779975);
nor I_45734 (I780009,I779927,I779992);
DFFARX1 I_45735 (I780009,I2507,I779616,I779602,);
nor I_45736 (I780040,I779642,I779975);
DFFARX1 I_45737 (I780040,I2507,I779616,I779587,);
nor I_45738 (I780071,I779919,I779975);
not I_45739 (I780088,I780071);
nand I_45740 (I779596,I780088,I779944);
not I_45741 (I780143,I2514);
DFFARX1 I_45742 (I1306517,I2507,I780143,I780169,);
not I_45743 (I780177,I780169);
nand I_45744 (I780194,I1306514,I1306523);
and I_45745 (I780211,I780194,I1306502);
DFFARX1 I_45746 (I780211,I2507,I780143,I780237,);
DFFARX1 I_45747 (I780237,I2507,I780143,I780132,);
DFFARX1 I_45748 (I1306505,I2507,I780143,I780268,);
nand I_45749 (I780276,I780268,I1306520);
not I_45750 (I780293,I780276);
DFFARX1 I_45751 (I780293,I2507,I780143,I780319,);
not I_45752 (I780327,I780319);
nor I_45753 (I780135,I780177,I780327);
DFFARX1 I_45754 (I1306526,I2507,I780143,I780367,);
nor I_45755 (I780126,I780367,I780237);
nor I_45756 (I780117,I780367,I780293);
nand I_45757 (I780403,I1306508,I1306529);
and I_45758 (I780420,I780403,I1306511);
DFFARX1 I_45759 (I780420,I2507,I780143,I780446,);
not I_45760 (I780454,I780446);
nand I_45761 (I780471,I780454,I780367);
nand I_45762 (I780120,I780454,I780276);
nor I_45763 (I780502,I1306502,I1306529);
and I_45764 (I780519,I780367,I780502);
nor I_45765 (I780536,I780454,I780519);
DFFARX1 I_45766 (I780536,I2507,I780143,I780129,);
nor I_45767 (I780567,I780169,I780502);
DFFARX1 I_45768 (I780567,I2507,I780143,I780114,);
nor I_45769 (I780598,I780446,I780502);
not I_45770 (I780615,I780598);
nand I_45771 (I780123,I780615,I780471);
not I_45772 (I780670,I2514);
DFFARX1 I_45773 (I128137,I2507,I780670,I780696,);
not I_45774 (I780704,I780696);
nand I_45775 (I780721,I128113,I128122);
and I_45776 (I780738,I780721,I128116);
DFFARX1 I_45777 (I780738,I2507,I780670,I780764,);
DFFARX1 I_45778 (I780764,I2507,I780670,I780659,);
DFFARX1 I_45779 (I128134,I2507,I780670,I780795,);
nand I_45780 (I780803,I780795,I128125);
not I_45781 (I780820,I780803);
DFFARX1 I_45782 (I780820,I2507,I780670,I780846,);
not I_45783 (I780854,I780846);
nor I_45784 (I780662,I780704,I780854);
DFFARX1 I_45785 (I128119,I2507,I780670,I780894,);
nor I_45786 (I780653,I780894,I780764);
nor I_45787 (I780644,I780894,I780820);
nand I_45788 (I780930,I128131,I128128);
and I_45789 (I780947,I780930,I128116);
DFFARX1 I_45790 (I780947,I2507,I780670,I780973,);
not I_45791 (I780981,I780973);
nand I_45792 (I780998,I780981,I780894);
nand I_45793 (I780647,I780981,I780803);
nor I_45794 (I781029,I128113,I128128);
and I_45795 (I781046,I780894,I781029);
nor I_45796 (I781063,I780981,I781046);
DFFARX1 I_45797 (I781063,I2507,I780670,I780656,);
nor I_45798 (I781094,I780696,I781029);
DFFARX1 I_45799 (I781094,I2507,I780670,I780641,);
nor I_45800 (I781125,I780973,I781029);
not I_45801 (I781142,I781125);
nand I_45802 (I780650,I781142,I780998);
not I_45803 (I781197,I2514);
DFFARX1 I_45804 (I1391007,I2507,I781197,I781223,);
not I_45805 (I781231,I781223);
nand I_45806 (I781248,I1391004,I1391013);
and I_45807 (I781265,I781248,I1390992);
DFFARX1 I_45808 (I781265,I2507,I781197,I781291,);
DFFARX1 I_45809 (I781291,I2507,I781197,I781186,);
DFFARX1 I_45810 (I1390995,I2507,I781197,I781322,);
nand I_45811 (I781330,I781322,I1391010);
not I_45812 (I781347,I781330);
DFFARX1 I_45813 (I781347,I2507,I781197,I781373,);
not I_45814 (I781381,I781373);
nor I_45815 (I781189,I781231,I781381);
DFFARX1 I_45816 (I1391016,I2507,I781197,I781421,);
nor I_45817 (I781180,I781421,I781291);
nor I_45818 (I781171,I781421,I781347);
nand I_45819 (I781457,I1390998,I1391019);
and I_45820 (I781474,I781457,I1391001);
DFFARX1 I_45821 (I781474,I2507,I781197,I781500,);
not I_45822 (I781508,I781500);
nand I_45823 (I781525,I781508,I781421);
nand I_45824 (I781174,I781508,I781330);
nor I_45825 (I781556,I1390992,I1391019);
and I_45826 (I781573,I781421,I781556);
nor I_45827 (I781590,I781508,I781573);
DFFARX1 I_45828 (I781590,I2507,I781197,I781183,);
nor I_45829 (I781621,I781223,I781556);
DFFARX1 I_45830 (I781621,I2507,I781197,I781168,);
nor I_45831 (I781652,I781500,I781556);
not I_45832 (I781669,I781652);
nand I_45833 (I781177,I781669,I781525);
not I_45834 (I781724,I2514);
DFFARX1 I_45835 (I1216142,I2507,I781724,I781750,);
not I_45836 (I781758,I781750);
nand I_45837 (I781775,I1216148,I1216130);
and I_45838 (I781792,I781775,I1216139);
DFFARX1 I_45839 (I781792,I2507,I781724,I781818,);
DFFARX1 I_45840 (I781818,I2507,I781724,I781713,);
DFFARX1 I_45841 (I1216145,I2507,I781724,I781849,);
nand I_45842 (I781857,I781849,I1216133);
not I_45843 (I781874,I781857);
DFFARX1 I_45844 (I781874,I2507,I781724,I781900,);
not I_45845 (I781908,I781900);
nor I_45846 (I781716,I781758,I781908);
DFFARX1 I_45847 (I1216151,I2507,I781724,I781948,);
nor I_45848 (I781707,I781948,I781818);
nor I_45849 (I781698,I781948,I781874);
nand I_45850 (I781984,I1216130,I1216136);
and I_45851 (I782001,I781984,I1216154);
DFFARX1 I_45852 (I782001,I2507,I781724,I782027,);
not I_45853 (I782035,I782027);
nand I_45854 (I782052,I782035,I781948);
nand I_45855 (I781701,I782035,I781857);
nor I_45856 (I782083,I1216133,I1216136);
and I_45857 (I782100,I781948,I782083);
nor I_45858 (I782117,I782035,I782100);
DFFARX1 I_45859 (I782117,I2507,I781724,I781710,);
nor I_45860 (I782148,I781750,I782083);
DFFARX1 I_45861 (I782148,I2507,I781724,I781695,);
nor I_45862 (I782179,I782027,I782083);
not I_45863 (I782196,I782179);
nand I_45864 (I781704,I782196,I782052);
not I_45865 (I782251,I2514);
DFFARX1 I_45866 (I950236,I2507,I782251,I782277,);
not I_45867 (I782285,I782277);
nand I_45868 (I782302,I950251,I950233);
and I_45869 (I782319,I782302,I950233);
DFFARX1 I_45870 (I782319,I2507,I782251,I782345,);
DFFARX1 I_45871 (I782345,I2507,I782251,I782240,);
DFFARX1 I_45872 (I950242,I2507,I782251,I782376,);
nand I_45873 (I782384,I782376,I950260);
not I_45874 (I782401,I782384);
DFFARX1 I_45875 (I782401,I2507,I782251,I782427,);
not I_45876 (I782435,I782427);
nor I_45877 (I782243,I782285,I782435);
DFFARX1 I_45878 (I950257,I2507,I782251,I782475,);
nor I_45879 (I782234,I782475,I782345);
nor I_45880 (I782225,I782475,I782401);
nand I_45881 (I782511,I950254,I950245);
and I_45882 (I782528,I782511,I950239);
DFFARX1 I_45883 (I782528,I2507,I782251,I782554,);
not I_45884 (I782562,I782554);
nand I_45885 (I782579,I782562,I782475);
nand I_45886 (I782228,I782562,I782384);
nor I_45887 (I782610,I950248,I950245);
and I_45888 (I782627,I782475,I782610);
nor I_45889 (I782644,I782562,I782627);
DFFARX1 I_45890 (I782644,I2507,I782251,I782237,);
nor I_45891 (I782675,I782277,I782610);
DFFARX1 I_45892 (I782675,I2507,I782251,I782222,);
nor I_45893 (I782706,I782554,I782610);
not I_45894 (I782723,I782706);
nand I_45895 (I782231,I782723,I782579);
not I_45896 (I782778,I2514);
DFFARX1 I_45897 (I767126,I2507,I782778,I782804,);
not I_45898 (I782812,I782804);
nand I_45899 (I782829,I767129,I767126);
and I_45900 (I782846,I782829,I767138);
DFFARX1 I_45901 (I782846,I2507,I782778,I782872,);
DFFARX1 I_45902 (I782872,I2507,I782778,I782767,);
DFFARX1 I_45903 (I767135,I2507,I782778,I782903,);
nand I_45904 (I782911,I782903,I767141);
not I_45905 (I782928,I782911);
DFFARX1 I_45906 (I782928,I2507,I782778,I782954,);
not I_45907 (I782962,I782954);
nor I_45908 (I782770,I782812,I782962);
DFFARX1 I_45909 (I767150,I2507,I782778,I783002,);
nor I_45910 (I782761,I783002,I782872);
nor I_45911 (I782752,I783002,I782928);
nand I_45912 (I783038,I767144,I767132);
and I_45913 (I783055,I783038,I767129);
DFFARX1 I_45914 (I783055,I2507,I782778,I783081,);
not I_45915 (I783089,I783081);
nand I_45916 (I783106,I783089,I783002);
nand I_45917 (I782755,I783089,I782911);
nor I_45918 (I783137,I767147,I767132);
and I_45919 (I783154,I783002,I783137);
nor I_45920 (I783171,I783089,I783154);
DFFARX1 I_45921 (I783171,I2507,I782778,I782764,);
nor I_45922 (I783202,I782804,I783137);
DFFARX1 I_45923 (I783202,I2507,I782778,I782749,);
nor I_45924 (I783233,I783081,I783137);
not I_45925 (I783250,I783233);
nand I_45926 (I782758,I783250,I783106);
not I_45927 (I783305,I2514);
DFFARX1 I_45928 (I345059,I2507,I783305,I783331,);
not I_45929 (I783339,I783331);
nand I_45930 (I783356,I345050,I345050);
and I_45931 (I783373,I783356,I345068);
DFFARX1 I_45932 (I783373,I2507,I783305,I783399,);
DFFARX1 I_45933 (I783399,I2507,I783305,I783294,);
DFFARX1 I_45934 (I345071,I2507,I783305,I783430,);
nand I_45935 (I783438,I783430,I345053);
not I_45936 (I783455,I783438);
DFFARX1 I_45937 (I783455,I2507,I783305,I783481,);
not I_45938 (I783489,I783481);
nor I_45939 (I783297,I783339,I783489);
DFFARX1 I_45940 (I345065,I2507,I783305,I783529,);
nor I_45941 (I783288,I783529,I783399);
nor I_45942 (I783279,I783529,I783455);
nand I_45943 (I783565,I345077,I345056);
and I_45944 (I783582,I783565,I345062);
DFFARX1 I_45945 (I783582,I2507,I783305,I783608,);
not I_45946 (I783616,I783608);
nand I_45947 (I783633,I783616,I783529);
nand I_45948 (I783282,I783616,I783438);
nor I_45949 (I783664,I345074,I345056);
and I_45950 (I783681,I783529,I783664);
nor I_45951 (I783698,I783616,I783681);
DFFARX1 I_45952 (I783698,I2507,I783305,I783291,);
nor I_45953 (I783729,I783331,I783664);
DFFARX1 I_45954 (I783729,I2507,I783305,I783276,);
nor I_45955 (I783760,I783608,I783664);
not I_45956 (I783777,I783760);
nand I_45957 (I783285,I783777,I783633);
not I_45958 (I783832,I2514);
DFFARX1 I_45959 (I1361257,I2507,I783832,I783858,);
not I_45960 (I783866,I783858);
nand I_45961 (I783883,I1361254,I1361263);
and I_45962 (I783900,I783883,I1361242);
DFFARX1 I_45963 (I783900,I2507,I783832,I783926,);
DFFARX1 I_45964 (I783926,I2507,I783832,I783821,);
DFFARX1 I_45965 (I1361245,I2507,I783832,I783957,);
nand I_45966 (I783965,I783957,I1361260);
not I_45967 (I783982,I783965);
DFFARX1 I_45968 (I783982,I2507,I783832,I784008,);
not I_45969 (I784016,I784008);
nor I_45970 (I783824,I783866,I784016);
DFFARX1 I_45971 (I1361266,I2507,I783832,I784056,);
nor I_45972 (I783815,I784056,I783926);
nor I_45973 (I783806,I784056,I783982);
nand I_45974 (I784092,I1361248,I1361269);
and I_45975 (I784109,I784092,I1361251);
DFFARX1 I_45976 (I784109,I2507,I783832,I784135,);
not I_45977 (I784143,I784135);
nand I_45978 (I784160,I784143,I784056);
nand I_45979 (I783809,I784143,I783965);
nor I_45980 (I784191,I1361242,I1361269);
and I_45981 (I784208,I784056,I784191);
nor I_45982 (I784225,I784143,I784208);
DFFARX1 I_45983 (I784225,I2507,I783832,I783818,);
nor I_45984 (I784256,I783858,I784191);
DFFARX1 I_45985 (I784256,I2507,I783832,I783803,);
nor I_45986 (I784287,I784135,I784191);
not I_45987 (I784304,I784287);
nand I_45988 (I783812,I784304,I784160);
not I_45989 (I784359,I2514);
DFFARX1 I_45990 (I1330317,I2507,I784359,I784385,);
not I_45991 (I784393,I784385);
nand I_45992 (I784410,I1330314,I1330323);
and I_45993 (I784427,I784410,I1330302);
DFFARX1 I_45994 (I784427,I2507,I784359,I784453,);
DFFARX1 I_45995 (I784453,I2507,I784359,I784348,);
DFFARX1 I_45996 (I1330305,I2507,I784359,I784484,);
nand I_45997 (I784492,I784484,I1330320);
not I_45998 (I784509,I784492);
DFFARX1 I_45999 (I784509,I2507,I784359,I784535,);
not I_46000 (I784543,I784535);
nor I_46001 (I784351,I784393,I784543);
DFFARX1 I_46002 (I1330326,I2507,I784359,I784583,);
nor I_46003 (I784342,I784583,I784453);
nor I_46004 (I784333,I784583,I784509);
nand I_46005 (I784619,I1330308,I1330329);
and I_46006 (I784636,I784619,I1330311);
DFFARX1 I_46007 (I784636,I2507,I784359,I784662,);
not I_46008 (I784670,I784662);
nand I_46009 (I784687,I784670,I784583);
nand I_46010 (I784336,I784670,I784492);
nor I_46011 (I784718,I1330302,I1330329);
and I_46012 (I784735,I784583,I784718);
nor I_46013 (I784752,I784670,I784735);
DFFARX1 I_46014 (I784752,I2507,I784359,I784345,);
nor I_46015 (I784783,I784385,I784718);
DFFARX1 I_46016 (I784783,I2507,I784359,I784330,);
nor I_46017 (I784814,I784662,I784718);
not I_46018 (I784831,I784814);
nand I_46019 (I784339,I784831,I784687);
not I_46020 (I784886,I2514);
DFFARX1 I_46021 (I1238990,I2507,I784886,I784912,);
not I_46022 (I784920,I784912);
nand I_46023 (I784937,I1238996,I1238978);
and I_46024 (I784954,I784937,I1238987);
DFFARX1 I_46025 (I784954,I2507,I784886,I784980,);
DFFARX1 I_46026 (I784980,I2507,I784886,I784875,);
DFFARX1 I_46027 (I1238993,I2507,I784886,I785011,);
nand I_46028 (I785019,I785011,I1238981);
not I_46029 (I785036,I785019);
DFFARX1 I_46030 (I785036,I2507,I784886,I785062,);
not I_46031 (I785070,I785062);
nor I_46032 (I784878,I784920,I785070);
DFFARX1 I_46033 (I1238999,I2507,I784886,I785110,);
nor I_46034 (I784869,I785110,I784980);
nor I_46035 (I784860,I785110,I785036);
nand I_46036 (I785146,I1238978,I1238984);
and I_46037 (I785163,I785146,I1239002);
DFFARX1 I_46038 (I785163,I2507,I784886,I785189,);
not I_46039 (I785197,I785189);
nand I_46040 (I785214,I785197,I785110);
nand I_46041 (I784863,I785197,I785019);
nor I_46042 (I785245,I1238981,I1238984);
and I_46043 (I785262,I785110,I785245);
nor I_46044 (I785279,I785197,I785262);
DFFARX1 I_46045 (I785279,I2507,I784886,I784872,);
nor I_46046 (I785310,I784912,I785245);
DFFARX1 I_46047 (I785310,I2507,I784886,I784857,);
nor I_46048 (I785341,I785189,I785245);
not I_46049 (I785358,I785341);
nand I_46050 (I784866,I785358,I785214);
not I_46051 (I785413,I2514);
DFFARX1 I_46052 (I327141,I2507,I785413,I785439,);
not I_46053 (I785447,I785439);
nand I_46054 (I785464,I327132,I327132);
and I_46055 (I785481,I785464,I327150);
DFFARX1 I_46056 (I785481,I2507,I785413,I785507,);
DFFARX1 I_46057 (I785507,I2507,I785413,I785402,);
DFFARX1 I_46058 (I327153,I2507,I785413,I785538,);
nand I_46059 (I785546,I785538,I327135);
not I_46060 (I785563,I785546);
DFFARX1 I_46061 (I785563,I2507,I785413,I785589,);
not I_46062 (I785597,I785589);
nor I_46063 (I785405,I785447,I785597);
DFFARX1 I_46064 (I327147,I2507,I785413,I785637,);
nor I_46065 (I785396,I785637,I785507);
nor I_46066 (I785387,I785637,I785563);
nand I_46067 (I785673,I327159,I327138);
and I_46068 (I785690,I785673,I327144);
DFFARX1 I_46069 (I785690,I2507,I785413,I785716,);
not I_46070 (I785724,I785716);
nand I_46071 (I785741,I785724,I785637);
nand I_46072 (I785390,I785724,I785546);
nor I_46073 (I785772,I327156,I327138);
and I_46074 (I785789,I785637,I785772);
nor I_46075 (I785806,I785724,I785789);
DFFARX1 I_46076 (I785806,I2507,I785413,I785399,);
nor I_46077 (I785837,I785439,I785772);
DFFARX1 I_46078 (I785837,I2507,I785413,I785384,);
nor I_46079 (I785868,I785716,I785772);
not I_46080 (I785885,I785868);
nand I_46081 (I785393,I785885,I785741);
not I_46082 (I785940,I2514);
DFFARX1 I_46083 (I122340,I2507,I785940,I785966,);
not I_46084 (I785974,I785966);
nand I_46085 (I785991,I122316,I122325);
and I_46086 (I786008,I785991,I122319);
DFFARX1 I_46087 (I786008,I2507,I785940,I786034,);
DFFARX1 I_46088 (I786034,I2507,I785940,I785929,);
DFFARX1 I_46089 (I122337,I2507,I785940,I786065,);
nand I_46090 (I786073,I786065,I122328);
not I_46091 (I786090,I786073);
DFFARX1 I_46092 (I786090,I2507,I785940,I786116,);
not I_46093 (I786124,I786116);
nor I_46094 (I785932,I785974,I786124);
DFFARX1 I_46095 (I122322,I2507,I785940,I786164,);
nor I_46096 (I785923,I786164,I786034);
nor I_46097 (I785914,I786164,I786090);
nand I_46098 (I786200,I122334,I122331);
and I_46099 (I786217,I786200,I122319);
DFFARX1 I_46100 (I786217,I2507,I785940,I786243,);
not I_46101 (I786251,I786243);
nand I_46102 (I786268,I786251,I786164);
nand I_46103 (I785917,I786251,I786073);
nor I_46104 (I786299,I122316,I122331);
and I_46105 (I786316,I786164,I786299);
nor I_46106 (I786333,I786251,I786316);
DFFARX1 I_46107 (I786333,I2507,I785940,I785926,);
nor I_46108 (I786364,I785966,I786299);
DFFARX1 I_46109 (I786364,I2507,I785940,I785911,);
nor I_46110 (I786395,I786243,I786299);
not I_46111 (I786412,I786395);
nand I_46112 (I785920,I786412,I786268);
not I_46113 (I786467,I2514);
DFFARX1 I_46114 (I311331,I2507,I786467,I786493,);
not I_46115 (I786501,I786493);
nand I_46116 (I786518,I311322,I311322);
and I_46117 (I786535,I786518,I311340);
DFFARX1 I_46118 (I786535,I2507,I786467,I786561,);
DFFARX1 I_46119 (I786561,I2507,I786467,I786456,);
DFFARX1 I_46120 (I311343,I2507,I786467,I786592,);
nand I_46121 (I786600,I786592,I311325);
not I_46122 (I786617,I786600);
DFFARX1 I_46123 (I786617,I2507,I786467,I786643,);
not I_46124 (I786651,I786643);
nor I_46125 (I786459,I786501,I786651);
DFFARX1 I_46126 (I311337,I2507,I786467,I786691,);
nor I_46127 (I786450,I786691,I786561);
nor I_46128 (I786441,I786691,I786617);
nand I_46129 (I786727,I311349,I311328);
and I_46130 (I786744,I786727,I311334);
DFFARX1 I_46131 (I786744,I2507,I786467,I786770,);
not I_46132 (I786778,I786770);
nand I_46133 (I786795,I786778,I786691);
nand I_46134 (I786444,I786778,I786600);
nor I_46135 (I786826,I311346,I311328);
and I_46136 (I786843,I786691,I786826);
nor I_46137 (I786860,I786778,I786843);
DFFARX1 I_46138 (I786860,I2507,I786467,I786453,);
nor I_46139 (I786891,I786493,I786826);
DFFARX1 I_46140 (I786891,I2507,I786467,I786438,);
nor I_46141 (I786922,I786770,I786826);
not I_46142 (I786939,I786922);
nand I_46143 (I786447,I786939,I786795);
not I_46144 (I786994,I2514);
DFFARX1 I_46145 (I1349357,I2507,I786994,I787020,);
not I_46146 (I787028,I787020);
nand I_46147 (I787045,I1349354,I1349363);
and I_46148 (I787062,I787045,I1349342);
DFFARX1 I_46149 (I787062,I2507,I786994,I787088,);
DFFARX1 I_46150 (I787088,I2507,I786994,I786983,);
DFFARX1 I_46151 (I1349345,I2507,I786994,I787119,);
nand I_46152 (I787127,I787119,I1349360);
not I_46153 (I787144,I787127);
DFFARX1 I_46154 (I787144,I2507,I786994,I787170,);
not I_46155 (I787178,I787170);
nor I_46156 (I786986,I787028,I787178);
DFFARX1 I_46157 (I1349366,I2507,I786994,I787218,);
nor I_46158 (I786977,I787218,I787088);
nor I_46159 (I786968,I787218,I787144);
nand I_46160 (I787254,I1349348,I1349369);
and I_46161 (I787271,I787254,I1349351);
DFFARX1 I_46162 (I787271,I2507,I786994,I787297,);
not I_46163 (I787305,I787297);
nand I_46164 (I787322,I787305,I787218);
nand I_46165 (I786971,I787305,I787127);
nor I_46166 (I787353,I1349342,I1349369);
and I_46167 (I787370,I787218,I787353);
nor I_46168 (I787387,I787305,I787370);
DFFARX1 I_46169 (I787387,I2507,I786994,I786980,);
nor I_46170 (I787418,I787020,I787353);
DFFARX1 I_46171 (I787418,I2507,I786994,I786965,);
nor I_46172 (I787449,I787297,I787353);
not I_46173 (I787466,I787449);
nand I_46174 (I786974,I787466,I787322);
not I_46175 (I787521,I2514);
DFFARX1 I_46176 (I1236814,I2507,I787521,I787547,);
not I_46177 (I787555,I787547);
nand I_46178 (I787572,I1236820,I1236802);
and I_46179 (I787589,I787572,I1236811);
DFFARX1 I_46180 (I787589,I2507,I787521,I787615,);
DFFARX1 I_46181 (I787615,I2507,I787521,I787510,);
DFFARX1 I_46182 (I1236817,I2507,I787521,I787646,);
nand I_46183 (I787654,I787646,I1236805);
not I_46184 (I787671,I787654);
DFFARX1 I_46185 (I787671,I2507,I787521,I787697,);
not I_46186 (I787705,I787697);
nor I_46187 (I787513,I787555,I787705);
DFFARX1 I_46188 (I1236823,I2507,I787521,I787745,);
nor I_46189 (I787504,I787745,I787615);
nor I_46190 (I787495,I787745,I787671);
nand I_46191 (I787781,I1236802,I1236808);
and I_46192 (I787798,I787781,I1236826);
DFFARX1 I_46193 (I787798,I2507,I787521,I787824,);
not I_46194 (I787832,I787824);
nand I_46195 (I787849,I787832,I787745);
nand I_46196 (I787498,I787832,I787654);
nor I_46197 (I787880,I1236805,I1236808);
and I_46198 (I787897,I787745,I787880);
nor I_46199 (I787914,I787832,I787897);
DFFARX1 I_46200 (I787914,I2507,I787521,I787507,);
nor I_46201 (I787945,I787547,I787880);
DFFARX1 I_46202 (I787945,I2507,I787521,I787492,);
nor I_46203 (I787976,I787824,I787880);
not I_46204 (I787993,I787976);
nand I_46205 (I787501,I787993,I787849);
not I_46206 (I788048,I2514);
DFFARX1 I_46207 (I693720,I2507,I788048,I788074,);
not I_46208 (I788082,I788074);
nand I_46209 (I788099,I693723,I693720);
and I_46210 (I788116,I788099,I693732);
DFFARX1 I_46211 (I788116,I2507,I788048,I788142,);
DFFARX1 I_46212 (I788142,I2507,I788048,I788037,);
DFFARX1 I_46213 (I693729,I2507,I788048,I788173,);
nand I_46214 (I788181,I788173,I693735);
not I_46215 (I788198,I788181);
DFFARX1 I_46216 (I788198,I2507,I788048,I788224,);
not I_46217 (I788232,I788224);
nor I_46218 (I788040,I788082,I788232);
DFFARX1 I_46219 (I693744,I2507,I788048,I788272,);
nor I_46220 (I788031,I788272,I788142);
nor I_46221 (I788022,I788272,I788198);
nand I_46222 (I788308,I693738,I693726);
and I_46223 (I788325,I788308,I693723);
DFFARX1 I_46224 (I788325,I2507,I788048,I788351,);
not I_46225 (I788359,I788351);
nand I_46226 (I788376,I788359,I788272);
nand I_46227 (I788025,I788359,I788181);
nor I_46228 (I788407,I693741,I693726);
and I_46229 (I788424,I788272,I788407);
nor I_46230 (I788441,I788359,I788424);
DFFARX1 I_46231 (I788441,I2507,I788048,I788034,);
nor I_46232 (I788472,I788074,I788407);
DFFARX1 I_46233 (I788472,I2507,I788048,I788019,);
nor I_46234 (I788503,I788351,I788407);
not I_46235 (I788520,I788503);
nand I_46236 (I788028,I788520,I788376);
not I_46237 (I788575,I2514);
DFFARX1 I_46238 (I1246062,I2507,I788575,I788601,);
not I_46239 (I788609,I788601);
nand I_46240 (I788626,I1246068,I1246050);
and I_46241 (I788643,I788626,I1246059);
DFFARX1 I_46242 (I788643,I2507,I788575,I788669,);
DFFARX1 I_46243 (I788669,I2507,I788575,I788564,);
DFFARX1 I_46244 (I1246065,I2507,I788575,I788700,);
nand I_46245 (I788708,I788700,I1246053);
not I_46246 (I788725,I788708);
DFFARX1 I_46247 (I788725,I2507,I788575,I788751,);
not I_46248 (I788759,I788751);
nor I_46249 (I788567,I788609,I788759);
DFFARX1 I_46250 (I1246071,I2507,I788575,I788799,);
nor I_46251 (I788558,I788799,I788669);
nor I_46252 (I788549,I788799,I788725);
nand I_46253 (I788835,I1246050,I1246056);
and I_46254 (I788852,I788835,I1246074);
DFFARX1 I_46255 (I788852,I2507,I788575,I788878,);
not I_46256 (I788886,I788878);
nand I_46257 (I788903,I788886,I788799);
nand I_46258 (I788552,I788886,I788708);
nor I_46259 (I788934,I1246053,I1246056);
and I_46260 (I788951,I788799,I788934);
nor I_46261 (I788968,I788886,I788951);
DFFARX1 I_46262 (I788968,I2507,I788575,I788561,);
nor I_46263 (I788999,I788601,I788934);
DFFARX1 I_46264 (I788999,I2507,I788575,I788546,);
nor I_46265 (I789030,I788878,I788934);
not I_46266 (I789047,I789030);
nand I_46267 (I788555,I789047,I788903);
not I_46268 (I789102,I2514);
DFFARX1 I_46269 (I1304791,I2507,I789102,I789128,);
not I_46270 (I789136,I789128);
nand I_46271 (I789153,I1304785,I1304803);
and I_46272 (I789170,I789153,I1304788);
DFFARX1 I_46273 (I789170,I2507,I789102,I789196,);
DFFARX1 I_46274 (I789196,I2507,I789102,I789091,);
DFFARX1 I_46275 (I1304809,I2507,I789102,I789227,);
nand I_46276 (I789235,I789227,I1304794);
not I_46277 (I789252,I789235);
DFFARX1 I_46278 (I789252,I2507,I789102,I789278,);
not I_46279 (I789286,I789278);
nor I_46280 (I789094,I789136,I789286);
DFFARX1 I_46281 (I1304806,I2507,I789102,I789326,);
nor I_46282 (I789085,I789326,I789196);
nor I_46283 (I789076,I789326,I789252);
nand I_46284 (I789362,I1304797,I1304812);
and I_46285 (I789379,I789362,I1304800);
DFFARX1 I_46286 (I789379,I2507,I789102,I789405,);
not I_46287 (I789413,I789405);
nand I_46288 (I789430,I789413,I789326);
nand I_46289 (I789079,I789413,I789235);
nor I_46290 (I789461,I1304785,I1304812);
and I_46291 (I789478,I789326,I789461);
nor I_46292 (I789495,I789413,I789478);
DFFARX1 I_46293 (I789495,I2507,I789102,I789088,);
nor I_46294 (I789526,I789128,I789461);
DFFARX1 I_46295 (I789526,I2507,I789102,I789073,);
nor I_46296 (I789557,I789405,I789461);
not I_46297 (I789574,I789557);
nand I_46298 (I789082,I789574,I789430);
not I_46299 (I789629,I2514);
DFFARX1 I_46300 (I395733,I2507,I789629,I789655,);
not I_46301 (I789663,I789655);
nand I_46302 (I789680,I395730,I395739);
and I_46303 (I789697,I789680,I395748);
DFFARX1 I_46304 (I789697,I2507,I789629,I789723,);
DFFARX1 I_46305 (I789723,I2507,I789629,I789618,);
DFFARX1 I_46306 (I395751,I2507,I789629,I789754,);
nand I_46307 (I789762,I789754,I395754);
not I_46308 (I789779,I789762);
DFFARX1 I_46309 (I789779,I2507,I789629,I789805,);
not I_46310 (I789813,I789805);
nor I_46311 (I789621,I789663,I789813);
DFFARX1 I_46312 (I395727,I2507,I789629,I789853,);
nor I_46313 (I789612,I789853,I789723);
nor I_46314 (I789603,I789853,I789779);
nand I_46315 (I789889,I395742,I395745);
and I_46316 (I789906,I789889,I395736);
DFFARX1 I_46317 (I789906,I2507,I789629,I789932,);
not I_46318 (I789940,I789932);
nand I_46319 (I789957,I789940,I789853);
nand I_46320 (I789606,I789940,I789762);
nor I_46321 (I789988,I395727,I395745);
and I_46322 (I790005,I789853,I789988);
nor I_46323 (I790022,I789940,I790005);
DFFARX1 I_46324 (I790022,I2507,I789629,I789615,);
nor I_46325 (I790053,I789655,I789988);
DFFARX1 I_46326 (I790053,I2507,I789629,I789600,);
nor I_46327 (I790084,I789932,I789988);
not I_46328 (I790101,I790084);
nand I_46329 (I789609,I790101,I789957);
not I_46330 (I790156,I2514);
DFFARX1 I_46331 (I197836,I2507,I790156,I790182,);
not I_46332 (I790190,I790182);
nand I_46333 (I790207,I197833,I197851);
and I_46334 (I790224,I790207,I197842);
DFFARX1 I_46335 (I790224,I2507,I790156,I790250,);
DFFARX1 I_46336 (I790250,I2507,I790156,I790145,);
DFFARX1 I_46337 (I197848,I2507,I790156,I790281,);
nand I_46338 (I790289,I790281,I197845);
not I_46339 (I790306,I790289);
DFFARX1 I_46340 (I790306,I2507,I790156,I790332,);
not I_46341 (I790340,I790332);
nor I_46342 (I790148,I790190,I790340);
DFFARX1 I_46343 (I197839,I2507,I790156,I790380,);
nor I_46344 (I790139,I790380,I790250);
nor I_46345 (I790130,I790380,I790306);
nand I_46346 (I790416,I197830,I197854);
and I_46347 (I790433,I790416,I197833);
DFFARX1 I_46348 (I790433,I2507,I790156,I790459,);
not I_46349 (I790467,I790459);
nand I_46350 (I790484,I790467,I790380);
nand I_46351 (I790133,I790467,I790289);
nor I_46352 (I790515,I197830,I197854);
and I_46353 (I790532,I790380,I790515);
nor I_46354 (I790549,I790467,I790532);
DFFARX1 I_46355 (I790549,I2507,I790156,I790142,);
nor I_46356 (I790580,I790182,I790515);
DFFARX1 I_46357 (I790580,I2507,I790156,I790127,);
nor I_46358 (I790611,I790459,I790515);
not I_46359 (I790628,I790611);
nand I_46360 (I790136,I790628,I790484);
not I_46361 (I790683,I2514);
DFFARX1 I_46362 (I507185,I2507,I790683,I790709,);
not I_46363 (I790717,I790709);
nand I_46364 (I790734,I507203,I507194);
and I_46365 (I790751,I790734,I507197);
DFFARX1 I_46366 (I790751,I2507,I790683,I790777,);
DFFARX1 I_46367 (I790777,I2507,I790683,I790672,);
DFFARX1 I_46368 (I507191,I2507,I790683,I790808,);
nand I_46369 (I790816,I790808,I507182);
not I_46370 (I790833,I790816);
DFFARX1 I_46371 (I790833,I2507,I790683,I790859,);
not I_46372 (I790867,I790859);
nor I_46373 (I790675,I790717,I790867);
DFFARX1 I_46374 (I507188,I2507,I790683,I790907,);
nor I_46375 (I790666,I790907,I790777);
nor I_46376 (I790657,I790907,I790833);
nand I_46377 (I790943,I507182,I507179);
and I_46378 (I790960,I790943,I507200);
DFFARX1 I_46379 (I790960,I2507,I790683,I790986,);
not I_46380 (I790994,I790986);
nand I_46381 (I791011,I790994,I790907);
nand I_46382 (I790660,I790994,I790816);
nor I_46383 (I791042,I507179,I507179);
and I_46384 (I791059,I790907,I791042);
nor I_46385 (I791076,I790994,I791059);
DFFARX1 I_46386 (I791076,I2507,I790683,I790669,);
nor I_46387 (I791107,I790709,I791042);
DFFARX1 I_46388 (I791107,I2507,I790683,I790654,);
nor I_46389 (I791138,I790986,I791042);
not I_46390 (I791155,I791138);
nand I_46391 (I790663,I791155,I791011);
not I_46392 (I791210,I2514);
DFFARX1 I_46393 (I187721,I2507,I791210,I791236,);
not I_46394 (I791244,I791236);
nand I_46395 (I791261,I187718,I187736);
and I_46396 (I791278,I791261,I187727);
DFFARX1 I_46397 (I791278,I2507,I791210,I791304,);
DFFARX1 I_46398 (I791304,I2507,I791210,I791199,);
DFFARX1 I_46399 (I187733,I2507,I791210,I791335,);
nand I_46400 (I791343,I791335,I187730);
not I_46401 (I791360,I791343);
DFFARX1 I_46402 (I791360,I2507,I791210,I791386,);
not I_46403 (I791394,I791386);
nor I_46404 (I791202,I791244,I791394);
DFFARX1 I_46405 (I187724,I2507,I791210,I791434,);
nor I_46406 (I791193,I791434,I791304);
nor I_46407 (I791184,I791434,I791360);
nand I_46408 (I791470,I187715,I187739);
and I_46409 (I791487,I791470,I187718);
DFFARX1 I_46410 (I791487,I2507,I791210,I791513,);
not I_46411 (I791521,I791513);
nand I_46412 (I791538,I791521,I791434);
nand I_46413 (I791187,I791521,I791343);
nor I_46414 (I791569,I187715,I187739);
and I_46415 (I791586,I791434,I791569);
nor I_46416 (I791603,I791521,I791586);
DFFARX1 I_46417 (I791603,I2507,I791210,I791196,);
nor I_46418 (I791634,I791236,I791569);
DFFARX1 I_46419 (I791634,I2507,I791210,I791181,);
nor I_46420 (I791665,I791513,I791569);
not I_46421 (I791682,I791665);
nand I_46422 (I791190,I791682,I791538);
not I_46423 (I791737,I2514);
DFFARX1 I_46424 (I928918,I2507,I791737,I791763,);
not I_46425 (I791771,I791763);
nand I_46426 (I791788,I928933,I928915);
and I_46427 (I791805,I791788,I928915);
DFFARX1 I_46428 (I791805,I2507,I791737,I791831,);
DFFARX1 I_46429 (I791831,I2507,I791737,I791726,);
DFFARX1 I_46430 (I928924,I2507,I791737,I791862,);
nand I_46431 (I791870,I791862,I928942);
not I_46432 (I791887,I791870);
DFFARX1 I_46433 (I791887,I2507,I791737,I791913,);
not I_46434 (I791921,I791913);
nor I_46435 (I791729,I791771,I791921);
DFFARX1 I_46436 (I928939,I2507,I791737,I791961,);
nor I_46437 (I791720,I791961,I791831);
nor I_46438 (I791711,I791961,I791887);
nand I_46439 (I791997,I928936,I928927);
and I_46440 (I792014,I791997,I928921);
DFFARX1 I_46441 (I792014,I2507,I791737,I792040,);
not I_46442 (I792048,I792040);
nand I_46443 (I792065,I792048,I791961);
nand I_46444 (I791714,I792048,I791870);
nor I_46445 (I792096,I928930,I928927);
and I_46446 (I792113,I791961,I792096);
nor I_46447 (I792130,I792048,I792113);
DFFARX1 I_46448 (I792130,I2507,I791737,I791723,);
nor I_46449 (I792161,I791763,I792096);
DFFARX1 I_46450 (I792161,I2507,I791737,I791708,);
nor I_46451 (I792192,I792040,I792096);
not I_46452 (I792209,I792192);
nand I_46453 (I791717,I792209,I792065);
not I_46454 (I792264,I2514);
DFFARX1 I_46455 (I27992,I2507,I792264,I792290,);
not I_46456 (I792298,I792290);
nand I_46457 (I792315,I28004,I28007);
and I_46458 (I792332,I792315,I27983);
DFFARX1 I_46459 (I792332,I2507,I792264,I792358,);
DFFARX1 I_46460 (I792358,I2507,I792264,I792253,);
DFFARX1 I_46461 (I28001,I2507,I792264,I792389,);
nand I_46462 (I792397,I792389,I27989);
not I_46463 (I792414,I792397);
DFFARX1 I_46464 (I792414,I2507,I792264,I792440,);
not I_46465 (I792448,I792440);
nor I_46466 (I792256,I792298,I792448);
DFFARX1 I_46467 (I27986,I2507,I792264,I792488,);
nor I_46468 (I792247,I792488,I792358);
nor I_46469 (I792238,I792488,I792414);
nand I_46470 (I792524,I27995,I27986);
and I_46471 (I792541,I792524,I27983);
DFFARX1 I_46472 (I792541,I2507,I792264,I792567,);
not I_46473 (I792575,I792567);
nand I_46474 (I792592,I792575,I792488);
nand I_46475 (I792241,I792575,I792397);
nor I_46476 (I792623,I27998,I27986);
and I_46477 (I792640,I792488,I792623);
nor I_46478 (I792657,I792575,I792640);
DFFARX1 I_46479 (I792657,I2507,I792264,I792250,);
nor I_46480 (I792688,I792290,I792623);
DFFARX1 I_46481 (I792688,I2507,I792264,I792235,);
nor I_46482 (I792719,I792567,I792623);
not I_46483 (I792736,I792719);
nand I_46484 (I792244,I792736,I792592);
not I_46485 (I792791,I2514);
DFFARX1 I_46486 (I140734,I2507,I792791,I792817,);
not I_46487 (I792825,I792817);
nand I_46488 (I792842,I140710,I140728);
and I_46489 (I792859,I792842,I140716);
DFFARX1 I_46490 (I792859,I2507,I792791,I792885,);
DFFARX1 I_46491 (I792885,I2507,I792791,I792780,);
DFFARX1 I_46492 (I140725,I2507,I792791,I792916,);
nand I_46493 (I792924,I792916,I140731);
not I_46494 (I792941,I792924);
DFFARX1 I_46495 (I792941,I2507,I792791,I792967,);
not I_46496 (I792975,I792967);
nor I_46497 (I792783,I792825,I792975);
DFFARX1 I_46498 (I140710,I2507,I792791,I793015,);
nor I_46499 (I792774,I793015,I792885);
nor I_46500 (I792765,I793015,I792941);
nand I_46501 (I793051,I140722,I140713);
and I_46502 (I793068,I793051,I140737);
DFFARX1 I_46503 (I793068,I2507,I792791,I793094,);
not I_46504 (I793102,I793094);
nand I_46505 (I793119,I793102,I793015);
nand I_46506 (I792768,I793102,I792924);
nor I_46507 (I793150,I140719,I140713);
and I_46508 (I793167,I793015,I793150);
nor I_46509 (I793184,I793102,I793167);
DFFARX1 I_46510 (I793184,I2507,I792791,I792777,);
nor I_46511 (I793215,I792817,I793150);
DFFARX1 I_46512 (I793215,I2507,I792791,I792762,);
nor I_46513 (I793246,I793094,I793150);
not I_46514 (I793263,I793246);
nand I_46515 (I792771,I793263,I793119);
not I_46516 (I793318,I2514);
DFFARX1 I_46517 (I625531,I2507,I793318,I793344,);
not I_46518 (I793352,I793344);
nand I_46519 (I793369,I625516,I625537);
and I_46520 (I793386,I793369,I625525);
DFFARX1 I_46521 (I793386,I2507,I793318,I793412,);
DFFARX1 I_46522 (I793412,I2507,I793318,I793307,);
DFFARX1 I_46523 (I625519,I2507,I793318,I793443,);
nand I_46524 (I793451,I793443,I625528);
not I_46525 (I793468,I793451);
DFFARX1 I_46526 (I793468,I2507,I793318,I793494,);
not I_46527 (I793502,I793494);
nor I_46528 (I793310,I793352,I793502);
DFFARX1 I_46529 (I625534,I2507,I793318,I793542,);
nor I_46530 (I793301,I793542,I793412);
nor I_46531 (I793292,I793542,I793468);
nand I_46532 (I793578,I625516,I625519);
and I_46533 (I793595,I793578,I625540);
DFFARX1 I_46534 (I793595,I2507,I793318,I793621,);
not I_46535 (I793629,I793621);
nand I_46536 (I793646,I793629,I793542);
nand I_46537 (I793295,I793629,I793451);
nor I_46538 (I793677,I625522,I625519);
and I_46539 (I793694,I793542,I793677);
nor I_46540 (I793711,I793629,I793694);
DFFARX1 I_46541 (I793711,I2507,I793318,I793304,);
nor I_46542 (I793742,I793344,I793677);
DFFARX1 I_46543 (I793742,I2507,I793318,I793289,);
nor I_46544 (I793773,I793621,I793677);
not I_46545 (I793790,I793773);
nand I_46546 (I793298,I793790,I793646);
not I_46547 (I793845,I2514);
DFFARX1 I_46548 (I7292,I2507,I793845,I793871,);
not I_46549 (I793879,I793871);
nand I_46550 (I793896,I7298,I7280);
and I_46551 (I793913,I793896,I7289);
DFFARX1 I_46552 (I793913,I2507,I793845,I793939,);
DFFARX1 I_46553 (I793939,I2507,I793845,I793834,);
DFFARX1 I_46554 (I7280,I2507,I793845,I793970,);
nand I_46555 (I793978,I793970,I7283);
not I_46556 (I793995,I793978);
DFFARX1 I_46557 (I793995,I2507,I793845,I794021,);
not I_46558 (I794029,I794021);
nor I_46559 (I793837,I793879,I794029);
DFFARX1 I_46560 (I7283,I2507,I793845,I794069,);
nor I_46561 (I793828,I794069,I793939);
nor I_46562 (I793819,I794069,I793995);
nand I_46563 (I794105,I7286,I7295);
and I_46564 (I794122,I794105,I7277);
DFFARX1 I_46565 (I794122,I2507,I793845,I794148,);
not I_46566 (I794156,I794148);
nand I_46567 (I794173,I794156,I794069);
nand I_46568 (I793822,I794156,I793978);
nor I_46569 (I794204,I7277,I7295);
and I_46570 (I794221,I794069,I794204);
nor I_46571 (I794238,I794156,I794221);
DFFARX1 I_46572 (I794238,I2507,I793845,I793831,);
nor I_46573 (I794269,I793871,I794204);
DFFARX1 I_46574 (I794269,I2507,I793845,I793816,);
nor I_46575 (I794300,I794148,I794204);
not I_46576 (I794317,I794300);
nand I_46577 (I793825,I794317,I794173);
not I_46578 (I794372,I2514);
DFFARX1 I_46579 (I550969,I2507,I794372,I794398,);
not I_46580 (I794406,I794398);
nand I_46581 (I794423,I550954,I550975);
and I_46582 (I794440,I794423,I550963);
DFFARX1 I_46583 (I794440,I2507,I794372,I794466,);
DFFARX1 I_46584 (I794466,I2507,I794372,I794361,);
DFFARX1 I_46585 (I550957,I2507,I794372,I794497,);
nand I_46586 (I794505,I794497,I550966);
not I_46587 (I794522,I794505);
DFFARX1 I_46588 (I794522,I2507,I794372,I794548,);
not I_46589 (I794556,I794548);
nor I_46590 (I794364,I794406,I794556);
DFFARX1 I_46591 (I550972,I2507,I794372,I794596,);
nor I_46592 (I794355,I794596,I794466);
nor I_46593 (I794346,I794596,I794522);
nand I_46594 (I794632,I550954,I550957);
and I_46595 (I794649,I794632,I550978);
DFFARX1 I_46596 (I794649,I2507,I794372,I794675,);
not I_46597 (I794683,I794675);
nand I_46598 (I794700,I794683,I794596);
nand I_46599 (I794349,I794683,I794505);
nor I_46600 (I794731,I550960,I550957);
and I_46601 (I794748,I794596,I794731);
nor I_46602 (I794765,I794683,I794748);
DFFARX1 I_46603 (I794765,I2507,I794372,I794358,);
nor I_46604 (I794796,I794398,I794731);
DFFARX1 I_46605 (I794796,I2507,I794372,I794343,);
nor I_46606 (I794827,I794675,I794731);
not I_46607 (I794844,I794827);
nand I_46608 (I794352,I794844,I794700);
not I_46609 (I794899,I2514);
DFFARX1 I_46610 (I348221,I2507,I794899,I794925,);
not I_46611 (I794933,I794925);
nand I_46612 (I794950,I348212,I348212);
and I_46613 (I794967,I794950,I348230);
DFFARX1 I_46614 (I794967,I2507,I794899,I794993,);
DFFARX1 I_46615 (I794993,I2507,I794899,I794888,);
DFFARX1 I_46616 (I348233,I2507,I794899,I795024,);
nand I_46617 (I795032,I795024,I348215);
not I_46618 (I795049,I795032);
DFFARX1 I_46619 (I795049,I2507,I794899,I795075,);
not I_46620 (I795083,I795075);
nor I_46621 (I794891,I794933,I795083);
DFFARX1 I_46622 (I348227,I2507,I794899,I795123,);
nor I_46623 (I794882,I795123,I794993);
nor I_46624 (I794873,I795123,I795049);
nand I_46625 (I795159,I348239,I348218);
and I_46626 (I795176,I795159,I348224);
DFFARX1 I_46627 (I795176,I2507,I794899,I795202,);
not I_46628 (I795210,I795202);
nand I_46629 (I795227,I795210,I795123);
nand I_46630 (I794876,I795210,I795032);
nor I_46631 (I795258,I348236,I348218);
and I_46632 (I795275,I795123,I795258);
nor I_46633 (I795292,I795210,I795275);
DFFARX1 I_46634 (I795292,I2507,I794899,I794885,);
nor I_46635 (I795323,I794925,I795258);
DFFARX1 I_46636 (I795323,I2507,I794899,I794870,);
nor I_46637 (I795354,I795202,I795258);
not I_46638 (I795371,I795354);
nand I_46639 (I794879,I795371,I795227);
not I_46640 (I795426,I2514);
DFFARX1 I_46641 (I292886,I2507,I795426,I795452,);
not I_46642 (I795460,I795452);
nand I_46643 (I795477,I292877,I292877);
and I_46644 (I795494,I795477,I292895);
DFFARX1 I_46645 (I795494,I2507,I795426,I795520,);
DFFARX1 I_46646 (I795520,I2507,I795426,I795415,);
DFFARX1 I_46647 (I292898,I2507,I795426,I795551,);
nand I_46648 (I795559,I795551,I292880);
not I_46649 (I795576,I795559);
DFFARX1 I_46650 (I795576,I2507,I795426,I795602,);
not I_46651 (I795610,I795602);
nor I_46652 (I795418,I795460,I795610);
DFFARX1 I_46653 (I292892,I2507,I795426,I795650,);
nor I_46654 (I795409,I795650,I795520);
nor I_46655 (I795400,I795650,I795576);
nand I_46656 (I795686,I292904,I292883);
and I_46657 (I795703,I795686,I292889);
DFFARX1 I_46658 (I795703,I2507,I795426,I795729,);
not I_46659 (I795737,I795729);
nand I_46660 (I795754,I795737,I795650);
nand I_46661 (I795403,I795737,I795559);
nor I_46662 (I795785,I292901,I292883);
and I_46663 (I795802,I795650,I795785);
nor I_46664 (I795819,I795737,I795802);
DFFARX1 I_46665 (I795819,I2507,I795426,I795412,);
nor I_46666 (I795850,I795452,I795785);
DFFARX1 I_46667 (I795850,I2507,I795426,I795397,);
nor I_46668 (I795881,I795729,I795785);
not I_46669 (I795898,I795881);
nand I_46670 (I795406,I795898,I795754);
not I_46671 (I795953,I2514);
DFFARX1 I_46672 (I1178612,I2507,I795953,I795979,);
not I_46673 (I795987,I795979);
nand I_46674 (I796004,I1178594,I1178594);
and I_46675 (I796021,I796004,I1178600);
DFFARX1 I_46676 (I796021,I2507,I795953,I796047,);
DFFARX1 I_46677 (I796047,I2507,I795953,I795942,);
DFFARX1 I_46678 (I1178597,I2507,I795953,I796078,);
nand I_46679 (I796086,I796078,I1178606);
not I_46680 (I796103,I796086);
DFFARX1 I_46681 (I796103,I2507,I795953,I796129,);
not I_46682 (I796137,I796129);
nor I_46683 (I795945,I795987,I796137);
DFFARX1 I_46684 (I1178618,I2507,I795953,I796177,);
nor I_46685 (I795936,I796177,I796047);
nor I_46686 (I795927,I796177,I796103);
nand I_46687 (I796213,I1178609,I1178603);
and I_46688 (I796230,I796213,I1178597);
DFFARX1 I_46689 (I796230,I2507,I795953,I796256,);
not I_46690 (I796264,I796256);
nand I_46691 (I796281,I796264,I796177);
nand I_46692 (I795930,I796264,I796086);
nor I_46693 (I796312,I1178615,I1178603);
and I_46694 (I796329,I796177,I796312);
nor I_46695 (I796346,I796264,I796329);
DFFARX1 I_46696 (I796346,I2507,I795953,I795939,);
nor I_46697 (I796377,I795979,I796312);
DFFARX1 I_46698 (I796377,I2507,I795953,I795924,);
nor I_46699 (I796408,I796256,I796312);
not I_46700 (I796425,I796408);
nand I_46701 (I795933,I796425,I796281);
not I_46702 (I796480,I2514);
DFFARX1 I_46703 (I485493,I2507,I796480,I796506,);
not I_46704 (I796514,I796506);
nand I_46705 (I796531,I485490,I485499);
and I_46706 (I796548,I796531,I485508);
DFFARX1 I_46707 (I796548,I2507,I796480,I796574,);
DFFARX1 I_46708 (I796574,I2507,I796480,I796469,);
DFFARX1 I_46709 (I485511,I2507,I796480,I796605,);
nand I_46710 (I796613,I796605,I485514);
not I_46711 (I796630,I796613);
DFFARX1 I_46712 (I796630,I2507,I796480,I796656,);
not I_46713 (I796664,I796656);
nor I_46714 (I796472,I796514,I796664);
DFFARX1 I_46715 (I485487,I2507,I796480,I796704,);
nor I_46716 (I796463,I796704,I796574);
nor I_46717 (I796454,I796704,I796630);
nand I_46718 (I796740,I485502,I485505);
and I_46719 (I796757,I796740,I485496);
DFFARX1 I_46720 (I796757,I2507,I796480,I796783,);
not I_46721 (I796791,I796783);
nand I_46722 (I796808,I796791,I796704);
nand I_46723 (I796457,I796791,I796613);
nor I_46724 (I796839,I485487,I485505);
and I_46725 (I796856,I796704,I796839);
nor I_46726 (I796873,I796791,I796856);
DFFARX1 I_46727 (I796873,I2507,I796480,I796466,);
nor I_46728 (I796904,I796506,I796839);
DFFARX1 I_46729 (I796904,I2507,I796480,I796451,);
nor I_46730 (I796935,I796783,I796839);
not I_46731 (I796952,I796935);
nand I_46732 (I796460,I796952,I796808);
not I_46733 (I797007,I2514);
DFFARX1 I_46734 (I1215054,I2507,I797007,I797033,);
not I_46735 (I797041,I797033);
nand I_46736 (I797058,I1215060,I1215042);
and I_46737 (I797075,I797058,I1215051);
DFFARX1 I_46738 (I797075,I2507,I797007,I797101,);
DFFARX1 I_46739 (I797101,I2507,I797007,I796996,);
DFFARX1 I_46740 (I1215057,I2507,I797007,I797132,);
nand I_46741 (I797140,I797132,I1215045);
not I_46742 (I797157,I797140);
DFFARX1 I_46743 (I797157,I2507,I797007,I797183,);
not I_46744 (I797191,I797183);
nor I_46745 (I796999,I797041,I797191);
DFFARX1 I_46746 (I1215063,I2507,I797007,I797231,);
nor I_46747 (I796990,I797231,I797101);
nor I_46748 (I796981,I797231,I797157);
nand I_46749 (I797267,I1215042,I1215048);
and I_46750 (I797284,I797267,I1215066);
DFFARX1 I_46751 (I797284,I2507,I797007,I797310,);
not I_46752 (I797318,I797310);
nand I_46753 (I797335,I797318,I797231);
nand I_46754 (I796984,I797318,I797140);
nor I_46755 (I797366,I1215045,I1215048);
and I_46756 (I797383,I797231,I797366);
nor I_46757 (I797400,I797318,I797383);
DFFARX1 I_46758 (I797400,I2507,I797007,I796993,);
nor I_46759 (I797431,I797033,I797366);
DFFARX1 I_46760 (I797431,I2507,I797007,I796978,);
nor I_46761 (I797462,I797310,I797366);
not I_46762 (I797479,I797462);
nand I_46763 (I796987,I797479,I797335);
not I_46764 (I797534,I2514);
DFFARX1 I_46765 (I583337,I2507,I797534,I797560,);
not I_46766 (I797568,I797560);
nand I_46767 (I797585,I583322,I583343);
and I_46768 (I797602,I797585,I583331);
DFFARX1 I_46769 (I797602,I2507,I797534,I797628,);
DFFARX1 I_46770 (I797628,I2507,I797534,I797523,);
DFFARX1 I_46771 (I583325,I2507,I797534,I797659,);
nand I_46772 (I797667,I797659,I583334);
not I_46773 (I797684,I797667);
DFFARX1 I_46774 (I797684,I2507,I797534,I797710,);
not I_46775 (I797718,I797710);
nor I_46776 (I797526,I797568,I797718);
DFFARX1 I_46777 (I583340,I2507,I797534,I797758,);
nor I_46778 (I797517,I797758,I797628);
nor I_46779 (I797508,I797758,I797684);
nand I_46780 (I797794,I583322,I583325);
and I_46781 (I797811,I797794,I583346);
DFFARX1 I_46782 (I797811,I2507,I797534,I797837,);
not I_46783 (I797845,I797837);
nand I_46784 (I797862,I797845,I797758);
nand I_46785 (I797511,I797845,I797667);
nor I_46786 (I797893,I583328,I583325);
and I_46787 (I797910,I797758,I797893);
nor I_46788 (I797927,I797845,I797910);
DFFARX1 I_46789 (I797927,I2507,I797534,I797520,);
nor I_46790 (I797958,I797560,I797893);
DFFARX1 I_46791 (I797958,I2507,I797534,I797505,);
nor I_46792 (I797989,I797837,I797893);
not I_46793 (I798006,I797989);
nand I_46794 (I797514,I798006,I797862);
not I_46795 (I798061,I2514);
DFFARX1 I_46796 (I995456,I2507,I798061,I798087,);
not I_46797 (I798095,I798087);
nand I_46798 (I798112,I995471,I995453);
and I_46799 (I798129,I798112,I995453);
DFFARX1 I_46800 (I798129,I2507,I798061,I798155,);
DFFARX1 I_46801 (I798155,I2507,I798061,I798050,);
DFFARX1 I_46802 (I995462,I2507,I798061,I798186,);
nand I_46803 (I798194,I798186,I995480);
not I_46804 (I798211,I798194);
DFFARX1 I_46805 (I798211,I2507,I798061,I798237,);
not I_46806 (I798245,I798237);
nor I_46807 (I798053,I798095,I798245);
DFFARX1 I_46808 (I995477,I2507,I798061,I798285,);
nor I_46809 (I798044,I798285,I798155);
nor I_46810 (I798035,I798285,I798211);
nand I_46811 (I798321,I995474,I995465);
and I_46812 (I798338,I798321,I995459);
DFFARX1 I_46813 (I798338,I2507,I798061,I798364,);
not I_46814 (I798372,I798364);
nand I_46815 (I798389,I798372,I798285);
nand I_46816 (I798038,I798372,I798194);
nor I_46817 (I798420,I995468,I995465);
and I_46818 (I798437,I798285,I798420);
nor I_46819 (I798454,I798372,I798437);
DFFARX1 I_46820 (I798454,I2507,I798061,I798047,);
nor I_46821 (I798485,I798087,I798420);
DFFARX1 I_46822 (I798485,I2507,I798061,I798032,);
nor I_46823 (I798516,I798364,I798420);
not I_46824 (I798533,I798516);
nand I_46825 (I798041,I798533,I798389);
not I_46826 (I798588,I2514);
DFFARX1 I_46827 (I654416,I2507,I798588,I798614,);
not I_46828 (I798622,I798614);
nand I_46829 (I798639,I654419,I654416);
and I_46830 (I798656,I798639,I654428);
DFFARX1 I_46831 (I798656,I2507,I798588,I798682,);
DFFARX1 I_46832 (I798682,I2507,I798588,I798577,);
DFFARX1 I_46833 (I654425,I2507,I798588,I798713,);
nand I_46834 (I798721,I798713,I654431);
not I_46835 (I798738,I798721);
DFFARX1 I_46836 (I798738,I2507,I798588,I798764,);
not I_46837 (I798772,I798764);
nor I_46838 (I798580,I798622,I798772);
DFFARX1 I_46839 (I654440,I2507,I798588,I798812,);
nor I_46840 (I798571,I798812,I798682);
nor I_46841 (I798562,I798812,I798738);
nand I_46842 (I798848,I654434,I654422);
and I_46843 (I798865,I798848,I654419);
DFFARX1 I_46844 (I798865,I2507,I798588,I798891,);
not I_46845 (I798899,I798891);
nand I_46846 (I798916,I798899,I798812);
nand I_46847 (I798565,I798899,I798721);
nor I_46848 (I798947,I654437,I654422);
and I_46849 (I798964,I798812,I798947);
nor I_46850 (I798981,I798899,I798964);
DFFARX1 I_46851 (I798981,I2507,I798588,I798574,);
nor I_46852 (I799012,I798614,I798947);
DFFARX1 I_46853 (I799012,I2507,I798588,I798559,);
nor I_46854 (I799043,I798891,I798947);
not I_46855 (I799060,I799043);
nand I_46856 (I798568,I799060,I798916);
not I_46857 (I799115,I2514);
DFFARX1 I_46858 (I1027541,I2507,I799115,I799141,);
not I_46859 (I799149,I799141);
nand I_46860 (I799166,I1027550,I1027538);
and I_46861 (I799183,I799166,I1027535);
DFFARX1 I_46862 (I799183,I2507,I799115,I799209,);
DFFARX1 I_46863 (I799209,I2507,I799115,I799104,);
DFFARX1 I_46864 (I1027535,I2507,I799115,I799240,);
nand I_46865 (I799248,I799240,I1027532);
not I_46866 (I799265,I799248);
DFFARX1 I_46867 (I799265,I2507,I799115,I799291,);
not I_46868 (I799299,I799291);
nor I_46869 (I799107,I799149,I799299);
DFFARX1 I_46870 (I1027538,I2507,I799115,I799339,);
nor I_46871 (I799098,I799339,I799209);
nor I_46872 (I799089,I799339,I799265);
nand I_46873 (I799375,I1027553,I1027544);
and I_46874 (I799392,I799375,I1027547);
DFFARX1 I_46875 (I799392,I2507,I799115,I799418,);
not I_46876 (I799426,I799418);
nand I_46877 (I799443,I799426,I799339);
nand I_46878 (I799092,I799426,I799248);
nor I_46879 (I799474,I1027532,I1027544);
and I_46880 (I799491,I799339,I799474);
nor I_46881 (I799508,I799426,I799491);
DFFARX1 I_46882 (I799508,I2507,I799115,I799101,);
nor I_46883 (I799539,I799141,I799474);
DFFARX1 I_46884 (I799539,I2507,I799115,I799086,);
nor I_46885 (I799570,I799418,I799474);
not I_46886 (I799587,I799570);
nand I_46887 (I799095,I799587,I799443);
not I_46888 (I799642,I2514);
DFFARX1 I_46889 (I250726,I2507,I799642,I799668,);
not I_46890 (I799676,I799668);
nand I_46891 (I799693,I250717,I250717);
and I_46892 (I799710,I799693,I250735);
DFFARX1 I_46893 (I799710,I2507,I799642,I799736,);
DFFARX1 I_46894 (I799736,I2507,I799642,I799631,);
DFFARX1 I_46895 (I250738,I2507,I799642,I799767,);
nand I_46896 (I799775,I799767,I250720);
not I_46897 (I799792,I799775);
DFFARX1 I_46898 (I799792,I2507,I799642,I799818,);
not I_46899 (I799826,I799818);
nor I_46900 (I799634,I799676,I799826);
DFFARX1 I_46901 (I250732,I2507,I799642,I799866,);
nor I_46902 (I799625,I799866,I799736);
nor I_46903 (I799616,I799866,I799792);
nand I_46904 (I799902,I250744,I250723);
and I_46905 (I799919,I799902,I250729);
DFFARX1 I_46906 (I799919,I2507,I799642,I799945,);
not I_46907 (I799953,I799945);
nand I_46908 (I799970,I799953,I799866);
nand I_46909 (I799619,I799953,I799775);
nor I_46910 (I800001,I250741,I250723);
and I_46911 (I800018,I799866,I800001);
nor I_46912 (I800035,I799953,I800018);
DFFARX1 I_46913 (I800035,I2507,I799642,I799628,);
nor I_46914 (I800066,I799668,I800001);
DFFARX1 I_46915 (I800066,I2507,I799642,I799613,);
nor I_46916 (I800097,I799945,I800001);
not I_46917 (I800114,I800097);
nand I_46918 (I799622,I800114,I799970);
not I_46919 (I800169,I2514);
DFFARX1 I_46920 (I1104628,I2507,I800169,I800195,);
not I_46921 (I800203,I800195);
nand I_46922 (I800220,I1104610,I1104610);
and I_46923 (I800237,I800220,I1104616);
DFFARX1 I_46924 (I800237,I2507,I800169,I800263,);
DFFARX1 I_46925 (I800263,I2507,I800169,I800158,);
DFFARX1 I_46926 (I1104613,I2507,I800169,I800294,);
nand I_46927 (I800302,I800294,I1104622);
not I_46928 (I800319,I800302);
DFFARX1 I_46929 (I800319,I2507,I800169,I800345,);
not I_46930 (I800353,I800345);
nor I_46931 (I800161,I800203,I800353);
DFFARX1 I_46932 (I1104634,I2507,I800169,I800393,);
nor I_46933 (I800152,I800393,I800263);
nor I_46934 (I800143,I800393,I800319);
nand I_46935 (I800429,I1104625,I1104619);
and I_46936 (I800446,I800429,I1104613);
DFFARX1 I_46937 (I800446,I2507,I800169,I800472,);
not I_46938 (I800480,I800472);
nand I_46939 (I800497,I800480,I800393);
nand I_46940 (I800146,I800480,I800302);
nor I_46941 (I800528,I1104631,I1104619);
and I_46942 (I800545,I800393,I800528);
nor I_46943 (I800562,I800480,I800545);
DFFARX1 I_46944 (I800562,I2507,I800169,I800155,);
nor I_46945 (I800593,I800195,I800528);
DFFARX1 I_46946 (I800593,I2507,I800169,I800140,);
nor I_46947 (I800624,I800472,I800528);
not I_46948 (I800641,I800624);
nand I_46949 (I800149,I800641,I800497);
not I_46950 (I800696,I2514);
DFFARX1 I_46951 (I999978,I2507,I800696,I800722,);
not I_46952 (I800730,I800722);
nand I_46953 (I800747,I999993,I999975);
and I_46954 (I800764,I800747,I999975);
DFFARX1 I_46955 (I800764,I2507,I800696,I800790,);
DFFARX1 I_46956 (I800790,I2507,I800696,I800685,);
DFFARX1 I_46957 (I999984,I2507,I800696,I800821,);
nand I_46958 (I800829,I800821,I1000002);
not I_46959 (I800846,I800829);
DFFARX1 I_46960 (I800846,I2507,I800696,I800872,);
not I_46961 (I800880,I800872);
nor I_46962 (I800688,I800730,I800880);
DFFARX1 I_46963 (I999999,I2507,I800696,I800920,);
nor I_46964 (I800679,I800920,I800790);
nor I_46965 (I800670,I800920,I800846);
nand I_46966 (I800956,I999996,I999987);
and I_46967 (I800973,I800956,I999981);
DFFARX1 I_46968 (I800973,I2507,I800696,I800999,);
not I_46969 (I801007,I800999);
nand I_46970 (I801024,I801007,I800920);
nand I_46971 (I800673,I801007,I800829);
nor I_46972 (I801055,I999990,I999987);
and I_46973 (I801072,I800920,I801055);
nor I_46974 (I801089,I801007,I801072);
DFFARX1 I_46975 (I801089,I2507,I800696,I800682,);
nor I_46976 (I801120,I800722,I801055);
DFFARX1 I_46977 (I801120,I2507,I800696,I800667,);
nor I_46978 (I801151,I800999,I801055);
not I_46979 (I801168,I801151);
nand I_46980 (I800676,I801168,I801024);
not I_46981 (I801223,I2514);
DFFARX1 I_46982 (I726088,I2507,I801223,I801249,);
not I_46983 (I801257,I801249);
nand I_46984 (I801274,I726091,I726088);
and I_46985 (I801291,I801274,I726100);
DFFARX1 I_46986 (I801291,I2507,I801223,I801317,);
DFFARX1 I_46987 (I801317,I2507,I801223,I801212,);
DFFARX1 I_46988 (I726097,I2507,I801223,I801348,);
nand I_46989 (I801356,I801348,I726103);
not I_46990 (I801373,I801356);
DFFARX1 I_46991 (I801373,I2507,I801223,I801399,);
not I_46992 (I801407,I801399);
nor I_46993 (I801215,I801257,I801407);
DFFARX1 I_46994 (I726112,I2507,I801223,I801447,);
nor I_46995 (I801206,I801447,I801317);
nor I_46996 (I801197,I801447,I801373);
nand I_46997 (I801483,I726106,I726094);
and I_46998 (I801500,I801483,I726091);
DFFARX1 I_46999 (I801500,I2507,I801223,I801526,);
not I_47000 (I801534,I801526);
nand I_47001 (I801551,I801534,I801447);
nand I_47002 (I801200,I801534,I801356);
nor I_47003 (I801582,I726109,I726094);
and I_47004 (I801599,I801447,I801582);
nor I_47005 (I801616,I801534,I801599);
DFFARX1 I_47006 (I801616,I2507,I801223,I801209,);
nor I_47007 (I801647,I801249,I801582);
DFFARX1 I_47008 (I801647,I2507,I801223,I801194,);
nor I_47009 (I801678,I801526,I801582);
not I_47010 (I801695,I801678);
nand I_47011 (I801203,I801695,I801551);
not I_47012 (I801750,I2514);
DFFARX1 I_47013 (I298156,I2507,I801750,I801776,);
not I_47014 (I801784,I801776);
nand I_47015 (I801801,I298147,I298147);
and I_47016 (I801818,I801801,I298165);
DFFARX1 I_47017 (I801818,I2507,I801750,I801844,);
DFFARX1 I_47018 (I801844,I2507,I801750,I801739,);
DFFARX1 I_47019 (I298168,I2507,I801750,I801875,);
nand I_47020 (I801883,I801875,I298150);
not I_47021 (I801900,I801883);
DFFARX1 I_47022 (I801900,I2507,I801750,I801926,);
not I_47023 (I801934,I801926);
nor I_47024 (I801742,I801784,I801934);
DFFARX1 I_47025 (I298162,I2507,I801750,I801974,);
nor I_47026 (I801733,I801974,I801844);
nor I_47027 (I801724,I801974,I801900);
nand I_47028 (I802010,I298174,I298153);
and I_47029 (I802027,I802010,I298159);
DFFARX1 I_47030 (I802027,I2507,I801750,I802053,);
not I_47031 (I802061,I802053);
nand I_47032 (I802078,I802061,I801974);
nand I_47033 (I801727,I802061,I801883);
nor I_47034 (I802109,I298171,I298153);
and I_47035 (I802126,I801974,I802109);
nor I_47036 (I802143,I802061,I802126);
DFFARX1 I_47037 (I802143,I2507,I801750,I801736,);
nor I_47038 (I802174,I801776,I802109);
DFFARX1 I_47039 (I802174,I2507,I801750,I801721,);
nor I_47040 (I802205,I802053,I802109);
not I_47041 (I802222,I802205);
nand I_47042 (I801730,I802222,I802078);
not I_47043 (I802277,I2514);
DFFARX1 I_47044 (I389205,I2507,I802277,I802303,);
not I_47045 (I802311,I802303);
nand I_47046 (I802328,I389202,I389211);
and I_47047 (I802345,I802328,I389220);
DFFARX1 I_47048 (I802345,I2507,I802277,I802371,);
DFFARX1 I_47049 (I802371,I2507,I802277,I802266,);
DFFARX1 I_47050 (I389223,I2507,I802277,I802402,);
nand I_47051 (I802410,I802402,I389226);
not I_47052 (I802427,I802410);
DFFARX1 I_47053 (I802427,I2507,I802277,I802453,);
not I_47054 (I802461,I802453);
nor I_47055 (I802269,I802311,I802461);
DFFARX1 I_47056 (I389199,I2507,I802277,I802501,);
nor I_47057 (I802260,I802501,I802371);
nor I_47058 (I802251,I802501,I802427);
nand I_47059 (I802537,I389214,I389217);
and I_47060 (I802554,I802537,I389208);
DFFARX1 I_47061 (I802554,I2507,I802277,I802580,);
not I_47062 (I802588,I802580);
nand I_47063 (I802605,I802588,I802501);
nand I_47064 (I802254,I802588,I802410);
nor I_47065 (I802636,I389199,I389217);
and I_47066 (I802653,I802501,I802636);
nor I_47067 (I802670,I802588,I802653);
DFFARX1 I_47068 (I802670,I2507,I802277,I802263,);
nor I_47069 (I802701,I802303,I802636);
DFFARX1 I_47070 (I802701,I2507,I802277,I802248,);
nor I_47071 (I802732,I802580,I802636);
not I_47072 (I802749,I802732);
nand I_47073 (I802257,I802749,I802605);
not I_47074 (I802804,I2514);
DFFARX1 I_47075 (I409877,I2507,I802804,I802830,);
not I_47076 (I802838,I802830);
nand I_47077 (I802855,I409874,I409883);
and I_47078 (I802872,I802855,I409892);
DFFARX1 I_47079 (I802872,I2507,I802804,I802898,);
DFFARX1 I_47080 (I802898,I2507,I802804,I802793,);
DFFARX1 I_47081 (I409895,I2507,I802804,I802929,);
nand I_47082 (I802937,I802929,I409898);
not I_47083 (I802954,I802937);
DFFARX1 I_47084 (I802954,I2507,I802804,I802980,);
not I_47085 (I802988,I802980);
nor I_47086 (I802796,I802838,I802988);
DFFARX1 I_47087 (I409871,I2507,I802804,I803028,);
nor I_47088 (I802787,I803028,I802898);
nor I_47089 (I802778,I803028,I802954);
nand I_47090 (I803064,I409886,I409889);
and I_47091 (I803081,I803064,I409880);
DFFARX1 I_47092 (I803081,I2507,I802804,I803107,);
not I_47093 (I803115,I803107);
nand I_47094 (I803132,I803115,I803028);
nand I_47095 (I802781,I803115,I802937);
nor I_47096 (I803163,I409871,I409889);
and I_47097 (I803180,I803028,I803163);
nor I_47098 (I803197,I803115,I803180);
DFFARX1 I_47099 (I803197,I2507,I802804,I802790,);
nor I_47100 (I803228,I802830,I803163);
DFFARX1 I_47101 (I803228,I2507,I802804,I802775,);
nor I_47102 (I803259,I803107,I803163);
not I_47103 (I803276,I803259);
nand I_47104 (I802784,I803276,I803132);
not I_47105 (I803331,I2514);
DFFARX1 I_47106 (I278657,I2507,I803331,I803357,);
not I_47107 (I803365,I803357);
nand I_47108 (I803382,I278648,I278648);
and I_47109 (I803399,I803382,I278666);
DFFARX1 I_47110 (I803399,I2507,I803331,I803425,);
DFFARX1 I_47111 (I803425,I2507,I803331,I803320,);
DFFARX1 I_47112 (I278669,I2507,I803331,I803456,);
nand I_47113 (I803464,I803456,I278651);
not I_47114 (I803481,I803464);
DFFARX1 I_47115 (I803481,I2507,I803331,I803507,);
not I_47116 (I803515,I803507);
nor I_47117 (I803323,I803365,I803515);
DFFARX1 I_47118 (I278663,I2507,I803331,I803555,);
nor I_47119 (I803314,I803555,I803425);
nor I_47120 (I803305,I803555,I803481);
nand I_47121 (I803591,I278675,I278654);
and I_47122 (I803608,I803591,I278660);
DFFARX1 I_47123 (I803608,I2507,I803331,I803634,);
not I_47124 (I803642,I803634);
nand I_47125 (I803659,I803642,I803555);
nand I_47126 (I803308,I803642,I803464);
nor I_47127 (I803690,I278672,I278654);
and I_47128 (I803707,I803555,I803690);
nor I_47129 (I803724,I803642,I803707);
DFFARX1 I_47130 (I803724,I2507,I803331,I803317,);
nor I_47131 (I803755,I803357,I803690);
DFFARX1 I_47132 (I803755,I2507,I803331,I803302,);
nor I_47133 (I803786,I803634,I803690);
not I_47134 (I803803,I803786);
nand I_47135 (I803311,I803803,I803659);
not I_47136 (I803858,I2514);
DFFARX1 I_47137 (I754988,I2507,I803858,I803884,);
not I_47138 (I803892,I803884);
nand I_47139 (I803909,I754991,I754988);
and I_47140 (I803926,I803909,I755000);
DFFARX1 I_47141 (I803926,I2507,I803858,I803952,);
DFFARX1 I_47142 (I803952,I2507,I803858,I803847,);
DFFARX1 I_47143 (I754997,I2507,I803858,I803983,);
nand I_47144 (I803991,I803983,I755003);
not I_47145 (I804008,I803991);
DFFARX1 I_47146 (I804008,I2507,I803858,I804034,);
not I_47147 (I804042,I804034);
nor I_47148 (I803850,I803892,I804042);
DFFARX1 I_47149 (I755012,I2507,I803858,I804082,);
nor I_47150 (I803841,I804082,I803952);
nor I_47151 (I803832,I804082,I804008);
nand I_47152 (I804118,I755006,I754994);
and I_47153 (I804135,I804118,I754991);
DFFARX1 I_47154 (I804135,I2507,I803858,I804161,);
not I_47155 (I804169,I804161);
nand I_47156 (I804186,I804169,I804082);
nand I_47157 (I803835,I804169,I803991);
nor I_47158 (I804217,I755009,I754994);
and I_47159 (I804234,I804082,I804217);
nor I_47160 (I804251,I804169,I804234);
DFFARX1 I_47161 (I804251,I2507,I803858,I803844,);
nor I_47162 (I804282,I803884,I804217);
DFFARX1 I_47163 (I804282,I2507,I803858,I803829,);
nor I_47164 (I804313,I804161,I804217);
not I_47165 (I804330,I804313);
nand I_47166 (I803838,I804330,I804186);
not I_47167 (I804385,I2514);
DFFARX1 I_47168 (I1279048,I2507,I804385,I804411,);
not I_47169 (I804419,I804411);
nand I_47170 (I804436,I1279030,I1279033);
and I_47171 (I804453,I804436,I1279045);
DFFARX1 I_47172 (I804453,I2507,I804385,I804479,);
DFFARX1 I_47173 (I804479,I2507,I804385,I804374,);
DFFARX1 I_47174 (I1279054,I2507,I804385,I804510,);
nand I_47175 (I804518,I804510,I1279039);
not I_47176 (I804535,I804518);
DFFARX1 I_47177 (I804535,I2507,I804385,I804561,);
not I_47178 (I804569,I804561);
nor I_47179 (I804377,I804419,I804569);
DFFARX1 I_47180 (I1279051,I2507,I804385,I804609,);
nor I_47181 (I804368,I804609,I804479);
nor I_47182 (I804359,I804609,I804535);
nand I_47183 (I804645,I1279042,I1279036);
and I_47184 (I804662,I804645,I1279030);
DFFARX1 I_47185 (I804662,I2507,I804385,I804688,);
not I_47186 (I804696,I804688);
nand I_47187 (I804713,I804696,I804609);
nand I_47188 (I804362,I804696,I804518);
nor I_47189 (I804744,I1279033,I1279036);
and I_47190 (I804761,I804609,I804744);
nor I_47191 (I804778,I804696,I804761);
DFFARX1 I_47192 (I804778,I2507,I804385,I804371,);
nor I_47193 (I804809,I804411,I804744);
DFFARX1 I_47194 (I804809,I2507,I804385,I804356,);
nor I_47195 (I804840,I804688,I804744);
not I_47196 (I804857,I804840);
nand I_47197 (I804365,I804857,I804713);
not I_47198 (I804912,I2514);
DFFARX1 I_47199 (I1272690,I2507,I804912,I804938,);
not I_47200 (I804946,I804938);
nand I_47201 (I804963,I1272672,I1272675);
and I_47202 (I804980,I804963,I1272687);
DFFARX1 I_47203 (I804980,I2507,I804912,I805006,);
DFFARX1 I_47204 (I805006,I2507,I804912,I804901,);
DFFARX1 I_47205 (I1272696,I2507,I804912,I805037,);
nand I_47206 (I805045,I805037,I1272681);
not I_47207 (I805062,I805045);
DFFARX1 I_47208 (I805062,I2507,I804912,I805088,);
not I_47209 (I805096,I805088);
nor I_47210 (I804904,I804946,I805096);
DFFARX1 I_47211 (I1272693,I2507,I804912,I805136,);
nor I_47212 (I804895,I805136,I805006);
nor I_47213 (I804886,I805136,I805062);
nand I_47214 (I805172,I1272684,I1272678);
and I_47215 (I805189,I805172,I1272672);
DFFARX1 I_47216 (I805189,I2507,I804912,I805215,);
not I_47217 (I805223,I805215);
nand I_47218 (I805240,I805223,I805136);
nand I_47219 (I804889,I805223,I805045);
nor I_47220 (I805271,I1272675,I1272678);
and I_47221 (I805288,I805136,I805271);
nor I_47222 (I805305,I805223,I805288);
DFFARX1 I_47223 (I805305,I2507,I804912,I804898,);
nor I_47224 (I805336,I804938,I805271);
DFFARX1 I_47225 (I805336,I2507,I804912,I804883,);
nor I_47226 (I805367,I805215,I805271);
not I_47227 (I805384,I805367);
nand I_47228 (I804892,I805384,I805240);
not I_47229 (I805439,I2514);
DFFARX1 I_47230 (I641700,I2507,I805439,I805465,);
not I_47231 (I805473,I805465);
nand I_47232 (I805490,I641703,I641700);
and I_47233 (I805507,I805490,I641712);
DFFARX1 I_47234 (I805507,I2507,I805439,I805533,);
DFFARX1 I_47235 (I805533,I2507,I805439,I805428,);
DFFARX1 I_47236 (I641709,I2507,I805439,I805564,);
nand I_47237 (I805572,I805564,I641715);
not I_47238 (I805589,I805572);
DFFARX1 I_47239 (I805589,I2507,I805439,I805615,);
not I_47240 (I805623,I805615);
nor I_47241 (I805431,I805473,I805623);
DFFARX1 I_47242 (I641724,I2507,I805439,I805663,);
nor I_47243 (I805422,I805663,I805533);
nor I_47244 (I805413,I805663,I805589);
nand I_47245 (I805699,I641718,I641706);
and I_47246 (I805716,I805699,I641703);
DFFARX1 I_47247 (I805716,I2507,I805439,I805742,);
not I_47248 (I805750,I805742);
nand I_47249 (I805767,I805750,I805663);
nand I_47250 (I805416,I805750,I805572);
nor I_47251 (I805798,I641721,I641706);
and I_47252 (I805815,I805663,I805798);
nor I_47253 (I805832,I805750,I805815);
DFFARX1 I_47254 (I805832,I2507,I805439,I805425,);
nor I_47255 (I805863,I805465,I805798);
DFFARX1 I_47256 (I805863,I2507,I805439,I805410,);
nor I_47257 (I805894,I805742,I805798);
not I_47258 (I805911,I805894);
nand I_47259 (I805419,I805911,I805767);
not I_47260 (I805966,I2514);
DFFARX1 I_47261 (I79653,I2507,I805966,I805992,);
not I_47262 (I806000,I805992);
nand I_47263 (I806017,I79629,I79638);
and I_47264 (I806034,I806017,I79632);
DFFARX1 I_47265 (I806034,I2507,I805966,I806060,);
DFFARX1 I_47266 (I806060,I2507,I805966,I805955,);
DFFARX1 I_47267 (I79650,I2507,I805966,I806091,);
nand I_47268 (I806099,I806091,I79641);
not I_47269 (I806116,I806099);
DFFARX1 I_47270 (I806116,I2507,I805966,I806142,);
not I_47271 (I806150,I806142);
nor I_47272 (I805958,I806000,I806150);
DFFARX1 I_47273 (I79635,I2507,I805966,I806190,);
nor I_47274 (I805949,I806190,I806060);
nor I_47275 (I805940,I806190,I806116);
nand I_47276 (I806226,I79647,I79644);
and I_47277 (I806243,I806226,I79632);
DFFARX1 I_47278 (I806243,I2507,I805966,I806269,);
not I_47279 (I806277,I806269);
nand I_47280 (I806294,I806277,I806190);
nand I_47281 (I805943,I806277,I806099);
nor I_47282 (I806325,I79629,I79644);
and I_47283 (I806342,I806190,I806325);
nor I_47284 (I806359,I806277,I806342);
DFFARX1 I_47285 (I806359,I2507,I805966,I805952,);
nor I_47286 (I806390,I805992,I806325);
DFFARX1 I_47287 (I806390,I2507,I805966,I805937,);
nor I_47288 (I806421,I806269,I806325);
not I_47289 (I806438,I806421);
nand I_47290 (I805946,I806438,I806294);
not I_47291 (I806493,I2514);
DFFARX1 I_47292 (I344005,I2507,I806493,I806519,);
not I_47293 (I806527,I806519);
nand I_47294 (I806544,I343996,I343996);
and I_47295 (I806561,I806544,I344014);
DFFARX1 I_47296 (I806561,I2507,I806493,I806587,);
DFFARX1 I_47297 (I806587,I2507,I806493,I806482,);
DFFARX1 I_47298 (I344017,I2507,I806493,I806618,);
nand I_47299 (I806626,I806618,I343999);
not I_47300 (I806643,I806626);
DFFARX1 I_47301 (I806643,I2507,I806493,I806669,);
not I_47302 (I806677,I806669);
nor I_47303 (I806485,I806527,I806677);
DFFARX1 I_47304 (I344011,I2507,I806493,I806717,);
nor I_47305 (I806476,I806717,I806587);
nor I_47306 (I806467,I806717,I806643);
nand I_47307 (I806753,I344023,I344002);
and I_47308 (I806770,I806753,I344008);
DFFARX1 I_47309 (I806770,I2507,I806493,I806796,);
not I_47310 (I806804,I806796);
nand I_47311 (I806821,I806804,I806717);
nand I_47312 (I806470,I806804,I806626);
nor I_47313 (I806852,I344020,I344002);
and I_47314 (I806869,I806717,I806852);
nor I_47315 (I806886,I806804,I806869);
DFFARX1 I_47316 (I806886,I2507,I806493,I806479,);
nor I_47317 (I806917,I806519,I806852);
DFFARX1 I_47318 (I806917,I2507,I806493,I806464,);
nor I_47319 (I806948,I806796,I806852);
not I_47320 (I806965,I806948);
nand I_47321 (I806473,I806965,I806821);
not I_47322 (I807020,I2514);
DFFARX1 I_47323 (I145494,I2507,I807020,I807046,);
not I_47324 (I807054,I807046);
nand I_47325 (I807071,I145470,I145488);
and I_47326 (I807088,I807071,I145476);
DFFARX1 I_47327 (I807088,I2507,I807020,I807114,);
DFFARX1 I_47328 (I807114,I2507,I807020,I807009,);
DFFARX1 I_47329 (I145485,I2507,I807020,I807145,);
nand I_47330 (I807153,I807145,I145491);
not I_47331 (I807170,I807153);
DFFARX1 I_47332 (I807170,I2507,I807020,I807196,);
not I_47333 (I807204,I807196);
nor I_47334 (I807012,I807054,I807204);
DFFARX1 I_47335 (I145470,I2507,I807020,I807244,);
nor I_47336 (I807003,I807244,I807114);
nor I_47337 (I806994,I807244,I807170);
nand I_47338 (I807280,I145482,I145473);
and I_47339 (I807297,I807280,I145497);
DFFARX1 I_47340 (I807297,I2507,I807020,I807323,);
not I_47341 (I807331,I807323);
nand I_47342 (I807348,I807331,I807244);
nand I_47343 (I806997,I807331,I807153);
nor I_47344 (I807379,I145479,I145473);
and I_47345 (I807396,I807244,I807379);
nor I_47346 (I807413,I807331,I807396);
DFFARX1 I_47347 (I807413,I2507,I807020,I807006,);
nor I_47348 (I807444,I807046,I807379);
DFFARX1 I_47349 (I807444,I2507,I807020,I806991,);
nor I_47350 (I807475,I807323,I807379);
not I_47351 (I807492,I807475);
nand I_47352 (I807000,I807492,I807348);
not I_47353 (I807547,I2514);
DFFARX1 I_47354 (I1339242,I2507,I807547,I807573,);
not I_47355 (I807581,I807573);
nand I_47356 (I807598,I1339239,I1339248);
and I_47357 (I807615,I807598,I1339227);
DFFARX1 I_47358 (I807615,I2507,I807547,I807641,);
DFFARX1 I_47359 (I807641,I2507,I807547,I807536,);
DFFARX1 I_47360 (I1339230,I2507,I807547,I807672,);
nand I_47361 (I807680,I807672,I1339245);
not I_47362 (I807697,I807680);
DFFARX1 I_47363 (I807697,I2507,I807547,I807723,);
not I_47364 (I807731,I807723);
nor I_47365 (I807539,I807581,I807731);
DFFARX1 I_47366 (I1339251,I2507,I807547,I807771,);
nor I_47367 (I807530,I807771,I807641);
nor I_47368 (I807521,I807771,I807697);
nand I_47369 (I807807,I1339233,I1339254);
and I_47370 (I807824,I807807,I1339236);
DFFARX1 I_47371 (I807824,I2507,I807547,I807850,);
not I_47372 (I807858,I807850);
nand I_47373 (I807875,I807858,I807771);
nand I_47374 (I807524,I807858,I807680);
nor I_47375 (I807906,I1339227,I1339254);
and I_47376 (I807923,I807771,I807906);
nor I_47377 (I807940,I807858,I807923);
DFFARX1 I_47378 (I807940,I2507,I807547,I807533,);
nor I_47379 (I807971,I807573,I807906);
DFFARX1 I_47380 (I807971,I2507,I807547,I807518,);
nor I_47381 (I808002,I807850,I807906);
not I_47382 (I808019,I808002);
nand I_47383 (I807527,I808019,I807875);
not I_47384 (I808074,I2514);
DFFARX1 I_47385 (I267590,I2507,I808074,I808100,);
not I_47386 (I808108,I808100);
nand I_47387 (I808125,I267581,I267581);
and I_47388 (I808142,I808125,I267599);
DFFARX1 I_47389 (I808142,I2507,I808074,I808168,);
DFFARX1 I_47390 (I808168,I2507,I808074,I808063,);
DFFARX1 I_47391 (I267602,I2507,I808074,I808199,);
nand I_47392 (I808207,I808199,I267584);
not I_47393 (I808224,I808207);
DFFARX1 I_47394 (I808224,I2507,I808074,I808250,);
not I_47395 (I808258,I808250);
nor I_47396 (I808066,I808108,I808258);
DFFARX1 I_47397 (I267596,I2507,I808074,I808298,);
nor I_47398 (I808057,I808298,I808168);
nor I_47399 (I808048,I808298,I808224);
nand I_47400 (I808334,I267608,I267587);
and I_47401 (I808351,I808334,I267593);
DFFARX1 I_47402 (I808351,I2507,I808074,I808377,);
not I_47403 (I808385,I808377);
nand I_47404 (I808402,I808385,I808298);
nand I_47405 (I808051,I808385,I808207);
nor I_47406 (I808433,I267605,I267587);
and I_47407 (I808450,I808298,I808433);
nor I_47408 (I808467,I808385,I808450);
DFFARX1 I_47409 (I808467,I2507,I808074,I808060,);
nor I_47410 (I808498,I808100,I808433);
DFFARX1 I_47411 (I808498,I2507,I808074,I808045,);
nor I_47412 (I808529,I808377,I808433);
not I_47413 (I808546,I808529);
nand I_47414 (I808054,I808546,I808402);
not I_47415 (I808601,I2514);
DFFARX1 I_47416 (I1127170,I2507,I808601,I808627,);
not I_47417 (I808635,I808627);
nand I_47418 (I808652,I1127152,I1127152);
and I_47419 (I808669,I808652,I1127158);
DFFARX1 I_47420 (I808669,I2507,I808601,I808695,);
DFFARX1 I_47421 (I808695,I2507,I808601,I808590,);
DFFARX1 I_47422 (I1127155,I2507,I808601,I808726,);
nand I_47423 (I808734,I808726,I1127164);
not I_47424 (I808751,I808734);
DFFARX1 I_47425 (I808751,I2507,I808601,I808777,);
not I_47426 (I808785,I808777);
nor I_47427 (I808593,I808635,I808785);
DFFARX1 I_47428 (I1127176,I2507,I808601,I808825,);
nor I_47429 (I808584,I808825,I808695);
nor I_47430 (I808575,I808825,I808751);
nand I_47431 (I808861,I1127167,I1127161);
and I_47432 (I808878,I808861,I1127155);
DFFARX1 I_47433 (I808878,I2507,I808601,I808904,);
not I_47434 (I808912,I808904);
nand I_47435 (I808929,I808912,I808825);
nand I_47436 (I808578,I808912,I808734);
nor I_47437 (I808960,I1127173,I1127161);
and I_47438 (I808977,I808825,I808960);
nor I_47439 (I808994,I808912,I808977);
DFFARX1 I_47440 (I808994,I2507,I808601,I808587,);
nor I_47441 (I809025,I808627,I808960);
DFFARX1 I_47442 (I809025,I2507,I808601,I808572,);
nor I_47443 (I809056,I808904,I808960);
not I_47444 (I809073,I809056);
nand I_47445 (I808581,I809073,I808929);
not I_47446 (I809128,I2514);
DFFARX1 I_47447 (I716840,I2507,I809128,I809154,);
not I_47448 (I809162,I809154);
nand I_47449 (I809179,I716843,I716840);
and I_47450 (I809196,I809179,I716852);
DFFARX1 I_47451 (I809196,I2507,I809128,I809222,);
DFFARX1 I_47452 (I809222,I2507,I809128,I809117,);
DFFARX1 I_47453 (I716849,I2507,I809128,I809253,);
nand I_47454 (I809261,I809253,I716855);
not I_47455 (I809278,I809261);
DFFARX1 I_47456 (I809278,I2507,I809128,I809304,);
not I_47457 (I809312,I809304);
nor I_47458 (I809120,I809162,I809312);
DFFARX1 I_47459 (I716864,I2507,I809128,I809352,);
nor I_47460 (I809111,I809352,I809222);
nor I_47461 (I809102,I809352,I809278);
nand I_47462 (I809388,I716858,I716846);
and I_47463 (I809405,I809388,I716843);
DFFARX1 I_47464 (I809405,I2507,I809128,I809431,);
not I_47465 (I809439,I809431);
nand I_47466 (I809456,I809439,I809352);
nand I_47467 (I809105,I809439,I809261);
nor I_47468 (I809487,I716861,I716846);
and I_47469 (I809504,I809352,I809487);
nor I_47470 (I809521,I809439,I809504);
DFFARX1 I_47471 (I809521,I2507,I809128,I809114,);
nor I_47472 (I809552,I809154,I809487);
DFFARX1 I_47473 (I809552,I2507,I809128,I809099,);
nor I_47474 (I809583,I809431,I809487);
not I_47475 (I809600,I809583);
nand I_47476 (I809108,I809600,I809456);
not I_47477 (I809655,I2514);
DFFARX1 I_47478 (I568309,I2507,I809655,I809681,);
not I_47479 (I809689,I809681);
nand I_47480 (I809706,I568294,I568315);
and I_47481 (I809723,I809706,I568303);
DFFARX1 I_47482 (I809723,I2507,I809655,I809749,);
DFFARX1 I_47483 (I809749,I2507,I809655,I809644,);
DFFARX1 I_47484 (I568297,I2507,I809655,I809780,);
nand I_47485 (I809788,I809780,I568306);
not I_47486 (I809805,I809788);
DFFARX1 I_47487 (I809805,I2507,I809655,I809831,);
not I_47488 (I809839,I809831);
nor I_47489 (I809647,I809689,I809839);
DFFARX1 I_47490 (I568312,I2507,I809655,I809879,);
nor I_47491 (I809638,I809879,I809749);
nor I_47492 (I809629,I809879,I809805);
nand I_47493 (I809915,I568294,I568297);
and I_47494 (I809932,I809915,I568318);
DFFARX1 I_47495 (I809932,I2507,I809655,I809958,);
not I_47496 (I809966,I809958);
nand I_47497 (I809983,I809966,I809879);
nand I_47498 (I809632,I809966,I809788);
nor I_47499 (I810014,I568300,I568297);
and I_47500 (I810031,I809879,I810014);
nor I_47501 (I810048,I809966,I810031);
DFFARX1 I_47502 (I810048,I2507,I809655,I809641,);
nor I_47503 (I810079,I809681,I810014);
DFFARX1 I_47504 (I810079,I2507,I809655,I809626,);
nor I_47505 (I810110,I809958,I810014);
not I_47506 (I810127,I810110);
nand I_47507 (I809635,I810127,I809983);
not I_47508 (I810182,I2514);
DFFARX1 I_47509 (I556749,I2507,I810182,I810208,);
not I_47510 (I810216,I810208);
nand I_47511 (I810233,I556734,I556755);
and I_47512 (I810250,I810233,I556743);
DFFARX1 I_47513 (I810250,I2507,I810182,I810276,);
DFFARX1 I_47514 (I810276,I2507,I810182,I810171,);
DFFARX1 I_47515 (I556737,I2507,I810182,I810307,);
nand I_47516 (I810315,I810307,I556746);
not I_47517 (I810332,I810315);
DFFARX1 I_47518 (I810332,I2507,I810182,I810358,);
not I_47519 (I810366,I810358);
nor I_47520 (I810174,I810216,I810366);
DFFARX1 I_47521 (I556752,I2507,I810182,I810406,);
nor I_47522 (I810165,I810406,I810276);
nor I_47523 (I810156,I810406,I810332);
nand I_47524 (I810442,I556734,I556737);
and I_47525 (I810459,I810442,I556758);
DFFARX1 I_47526 (I810459,I2507,I810182,I810485,);
not I_47527 (I810493,I810485);
nand I_47528 (I810510,I810493,I810406);
nand I_47529 (I810159,I810493,I810315);
nor I_47530 (I810541,I556740,I556737);
and I_47531 (I810558,I810406,I810541);
nor I_47532 (I810575,I810493,I810558);
DFFARX1 I_47533 (I810575,I2507,I810182,I810168,);
nor I_47534 (I810606,I810208,I810541);
DFFARX1 I_47535 (I810606,I2507,I810182,I810153,);
nor I_47536 (I810637,I810485,I810541);
not I_47537 (I810654,I810637);
nand I_47538 (I810162,I810654,I810510);
not I_47539 (I810709,I2514);
DFFARX1 I_47540 (I77545,I2507,I810709,I810735,);
not I_47541 (I810743,I810735);
nand I_47542 (I810760,I77521,I77530);
and I_47543 (I810777,I810760,I77524);
DFFARX1 I_47544 (I810777,I2507,I810709,I810803,);
DFFARX1 I_47545 (I810803,I2507,I810709,I810698,);
DFFARX1 I_47546 (I77542,I2507,I810709,I810834,);
nand I_47547 (I810842,I810834,I77533);
not I_47548 (I810859,I810842);
DFFARX1 I_47549 (I810859,I2507,I810709,I810885,);
not I_47550 (I810893,I810885);
nor I_47551 (I810701,I810743,I810893);
DFFARX1 I_47552 (I77527,I2507,I810709,I810933,);
nor I_47553 (I810692,I810933,I810803);
nor I_47554 (I810683,I810933,I810859);
nand I_47555 (I810969,I77539,I77536);
and I_47556 (I810986,I810969,I77524);
DFFARX1 I_47557 (I810986,I2507,I810709,I811012,);
not I_47558 (I811020,I811012);
nand I_47559 (I811037,I811020,I810933);
nand I_47560 (I810686,I811020,I810842);
nor I_47561 (I811068,I77521,I77536);
and I_47562 (I811085,I810933,I811068);
nor I_47563 (I811102,I811020,I811085);
DFFARX1 I_47564 (I811102,I2507,I810709,I810695,);
nor I_47565 (I811133,I810735,I811068);
DFFARX1 I_47566 (I811133,I2507,I810709,I810680,);
nor I_47567 (I811164,I811012,I811068);
not I_47568 (I811181,I811164);
nand I_47569 (I810689,I811181,I811037);
not I_47570 (I811236,I2514);
DFFARX1 I_47571 (I644012,I2507,I811236,I811262,);
not I_47572 (I811270,I811262);
nand I_47573 (I811287,I644015,I644012);
and I_47574 (I811304,I811287,I644024);
DFFARX1 I_47575 (I811304,I2507,I811236,I811330,);
DFFARX1 I_47576 (I811330,I2507,I811236,I811225,);
DFFARX1 I_47577 (I644021,I2507,I811236,I811361,);
nand I_47578 (I811369,I811361,I644027);
not I_47579 (I811386,I811369);
DFFARX1 I_47580 (I811386,I2507,I811236,I811412,);
not I_47581 (I811420,I811412);
nor I_47582 (I811228,I811270,I811420);
DFFARX1 I_47583 (I644036,I2507,I811236,I811460,);
nor I_47584 (I811219,I811460,I811330);
nor I_47585 (I811210,I811460,I811386);
nand I_47586 (I811496,I644030,I644018);
and I_47587 (I811513,I811496,I644015);
DFFARX1 I_47588 (I811513,I2507,I811236,I811539,);
not I_47589 (I811547,I811539);
nand I_47590 (I811564,I811547,I811460);
nand I_47591 (I811213,I811547,I811369);
nor I_47592 (I811595,I644033,I644018);
and I_47593 (I811612,I811460,I811595);
nor I_47594 (I811629,I811547,I811612);
DFFARX1 I_47595 (I811629,I2507,I811236,I811222,);
nor I_47596 (I811660,I811262,I811595);
DFFARX1 I_47597 (I811660,I2507,I811236,I811207,);
nor I_47598 (I811691,I811539,I811595);
not I_47599 (I811708,I811691);
nand I_47600 (I811216,I811708,I811564);
not I_47601 (I811763,I2514);
DFFARX1 I_47602 (I600099,I2507,I811763,I811789,);
not I_47603 (I811797,I811789);
nand I_47604 (I811814,I600084,I600105);
and I_47605 (I811831,I811814,I600093);
DFFARX1 I_47606 (I811831,I2507,I811763,I811857,);
DFFARX1 I_47607 (I811857,I2507,I811763,I811752,);
DFFARX1 I_47608 (I600087,I2507,I811763,I811888,);
nand I_47609 (I811896,I811888,I600096);
not I_47610 (I811913,I811896);
DFFARX1 I_47611 (I811913,I2507,I811763,I811939,);
not I_47612 (I811947,I811939);
nor I_47613 (I811755,I811797,I811947);
DFFARX1 I_47614 (I600102,I2507,I811763,I811987,);
nor I_47615 (I811746,I811987,I811857);
nor I_47616 (I811737,I811987,I811913);
nand I_47617 (I812023,I600084,I600087);
and I_47618 (I812040,I812023,I600108);
DFFARX1 I_47619 (I812040,I2507,I811763,I812066,);
not I_47620 (I812074,I812066);
nand I_47621 (I812091,I812074,I811987);
nand I_47622 (I811740,I812074,I811896);
nor I_47623 (I812122,I600090,I600087);
and I_47624 (I812139,I811987,I812122);
nor I_47625 (I812156,I812074,I812139);
DFFARX1 I_47626 (I812156,I2507,I811763,I811749,);
nor I_47627 (I812187,I811789,I812122);
DFFARX1 I_47628 (I812187,I2507,I811763,I811734,);
nor I_47629 (I812218,I812066,I812122);
not I_47630 (I812235,I812218);
nand I_47631 (I811743,I812235,I812091);
not I_47632 (I812290,I2514);
DFFARX1 I_47633 (I1112142,I2507,I812290,I812316,);
not I_47634 (I812324,I812316);
nand I_47635 (I812341,I1112124,I1112124);
and I_47636 (I812358,I812341,I1112130);
DFFARX1 I_47637 (I812358,I2507,I812290,I812384,);
DFFARX1 I_47638 (I812384,I2507,I812290,I812279,);
DFFARX1 I_47639 (I1112127,I2507,I812290,I812415,);
nand I_47640 (I812423,I812415,I1112136);
not I_47641 (I812440,I812423);
DFFARX1 I_47642 (I812440,I2507,I812290,I812466,);
not I_47643 (I812474,I812466);
nor I_47644 (I812282,I812324,I812474);
DFFARX1 I_47645 (I1112148,I2507,I812290,I812514,);
nor I_47646 (I812273,I812514,I812384);
nor I_47647 (I812264,I812514,I812440);
nand I_47648 (I812550,I1112139,I1112133);
and I_47649 (I812567,I812550,I1112127);
DFFARX1 I_47650 (I812567,I2507,I812290,I812593,);
not I_47651 (I812601,I812593);
nand I_47652 (I812618,I812601,I812514);
nand I_47653 (I812267,I812601,I812423);
nor I_47654 (I812649,I1112145,I1112133);
and I_47655 (I812666,I812514,I812649);
nor I_47656 (I812683,I812601,I812666);
DFFARX1 I_47657 (I812683,I2507,I812290,I812276,);
nor I_47658 (I812714,I812316,I812649);
DFFARX1 I_47659 (I812714,I2507,I812290,I812261,);
nor I_47660 (I812745,I812593,I812649);
not I_47661 (I812762,I812745);
nand I_47662 (I812270,I812762,I812618);
not I_47663 (I812817,I2514);
DFFARX1 I_47664 (I520275,I2507,I812817,I812843,);
not I_47665 (I812851,I812843);
nand I_47666 (I812868,I520293,I520284);
and I_47667 (I812885,I812868,I520287);
DFFARX1 I_47668 (I812885,I2507,I812817,I812911,);
DFFARX1 I_47669 (I812911,I2507,I812817,I812806,);
DFFARX1 I_47670 (I520281,I2507,I812817,I812942,);
nand I_47671 (I812950,I812942,I520272);
not I_47672 (I812967,I812950);
DFFARX1 I_47673 (I812967,I2507,I812817,I812993,);
not I_47674 (I813001,I812993);
nor I_47675 (I812809,I812851,I813001);
DFFARX1 I_47676 (I520278,I2507,I812817,I813041,);
nor I_47677 (I812800,I813041,I812911);
nor I_47678 (I812791,I813041,I812967);
nand I_47679 (I813077,I520272,I520269);
and I_47680 (I813094,I813077,I520290);
DFFARX1 I_47681 (I813094,I2507,I812817,I813120,);
not I_47682 (I813128,I813120);
nand I_47683 (I813145,I813128,I813041);
nand I_47684 (I812794,I813128,I812950);
nor I_47685 (I813176,I520269,I520269);
and I_47686 (I813193,I813041,I813176);
nor I_47687 (I813210,I813128,I813193);
DFFARX1 I_47688 (I813210,I2507,I812817,I812803,);
nor I_47689 (I813241,I812843,I813176);
DFFARX1 I_47690 (I813241,I2507,I812817,I812788,);
nor I_47691 (I813272,I813120,I813176);
not I_47692 (I813289,I813272);
nand I_47693 (I812797,I813289,I813145);
not I_47694 (I813344,I2514);
DFFARX1 I_47695 (I729556,I2507,I813344,I813370,);
not I_47696 (I813378,I813370);
nand I_47697 (I813395,I729559,I729556);
and I_47698 (I813412,I813395,I729568);
DFFARX1 I_47699 (I813412,I2507,I813344,I813438,);
DFFARX1 I_47700 (I813438,I2507,I813344,I813333,);
DFFARX1 I_47701 (I729565,I2507,I813344,I813469,);
nand I_47702 (I813477,I813469,I729571);
not I_47703 (I813494,I813477);
DFFARX1 I_47704 (I813494,I2507,I813344,I813520,);
not I_47705 (I813528,I813520);
nor I_47706 (I813336,I813378,I813528);
DFFARX1 I_47707 (I729580,I2507,I813344,I813568,);
nor I_47708 (I813327,I813568,I813438);
nor I_47709 (I813318,I813568,I813494);
nand I_47710 (I813604,I729574,I729562);
and I_47711 (I813621,I813604,I729559);
DFFARX1 I_47712 (I813621,I2507,I813344,I813647,);
not I_47713 (I813655,I813647);
nand I_47714 (I813672,I813655,I813568);
nand I_47715 (I813321,I813655,I813477);
nor I_47716 (I813703,I729577,I729562);
and I_47717 (I813720,I813568,I813703);
nor I_47718 (I813737,I813655,I813720);
DFFARX1 I_47719 (I813737,I2507,I813344,I813330,);
nor I_47720 (I813768,I813370,I813703);
DFFARX1 I_47721 (I813768,I2507,I813344,I813315,);
nor I_47722 (I813799,I813647,I813703);
not I_47723 (I813816,I813799);
nand I_47724 (I813324,I813816,I813672);
not I_47725 (I813871,I2514);
DFFARX1 I_47726 (I1160116,I2507,I813871,I813897,);
not I_47727 (I813905,I813897);
nand I_47728 (I813922,I1160098,I1160098);
and I_47729 (I813939,I813922,I1160104);
DFFARX1 I_47730 (I813939,I2507,I813871,I813965,);
DFFARX1 I_47731 (I813965,I2507,I813871,I813860,);
DFFARX1 I_47732 (I1160101,I2507,I813871,I813996,);
nand I_47733 (I814004,I813996,I1160110);
not I_47734 (I814021,I814004);
DFFARX1 I_47735 (I814021,I2507,I813871,I814047,);
not I_47736 (I814055,I814047);
nor I_47737 (I813863,I813905,I814055);
DFFARX1 I_47738 (I1160122,I2507,I813871,I814095,);
nor I_47739 (I813854,I814095,I813965);
nor I_47740 (I813845,I814095,I814021);
nand I_47741 (I814131,I1160113,I1160107);
and I_47742 (I814148,I814131,I1160101);
DFFARX1 I_47743 (I814148,I2507,I813871,I814174,);
not I_47744 (I814182,I814174);
nand I_47745 (I814199,I814182,I814095);
nand I_47746 (I813848,I814182,I814004);
nor I_47747 (I814230,I1160119,I1160107);
and I_47748 (I814247,I814095,I814230);
nor I_47749 (I814264,I814182,I814247);
DFFARX1 I_47750 (I814264,I2507,I813871,I813857,);
nor I_47751 (I814295,I813897,I814230);
DFFARX1 I_47752 (I814295,I2507,I813871,I813842,);
nor I_47753 (I814326,I814174,I814230);
not I_47754 (I814343,I814326);
nand I_47755 (I813851,I814343,I814199);
not I_47756 (I814398,I2514);
DFFARX1 I_47757 (I490389,I2507,I814398,I814424,);
not I_47758 (I814432,I814424);
nand I_47759 (I814449,I490386,I490395);
and I_47760 (I814466,I814449,I490404);
DFFARX1 I_47761 (I814466,I2507,I814398,I814492,);
DFFARX1 I_47762 (I814492,I2507,I814398,I814387,);
DFFARX1 I_47763 (I490407,I2507,I814398,I814523,);
nand I_47764 (I814531,I814523,I490410);
not I_47765 (I814548,I814531);
DFFARX1 I_47766 (I814548,I2507,I814398,I814574,);
not I_47767 (I814582,I814574);
nor I_47768 (I814390,I814432,I814582);
DFFARX1 I_47769 (I490383,I2507,I814398,I814622,);
nor I_47770 (I814381,I814622,I814492);
nor I_47771 (I814372,I814622,I814548);
nand I_47772 (I814658,I490398,I490401);
and I_47773 (I814675,I814658,I490392);
DFFARX1 I_47774 (I814675,I2507,I814398,I814701,);
not I_47775 (I814709,I814701);
nand I_47776 (I814726,I814709,I814622);
nand I_47777 (I814375,I814709,I814531);
nor I_47778 (I814757,I490383,I490401);
and I_47779 (I814774,I814622,I814757);
nor I_47780 (I814791,I814709,I814774);
DFFARX1 I_47781 (I814791,I2507,I814398,I814384,);
nor I_47782 (I814822,I814424,I814757);
DFFARX1 I_47783 (I814822,I2507,I814398,I814369,);
nor I_47784 (I814853,I814701,I814757);
not I_47785 (I814870,I814853);
nand I_47786 (I814378,I814870,I814726);
not I_47787 (I814925,I2514);
DFFARX1 I_47788 (I1100004,I2507,I814925,I814951,);
not I_47789 (I814959,I814951);
nand I_47790 (I814976,I1099986,I1099986);
and I_47791 (I814993,I814976,I1099992);
DFFARX1 I_47792 (I814993,I2507,I814925,I815019,);
DFFARX1 I_47793 (I815019,I2507,I814925,I814914,);
DFFARX1 I_47794 (I1099989,I2507,I814925,I815050,);
nand I_47795 (I815058,I815050,I1099998);
not I_47796 (I815075,I815058);
DFFARX1 I_47797 (I815075,I2507,I814925,I815101,);
not I_47798 (I815109,I815101);
nor I_47799 (I814917,I814959,I815109);
DFFARX1 I_47800 (I1100010,I2507,I814925,I815149,);
nor I_47801 (I814908,I815149,I815019);
nor I_47802 (I814899,I815149,I815075);
nand I_47803 (I815185,I1100001,I1099995);
and I_47804 (I815202,I815185,I1099989);
DFFARX1 I_47805 (I815202,I2507,I814925,I815228,);
not I_47806 (I815236,I815228);
nand I_47807 (I815253,I815236,I815149);
nand I_47808 (I814902,I815236,I815058);
nor I_47809 (I815284,I1100007,I1099995);
and I_47810 (I815301,I815149,I815284);
nor I_47811 (I815318,I815236,I815301);
DFFARX1 I_47812 (I815318,I2507,I814925,I814911,);
nor I_47813 (I815349,I814951,I815284);
DFFARX1 I_47814 (I815349,I2507,I814925,I814896,);
nor I_47815 (I815380,I815228,I815284);
not I_47816 (I815397,I815380);
nand I_47817 (I814905,I815397,I815253);
not I_47818 (I815452,I2514);
DFFARX1 I_47819 (I72275,I2507,I815452,I815478,);
not I_47820 (I815486,I815478);
nand I_47821 (I815503,I72251,I72260);
and I_47822 (I815520,I815503,I72254);
DFFARX1 I_47823 (I815520,I2507,I815452,I815546,);
DFFARX1 I_47824 (I815546,I2507,I815452,I815441,);
DFFARX1 I_47825 (I72272,I2507,I815452,I815577,);
nand I_47826 (I815585,I815577,I72263);
not I_47827 (I815602,I815585);
DFFARX1 I_47828 (I815602,I2507,I815452,I815628,);
not I_47829 (I815636,I815628);
nor I_47830 (I815444,I815486,I815636);
DFFARX1 I_47831 (I72257,I2507,I815452,I815676,);
nor I_47832 (I815435,I815676,I815546);
nor I_47833 (I815426,I815676,I815602);
nand I_47834 (I815712,I72269,I72266);
and I_47835 (I815729,I815712,I72254);
DFFARX1 I_47836 (I815729,I2507,I815452,I815755,);
not I_47837 (I815763,I815755);
nand I_47838 (I815780,I815763,I815676);
nand I_47839 (I815429,I815763,I815585);
nor I_47840 (I815811,I72251,I72266);
and I_47841 (I815828,I815676,I815811);
nor I_47842 (I815845,I815763,I815828);
DFFARX1 I_47843 (I815845,I2507,I815452,I815438,);
nor I_47844 (I815876,I815478,I815811);
DFFARX1 I_47845 (I815876,I2507,I815452,I815423,);
nor I_47846 (I815907,I815755,I815811);
not I_47847 (I815924,I815907);
nand I_47848 (I815432,I815924,I815780);
not I_47849 (I815979,I2514);
DFFARX1 I_47850 (I585071,I2507,I815979,I816005,);
not I_47851 (I816013,I816005);
nand I_47852 (I816030,I585056,I585077);
and I_47853 (I816047,I816030,I585065);
DFFARX1 I_47854 (I816047,I2507,I815979,I816073,);
DFFARX1 I_47855 (I816073,I2507,I815979,I815968,);
DFFARX1 I_47856 (I585059,I2507,I815979,I816104,);
nand I_47857 (I816112,I816104,I585068);
not I_47858 (I816129,I816112);
DFFARX1 I_47859 (I816129,I2507,I815979,I816155,);
not I_47860 (I816163,I816155);
nor I_47861 (I815971,I816013,I816163);
DFFARX1 I_47862 (I585074,I2507,I815979,I816203,);
nor I_47863 (I815962,I816203,I816073);
nor I_47864 (I815953,I816203,I816129);
nand I_47865 (I816239,I585056,I585059);
and I_47866 (I816256,I816239,I585080);
DFFARX1 I_47867 (I816256,I2507,I815979,I816282,);
not I_47868 (I816290,I816282);
nand I_47869 (I816307,I816290,I816203);
nand I_47870 (I815956,I816290,I816112);
nor I_47871 (I816338,I585062,I585059);
and I_47872 (I816355,I816203,I816338);
nor I_47873 (I816372,I816290,I816355);
DFFARX1 I_47874 (I816372,I2507,I815979,I815965,);
nor I_47875 (I816403,I816005,I816338);
DFFARX1 I_47876 (I816403,I2507,I815979,I815950,);
nor I_47877 (I816434,I816282,I816338);
not I_47878 (I816451,I816434);
nand I_47879 (I815959,I816451,I816307);
not I_47880 (I816506,I2514);
DFFARX1 I_47881 (I751520,I2507,I816506,I816532,);
not I_47882 (I816540,I816532);
nand I_47883 (I816557,I751523,I751520);
and I_47884 (I816574,I816557,I751532);
DFFARX1 I_47885 (I816574,I2507,I816506,I816600,);
DFFARX1 I_47886 (I816600,I2507,I816506,I816495,);
DFFARX1 I_47887 (I751529,I2507,I816506,I816631,);
nand I_47888 (I816639,I816631,I751535);
not I_47889 (I816656,I816639);
DFFARX1 I_47890 (I816656,I2507,I816506,I816682,);
not I_47891 (I816690,I816682);
nor I_47892 (I816498,I816540,I816690);
DFFARX1 I_47893 (I751544,I2507,I816506,I816730,);
nor I_47894 (I816489,I816730,I816600);
nor I_47895 (I816480,I816730,I816656);
nand I_47896 (I816766,I751538,I751526);
and I_47897 (I816783,I816766,I751523);
DFFARX1 I_47898 (I816783,I2507,I816506,I816809,);
not I_47899 (I816817,I816809);
nand I_47900 (I816834,I816817,I816730);
nand I_47901 (I816483,I816817,I816639);
nor I_47902 (I816865,I751541,I751526);
and I_47903 (I816882,I816730,I816865);
nor I_47904 (I816899,I816817,I816882);
DFFARX1 I_47905 (I816899,I2507,I816506,I816492,);
nor I_47906 (I816930,I816532,I816865);
DFFARX1 I_47907 (I816930,I2507,I816506,I816477,);
nor I_47908 (I816961,I816809,I816865);
not I_47909 (I816978,I816961);
nand I_47910 (I816486,I816978,I816834);
not I_47911 (I817033,I2514);
DFFARX1 I_47912 (I636498,I2507,I817033,I817059,);
not I_47913 (I817067,I817059);
nand I_47914 (I817084,I636501,I636498);
and I_47915 (I817101,I817084,I636510);
DFFARX1 I_47916 (I817101,I2507,I817033,I817127,);
DFFARX1 I_47917 (I817127,I2507,I817033,I817022,);
DFFARX1 I_47918 (I636507,I2507,I817033,I817158,);
nand I_47919 (I817166,I817158,I636513);
not I_47920 (I817183,I817166);
DFFARX1 I_47921 (I817183,I2507,I817033,I817209,);
not I_47922 (I817217,I817209);
nor I_47923 (I817025,I817067,I817217);
DFFARX1 I_47924 (I636522,I2507,I817033,I817257,);
nor I_47925 (I817016,I817257,I817127);
nor I_47926 (I817007,I817257,I817183);
nand I_47927 (I817293,I636516,I636504);
and I_47928 (I817310,I817293,I636501);
DFFARX1 I_47929 (I817310,I2507,I817033,I817336,);
not I_47930 (I817344,I817336);
nand I_47931 (I817361,I817344,I817257);
nand I_47932 (I817010,I817344,I817166);
nor I_47933 (I817392,I636519,I636504);
and I_47934 (I817409,I817257,I817392);
nor I_47935 (I817426,I817344,I817409);
DFFARX1 I_47936 (I817426,I2507,I817033,I817019,);
nor I_47937 (I817457,I817059,I817392);
DFFARX1 I_47938 (I817457,I2507,I817033,I817004,);
nor I_47939 (I817488,I817336,I817392);
not I_47940 (I817505,I817488);
nand I_47941 (I817013,I817505,I817361);
not I_47942 (I817560,I2514);
DFFARX1 I_47943 (I520870,I2507,I817560,I817586,);
not I_47944 (I817594,I817586);
nand I_47945 (I817611,I520888,I520879);
and I_47946 (I817628,I817611,I520882);
DFFARX1 I_47947 (I817628,I2507,I817560,I817654,);
DFFARX1 I_47948 (I817654,I2507,I817560,I817549,);
DFFARX1 I_47949 (I520876,I2507,I817560,I817685,);
nand I_47950 (I817693,I817685,I520867);
not I_47951 (I817710,I817693);
DFFARX1 I_47952 (I817710,I2507,I817560,I817736,);
not I_47953 (I817744,I817736);
nor I_47954 (I817552,I817594,I817744);
DFFARX1 I_47955 (I520873,I2507,I817560,I817784,);
nor I_47956 (I817543,I817784,I817654);
nor I_47957 (I817534,I817784,I817710);
nand I_47958 (I817820,I520867,I520864);
and I_47959 (I817837,I817820,I520885);
DFFARX1 I_47960 (I817837,I2507,I817560,I817863,);
not I_47961 (I817871,I817863);
nand I_47962 (I817888,I817871,I817784);
nand I_47963 (I817537,I817871,I817693);
nor I_47964 (I817919,I520864,I520864);
and I_47965 (I817936,I817784,I817919);
nor I_47966 (I817953,I817871,I817936);
DFFARX1 I_47967 (I817953,I2507,I817560,I817546,);
nor I_47968 (I817984,I817586,I817919);
DFFARX1 I_47969 (I817984,I2507,I817560,I817531,);
nor I_47970 (I818015,I817863,I817919);
not I_47971 (I818032,I818015);
nand I_47972 (I817540,I818032,I817888);
not I_47973 (I818087,I2514);
DFFARX1 I_47974 (I464821,I2507,I818087,I818113,);
not I_47975 (I818121,I818113);
nand I_47976 (I818138,I464818,I464827);
and I_47977 (I818155,I818138,I464836);
DFFARX1 I_47978 (I818155,I2507,I818087,I818181,);
DFFARX1 I_47979 (I818181,I2507,I818087,I818076,);
DFFARX1 I_47980 (I464839,I2507,I818087,I818212,);
nand I_47981 (I818220,I818212,I464842);
not I_47982 (I818237,I818220);
DFFARX1 I_47983 (I818237,I2507,I818087,I818263,);
not I_47984 (I818271,I818263);
nor I_47985 (I818079,I818121,I818271);
DFFARX1 I_47986 (I464815,I2507,I818087,I818311,);
nor I_47987 (I818070,I818311,I818181);
nor I_47988 (I818061,I818311,I818237);
nand I_47989 (I818347,I464830,I464833);
and I_47990 (I818364,I818347,I464824);
DFFARX1 I_47991 (I818364,I2507,I818087,I818390,);
not I_47992 (I818398,I818390);
nand I_47993 (I818415,I818398,I818311);
nand I_47994 (I818064,I818398,I818220);
nor I_47995 (I818446,I464815,I464833);
and I_47996 (I818463,I818311,I818446);
nor I_47997 (I818480,I818398,I818463);
DFFARX1 I_47998 (I818480,I2507,I818087,I818073,);
nor I_47999 (I818511,I818113,I818446);
DFFARX1 I_48000 (I818511,I2507,I818087,I818058,);
nor I_48001 (I818542,I818390,I818446);
not I_48002 (I818559,I818542);
nand I_48003 (I818067,I818559,I818415);
not I_48004 (I818614,I2514);
DFFARX1 I_48005 (I557905,I2507,I818614,I818640,);
not I_48006 (I818648,I818640);
nand I_48007 (I818665,I557890,I557911);
and I_48008 (I818682,I818665,I557899);
DFFARX1 I_48009 (I818682,I2507,I818614,I818708,);
DFFARX1 I_48010 (I818708,I2507,I818614,I818603,);
DFFARX1 I_48011 (I557893,I2507,I818614,I818739,);
nand I_48012 (I818747,I818739,I557902);
not I_48013 (I818764,I818747);
DFFARX1 I_48014 (I818764,I2507,I818614,I818790,);
not I_48015 (I818798,I818790);
nor I_48016 (I818606,I818648,I818798);
DFFARX1 I_48017 (I557908,I2507,I818614,I818838,);
nor I_48018 (I818597,I818838,I818708);
nor I_48019 (I818588,I818838,I818764);
nand I_48020 (I818874,I557890,I557893);
and I_48021 (I818891,I818874,I557914);
DFFARX1 I_48022 (I818891,I2507,I818614,I818917,);
not I_48023 (I818925,I818917);
nand I_48024 (I818942,I818925,I818838);
nand I_48025 (I818591,I818925,I818747);
nor I_48026 (I818973,I557896,I557893);
and I_48027 (I818990,I818838,I818973);
nor I_48028 (I819007,I818925,I818990);
DFFARX1 I_48029 (I819007,I2507,I818614,I818600,);
nor I_48030 (I819038,I818640,I818973);
DFFARX1 I_48031 (I819038,I2507,I818614,I818585,);
nor I_48032 (I819069,I818917,I818973);
not I_48033 (I819086,I819069);
nand I_48034 (I818594,I819086,I818942);
not I_48035 (I819141,I2514);
DFFARX1 I_48036 (I335046,I2507,I819141,I819167,);
not I_48037 (I819175,I819167);
nand I_48038 (I819192,I335037,I335037);
and I_48039 (I819209,I819192,I335055);
DFFARX1 I_48040 (I819209,I2507,I819141,I819235,);
DFFARX1 I_48041 (I819235,I2507,I819141,I819130,);
DFFARX1 I_48042 (I335058,I2507,I819141,I819266,);
nand I_48043 (I819274,I819266,I335040);
not I_48044 (I819291,I819274);
DFFARX1 I_48045 (I819291,I2507,I819141,I819317,);
not I_48046 (I819325,I819317);
nor I_48047 (I819133,I819175,I819325);
DFFARX1 I_48048 (I335052,I2507,I819141,I819365,);
nor I_48049 (I819124,I819365,I819235);
nor I_48050 (I819115,I819365,I819291);
nand I_48051 (I819401,I335064,I335043);
and I_48052 (I819418,I819401,I335049);
DFFARX1 I_48053 (I819418,I2507,I819141,I819444,);
not I_48054 (I819452,I819444);
nand I_48055 (I819469,I819452,I819365);
nand I_48056 (I819118,I819452,I819274);
nor I_48057 (I819500,I335061,I335043);
and I_48058 (I819517,I819365,I819500);
nor I_48059 (I819534,I819452,I819517);
DFFARX1 I_48060 (I819534,I2507,I819141,I819127,);
nor I_48061 (I819565,I819167,I819500);
DFFARX1 I_48062 (I819565,I2507,I819141,I819112,);
nor I_48063 (I819596,I819444,I819500);
not I_48064 (I819613,I819596);
nand I_48065 (I819121,I819613,I819469);
not I_48066 (I819668,I2514);
DFFARX1 I_48067 (I593163,I2507,I819668,I819694,);
not I_48068 (I819702,I819694);
nand I_48069 (I819719,I593148,I593169);
and I_48070 (I819736,I819719,I593157);
DFFARX1 I_48071 (I819736,I2507,I819668,I819762,);
DFFARX1 I_48072 (I819762,I2507,I819668,I819657,);
DFFARX1 I_48073 (I593151,I2507,I819668,I819793,);
nand I_48074 (I819801,I819793,I593160);
not I_48075 (I819818,I819801);
DFFARX1 I_48076 (I819818,I2507,I819668,I819844,);
not I_48077 (I819852,I819844);
nor I_48078 (I819660,I819702,I819852);
DFFARX1 I_48079 (I593166,I2507,I819668,I819892,);
nor I_48080 (I819651,I819892,I819762);
nor I_48081 (I819642,I819892,I819818);
nand I_48082 (I819928,I593148,I593151);
and I_48083 (I819945,I819928,I593172);
DFFARX1 I_48084 (I819945,I2507,I819668,I819971,);
not I_48085 (I819979,I819971);
nand I_48086 (I819996,I819979,I819892);
nand I_48087 (I819645,I819979,I819801);
nor I_48088 (I820027,I593154,I593151);
and I_48089 (I820044,I819892,I820027);
nor I_48090 (I820061,I819979,I820044);
DFFARX1 I_48091 (I820061,I2507,I819668,I819654,);
nor I_48092 (I820092,I819694,I820027);
DFFARX1 I_48093 (I820092,I2507,I819668,I819639,);
nor I_48094 (I820123,I819971,I820027);
not I_48095 (I820140,I820123);
nand I_48096 (I819648,I820140,I819996);
not I_48097 (I820195,I2514);
DFFARX1 I_48098 (I65424,I2507,I820195,I820221,);
not I_48099 (I820229,I820221);
nand I_48100 (I820246,I65400,I65409);
and I_48101 (I820263,I820246,I65403);
DFFARX1 I_48102 (I820263,I2507,I820195,I820289,);
DFFARX1 I_48103 (I820289,I2507,I820195,I820184,);
DFFARX1 I_48104 (I65421,I2507,I820195,I820320,);
nand I_48105 (I820328,I820320,I65412);
not I_48106 (I820345,I820328);
DFFARX1 I_48107 (I820345,I2507,I820195,I820371,);
not I_48108 (I820379,I820371);
nor I_48109 (I820187,I820229,I820379);
DFFARX1 I_48110 (I65406,I2507,I820195,I820419,);
nor I_48111 (I820178,I820419,I820289);
nor I_48112 (I820169,I820419,I820345);
nand I_48113 (I820455,I65418,I65415);
and I_48114 (I820472,I820455,I65403);
DFFARX1 I_48115 (I820472,I2507,I820195,I820498,);
not I_48116 (I820506,I820498);
nand I_48117 (I820523,I820506,I820419);
nand I_48118 (I820172,I820506,I820328);
nor I_48119 (I820554,I65400,I65415);
and I_48120 (I820571,I820419,I820554);
nor I_48121 (I820588,I820506,I820571);
DFFARX1 I_48122 (I820588,I2507,I820195,I820181,);
nor I_48123 (I820619,I820221,I820554);
DFFARX1 I_48124 (I820619,I2507,I820195,I820166,);
nor I_48125 (I820650,I820498,I820554);
not I_48126 (I820667,I820650);
nand I_48127 (I820175,I820667,I820523);
not I_48128 (I820722,I2514);
DFFARX1 I_48129 (I63843,I2507,I820722,I820748,);
not I_48130 (I820756,I820748);
nand I_48131 (I820773,I63819,I63828);
and I_48132 (I820790,I820773,I63822);
DFFARX1 I_48133 (I820790,I2507,I820722,I820816,);
DFFARX1 I_48134 (I820816,I2507,I820722,I820711,);
DFFARX1 I_48135 (I63840,I2507,I820722,I820847,);
nand I_48136 (I820855,I820847,I63831);
not I_48137 (I820872,I820855);
DFFARX1 I_48138 (I820872,I2507,I820722,I820898,);
not I_48139 (I820906,I820898);
nor I_48140 (I820714,I820756,I820906);
DFFARX1 I_48141 (I63825,I2507,I820722,I820946,);
nor I_48142 (I820705,I820946,I820816);
nor I_48143 (I820696,I820946,I820872);
nand I_48144 (I820982,I63837,I63834);
and I_48145 (I820999,I820982,I63822);
DFFARX1 I_48146 (I820999,I2507,I820722,I821025,);
not I_48147 (I821033,I821025);
nand I_48148 (I821050,I821033,I820946);
nand I_48149 (I820699,I821033,I820855);
nor I_48150 (I821081,I63819,I63834);
and I_48151 (I821098,I820946,I821081);
nor I_48152 (I821115,I821033,I821098);
DFFARX1 I_48153 (I821115,I2507,I820722,I820708,);
nor I_48154 (I821146,I820748,I821081);
DFFARX1 I_48155 (I821146,I2507,I820722,I820693,);
nor I_48156 (I821177,I821025,I821081);
not I_48157 (I821194,I821177);
nand I_48158 (I820702,I821194,I821050);
not I_48159 (I821249,I2514);
DFFARX1 I_48160 (I57519,I2507,I821249,I821275,);
not I_48161 (I821283,I821275);
nand I_48162 (I821300,I57495,I57504);
and I_48163 (I821317,I821300,I57498);
DFFARX1 I_48164 (I821317,I2507,I821249,I821343,);
DFFARX1 I_48165 (I821343,I2507,I821249,I821238,);
DFFARX1 I_48166 (I57516,I2507,I821249,I821374,);
nand I_48167 (I821382,I821374,I57507);
not I_48168 (I821399,I821382);
DFFARX1 I_48169 (I821399,I2507,I821249,I821425,);
not I_48170 (I821433,I821425);
nor I_48171 (I821241,I821283,I821433);
DFFARX1 I_48172 (I57501,I2507,I821249,I821473,);
nor I_48173 (I821232,I821473,I821343);
nor I_48174 (I821223,I821473,I821399);
nand I_48175 (I821509,I57513,I57510);
and I_48176 (I821526,I821509,I57498);
DFFARX1 I_48177 (I821526,I2507,I821249,I821552,);
not I_48178 (I821560,I821552);
nand I_48179 (I821577,I821560,I821473);
nand I_48180 (I821226,I821560,I821382);
nor I_48181 (I821608,I57495,I57510);
and I_48182 (I821625,I821473,I821608);
nor I_48183 (I821642,I821560,I821625);
DFFARX1 I_48184 (I821642,I2507,I821249,I821235,);
nor I_48185 (I821673,I821275,I821608);
DFFARX1 I_48186 (I821673,I2507,I821249,I821220,);
nor I_48187 (I821704,I821552,I821608);
not I_48188 (I821721,I821704);
nand I_48189 (I821229,I821721,I821577);
not I_48190 (I821776,I2514);
DFFARX1 I_48191 (I897910,I2507,I821776,I821802,);
not I_48192 (I821810,I821802);
nand I_48193 (I821827,I897925,I897907);
and I_48194 (I821844,I821827,I897907);
DFFARX1 I_48195 (I821844,I2507,I821776,I821870,);
DFFARX1 I_48196 (I821870,I2507,I821776,I821765,);
DFFARX1 I_48197 (I897916,I2507,I821776,I821901,);
nand I_48198 (I821909,I821901,I897934);
not I_48199 (I821926,I821909);
DFFARX1 I_48200 (I821926,I2507,I821776,I821952,);
not I_48201 (I821960,I821952);
nor I_48202 (I821768,I821810,I821960);
DFFARX1 I_48203 (I897931,I2507,I821776,I822000,);
nor I_48204 (I821759,I822000,I821870);
nor I_48205 (I821750,I822000,I821926);
nand I_48206 (I822036,I897928,I897919);
and I_48207 (I822053,I822036,I897913);
DFFARX1 I_48208 (I822053,I2507,I821776,I822079,);
not I_48209 (I822087,I822079);
nand I_48210 (I822104,I822087,I822000);
nand I_48211 (I821753,I822087,I821909);
nor I_48212 (I822135,I897922,I897919);
and I_48213 (I822152,I822000,I822135);
nor I_48214 (I822169,I822087,I822152);
DFFARX1 I_48215 (I822169,I2507,I821776,I821762,);
nor I_48216 (I822200,I821802,I822135);
DFFARX1 I_48217 (I822200,I2507,I821776,I821747,);
nor I_48218 (I822231,I822079,I822135);
not I_48219 (I822248,I822231);
nand I_48220 (I821756,I822248,I822104);
not I_48221 (I822303,I2514);
DFFARX1 I_48222 (I465909,I2507,I822303,I822329,);
not I_48223 (I822337,I822329);
nand I_48224 (I822354,I465906,I465915);
and I_48225 (I822371,I822354,I465924);
DFFARX1 I_48226 (I822371,I2507,I822303,I822397,);
DFFARX1 I_48227 (I822397,I2507,I822303,I822292,);
DFFARX1 I_48228 (I465927,I2507,I822303,I822428,);
nand I_48229 (I822436,I822428,I465930);
not I_48230 (I822453,I822436);
DFFARX1 I_48231 (I822453,I2507,I822303,I822479,);
not I_48232 (I822487,I822479);
nor I_48233 (I822295,I822337,I822487);
DFFARX1 I_48234 (I465903,I2507,I822303,I822527,);
nor I_48235 (I822286,I822527,I822397);
nor I_48236 (I822277,I822527,I822453);
nand I_48237 (I822563,I465918,I465921);
and I_48238 (I822580,I822563,I465912);
DFFARX1 I_48239 (I822580,I2507,I822303,I822606,);
not I_48240 (I822614,I822606);
nand I_48241 (I822631,I822614,I822527);
nand I_48242 (I822280,I822614,I822436);
nor I_48243 (I822662,I465903,I465921);
and I_48244 (I822679,I822527,I822662);
nor I_48245 (I822696,I822614,I822679);
DFFARX1 I_48246 (I822696,I2507,I822303,I822289,);
nor I_48247 (I822727,I822329,I822662);
DFFARX1 I_48248 (I822727,I2507,I822303,I822274,);
nor I_48249 (I822758,I822606,I822662);
not I_48250 (I822775,I822758);
nand I_48251 (I822283,I822775,I822631);
not I_48252 (I822830,I2514);
DFFARX1 I_48253 (I449589,I2507,I822830,I822856,);
not I_48254 (I822864,I822856);
nand I_48255 (I822881,I449586,I449595);
and I_48256 (I822898,I822881,I449604);
DFFARX1 I_48257 (I822898,I2507,I822830,I822924,);
DFFARX1 I_48258 (I822924,I2507,I822830,I822819,);
DFFARX1 I_48259 (I449607,I2507,I822830,I822955,);
nand I_48260 (I822963,I822955,I449610);
not I_48261 (I822980,I822963);
DFFARX1 I_48262 (I822980,I2507,I822830,I823006,);
not I_48263 (I823014,I823006);
nor I_48264 (I822822,I822864,I823014);
DFFARX1 I_48265 (I449583,I2507,I822830,I823054,);
nor I_48266 (I822813,I823054,I822924);
nor I_48267 (I822804,I823054,I822980);
nand I_48268 (I823090,I449598,I449601);
and I_48269 (I823107,I823090,I449592);
DFFARX1 I_48270 (I823107,I2507,I822830,I823133,);
not I_48271 (I823141,I823133);
nand I_48272 (I823158,I823141,I823054);
nand I_48273 (I822807,I823141,I822963);
nor I_48274 (I823189,I449583,I449601);
and I_48275 (I823206,I823054,I823189);
nor I_48276 (I823223,I823141,I823206);
DFFARX1 I_48277 (I823223,I2507,I822830,I822816,);
nor I_48278 (I823254,I822856,I823189);
DFFARX1 I_48279 (I823254,I2507,I822830,I822801,);
nor I_48280 (I823285,I823133,I823189);
not I_48281 (I823302,I823285);
nand I_48282 (I822810,I823302,I823158);
not I_48283 (I823357,I2514);
DFFARX1 I_48284 (I1282516,I2507,I823357,I823383,);
not I_48285 (I823391,I823383);
nand I_48286 (I823408,I1282498,I1282501);
and I_48287 (I823425,I823408,I1282513);
DFFARX1 I_48288 (I823425,I2507,I823357,I823451,);
DFFARX1 I_48289 (I823451,I2507,I823357,I823346,);
DFFARX1 I_48290 (I1282522,I2507,I823357,I823482,);
nand I_48291 (I823490,I823482,I1282507);
not I_48292 (I823507,I823490);
DFFARX1 I_48293 (I823507,I2507,I823357,I823533,);
not I_48294 (I823541,I823533);
nor I_48295 (I823349,I823391,I823541);
DFFARX1 I_48296 (I1282519,I2507,I823357,I823581,);
nor I_48297 (I823340,I823581,I823451);
nor I_48298 (I823331,I823581,I823507);
nand I_48299 (I823617,I1282510,I1282504);
and I_48300 (I823634,I823617,I1282498);
DFFARX1 I_48301 (I823634,I2507,I823357,I823660,);
not I_48302 (I823668,I823660);
nand I_48303 (I823685,I823668,I823581);
nand I_48304 (I823334,I823668,I823490);
nor I_48305 (I823716,I1282501,I1282504);
and I_48306 (I823733,I823581,I823716);
nor I_48307 (I823750,I823668,I823733);
DFFARX1 I_48308 (I823750,I2507,I823357,I823343,);
nor I_48309 (I823781,I823383,I823716);
DFFARX1 I_48310 (I823781,I2507,I823357,I823328,);
nor I_48311 (I823812,I823660,I823716);
not I_48312 (I823829,I823812);
nand I_48313 (I823337,I823829,I823685);
not I_48314 (I823884,I2514);
DFFARX1 I_48315 (I594897,I2507,I823884,I823910,);
not I_48316 (I823918,I823910);
nand I_48317 (I823935,I594882,I594903);
and I_48318 (I823952,I823935,I594891);
DFFARX1 I_48319 (I823952,I2507,I823884,I823978,);
DFFARX1 I_48320 (I823978,I2507,I823884,I823873,);
DFFARX1 I_48321 (I594885,I2507,I823884,I824009,);
nand I_48322 (I824017,I824009,I594894);
not I_48323 (I824034,I824017);
DFFARX1 I_48324 (I824034,I2507,I823884,I824060,);
not I_48325 (I824068,I824060);
nor I_48326 (I823876,I823918,I824068);
DFFARX1 I_48327 (I594900,I2507,I823884,I824108,);
nor I_48328 (I823867,I824108,I823978);
nor I_48329 (I823858,I824108,I824034);
nand I_48330 (I824144,I594882,I594885);
and I_48331 (I824161,I824144,I594906);
DFFARX1 I_48332 (I824161,I2507,I823884,I824187,);
not I_48333 (I824195,I824187);
nand I_48334 (I824212,I824195,I824108);
nand I_48335 (I823861,I824195,I824017);
nor I_48336 (I824243,I594888,I594885);
and I_48337 (I824260,I824108,I824243);
nor I_48338 (I824277,I824195,I824260);
DFFARX1 I_48339 (I824277,I2507,I823884,I823870,);
nor I_48340 (I824308,I823910,I824243);
DFFARX1 I_48341 (I824308,I2507,I823884,I823855,);
nor I_48342 (I824339,I824187,I824243);
not I_48343 (I824356,I824339);
nand I_48344 (I823864,I824356,I824212);
not I_48345 (I824411,I2514);
DFFARX1 I_48346 (I1136996,I2507,I824411,I824437,);
not I_48347 (I824445,I824437);
nand I_48348 (I824462,I1136978,I1136978);
and I_48349 (I824479,I824462,I1136984);
DFFARX1 I_48350 (I824479,I2507,I824411,I824505,);
DFFARX1 I_48351 (I824505,I2507,I824411,I824400,);
DFFARX1 I_48352 (I1136981,I2507,I824411,I824536,);
nand I_48353 (I824544,I824536,I1136990);
not I_48354 (I824561,I824544);
DFFARX1 I_48355 (I824561,I2507,I824411,I824587,);
not I_48356 (I824595,I824587);
nor I_48357 (I824403,I824445,I824595);
DFFARX1 I_48358 (I1137002,I2507,I824411,I824635,);
nor I_48359 (I824394,I824635,I824505);
nor I_48360 (I824385,I824635,I824561);
nand I_48361 (I824671,I1136993,I1136987);
and I_48362 (I824688,I824671,I1136981);
DFFARX1 I_48363 (I824688,I2507,I824411,I824714,);
not I_48364 (I824722,I824714);
nand I_48365 (I824739,I824722,I824635);
nand I_48366 (I824388,I824722,I824544);
nor I_48367 (I824770,I1136999,I1136987);
and I_48368 (I824787,I824635,I824770);
nor I_48369 (I824804,I824722,I824787);
DFFARX1 I_48370 (I824804,I2507,I824411,I824397,);
nor I_48371 (I824835,I824437,I824770);
DFFARX1 I_48372 (I824835,I2507,I824411,I824382,);
nor I_48373 (I824866,I824714,I824770);
not I_48374 (I824883,I824866);
nand I_48375 (I824391,I824883,I824739);
not I_48376 (I824938,I2514);
DFFARX1 I_48377 (I948298,I2507,I824938,I824964,);
not I_48378 (I824972,I824964);
nand I_48379 (I824989,I948313,I948295);
and I_48380 (I825006,I824989,I948295);
DFFARX1 I_48381 (I825006,I2507,I824938,I825032,);
DFFARX1 I_48382 (I825032,I2507,I824938,I824927,);
DFFARX1 I_48383 (I948304,I2507,I824938,I825063,);
nand I_48384 (I825071,I825063,I948322);
not I_48385 (I825088,I825071);
DFFARX1 I_48386 (I825088,I2507,I824938,I825114,);
not I_48387 (I825122,I825114);
nor I_48388 (I824930,I824972,I825122);
DFFARX1 I_48389 (I948319,I2507,I824938,I825162,);
nor I_48390 (I824921,I825162,I825032);
nor I_48391 (I824912,I825162,I825088);
nand I_48392 (I825198,I948316,I948307);
and I_48393 (I825215,I825198,I948301);
DFFARX1 I_48394 (I825215,I2507,I824938,I825241,);
not I_48395 (I825249,I825241);
nand I_48396 (I825266,I825249,I825162);
nand I_48397 (I824915,I825249,I825071);
nor I_48398 (I825297,I948310,I948307);
and I_48399 (I825314,I825162,I825297);
nor I_48400 (I825331,I825249,I825314);
DFFARX1 I_48401 (I825331,I2507,I824938,I824924,);
nor I_48402 (I825362,I824964,I825297);
DFFARX1 I_48403 (I825362,I2507,I824938,I824909,);
nor I_48404 (I825393,I825241,I825297);
not I_48405 (I825410,I825393);
nand I_48406 (I824918,I825410,I825266);
not I_48407 (I825465,I2514);
DFFARX1 I_48408 (I1324367,I2507,I825465,I825491,);
not I_48409 (I825499,I825491);
nand I_48410 (I825516,I1324364,I1324373);
and I_48411 (I825533,I825516,I1324352);
DFFARX1 I_48412 (I825533,I2507,I825465,I825559,);
DFFARX1 I_48413 (I825559,I2507,I825465,I825454,);
DFFARX1 I_48414 (I1324355,I2507,I825465,I825590,);
nand I_48415 (I825598,I825590,I1324370);
not I_48416 (I825615,I825598);
DFFARX1 I_48417 (I825615,I2507,I825465,I825641,);
not I_48418 (I825649,I825641);
nor I_48419 (I825457,I825499,I825649);
DFFARX1 I_48420 (I1324376,I2507,I825465,I825689,);
nor I_48421 (I825448,I825689,I825559);
nor I_48422 (I825439,I825689,I825615);
nand I_48423 (I825725,I1324358,I1324379);
and I_48424 (I825742,I825725,I1324361);
DFFARX1 I_48425 (I825742,I2507,I825465,I825768,);
not I_48426 (I825776,I825768);
nand I_48427 (I825793,I825776,I825689);
nand I_48428 (I825442,I825776,I825598);
nor I_48429 (I825824,I1324352,I1324379);
and I_48430 (I825841,I825689,I825824);
nor I_48431 (I825858,I825776,I825841);
DFFARX1 I_48432 (I825858,I2507,I825465,I825451,);
nor I_48433 (I825889,I825491,I825824);
DFFARX1 I_48434 (I825889,I2507,I825465,I825436,);
nor I_48435 (I825920,I825768,I825824);
not I_48436 (I825937,I825920);
nand I_48437 (I825445,I825937,I825793);
not I_48438 (I825992,I2514);
DFFARX1 I_48439 (I1047737,I2507,I825992,I826018,);
not I_48440 (I826026,I826018);
nand I_48441 (I826043,I1047746,I1047734);
and I_48442 (I826060,I826043,I1047731);
DFFARX1 I_48443 (I826060,I2507,I825992,I826086,);
DFFARX1 I_48444 (I826086,I2507,I825992,I825981,);
DFFARX1 I_48445 (I1047731,I2507,I825992,I826117,);
nand I_48446 (I826125,I826117,I1047728);
not I_48447 (I826142,I826125);
DFFARX1 I_48448 (I826142,I2507,I825992,I826168,);
not I_48449 (I826176,I826168);
nor I_48450 (I825984,I826026,I826176);
DFFARX1 I_48451 (I1047734,I2507,I825992,I826216,);
nor I_48452 (I825975,I826216,I826086);
nor I_48453 (I825966,I826216,I826142);
nand I_48454 (I826252,I1047749,I1047740);
and I_48455 (I826269,I826252,I1047743);
DFFARX1 I_48456 (I826269,I2507,I825992,I826295,);
not I_48457 (I826303,I826295);
nand I_48458 (I826320,I826303,I826216);
nand I_48459 (I825969,I826303,I826125);
nor I_48460 (I826351,I1047728,I1047740);
and I_48461 (I826368,I826216,I826351);
nor I_48462 (I826385,I826303,I826368);
DFFARX1 I_48463 (I826385,I2507,I825992,I825978,);
nor I_48464 (I826416,I826018,I826351);
DFFARX1 I_48465 (I826416,I2507,I825992,I825963,);
nor I_48466 (I826447,I826295,I826351);
not I_48467 (I826464,I826447);
nand I_48468 (I825972,I826464,I826320);
not I_48469 (I826519,I2514);
DFFARX1 I_48470 (I344532,I2507,I826519,I826545,);
not I_48471 (I826553,I826545);
nand I_48472 (I826570,I344523,I344523);
and I_48473 (I826587,I826570,I344541);
DFFARX1 I_48474 (I826587,I2507,I826519,I826613,);
DFFARX1 I_48475 (I826613,I2507,I826519,I826508,);
DFFARX1 I_48476 (I344544,I2507,I826519,I826644,);
nand I_48477 (I826652,I826644,I344526);
not I_48478 (I826669,I826652);
DFFARX1 I_48479 (I826669,I2507,I826519,I826695,);
not I_48480 (I826703,I826695);
nor I_48481 (I826511,I826553,I826703);
DFFARX1 I_48482 (I344538,I2507,I826519,I826743,);
nor I_48483 (I826502,I826743,I826613);
nor I_48484 (I826493,I826743,I826669);
nand I_48485 (I826779,I344550,I344529);
and I_48486 (I826796,I826779,I344535);
DFFARX1 I_48487 (I826796,I2507,I826519,I826822,);
not I_48488 (I826830,I826822);
nand I_48489 (I826847,I826830,I826743);
nand I_48490 (I826496,I826830,I826652);
nor I_48491 (I826878,I344547,I344529);
and I_48492 (I826895,I826743,I826878);
nor I_48493 (I826912,I826830,I826895);
DFFARX1 I_48494 (I826912,I2507,I826519,I826505,);
nor I_48495 (I826943,I826545,I826878);
DFFARX1 I_48496 (I826943,I2507,I826519,I826490,);
nor I_48497 (I826974,I826822,I826878);
not I_48498 (I826991,I826974);
nand I_48499 (I826499,I826991,I826847);
not I_48500 (I827046,I2514);
DFFARX1 I_48501 (I1163584,I2507,I827046,I827072,);
not I_48502 (I827080,I827072);
nand I_48503 (I827097,I1163566,I1163566);
and I_48504 (I827114,I827097,I1163572);
DFFARX1 I_48505 (I827114,I2507,I827046,I827140,);
DFFARX1 I_48506 (I827140,I2507,I827046,I827035,);
DFFARX1 I_48507 (I1163569,I2507,I827046,I827171,);
nand I_48508 (I827179,I827171,I1163578);
not I_48509 (I827196,I827179);
DFFARX1 I_48510 (I827196,I2507,I827046,I827222,);
not I_48511 (I827230,I827222);
nor I_48512 (I827038,I827080,I827230);
DFFARX1 I_48513 (I1163590,I2507,I827046,I827270,);
nor I_48514 (I827029,I827270,I827140);
nor I_48515 (I827020,I827270,I827196);
nand I_48516 (I827306,I1163581,I1163575);
and I_48517 (I827323,I827306,I1163569);
DFFARX1 I_48518 (I827323,I2507,I827046,I827349,);
not I_48519 (I827357,I827349);
nand I_48520 (I827374,I827357,I827270);
nand I_48521 (I827023,I827357,I827179);
nor I_48522 (I827405,I1163587,I1163575);
and I_48523 (I827422,I827270,I827405);
nor I_48524 (I827439,I827357,I827422);
DFFARX1 I_48525 (I827439,I2507,I827046,I827032,);
nor I_48526 (I827470,I827072,I827405);
DFFARX1 I_48527 (I827470,I2507,I827046,I827017,);
nor I_48528 (I827501,I827349,I827405);
not I_48529 (I827518,I827501);
nand I_48530 (I827026,I827518,I827374);
not I_48531 (I827573,I2514);
DFFARX1 I_48532 (I702390,I2507,I827573,I827599,);
not I_48533 (I827607,I827599);
nand I_48534 (I827624,I702393,I702390);
and I_48535 (I827641,I827624,I702402);
DFFARX1 I_48536 (I827641,I2507,I827573,I827667,);
DFFARX1 I_48537 (I827667,I2507,I827573,I827562,);
DFFARX1 I_48538 (I702399,I2507,I827573,I827698,);
nand I_48539 (I827706,I827698,I702405);
not I_48540 (I827723,I827706);
DFFARX1 I_48541 (I827723,I2507,I827573,I827749,);
not I_48542 (I827757,I827749);
nor I_48543 (I827565,I827607,I827757);
DFFARX1 I_48544 (I702414,I2507,I827573,I827797,);
nor I_48545 (I827556,I827797,I827667);
nor I_48546 (I827547,I827797,I827723);
nand I_48547 (I827833,I702408,I702396);
and I_48548 (I827850,I827833,I702393);
DFFARX1 I_48549 (I827850,I2507,I827573,I827876,);
not I_48550 (I827884,I827876);
nand I_48551 (I827901,I827884,I827797);
nand I_48552 (I827550,I827884,I827706);
nor I_48553 (I827932,I702411,I702396);
and I_48554 (I827949,I827797,I827932);
nor I_48555 (I827966,I827884,I827949);
DFFARX1 I_48556 (I827966,I2507,I827573,I827559,);
nor I_48557 (I827997,I827599,I827932);
DFFARX1 I_48558 (I827997,I2507,I827573,I827544,);
nor I_48559 (I828028,I827876,I827932);
not I_48560 (I828045,I828028);
nand I_48561 (I827553,I828045,I827901);
not I_48562 (I828100,I2514);
DFFARX1 I_48563 (I980598,I2507,I828100,I828126,);
not I_48564 (I828134,I828126);
nand I_48565 (I828151,I980613,I980595);
and I_48566 (I828168,I828151,I980595);
DFFARX1 I_48567 (I828168,I2507,I828100,I828194,);
DFFARX1 I_48568 (I828194,I2507,I828100,I828089,);
DFFARX1 I_48569 (I980604,I2507,I828100,I828225,);
nand I_48570 (I828233,I828225,I980622);
not I_48571 (I828250,I828233);
DFFARX1 I_48572 (I828250,I2507,I828100,I828276,);
not I_48573 (I828284,I828276);
nor I_48574 (I828092,I828134,I828284);
DFFARX1 I_48575 (I980619,I2507,I828100,I828324,);
nor I_48576 (I828083,I828324,I828194);
nor I_48577 (I828074,I828324,I828250);
nand I_48578 (I828360,I980616,I980607);
and I_48579 (I828377,I828360,I980601);
DFFARX1 I_48580 (I828377,I2507,I828100,I828403,);
not I_48581 (I828411,I828403);
nand I_48582 (I828428,I828411,I828324);
nand I_48583 (I828077,I828411,I828233);
nor I_48584 (I828459,I980610,I980607);
and I_48585 (I828476,I828324,I828459);
nor I_48586 (I828493,I828411,I828476);
DFFARX1 I_48587 (I828493,I2507,I828100,I828086,);
nor I_48588 (I828524,I828126,I828459);
DFFARX1 I_48589 (I828524,I2507,I828100,I828071,);
nor I_48590 (I828555,I828403,I828459);
not I_48591 (I828572,I828555);
nand I_48592 (I828080,I828572,I828428);
not I_48593 (I828627,I2514);
DFFARX1 I_48594 (I459925,I2507,I828627,I828653,);
not I_48595 (I828661,I828653);
nand I_48596 (I828678,I459922,I459931);
and I_48597 (I828695,I828678,I459940);
DFFARX1 I_48598 (I828695,I2507,I828627,I828721,);
DFFARX1 I_48599 (I828721,I2507,I828627,I828616,);
DFFARX1 I_48600 (I459943,I2507,I828627,I828752,);
nand I_48601 (I828760,I828752,I459946);
not I_48602 (I828777,I828760);
DFFARX1 I_48603 (I828777,I2507,I828627,I828803,);
not I_48604 (I828811,I828803);
nor I_48605 (I828619,I828661,I828811);
DFFARX1 I_48606 (I459919,I2507,I828627,I828851,);
nor I_48607 (I828610,I828851,I828721);
nor I_48608 (I828601,I828851,I828777);
nand I_48609 (I828887,I459934,I459937);
and I_48610 (I828904,I828887,I459928);
DFFARX1 I_48611 (I828904,I2507,I828627,I828930,);
not I_48612 (I828938,I828930);
nand I_48613 (I828955,I828938,I828851);
nand I_48614 (I828604,I828938,I828760);
nor I_48615 (I828986,I459919,I459937);
and I_48616 (I829003,I828851,I828986);
nor I_48617 (I829020,I828938,I829003);
DFFARX1 I_48618 (I829020,I2507,I828627,I828613,);
nor I_48619 (I829051,I828653,I828986);
DFFARX1 I_48620 (I829051,I2507,I828627,I828598,);
nor I_48621 (I829082,I828930,I828986);
not I_48622 (I829099,I829082);
nand I_48623 (I828607,I829099,I828955);
not I_48624 (I829154,I2514);
DFFARX1 I_48625 (I1143354,I2507,I829154,I829180,);
not I_48626 (I829188,I829180);
nand I_48627 (I829205,I1143336,I1143336);
and I_48628 (I829222,I829205,I1143342);
DFFARX1 I_48629 (I829222,I2507,I829154,I829248,);
DFFARX1 I_48630 (I829248,I2507,I829154,I829143,);
DFFARX1 I_48631 (I1143339,I2507,I829154,I829279,);
nand I_48632 (I829287,I829279,I1143348);
not I_48633 (I829304,I829287);
DFFARX1 I_48634 (I829304,I2507,I829154,I829330,);
not I_48635 (I829338,I829330);
nor I_48636 (I829146,I829188,I829338);
DFFARX1 I_48637 (I1143360,I2507,I829154,I829378,);
nor I_48638 (I829137,I829378,I829248);
nor I_48639 (I829128,I829378,I829304);
nand I_48640 (I829414,I1143351,I1143345);
and I_48641 (I829431,I829414,I1143339);
DFFARX1 I_48642 (I829431,I2507,I829154,I829457,);
not I_48643 (I829465,I829457);
nand I_48644 (I829482,I829465,I829378);
nand I_48645 (I829131,I829465,I829287);
nor I_48646 (I829513,I1143357,I1143345);
and I_48647 (I829530,I829378,I829513);
nor I_48648 (I829547,I829465,I829530);
DFFARX1 I_48649 (I829547,I2507,I829154,I829140,);
nor I_48650 (I829578,I829180,I829513);
DFFARX1 I_48651 (I829578,I2507,I829154,I829125,);
nor I_48652 (I829609,I829457,I829513);
not I_48653 (I829626,I829609);
nand I_48654 (I829134,I829626,I829482);
not I_48655 (I829681,I2514);
DFFARX1 I_48656 (I1070526,I2507,I829681,I829707,);
not I_48657 (I829715,I829707);
nand I_48658 (I829732,I1070508,I1070508);
and I_48659 (I829749,I829732,I1070514);
DFFARX1 I_48660 (I829749,I2507,I829681,I829775,);
DFFARX1 I_48661 (I829775,I2507,I829681,I829670,);
DFFARX1 I_48662 (I1070511,I2507,I829681,I829806,);
nand I_48663 (I829814,I829806,I1070520);
not I_48664 (I829831,I829814);
DFFARX1 I_48665 (I829831,I2507,I829681,I829857,);
not I_48666 (I829865,I829857);
nor I_48667 (I829673,I829715,I829865);
DFFARX1 I_48668 (I1070532,I2507,I829681,I829905,);
nor I_48669 (I829664,I829905,I829775);
nor I_48670 (I829655,I829905,I829831);
nand I_48671 (I829941,I1070523,I1070517);
and I_48672 (I829958,I829941,I1070511);
DFFARX1 I_48673 (I829958,I2507,I829681,I829984,);
not I_48674 (I829992,I829984);
nand I_48675 (I830009,I829992,I829905);
nand I_48676 (I829658,I829992,I829814);
nor I_48677 (I830040,I1070529,I1070517);
and I_48678 (I830057,I829905,I830040);
nor I_48679 (I830074,I829992,I830057);
DFFARX1 I_48680 (I830074,I2507,I829681,I829667,);
nor I_48681 (I830105,I829707,I830040);
DFFARX1 I_48682 (I830105,I2507,I829681,I829652,);
nor I_48683 (I830136,I829984,I830040);
not I_48684 (I830153,I830136);
nand I_48685 (I829661,I830153,I830009);
not I_48686 (I830208,I2514);
DFFARX1 I_48687 (I1284250,I2507,I830208,I830234,);
not I_48688 (I830242,I830234);
nand I_48689 (I830259,I1284232,I1284235);
and I_48690 (I830276,I830259,I1284247);
DFFARX1 I_48691 (I830276,I2507,I830208,I830302,);
DFFARX1 I_48692 (I830302,I2507,I830208,I830197,);
DFFARX1 I_48693 (I1284256,I2507,I830208,I830333,);
nand I_48694 (I830341,I830333,I1284241);
not I_48695 (I830358,I830341);
DFFARX1 I_48696 (I830358,I2507,I830208,I830384,);
not I_48697 (I830392,I830384);
nor I_48698 (I830200,I830242,I830392);
DFFARX1 I_48699 (I1284253,I2507,I830208,I830432,);
nor I_48700 (I830191,I830432,I830302);
nor I_48701 (I830182,I830432,I830358);
nand I_48702 (I830468,I1284244,I1284238);
and I_48703 (I830485,I830468,I1284232);
DFFARX1 I_48704 (I830485,I2507,I830208,I830511,);
not I_48705 (I830519,I830511);
nand I_48706 (I830536,I830519,I830432);
nand I_48707 (I830185,I830519,I830341);
nor I_48708 (I830567,I1284235,I1284238);
and I_48709 (I830584,I830432,I830567);
nor I_48710 (I830601,I830519,I830584);
DFFARX1 I_48711 (I830601,I2507,I830208,I830194,);
nor I_48712 (I830632,I830234,I830567);
DFFARX1 I_48713 (I830632,I2507,I830208,I830179,);
nor I_48714 (I830663,I830511,I830567);
not I_48715 (I830680,I830663);
nand I_48716 (I830188,I830680,I830536);
not I_48717 (I830735,I2514);
DFFARX1 I_48718 (I1064746,I2507,I830735,I830761,);
not I_48719 (I830769,I830761);
nand I_48720 (I830786,I1064728,I1064728);
and I_48721 (I830803,I830786,I1064734);
DFFARX1 I_48722 (I830803,I2507,I830735,I830829,);
DFFARX1 I_48723 (I830829,I2507,I830735,I830724,);
DFFARX1 I_48724 (I1064731,I2507,I830735,I830860,);
nand I_48725 (I830868,I830860,I1064740);
not I_48726 (I830885,I830868);
DFFARX1 I_48727 (I830885,I2507,I830735,I830911,);
not I_48728 (I830919,I830911);
nor I_48729 (I830727,I830769,I830919);
DFFARX1 I_48730 (I1064752,I2507,I830735,I830959,);
nor I_48731 (I830718,I830959,I830829);
nor I_48732 (I830709,I830959,I830885);
nand I_48733 (I830995,I1064743,I1064737);
and I_48734 (I831012,I830995,I1064731);
DFFARX1 I_48735 (I831012,I2507,I830735,I831038,);
not I_48736 (I831046,I831038);
nand I_48737 (I831063,I831046,I830959);
nand I_48738 (I830712,I831046,I830868);
nor I_48739 (I831094,I1064749,I1064737);
and I_48740 (I831111,I830959,I831094);
nor I_48741 (I831128,I831046,I831111);
DFFARX1 I_48742 (I831128,I2507,I830735,I830721,);
nor I_48743 (I831159,I830761,I831094);
DFFARX1 I_48744 (I831159,I2507,I830735,I830706,);
nor I_48745 (I831190,I831038,I831094);
not I_48746 (I831207,I831190);
nand I_48747 (I830715,I831207,I831063);
not I_48748 (I831262,I2514);
DFFARX1 I_48749 (I649792,I2507,I831262,I831288,);
not I_48750 (I831296,I831288);
nand I_48751 (I831313,I649795,I649792);
and I_48752 (I831330,I831313,I649804);
DFFARX1 I_48753 (I831330,I2507,I831262,I831356,);
DFFARX1 I_48754 (I831356,I2507,I831262,I831251,);
DFFARX1 I_48755 (I649801,I2507,I831262,I831387,);
nand I_48756 (I831395,I831387,I649807);
not I_48757 (I831412,I831395);
DFFARX1 I_48758 (I831412,I2507,I831262,I831438,);
not I_48759 (I831446,I831438);
nor I_48760 (I831254,I831296,I831446);
DFFARX1 I_48761 (I649816,I2507,I831262,I831486,);
nor I_48762 (I831245,I831486,I831356);
nor I_48763 (I831236,I831486,I831412);
nand I_48764 (I831522,I649810,I649798);
and I_48765 (I831539,I831522,I649795);
DFFARX1 I_48766 (I831539,I2507,I831262,I831565,);
not I_48767 (I831573,I831565);
nand I_48768 (I831590,I831573,I831486);
nand I_48769 (I831239,I831573,I831395);
nor I_48770 (I831621,I649813,I649798);
and I_48771 (I831638,I831486,I831621);
nor I_48772 (I831655,I831573,I831638);
DFFARX1 I_48773 (I831655,I2507,I831262,I831248,);
nor I_48774 (I831686,I831288,I831621);
DFFARX1 I_48775 (I831686,I2507,I831262,I831233,);
nor I_48776 (I831717,I831565,I831621);
not I_48777 (I831734,I831717);
nand I_48778 (I831242,I831734,I831590);
not I_48779 (I831789,I2514);
DFFARX1 I_48780 (I898556,I2507,I831789,I831815,);
not I_48781 (I831823,I831815);
nand I_48782 (I831840,I898571,I898553);
and I_48783 (I831857,I831840,I898553);
DFFARX1 I_48784 (I831857,I2507,I831789,I831883,);
DFFARX1 I_48785 (I831883,I2507,I831789,I831778,);
DFFARX1 I_48786 (I898562,I2507,I831789,I831914,);
nand I_48787 (I831922,I831914,I898580);
not I_48788 (I831939,I831922);
DFFARX1 I_48789 (I831939,I2507,I831789,I831965,);
not I_48790 (I831973,I831965);
nor I_48791 (I831781,I831823,I831973);
DFFARX1 I_48792 (I898577,I2507,I831789,I832013,);
nor I_48793 (I831772,I832013,I831883);
nor I_48794 (I831763,I832013,I831939);
nand I_48795 (I832049,I898574,I898565);
and I_48796 (I832066,I832049,I898559);
DFFARX1 I_48797 (I832066,I2507,I831789,I832092,);
not I_48798 (I832100,I832092);
nand I_48799 (I832117,I832100,I832013);
nand I_48800 (I831766,I832100,I831922);
nor I_48801 (I832148,I898568,I898565);
and I_48802 (I832165,I832013,I832148);
nor I_48803 (I832182,I832100,I832165);
DFFARX1 I_48804 (I832182,I2507,I831789,I831775,);
nor I_48805 (I832213,I831815,I832148);
DFFARX1 I_48806 (I832213,I2507,I831789,I831760,);
nor I_48807 (I832244,I832092,I832148);
not I_48808 (I832261,I832244);
nand I_48809 (I831769,I832261,I832117);
not I_48810 (I832316,I2514);
DFFARX1 I_48811 (I328722,I2507,I832316,I832342,);
not I_48812 (I832350,I832342);
nand I_48813 (I832367,I328713,I328713);
and I_48814 (I832384,I832367,I328731);
DFFARX1 I_48815 (I832384,I2507,I832316,I832410,);
DFFARX1 I_48816 (I832410,I2507,I832316,I832305,);
DFFARX1 I_48817 (I328734,I2507,I832316,I832441,);
nand I_48818 (I832449,I832441,I328716);
not I_48819 (I832466,I832449);
DFFARX1 I_48820 (I832466,I2507,I832316,I832492,);
not I_48821 (I832500,I832492);
nor I_48822 (I832308,I832350,I832500);
DFFARX1 I_48823 (I328728,I2507,I832316,I832540,);
nor I_48824 (I832299,I832540,I832410);
nor I_48825 (I832290,I832540,I832466);
nand I_48826 (I832576,I328740,I328719);
and I_48827 (I832593,I832576,I328725);
DFFARX1 I_48828 (I832593,I2507,I832316,I832619,);
not I_48829 (I832627,I832619);
nand I_48830 (I832644,I832627,I832540);
nand I_48831 (I832293,I832627,I832449);
nor I_48832 (I832675,I328737,I328719);
and I_48833 (I832692,I832540,I832675);
nor I_48834 (I832709,I832627,I832692);
DFFARX1 I_48835 (I832709,I2507,I832316,I832302,);
nor I_48836 (I832740,I832342,I832675);
DFFARX1 I_48837 (I832740,I2507,I832316,I832287,);
nor I_48838 (I832771,I832619,I832675);
not I_48839 (I832788,I832771);
nand I_48840 (I832296,I832788,I832644);
not I_48841 (I832843,I2514);
DFFARX1 I_48842 (I570621,I2507,I832843,I832869,);
not I_48843 (I832877,I832869);
nand I_48844 (I832894,I570606,I570627);
and I_48845 (I832911,I832894,I570615);
DFFARX1 I_48846 (I832911,I2507,I832843,I832937,);
DFFARX1 I_48847 (I832937,I2507,I832843,I832832,);
DFFARX1 I_48848 (I570609,I2507,I832843,I832968,);
nand I_48849 (I832976,I832968,I570618);
not I_48850 (I832993,I832976);
DFFARX1 I_48851 (I832993,I2507,I832843,I833019,);
not I_48852 (I833027,I833019);
nor I_48853 (I832835,I832877,I833027);
DFFARX1 I_48854 (I570624,I2507,I832843,I833067,);
nor I_48855 (I832826,I833067,I832937);
nor I_48856 (I832817,I833067,I832993);
nand I_48857 (I833103,I570606,I570609);
and I_48858 (I833120,I833103,I570630);
DFFARX1 I_48859 (I833120,I2507,I832843,I833146,);
not I_48860 (I833154,I833146);
nand I_48861 (I833171,I833154,I833067);
nand I_48862 (I832820,I833154,I832976);
nor I_48863 (I833202,I570612,I570609);
and I_48864 (I833219,I833067,I833202);
nor I_48865 (I833236,I833154,I833219);
DFFARX1 I_48866 (I833236,I2507,I832843,I832829,);
nor I_48867 (I833267,I832869,I833202);
DFFARX1 I_48868 (I833267,I2507,I832843,I832814,);
nor I_48869 (I833298,I833146,I833202);
not I_48870 (I833315,I833298);
nand I_48871 (I832823,I833315,I833171);
not I_48872 (I833370,I2514);
DFFARX1 I_48873 (I1315442,I2507,I833370,I833396,);
not I_48874 (I833404,I833396);
nand I_48875 (I833421,I1315439,I1315448);
and I_48876 (I833438,I833421,I1315427);
DFFARX1 I_48877 (I833438,I2507,I833370,I833464,);
DFFARX1 I_48878 (I833464,I2507,I833370,I833359,);
DFFARX1 I_48879 (I1315430,I2507,I833370,I833495,);
nand I_48880 (I833503,I833495,I1315445);
not I_48881 (I833520,I833503);
DFFARX1 I_48882 (I833520,I2507,I833370,I833546,);
not I_48883 (I833554,I833546);
nor I_48884 (I833362,I833404,I833554);
DFFARX1 I_48885 (I1315451,I2507,I833370,I833594,);
nor I_48886 (I833353,I833594,I833464);
nor I_48887 (I833344,I833594,I833520);
nand I_48888 (I833630,I1315433,I1315454);
and I_48889 (I833647,I833630,I1315436);
DFFARX1 I_48890 (I833647,I2507,I833370,I833673,);
not I_48891 (I833681,I833673);
nand I_48892 (I833698,I833681,I833594);
nand I_48893 (I833347,I833681,I833503);
nor I_48894 (I833729,I1315427,I1315454);
and I_48895 (I833746,I833594,I833729);
nor I_48896 (I833763,I833681,I833746);
DFFARX1 I_48897 (I833763,I2507,I833370,I833356,);
nor I_48898 (I833794,I833396,I833729);
DFFARX1 I_48899 (I833794,I2507,I833370,I833341,);
nor I_48900 (I833825,I833673,I833729);
not I_48901 (I833842,I833825);
nand I_48902 (I833350,I833842,I833698);
not I_48903 (I833897,I2514);
DFFARX1 I_48904 (I1354117,I2507,I833897,I833923,);
not I_48905 (I833931,I833923);
nand I_48906 (I833948,I1354114,I1354123);
and I_48907 (I833965,I833948,I1354102);
DFFARX1 I_48908 (I833965,I2507,I833897,I833991,);
DFFARX1 I_48909 (I833991,I2507,I833897,I833886,);
DFFARX1 I_48910 (I1354105,I2507,I833897,I834022,);
nand I_48911 (I834030,I834022,I1354120);
not I_48912 (I834047,I834030);
DFFARX1 I_48913 (I834047,I2507,I833897,I834073,);
not I_48914 (I834081,I834073);
nor I_48915 (I833889,I833931,I834081);
DFFARX1 I_48916 (I1354126,I2507,I833897,I834121,);
nor I_48917 (I833880,I834121,I833991);
nor I_48918 (I833871,I834121,I834047);
nand I_48919 (I834157,I1354108,I1354129);
and I_48920 (I834174,I834157,I1354111);
DFFARX1 I_48921 (I834174,I2507,I833897,I834200,);
not I_48922 (I834208,I834200);
nand I_48923 (I834225,I834208,I834121);
nand I_48924 (I833874,I834208,I834030);
nor I_48925 (I834256,I1354102,I1354129);
and I_48926 (I834273,I834121,I834256);
nor I_48927 (I834290,I834208,I834273);
DFFARX1 I_48928 (I834290,I2507,I833897,I833883,);
nor I_48929 (I834321,I833923,I834256);
DFFARX1 I_48930 (I834321,I2507,I833897,I833868,);
nor I_48931 (I834352,I834200,I834256);
not I_48932 (I834369,I834352);
nand I_48933 (I833877,I834369,I834225);
not I_48934 (I834424,I2514);
DFFARX1 I_48935 (I243056,I2507,I834424,I834450,);
not I_48936 (I834458,I834450);
nand I_48937 (I834475,I243053,I243071);
and I_48938 (I834492,I834475,I243062);
DFFARX1 I_48939 (I834492,I2507,I834424,I834518,);
DFFARX1 I_48940 (I834518,I2507,I834424,I834413,);
DFFARX1 I_48941 (I243068,I2507,I834424,I834549,);
nand I_48942 (I834557,I834549,I243065);
not I_48943 (I834574,I834557);
DFFARX1 I_48944 (I834574,I2507,I834424,I834600,);
not I_48945 (I834608,I834600);
nor I_48946 (I834416,I834458,I834608);
DFFARX1 I_48947 (I243059,I2507,I834424,I834648,);
nor I_48948 (I834407,I834648,I834518);
nor I_48949 (I834398,I834648,I834574);
nand I_48950 (I834684,I243050,I243074);
and I_48951 (I834701,I834684,I243053);
DFFARX1 I_48952 (I834701,I2507,I834424,I834727,);
not I_48953 (I834735,I834727);
nand I_48954 (I834752,I834735,I834648);
nand I_48955 (I834401,I834735,I834557);
nor I_48956 (I834783,I243050,I243074);
and I_48957 (I834800,I834648,I834783);
nor I_48958 (I834817,I834735,I834800);
DFFARX1 I_48959 (I834817,I2507,I834424,I834410,);
nor I_48960 (I834848,I834450,I834783);
DFFARX1 I_48961 (I834848,I2507,I834424,I834395,);
nor I_48962 (I834879,I834727,I834783);
not I_48963 (I834896,I834879);
nand I_48964 (I834404,I834896,I834752);
not I_48965 (I834951,I2514);
DFFARX1 I_48966 (I1264020,I2507,I834951,I834977,);
not I_48967 (I834985,I834977);
nand I_48968 (I835002,I1264002,I1264005);
and I_48969 (I835019,I835002,I1264017);
DFFARX1 I_48970 (I835019,I2507,I834951,I835045,);
DFFARX1 I_48971 (I835045,I2507,I834951,I834940,);
DFFARX1 I_48972 (I1264026,I2507,I834951,I835076,);
nand I_48973 (I835084,I835076,I1264011);
not I_48974 (I835101,I835084);
DFFARX1 I_48975 (I835101,I2507,I834951,I835127,);
not I_48976 (I835135,I835127);
nor I_48977 (I834943,I834985,I835135);
DFFARX1 I_48978 (I1264023,I2507,I834951,I835175,);
nor I_48979 (I834934,I835175,I835045);
nor I_48980 (I834925,I835175,I835101);
nand I_48981 (I835211,I1264014,I1264008);
and I_48982 (I835228,I835211,I1264002);
DFFARX1 I_48983 (I835228,I2507,I834951,I835254,);
not I_48984 (I835262,I835254);
nand I_48985 (I835279,I835262,I835175);
nand I_48986 (I834928,I835262,I835084);
nor I_48987 (I835310,I1264005,I1264008);
and I_48988 (I835327,I835175,I835310);
nor I_48989 (I835344,I835262,I835327);
DFFARX1 I_48990 (I835344,I2507,I834951,I834937,);
nor I_48991 (I835375,I834977,I835310);
DFFARX1 I_48992 (I835375,I2507,I834951,I834922,);
nor I_48993 (I835406,I835254,I835310);
not I_48994 (I835423,I835406);
nand I_48995 (I834931,I835423,I835279);
not I_48996 (I835478,I2514);
DFFARX1 I_48997 (I177606,I2507,I835478,I835504,);
not I_48998 (I835512,I835504);
nand I_48999 (I835529,I177603,I177621);
and I_49000 (I835546,I835529,I177612);
DFFARX1 I_49001 (I835546,I2507,I835478,I835572,);
DFFARX1 I_49002 (I835572,I2507,I835478,I835467,);
DFFARX1 I_49003 (I177618,I2507,I835478,I835603,);
nand I_49004 (I835611,I835603,I177615);
not I_49005 (I835628,I835611);
DFFARX1 I_49006 (I835628,I2507,I835478,I835654,);
not I_49007 (I835662,I835654);
nor I_49008 (I835470,I835512,I835662);
DFFARX1 I_49009 (I177609,I2507,I835478,I835702,);
nor I_49010 (I835461,I835702,I835572);
nor I_49011 (I835452,I835702,I835628);
nand I_49012 (I835738,I177600,I177624);
and I_49013 (I835755,I835738,I177603);
DFFARX1 I_49014 (I835755,I2507,I835478,I835781,);
not I_49015 (I835789,I835781);
nand I_49016 (I835806,I835789,I835702);
nand I_49017 (I835455,I835789,I835611);
nor I_49018 (I835837,I177600,I177624);
and I_49019 (I835854,I835702,I835837);
nor I_49020 (I835871,I835789,I835854);
DFFARX1 I_49021 (I835871,I2507,I835478,I835464,);
nor I_49022 (I835902,I835504,I835837);
DFFARX1 I_49023 (I835902,I2507,I835478,I835449,);
nor I_49024 (I835933,I835781,I835837);
not I_49025 (I835950,I835933);
nand I_49026 (I835458,I835950,I835806);
not I_49027 (I836005,I2514);
DFFARX1 I_49028 (I1035395,I2507,I836005,I836031,);
not I_49029 (I836039,I836031);
nand I_49030 (I836056,I1035404,I1035392);
and I_49031 (I836073,I836056,I1035389);
DFFARX1 I_49032 (I836073,I2507,I836005,I836099,);
DFFARX1 I_49033 (I836099,I2507,I836005,I835994,);
DFFARX1 I_49034 (I1035389,I2507,I836005,I836130,);
nand I_49035 (I836138,I836130,I1035386);
not I_49036 (I836155,I836138);
DFFARX1 I_49037 (I836155,I2507,I836005,I836181,);
not I_49038 (I836189,I836181);
nor I_49039 (I835997,I836039,I836189);
DFFARX1 I_49040 (I1035392,I2507,I836005,I836229,);
nor I_49041 (I835988,I836229,I836099);
nor I_49042 (I835979,I836229,I836155);
nand I_49043 (I836265,I1035407,I1035398);
and I_49044 (I836282,I836265,I1035401);
DFFARX1 I_49045 (I836282,I2507,I836005,I836308,);
not I_49046 (I836316,I836308);
nand I_49047 (I836333,I836316,I836229);
nand I_49048 (I835982,I836316,I836138);
nor I_49049 (I836364,I1035386,I1035398);
and I_49050 (I836381,I836229,I836364);
nor I_49051 (I836398,I836316,I836381);
DFFARX1 I_49052 (I836398,I2507,I836005,I835991,);
nor I_49053 (I836429,I836031,I836364);
DFFARX1 I_49054 (I836429,I2507,I836005,I835976,);
nor I_49055 (I836460,I836308,I836364);
not I_49056 (I836477,I836460);
nand I_49057 (I835985,I836477,I836333);
not I_49058 (I836532,I2514);
DFFARX1 I_49059 (I367193,I2507,I836532,I836558,);
not I_49060 (I836566,I836558);
nand I_49061 (I836583,I367184,I367184);
and I_49062 (I836600,I836583,I367202);
DFFARX1 I_49063 (I836600,I2507,I836532,I836626,);
DFFARX1 I_49064 (I836626,I2507,I836532,I836521,);
DFFARX1 I_49065 (I367205,I2507,I836532,I836657,);
nand I_49066 (I836665,I836657,I367187);
not I_49067 (I836682,I836665);
DFFARX1 I_49068 (I836682,I2507,I836532,I836708,);
not I_49069 (I836716,I836708);
nor I_49070 (I836524,I836566,I836716);
DFFARX1 I_49071 (I367199,I2507,I836532,I836756,);
nor I_49072 (I836515,I836756,I836626);
nor I_49073 (I836506,I836756,I836682);
nand I_49074 (I836792,I367211,I367190);
and I_49075 (I836809,I836792,I367196);
DFFARX1 I_49076 (I836809,I2507,I836532,I836835,);
not I_49077 (I836843,I836835);
nand I_49078 (I836860,I836843,I836756);
nand I_49079 (I836509,I836843,I836665);
nor I_49080 (I836891,I367208,I367190);
and I_49081 (I836908,I836756,I836891);
nor I_49082 (I836925,I836843,I836908);
DFFARX1 I_49083 (I836925,I2507,I836532,I836518,);
nor I_49084 (I836956,I836558,I836891);
DFFARX1 I_49085 (I836956,I2507,I836532,I836503,);
nor I_49086 (I836987,I836835,I836891);
not I_49087 (I837004,I836987);
nand I_49088 (I836512,I837004,I836860);
not I_49089 (I837059,I2514);
DFFARX1 I_49090 (I921166,I2507,I837059,I837085,);
not I_49091 (I837093,I837085);
nand I_49092 (I837110,I921181,I921163);
and I_49093 (I837127,I837110,I921163);
DFFARX1 I_49094 (I837127,I2507,I837059,I837153,);
DFFARX1 I_49095 (I837153,I2507,I837059,I837048,);
DFFARX1 I_49096 (I921172,I2507,I837059,I837184,);
nand I_49097 (I837192,I837184,I921190);
not I_49098 (I837209,I837192);
DFFARX1 I_49099 (I837209,I2507,I837059,I837235,);
not I_49100 (I837243,I837235);
nor I_49101 (I837051,I837093,I837243);
DFFARX1 I_49102 (I921187,I2507,I837059,I837283,);
nor I_49103 (I837042,I837283,I837153);
nor I_49104 (I837033,I837283,I837209);
nand I_49105 (I837319,I921184,I921175);
and I_49106 (I837336,I837319,I921169);
DFFARX1 I_49107 (I837336,I2507,I837059,I837362,);
not I_49108 (I837370,I837362);
nand I_49109 (I837387,I837370,I837283);
nand I_49110 (I837036,I837370,I837192);
nor I_49111 (I837418,I921178,I921175);
and I_49112 (I837435,I837283,I837418);
nor I_49113 (I837452,I837370,I837435);
DFFARX1 I_49114 (I837452,I2507,I837059,I837045,);
nor I_49115 (I837483,I837085,I837418);
DFFARX1 I_49116 (I837483,I2507,I837059,I837030,);
nor I_49117 (I837514,I837362,I837418);
not I_49118 (I837531,I837514);
nand I_49119 (I837039,I837531,I837387);
not I_49120 (I837586,I2514);
DFFARX1 I_49121 (I311858,I2507,I837586,I837612,);
not I_49122 (I837620,I837612);
nand I_49123 (I837637,I311849,I311849);
and I_49124 (I837654,I837637,I311867);
DFFARX1 I_49125 (I837654,I2507,I837586,I837680,);
DFFARX1 I_49126 (I837680,I2507,I837586,I837575,);
DFFARX1 I_49127 (I311870,I2507,I837586,I837711,);
nand I_49128 (I837719,I837711,I311852);
not I_49129 (I837736,I837719);
DFFARX1 I_49130 (I837736,I2507,I837586,I837762,);
not I_49131 (I837770,I837762);
nor I_49132 (I837578,I837620,I837770);
DFFARX1 I_49133 (I311864,I2507,I837586,I837810,);
nor I_49134 (I837569,I837810,I837680);
nor I_49135 (I837560,I837810,I837736);
nand I_49136 (I837846,I311876,I311855);
and I_49137 (I837863,I837846,I311861);
DFFARX1 I_49138 (I837863,I2507,I837586,I837889,);
not I_49139 (I837897,I837889);
nand I_49140 (I837914,I837897,I837810);
nand I_49141 (I837563,I837897,I837719);
nor I_49142 (I837945,I311873,I311855);
and I_49143 (I837962,I837810,I837945);
nor I_49144 (I837979,I837897,I837962);
DFFARX1 I_49145 (I837979,I2507,I837586,I837572,);
nor I_49146 (I838010,I837612,I837945);
DFFARX1 I_49147 (I838010,I2507,I837586,I837557,);
nor I_49148 (I838041,I837889,I837945);
not I_49149 (I838058,I838041);
nand I_49150 (I837566,I838058,I837914);
not I_49151 (I838113,I2514);
DFFARX1 I_49152 (I302899,I2507,I838113,I838139,);
not I_49153 (I838147,I838139);
nand I_49154 (I838164,I302890,I302890);
and I_49155 (I838181,I838164,I302908);
DFFARX1 I_49156 (I838181,I2507,I838113,I838207,);
DFFARX1 I_49157 (I838207,I2507,I838113,I838102,);
DFFARX1 I_49158 (I302911,I2507,I838113,I838238,);
nand I_49159 (I838246,I838238,I302893);
not I_49160 (I838263,I838246);
DFFARX1 I_49161 (I838263,I2507,I838113,I838289,);
not I_49162 (I838297,I838289);
nor I_49163 (I838105,I838147,I838297);
DFFARX1 I_49164 (I302905,I2507,I838113,I838337,);
nor I_49165 (I838096,I838337,I838207);
nor I_49166 (I838087,I838337,I838263);
nand I_49167 (I838373,I302917,I302896);
and I_49168 (I838390,I838373,I302902);
DFFARX1 I_49169 (I838390,I2507,I838113,I838416,);
not I_49170 (I838424,I838416);
nand I_49171 (I838441,I838424,I838337);
nand I_49172 (I838090,I838424,I838246);
nor I_49173 (I838472,I302914,I302896);
and I_49174 (I838489,I838337,I838472);
nor I_49175 (I838506,I838424,I838489);
DFFARX1 I_49176 (I838506,I2507,I838113,I838099,);
nor I_49177 (I838537,I838139,I838472);
DFFARX1 I_49178 (I838537,I2507,I838113,I838084,);
nor I_49179 (I838568,I838416,I838472);
not I_49180 (I838585,I838568);
nand I_49181 (I838093,I838585,I838441);
not I_49182 (I838640,I2514);
DFFARX1 I_49183 (I722620,I2507,I838640,I838666,);
not I_49184 (I838674,I838666);
nand I_49185 (I838691,I722623,I722620);
and I_49186 (I838708,I838691,I722632);
DFFARX1 I_49187 (I838708,I2507,I838640,I838734,);
DFFARX1 I_49188 (I838734,I2507,I838640,I838629,);
DFFARX1 I_49189 (I722629,I2507,I838640,I838765,);
nand I_49190 (I838773,I838765,I722635);
not I_49191 (I838790,I838773);
DFFARX1 I_49192 (I838790,I2507,I838640,I838816,);
not I_49193 (I838824,I838816);
nor I_49194 (I838632,I838674,I838824);
DFFARX1 I_49195 (I722644,I2507,I838640,I838864,);
nor I_49196 (I838623,I838864,I838734);
nor I_49197 (I838614,I838864,I838790);
nand I_49198 (I838900,I722638,I722626);
and I_49199 (I838917,I838900,I722623);
DFFARX1 I_49200 (I838917,I2507,I838640,I838943,);
not I_49201 (I838951,I838943);
nand I_49202 (I838968,I838951,I838864);
nand I_49203 (I838617,I838951,I838773);
nor I_49204 (I838999,I722641,I722626);
and I_49205 (I839016,I838864,I838999);
nor I_49206 (I839033,I838951,I839016);
DFFARX1 I_49207 (I839033,I2507,I838640,I838626,);
nor I_49208 (I839064,I838666,I838999);
DFFARX1 I_49209 (I839064,I2507,I838640,I838611,);
nor I_49210 (I839095,I838943,I838999);
not I_49211 (I839112,I839095);
nand I_49212 (I838620,I839112,I838968);
not I_49213 (I839167,I2514);
DFFARX1 I_49214 (I1392197,I2507,I839167,I839193,);
not I_49215 (I839201,I839193);
nand I_49216 (I839218,I1392194,I1392203);
and I_49217 (I839235,I839218,I1392182);
DFFARX1 I_49218 (I839235,I2507,I839167,I839261,);
DFFARX1 I_49219 (I839261,I2507,I839167,I839156,);
DFFARX1 I_49220 (I1392185,I2507,I839167,I839292,);
nand I_49221 (I839300,I839292,I1392200);
not I_49222 (I839317,I839300);
DFFARX1 I_49223 (I839317,I2507,I839167,I839343,);
not I_49224 (I839351,I839343);
nor I_49225 (I839159,I839201,I839351);
DFFARX1 I_49226 (I1392206,I2507,I839167,I839391,);
nor I_49227 (I839150,I839391,I839261);
nor I_49228 (I839141,I839391,I839317);
nand I_49229 (I839427,I1392188,I1392209);
and I_49230 (I839444,I839427,I1392191);
DFFARX1 I_49231 (I839444,I2507,I839167,I839470,);
not I_49232 (I839478,I839470);
nand I_49233 (I839495,I839478,I839391);
nand I_49234 (I839144,I839478,I839300);
nor I_49235 (I839526,I1392182,I1392209);
and I_49236 (I839543,I839391,I839526);
nor I_49237 (I839560,I839478,I839543);
DFFARX1 I_49238 (I839560,I2507,I839167,I839153,);
nor I_49239 (I839591,I839193,I839526);
DFFARX1 I_49240 (I839591,I2507,I839167,I839138,);
nor I_49241 (I839622,I839470,I839526);
not I_49242 (I839639,I839622);
nand I_49243 (I839147,I839639,I839495);
not I_49244 (I839694,I2514);
DFFARX1 I_49245 (I279184,I2507,I839694,I839720,);
not I_49246 (I839728,I839720);
nand I_49247 (I839745,I279175,I279175);
and I_49248 (I839762,I839745,I279193);
DFFARX1 I_49249 (I839762,I2507,I839694,I839788,);
DFFARX1 I_49250 (I839788,I2507,I839694,I839683,);
DFFARX1 I_49251 (I279196,I2507,I839694,I839819,);
nand I_49252 (I839827,I839819,I279178);
not I_49253 (I839844,I839827);
DFFARX1 I_49254 (I839844,I2507,I839694,I839870,);
not I_49255 (I839878,I839870);
nor I_49256 (I839686,I839728,I839878);
DFFARX1 I_49257 (I279190,I2507,I839694,I839918,);
nor I_49258 (I839677,I839918,I839788);
nor I_49259 (I839668,I839918,I839844);
nand I_49260 (I839954,I279202,I279181);
and I_49261 (I839971,I839954,I279187);
DFFARX1 I_49262 (I839971,I2507,I839694,I839997,);
not I_49263 (I840005,I839997);
nand I_49264 (I840022,I840005,I839918);
nand I_49265 (I839671,I840005,I839827);
nor I_49266 (I840053,I279199,I279181);
and I_49267 (I840070,I839918,I840053);
nor I_49268 (I840087,I840005,I840070);
DFFARX1 I_49269 (I840087,I2507,I839694,I839680,);
nor I_49270 (I840118,I839720,I840053);
DFFARX1 I_49271 (I840118,I2507,I839694,I839665,);
nor I_49272 (I840149,I839997,I840053);
not I_49273 (I840166,I840149);
nand I_49274 (I839674,I840166,I840022);
not I_49275 (I840221,I2514);
DFFARX1 I_49276 (I313439,I2507,I840221,I840247,);
not I_49277 (I840255,I840247);
nand I_49278 (I840272,I313430,I313430);
and I_49279 (I840289,I840272,I313448);
DFFARX1 I_49280 (I840289,I2507,I840221,I840315,);
DFFARX1 I_49281 (I840315,I2507,I840221,I840210,);
DFFARX1 I_49282 (I313451,I2507,I840221,I840346,);
nand I_49283 (I840354,I840346,I313433);
not I_49284 (I840371,I840354);
DFFARX1 I_49285 (I840371,I2507,I840221,I840397,);
not I_49286 (I840405,I840397);
nor I_49287 (I840213,I840255,I840405);
DFFARX1 I_49288 (I313445,I2507,I840221,I840445,);
nor I_49289 (I840204,I840445,I840315);
nor I_49290 (I840195,I840445,I840371);
nand I_49291 (I840481,I313457,I313436);
and I_49292 (I840498,I840481,I313442);
DFFARX1 I_49293 (I840498,I2507,I840221,I840524,);
not I_49294 (I840532,I840524);
nand I_49295 (I840549,I840532,I840445);
nand I_49296 (I840198,I840532,I840354);
nor I_49297 (I840580,I313454,I313436);
and I_49298 (I840597,I840445,I840580);
nor I_49299 (I840614,I840532,I840597);
DFFARX1 I_49300 (I840614,I2507,I840221,I840207,);
nor I_49301 (I840645,I840247,I840580);
DFFARX1 I_49302 (I840645,I2507,I840221,I840192,);
nor I_49303 (I840676,I840524,I840580);
not I_49304 (I840693,I840676);
nand I_49305 (I840201,I840693,I840549);
not I_49306 (I840748,I2514);
DFFARX1 I_49307 (I1350547,I2507,I840748,I840774,);
not I_49308 (I840782,I840774);
nand I_49309 (I840799,I1350544,I1350553);
and I_49310 (I840816,I840799,I1350532);
DFFARX1 I_49311 (I840816,I2507,I840748,I840842,);
DFFARX1 I_49312 (I840842,I2507,I840748,I840737,);
DFFARX1 I_49313 (I1350535,I2507,I840748,I840873,);
nand I_49314 (I840881,I840873,I1350550);
not I_49315 (I840898,I840881);
DFFARX1 I_49316 (I840898,I2507,I840748,I840924,);
not I_49317 (I840932,I840924);
nor I_49318 (I840740,I840782,I840932);
DFFARX1 I_49319 (I1350556,I2507,I840748,I840972,);
nor I_49320 (I840731,I840972,I840842);
nor I_49321 (I840722,I840972,I840898);
nand I_49322 (I841008,I1350538,I1350559);
and I_49323 (I841025,I841008,I1350541);
DFFARX1 I_49324 (I841025,I2507,I840748,I841051,);
not I_49325 (I841059,I841051);
nand I_49326 (I841076,I841059,I840972);
nand I_49327 (I840725,I841059,I840881);
nor I_49328 (I841107,I1350532,I1350559);
and I_49329 (I841124,I840972,I841107);
nor I_49330 (I841141,I841059,I841124);
DFFARX1 I_49331 (I841141,I2507,I840748,I840734,);
nor I_49332 (I841172,I840774,I841107);
DFFARX1 I_49333 (I841172,I2507,I840748,I840719,);
nor I_49334 (I841203,I841051,I841107);
not I_49335 (I841220,I841203);
nand I_49336 (I840728,I841220,I841076);
not I_49337 (I841275,I2514);
DFFARX1 I_49338 (I76491,I2507,I841275,I841301,);
not I_49339 (I841309,I841301);
nand I_49340 (I841326,I76467,I76476);
and I_49341 (I841343,I841326,I76470);
DFFARX1 I_49342 (I841343,I2507,I841275,I841369,);
DFFARX1 I_49343 (I841369,I2507,I841275,I841264,);
DFFARX1 I_49344 (I76488,I2507,I841275,I841400,);
nand I_49345 (I841408,I841400,I76479);
not I_49346 (I841425,I841408);
DFFARX1 I_49347 (I841425,I2507,I841275,I841451,);
not I_49348 (I841459,I841451);
nor I_49349 (I841267,I841309,I841459);
DFFARX1 I_49350 (I76473,I2507,I841275,I841499,);
nor I_49351 (I841258,I841499,I841369);
nor I_49352 (I841249,I841499,I841425);
nand I_49353 (I841535,I76485,I76482);
and I_49354 (I841552,I841535,I76470);
DFFARX1 I_49355 (I841552,I2507,I841275,I841578,);
not I_49356 (I841586,I841578);
nand I_49357 (I841603,I841586,I841499);
nand I_49358 (I841252,I841586,I841408);
nor I_49359 (I841634,I76467,I76482);
and I_49360 (I841651,I841499,I841634);
nor I_49361 (I841668,I841586,I841651);
DFFARX1 I_49362 (I841668,I2507,I841275,I841261,);
nor I_49363 (I841699,I841301,I841634);
DFFARX1 I_49364 (I841699,I2507,I841275,I841246,);
nor I_49365 (I841730,I841578,I841634);
not I_49366 (I841747,I841730);
nand I_49367 (I841255,I841747,I841603);
not I_49368 (I841802,I2514);
DFFARX1 I_49369 (I172251,I2507,I841802,I841828,);
not I_49370 (I841836,I841828);
nand I_49371 (I841853,I172248,I172266);
and I_49372 (I841870,I841853,I172257);
DFFARX1 I_49373 (I841870,I2507,I841802,I841896,);
DFFARX1 I_49374 (I841896,I2507,I841802,I841791,);
DFFARX1 I_49375 (I172263,I2507,I841802,I841927,);
nand I_49376 (I841935,I841927,I172260);
not I_49377 (I841952,I841935);
DFFARX1 I_49378 (I841952,I2507,I841802,I841978,);
not I_49379 (I841986,I841978);
nor I_49380 (I841794,I841836,I841986);
DFFARX1 I_49381 (I172254,I2507,I841802,I842026,);
nor I_49382 (I841785,I842026,I841896);
nor I_49383 (I841776,I842026,I841952);
nand I_49384 (I842062,I172245,I172269);
and I_49385 (I842079,I842062,I172248);
DFFARX1 I_49386 (I842079,I2507,I841802,I842105,);
not I_49387 (I842113,I842105);
nand I_49388 (I842130,I842113,I842026);
nand I_49389 (I841779,I842113,I841935);
nor I_49390 (I842161,I172245,I172269);
and I_49391 (I842178,I842026,I842161);
nor I_49392 (I842195,I842113,I842178);
DFFARX1 I_49393 (I842195,I2507,I841802,I841788,);
nor I_49394 (I842226,I841828,I842161);
DFFARX1 I_49395 (I842226,I2507,I841802,I841773,);
nor I_49396 (I842257,I842105,I842161);
not I_49397 (I842274,I842257);
nand I_49398 (I841782,I842274,I842130);
not I_49399 (I842329,I2514);
DFFARX1 I_49400 (I1219406,I2507,I842329,I842355,);
not I_49401 (I842363,I842355);
nand I_49402 (I842380,I1219412,I1219394);
and I_49403 (I842397,I842380,I1219403);
DFFARX1 I_49404 (I842397,I2507,I842329,I842423,);
DFFARX1 I_49405 (I842423,I2507,I842329,I842318,);
DFFARX1 I_49406 (I1219409,I2507,I842329,I842454,);
nand I_49407 (I842462,I842454,I1219397);
not I_49408 (I842479,I842462);
DFFARX1 I_49409 (I842479,I2507,I842329,I842505,);
not I_49410 (I842513,I842505);
nor I_49411 (I842321,I842363,I842513);
DFFARX1 I_49412 (I1219415,I2507,I842329,I842553,);
nor I_49413 (I842312,I842553,I842423);
nor I_49414 (I842303,I842553,I842479);
nand I_49415 (I842589,I1219394,I1219400);
and I_49416 (I842606,I842589,I1219418);
DFFARX1 I_49417 (I842606,I2507,I842329,I842632,);
not I_49418 (I842640,I842632);
nand I_49419 (I842657,I842640,I842553);
nand I_49420 (I842306,I842640,I842462);
nor I_49421 (I842688,I1219397,I1219400);
and I_49422 (I842705,I842553,I842688);
nor I_49423 (I842722,I842640,I842705);
DFFARX1 I_49424 (I842722,I2507,I842329,I842315,);
nor I_49425 (I842753,I842355,I842688);
DFFARX1 I_49426 (I842753,I2507,I842329,I842300,);
nor I_49427 (I842784,I842632,I842688);
not I_49428 (I842801,I842784);
nand I_49429 (I842309,I842801,I842657);
not I_49430 (I842856,I2514);
DFFARX1 I_49431 (I455029,I2507,I842856,I842882,);
not I_49432 (I842890,I842882);
nand I_49433 (I842907,I455026,I455035);
and I_49434 (I842924,I842907,I455044);
DFFARX1 I_49435 (I842924,I2507,I842856,I842950,);
DFFARX1 I_49436 (I842950,I2507,I842856,I842845,);
DFFARX1 I_49437 (I455047,I2507,I842856,I842981,);
nand I_49438 (I842989,I842981,I455050);
not I_49439 (I843006,I842989);
DFFARX1 I_49440 (I843006,I2507,I842856,I843032,);
not I_49441 (I843040,I843032);
nor I_49442 (I842848,I842890,I843040);
DFFARX1 I_49443 (I455023,I2507,I842856,I843080,);
nor I_49444 (I842839,I843080,I842950);
nor I_49445 (I842830,I843080,I843006);
nand I_49446 (I843116,I455038,I455041);
and I_49447 (I843133,I843116,I455032);
DFFARX1 I_49448 (I843133,I2507,I842856,I843159,);
not I_49449 (I843167,I843159);
nand I_49450 (I843184,I843167,I843080);
nand I_49451 (I842833,I843167,I842989);
nor I_49452 (I843215,I455023,I455041);
and I_49453 (I843232,I843080,I843215);
nor I_49454 (I843249,I843167,I843232);
DFFARX1 I_49455 (I843249,I2507,I842856,I842842,);
nor I_49456 (I843280,I842882,I843215);
DFFARX1 I_49457 (I843280,I2507,I842856,I842827,);
nor I_49458 (I843311,I843159,I843215);
not I_49459 (I843328,I843311);
nand I_49460 (I842836,I843328,I843184);
not I_49461 (I843383,I2514);
DFFARX1 I_49462 (I255996,I2507,I843383,I843409,);
not I_49463 (I843417,I843409);
nand I_49464 (I843434,I255987,I255987);
and I_49465 (I843451,I843434,I256005);
DFFARX1 I_49466 (I843451,I2507,I843383,I843477,);
DFFARX1 I_49467 (I843477,I2507,I843383,I843372,);
DFFARX1 I_49468 (I256008,I2507,I843383,I843508,);
nand I_49469 (I843516,I843508,I255990);
not I_49470 (I843533,I843516);
DFFARX1 I_49471 (I843533,I2507,I843383,I843559,);
not I_49472 (I843567,I843559);
nor I_49473 (I843375,I843417,I843567);
DFFARX1 I_49474 (I256002,I2507,I843383,I843607,);
nor I_49475 (I843366,I843607,I843477);
nor I_49476 (I843357,I843607,I843533);
nand I_49477 (I843643,I256014,I255993);
and I_49478 (I843660,I843643,I255999);
DFFARX1 I_49479 (I843660,I2507,I843383,I843686,);
not I_49480 (I843694,I843686);
nand I_49481 (I843711,I843694,I843607);
nand I_49482 (I843360,I843694,I843516);
nor I_49483 (I843742,I256011,I255993);
and I_49484 (I843759,I843607,I843742);
nor I_49485 (I843776,I843694,I843759);
DFFARX1 I_49486 (I843776,I2507,I843383,I843369,);
nor I_49487 (I843807,I843409,I843742);
DFFARX1 I_49488 (I843807,I2507,I843383,I843354,);
nor I_49489 (I843838,I843686,I843742);
not I_49490 (I843855,I843838);
nand I_49491 (I843363,I843855,I843711);
not I_49492 (I843910,I2514);
DFFARX1 I_49493 (I1049420,I2507,I843910,I843936,);
not I_49494 (I843944,I843936);
nand I_49495 (I843961,I1049429,I1049417);
and I_49496 (I843978,I843961,I1049414);
DFFARX1 I_49497 (I843978,I2507,I843910,I844004,);
DFFARX1 I_49498 (I844004,I2507,I843910,I843899,);
DFFARX1 I_49499 (I1049414,I2507,I843910,I844035,);
nand I_49500 (I844043,I844035,I1049411);
not I_49501 (I844060,I844043);
DFFARX1 I_49502 (I844060,I2507,I843910,I844086,);
not I_49503 (I844094,I844086);
nor I_49504 (I843902,I843944,I844094);
DFFARX1 I_49505 (I1049417,I2507,I843910,I844134,);
nor I_49506 (I843893,I844134,I844004);
nor I_49507 (I843884,I844134,I844060);
nand I_49508 (I844170,I1049432,I1049423);
and I_49509 (I844187,I844170,I1049426);
DFFARX1 I_49510 (I844187,I2507,I843910,I844213,);
not I_49511 (I844221,I844213);
nand I_49512 (I844238,I844221,I844134);
nand I_49513 (I843887,I844221,I844043);
nor I_49514 (I844269,I1049411,I1049423);
and I_49515 (I844286,I844134,I844269);
nor I_49516 (I844303,I844221,I844286);
DFFARX1 I_49517 (I844303,I2507,I843910,I843896,);
nor I_49518 (I844334,I843936,I844269);
DFFARX1 I_49519 (I844334,I2507,I843910,I843881,);
nor I_49520 (I844365,I844213,I844269);
not I_49521 (I844382,I844365);
nand I_49522 (I843890,I844382,I844238);
not I_49523 (I844437,I2514);
DFFARX1 I_49524 (I19560,I2507,I844437,I844463,);
not I_49525 (I844471,I844463);
nand I_49526 (I844488,I19572,I19575);
and I_49527 (I844505,I844488,I19551);
DFFARX1 I_49528 (I844505,I2507,I844437,I844531,);
DFFARX1 I_49529 (I844531,I2507,I844437,I844426,);
DFFARX1 I_49530 (I19569,I2507,I844437,I844562,);
nand I_49531 (I844570,I844562,I19557);
not I_49532 (I844587,I844570);
DFFARX1 I_49533 (I844587,I2507,I844437,I844613,);
not I_49534 (I844621,I844613);
nor I_49535 (I844429,I844471,I844621);
DFFARX1 I_49536 (I19554,I2507,I844437,I844661,);
nor I_49537 (I844420,I844661,I844531);
nor I_49538 (I844411,I844661,I844587);
nand I_49539 (I844697,I19563,I19554);
and I_49540 (I844714,I844697,I19551);
DFFARX1 I_49541 (I844714,I2507,I844437,I844740,);
not I_49542 (I844748,I844740);
nand I_49543 (I844765,I844748,I844661);
nand I_49544 (I844414,I844748,I844570);
nor I_49545 (I844796,I19566,I19554);
and I_49546 (I844813,I844661,I844796);
nor I_49547 (I844830,I844748,I844813);
DFFARX1 I_49548 (I844830,I2507,I844437,I844423,);
nor I_49549 (I844861,I844463,I844796);
DFFARX1 I_49550 (I844861,I2507,I844437,I844408,);
nor I_49551 (I844892,I844740,I844796);
not I_49552 (I844909,I844892);
nand I_49553 (I844417,I844909,I844765);
not I_49554 (I844964,I2514);
DFFARX1 I_49555 (I681582,I2507,I844964,I844990,);
not I_49556 (I844998,I844990);
nand I_49557 (I845015,I681585,I681582);
and I_49558 (I845032,I845015,I681594);
DFFARX1 I_49559 (I845032,I2507,I844964,I845058,);
DFFARX1 I_49560 (I845058,I2507,I844964,I844953,);
DFFARX1 I_49561 (I681591,I2507,I844964,I845089,);
nand I_49562 (I845097,I845089,I681597);
not I_49563 (I845114,I845097);
DFFARX1 I_49564 (I845114,I2507,I844964,I845140,);
not I_49565 (I845148,I845140);
nor I_49566 (I844956,I844998,I845148);
DFFARX1 I_49567 (I681606,I2507,I844964,I845188,);
nor I_49568 (I844947,I845188,I845058);
nor I_49569 (I844938,I845188,I845114);
nand I_49570 (I845224,I681600,I681588);
and I_49571 (I845241,I845224,I681585);
DFFARX1 I_49572 (I845241,I2507,I844964,I845267,);
not I_49573 (I845275,I845267);
nand I_49574 (I845292,I845275,I845188);
nand I_49575 (I844941,I845275,I845097);
nor I_49576 (I845323,I681603,I681588);
and I_49577 (I845340,I845188,I845323);
nor I_49578 (I845357,I845275,I845340);
DFFARX1 I_49579 (I845357,I2507,I844964,I844950,);
nor I_49580 (I845388,I844990,I845323);
DFFARX1 I_49581 (I845388,I2507,I844964,I844935,);
nor I_49582 (I845419,I845267,I845323);
not I_49583 (I845436,I845419);
nand I_49584 (I844944,I845436,I845292);
not I_49585 (I845491,I2514);
DFFARX1 I_49586 (I363504,I2507,I845491,I845517,);
not I_49587 (I845525,I845517);
nand I_49588 (I845542,I363495,I363495);
and I_49589 (I845559,I845542,I363513);
DFFARX1 I_49590 (I845559,I2507,I845491,I845585,);
DFFARX1 I_49591 (I845585,I2507,I845491,I845480,);
DFFARX1 I_49592 (I363516,I2507,I845491,I845616,);
nand I_49593 (I845624,I845616,I363498);
not I_49594 (I845641,I845624);
DFFARX1 I_49595 (I845641,I2507,I845491,I845667,);
not I_49596 (I845675,I845667);
nor I_49597 (I845483,I845525,I845675);
DFFARX1 I_49598 (I363510,I2507,I845491,I845715,);
nor I_49599 (I845474,I845715,I845585);
nor I_49600 (I845465,I845715,I845641);
nand I_49601 (I845751,I363522,I363501);
and I_49602 (I845768,I845751,I363507);
DFFARX1 I_49603 (I845768,I2507,I845491,I845794,);
not I_49604 (I845802,I845794);
nand I_49605 (I845819,I845802,I845715);
nand I_49606 (I845468,I845802,I845624);
nor I_49607 (I845850,I363519,I363501);
and I_49608 (I845867,I845715,I845850);
nor I_49609 (I845884,I845802,I845867);
DFFARX1 I_49610 (I845884,I2507,I845491,I845477,);
nor I_49611 (I845915,I845517,I845850);
DFFARX1 I_49612 (I845915,I2507,I845491,I845462,);
nor I_49613 (I845946,I845794,I845850);
not I_49614 (I845963,I845946);
nand I_49615 (I845471,I845963,I845819);
not I_49616 (I846018,I2514);
DFFARX1 I_49617 (I1279626,I2507,I846018,I846044,);
not I_49618 (I846052,I846044);
nand I_49619 (I846069,I1279608,I1279611);
and I_49620 (I846086,I846069,I1279623);
DFFARX1 I_49621 (I846086,I2507,I846018,I846112,);
DFFARX1 I_49622 (I846112,I2507,I846018,I846007,);
DFFARX1 I_49623 (I1279632,I2507,I846018,I846143,);
nand I_49624 (I846151,I846143,I1279617);
not I_49625 (I846168,I846151);
DFFARX1 I_49626 (I846168,I2507,I846018,I846194,);
not I_49627 (I846202,I846194);
nor I_49628 (I846010,I846052,I846202);
DFFARX1 I_49629 (I1279629,I2507,I846018,I846242,);
nor I_49630 (I846001,I846242,I846112);
nor I_49631 (I845992,I846242,I846168);
nand I_49632 (I846278,I1279620,I1279614);
and I_49633 (I846295,I846278,I1279608);
DFFARX1 I_49634 (I846295,I2507,I846018,I846321,);
not I_49635 (I846329,I846321);
nand I_49636 (I846346,I846329,I846242);
nand I_49637 (I845995,I846329,I846151);
nor I_49638 (I846377,I1279611,I1279614);
and I_49639 (I846394,I846242,I846377);
nor I_49640 (I846411,I846329,I846394);
DFFARX1 I_49641 (I846411,I2507,I846018,I846004,);
nor I_49642 (I846442,I846044,I846377);
DFFARX1 I_49643 (I846442,I2507,I846018,I845989,);
nor I_49644 (I846473,I846321,I846377);
not I_49645 (I846490,I846473);
nand I_49646 (I845998,I846490,I846346);
not I_49647 (I846545,I2514);
DFFARX1 I_49648 (I720886,I2507,I846545,I846571,);
not I_49649 (I846579,I846571);
nand I_49650 (I846596,I720889,I720886);
and I_49651 (I846613,I846596,I720898);
DFFARX1 I_49652 (I846613,I2507,I846545,I846639,);
DFFARX1 I_49653 (I846639,I2507,I846545,I846534,);
DFFARX1 I_49654 (I720895,I2507,I846545,I846670,);
nand I_49655 (I846678,I846670,I720901);
not I_49656 (I846695,I846678);
DFFARX1 I_49657 (I846695,I2507,I846545,I846721,);
not I_49658 (I846729,I846721);
nor I_49659 (I846537,I846579,I846729);
DFFARX1 I_49660 (I720910,I2507,I846545,I846769,);
nor I_49661 (I846528,I846769,I846639);
nor I_49662 (I846519,I846769,I846695);
nand I_49663 (I846805,I720904,I720892);
and I_49664 (I846822,I846805,I720889);
DFFARX1 I_49665 (I846822,I2507,I846545,I846848,);
not I_49666 (I846856,I846848);
nand I_49667 (I846873,I846856,I846769);
nand I_49668 (I846522,I846856,I846678);
nor I_49669 (I846904,I720907,I720892);
and I_49670 (I846921,I846769,I846904);
nor I_49671 (I846938,I846856,I846921);
DFFARX1 I_49672 (I846938,I2507,I846545,I846531,);
nor I_49673 (I846969,I846571,I846904);
DFFARX1 I_49674 (I846969,I2507,I846545,I846516,);
nor I_49675 (I847000,I846848,I846904);
not I_49676 (I847017,I847000);
nand I_49677 (I846525,I847017,I846873);
not I_49678 (I847072,I2514);
DFFARX1 I_49679 (I271806,I2507,I847072,I847098,);
not I_49680 (I847106,I847098);
nand I_49681 (I847123,I271797,I271797);
and I_49682 (I847140,I847123,I271815);
DFFARX1 I_49683 (I847140,I2507,I847072,I847166,);
DFFARX1 I_49684 (I847166,I2507,I847072,I847061,);
DFFARX1 I_49685 (I271818,I2507,I847072,I847197,);
nand I_49686 (I847205,I847197,I271800);
not I_49687 (I847222,I847205);
DFFARX1 I_49688 (I847222,I2507,I847072,I847248,);
not I_49689 (I847256,I847248);
nor I_49690 (I847064,I847106,I847256);
DFFARX1 I_49691 (I271812,I2507,I847072,I847296,);
nor I_49692 (I847055,I847296,I847166);
nor I_49693 (I847046,I847296,I847222);
nand I_49694 (I847332,I271824,I271803);
and I_49695 (I847349,I847332,I271809);
DFFARX1 I_49696 (I847349,I2507,I847072,I847375,);
not I_49697 (I847383,I847375);
nand I_49698 (I847400,I847383,I847296);
nand I_49699 (I847049,I847383,I847205);
nor I_49700 (I847431,I271821,I271803);
and I_49701 (I847448,I847296,I847431);
nor I_49702 (I847465,I847383,I847448);
DFFARX1 I_49703 (I847465,I2507,I847072,I847058,);
nor I_49704 (I847496,I847098,I847431);
DFFARX1 I_49705 (I847496,I2507,I847072,I847043,);
nor I_49706 (I847527,I847375,I847431);
not I_49707 (I847544,I847527);
nand I_49708 (I847052,I847544,I847400);
not I_49709 (I847599,I2514);
DFFARX1 I_49710 (I471349,I2507,I847599,I847625,);
not I_49711 (I847633,I847625);
nand I_49712 (I847650,I471346,I471355);
and I_49713 (I847667,I847650,I471364);
DFFARX1 I_49714 (I847667,I2507,I847599,I847693,);
DFFARX1 I_49715 (I847693,I2507,I847599,I847588,);
DFFARX1 I_49716 (I471367,I2507,I847599,I847724,);
nand I_49717 (I847732,I847724,I471370);
not I_49718 (I847749,I847732);
DFFARX1 I_49719 (I847749,I2507,I847599,I847775,);
not I_49720 (I847783,I847775);
nor I_49721 (I847591,I847633,I847783);
DFFARX1 I_49722 (I471343,I2507,I847599,I847823,);
nor I_49723 (I847582,I847823,I847693);
nor I_49724 (I847573,I847823,I847749);
nand I_49725 (I847859,I471358,I471361);
and I_49726 (I847876,I847859,I471352);
DFFARX1 I_49727 (I847876,I2507,I847599,I847902,);
not I_49728 (I847910,I847902);
nand I_49729 (I847927,I847910,I847823);
nand I_49730 (I847576,I847910,I847732);
nor I_49731 (I847958,I471343,I471361);
and I_49732 (I847975,I847823,I847958);
nor I_49733 (I847992,I847910,I847975);
DFFARX1 I_49734 (I847992,I2507,I847599,I847585,);
nor I_49735 (I848023,I847625,I847958);
DFFARX1 I_49736 (I848023,I2507,I847599,I847570,);
nor I_49737 (I848054,I847902,I847958);
not I_49738 (I848071,I848054);
nand I_49739 (I847579,I848071,I847927);
not I_49740 (I848126,I2514);
DFFARX1 I_49741 (I771750,I2507,I848126,I848152,);
not I_49742 (I848160,I848152);
nand I_49743 (I848177,I771753,I771750);
and I_49744 (I848194,I848177,I771762);
DFFARX1 I_49745 (I848194,I2507,I848126,I848220,);
DFFARX1 I_49746 (I848220,I2507,I848126,I848115,);
DFFARX1 I_49747 (I771759,I2507,I848126,I848251,);
nand I_49748 (I848259,I848251,I771765);
not I_49749 (I848276,I848259);
DFFARX1 I_49750 (I848276,I2507,I848126,I848302,);
not I_49751 (I848310,I848302);
nor I_49752 (I848118,I848160,I848310);
DFFARX1 I_49753 (I771774,I2507,I848126,I848350,);
nor I_49754 (I848109,I848350,I848220);
nor I_49755 (I848100,I848350,I848276);
nand I_49756 (I848386,I771768,I771756);
and I_49757 (I848403,I848386,I771753);
DFFARX1 I_49758 (I848403,I2507,I848126,I848429,);
not I_49759 (I848437,I848429);
nand I_49760 (I848454,I848437,I848350);
nand I_49761 (I848103,I848437,I848259);
nor I_49762 (I848485,I771771,I771756);
and I_49763 (I848502,I848350,I848485);
nor I_49764 (I848519,I848437,I848502);
DFFARX1 I_49765 (I848519,I2507,I848126,I848112,);
nor I_49766 (I848550,I848152,I848485);
DFFARX1 I_49767 (I848550,I2507,I848126,I848097,);
nor I_49768 (I848581,I848429,I848485);
not I_49769 (I848598,I848581);
nand I_49770 (I848106,I848598,I848454);
not I_49771 (I848653,I2514);
DFFARX1 I_49772 (I357707,I2507,I848653,I848679,);
not I_49773 (I848687,I848679);
nand I_49774 (I848704,I357698,I357698);
and I_49775 (I848721,I848704,I357716);
DFFARX1 I_49776 (I848721,I2507,I848653,I848747,);
DFFARX1 I_49777 (I848747,I2507,I848653,I848642,);
DFFARX1 I_49778 (I357719,I2507,I848653,I848778,);
nand I_49779 (I848786,I848778,I357701);
not I_49780 (I848803,I848786);
DFFARX1 I_49781 (I848803,I2507,I848653,I848829,);
not I_49782 (I848837,I848829);
nor I_49783 (I848645,I848687,I848837);
DFFARX1 I_49784 (I357713,I2507,I848653,I848877,);
nor I_49785 (I848636,I848877,I848747);
nor I_49786 (I848627,I848877,I848803);
nand I_49787 (I848913,I357725,I357704);
and I_49788 (I848930,I848913,I357710);
DFFARX1 I_49789 (I848930,I2507,I848653,I848956,);
not I_49790 (I848964,I848956);
nand I_49791 (I848981,I848964,I848877);
nand I_49792 (I848630,I848964,I848786);
nor I_49793 (I849012,I357722,I357704);
and I_49794 (I849029,I848877,I849012);
nor I_49795 (I849046,I848964,I849029);
DFFARX1 I_49796 (I849046,I2507,I848653,I848639,);
nor I_49797 (I849077,I848679,I849012);
DFFARX1 I_49798 (I849077,I2507,I848653,I848624,);
nor I_49799 (I849108,I848956,I849012);
not I_49800 (I849125,I849108);
nand I_49801 (I848633,I849125,I848981);
not I_49802 (I849180,I2514);
DFFARX1 I_49803 (I1204622,I2507,I849180,I849206,);
not I_49804 (I849214,I849206);
nand I_49805 (I849231,I1204604,I1204604);
and I_49806 (I849248,I849231,I1204610);
DFFARX1 I_49807 (I849248,I2507,I849180,I849274,);
DFFARX1 I_49808 (I849274,I2507,I849180,I849169,);
DFFARX1 I_49809 (I1204607,I2507,I849180,I849305,);
nand I_49810 (I849313,I849305,I1204616);
not I_49811 (I849330,I849313);
DFFARX1 I_49812 (I849330,I2507,I849180,I849356,);
not I_49813 (I849364,I849356);
nor I_49814 (I849172,I849214,I849364);
DFFARX1 I_49815 (I1204628,I2507,I849180,I849404,);
nor I_49816 (I849163,I849404,I849274);
nor I_49817 (I849154,I849404,I849330);
nand I_49818 (I849440,I1204619,I1204613);
and I_49819 (I849457,I849440,I1204607);
DFFARX1 I_49820 (I849457,I2507,I849180,I849483,);
not I_49821 (I849491,I849483);
nand I_49822 (I849508,I849491,I849404);
nand I_49823 (I849157,I849491,I849313);
nor I_49824 (I849539,I1204625,I1204613);
and I_49825 (I849556,I849404,I849539);
nor I_49826 (I849573,I849491,I849556);
DFFARX1 I_49827 (I849573,I2507,I849180,I849166,);
nor I_49828 (I849604,I849206,I849539);
DFFARX1 I_49829 (I849604,I2507,I849180,I849151,);
nor I_49830 (I849635,I849483,I849539);
not I_49831 (I849652,I849635);
nand I_49832 (I849160,I849652,I849508);
not I_49833 (I849707,I2514);
DFFARX1 I_49834 (I475157,I2507,I849707,I849733,);
not I_49835 (I849741,I849733);
nand I_49836 (I849758,I475154,I475163);
and I_49837 (I849775,I849758,I475172);
DFFARX1 I_49838 (I849775,I2507,I849707,I849801,);
DFFARX1 I_49839 (I849801,I2507,I849707,I849696,);
DFFARX1 I_49840 (I475175,I2507,I849707,I849832,);
nand I_49841 (I849840,I849832,I475178);
not I_49842 (I849857,I849840);
DFFARX1 I_49843 (I849857,I2507,I849707,I849883,);
not I_49844 (I849891,I849883);
nor I_49845 (I849699,I849741,I849891);
DFFARX1 I_49846 (I475151,I2507,I849707,I849931,);
nor I_49847 (I849690,I849931,I849801);
nor I_49848 (I849681,I849931,I849857);
nand I_49849 (I849967,I475166,I475169);
and I_49850 (I849984,I849967,I475160);
DFFARX1 I_49851 (I849984,I2507,I849707,I850010,);
not I_49852 (I850018,I850010);
nand I_49853 (I850035,I850018,I849931);
nand I_49854 (I849684,I850018,I849840);
nor I_49855 (I850066,I475151,I475169);
and I_49856 (I850083,I849931,I850066);
nor I_49857 (I850100,I850018,I850083);
DFFARX1 I_49858 (I850100,I2507,I849707,I849693,);
nor I_49859 (I850131,I849733,I850066);
DFFARX1 I_49860 (I850131,I2507,I849707,I849678,);
nor I_49861 (I850162,I850010,I850066);
not I_49862 (I850179,I850162);
nand I_49863 (I849687,I850179,I850035);
not I_49864 (I850234,I2514);
DFFARX1 I_49865 (I446869,I2507,I850234,I850260,);
not I_49866 (I850268,I850260);
nand I_49867 (I850285,I446866,I446875);
and I_49868 (I850302,I850285,I446884);
DFFARX1 I_49869 (I850302,I2507,I850234,I850328,);
DFFARX1 I_49870 (I850328,I2507,I850234,I850223,);
DFFARX1 I_49871 (I446887,I2507,I850234,I850359,);
nand I_49872 (I850367,I850359,I446890);
not I_49873 (I850384,I850367);
DFFARX1 I_49874 (I850384,I2507,I850234,I850410,);
not I_49875 (I850418,I850410);
nor I_49876 (I850226,I850268,I850418);
DFFARX1 I_49877 (I446863,I2507,I850234,I850458,);
nor I_49878 (I850217,I850458,I850328);
nor I_49879 (I850208,I850458,I850384);
nand I_49880 (I850494,I446878,I446881);
and I_49881 (I850511,I850494,I446872);
DFFARX1 I_49882 (I850511,I2507,I850234,I850537,);
not I_49883 (I850545,I850537);
nand I_49884 (I850562,I850545,I850458);
nand I_49885 (I850211,I850545,I850367);
nor I_49886 (I850593,I446863,I446881);
and I_49887 (I850610,I850458,I850593);
nor I_49888 (I850627,I850545,I850610);
DFFARX1 I_49889 (I850627,I2507,I850234,I850220,);
nor I_49890 (I850658,I850260,I850593);
DFFARX1 I_49891 (I850658,I2507,I850234,I850205,);
nor I_49892 (I850689,I850537,I850593);
not I_49893 (I850706,I850689);
nand I_49894 (I850214,I850706,I850562);
not I_49895 (I850761,I2514);
DFFARX1 I_49896 (I44856,I2507,I850761,I850787,);
not I_49897 (I850795,I850787);
nand I_49898 (I850812,I44868,I44871);
and I_49899 (I850829,I850812,I44847);
DFFARX1 I_49900 (I850829,I2507,I850761,I850855,);
DFFARX1 I_49901 (I850855,I2507,I850761,I850750,);
DFFARX1 I_49902 (I44865,I2507,I850761,I850886,);
nand I_49903 (I850894,I850886,I44853);
not I_49904 (I850911,I850894);
DFFARX1 I_49905 (I850911,I2507,I850761,I850937,);
not I_49906 (I850945,I850937);
nor I_49907 (I850753,I850795,I850945);
DFFARX1 I_49908 (I44850,I2507,I850761,I850985,);
nor I_49909 (I850744,I850985,I850855);
nor I_49910 (I850735,I850985,I850911);
nand I_49911 (I851021,I44859,I44850);
and I_49912 (I851038,I851021,I44847);
DFFARX1 I_49913 (I851038,I2507,I850761,I851064,);
not I_49914 (I851072,I851064);
nand I_49915 (I851089,I851072,I850985);
nand I_49916 (I850738,I851072,I850894);
nor I_49917 (I851120,I44862,I44850);
and I_49918 (I851137,I850985,I851120);
nor I_49919 (I851154,I851072,I851137);
DFFARX1 I_49920 (I851154,I2507,I850761,I850747,);
nor I_49921 (I851185,I850787,I851120);
DFFARX1 I_49922 (I851185,I2507,I850761,I850732,);
nor I_49923 (I851216,I851064,I851120);
not I_49924 (I851233,I851216);
nand I_49925 (I850741,I851233,I851089);
not I_49926 (I851288,I2514);
DFFARX1 I_49927 (I1265176,I2507,I851288,I851314,);
not I_49928 (I851322,I851314);
nand I_49929 (I851339,I1265158,I1265161);
and I_49930 (I851356,I851339,I1265173);
DFFARX1 I_49931 (I851356,I2507,I851288,I851382,);
DFFARX1 I_49932 (I851382,I2507,I851288,I851277,);
DFFARX1 I_49933 (I1265182,I2507,I851288,I851413,);
nand I_49934 (I851421,I851413,I1265167);
not I_49935 (I851438,I851421);
DFFARX1 I_49936 (I851438,I2507,I851288,I851464,);
not I_49937 (I851472,I851464);
nor I_49938 (I851280,I851322,I851472);
DFFARX1 I_49939 (I1265179,I2507,I851288,I851512,);
nor I_49940 (I851271,I851512,I851382);
nor I_49941 (I851262,I851512,I851438);
nand I_49942 (I851548,I1265170,I1265164);
and I_49943 (I851565,I851548,I1265158);
DFFARX1 I_49944 (I851565,I2507,I851288,I851591,);
not I_49945 (I851599,I851591);
nand I_49946 (I851616,I851599,I851512);
nand I_49947 (I851265,I851599,I851421);
nor I_49948 (I851647,I1265161,I1265164);
and I_49949 (I851664,I851512,I851647);
nor I_49950 (I851681,I851599,I851664);
DFFARX1 I_49951 (I851681,I2507,I851288,I851274,);
nor I_49952 (I851712,I851314,I851647);
DFFARX1 I_49953 (I851712,I2507,I851288,I851259,);
nor I_49954 (I851743,I851591,I851647);
not I_49955 (I851760,I851743);
nand I_49956 (I851268,I851760,I851616);
not I_49957 (I851815,I2514);
DFFARX1 I_49958 (I702968,I2507,I851815,I851841,);
not I_49959 (I851849,I851841);
nand I_49960 (I851866,I702971,I702968);
and I_49961 (I851883,I851866,I702980);
DFFARX1 I_49962 (I851883,I2507,I851815,I851909,);
DFFARX1 I_49963 (I851909,I2507,I851815,I851804,);
DFFARX1 I_49964 (I702977,I2507,I851815,I851940,);
nand I_49965 (I851948,I851940,I702983);
not I_49966 (I851965,I851948);
DFFARX1 I_49967 (I851965,I2507,I851815,I851991,);
not I_49968 (I851999,I851991);
nor I_49969 (I851807,I851849,I851999);
DFFARX1 I_49970 (I702992,I2507,I851815,I852039,);
nor I_49971 (I851798,I852039,I851909);
nor I_49972 (I851789,I852039,I851965);
nand I_49973 (I852075,I702986,I702974);
and I_49974 (I852092,I852075,I702971);
DFFARX1 I_49975 (I852092,I2507,I851815,I852118,);
not I_49976 (I852126,I852118);
nand I_49977 (I852143,I852126,I852039);
nand I_49978 (I851792,I852126,I851948);
nor I_49979 (I852174,I702989,I702974);
and I_49980 (I852191,I852039,I852174);
nor I_49981 (I852208,I852126,I852191);
DFFARX1 I_49982 (I852208,I2507,I851815,I851801,);
nor I_49983 (I852239,I851841,I852174);
DFFARX1 I_49984 (I852239,I2507,I851815,I851786,);
nor I_49985 (I852270,I852118,I852174);
not I_49986 (I852287,I852270);
nand I_49987 (I851795,I852287,I852143);
not I_49988 (I852342,I2514);
DFFARX1 I_49989 (I276022,I2507,I852342,I852368,);
not I_49990 (I852376,I852368);
nand I_49991 (I852393,I276013,I276013);
and I_49992 (I852410,I852393,I276031);
DFFARX1 I_49993 (I852410,I2507,I852342,I852436,);
DFFARX1 I_49994 (I852436,I2507,I852342,I852331,);
DFFARX1 I_49995 (I276034,I2507,I852342,I852467,);
nand I_49996 (I852475,I852467,I276016);
not I_49997 (I852492,I852475);
DFFARX1 I_49998 (I852492,I2507,I852342,I852518,);
not I_49999 (I852526,I852518);
nor I_50000 (I852334,I852376,I852526);
DFFARX1 I_50001 (I276028,I2507,I852342,I852566,);
nor I_50002 (I852325,I852566,I852436);
nor I_50003 (I852316,I852566,I852492);
nand I_50004 (I852602,I276040,I276019);
and I_50005 (I852619,I852602,I276025);
DFFARX1 I_50006 (I852619,I2507,I852342,I852645,);
not I_50007 (I852653,I852645);
nand I_50008 (I852670,I852653,I852566);
nand I_50009 (I852319,I852653,I852475);
nor I_50010 (I852701,I276037,I276019);
and I_50011 (I852718,I852566,I852701);
nor I_50012 (I852735,I852653,I852718);
DFFARX1 I_50013 (I852735,I2507,I852342,I852328,);
nor I_50014 (I852766,I852368,I852701);
DFFARX1 I_50015 (I852766,I2507,I852342,I852313,);
nor I_50016 (I852797,I852645,I852701);
not I_50017 (I852814,I852797);
nand I_50018 (I852322,I852814,I852670);
not I_50019 (I852869,I2514);
DFFARX1 I_50020 (I1075150,I2507,I852869,I852895,);
not I_50021 (I852903,I852895);
nand I_50022 (I852920,I1075132,I1075132);
and I_50023 (I852937,I852920,I1075138);
DFFARX1 I_50024 (I852937,I2507,I852869,I852963,);
DFFARX1 I_50025 (I852963,I2507,I852869,I852858,);
DFFARX1 I_50026 (I1075135,I2507,I852869,I852994,);
nand I_50027 (I853002,I852994,I1075144);
not I_50028 (I853019,I853002);
DFFARX1 I_50029 (I853019,I2507,I852869,I853045,);
not I_50030 (I853053,I853045);
nor I_50031 (I852861,I852903,I853053);
DFFARX1 I_50032 (I1075156,I2507,I852869,I853093,);
nor I_50033 (I852852,I853093,I852963);
nor I_50034 (I852843,I853093,I853019);
nand I_50035 (I853129,I1075147,I1075141);
and I_50036 (I853146,I853129,I1075135);
DFFARX1 I_50037 (I853146,I2507,I852869,I853172,);
not I_50038 (I853180,I853172);
nand I_50039 (I853197,I853180,I853093);
nand I_50040 (I852846,I853180,I853002);
nor I_50041 (I853228,I1075153,I1075141);
and I_50042 (I853245,I853093,I853228);
nor I_50043 (I853262,I853180,I853245);
DFFARX1 I_50044 (I853262,I2507,I852869,I852855,);
nor I_50045 (I853293,I852895,I853228);
DFFARX1 I_50046 (I853293,I2507,I852869,I852840,);
nor I_50047 (I853324,I853172,I853228);
not I_50048 (I853341,I853324);
nand I_50049 (I852849,I853341,I853197);
not I_50050 (I853396,I2514);
DFFARX1 I_50051 (I774062,I2507,I853396,I853422,);
not I_50052 (I853430,I853422);
nand I_50053 (I853447,I774065,I774062);
and I_50054 (I853464,I853447,I774074);
DFFARX1 I_50055 (I853464,I2507,I853396,I853490,);
DFFARX1 I_50056 (I853490,I2507,I853396,I853385,);
DFFARX1 I_50057 (I774071,I2507,I853396,I853521,);
nand I_50058 (I853529,I853521,I774077);
not I_50059 (I853546,I853529);
DFFARX1 I_50060 (I853546,I2507,I853396,I853572,);
not I_50061 (I853580,I853572);
nor I_50062 (I853388,I853430,I853580);
DFFARX1 I_50063 (I774086,I2507,I853396,I853620,);
nor I_50064 (I853379,I853620,I853490);
nor I_50065 (I853370,I853620,I853546);
nand I_50066 (I853656,I774080,I774068);
and I_50067 (I853673,I853656,I774065);
DFFARX1 I_50068 (I853673,I2507,I853396,I853699,);
not I_50069 (I853707,I853699);
nand I_50070 (I853724,I853707,I853620);
nand I_50071 (I853373,I853707,I853529);
nor I_50072 (I853755,I774083,I774068);
and I_50073 (I853772,I853620,I853755);
nor I_50074 (I853789,I853707,I853772);
DFFARX1 I_50075 (I853789,I2507,I853396,I853382,);
nor I_50076 (I853820,I853422,I853755);
DFFARX1 I_50077 (I853820,I2507,I853396,I853367,);
nor I_50078 (I853851,I853699,I853755);
not I_50079 (I853868,I853851);
nand I_50080 (I853376,I853868,I853724);
not I_50081 (I853923,I2514);
DFFARX1 I_50082 (I708748,I2507,I853923,I853949,);
not I_50083 (I853957,I853949);
nand I_50084 (I853974,I708751,I708748);
and I_50085 (I853991,I853974,I708760);
DFFARX1 I_50086 (I853991,I2507,I853923,I854017,);
DFFARX1 I_50087 (I854017,I2507,I853923,I853912,);
DFFARX1 I_50088 (I708757,I2507,I853923,I854048,);
nand I_50089 (I854056,I854048,I708763);
not I_50090 (I854073,I854056);
DFFARX1 I_50091 (I854073,I2507,I853923,I854099,);
not I_50092 (I854107,I854099);
nor I_50093 (I853915,I853957,I854107);
DFFARX1 I_50094 (I708772,I2507,I853923,I854147,);
nor I_50095 (I853906,I854147,I854017);
nor I_50096 (I853897,I854147,I854073);
nand I_50097 (I854183,I708766,I708754);
and I_50098 (I854200,I854183,I708751);
DFFARX1 I_50099 (I854200,I2507,I853923,I854226,);
not I_50100 (I854234,I854226);
nand I_50101 (I854251,I854234,I854147);
nand I_50102 (I853900,I854234,I854056);
nor I_50103 (I854282,I708769,I708754);
and I_50104 (I854299,I854147,I854282);
nor I_50105 (I854316,I854234,I854299);
DFFARX1 I_50106 (I854316,I2507,I853923,I853909,);
nor I_50107 (I854347,I853949,I854282);
DFFARX1 I_50108 (I854347,I2507,I853923,I853894,);
nor I_50109 (I854378,I854226,I854282);
not I_50110 (I854395,I854378);
nand I_50111 (I853903,I854395,I854251);
not I_50112 (I854450,I2514);
DFFARX1 I_50113 (I1380892,I2507,I854450,I854476,);
not I_50114 (I854484,I854476);
nand I_50115 (I854501,I1380889,I1380898);
and I_50116 (I854518,I854501,I1380877);
DFFARX1 I_50117 (I854518,I2507,I854450,I854544,);
DFFARX1 I_50118 (I854544,I2507,I854450,I854439,);
DFFARX1 I_50119 (I1380880,I2507,I854450,I854575,);
nand I_50120 (I854583,I854575,I1380895);
not I_50121 (I854600,I854583);
DFFARX1 I_50122 (I854600,I2507,I854450,I854626,);
not I_50123 (I854634,I854626);
nor I_50124 (I854442,I854484,I854634);
DFFARX1 I_50125 (I1380901,I2507,I854450,I854674,);
nor I_50126 (I854433,I854674,I854544);
nor I_50127 (I854424,I854674,I854600);
nand I_50128 (I854710,I1380883,I1380904);
and I_50129 (I854727,I854710,I1380886);
DFFARX1 I_50130 (I854727,I2507,I854450,I854753,);
not I_50131 (I854761,I854753);
nand I_50132 (I854778,I854761,I854674);
nand I_50133 (I854427,I854761,I854583);
nor I_50134 (I854809,I1380877,I1380904);
and I_50135 (I854826,I854674,I854809);
nor I_50136 (I854843,I854761,I854826);
DFFARX1 I_50137 (I854843,I2507,I854450,I854436,);
nor I_50138 (I854874,I854476,I854809);
DFFARX1 I_50139 (I854874,I2507,I854450,I854421,);
nor I_50140 (I854905,I854753,I854809);
not I_50141 (I854922,I854905);
nand I_50142 (I854430,I854922,I854778);
not I_50143 (I854977,I2514);
DFFARX1 I_50144 (I456661,I2507,I854977,I855003,);
not I_50145 (I855011,I855003);
nand I_50146 (I855028,I456658,I456667);
and I_50147 (I855045,I855028,I456676);
DFFARX1 I_50148 (I855045,I2507,I854977,I855071,);
DFFARX1 I_50149 (I855071,I2507,I854977,I854966,);
DFFARX1 I_50150 (I456679,I2507,I854977,I855102,);
nand I_50151 (I855110,I855102,I456682);
not I_50152 (I855127,I855110);
DFFARX1 I_50153 (I855127,I2507,I854977,I855153,);
not I_50154 (I855161,I855153);
nor I_50155 (I854969,I855011,I855161);
DFFARX1 I_50156 (I456655,I2507,I854977,I855201,);
nor I_50157 (I854960,I855201,I855071);
nor I_50158 (I854951,I855201,I855127);
nand I_50159 (I855237,I456670,I456673);
and I_50160 (I855254,I855237,I456664);
DFFARX1 I_50161 (I855254,I2507,I854977,I855280,);
not I_50162 (I855288,I855280);
nand I_50163 (I855305,I855288,I855201);
nand I_50164 (I854954,I855288,I855110);
nor I_50165 (I855336,I456655,I456673);
and I_50166 (I855353,I855201,I855336);
nor I_50167 (I855370,I855288,I855353);
DFFARX1 I_50168 (I855370,I2507,I854977,I854963,);
nor I_50169 (I855401,I855003,I855336);
DFFARX1 I_50170 (I855401,I2507,I854977,I854948,);
nor I_50171 (I855432,I855280,I855336);
not I_50172 (I855449,I855432);
nand I_50173 (I854957,I855449,I855305);
not I_50174 (I855504,I2514);
DFFARX1 I_50175 (I484405,I2507,I855504,I855530,);
not I_50176 (I855538,I855530);
nand I_50177 (I855555,I484402,I484411);
and I_50178 (I855572,I855555,I484420);
DFFARX1 I_50179 (I855572,I2507,I855504,I855598,);
DFFARX1 I_50180 (I855598,I2507,I855504,I855493,);
DFFARX1 I_50181 (I484423,I2507,I855504,I855629,);
nand I_50182 (I855637,I855629,I484426);
not I_50183 (I855654,I855637);
DFFARX1 I_50184 (I855654,I2507,I855504,I855680,);
not I_50185 (I855688,I855680);
nor I_50186 (I855496,I855538,I855688);
DFFARX1 I_50187 (I484399,I2507,I855504,I855728,);
nor I_50188 (I855487,I855728,I855598);
nor I_50189 (I855478,I855728,I855654);
nand I_50190 (I855764,I484414,I484417);
and I_50191 (I855781,I855764,I484408);
DFFARX1 I_50192 (I855781,I2507,I855504,I855807,);
not I_50193 (I855815,I855807);
nand I_50194 (I855832,I855815,I855728);
nand I_50195 (I855481,I855815,I855637);
nor I_50196 (I855863,I484399,I484417);
and I_50197 (I855880,I855728,I855863);
nor I_50198 (I855897,I855815,I855880);
DFFARX1 I_50199 (I855897,I2507,I855504,I855490,);
nor I_50200 (I855928,I855530,I855863);
DFFARX1 I_50201 (I855928,I2507,I855504,I855475,);
nor I_50202 (I855959,I855807,I855863);
not I_50203 (I855976,I855959);
nand I_50204 (I855484,I855976,I855832);
not I_50205 (I856031,I2514);
DFFARX1 I_50206 (I1183236,I2507,I856031,I856057,);
not I_50207 (I856065,I856057);
nand I_50208 (I856082,I1183218,I1183218);
and I_50209 (I856099,I856082,I1183224);
DFFARX1 I_50210 (I856099,I2507,I856031,I856125,);
DFFARX1 I_50211 (I856125,I2507,I856031,I856020,);
DFFARX1 I_50212 (I1183221,I2507,I856031,I856156,);
nand I_50213 (I856164,I856156,I1183230);
not I_50214 (I856181,I856164);
DFFARX1 I_50215 (I856181,I2507,I856031,I856207,);
not I_50216 (I856215,I856207);
nor I_50217 (I856023,I856065,I856215);
DFFARX1 I_50218 (I1183242,I2507,I856031,I856255,);
nor I_50219 (I856014,I856255,I856125);
nor I_50220 (I856005,I856255,I856181);
nand I_50221 (I856291,I1183233,I1183227);
and I_50222 (I856308,I856291,I1183221);
DFFARX1 I_50223 (I856308,I2507,I856031,I856334,);
not I_50224 (I856342,I856334);
nand I_50225 (I856359,I856342,I856255);
nand I_50226 (I856008,I856342,I856164);
nor I_50227 (I856390,I1183239,I1183227);
and I_50228 (I856407,I856255,I856390);
nor I_50229 (I856424,I856342,I856407);
DFFARX1 I_50230 (I856424,I2507,I856031,I856017,);
nor I_50231 (I856455,I856057,I856390);
DFFARX1 I_50232 (I856455,I2507,I856031,I856002,);
nor I_50233 (I856486,I856334,I856390);
not I_50234 (I856503,I856486);
nand I_50235 (I856011,I856503,I856359);
not I_50236 (I856558,I2514);
DFFARX1 I_50237 (I766548,I2507,I856558,I856584,);
not I_50238 (I856592,I856584);
nand I_50239 (I856609,I766551,I766548);
and I_50240 (I856626,I856609,I766560);
DFFARX1 I_50241 (I856626,I2507,I856558,I856652,);
DFFARX1 I_50242 (I856652,I2507,I856558,I856547,);
DFFARX1 I_50243 (I766557,I2507,I856558,I856683,);
nand I_50244 (I856691,I856683,I766563);
not I_50245 (I856708,I856691);
DFFARX1 I_50246 (I856708,I2507,I856558,I856734,);
not I_50247 (I856742,I856734);
nor I_50248 (I856550,I856592,I856742);
DFFARX1 I_50249 (I766572,I2507,I856558,I856782,);
nor I_50250 (I856541,I856782,I856652);
nor I_50251 (I856532,I856782,I856708);
nand I_50252 (I856818,I766566,I766554);
and I_50253 (I856835,I856818,I766551);
DFFARX1 I_50254 (I856835,I2507,I856558,I856861,);
not I_50255 (I856869,I856861);
nand I_50256 (I856886,I856869,I856782);
nand I_50257 (I856535,I856869,I856691);
nor I_50258 (I856917,I766569,I766554);
and I_50259 (I856934,I856782,I856917);
nor I_50260 (I856951,I856869,I856934);
DFFARX1 I_50261 (I856951,I2507,I856558,I856544,);
nor I_50262 (I856982,I856584,I856917);
DFFARX1 I_50263 (I856982,I2507,I856558,I856529,);
nor I_50264 (I857013,I856861,I856917);
not I_50265 (I857030,I857013);
nand I_50266 (I856538,I857030,I856886);
not I_50267 (I857085,I2514);
DFFARX1 I_50268 (I978014,I2507,I857085,I857111,);
not I_50269 (I857119,I857111);
nand I_50270 (I857136,I978029,I978011);
and I_50271 (I857153,I857136,I978011);
DFFARX1 I_50272 (I857153,I2507,I857085,I857179,);
DFFARX1 I_50273 (I857179,I2507,I857085,I857074,);
DFFARX1 I_50274 (I978020,I2507,I857085,I857210,);
nand I_50275 (I857218,I857210,I978038);
not I_50276 (I857235,I857218);
DFFARX1 I_50277 (I857235,I2507,I857085,I857261,);
not I_50278 (I857269,I857261);
nor I_50279 (I857077,I857119,I857269);
DFFARX1 I_50280 (I978035,I2507,I857085,I857309,);
nor I_50281 (I857068,I857309,I857179);
nor I_50282 (I857059,I857309,I857235);
nand I_50283 (I857345,I978032,I978023);
and I_50284 (I857362,I857345,I978017);
DFFARX1 I_50285 (I857362,I2507,I857085,I857388,);
not I_50286 (I857396,I857388);
nand I_50287 (I857413,I857396,I857309);
nand I_50288 (I857062,I857396,I857218);
nor I_50289 (I857444,I978026,I978023);
and I_50290 (I857461,I857309,I857444);
nor I_50291 (I857478,I857396,I857461);
DFFARX1 I_50292 (I857478,I2507,I857085,I857071,);
nor I_50293 (I857509,I857111,I857444);
DFFARX1 I_50294 (I857509,I2507,I857085,I857056,);
nor I_50295 (I857540,I857388,I857444);
not I_50296 (I857557,I857540);
nand I_50297 (I857065,I857557,I857413);
not I_50298 (I857612,I2514);
DFFARX1 I_50299 (I997394,I2507,I857612,I857638,);
not I_50300 (I857646,I857638);
nand I_50301 (I857663,I997409,I997391);
and I_50302 (I857680,I857663,I997391);
DFFARX1 I_50303 (I857680,I2507,I857612,I857706,);
DFFARX1 I_50304 (I857706,I2507,I857612,I857601,);
DFFARX1 I_50305 (I997400,I2507,I857612,I857737,);
nand I_50306 (I857745,I857737,I997418);
not I_50307 (I857762,I857745);
DFFARX1 I_50308 (I857762,I2507,I857612,I857788,);
not I_50309 (I857796,I857788);
nor I_50310 (I857604,I857646,I857796);
DFFARX1 I_50311 (I997415,I2507,I857612,I857836,);
nor I_50312 (I857595,I857836,I857706);
nor I_50313 (I857586,I857836,I857762);
nand I_50314 (I857872,I997412,I997403);
and I_50315 (I857889,I857872,I997397);
DFFARX1 I_50316 (I857889,I2507,I857612,I857915,);
not I_50317 (I857923,I857915);
nand I_50318 (I857940,I857923,I857836);
nand I_50319 (I857589,I857923,I857745);
nor I_50320 (I857971,I997406,I997403);
and I_50321 (I857988,I857836,I857971);
nor I_50322 (I858005,I857923,I857988);
DFFARX1 I_50323 (I858005,I2507,I857612,I857598,);
nor I_50324 (I858036,I857638,I857971);
DFFARX1 I_50325 (I858036,I2507,I857612,I857583,);
nor I_50326 (I858067,I857915,I857971);
not I_50327 (I858084,I858067);
nand I_50328 (I857592,I858084,I857940);
not I_50329 (I858139,I2514);
DFFARX1 I_50330 (I1015199,I2507,I858139,I858165,);
not I_50331 (I858173,I858165);
nand I_50332 (I858190,I1015208,I1015196);
and I_50333 (I858207,I858190,I1015193);
DFFARX1 I_50334 (I858207,I2507,I858139,I858233,);
DFFARX1 I_50335 (I858233,I2507,I858139,I858128,);
DFFARX1 I_50336 (I1015193,I2507,I858139,I858264,);
nand I_50337 (I858272,I858264,I1015190);
not I_50338 (I858289,I858272);
DFFARX1 I_50339 (I858289,I2507,I858139,I858315,);
not I_50340 (I858323,I858315);
nor I_50341 (I858131,I858173,I858323);
DFFARX1 I_50342 (I1015196,I2507,I858139,I858363,);
nor I_50343 (I858122,I858363,I858233);
nor I_50344 (I858113,I858363,I858289);
nand I_50345 (I858399,I1015211,I1015202);
and I_50346 (I858416,I858399,I1015205);
DFFARX1 I_50347 (I858416,I2507,I858139,I858442,);
not I_50348 (I858450,I858442);
nand I_50349 (I858467,I858450,I858363);
nand I_50350 (I858116,I858450,I858272);
nor I_50351 (I858498,I1015190,I1015202);
and I_50352 (I858515,I858363,I858498);
nor I_50353 (I858532,I858450,I858515);
DFFARX1 I_50354 (I858532,I2507,I858139,I858125,);
nor I_50355 (I858563,I858165,I858498);
DFFARX1 I_50356 (I858563,I2507,I858139,I858110,);
nor I_50357 (I858594,I858442,I858498);
not I_50358 (I858611,I858594);
nand I_50359 (I858119,I858611,I858467);
not I_50360 (I858666,I2514);
DFFARX1 I_50361 (I741116,I2507,I858666,I858692,);
not I_50362 (I858700,I858692);
nand I_50363 (I858717,I741119,I741116);
and I_50364 (I858734,I858717,I741128);
DFFARX1 I_50365 (I858734,I2507,I858666,I858760,);
DFFARX1 I_50366 (I858760,I2507,I858666,I858655,);
DFFARX1 I_50367 (I741125,I2507,I858666,I858791,);
nand I_50368 (I858799,I858791,I741131);
not I_50369 (I858816,I858799);
DFFARX1 I_50370 (I858816,I2507,I858666,I858842,);
not I_50371 (I858850,I858842);
nor I_50372 (I858658,I858700,I858850);
DFFARX1 I_50373 (I741140,I2507,I858666,I858890,);
nor I_50374 (I858649,I858890,I858760);
nor I_50375 (I858640,I858890,I858816);
nand I_50376 (I858926,I741134,I741122);
and I_50377 (I858943,I858926,I741119);
DFFARX1 I_50378 (I858943,I2507,I858666,I858969,);
not I_50379 (I858977,I858969);
nand I_50380 (I858994,I858977,I858890);
nand I_50381 (I858643,I858977,I858799);
nor I_50382 (I859025,I741137,I741122);
and I_50383 (I859042,I858890,I859025);
nor I_50384 (I859059,I858977,I859042);
DFFARX1 I_50385 (I859059,I2507,I858666,I858652,);
nor I_50386 (I859090,I858692,I859025);
DFFARX1 I_50387 (I859090,I2507,I858666,I858637,);
nor I_50388 (I859121,I858969,I859025);
not I_50389 (I859138,I859121);
nand I_50390 (I858646,I859138,I858994);
not I_50391 (I859193,I2514);
DFFARX1 I_50392 (I890804,I2507,I859193,I859219,);
not I_50393 (I859227,I859219);
nand I_50394 (I859244,I890819,I890801);
and I_50395 (I859261,I859244,I890801);
DFFARX1 I_50396 (I859261,I2507,I859193,I859287,);
DFFARX1 I_50397 (I859287,I2507,I859193,I859182,);
DFFARX1 I_50398 (I890810,I2507,I859193,I859318,);
nand I_50399 (I859326,I859318,I890828);
not I_50400 (I859343,I859326);
DFFARX1 I_50401 (I859343,I2507,I859193,I859369,);
not I_50402 (I859377,I859369);
nor I_50403 (I859185,I859227,I859377);
DFFARX1 I_50404 (I890825,I2507,I859193,I859417,);
nor I_50405 (I859176,I859417,I859287);
nor I_50406 (I859167,I859417,I859343);
nand I_50407 (I859453,I890822,I890813);
and I_50408 (I859470,I859453,I890807);
DFFARX1 I_50409 (I859470,I2507,I859193,I859496,);
not I_50410 (I859504,I859496);
nand I_50411 (I859521,I859504,I859417);
nand I_50412 (I859170,I859504,I859326);
nor I_50413 (I859552,I890816,I890813);
and I_50414 (I859569,I859417,I859552);
nor I_50415 (I859586,I859504,I859569);
DFFARX1 I_50416 (I859586,I2507,I859193,I859179,);
nor I_50417 (I859617,I859219,I859552);
DFFARX1 I_50418 (I859617,I2507,I859193,I859164,);
nor I_50419 (I859648,I859496,I859552);
not I_50420 (I859665,I859648);
nand I_50421 (I859173,I859665,I859521);
not I_50422 (I859720,I2514);
DFFARX1 I_50423 (I260212,I2507,I859720,I859746,);
not I_50424 (I859754,I859746);
nand I_50425 (I859771,I260203,I260203);
and I_50426 (I859788,I859771,I260221);
DFFARX1 I_50427 (I859788,I2507,I859720,I859814,);
DFFARX1 I_50428 (I859814,I2507,I859720,I859709,);
DFFARX1 I_50429 (I260224,I2507,I859720,I859845,);
nand I_50430 (I859853,I859845,I260206);
not I_50431 (I859870,I859853);
DFFARX1 I_50432 (I859870,I2507,I859720,I859896,);
not I_50433 (I859904,I859896);
nor I_50434 (I859712,I859754,I859904);
DFFARX1 I_50435 (I260218,I2507,I859720,I859944,);
nor I_50436 (I859703,I859944,I859814);
nor I_50437 (I859694,I859944,I859870);
nand I_50438 (I859980,I260230,I260209);
and I_50439 (I859997,I859980,I260215);
DFFARX1 I_50440 (I859997,I2507,I859720,I860023,);
not I_50441 (I860031,I860023);
nand I_50442 (I860048,I860031,I859944);
nand I_50443 (I859697,I860031,I859853);
nor I_50444 (I860079,I260227,I260209);
and I_50445 (I860096,I859944,I860079);
nor I_50446 (I860113,I860031,I860096);
DFFARX1 I_50447 (I860113,I2507,I859720,I859706,);
nor I_50448 (I860144,I859746,I860079);
DFFARX1 I_50449 (I860144,I2507,I859720,I859691,);
nor I_50450 (I860175,I860023,I860079);
not I_50451 (I860192,I860175);
nand I_50452 (I859700,I860192,I860048);
not I_50453 (I860247,I2514);
DFFARX1 I_50454 (I231156,I2507,I860247,I860273,);
not I_50455 (I860281,I860273);
nand I_50456 (I860298,I231153,I231171);
and I_50457 (I860315,I860298,I231162);
DFFARX1 I_50458 (I860315,I2507,I860247,I860341,);
DFFARX1 I_50459 (I860341,I2507,I860247,I860236,);
DFFARX1 I_50460 (I231168,I2507,I860247,I860372,);
nand I_50461 (I860380,I860372,I231165);
not I_50462 (I860397,I860380);
DFFARX1 I_50463 (I860397,I2507,I860247,I860423,);
not I_50464 (I860431,I860423);
nor I_50465 (I860239,I860281,I860431);
DFFARX1 I_50466 (I231159,I2507,I860247,I860471,);
nor I_50467 (I860230,I860471,I860341);
nor I_50468 (I860221,I860471,I860397);
nand I_50469 (I860507,I231150,I231174);
and I_50470 (I860524,I860507,I231153);
DFFARX1 I_50471 (I860524,I2507,I860247,I860550,);
not I_50472 (I860558,I860550);
nand I_50473 (I860575,I860558,I860471);
nand I_50474 (I860224,I860558,I860380);
nor I_50475 (I860606,I231150,I231174);
and I_50476 (I860623,I860471,I860606);
nor I_50477 (I860640,I860558,I860623);
DFFARX1 I_50478 (I860640,I2507,I860247,I860233,);
nor I_50479 (I860671,I860273,I860606);
DFFARX1 I_50480 (I860671,I2507,I860247,I860218,);
nor I_50481 (I860702,I860550,I860606);
not I_50482 (I860719,I860702);
nand I_50483 (I860227,I860719,I860575);
not I_50484 (I860774,I2514);
DFFARX1 I_50485 (I923104,I2507,I860774,I860800,);
not I_50486 (I860808,I860800);
nand I_50487 (I860825,I923119,I923101);
and I_50488 (I860842,I860825,I923101);
DFFARX1 I_50489 (I860842,I2507,I860774,I860868,);
DFFARX1 I_50490 (I860868,I2507,I860774,I860763,);
DFFARX1 I_50491 (I923110,I2507,I860774,I860899,);
nand I_50492 (I860907,I860899,I923128);
not I_50493 (I860924,I860907);
DFFARX1 I_50494 (I860924,I2507,I860774,I860950,);
not I_50495 (I860958,I860950);
nor I_50496 (I860766,I860808,I860958);
DFFARX1 I_50497 (I923125,I2507,I860774,I860998,);
nor I_50498 (I860757,I860998,I860868);
nor I_50499 (I860748,I860998,I860924);
nand I_50500 (I861034,I923122,I923113);
and I_50501 (I861051,I861034,I923107);
DFFARX1 I_50502 (I861051,I2507,I860774,I861077,);
not I_50503 (I861085,I861077);
nand I_50504 (I861102,I861085,I860998);
nand I_50505 (I860751,I861085,I860907);
nor I_50506 (I861133,I923116,I923113);
and I_50507 (I861150,I860998,I861133);
nor I_50508 (I861167,I861085,I861150);
DFFARX1 I_50509 (I861167,I2507,I860774,I860760,);
nor I_50510 (I861198,I860800,I861133);
DFFARX1 I_50511 (I861198,I2507,I860774,I860745,);
nor I_50512 (I861229,I861077,I861133);
not I_50513 (I861246,I861229);
nand I_50514 (I860754,I861246,I861102);
not I_50515 (I861301,I2514);
DFFARX1 I_50516 (I432725,I2507,I861301,I861327,);
not I_50517 (I861335,I861327);
nand I_50518 (I861352,I432722,I432731);
and I_50519 (I861369,I861352,I432740);
DFFARX1 I_50520 (I861369,I2507,I861301,I861395,);
DFFARX1 I_50521 (I861395,I2507,I861301,I861290,);
DFFARX1 I_50522 (I432743,I2507,I861301,I861426,);
nand I_50523 (I861434,I861426,I432746);
not I_50524 (I861451,I861434);
DFFARX1 I_50525 (I861451,I2507,I861301,I861477,);
not I_50526 (I861485,I861477);
nor I_50527 (I861293,I861335,I861485);
DFFARX1 I_50528 (I432719,I2507,I861301,I861525,);
nor I_50529 (I861284,I861525,I861395);
nor I_50530 (I861275,I861525,I861451);
nand I_50531 (I861561,I432734,I432737);
and I_50532 (I861578,I861561,I432728);
DFFARX1 I_50533 (I861578,I2507,I861301,I861604,);
not I_50534 (I861612,I861604);
nand I_50535 (I861629,I861612,I861525);
nand I_50536 (I861278,I861612,I861434);
nor I_50537 (I861660,I432719,I432737);
and I_50538 (I861677,I861525,I861660);
nor I_50539 (I861694,I861612,I861677);
DFFARX1 I_50540 (I861694,I2507,I861301,I861287,);
nor I_50541 (I861725,I861327,I861660);
DFFARX1 I_50542 (I861725,I2507,I861301,I861272,);
nor I_50543 (I861756,I861604,I861660);
not I_50544 (I861773,I861756);
nand I_50545 (I861281,I861773,I861629);
not I_50546 (I861828,I2514);
DFFARX1 I_50547 (I1142776,I2507,I861828,I861854,);
not I_50548 (I861862,I861854);
nand I_50549 (I861879,I1142758,I1142758);
and I_50550 (I861896,I861879,I1142764);
DFFARX1 I_50551 (I861896,I2507,I861828,I861922,);
DFFARX1 I_50552 (I861922,I2507,I861828,I861817,);
DFFARX1 I_50553 (I1142761,I2507,I861828,I861953,);
nand I_50554 (I861961,I861953,I1142770);
not I_50555 (I861978,I861961);
DFFARX1 I_50556 (I861978,I2507,I861828,I862004,);
not I_50557 (I862012,I862004);
nor I_50558 (I861820,I861862,I862012);
DFFARX1 I_50559 (I1142782,I2507,I861828,I862052,);
nor I_50560 (I861811,I862052,I861922);
nor I_50561 (I861802,I862052,I861978);
nand I_50562 (I862088,I1142773,I1142767);
and I_50563 (I862105,I862088,I1142761);
DFFARX1 I_50564 (I862105,I2507,I861828,I862131,);
not I_50565 (I862139,I862131);
nand I_50566 (I862156,I862139,I862052);
nand I_50567 (I861805,I862139,I861961);
nor I_50568 (I862187,I1142779,I1142767);
and I_50569 (I862204,I862052,I862187);
nor I_50570 (I862221,I862139,I862204);
DFFARX1 I_50571 (I862221,I2507,I861828,I861814,);
nor I_50572 (I862252,I861854,I862187);
DFFARX1 I_50573 (I862252,I2507,I861828,I861799,);
nor I_50574 (I862283,I862131,I862187);
not I_50575 (I862300,I862283);
nand I_50576 (I861808,I862300,I862156);
not I_50577 (I862355,I2514);
DFFARX1 I_50578 (I1028663,I2507,I862355,I862381,);
not I_50579 (I862389,I862381);
nand I_50580 (I862406,I1028672,I1028660);
and I_50581 (I862423,I862406,I1028657);
DFFARX1 I_50582 (I862423,I2507,I862355,I862449,);
DFFARX1 I_50583 (I862449,I2507,I862355,I862344,);
DFFARX1 I_50584 (I1028657,I2507,I862355,I862480,);
nand I_50585 (I862488,I862480,I1028654);
not I_50586 (I862505,I862488);
DFFARX1 I_50587 (I862505,I2507,I862355,I862531,);
not I_50588 (I862539,I862531);
nor I_50589 (I862347,I862389,I862539);
DFFARX1 I_50590 (I1028660,I2507,I862355,I862579,);
nor I_50591 (I862338,I862579,I862449);
nor I_50592 (I862329,I862579,I862505);
nand I_50593 (I862615,I1028675,I1028666);
and I_50594 (I862632,I862615,I1028669);
DFFARX1 I_50595 (I862632,I2507,I862355,I862658,);
not I_50596 (I862666,I862658);
nand I_50597 (I862683,I862666,I862579);
nand I_50598 (I862332,I862666,I862488);
nor I_50599 (I862714,I1028654,I1028666);
and I_50600 (I862731,I862579,I862714);
nor I_50601 (I862748,I862666,I862731);
DFFARX1 I_50602 (I862748,I2507,I862355,I862341,);
nor I_50603 (I862779,I862381,I862714);
DFFARX1 I_50604 (I862779,I2507,I862355,I862326,);
nor I_50605 (I862810,I862658,I862714);
not I_50606 (I862827,I862810);
nand I_50607 (I862335,I862827,I862683);
not I_50608 (I862882,I2514);
DFFARX1 I_50609 (I6697,I2507,I862882,I862908,);
not I_50610 (I862916,I862908);
nand I_50611 (I862933,I6703,I6685);
and I_50612 (I862950,I862933,I6694);
DFFARX1 I_50613 (I862950,I2507,I862882,I862976,);
DFFARX1 I_50614 (I862976,I2507,I862882,I862871,);
DFFARX1 I_50615 (I6685,I2507,I862882,I863007,);
nand I_50616 (I863015,I863007,I6688);
not I_50617 (I863032,I863015);
DFFARX1 I_50618 (I863032,I2507,I862882,I863058,);
not I_50619 (I863066,I863058);
nor I_50620 (I862874,I862916,I863066);
DFFARX1 I_50621 (I6688,I2507,I862882,I863106,);
nor I_50622 (I862865,I863106,I862976);
nor I_50623 (I862856,I863106,I863032);
nand I_50624 (I863142,I6691,I6700);
and I_50625 (I863159,I863142,I6682);
DFFARX1 I_50626 (I863159,I2507,I862882,I863185,);
not I_50627 (I863193,I863185);
nand I_50628 (I863210,I863193,I863106);
nand I_50629 (I862859,I863193,I863015);
nor I_50630 (I863241,I6682,I6700);
and I_50631 (I863258,I863106,I863241);
nor I_50632 (I863275,I863193,I863258);
DFFARX1 I_50633 (I863275,I2507,I862882,I862868,);
nor I_50634 (I863306,I862908,I863241);
DFFARX1 I_50635 (I863306,I2507,I862882,I862853,);
nor I_50636 (I863337,I863185,I863241);
not I_50637 (I863354,I863337);
nand I_50638 (I862862,I863354,I863210);
not I_50639 (I863409,I2514);
DFFARX1 I_50640 (I463733,I2507,I863409,I863435,);
not I_50641 (I863443,I863435);
nand I_50642 (I863460,I463730,I463739);
and I_50643 (I863477,I863460,I463748);
DFFARX1 I_50644 (I863477,I2507,I863409,I863503,);
DFFARX1 I_50645 (I863503,I2507,I863409,I863398,);
DFFARX1 I_50646 (I463751,I2507,I863409,I863534,);
nand I_50647 (I863542,I863534,I463754);
not I_50648 (I863559,I863542);
DFFARX1 I_50649 (I863559,I2507,I863409,I863585,);
not I_50650 (I863593,I863585);
nor I_50651 (I863401,I863443,I863593);
DFFARX1 I_50652 (I463727,I2507,I863409,I863633,);
nor I_50653 (I863392,I863633,I863503);
nor I_50654 (I863383,I863633,I863559);
nand I_50655 (I863669,I463742,I463745);
and I_50656 (I863686,I863669,I463736);
DFFARX1 I_50657 (I863686,I2507,I863409,I863712,);
not I_50658 (I863720,I863712);
nand I_50659 (I863737,I863720,I863633);
nand I_50660 (I863386,I863720,I863542);
nor I_50661 (I863768,I463727,I463745);
and I_50662 (I863785,I863633,I863768);
nor I_50663 (I863802,I863720,I863785);
DFFARX1 I_50664 (I863802,I2507,I863409,I863395,);
nor I_50665 (I863833,I863435,I863768);
DFFARX1 I_50666 (I863833,I2507,I863409,I863380,);
nor I_50667 (I863864,I863712,I863768);
not I_50668 (I863881,I863864);
nand I_50669 (I863389,I863881,I863737);
not I_50670 (I863936,I2514);
DFFARX1 I_50671 (I1301986,I2507,I863936,I863962,);
not I_50672 (I863970,I863962);
nand I_50673 (I863987,I1301980,I1301998);
and I_50674 (I864004,I863987,I1301983);
DFFARX1 I_50675 (I864004,I2507,I863936,I864030,);
DFFARX1 I_50676 (I864030,I2507,I863936,I863925,);
DFFARX1 I_50677 (I1302004,I2507,I863936,I864061,);
nand I_50678 (I864069,I864061,I1301989);
not I_50679 (I864086,I864069);
DFFARX1 I_50680 (I864086,I2507,I863936,I864112,);
not I_50681 (I864120,I864112);
nor I_50682 (I863928,I863970,I864120);
DFFARX1 I_50683 (I1302001,I2507,I863936,I864160,);
nor I_50684 (I863919,I864160,I864030);
nor I_50685 (I863910,I864160,I864086);
nand I_50686 (I864196,I1301992,I1302007);
and I_50687 (I864213,I864196,I1301995);
DFFARX1 I_50688 (I864213,I2507,I863936,I864239,);
not I_50689 (I864247,I864239);
nand I_50690 (I864264,I864247,I864160);
nand I_50691 (I863913,I864247,I864069);
nor I_50692 (I864295,I1301980,I1302007);
and I_50693 (I864312,I864160,I864295);
nor I_50694 (I864329,I864247,I864312);
DFFARX1 I_50695 (I864329,I2507,I863936,I863922,);
nor I_50696 (I864360,I863962,I864295);
DFFARX1 I_50697 (I864360,I2507,I863936,I863907,);
nor I_50698 (I864391,I864239,I864295);
not I_50699 (I864408,I864391);
nand I_50700 (I863916,I864408,I864264);
not I_50701 (I864463,I2514);
DFFARX1 I_50702 (I1249326,I2507,I864463,I864489,);
not I_50703 (I864497,I864489);
nand I_50704 (I864514,I1249332,I1249314);
and I_50705 (I864531,I864514,I1249323);
DFFARX1 I_50706 (I864531,I2507,I864463,I864557,);
DFFARX1 I_50707 (I864557,I2507,I864463,I864452,);
DFFARX1 I_50708 (I1249329,I2507,I864463,I864588,);
nand I_50709 (I864596,I864588,I1249317);
not I_50710 (I864613,I864596);
DFFARX1 I_50711 (I864613,I2507,I864463,I864639,);
not I_50712 (I864647,I864639);
nor I_50713 (I864455,I864497,I864647);
DFFARX1 I_50714 (I1249335,I2507,I864463,I864687,);
nor I_50715 (I864446,I864687,I864557);
nor I_50716 (I864437,I864687,I864613);
nand I_50717 (I864723,I1249314,I1249320);
and I_50718 (I864740,I864723,I1249338);
DFFARX1 I_50719 (I864740,I2507,I864463,I864766,);
not I_50720 (I864774,I864766);
nand I_50721 (I864791,I864774,I864687);
nand I_50722 (I864440,I864774,I864596);
nor I_50723 (I864822,I1249317,I1249320);
and I_50724 (I864839,I864687,I864822);
nor I_50725 (I864856,I864774,I864839);
DFFARX1 I_50726 (I864856,I2507,I864463,I864449,);
nor I_50727 (I864887,I864489,I864822);
DFFARX1 I_50728 (I864887,I2507,I864463,I864434,);
nor I_50729 (I864918,I864766,I864822);
not I_50730 (I864935,I864918);
nand I_50731 (I864443,I864935,I864791);
not I_50732 (I864990,I2514);
DFFARX1 I_50733 (I656150,I2507,I864990,I865016,);
not I_50734 (I865024,I865016);
nand I_50735 (I865041,I656153,I656150);
and I_50736 (I865058,I865041,I656162);
DFFARX1 I_50737 (I865058,I2507,I864990,I865084,);
DFFARX1 I_50738 (I865084,I2507,I864990,I864979,);
DFFARX1 I_50739 (I656159,I2507,I864990,I865115,);
nand I_50740 (I865123,I865115,I656165);
not I_50741 (I865140,I865123);
DFFARX1 I_50742 (I865140,I2507,I864990,I865166,);
not I_50743 (I865174,I865166);
nor I_50744 (I864982,I865024,I865174);
DFFARX1 I_50745 (I656174,I2507,I864990,I865214,);
nor I_50746 (I864973,I865214,I865084);
nor I_50747 (I864964,I865214,I865140);
nand I_50748 (I865250,I656168,I656156);
and I_50749 (I865267,I865250,I656153);
DFFARX1 I_50750 (I865267,I2507,I864990,I865293,);
not I_50751 (I865301,I865293);
nand I_50752 (I865318,I865301,I865214);
nand I_50753 (I864967,I865301,I865123);
nor I_50754 (I865349,I656171,I656156);
and I_50755 (I865366,I865214,I865349);
nor I_50756 (I865383,I865301,I865366);
DFFARX1 I_50757 (I865383,I2507,I864990,I864976,);
nor I_50758 (I865414,I865016,I865349);
DFFARX1 I_50759 (I865414,I2507,I864990,I864961,);
nor I_50760 (I865445,I865293,I865349);
not I_50761 (I865462,I865445);
nand I_50762 (I864970,I865462,I865318);
not I_50763 (I865517,I2514);
DFFARX1 I_50764 (I1193640,I2507,I865517,I865543,);
not I_50765 (I865551,I865543);
nand I_50766 (I865568,I1193622,I1193622);
and I_50767 (I865585,I865568,I1193628);
DFFARX1 I_50768 (I865585,I2507,I865517,I865611,);
DFFARX1 I_50769 (I865611,I2507,I865517,I865506,);
DFFARX1 I_50770 (I1193625,I2507,I865517,I865642,);
nand I_50771 (I865650,I865642,I1193634);
not I_50772 (I865667,I865650);
DFFARX1 I_50773 (I865667,I2507,I865517,I865693,);
not I_50774 (I865701,I865693);
nor I_50775 (I865509,I865551,I865701);
DFFARX1 I_50776 (I1193646,I2507,I865517,I865741,);
nor I_50777 (I865500,I865741,I865611);
nor I_50778 (I865491,I865741,I865667);
nand I_50779 (I865777,I1193637,I1193631);
and I_50780 (I865794,I865777,I1193625);
DFFARX1 I_50781 (I865794,I2507,I865517,I865820,);
not I_50782 (I865828,I865820);
nand I_50783 (I865845,I865828,I865741);
nand I_50784 (I865494,I865828,I865650);
nor I_50785 (I865876,I1193643,I1193631);
and I_50786 (I865893,I865741,I865876);
nor I_50787 (I865910,I865828,I865893);
DFFARX1 I_50788 (I865910,I2507,I865517,I865503,);
nor I_50789 (I865941,I865543,I865876);
DFFARX1 I_50790 (I865941,I2507,I865517,I865488,);
nor I_50791 (I865972,I865820,I865876);
not I_50792 (I865989,I865972);
nand I_50793 (I865497,I865989,I865845);
not I_50794 (I866044,I2514);
DFFARX1 I_50795 (I116016,I2507,I866044,I866070,);
not I_50796 (I866078,I866070);
nand I_50797 (I866095,I115992,I116001);
and I_50798 (I866112,I866095,I115995);
DFFARX1 I_50799 (I866112,I2507,I866044,I866138,);
DFFARX1 I_50800 (I866138,I2507,I866044,I866033,);
DFFARX1 I_50801 (I116013,I2507,I866044,I866169,);
nand I_50802 (I866177,I866169,I116004);
not I_50803 (I866194,I866177);
DFFARX1 I_50804 (I866194,I2507,I866044,I866220,);
not I_50805 (I866228,I866220);
nor I_50806 (I866036,I866078,I866228);
DFFARX1 I_50807 (I115998,I2507,I866044,I866268,);
nor I_50808 (I866027,I866268,I866138);
nor I_50809 (I866018,I866268,I866194);
nand I_50810 (I866304,I116010,I116007);
and I_50811 (I866321,I866304,I115995);
DFFARX1 I_50812 (I866321,I2507,I866044,I866347,);
not I_50813 (I866355,I866347);
nand I_50814 (I866372,I866355,I866268);
nand I_50815 (I866021,I866355,I866177);
nor I_50816 (I866403,I115992,I116007);
and I_50817 (I866420,I866268,I866403);
nor I_50818 (I866437,I866355,I866420);
DFFARX1 I_50819 (I866437,I2507,I866044,I866030,);
nor I_50820 (I866468,I866070,I866403);
DFFARX1 I_50821 (I866468,I2507,I866044,I866015,);
nor I_50822 (I866499,I866347,I866403);
not I_50823 (I866516,I866499);
nand I_50824 (I866024,I866516,I866372);
not I_50825 (I866571,I2514);
DFFARX1 I_50826 (I1131216,I2507,I866571,I866597,);
not I_50827 (I866605,I866597);
nand I_50828 (I866622,I1131198,I1131198);
and I_50829 (I866639,I866622,I1131204);
DFFARX1 I_50830 (I866639,I2507,I866571,I866665,);
DFFARX1 I_50831 (I866665,I2507,I866571,I866560,);
DFFARX1 I_50832 (I1131201,I2507,I866571,I866696,);
nand I_50833 (I866704,I866696,I1131210);
not I_50834 (I866721,I866704);
DFFARX1 I_50835 (I866721,I2507,I866571,I866747,);
not I_50836 (I866755,I866747);
nor I_50837 (I866563,I866605,I866755);
DFFARX1 I_50838 (I1131222,I2507,I866571,I866795,);
nor I_50839 (I866554,I866795,I866665);
nor I_50840 (I866545,I866795,I866721);
nand I_50841 (I866831,I1131213,I1131207);
and I_50842 (I866848,I866831,I1131201);
DFFARX1 I_50843 (I866848,I2507,I866571,I866874,);
not I_50844 (I866882,I866874);
nand I_50845 (I866899,I866882,I866795);
nand I_50846 (I866548,I866882,I866704);
nor I_50847 (I866930,I1131219,I1131207);
and I_50848 (I866947,I866795,I866930);
nor I_50849 (I866964,I866882,I866947);
DFFARX1 I_50850 (I866964,I2507,I866571,I866557,);
nor I_50851 (I866995,I866597,I866930);
DFFARX1 I_50852 (I866995,I2507,I866571,I866542,);
nor I_50853 (I867026,I866874,I866930);
not I_50854 (I867043,I867026);
nand I_50855 (I866551,I867043,I866899);
not I_50856 (I867098,I2514);
DFFARX1 I_50857 (I336100,I2507,I867098,I867124,);
not I_50858 (I867132,I867124);
nand I_50859 (I867149,I336091,I336091);
and I_50860 (I867166,I867149,I336109);
DFFARX1 I_50861 (I867166,I2507,I867098,I867192,);
DFFARX1 I_50862 (I867192,I2507,I867098,I867087,);
DFFARX1 I_50863 (I336112,I2507,I867098,I867223,);
nand I_50864 (I867231,I867223,I336094);
not I_50865 (I867248,I867231);
DFFARX1 I_50866 (I867248,I2507,I867098,I867274,);
not I_50867 (I867282,I867274);
nor I_50868 (I867090,I867132,I867282);
DFFARX1 I_50869 (I336106,I2507,I867098,I867322,);
nor I_50870 (I867081,I867322,I867192);
nor I_50871 (I867072,I867322,I867248);
nand I_50872 (I867358,I336118,I336097);
and I_50873 (I867375,I867358,I336103);
DFFARX1 I_50874 (I867375,I2507,I867098,I867401,);
not I_50875 (I867409,I867401);
nand I_50876 (I867426,I867409,I867322);
nand I_50877 (I867075,I867409,I867231);
nor I_50878 (I867457,I336115,I336097);
and I_50879 (I867474,I867322,I867457);
nor I_50880 (I867491,I867409,I867474);
DFFARX1 I_50881 (I867491,I2507,I867098,I867084,);
nor I_50882 (I867522,I867124,I867457);
DFFARX1 I_50883 (I867522,I2507,I867098,I867069,);
nor I_50884 (I867553,I867401,I867457);
not I_50885 (I867570,I867553);
nand I_50886 (I867078,I867570,I867426);
not I_50887 (I867625,I2514);
DFFARX1 I_50888 (I571777,I2507,I867625,I867651,);
not I_50889 (I867659,I867651);
nand I_50890 (I867676,I571762,I571783);
and I_50891 (I867693,I867676,I571771);
DFFARX1 I_50892 (I867693,I2507,I867625,I867719,);
DFFARX1 I_50893 (I867719,I2507,I867625,I867614,);
DFFARX1 I_50894 (I571765,I2507,I867625,I867750,);
nand I_50895 (I867758,I867750,I571774);
not I_50896 (I867775,I867758);
DFFARX1 I_50897 (I867775,I2507,I867625,I867801,);
not I_50898 (I867809,I867801);
nor I_50899 (I867617,I867659,I867809);
DFFARX1 I_50900 (I571780,I2507,I867625,I867849,);
nor I_50901 (I867608,I867849,I867719);
nor I_50902 (I867599,I867849,I867775);
nand I_50903 (I867885,I571762,I571765);
and I_50904 (I867902,I867885,I571786);
DFFARX1 I_50905 (I867902,I2507,I867625,I867928,);
not I_50906 (I867936,I867928);
nand I_50907 (I867953,I867936,I867849);
nand I_50908 (I867602,I867936,I867758);
nor I_50909 (I867984,I571768,I571765);
and I_50910 (I868001,I867849,I867984);
nor I_50911 (I868018,I867936,I868001);
DFFARX1 I_50912 (I868018,I2507,I867625,I867611,);
nor I_50913 (I868049,I867651,I867984);
DFFARX1 I_50914 (I868049,I2507,I867625,I867596,);
nor I_50915 (I868080,I867928,I867984);
not I_50916 (I868097,I868080);
nand I_50917 (I867605,I868097,I867953);
not I_50918 (I868152,I2514);
DFFARX1 I_50919 (I215686,I2507,I868152,I868178,);
not I_50920 (I868186,I868178);
nand I_50921 (I868203,I215683,I215701);
and I_50922 (I868220,I868203,I215692);
DFFARX1 I_50923 (I868220,I2507,I868152,I868246,);
DFFARX1 I_50924 (I868246,I2507,I868152,I868141,);
DFFARX1 I_50925 (I215698,I2507,I868152,I868277,);
nand I_50926 (I868285,I868277,I215695);
not I_50927 (I868302,I868285);
DFFARX1 I_50928 (I868302,I2507,I868152,I868328,);
not I_50929 (I868336,I868328);
nor I_50930 (I868144,I868186,I868336);
DFFARX1 I_50931 (I215689,I2507,I868152,I868376,);
nor I_50932 (I868135,I868376,I868246);
nor I_50933 (I868126,I868376,I868302);
nand I_50934 (I868412,I215680,I215704);
and I_50935 (I868429,I868412,I215683);
DFFARX1 I_50936 (I868429,I2507,I868152,I868455,);
not I_50937 (I868463,I868455);
nand I_50938 (I868480,I868463,I868376);
nand I_50939 (I868129,I868463,I868285);
nor I_50940 (I868511,I215680,I215704);
and I_50941 (I868528,I868376,I868511);
nor I_50942 (I868545,I868463,I868528);
DFFARX1 I_50943 (I868545,I2507,I868152,I868138,);
nor I_50944 (I868576,I868178,I868511);
DFFARX1 I_50945 (I868576,I2507,I868152,I868123,);
nor I_50946 (I868607,I868455,I868511);
not I_50947 (I868624,I868607);
nand I_50948 (I868132,I868624,I868480);
not I_50949 (I868679,I2514);
DFFARX1 I_50950 (I1371372,I2507,I868679,I868705,);
not I_50951 (I868713,I868705);
nand I_50952 (I868730,I1371369,I1371378);
and I_50953 (I868747,I868730,I1371357);
DFFARX1 I_50954 (I868747,I2507,I868679,I868773,);
DFFARX1 I_50955 (I868773,I2507,I868679,I868668,);
DFFARX1 I_50956 (I1371360,I2507,I868679,I868804,);
nand I_50957 (I868812,I868804,I1371375);
not I_50958 (I868829,I868812);
DFFARX1 I_50959 (I868829,I2507,I868679,I868855,);
not I_50960 (I868863,I868855);
nor I_50961 (I868671,I868713,I868863);
DFFARX1 I_50962 (I1371381,I2507,I868679,I868903,);
nor I_50963 (I868662,I868903,I868773);
nor I_50964 (I868653,I868903,I868829);
nand I_50965 (I868939,I1371363,I1371384);
and I_50966 (I868956,I868939,I1371366);
DFFARX1 I_50967 (I868956,I2507,I868679,I868982,);
not I_50968 (I868990,I868982);
nand I_50969 (I869007,I868990,I868903);
nand I_50970 (I868656,I868990,I868812);
nor I_50971 (I869038,I1371357,I1371384);
and I_50972 (I869055,I868903,I869038);
nor I_50973 (I869072,I868990,I869055);
DFFARX1 I_50974 (I869072,I2507,I868679,I868665,);
nor I_50975 (I869103,I868705,I869038);
DFFARX1 I_50976 (I869103,I2507,I868679,I868650,);
nor I_50977 (I869134,I868982,I869038);
not I_50978 (I869151,I869134);
nand I_50979 (I868659,I869151,I869007);
not I_50980 (I869206,I2514);
DFFARX1 I_50981 (I339262,I2507,I869206,I869232,);
not I_50982 (I869240,I869232);
nand I_50983 (I869257,I339253,I339253);
and I_50984 (I869274,I869257,I339271);
DFFARX1 I_50985 (I869274,I2507,I869206,I869300,);
DFFARX1 I_50986 (I869300,I2507,I869206,I869195,);
DFFARX1 I_50987 (I339274,I2507,I869206,I869331,);
nand I_50988 (I869339,I869331,I339256);
not I_50989 (I869356,I869339);
DFFARX1 I_50990 (I869356,I2507,I869206,I869382,);
not I_50991 (I869390,I869382);
nor I_50992 (I869198,I869240,I869390);
DFFARX1 I_50993 (I339268,I2507,I869206,I869430,);
nor I_50994 (I869189,I869430,I869300);
nor I_50995 (I869180,I869430,I869356);
nand I_50996 (I869466,I339280,I339259);
and I_50997 (I869483,I869466,I339265);
DFFARX1 I_50998 (I869483,I2507,I869206,I869509,);
not I_50999 (I869517,I869509);
nand I_51000 (I869534,I869517,I869430);
nand I_51001 (I869183,I869517,I869339);
nor I_51002 (I869565,I339277,I339259);
and I_51003 (I869582,I869430,I869565);
nor I_51004 (I869599,I869517,I869582);
DFFARX1 I_51005 (I869599,I2507,I869206,I869192,);
nor I_51006 (I869630,I869232,I869565);
DFFARX1 I_51007 (I869630,I2507,I869206,I869177,);
nor I_51008 (I869661,I869509,I869565);
not I_51009 (I869678,I869661);
nand I_51010 (I869186,I869678,I869534);
not I_51011 (I869733,I2514);
DFFARX1 I_51012 (I173441,I2507,I869733,I869759,);
not I_51013 (I869767,I869759);
nand I_51014 (I869784,I173438,I173456);
and I_51015 (I869801,I869784,I173447);
DFFARX1 I_51016 (I869801,I2507,I869733,I869827,);
DFFARX1 I_51017 (I869827,I2507,I869733,I869722,);
DFFARX1 I_51018 (I173453,I2507,I869733,I869858,);
nand I_51019 (I869866,I869858,I173450);
not I_51020 (I869883,I869866);
DFFARX1 I_51021 (I869883,I2507,I869733,I869909,);
not I_51022 (I869917,I869909);
nor I_51023 (I869725,I869767,I869917);
DFFARX1 I_51024 (I173444,I2507,I869733,I869957,);
nor I_51025 (I869716,I869957,I869827);
nor I_51026 (I869707,I869957,I869883);
nand I_51027 (I869993,I173435,I173459);
and I_51028 (I870010,I869993,I173438);
DFFARX1 I_51029 (I870010,I2507,I869733,I870036,);
not I_51030 (I870044,I870036);
nand I_51031 (I870061,I870044,I869957);
nand I_51032 (I869710,I870044,I869866);
nor I_51033 (I870092,I173435,I173459);
and I_51034 (I870109,I869957,I870092);
nor I_51035 (I870126,I870044,I870109);
DFFARX1 I_51036 (I870126,I2507,I869733,I869719,);
nor I_51037 (I870157,I869759,I870092);
DFFARX1 I_51038 (I870157,I2507,I869733,I869704,);
nor I_51039 (I870188,I870036,I870092);
not I_51040 (I870205,I870188);
nand I_51041 (I869713,I870205,I870061);
not I_51042 (I870260,I2514);
DFFARX1 I_51043 (I578713,I2507,I870260,I870286,);
not I_51044 (I870294,I870286);
nand I_51045 (I870311,I578698,I578719);
and I_51046 (I870328,I870311,I578707);
DFFARX1 I_51047 (I870328,I2507,I870260,I870354,);
DFFARX1 I_51048 (I870354,I2507,I870260,I870249,);
DFFARX1 I_51049 (I578701,I2507,I870260,I870385,);
nand I_51050 (I870393,I870385,I578710);
not I_51051 (I870410,I870393);
DFFARX1 I_51052 (I870410,I2507,I870260,I870436,);
not I_51053 (I870444,I870436);
nor I_51054 (I870252,I870294,I870444);
DFFARX1 I_51055 (I578716,I2507,I870260,I870484,);
nor I_51056 (I870243,I870484,I870354);
nor I_51057 (I870234,I870484,I870410);
nand I_51058 (I870520,I578698,I578701);
and I_51059 (I870537,I870520,I578722);
DFFARX1 I_51060 (I870537,I2507,I870260,I870563,);
not I_51061 (I870571,I870563);
nand I_51062 (I870588,I870571,I870484);
nand I_51063 (I870237,I870571,I870393);
nor I_51064 (I870619,I578704,I578701);
and I_51065 (I870636,I870484,I870619);
nor I_51066 (I870653,I870571,I870636);
DFFARX1 I_51067 (I870653,I2507,I870260,I870246,);
nor I_51068 (I870684,I870286,I870619);
DFFARX1 I_51069 (I870684,I2507,I870260,I870231,);
nor I_51070 (I870715,I870563,I870619);
not I_51071 (I870732,I870715);
nand I_51072 (I870240,I870732,I870588);
not I_51073 (I870787,I2514);
DFFARX1 I_51074 (I623797,I2507,I870787,I870813,);
not I_51075 (I870821,I870813);
nand I_51076 (I870838,I623782,I623803);
and I_51077 (I870855,I870838,I623791);
DFFARX1 I_51078 (I870855,I2507,I870787,I870881,);
DFFARX1 I_51079 (I870881,I2507,I870787,I870776,);
DFFARX1 I_51080 (I623785,I2507,I870787,I870912,);
nand I_51081 (I870920,I870912,I623794);
not I_51082 (I870937,I870920);
DFFARX1 I_51083 (I870937,I2507,I870787,I870963,);
not I_51084 (I870971,I870963);
nor I_51085 (I870779,I870821,I870971);
DFFARX1 I_51086 (I623800,I2507,I870787,I871011,);
nor I_51087 (I870770,I871011,I870881);
nor I_51088 (I870761,I871011,I870937);
nand I_51089 (I871047,I623782,I623785);
and I_51090 (I871064,I871047,I623806);
DFFARX1 I_51091 (I871064,I2507,I870787,I871090,);
not I_51092 (I871098,I871090);
nand I_51093 (I871115,I871098,I871011);
nand I_51094 (I870764,I871098,I870920);
nor I_51095 (I871146,I623788,I623785);
and I_51096 (I871163,I871011,I871146);
nor I_51097 (I871180,I871098,I871163);
DFFARX1 I_51098 (I871180,I2507,I870787,I870773,);
nor I_51099 (I871211,I870813,I871146);
DFFARX1 I_51100 (I871211,I2507,I870787,I870758,);
nor I_51101 (I871242,I871090,I871146);
not I_51102 (I871259,I871242);
nand I_51103 (I870767,I871259,I871115);
not I_51104 (I871314,I2514);
DFFARX1 I_51105 (I1055591,I2507,I871314,I871340,);
not I_51106 (I871348,I871340);
nand I_51107 (I871365,I1055600,I1055588);
and I_51108 (I871382,I871365,I1055585);
DFFARX1 I_51109 (I871382,I2507,I871314,I871408,);
DFFARX1 I_51110 (I871408,I2507,I871314,I871303,);
DFFARX1 I_51111 (I1055585,I2507,I871314,I871439,);
nand I_51112 (I871447,I871439,I1055582);
not I_51113 (I871464,I871447);
DFFARX1 I_51114 (I871464,I2507,I871314,I871490,);
not I_51115 (I871498,I871490);
nor I_51116 (I871306,I871348,I871498);
DFFARX1 I_51117 (I1055588,I2507,I871314,I871538,);
nor I_51118 (I871297,I871538,I871408);
nor I_51119 (I871288,I871538,I871464);
nand I_51120 (I871574,I1055603,I1055594);
and I_51121 (I871591,I871574,I1055597);
DFFARX1 I_51122 (I871591,I2507,I871314,I871617,);
not I_51123 (I871625,I871617);
nand I_51124 (I871642,I871625,I871538);
nand I_51125 (I871291,I871625,I871447);
nor I_51126 (I871673,I1055582,I1055594);
and I_51127 (I871690,I871538,I871673);
nor I_51128 (I871707,I871625,I871690);
DFFARX1 I_51129 (I871707,I2507,I871314,I871300,);
nor I_51130 (I871738,I871340,I871673);
DFFARX1 I_51131 (I871738,I2507,I871314,I871285,);
nor I_51132 (I871769,I871617,I871673);
not I_51133 (I871786,I871769);
nand I_51134 (I871294,I871786,I871642);
not I_51135 (I871841,I2514);
DFFARX1 I_51136 (I193076,I2507,I871841,I871867,);
not I_51137 (I871875,I871867);
nand I_51138 (I871892,I193073,I193091);
and I_51139 (I871909,I871892,I193082);
DFFARX1 I_51140 (I871909,I2507,I871841,I871935,);
DFFARX1 I_51141 (I871935,I2507,I871841,I871830,);
DFFARX1 I_51142 (I193088,I2507,I871841,I871966,);
nand I_51143 (I871974,I871966,I193085);
not I_51144 (I871991,I871974);
DFFARX1 I_51145 (I871991,I2507,I871841,I872017,);
not I_51146 (I872025,I872017);
nor I_51147 (I871833,I871875,I872025);
DFFARX1 I_51148 (I193079,I2507,I871841,I872065,);
nor I_51149 (I871824,I872065,I871935);
nor I_51150 (I871815,I872065,I871991);
nand I_51151 (I872101,I193070,I193094);
and I_51152 (I872118,I872101,I193073);
DFFARX1 I_51153 (I872118,I2507,I871841,I872144,);
not I_51154 (I872152,I872144);
nand I_51155 (I872169,I872152,I872065);
nand I_51156 (I871818,I872152,I871974);
nor I_51157 (I872200,I193070,I193094);
and I_51158 (I872217,I872065,I872200);
nor I_51159 (I872234,I872152,I872217);
DFFARX1 I_51160 (I872234,I2507,I871841,I871827,);
nor I_51161 (I872265,I871867,I872200);
DFFARX1 I_51162 (I872265,I2507,I871841,I871812,);
nor I_51163 (I872296,I872144,I872200);
not I_51164 (I872313,I872296);
nand I_51165 (I871821,I872313,I872169);
not I_51166 (I872368,I2514);
DFFARX1 I_51167 (I655572,I2507,I872368,I872394,);
not I_51168 (I872402,I872394);
nand I_51169 (I872419,I655575,I655572);
and I_51170 (I872436,I872419,I655584);
DFFARX1 I_51171 (I872436,I2507,I872368,I872462,);
DFFARX1 I_51172 (I872462,I2507,I872368,I872357,);
DFFARX1 I_51173 (I655581,I2507,I872368,I872493,);
nand I_51174 (I872501,I872493,I655587);
not I_51175 (I872518,I872501);
DFFARX1 I_51176 (I872518,I2507,I872368,I872544,);
not I_51177 (I872552,I872544);
nor I_51178 (I872360,I872402,I872552);
DFFARX1 I_51179 (I655596,I2507,I872368,I872592,);
nor I_51180 (I872351,I872592,I872462);
nor I_51181 (I872342,I872592,I872518);
nand I_51182 (I872628,I655590,I655578);
and I_51183 (I872645,I872628,I655575);
DFFARX1 I_51184 (I872645,I2507,I872368,I872671,);
not I_51185 (I872679,I872671);
nand I_51186 (I872696,I872679,I872592);
nand I_51187 (I872345,I872679,I872501);
nor I_51188 (I872727,I655593,I655578);
and I_51189 (I872744,I872592,I872727);
nor I_51190 (I872761,I872679,I872744);
DFFARX1 I_51191 (I872761,I2507,I872368,I872354,);
nor I_51192 (I872792,I872394,I872727);
DFFARX1 I_51193 (I872792,I2507,I872368,I872339,);
nor I_51194 (I872823,I872671,I872727);
not I_51195 (I872840,I872823);
nand I_51196 (I872348,I872840,I872696);
not I_51197 (I872895,I2514);
DFFARX1 I_51198 (I684472,I2507,I872895,I872921,);
not I_51199 (I872929,I872921);
nand I_51200 (I872946,I684475,I684472);
and I_51201 (I872963,I872946,I684484);
DFFARX1 I_51202 (I872963,I2507,I872895,I872989,);
DFFARX1 I_51203 (I872989,I2507,I872895,I872884,);
DFFARX1 I_51204 (I684481,I2507,I872895,I873020,);
nand I_51205 (I873028,I873020,I684487);
not I_51206 (I873045,I873028);
DFFARX1 I_51207 (I873045,I2507,I872895,I873071,);
not I_51208 (I873079,I873071);
nor I_51209 (I872887,I872929,I873079);
DFFARX1 I_51210 (I684496,I2507,I872895,I873119,);
nor I_51211 (I872878,I873119,I872989);
nor I_51212 (I872869,I873119,I873045);
nand I_51213 (I873155,I684490,I684478);
and I_51214 (I873172,I873155,I684475);
DFFARX1 I_51215 (I873172,I2507,I872895,I873198,);
not I_51216 (I873206,I873198);
nand I_51217 (I873223,I873206,I873119);
nand I_51218 (I872872,I873206,I873028);
nor I_51219 (I873254,I684493,I684478);
and I_51220 (I873271,I873119,I873254);
nor I_51221 (I873288,I873206,I873271);
DFFARX1 I_51222 (I873288,I2507,I872895,I872881,);
nor I_51223 (I873319,I872921,I873254);
DFFARX1 I_51224 (I873319,I2507,I872895,I872866,);
nor I_51225 (I873350,I873198,I873254);
not I_51226 (I873367,I873350);
nand I_51227 (I872875,I873367,I873223);
not I_51228 (I873422,I2514);
DFFARX1 I_51229 (I962510,I2507,I873422,I873448,);
not I_51230 (I873456,I873448);
nand I_51231 (I873473,I962525,I962507);
and I_51232 (I873490,I873473,I962507);
DFFARX1 I_51233 (I873490,I2507,I873422,I873516,);
DFFARX1 I_51234 (I873516,I2507,I873422,I873411,);
DFFARX1 I_51235 (I962516,I2507,I873422,I873547,);
nand I_51236 (I873555,I873547,I962534);
not I_51237 (I873572,I873555);
DFFARX1 I_51238 (I873572,I2507,I873422,I873598,);
not I_51239 (I873606,I873598);
nor I_51240 (I873414,I873456,I873606);
DFFARX1 I_51241 (I962531,I2507,I873422,I873646,);
nor I_51242 (I873405,I873646,I873516);
nor I_51243 (I873396,I873646,I873572);
nand I_51244 (I873682,I962528,I962519);
and I_51245 (I873699,I873682,I962513);
DFFARX1 I_51246 (I873699,I2507,I873422,I873725,);
not I_51247 (I873733,I873725);
nand I_51248 (I873750,I873733,I873646);
nand I_51249 (I873399,I873733,I873555);
nor I_51250 (I873781,I962522,I962519);
and I_51251 (I873798,I873646,I873781);
nor I_51252 (I873815,I873733,I873798);
DFFARX1 I_51253 (I873815,I2507,I873422,I873408,);
nor I_51254 (I873846,I873448,I873781);
DFFARX1 I_51255 (I873846,I2507,I873422,I873393,);
nor I_51256 (I873877,I873725,I873781);
not I_51257 (I873894,I873877);
nand I_51258 (I873402,I873894,I873750);
not I_51259 (I873949,I2514);
DFFARX1 I_51260 (I1361852,I2507,I873949,I873975,);
not I_51261 (I873983,I873975);
nand I_51262 (I874000,I1361849,I1361858);
and I_51263 (I874017,I874000,I1361837);
DFFARX1 I_51264 (I874017,I2507,I873949,I874043,);
DFFARX1 I_51265 (I874043,I2507,I873949,I873938,);
DFFARX1 I_51266 (I1361840,I2507,I873949,I874074,);
nand I_51267 (I874082,I874074,I1361855);
not I_51268 (I874099,I874082);
DFFARX1 I_51269 (I874099,I2507,I873949,I874125,);
not I_51270 (I874133,I874125);
nor I_51271 (I873941,I873983,I874133);
DFFARX1 I_51272 (I1361861,I2507,I873949,I874173,);
nor I_51273 (I873932,I874173,I874043);
nor I_51274 (I873923,I874173,I874099);
nand I_51275 (I874209,I1361843,I1361864);
and I_51276 (I874226,I874209,I1361846);
DFFARX1 I_51277 (I874226,I2507,I873949,I874252,);
not I_51278 (I874260,I874252);
nand I_51279 (I874277,I874260,I874173);
nand I_51280 (I873926,I874260,I874082);
nor I_51281 (I874308,I1361837,I1361864);
and I_51282 (I874325,I874173,I874308);
nor I_51283 (I874342,I874260,I874325);
DFFARX1 I_51284 (I874342,I2507,I873949,I873935,);
nor I_51285 (I874373,I873975,I874308);
DFFARX1 I_51286 (I874373,I2507,I873949,I873920,);
nor I_51287 (I874404,I874252,I874308);
not I_51288 (I874421,I874404);
nand I_51289 (I873929,I874421,I874277);
not I_51290 (I874476,I2514);
DFFARX1 I_51291 (I466453,I2507,I874476,I874502,);
not I_51292 (I874510,I874502);
nand I_51293 (I874527,I466450,I466459);
and I_51294 (I874544,I874527,I466468);
DFFARX1 I_51295 (I874544,I2507,I874476,I874570,);
DFFARX1 I_51296 (I874570,I2507,I874476,I874465,);
DFFARX1 I_51297 (I466471,I2507,I874476,I874601,);
nand I_51298 (I874609,I874601,I466474);
not I_51299 (I874626,I874609);
DFFARX1 I_51300 (I874626,I2507,I874476,I874652,);
not I_51301 (I874660,I874652);
nor I_51302 (I874468,I874510,I874660);
DFFARX1 I_51303 (I466447,I2507,I874476,I874700,);
nor I_51304 (I874459,I874700,I874570);
nor I_51305 (I874450,I874700,I874626);
nand I_51306 (I874736,I466462,I466465);
and I_51307 (I874753,I874736,I466456);
DFFARX1 I_51308 (I874753,I2507,I874476,I874779,);
not I_51309 (I874787,I874779);
nand I_51310 (I874804,I874787,I874700);
nand I_51311 (I874453,I874787,I874609);
nor I_51312 (I874835,I466447,I466465);
and I_51313 (I874852,I874700,I874835);
nor I_51314 (I874869,I874787,I874852);
DFFARX1 I_51315 (I874869,I2507,I874476,I874462,);
nor I_51316 (I874900,I874502,I874835);
DFFARX1 I_51317 (I874900,I2507,I874476,I874447,);
nor I_51318 (I874931,I874779,I874835);
not I_51319 (I874948,I874931);
nand I_51320 (I874456,I874948,I874804);
not I_51321 (I875003,I2514);
DFFARX1 I_51322 (I690830,I2507,I875003,I875029,);
not I_51323 (I875037,I875029);
nand I_51324 (I875054,I690833,I690830);
and I_51325 (I875071,I875054,I690842);
DFFARX1 I_51326 (I875071,I2507,I875003,I875097,);
DFFARX1 I_51327 (I875097,I2507,I875003,I874992,);
DFFARX1 I_51328 (I690839,I2507,I875003,I875128,);
nand I_51329 (I875136,I875128,I690845);
not I_51330 (I875153,I875136);
DFFARX1 I_51331 (I875153,I2507,I875003,I875179,);
not I_51332 (I875187,I875179);
nor I_51333 (I874995,I875037,I875187);
DFFARX1 I_51334 (I690854,I2507,I875003,I875227,);
nor I_51335 (I874986,I875227,I875097);
nor I_51336 (I874977,I875227,I875153);
nand I_51337 (I875263,I690848,I690836);
and I_51338 (I875280,I875263,I690833);
DFFARX1 I_51339 (I875280,I2507,I875003,I875306,);
not I_51340 (I875314,I875306);
nand I_51341 (I875331,I875314,I875227);
nand I_51342 (I874980,I875314,I875136);
nor I_51343 (I875362,I690851,I690836);
and I_51344 (I875379,I875227,I875362);
nor I_51345 (I875396,I875314,I875379);
DFFARX1 I_51346 (I875396,I2507,I875003,I874989,);
nor I_51347 (I875427,I875029,I875362);
DFFARX1 I_51348 (I875427,I2507,I875003,I874974,);
nor I_51349 (I875458,I875306,I875362);
not I_51350 (I875475,I875458);
nand I_51351 (I874983,I875475,I875331);
not I_51352 (I875530,I2514);
DFFARX1 I_51353 (I583915,I2507,I875530,I875556,);
not I_51354 (I875564,I875556);
nand I_51355 (I875581,I583900,I583921);
and I_51356 (I875598,I875581,I583909);
DFFARX1 I_51357 (I875598,I2507,I875530,I875624,);
DFFARX1 I_51358 (I875624,I2507,I875530,I875519,);
DFFARX1 I_51359 (I583903,I2507,I875530,I875655,);
nand I_51360 (I875663,I875655,I583912);
not I_51361 (I875680,I875663);
DFFARX1 I_51362 (I875680,I2507,I875530,I875706,);
not I_51363 (I875714,I875706);
nor I_51364 (I875522,I875564,I875714);
DFFARX1 I_51365 (I583918,I2507,I875530,I875754,);
nor I_51366 (I875513,I875754,I875624);
nor I_51367 (I875504,I875754,I875680);
nand I_51368 (I875790,I583900,I583903);
and I_51369 (I875807,I875790,I583924);
DFFARX1 I_51370 (I875807,I2507,I875530,I875833,);
not I_51371 (I875841,I875833);
nand I_51372 (I875858,I875841,I875754);
nand I_51373 (I875507,I875841,I875663);
nor I_51374 (I875889,I583906,I583903);
and I_51375 (I875906,I875754,I875889);
nor I_51376 (I875923,I875841,I875906);
DFFARX1 I_51377 (I875923,I2507,I875530,I875516,);
nor I_51378 (I875954,I875556,I875889);
DFFARX1 I_51379 (I875954,I2507,I875530,I875501,);
nor I_51380 (I875985,I875833,I875889);
not I_51381 (I876002,I875985);
nand I_51382 (I875510,I876002,I875858);
not I_51383 (I876057,I2514);
DFFARX1 I_51384 (I616283,I2507,I876057,I876083,);
not I_51385 (I876091,I876083);
nand I_51386 (I876108,I616268,I616289);
and I_51387 (I876125,I876108,I616277);
DFFARX1 I_51388 (I876125,I2507,I876057,I876151,);
DFFARX1 I_51389 (I876151,I2507,I876057,I876046,);
DFFARX1 I_51390 (I616271,I2507,I876057,I876182,);
nand I_51391 (I876190,I876182,I616280);
not I_51392 (I876207,I876190);
DFFARX1 I_51393 (I876207,I2507,I876057,I876233,);
not I_51394 (I876241,I876233);
nor I_51395 (I876049,I876091,I876241);
DFFARX1 I_51396 (I616286,I2507,I876057,I876281,);
nor I_51397 (I876040,I876281,I876151);
nor I_51398 (I876031,I876281,I876207);
nand I_51399 (I876317,I616268,I616271);
and I_51400 (I876334,I876317,I616292);
DFFARX1 I_51401 (I876334,I2507,I876057,I876360,);
not I_51402 (I876368,I876360);
nand I_51403 (I876385,I876368,I876281);
nand I_51404 (I876034,I876368,I876190);
nor I_51405 (I876416,I616274,I616271);
and I_51406 (I876433,I876281,I876416);
nor I_51407 (I876450,I876368,I876433);
DFFARX1 I_51408 (I876450,I2507,I876057,I876043,);
nor I_51409 (I876481,I876083,I876416);
DFFARX1 I_51410 (I876481,I2507,I876057,I876028,);
nor I_51411 (I876512,I876360,I876416);
not I_51412 (I876529,I876512);
nand I_51413 (I876037,I876529,I876385);
not I_51414 (I876584,I2514);
DFFARX1 I_51415 (I664820,I2507,I876584,I876610,);
not I_51416 (I876618,I876610);
nand I_51417 (I876635,I664823,I664820);
and I_51418 (I876652,I876635,I664832);
DFFARX1 I_51419 (I876652,I2507,I876584,I876678,);
DFFARX1 I_51420 (I876678,I2507,I876584,I876573,);
DFFARX1 I_51421 (I664829,I2507,I876584,I876709,);
nand I_51422 (I876717,I876709,I664835);
not I_51423 (I876734,I876717);
DFFARX1 I_51424 (I876734,I2507,I876584,I876760,);
not I_51425 (I876768,I876760);
nor I_51426 (I876576,I876618,I876768);
DFFARX1 I_51427 (I664844,I2507,I876584,I876808,);
nor I_51428 (I876567,I876808,I876678);
nor I_51429 (I876558,I876808,I876734);
nand I_51430 (I876844,I664838,I664826);
and I_51431 (I876861,I876844,I664823);
DFFARX1 I_51432 (I876861,I2507,I876584,I876887,);
not I_51433 (I876895,I876887);
nand I_51434 (I876912,I876895,I876808);
nand I_51435 (I876561,I876895,I876717);
nor I_51436 (I876943,I664841,I664826);
and I_51437 (I876960,I876808,I876943);
nor I_51438 (I876977,I876895,I876960);
DFFARX1 I_51439 (I876977,I2507,I876584,I876570,);
nor I_51440 (I877008,I876610,I876943);
DFFARX1 I_51441 (I877008,I2507,I876584,I876555,);
nor I_51442 (I877039,I876887,I876943);
not I_51443 (I877056,I877039);
nand I_51444 (I876564,I877056,I876912);
not I_51445 (I877111,I2514);
DFFARX1 I_51446 (I264428,I2507,I877111,I877137,);
not I_51447 (I877145,I877137);
nand I_51448 (I877162,I264419,I264419);
and I_51449 (I877179,I877162,I264437);
DFFARX1 I_51450 (I877179,I2507,I877111,I877205,);
DFFARX1 I_51451 (I877205,I2507,I877111,I877100,);
DFFARX1 I_51452 (I264440,I2507,I877111,I877236,);
nand I_51453 (I877244,I877236,I264422);
not I_51454 (I877261,I877244);
DFFARX1 I_51455 (I877261,I2507,I877111,I877287,);
not I_51456 (I877295,I877287);
nor I_51457 (I877103,I877145,I877295);
DFFARX1 I_51458 (I264434,I2507,I877111,I877335,);
nor I_51459 (I877094,I877335,I877205);
nor I_51460 (I877085,I877335,I877261);
nand I_51461 (I877371,I264446,I264425);
and I_51462 (I877388,I877371,I264431);
DFFARX1 I_51463 (I877388,I2507,I877111,I877414,);
not I_51464 (I877422,I877414);
nand I_51465 (I877439,I877422,I877335);
nand I_51466 (I877088,I877422,I877244);
nor I_51467 (I877470,I264443,I264425);
and I_51468 (I877487,I877335,I877470);
nor I_51469 (I877504,I877422,I877487);
DFFARX1 I_51470 (I877504,I2507,I877111,I877097,);
nor I_51471 (I877535,I877137,I877470);
DFFARX1 I_51472 (I877535,I2507,I877111,I877082,);
nor I_51473 (I877566,I877414,I877470);
not I_51474 (I877583,I877566);
nand I_51475 (I877091,I877583,I877439);
not I_51476 (I877638,I2514);
DFFARX1 I_51477 (I142519,I2507,I877638,I877664,);
not I_51478 (I877672,I877664);
nand I_51479 (I877689,I142495,I142513);
and I_51480 (I877706,I877689,I142501);
DFFARX1 I_51481 (I877706,I2507,I877638,I877732,);
DFFARX1 I_51482 (I877732,I2507,I877638,I877627,);
DFFARX1 I_51483 (I142510,I2507,I877638,I877763,);
nand I_51484 (I877771,I877763,I142516);
not I_51485 (I877788,I877771);
DFFARX1 I_51486 (I877788,I2507,I877638,I877814,);
not I_51487 (I877822,I877814);
nor I_51488 (I877630,I877672,I877822);
DFFARX1 I_51489 (I142495,I2507,I877638,I877862,);
nor I_51490 (I877621,I877862,I877732);
nor I_51491 (I877612,I877862,I877788);
nand I_51492 (I877898,I142507,I142498);
and I_51493 (I877915,I877898,I142522);
DFFARX1 I_51494 (I877915,I2507,I877638,I877941,);
not I_51495 (I877949,I877941);
nand I_51496 (I877966,I877949,I877862);
nand I_51497 (I877615,I877949,I877771);
nor I_51498 (I877997,I142504,I142498);
and I_51499 (I878014,I877862,I877997);
nor I_51500 (I878031,I877949,I878014);
DFFARX1 I_51501 (I878031,I2507,I877638,I877624,);
nor I_51502 (I878062,I877664,I877997);
DFFARX1 I_51503 (I878062,I2507,I877638,I877609,);
nor I_51504 (I878093,I877941,I877997);
not I_51505 (I878110,I878093);
nand I_51506 (I877618,I878110,I877966);
not I_51507 (I878165,I2514);
DFFARX1 I_51508 (I1128326,I2507,I878165,I878191,);
not I_51509 (I878199,I878191);
nand I_51510 (I878216,I1128308,I1128308);
and I_51511 (I878233,I878216,I1128314);
DFFARX1 I_51512 (I878233,I2507,I878165,I878259,);
DFFARX1 I_51513 (I878259,I2507,I878165,I878154,);
DFFARX1 I_51514 (I1128311,I2507,I878165,I878290,);
nand I_51515 (I878298,I878290,I1128320);
not I_51516 (I878315,I878298);
DFFARX1 I_51517 (I878315,I2507,I878165,I878341,);
not I_51518 (I878349,I878341);
nor I_51519 (I878157,I878199,I878349);
DFFARX1 I_51520 (I1128332,I2507,I878165,I878389,);
nor I_51521 (I878148,I878389,I878259);
nor I_51522 (I878139,I878389,I878315);
nand I_51523 (I878425,I1128323,I1128317);
and I_51524 (I878442,I878425,I1128311);
DFFARX1 I_51525 (I878442,I2507,I878165,I878468,);
not I_51526 (I878476,I878468);
nand I_51527 (I878493,I878476,I878389);
nand I_51528 (I878142,I878476,I878298);
nor I_51529 (I878524,I1128329,I1128317);
and I_51530 (I878541,I878389,I878524);
nor I_51531 (I878558,I878476,I878541);
DFFARX1 I_51532 (I878558,I2507,I878165,I878151,);
nor I_51533 (I878589,I878191,I878524);
DFFARX1 I_51534 (I878589,I2507,I878165,I878136,);
nor I_51535 (I878620,I878468,I878524);
not I_51536 (I878637,I878620);
nand I_51537 (I878145,I878637,I878493);
not I_51538 (I878692,I2514);
DFFARX1 I_51539 (I1093646,I2507,I878692,I878718,);
not I_51540 (I878726,I878718);
nand I_51541 (I878743,I1093628,I1093628);
and I_51542 (I878760,I878743,I1093634);
DFFARX1 I_51543 (I878760,I2507,I878692,I878786,);
DFFARX1 I_51544 (I878786,I2507,I878692,I878681,);
DFFARX1 I_51545 (I1093631,I2507,I878692,I878817,);
nand I_51546 (I878825,I878817,I1093640);
not I_51547 (I878842,I878825);
DFFARX1 I_51548 (I878842,I2507,I878692,I878868,);
not I_51549 (I878876,I878868);
nor I_51550 (I878684,I878726,I878876);
DFFARX1 I_51551 (I1093652,I2507,I878692,I878916,);
nor I_51552 (I878675,I878916,I878786);
nor I_51553 (I878666,I878916,I878842);
nand I_51554 (I878952,I1093643,I1093637);
and I_51555 (I878969,I878952,I1093631);
DFFARX1 I_51556 (I878969,I2507,I878692,I878995,);
not I_51557 (I879003,I878995);
nand I_51558 (I879020,I879003,I878916);
nand I_51559 (I878669,I879003,I878825);
nor I_51560 (I879051,I1093649,I1093637);
and I_51561 (I879068,I878916,I879051);
nor I_51562 (I879085,I879003,I879068);
DFFARX1 I_51563 (I879085,I2507,I878692,I878678,);
nor I_51564 (I879116,I878718,I879051);
DFFARX1 I_51565 (I879116,I2507,I878692,I878663,);
nor I_51566 (I879147,I878995,I879051);
not I_51567 (I879164,I879147);
nand I_51568 (I878672,I879164,I879020);
not I_51569 (I879219,I2514);
DFFARX1 I_51570 (I533365,I2507,I879219,I879245,);
not I_51571 (I879253,I879245);
nand I_51572 (I879270,I533383,I533374);
and I_51573 (I879287,I879270,I533377);
DFFARX1 I_51574 (I879287,I2507,I879219,I879313,);
DFFARX1 I_51575 (I879313,I2507,I879219,I879208,);
DFFARX1 I_51576 (I533371,I2507,I879219,I879344,);
nand I_51577 (I879352,I879344,I533362);
not I_51578 (I879369,I879352);
DFFARX1 I_51579 (I879369,I2507,I879219,I879395,);
not I_51580 (I879403,I879395);
nor I_51581 (I879211,I879253,I879403);
DFFARX1 I_51582 (I533368,I2507,I879219,I879443,);
nor I_51583 (I879202,I879443,I879313);
nor I_51584 (I879193,I879443,I879369);
nand I_51585 (I879479,I533362,I533359);
and I_51586 (I879496,I879479,I533380);
DFFARX1 I_51587 (I879496,I2507,I879219,I879522,);
not I_51588 (I879530,I879522);
nand I_51589 (I879547,I879530,I879443);
nand I_51590 (I879196,I879530,I879352);
nor I_51591 (I879578,I533359,I533359);
and I_51592 (I879595,I879443,I879578);
nor I_51593 (I879612,I879530,I879595);
DFFARX1 I_51594 (I879612,I2507,I879219,I879205,);
nor I_51595 (I879643,I879245,I879578);
DFFARX1 I_51596 (I879643,I2507,I879219,I879190,);
nor I_51597 (I879674,I879522,I879578);
not I_51598 (I879691,I879674);
nand I_51599 (I879199,I879691,I879547);
not I_51600 (I879746,I2514);
DFFARX1 I_51601 (I426741,I2507,I879746,I879772,);
not I_51602 (I879780,I879772);
nand I_51603 (I879797,I426738,I426747);
and I_51604 (I879814,I879797,I426756);
DFFARX1 I_51605 (I879814,I2507,I879746,I879840,);
DFFARX1 I_51606 (I879840,I2507,I879746,I879735,);
DFFARX1 I_51607 (I426759,I2507,I879746,I879871,);
nand I_51608 (I879879,I879871,I426762);
not I_51609 (I879896,I879879);
DFFARX1 I_51610 (I879896,I2507,I879746,I879922,);
not I_51611 (I879930,I879922);
nor I_51612 (I879738,I879780,I879930);
DFFARX1 I_51613 (I426735,I2507,I879746,I879970,);
nor I_51614 (I879729,I879970,I879840);
nor I_51615 (I879720,I879970,I879896);
nand I_51616 (I880006,I426750,I426753);
and I_51617 (I880023,I880006,I426744);
DFFARX1 I_51618 (I880023,I2507,I879746,I880049,);
not I_51619 (I880057,I880049);
nand I_51620 (I880074,I880057,I879970);
nand I_51621 (I879723,I880057,I879879);
nor I_51622 (I880105,I426735,I426753);
and I_51623 (I880122,I879970,I880105);
nor I_51624 (I880139,I880057,I880122);
DFFARX1 I_51625 (I880139,I2507,I879746,I879732,);
nor I_51626 (I880170,I879772,I880105);
DFFARX1 I_51627 (I880170,I2507,I879746,I879717,);
nor I_51628 (I880201,I880049,I880105);
not I_51629 (I880218,I880201);
nand I_51630 (I879726,I880218,I880074);
not I_51631 (I880273,I2514);
DFFARX1 I_51632 (I1121390,I2507,I880273,I880299,);
not I_51633 (I880307,I880299);
nand I_51634 (I880324,I1121372,I1121372);
and I_51635 (I880341,I880324,I1121378);
DFFARX1 I_51636 (I880341,I2507,I880273,I880367,);
DFFARX1 I_51637 (I880367,I2507,I880273,I880262,);
DFFARX1 I_51638 (I1121375,I2507,I880273,I880398,);
nand I_51639 (I880406,I880398,I1121384);
not I_51640 (I880423,I880406);
DFFARX1 I_51641 (I880423,I2507,I880273,I880449,);
not I_51642 (I880457,I880449);
nor I_51643 (I880265,I880307,I880457);
DFFARX1 I_51644 (I1121396,I2507,I880273,I880497,);
nor I_51645 (I880256,I880497,I880367);
nor I_51646 (I880247,I880497,I880423);
nand I_51647 (I880533,I1121387,I1121381);
and I_51648 (I880550,I880533,I1121375);
DFFARX1 I_51649 (I880550,I2507,I880273,I880576,);
not I_51650 (I880584,I880576);
nand I_51651 (I880601,I880584,I880497);
nand I_51652 (I880250,I880584,I880406);
nor I_51653 (I880632,I1121393,I1121381);
and I_51654 (I880649,I880497,I880632);
nor I_51655 (I880666,I880584,I880649);
DFFARX1 I_51656 (I880666,I2507,I880273,I880259,);
nor I_51657 (I880697,I880299,I880632);
DFFARX1 I_51658 (I880697,I2507,I880273,I880244,);
nor I_51659 (I880728,I880576,I880632);
not I_51660 (I880745,I880728);
nand I_51661 (I880253,I880745,I880601);
not I_51662 (I880800,I2514);
DFFARX1 I_51663 (I1285984,I2507,I880800,I880826,);
not I_51664 (I880834,I880826);
nand I_51665 (I880851,I1285966,I1285969);
and I_51666 (I880868,I880851,I1285981);
DFFARX1 I_51667 (I880868,I2507,I880800,I880894,);
DFFARX1 I_51668 (I880894,I2507,I880800,I880789,);
DFFARX1 I_51669 (I1285990,I2507,I880800,I880925,);
nand I_51670 (I880933,I880925,I1285975);
not I_51671 (I880950,I880933);
DFFARX1 I_51672 (I880950,I2507,I880800,I880976,);
not I_51673 (I880984,I880976);
nor I_51674 (I880792,I880834,I880984);
DFFARX1 I_51675 (I1285987,I2507,I880800,I881024,);
nor I_51676 (I880783,I881024,I880894);
nor I_51677 (I880774,I881024,I880950);
nand I_51678 (I881060,I1285978,I1285972);
and I_51679 (I881077,I881060,I1285966);
DFFARX1 I_51680 (I881077,I2507,I880800,I881103,);
not I_51681 (I881111,I881103);
nand I_51682 (I881128,I881111,I881024);
nand I_51683 (I880777,I881111,I880933);
nor I_51684 (I881159,I1285969,I1285972);
and I_51685 (I881176,I881024,I881159);
nor I_51686 (I881193,I881111,I881176);
DFFARX1 I_51687 (I881193,I2507,I880800,I880786,);
nor I_51688 (I881224,I880826,I881159);
DFFARX1 I_51689 (I881224,I2507,I880800,I880771,);
nor I_51690 (I881255,I881103,I881159);
not I_51691 (I881272,I881255);
nand I_51692 (I880780,I881272,I881128);
not I_51693 (I881327,I2514);
DFFARX1 I_51694 (I746318,I2507,I881327,I881353,);
not I_51695 (I881361,I881353);
nand I_51696 (I881378,I746321,I746318);
and I_51697 (I881395,I881378,I746330);
DFFARX1 I_51698 (I881395,I2507,I881327,I881421,);
DFFARX1 I_51699 (I881421,I2507,I881327,I881316,);
DFFARX1 I_51700 (I746327,I2507,I881327,I881452,);
nand I_51701 (I881460,I881452,I746333);
not I_51702 (I881477,I881460);
DFFARX1 I_51703 (I881477,I2507,I881327,I881503,);
not I_51704 (I881511,I881503);
nor I_51705 (I881319,I881361,I881511);
DFFARX1 I_51706 (I746342,I2507,I881327,I881551,);
nor I_51707 (I881310,I881551,I881421);
nor I_51708 (I881301,I881551,I881477);
nand I_51709 (I881587,I746336,I746324);
and I_51710 (I881604,I881587,I746321);
DFFARX1 I_51711 (I881604,I2507,I881327,I881630,);
not I_51712 (I881638,I881630);
nand I_51713 (I881655,I881638,I881551);
nand I_51714 (I881304,I881638,I881460);
nor I_51715 (I881686,I746339,I746324);
and I_51716 (I881703,I881551,I881686);
nor I_51717 (I881720,I881638,I881703);
DFFARX1 I_51718 (I881720,I2507,I881327,I881313,);
nor I_51719 (I881751,I881353,I881686);
DFFARX1 I_51720 (I881751,I2507,I881327,I881298,);
nor I_51721 (I881782,I881630,I881686);
not I_51722 (I881799,I881782);
nand I_51723 (I881307,I881799,I881655);
not I_51724 (I881854,I2514);
DFFARX1 I_51725 (I483861,I2507,I881854,I881880,);
not I_51726 (I881888,I881880);
nand I_51727 (I881905,I483858,I483867);
and I_51728 (I881922,I881905,I483876);
DFFARX1 I_51729 (I881922,I2507,I881854,I881948,);
DFFARX1 I_51730 (I881948,I2507,I881854,I881843,);
DFFARX1 I_51731 (I483879,I2507,I881854,I881979,);
nand I_51732 (I881987,I881979,I483882);
not I_51733 (I882004,I881987);
DFFARX1 I_51734 (I882004,I2507,I881854,I882030,);
not I_51735 (I882038,I882030);
nor I_51736 (I881846,I881888,I882038);
DFFARX1 I_51737 (I483855,I2507,I881854,I882078,);
nor I_51738 (I881837,I882078,I881948);
nor I_51739 (I881828,I882078,I882004);
nand I_51740 (I882114,I483870,I483873);
and I_51741 (I882131,I882114,I483864);
DFFARX1 I_51742 (I882131,I2507,I881854,I882157,);
not I_51743 (I882165,I882157);
nand I_51744 (I882182,I882165,I882078);
nand I_51745 (I881831,I882165,I881987);
nor I_51746 (I882213,I483855,I483873);
and I_51747 (I882230,I882078,I882213);
nor I_51748 (I882247,I882165,I882230);
DFFARX1 I_51749 (I882247,I2507,I881854,I881840,);
nor I_51750 (I882278,I881880,I882213);
DFFARX1 I_51751 (I882278,I2507,I881854,I881825,);
nor I_51752 (I882309,I882157,I882213);
not I_51753 (I882326,I882309);
nand I_51754 (I881834,I882326,I882182);
not I_51755 (I882381,I2514);
DFFARX1 I_51756 (I1072260,I2507,I882381,I882407,);
not I_51757 (I882415,I882407);
nand I_51758 (I882432,I1072242,I1072242);
and I_51759 (I882449,I882432,I1072248);
DFFARX1 I_51760 (I882449,I2507,I882381,I882475,);
DFFARX1 I_51761 (I882475,I2507,I882381,I882370,);
DFFARX1 I_51762 (I1072245,I2507,I882381,I882506,);
nand I_51763 (I882514,I882506,I1072254);
not I_51764 (I882531,I882514);
DFFARX1 I_51765 (I882531,I2507,I882381,I882557,);
not I_51766 (I882565,I882557);
nor I_51767 (I882373,I882415,I882565);
DFFARX1 I_51768 (I1072266,I2507,I882381,I882605,);
nor I_51769 (I882364,I882605,I882475);
nor I_51770 (I882355,I882605,I882531);
nand I_51771 (I882641,I1072257,I1072251);
and I_51772 (I882658,I882641,I1072245);
DFFARX1 I_51773 (I882658,I2507,I882381,I882684,);
not I_51774 (I882692,I882684);
nand I_51775 (I882709,I882692,I882605);
nand I_51776 (I882358,I882692,I882514);
nor I_51777 (I882740,I1072263,I1072251);
and I_51778 (I882757,I882605,I882740);
nor I_51779 (I882774,I882692,I882757);
DFFARX1 I_51780 (I882774,I2507,I882381,I882367,);
nor I_51781 (I882805,I882407,I882740);
DFFARX1 I_51782 (I882805,I2507,I882381,I882352,);
nor I_51783 (I882836,I882684,I882740);
not I_51784 (I882853,I882836);
nand I_51785 (I882361,I882853,I882709);
not I_51786 (I882908,I2514);
DFFARX1 I_51787 (I1277314,I2507,I882908,I882934,);
not I_51788 (I882942,I882934);
nand I_51789 (I882959,I1277296,I1277299);
and I_51790 (I882976,I882959,I1277311);
DFFARX1 I_51791 (I882976,I2507,I882908,I883002,);
DFFARX1 I_51792 (I883002,I2507,I882908,I882897,);
DFFARX1 I_51793 (I1277320,I2507,I882908,I883033,);
nand I_51794 (I883041,I883033,I1277305);
not I_51795 (I883058,I883041);
DFFARX1 I_51796 (I883058,I2507,I882908,I883084,);
not I_51797 (I883092,I883084);
nor I_51798 (I882900,I882942,I883092);
DFFARX1 I_51799 (I1277317,I2507,I882908,I883132,);
nor I_51800 (I882891,I883132,I883002);
nor I_51801 (I882882,I883132,I883058);
nand I_51802 (I883168,I1277308,I1277302);
and I_51803 (I883185,I883168,I1277296);
DFFARX1 I_51804 (I883185,I2507,I882908,I883211,);
not I_51805 (I883219,I883211);
nand I_51806 (I883236,I883219,I883132);
nand I_51807 (I882885,I883219,I883041);
nor I_51808 (I883267,I1277299,I1277302);
and I_51809 (I883284,I883132,I883267);
nor I_51810 (I883301,I883219,I883284);
DFFARX1 I_51811 (I883301,I2507,I882908,I882894,);
nor I_51812 (I883332,I882934,I883267);
DFFARX1 I_51813 (I883332,I2507,I882908,I882879,);
nor I_51814 (I883363,I883211,I883267);
not I_51815 (I883380,I883363);
nand I_51816 (I882888,I883380,I883236);
not I_51817 (I883435,I2514);
DFFARX1 I_51818 (I1331507,I2507,I883435,I883461,);
not I_51819 (I883469,I883461);
nand I_51820 (I883486,I1331504,I1331513);
and I_51821 (I883503,I883486,I1331492);
DFFARX1 I_51822 (I883503,I2507,I883435,I883529,);
DFFARX1 I_51823 (I883529,I2507,I883435,I883424,);
DFFARX1 I_51824 (I1331495,I2507,I883435,I883560,);
nand I_51825 (I883568,I883560,I1331510);
not I_51826 (I883585,I883568);
DFFARX1 I_51827 (I883585,I2507,I883435,I883611,);
not I_51828 (I883619,I883611);
nor I_51829 (I883427,I883469,I883619);
DFFARX1 I_51830 (I1331516,I2507,I883435,I883659,);
nor I_51831 (I883418,I883659,I883529);
nor I_51832 (I883409,I883659,I883585);
nand I_51833 (I883695,I1331498,I1331519);
and I_51834 (I883712,I883695,I1331501);
DFFARX1 I_51835 (I883712,I2507,I883435,I883738,);
not I_51836 (I883746,I883738);
nand I_51837 (I883763,I883746,I883659);
nand I_51838 (I883412,I883746,I883568);
nor I_51839 (I883794,I1331492,I1331519);
and I_51840 (I883811,I883659,I883794);
nor I_51841 (I883828,I883746,I883811);
DFFARX1 I_51842 (I883828,I2507,I883435,I883421,);
nor I_51843 (I883859,I883461,I883794);
DFFARX1 I_51844 (I883859,I2507,I883435,I883406,);
nor I_51845 (I883890,I883738,I883794);
not I_51846 (I883907,I883890);
nand I_51847 (I883415,I883907,I883763);
not I_51848 (I883962,I2514);
DFFARX1 I_51849 (I404981,I2507,I883962,I883988,);
not I_51850 (I883996,I883988);
nand I_51851 (I884013,I404978,I404987);
and I_51852 (I884030,I884013,I404996);
DFFARX1 I_51853 (I884030,I2507,I883962,I884056,);
DFFARX1 I_51854 (I884056,I2507,I883962,I883951,);
DFFARX1 I_51855 (I404999,I2507,I883962,I884087,);
nand I_51856 (I884095,I884087,I405002);
not I_51857 (I884112,I884095);
DFFARX1 I_51858 (I884112,I2507,I883962,I884138,);
not I_51859 (I884146,I884138);
nor I_51860 (I883954,I883996,I884146);
DFFARX1 I_51861 (I404975,I2507,I883962,I884186,);
nor I_51862 (I883945,I884186,I884056);
nor I_51863 (I883936,I884186,I884112);
nand I_51864 (I884222,I404990,I404993);
and I_51865 (I884239,I884222,I404984);
DFFARX1 I_51866 (I884239,I2507,I883962,I884265,);
not I_51867 (I884273,I884265);
nand I_51868 (I884290,I884273,I884186);
nand I_51869 (I883939,I884273,I884095);
nor I_51870 (I884321,I404975,I404993);
and I_51871 (I884338,I884186,I884321);
nor I_51872 (I884355,I884273,I884338);
DFFARX1 I_51873 (I884355,I2507,I883962,I883948,);
nor I_51874 (I884386,I883988,I884321);
DFFARX1 I_51875 (I884386,I2507,I883962,I883933,);
nor I_51876 (I884417,I884265,I884321);
not I_51877 (I884434,I884417);
nand I_51878 (I883942,I884434,I884290);
not I_51879 (I884489,I2514);
DFFARX1 I_51880 (I445237,I2507,I884489,I884515,);
not I_51881 (I884523,I884515);
nand I_51882 (I884540,I445234,I445243);
and I_51883 (I884557,I884540,I445252);
DFFARX1 I_51884 (I884557,I2507,I884489,I884583,);
DFFARX1 I_51885 (I884583,I2507,I884489,I884478,);
DFFARX1 I_51886 (I445255,I2507,I884489,I884614,);
nand I_51887 (I884622,I884614,I445258);
not I_51888 (I884639,I884622);
DFFARX1 I_51889 (I884639,I2507,I884489,I884665,);
not I_51890 (I884673,I884665);
nor I_51891 (I884481,I884523,I884673);
DFFARX1 I_51892 (I445231,I2507,I884489,I884713,);
nor I_51893 (I884472,I884713,I884583);
nor I_51894 (I884463,I884713,I884639);
nand I_51895 (I884749,I445246,I445249);
and I_51896 (I884766,I884749,I445240);
DFFARX1 I_51897 (I884766,I2507,I884489,I884792,);
not I_51898 (I884800,I884792);
nand I_51899 (I884817,I884800,I884713);
nand I_51900 (I884466,I884800,I884622);
nor I_51901 (I884848,I445231,I445249);
and I_51902 (I884865,I884713,I884848);
nor I_51903 (I884882,I884800,I884865);
DFFARX1 I_51904 (I884882,I2507,I884489,I884475,);
nor I_51905 (I884913,I884515,I884848);
DFFARX1 I_51906 (I884913,I2507,I884489,I884460,);
nor I_51907 (I884944,I884792,I884848);
not I_51908 (I884961,I884944);
nand I_51909 (I884469,I884961,I884817);
not I_51910 (I885022,I2514);
DFFARX1 I_51911 (I328186,I2507,I885022,I885048,);
DFFARX1 I_51912 (I328192,I2507,I885022,I885065,);
not I_51913 (I885073,I885065);
not I_51914 (I885090,I328213);
nor I_51915 (I885107,I885090,I328201);
not I_51916 (I885124,I328210);
nor I_51917 (I885141,I885107,I328195);
nor I_51918 (I885158,I885065,I885141);
DFFARX1 I_51919 (I885158,I2507,I885022,I885008,);
nor I_51920 (I885189,I328195,I328201);
nand I_51921 (I885206,I885189,I328213);
DFFARX1 I_51922 (I885206,I2507,I885022,I885011,);
nor I_51923 (I885237,I885124,I328195);
nand I_51924 (I885254,I885237,I328186);
nor I_51925 (I885271,I885048,I885254);
DFFARX1 I_51926 (I885271,I2507,I885022,I884987,);
not I_51927 (I885302,I885254);
nand I_51928 (I884999,I885065,I885302);
DFFARX1 I_51929 (I885254,I2507,I885022,I885342,);
not I_51930 (I885350,I885342);
not I_51931 (I885367,I328195);
not I_51932 (I885384,I328198);
nor I_51933 (I885401,I885384,I328210);
nor I_51934 (I885014,I885350,I885401);
nor I_51935 (I885432,I885384,I328207);
and I_51936 (I885449,I885432,I328189);
or I_51937 (I885466,I885449,I328204);
DFFARX1 I_51938 (I885466,I2507,I885022,I885492,);
nor I_51939 (I885002,I885492,I885048);
not I_51940 (I885514,I885492);
and I_51941 (I885531,I885514,I885048);
nor I_51942 (I884996,I885073,I885531);
nand I_51943 (I885562,I885514,I885124);
nor I_51944 (I884990,I885384,I885562);
nand I_51945 (I884993,I885514,I885302);
nand I_51946 (I885607,I885124,I328198);
nor I_51947 (I885005,I885367,I885607);
not I_51948 (I885668,I2514);
DFFARX1 I_51949 (I556159,I2507,I885668,I885694,);
DFFARX1 I_51950 (I556171,I2507,I885668,I885711,);
not I_51951 (I885719,I885711);
not I_51952 (I885736,I556180);
nor I_51953 (I885753,I885736,I556156);
not I_51954 (I885770,I556174);
nor I_51955 (I885787,I885753,I556168);
nor I_51956 (I885804,I885711,I885787);
DFFARX1 I_51957 (I885804,I2507,I885668,I885654,);
nor I_51958 (I885835,I556168,I556156);
nand I_51959 (I885852,I885835,I556180);
DFFARX1 I_51960 (I885852,I2507,I885668,I885657,);
nor I_51961 (I885883,I885770,I556168);
nand I_51962 (I885900,I885883,I556162);
nor I_51963 (I885917,I885694,I885900);
DFFARX1 I_51964 (I885917,I2507,I885668,I885633,);
not I_51965 (I885948,I885900);
nand I_51966 (I885645,I885711,I885948);
DFFARX1 I_51967 (I885900,I2507,I885668,I885988,);
not I_51968 (I885996,I885988);
not I_51969 (I886013,I556168);
not I_51970 (I886030,I556177);
nor I_51971 (I886047,I886030,I556174);
nor I_51972 (I885660,I885996,I886047);
nor I_51973 (I886078,I886030,I556159);
and I_51974 (I886095,I886078,I556156);
or I_51975 (I886112,I886095,I556165);
DFFARX1 I_51976 (I886112,I2507,I885668,I886138,);
nor I_51977 (I885648,I886138,I885694);
not I_51978 (I886160,I886138);
and I_51979 (I886177,I886160,I885694);
nor I_51980 (I885642,I885719,I886177);
nand I_51981 (I886208,I886160,I885770);
nor I_51982 (I885636,I886030,I886208);
nand I_51983 (I885639,I886160,I885948);
nand I_51984 (I886253,I885770,I556177);
nor I_51985 (I885651,I886013,I886253);
not I_51986 (I886314,I2514);
DFFARX1 I_51987 (I365076,I2507,I886314,I886340,);
DFFARX1 I_51988 (I365082,I2507,I886314,I886357,);
not I_51989 (I886365,I886357);
not I_51990 (I886382,I365103);
nor I_51991 (I886399,I886382,I365091);
not I_51992 (I886416,I365100);
nor I_51993 (I886433,I886399,I365085);
nor I_51994 (I886450,I886357,I886433);
DFFARX1 I_51995 (I886450,I2507,I886314,I886300,);
nor I_51996 (I886481,I365085,I365091);
nand I_51997 (I886498,I886481,I365103);
DFFARX1 I_51998 (I886498,I2507,I886314,I886303,);
nor I_51999 (I886529,I886416,I365085);
nand I_52000 (I886546,I886529,I365076);
nor I_52001 (I886563,I886340,I886546);
DFFARX1 I_52002 (I886563,I2507,I886314,I886279,);
not I_52003 (I886594,I886546);
nand I_52004 (I886291,I886357,I886594);
DFFARX1 I_52005 (I886546,I2507,I886314,I886634,);
not I_52006 (I886642,I886634);
not I_52007 (I886659,I365085);
not I_52008 (I886676,I365088);
nor I_52009 (I886693,I886676,I365100);
nor I_52010 (I886306,I886642,I886693);
nor I_52011 (I886724,I886676,I365097);
and I_52012 (I886741,I886724,I365079);
or I_52013 (I886758,I886741,I365094);
DFFARX1 I_52014 (I886758,I2507,I886314,I886784,);
nor I_52015 (I886294,I886784,I886340);
not I_52016 (I886806,I886784);
and I_52017 (I886823,I886806,I886340);
nor I_52018 (I886288,I886365,I886823);
nand I_52019 (I886854,I886806,I886416);
nor I_52020 (I886282,I886676,I886854);
nand I_52021 (I886285,I886806,I886594);
nand I_52022 (I886899,I886416,I365088);
nor I_52023 (I886297,I886659,I886899);
not I_52024 (I886960,I2514);
DFFARX1 I_52025 (I780120,I2507,I886960,I886986,);
DFFARX1 I_52026 (I780117,I2507,I886960,I887003,);
not I_52027 (I887011,I887003);
not I_52028 (I887028,I780117);
nor I_52029 (I887045,I887028,I780120);
not I_52030 (I887062,I780132);
nor I_52031 (I887079,I887045,I780126);
nor I_52032 (I887096,I887003,I887079);
DFFARX1 I_52033 (I887096,I2507,I886960,I886946,);
nor I_52034 (I887127,I780126,I780120);
nand I_52035 (I887144,I887127,I780117);
DFFARX1 I_52036 (I887144,I2507,I886960,I886949,);
nor I_52037 (I887175,I887062,I780126);
nand I_52038 (I887192,I887175,I780114);
nor I_52039 (I887209,I886986,I887192);
DFFARX1 I_52040 (I887209,I2507,I886960,I886925,);
not I_52041 (I887240,I887192);
nand I_52042 (I886937,I887003,I887240);
DFFARX1 I_52043 (I887192,I2507,I886960,I887280,);
not I_52044 (I887288,I887280);
not I_52045 (I887305,I780126);
not I_52046 (I887322,I780123);
nor I_52047 (I887339,I887322,I780132);
nor I_52048 (I886952,I887288,I887339);
nor I_52049 (I887370,I887322,I780129);
and I_52050 (I887387,I887370,I780135);
or I_52051 (I887404,I887387,I780114);
DFFARX1 I_52052 (I887404,I2507,I886960,I887430,);
nor I_52053 (I886940,I887430,I886986);
not I_52054 (I887452,I887430);
and I_52055 (I887469,I887452,I886986);
nor I_52056 (I886934,I887011,I887469);
nand I_52057 (I887500,I887452,I887062);
nor I_52058 (I886928,I887322,I887500);
nand I_52059 (I886931,I887452,I887240);
nand I_52060 (I887545,I887062,I780123);
nor I_52061 (I886943,I887305,I887545);
not I_52062 (I887606,I2514);
DFFARX1 I_52063 (I1357672,I2507,I887606,I887632,);
DFFARX1 I_52064 (I1357696,I2507,I887606,I887649,);
not I_52065 (I887657,I887649);
not I_52066 (I887674,I1357678);
nor I_52067 (I887691,I887674,I1357687);
not I_52068 (I887708,I1357672);
nor I_52069 (I887725,I887691,I1357693);
nor I_52070 (I887742,I887649,I887725);
DFFARX1 I_52071 (I887742,I2507,I887606,I887592,);
nor I_52072 (I887773,I1357693,I1357687);
nand I_52073 (I887790,I887773,I1357678);
DFFARX1 I_52074 (I887790,I2507,I887606,I887595,);
nor I_52075 (I887821,I887708,I1357693);
nand I_52076 (I887838,I887821,I1357690);
nor I_52077 (I887855,I887632,I887838);
DFFARX1 I_52078 (I887855,I2507,I887606,I887571,);
not I_52079 (I887886,I887838);
nand I_52080 (I887583,I887649,I887886);
DFFARX1 I_52081 (I887838,I2507,I887606,I887926,);
not I_52082 (I887934,I887926);
not I_52083 (I887951,I1357693);
not I_52084 (I887968,I1357684);
nor I_52085 (I887985,I887968,I1357672);
nor I_52086 (I887598,I887934,I887985);
nor I_52087 (I888016,I887968,I1357675);
and I_52088 (I888033,I888016,I1357699);
or I_52089 (I888050,I888033,I1357681);
DFFARX1 I_52090 (I888050,I2507,I887606,I888076,);
nor I_52091 (I887586,I888076,I887632);
not I_52092 (I888098,I888076);
and I_52093 (I888115,I888098,I887632);
nor I_52094 (I887580,I887657,I888115);
nand I_52095 (I888146,I888098,I887708);
nor I_52096 (I887574,I887968,I888146);
nand I_52097 (I887577,I888098,I887886);
nand I_52098 (I888191,I887708,I1357684);
nor I_52099 (I887589,I887951,I888191);
not I_52100 (I888252,I2514);
DFFARX1 I_52101 (I612225,I2507,I888252,I888278,);
DFFARX1 I_52102 (I612237,I2507,I888252,I888295,);
not I_52103 (I888303,I888295);
not I_52104 (I888320,I612246);
nor I_52105 (I888337,I888320,I612222);
not I_52106 (I888354,I612240);
nor I_52107 (I888371,I888337,I612234);
nor I_52108 (I888388,I888295,I888371);
DFFARX1 I_52109 (I888388,I2507,I888252,I888238,);
nor I_52110 (I888419,I612234,I612222);
nand I_52111 (I888436,I888419,I612246);
DFFARX1 I_52112 (I888436,I2507,I888252,I888241,);
nor I_52113 (I888467,I888354,I612234);
nand I_52114 (I888484,I888467,I612228);
nor I_52115 (I888501,I888278,I888484);
DFFARX1 I_52116 (I888501,I2507,I888252,I888217,);
not I_52117 (I888532,I888484);
nand I_52118 (I888229,I888295,I888532);
DFFARX1 I_52119 (I888484,I2507,I888252,I888572,);
not I_52120 (I888580,I888572);
not I_52121 (I888597,I612234);
not I_52122 (I888614,I612243);
nor I_52123 (I888631,I888614,I612240);
nor I_52124 (I888244,I888580,I888631);
nor I_52125 (I888662,I888614,I612225);
and I_52126 (I888679,I888662,I612222);
or I_52127 (I888696,I888679,I612231);
DFFARX1 I_52128 (I888696,I2507,I888252,I888722,);
nor I_52129 (I888232,I888722,I888278);
not I_52130 (I888744,I888722);
and I_52131 (I888761,I888744,I888278);
nor I_52132 (I888226,I888303,I888761);
nand I_52133 (I888792,I888744,I888354);
nor I_52134 (I888220,I888614,I888792);
nand I_52135 (I888223,I888744,I888532);
nand I_52136 (I888837,I888354,I612243);
nor I_52137 (I888235,I888597,I888837);
not I_52138 (I888898,I2514);
DFFARX1 I_52139 (I91750,I2507,I888898,I888924,);
DFFARX1 I_52140 (I91756,I2507,I888898,I888941,);
not I_52141 (I888949,I888941);
not I_52142 (I888966,I91774);
nor I_52143 (I888983,I888966,I91753);
not I_52144 (I889000,I91759);
nor I_52145 (I889017,I888983,I91765);
nor I_52146 (I889034,I888941,I889017);
DFFARX1 I_52147 (I889034,I2507,I888898,I888884,);
nor I_52148 (I889065,I91765,I91753);
nand I_52149 (I889082,I889065,I91774);
DFFARX1 I_52150 (I889082,I2507,I888898,I888887,);
nor I_52151 (I889113,I889000,I91765);
nand I_52152 (I889130,I889113,I91771);
nor I_52153 (I889147,I888924,I889130);
DFFARX1 I_52154 (I889147,I2507,I888898,I888863,);
not I_52155 (I889178,I889130);
nand I_52156 (I888875,I888941,I889178);
DFFARX1 I_52157 (I889130,I2507,I888898,I889218,);
not I_52158 (I889226,I889218);
not I_52159 (I889243,I91765);
not I_52160 (I889260,I91753);
nor I_52161 (I889277,I889260,I91759);
nor I_52162 (I888890,I889226,I889277);
nor I_52163 (I889308,I889260,I91762);
and I_52164 (I889325,I889308,I91750);
or I_52165 (I889342,I889325,I91768);
DFFARX1 I_52166 (I889342,I2507,I888898,I889368,);
nor I_52167 (I888878,I889368,I888924);
not I_52168 (I889390,I889368);
and I_52169 (I889407,I889390,I888924);
nor I_52170 (I888872,I888949,I889407);
nand I_52171 (I889438,I889390,I889000);
nor I_52172 (I888866,I889260,I889438);
nand I_52173 (I888869,I889390,I889178);
nand I_52174 (I889483,I889000,I91753);
nor I_52175 (I888881,I889243,I889483);
not I_52176 (I889544,I2514);
DFFARX1 I_52177 (I220446,I2507,I889544,I889570,);
DFFARX1 I_52178 (I220458,I2507,I889544,I889587,);
not I_52179 (I889595,I889587);
not I_52180 (I889612,I220464);
nor I_52181 (I889629,I889612,I220449);
not I_52182 (I889646,I220440);
nor I_52183 (I889663,I889629,I220461);
nor I_52184 (I889680,I889587,I889663);
DFFARX1 I_52185 (I889680,I2507,I889544,I889530,);
nor I_52186 (I889711,I220461,I220449);
nand I_52187 (I889728,I889711,I220464);
DFFARX1 I_52188 (I889728,I2507,I889544,I889533,);
nor I_52189 (I889759,I889646,I220461);
nand I_52190 (I889776,I889759,I220443);
nor I_52191 (I889793,I889570,I889776);
DFFARX1 I_52192 (I889793,I2507,I889544,I889509,);
not I_52193 (I889824,I889776);
nand I_52194 (I889521,I889587,I889824);
DFFARX1 I_52195 (I889776,I2507,I889544,I889864,);
not I_52196 (I889872,I889864);
not I_52197 (I889889,I220461);
not I_52198 (I889906,I220452);
nor I_52199 (I889923,I889906,I220440);
nor I_52200 (I889536,I889872,I889923);
nor I_52201 (I889954,I889906,I220455);
and I_52202 (I889971,I889954,I220443);
or I_52203 (I889988,I889971,I220440);
DFFARX1 I_52204 (I889988,I2507,I889544,I890014,);
nor I_52205 (I889524,I890014,I889570);
not I_52206 (I890036,I890014);
and I_52207 (I890053,I890036,I889570);
nor I_52208 (I889518,I889595,I890053);
nand I_52209 (I890084,I890036,I889646);
nor I_52210 (I889512,I889906,I890084);
nand I_52211 (I889515,I890036,I889824);
nand I_52212 (I890129,I889646,I220452);
nor I_52213 (I889527,I889889,I890129);
not I_52214 (I890190,I2514);
DFFARX1 I_52215 (I1133528,I2507,I890190,I890216,);
DFFARX1 I_52216 (I1133510,I2507,I890190,I890233,);
not I_52217 (I890241,I890233);
not I_52218 (I890258,I1133519);
nor I_52219 (I890275,I890258,I1133531);
not I_52220 (I890292,I1133513);
nor I_52221 (I890309,I890275,I1133522);
nor I_52222 (I890326,I890233,I890309);
DFFARX1 I_52223 (I890326,I2507,I890190,I890176,);
nor I_52224 (I890357,I1133522,I1133531);
nand I_52225 (I890374,I890357,I1133519);
DFFARX1 I_52226 (I890374,I2507,I890190,I890179,);
nor I_52227 (I890405,I890292,I1133522);
nand I_52228 (I890422,I890405,I1133534);
nor I_52229 (I890439,I890216,I890422);
DFFARX1 I_52230 (I890439,I2507,I890190,I890155,);
not I_52231 (I890470,I890422);
nand I_52232 (I890167,I890233,I890470);
DFFARX1 I_52233 (I890422,I2507,I890190,I890510,);
not I_52234 (I890518,I890510);
not I_52235 (I890535,I1133522);
not I_52236 (I890552,I1133510);
nor I_52237 (I890569,I890552,I1133513);
nor I_52238 (I890182,I890518,I890569);
nor I_52239 (I890600,I890552,I1133516);
and I_52240 (I890617,I890600,I1133525);
or I_52241 (I890634,I890617,I1133513);
DFFARX1 I_52242 (I890634,I2507,I890190,I890660,);
nor I_52243 (I890170,I890660,I890216);
not I_52244 (I890682,I890660);
and I_52245 (I890699,I890682,I890216);
nor I_52246 (I890164,I890241,I890699);
nand I_52247 (I890730,I890682,I890292);
nor I_52248 (I890158,I890552,I890730);
nand I_52249 (I890161,I890682,I890470);
nand I_52250 (I890775,I890292,I1133510);
nor I_52251 (I890173,I890535,I890775);
not I_52252 (I890836,I2514);
DFFARX1 I_52253 (I445781,I2507,I890836,I890862,);
DFFARX1 I_52254 (I445778,I2507,I890836,I890879,);
not I_52255 (I890887,I890879);
not I_52256 (I890904,I445793);
nor I_52257 (I890921,I890904,I445796);
not I_52258 (I890938,I445784);
nor I_52259 (I890955,I890921,I445790);
nor I_52260 (I890972,I890879,I890955);
DFFARX1 I_52261 (I890972,I2507,I890836,I890822,);
nor I_52262 (I891003,I445790,I445796);
nand I_52263 (I891020,I891003,I445793);
DFFARX1 I_52264 (I891020,I2507,I890836,I890825,);
nor I_52265 (I891051,I890938,I445790);
nand I_52266 (I891068,I891051,I445802);
nor I_52267 (I891085,I890862,I891068);
DFFARX1 I_52268 (I891085,I2507,I890836,I890801,);
not I_52269 (I891116,I891068);
nand I_52270 (I890813,I890879,I891116);
DFFARX1 I_52271 (I891068,I2507,I890836,I891156,);
not I_52272 (I891164,I891156);
not I_52273 (I891181,I445790);
not I_52274 (I891198,I445775);
nor I_52275 (I891215,I891198,I445784);
nor I_52276 (I890828,I891164,I891215);
nor I_52277 (I891246,I891198,I445787);
and I_52278 (I891263,I891246,I445775);
or I_52279 (I891280,I891263,I445799);
DFFARX1 I_52280 (I891280,I2507,I890836,I891306,);
nor I_52281 (I890816,I891306,I890862);
not I_52282 (I891328,I891306);
and I_52283 (I891345,I891328,I890862);
nor I_52284 (I890810,I890887,I891345);
nand I_52285 (I891376,I891328,I890938);
nor I_52286 (I890804,I891198,I891376);
nand I_52287 (I890807,I891328,I891116);
nand I_52288 (I891421,I890938,I445775);
nor I_52289 (I890819,I891181,I891421);
not I_52290 (I891482,I2514);
DFFARX1 I_52291 (I704130,I2507,I891482,I891508,);
DFFARX1 I_52292 (I704124,I2507,I891482,I891525,);
not I_52293 (I891533,I891525);
not I_52294 (I891550,I704139);
nor I_52295 (I891567,I891550,I704124);
not I_52296 (I891584,I704133);
nor I_52297 (I891601,I891567,I704142);
nor I_52298 (I891618,I891525,I891601);
DFFARX1 I_52299 (I891618,I2507,I891482,I891468,);
nor I_52300 (I891649,I704142,I704124);
nand I_52301 (I891666,I891649,I704139);
DFFARX1 I_52302 (I891666,I2507,I891482,I891471,);
nor I_52303 (I891697,I891584,I704142);
nand I_52304 (I891714,I891697,I704127);
nor I_52305 (I891731,I891508,I891714);
DFFARX1 I_52306 (I891731,I2507,I891482,I891447,);
not I_52307 (I891762,I891714);
nand I_52308 (I891459,I891525,I891762);
DFFARX1 I_52309 (I891714,I2507,I891482,I891802,);
not I_52310 (I891810,I891802);
not I_52311 (I891827,I704142);
not I_52312 (I891844,I704136);
nor I_52313 (I891861,I891844,I704133);
nor I_52314 (I891474,I891810,I891861);
nor I_52315 (I891892,I891844,I704145);
and I_52316 (I891909,I891892,I704148);
or I_52317 (I891926,I891909,I704127);
DFFARX1 I_52318 (I891926,I2507,I891482,I891952,);
nor I_52319 (I891462,I891952,I891508);
not I_52320 (I891974,I891952);
and I_52321 (I891991,I891974,I891508);
nor I_52322 (I891456,I891533,I891991);
nand I_52323 (I892022,I891974,I891584);
nor I_52324 (I891450,I891844,I892022);
nand I_52325 (I891453,I891974,I891762);
nand I_52326 (I892067,I891584,I704136);
nor I_52327 (I891465,I891827,I892067);
not I_52328 (I892128,I2514);
DFFARX1 I_52329 (I109668,I2507,I892128,I892154,);
DFFARX1 I_52330 (I109674,I2507,I892128,I892171,);
not I_52331 (I892179,I892171);
not I_52332 (I892196,I109692);
nor I_52333 (I892213,I892196,I109671);
not I_52334 (I892230,I109677);
nor I_52335 (I892247,I892213,I109683);
nor I_52336 (I892264,I892171,I892247);
DFFARX1 I_52337 (I892264,I2507,I892128,I892114,);
nor I_52338 (I892295,I109683,I109671);
nand I_52339 (I892312,I892295,I109692);
DFFARX1 I_52340 (I892312,I2507,I892128,I892117,);
nor I_52341 (I892343,I892230,I109683);
nand I_52342 (I892360,I892343,I109689);
nor I_52343 (I892377,I892154,I892360);
DFFARX1 I_52344 (I892377,I2507,I892128,I892093,);
not I_52345 (I892408,I892360);
nand I_52346 (I892105,I892171,I892408);
DFFARX1 I_52347 (I892360,I2507,I892128,I892448,);
not I_52348 (I892456,I892448);
not I_52349 (I892473,I109683);
not I_52350 (I892490,I109671);
nor I_52351 (I892507,I892490,I109677);
nor I_52352 (I892120,I892456,I892507);
nor I_52353 (I892538,I892490,I109680);
and I_52354 (I892555,I892538,I109668);
or I_52355 (I892572,I892555,I109686);
DFFARX1 I_52356 (I892572,I2507,I892128,I892598,);
nor I_52357 (I892108,I892598,I892154);
not I_52358 (I892620,I892598);
and I_52359 (I892637,I892620,I892154);
nor I_52360 (I892102,I892179,I892637);
nand I_52361 (I892668,I892620,I892230);
nor I_52362 (I892096,I892490,I892668);
nand I_52363 (I892099,I892620,I892408);
nand I_52364 (I892713,I892230,I109671);
nor I_52365 (I892111,I892473,I892713);
not I_52366 (I892774,I2514);
DFFARX1 I_52367 (I518487,I2507,I892774,I892800,);
DFFARX1 I_52368 (I518499,I2507,I892774,I892817,);
not I_52369 (I892825,I892817);
not I_52370 (I892842,I518484);
nor I_52371 (I892859,I892842,I518502);
not I_52372 (I892876,I518508);
nor I_52373 (I892893,I892859,I518490);
nor I_52374 (I892910,I892817,I892893);
DFFARX1 I_52375 (I892910,I2507,I892774,I892760,);
nor I_52376 (I892941,I518490,I518502);
nand I_52377 (I892958,I892941,I518484);
DFFARX1 I_52378 (I892958,I2507,I892774,I892763,);
nor I_52379 (I892989,I892876,I518490);
nand I_52380 (I893006,I892989,I518493);
nor I_52381 (I893023,I892800,I893006);
DFFARX1 I_52382 (I893023,I2507,I892774,I892739,);
not I_52383 (I893054,I893006);
nand I_52384 (I892751,I892817,I893054);
DFFARX1 I_52385 (I893006,I2507,I892774,I893094,);
not I_52386 (I893102,I893094);
not I_52387 (I893119,I518490);
not I_52388 (I893136,I518496);
nor I_52389 (I893153,I893136,I518508);
nor I_52390 (I892766,I893102,I893153);
nor I_52391 (I893184,I893136,I518505);
and I_52392 (I893201,I893184,I518484);
or I_52393 (I893218,I893201,I518487);
DFFARX1 I_52394 (I893218,I2507,I892774,I893244,);
nor I_52395 (I892754,I893244,I892800);
not I_52396 (I893266,I893244);
and I_52397 (I893283,I893266,I892800);
nor I_52398 (I892748,I892825,I893283);
nand I_52399 (I893314,I893266,I892876);
nor I_52400 (I892742,I893136,I893314);
nand I_52401 (I892745,I893266,I893054);
nand I_52402 (I893359,I892876,I518496);
nor I_52403 (I892757,I893119,I893359);
not I_52404 (I893420,I2514);
DFFARX1 I_52405 (I213901,I2507,I893420,I893446,);
DFFARX1 I_52406 (I213913,I2507,I893420,I893463,);
not I_52407 (I893471,I893463);
not I_52408 (I893488,I213919);
nor I_52409 (I893505,I893488,I213904);
not I_52410 (I893522,I213895);
nor I_52411 (I893539,I893505,I213916);
nor I_52412 (I893556,I893463,I893539);
DFFARX1 I_52413 (I893556,I2507,I893420,I893406,);
nor I_52414 (I893587,I213916,I213904);
nand I_52415 (I893604,I893587,I213919);
DFFARX1 I_52416 (I893604,I2507,I893420,I893409,);
nor I_52417 (I893635,I893522,I213916);
nand I_52418 (I893652,I893635,I213898);
nor I_52419 (I893669,I893446,I893652);
DFFARX1 I_52420 (I893669,I2507,I893420,I893385,);
not I_52421 (I893700,I893652);
nand I_52422 (I893397,I893463,I893700);
DFFARX1 I_52423 (I893652,I2507,I893420,I893740,);
not I_52424 (I893748,I893740);
not I_52425 (I893765,I213916);
not I_52426 (I893782,I213907);
nor I_52427 (I893799,I893782,I213895);
nor I_52428 (I893412,I893748,I893799);
nor I_52429 (I893830,I893782,I213910);
and I_52430 (I893847,I893830,I213898);
or I_52431 (I893864,I893847,I213895);
DFFARX1 I_52432 (I893864,I2507,I893420,I893890,);
nor I_52433 (I893400,I893890,I893446);
not I_52434 (I893912,I893890);
and I_52435 (I893929,I893912,I893446);
nor I_52436 (I893394,I893471,I893929);
nand I_52437 (I893960,I893912,I893522);
nor I_52438 (I893388,I893782,I893960);
nand I_52439 (I893391,I893912,I893700);
nand I_52440 (I894005,I893522,I213907);
nor I_52441 (I893403,I893765,I894005);
not I_52442 (I894066,I2514);
DFFARX1 I_52443 (I31145,I2507,I894066,I894092,);
DFFARX1 I_52444 (I31151,I2507,I894066,I894109,);
not I_52445 (I894117,I894109);
not I_52446 (I894134,I31145);
nor I_52447 (I894151,I894134,I31157);
not I_52448 (I894168,I31169);
nor I_52449 (I894185,I894151,I31163);
nor I_52450 (I894202,I894109,I894185);
DFFARX1 I_52451 (I894202,I2507,I894066,I894052,);
nor I_52452 (I894233,I31163,I31157);
nand I_52453 (I894250,I894233,I31145);
DFFARX1 I_52454 (I894250,I2507,I894066,I894055,);
nor I_52455 (I894281,I894168,I31163);
nand I_52456 (I894298,I894281,I31148);
nor I_52457 (I894315,I894092,I894298);
DFFARX1 I_52458 (I894315,I2507,I894066,I894031,);
not I_52459 (I894346,I894298);
nand I_52460 (I894043,I894109,I894346);
DFFARX1 I_52461 (I894298,I2507,I894066,I894386,);
not I_52462 (I894394,I894386);
not I_52463 (I894411,I31163);
not I_52464 (I894428,I31148);
nor I_52465 (I894445,I894428,I31169);
nor I_52466 (I894058,I894394,I894445);
nor I_52467 (I894476,I894428,I31166);
and I_52468 (I894493,I894476,I31160);
or I_52469 (I894510,I894493,I31154);
DFFARX1 I_52470 (I894510,I2507,I894066,I894536,);
nor I_52471 (I894046,I894536,I894092);
not I_52472 (I894558,I894536);
and I_52473 (I894575,I894558,I894092);
nor I_52474 (I894040,I894117,I894575);
nand I_52475 (I894606,I894558,I894168);
nor I_52476 (I894034,I894428,I894606);
nand I_52477 (I894037,I894558,I894346);
nand I_52478 (I894651,I894168,I31148);
nor I_52479 (I894049,I894411,I894651);
not I_52480 (I894712,I2514);
DFFARX1 I_52481 (I1185548,I2507,I894712,I894738,);
DFFARX1 I_52482 (I1185530,I2507,I894712,I894755,);
not I_52483 (I894763,I894755);
not I_52484 (I894780,I1185539);
nor I_52485 (I894797,I894780,I1185551);
not I_52486 (I894814,I1185533);
nor I_52487 (I894831,I894797,I1185542);
nor I_52488 (I894848,I894755,I894831);
DFFARX1 I_52489 (I894848,I2507,I894712,I894698,);
nor I_52490 (I894879,I1185542,I1185551);
nand I_52491 (I894896,I894879,I1185539);
DFFARX1 I_52492 (I894896,I2507,I894712,I894701,);
nor I_52493 (I894927,I894814,I1185542);
nand I_52494 (I894944,I894927,I1185554);
nor I_52495 (I894961,I894738,I894944);
DFFARX1 I_52496 (I894961,I2507,I894712,I894677,);
not I_52497 (I894992,I894944);
nand I_52498 (I894689,I894755,I894992);
DFFARX1 I_52499 (I894944,I2507,I894712,I895032,);
not I_52500 (I895040,I895032);
not I_52501 (I895057,I1185542);
not I_52502 (I895074,I1185530);
nor I_52503 (I895091,I895074,I1185533);
nor I_52504 (I894704,I895040,I895091);
nor I_52505 (I895122,I895074,I1185536);
and I_52506 (I895139,I895122,I1185545);
or I_52507 (I895156,I895139,I1185533);
DFFARX1 I_52508 (I895156,I2507,I894712,I895182,);
nor I_52509 (I894692,I895182,I894738);
not I_52510 (I895204,I895182);
and I_52511 (I895221,I895204,I894738);
nor I_52512 (I894686,I894763,I895221);
nand I_52513 (I895252,I895204,I894814);
nor I_52514 (I894680,I895074,I895252);
nand I_52515 (I894683,I895204,I894992);
nand I_52516 (I895297,I894814,I1185530);
nor I_52517 (I894695,I895057,I895297);
not I_52518 (I895358,I2514);
DFFARX1 I_52519 (I1033703,I2507,I895358,I895384,);
DFFARX1 I_52520 (I1033706,I2507,I895358,I895401,);
not I_52521 (I895409,I895401);
not I_52522 (I895426,I1033703);
nor I_52523 (I895443,I895426,I1033715);
not I_52524 (I895460,I1033724);
nor I_52525 (I895477,I895443,I1033712);
nor I_52526 (I895494,I895401,I895477);
DFFARX1 I_52527 (I895494,I2507,I895358,I895344,);
nor I_52528 (I895525,I1033712,I1033715);
nand I_52529 (I895542,I895525,I1033703);
DFFARX1 I_52530 (I895542,I2507,I895358,I895347,);
nor I_52531 (I895573,I895460,I1033712);
nand I_52532 (I895590,I895573,I1033718);
nor I_52533 (I895607,I895384,I895590);
DFFARX1 I_52534 (I895607,I2507,I895358,I895323,);
not I_52535 (I895638,I895590);
nand I_52536 (I895335,I895401,I895638);
DFFARX1 I_52537 (I895590,I2507,I895358,I895678,);
not I_52538 (I895686,I895678);
not I_52539 (I895703,I1033712);
not I_52540 (I895720,I1033709);
nor I_52541 (I895737,I895720,I1033724);
nor I_52542 (I895350,I895686,I895737);
nor I_52543 (I895768,I895720,I1033721);
and I_52544 (I895785,I895768,I1033709);
or I_52545 (I895802,I895785,I1033706);
DFFARX1 I_52546 (I895802,I2507,I895358,I895828,);
nor I_52547 (I895338,I895828,I895384);
not I_52548 (I895850,I895828);
and I_52549 (I895867,I895850,I895384);
nor I_52550 (I895332,I895409,I895867);
nand I_52551 (I895898,I895850,I895460);
nor I_52552 (I895326,I895720,I895898);
nand I_52553 (I895329,I895850,I895638);
nand I_52554 (I895943,I895460,I1033709);
nor I_52555 (I895341,I895703,I895943);
not I_52556 (I896004,I2514);
DFFARX1 I_52557 (I831766,I2507,I896004,I896030,);
DFFARX1 I_52558 (I831763,I2507,I896004,I896047,);
not I_52559 (I896055,I896047);
not I_52560 (I896072,I831763);
nor I_52561 (I896089,I896072,I831766);
not I_52562 (I896106,I831778);
nor I_52563 (I896123,I896089,I831772);
nor I_52564 (I896140,I896047,I896123);
DFFARX1 I_52565 (I896140,I2507,I896004,I895990,);
nor I_52566 (I896171,I831772,I831766);
nand I_52567 (I896188,I896171,I831763);
DFFARX1 I_52568 (I896188,I2507,I896004,I895993,);
nor I_52569 (I896219,I896106,I831772);
nand I_52570 (I896236,I896219,I831760);
nor I_52571 (I896253,I896030,I896236);
DFFARX1 I_52572 (I896253,I2507,I896004,I895969,);
not I_52573 (I896284,I896236);
nand I_52574 (I895981,I896047,I896284);
DFFARX1 I_52575 (I896236,I2507,I896004,I896324,);
not I_52576 (I896332,I896324);
not I_52577 (I896349,I831772);
not I_52578 (I896366,I831769);
nor I_52579 (I896383,I896366,I831778);
nor I_52580 (I895996,I896332,I896383);
nor I_52581 (I896414,I896366,I831775);
and I_52582 (I896431,I896414,I831781);
or I_52583 (I896448,I896431,I831760);
DFFARX1 I_52584 (I896448,I2507,I896004,I896474,);
nor I_52585 (I895984,I896474,I896030);
not I_52586 (I896496,I896474);
and I_52587 (I896513,I896496,I896030);
nor I_52588 (I895978,I896055,I896513);
nand I_52589 (I896544,I896496,I896106);
nor I_52590 (I895972,I896366,I896544);
nand I_52591 (I895975,I896496,I896284);
nand I_52592 (I896589,I896106,I831769);
nor I_52593 (I895987,I896349,I896589);
not I_52594 (I896650,I2514);
DFFARX1 I_52595 (I446325,I2507,I896650,I896676,);
DFFARX1 I_52596 (I446322,I2507,I896650,I896693,);
not I_52597 (I896701,I896693);
not I_52598 (I896718,I446337);
nor I_52599 (I896735,I896718,I446340);
not I_52600 (I896752,I446328);
nor I_52601 (I896769,I896735,I446334);
nor I_52602 (I896786,I896693,I896769);
DFFARX1 I_52603 (I896786,I2507,I896650,I896636,);
nor I_52604 (I896817,I446334,I446340);
nand I_52605 (I896834,I896817,I446337);
DFFARX1 I_52606 (I896834,I2507,I896650,I896639,);
nor I_52607 (I896865,I896752,I446334);
nand I_52608 (I896882,I896865,I446346);
nor I_52609 (I896899,I896676,I896882);
DFFARX1 I_52610 (I896899,I2507,I896650,I896615,);
not I_52611 (I896930,I896882);
nand I_52612 (I896627,I896693,I896930);
DFFARX1 I_52613 (I896882,I2507,I896650,I896970,);
not I_52614 (I896978,I896970);
not I_52615 (I896995,I446334);
not I_52616 (I897012,I446319);
nor I_52617 (I897029,I897012,I446328);
nor I_52618 (I896642,I896978,I897029);
nor I_52619 (I897060,I897012,I446331);
and I_52620 (I897077,I897060,I446319);
or I_52621 (I897094,I897077,I446343);
DFFARX1 I_52622 (I897094,I2507,I896650,I897120,);
nor I_52623 (I896630,I897120,I896676);
not I_52624 (I897142,I897120);
and I_52625 (I897159,I897142,I896676);
nor I_52626 (I896624,I896701,I897159);
nand I_52627 (I897190,I897142,I896752);
nor I_52628 (I896618,I897012,I897190);
nand I_52629 (I896621,I897142,I896930);
nand I_52630 (I897235,I896752,I446319);
nor I_52631 (I896633,I896995,I897235);
not I_52632 (I897296,I2514);
DFFARX1 I_52633 (I229966,I2507,I897296,I897322,);
DFFARX1 I_52634 (I229978,I2507,I897296,I897339,);
not I_52635 (I897347,I897339);
not I_52636 (I897364,I229984);
nor I_52637 (I897381,I897364,I229969);
not I_52638 (I897398,I229960);
nor I_52639 (I897415,I897381,I229981);
nor I_52640 (I897432,I897339,I897415);
DFFARX1 I_52641 (I897432,I2507,I897296,I897282,);
nor I_52642 (I897463,I229981,I229969);
nand I_52643 (I897480,I897463,I229984);
DFFARX1 I_52644 (I897480,I2507,I897296,I897285,);
nor I_52645 (I897511,I897398,I229981);
nand I_52646 (I897528,I897511,I229963);
nor I_52647 (I897545,I897322,I897528);
DFFARX1 I_52648 (I897545,I2507,I897296,I897261,);
not I_52649 (I897576,I897528);
nand I_52650 (I897273,I897339,I897576);
DFFARX1 I_52651 (I897528,I2507,I897296,I897616,);
not I_52652 (I897624,I897616);
not I_52653 (I897641,I229981);
not I_52654 (I897658,I229972);
nor I_52655 (I897675,I897658,I229960);
nor I_52656 (I897288,I897624,I897675);
nor I_52657 (I897706,I897658,I229975);
and I_52658 (I897723,I897706,I229963);
or I_52659 (I897740,I897723,I229960);
DFFARX1 I_52660 (I897740,I2507,I897296,I897766,);
nor I_52661 (I897276,I897766,I897322);
not I_52662 (I897788,I897766);
and I_52663 (I897805,I897788,I897322);
nor I_52664 (I897270,I897347,I897805);
nand I_52665 (I897836,I897788,I897398);
nor I_52666 (I897264,I897658,I897836);
nand I_52667 (I897267,I897788,I897576);
nand I_52668 (I897881,I897398,I229972);
nor I_52669 (I897279,I897641,I897881);
not I_52670 (I897942,I2514);
DFFARX1 I_52671 (I320808,I2507,I897942,I897968,);
DFFARX1 I_52672 (I320814,I2507,I897942,I897985,);
not I_52673 (I897993,I897985);
not I_52674 (I898010,I320835);
nor I_52675 (I898027,I898010,I320823);
not I_52676 (I898044,I320832);
nor I_52677 (I898061,I898027,I320817);
nor I_52678 (I898078,I897985,I898061);
DFFARX1 I_52679 (I898078,I2507,I897942,I897928,);
nor I_52680 (I898109,I320817,I320823);
nand I_52681 (I898126,I898109,I320835);
DFFARX1 I_52682 (I898126,I2507,I897942,I897931,);
nor I_52683 (I898157,I898044,I320817);
nand I_52684 (I898174,I898157,I320808);
nor I_52685 (I898191,I897968,I898174);
DFFARX1 I_52686 (I898191,I2507,I897942,I897907,);
not I_52687 (I898222,I898174);
nand I_52688 (I897919,I897985,I898222);
DFFARX1 I_52689 (I898174,I2507,I897942,I898262,);
not I_52690 (I898270,I898262);
not I_52691 (I898287,I320817);
not I_52692 (I898304,I320820);
nor I_52693 (I898321,I898304,I320832);
nor I_52694 (I897934,I898270,I898321);
nor I_52695 (I898352,I898304,I320829);
and I_52696 (I898369,I898352,I320811);
or I_52697 (I898386,I898369,I320826);
DFFARX1 I_52698 (I898386,I2507,I897942,I898412,);
nor I_52699 (I897922,I898412,I897968);
not I_52700 (I898434,I898412);
and I_52701 (I898451,I898434,I897968);
nor I_52702 (I897916,I897993,I898451);
nand I_52703 (I898482,I898434,I898044);
nor I_52704 (I897910,I898304,I898482);
nand I_52705 (I897913,I898434,I898222);
nand I_52706 (I898527,I898044,I320820);
nor I_52707 (I897925,I898287,I898527);
not I_52708 (I898588,I2514);
DFFARX1 I_52709 (I1173988,I2507,I898588,I898614,);
DFFARX1 I_52710 (I1173970,I2507,I898588,I898631,);
not I_52711 (I898639,I898631);
not I_52712 (I898656,I1173979);
nor I_52713 (I898673,I898656,I1173991);
not I_52714 (I898690,I1173973);
nor I_52715 (I898707,I898673,I1173982);
nor I_52716 (I898724,I898631,I898707);
DFFARX1 I_52717 (I898724,I2507,I898588,I898574,);
nor I_52718 (I898755,I1173982,I1173991);
nand I_52719 (I898772,I898755,I1173979);
DFFARX1 I_52720 (I898772,I2507,I898588,I898577,);
nor I_52721 (I898803,I898690,I1173982);
nand I_52722 (I898820,I898803,I1173994);
nor I_52723 (I898837,I898614,I898820);
DFFARX1 I_52724 (I898837,I2507,I898588,I898553,);
not I_52725 (I898868,I898820);
nand I_52726 (I898565,I898631,I898868);
DFFARX1 I_52727 (I898820,I2507,I898588,I898908,);
not I_52728 (I898916,I898908);
not I_52729 (I898933,I1173982);
not I_52730 (I898950,I1173970);
nor I_52731 (I898967,I898950,I1173973);
nor I_52732 (I898580,I898916,I898967);
nor I_52733 (I898998,I898950,I1173976);
and I_52734 (I899015,I898998,I1173985);
or I_52735 (I899032,I899015,I1173973);
DFFARX1 I_52736 (I899032,I2507,I898588,I899058,);
nor I_52737 (I898568,I899058,I898614);
not I_52738 (I899080,I899058);
and I_52739 (I899097,I899080,I898614);
nor I_52740 (I898562,I898639,I899097);
nand I_52741 (I899128,I899080,I898690);
nor I_52742 (I898556,I898950,I899128);
nand I_52743 (I898559,I899080,I898868);
nand I_52744 (I899173,I898690,I1173970);
nor I_52745 (I898571,I898933,I899173);
not I_52746 (I899234,I2514);
DFFARX1 I_52747 (I599509,I2507,I899234,I899260,);
DFFARX1 I_52748 (I599521,I2507,I899234,I899277,);
not I_52749 (I899285,I899277);
not I_52750 (I899302,I599530);
nor I_52751 (I899319,I899302,I599506);
not I_52752 (I899336,I599524);
nor I_52753 (I899353,I899319,I599518);
nor I_52754 (I899370,I899277,I899353);
DFFARX1 I_52755 (I899370,I2507,I899234,I899220,);
nor I_52756 (I899401,I599518,I599506);
nand I_52757 (I899418,I899401,I599530);
DFFARX1 I_52758 (I899418,I2507,I899234,I899223,);
nor I_52759 (I899449,I899336,I599518);
nand I_52760 (I899466,I899449,I599512);
nor I_52761 (I899483,I899260,I899466);
DFFARX1 I_52762 (I899483,I2507,I899234,I899199,);
not I_52763 (I899514,I899466);
nand I_52764 (I899211,I899277,I899514);
DFFARX1 I_52765 (I899466,I2507,I899234,I899554,);
not I_52766 (I899562,I899554);
not I_52767 (I899579,I599518);
not I_52768 (I899596,I599527);
nor I_52769 (I899613,I899596,I599524);
nor I_52770 (I899226,I899562,I899613);
nor I_52771 (I899644,I899596,I599509);
and I_52772 (I899661,I899644,I599506);
or I_52773 (I899678,I899661,I599515);
DFFARX1 I_52774 (I899678,I2507,I899234,I899704,);
nor I_52775 (I899214,I899704,I899260);
not I_52776 (I899726,I899704);
and I_52777 (I899743,I899726,I899260);
nor I_52778 (I899208,I899285,I899743);
nand I_52779 (I899774,I899726,I899336);
nor I_52780 (I899202,I899596,I899774);
nand I_52781 (I899205,I899726,I899514);
nand I_52782 (I899819,I899336,I599527);
nor I_52783 (I899217,I899579,I899819);
not I_52784 (I899880,I2514);
DFFARX1 I_52785 (I202001,I2507,I899880,I899906,);
DFFARX1 I_52786 (I202013,I2507,I899880,I899923,);
not I_52787 (I899931,I899923);
not I_52788 (I899948,I202019);
nor I_52789 (I899965,I899948,I202004);
not I_52790 (I899982,I201995);
nor I_52791 (I899999,I899965,I202016);
nor I_52792 (I900016,I899923,I899999);
DFFARX1 I_52793 (I900016,I2507,I899880,I899866,);
nor I_52794 (I900047,I202016,I202004);
nand I_52795 (I900064,I900047,I202019);
DFFARX1 I_52796 (I900064,I2507,I899880,I899869,);
nor I_52797 (I900095,I899982,I202016);
nand I_52798 (I900112,I900095,I201998);
nor I_52799 (I900129,I899906,I900112);
DFFARX1 I_52800 (I900129,I2507,I899880,I899845,);
not I_52801 (I900160,I900112);
nand I_52802 (I899857,I899923,I900160);
DFFARX1 I_52803 (I900112,I2507,I899880,I900200,);
not I_52804 (I900208,I900200);
not I_52805 (I900225,I202016);
not I_52806 (I900242,I202007);
nor I_52807 (I900259,I900242,I201995);
nor I_52808 (I899872,I900208,I900259);
nor I_52809 (I900290,I900242,I202010);
and I_52810 (I900307,I900290,I201998);
or I_52811 (I900324,I900307,I201995);
DFFARX1 I_52812 (I900324,I2507,I899880,I900350,);
nor I_52813 (I899860,I900350,I899906);
not I_52814 (I900372,I900350);
and I_52815 (I900389,I900372,I899906);
nor I_52816 (I899854,I899931,I900389);
nand I_52817 (I900420,I900372,I899982);
nor I_52818 (I899848,I900242,I900420);
nand I_52819 (I899851,I900372,I900160);
nand I_52820 (I900465,I899982,I202007);
nor I_52821 (I899863,I900225,I900465);
not I_52822 (I900526,I2514);
DFFARX1 I_52823 (I1220500,I2507,I900526,I900552,);
DFFARX1 I_52824 (I1220506,I2507,I900526,I900569,);
not I_52825 (I900577,I900569);
not I_52826 (I900594,I1220503);
nor I_52827 (I900611,I900594,I1220482);
not I_52828 (I900628,I1220485);
nor I_52829 (I900645,I900611,I1220491);
nor I_52830 (I900662,I900569,I900645);
DFFARX1 I_52831 (I900662,I2507,I900526,I900512,);
nor I_52832 (I900693,I1220491,I1220482);
nand I_52833 (I900710,I900693,I1220503);
DFFARX1 I_52834 (I900710,I2507,I900526,I900515,);
nor I_52835 (I900741,I900628,I1220491);
nand I_52836 (I900758,I900741,I1220485);
nor I_52837 (I900775,I900552,I900758);
DFFARX1 I_52838 (I900775,I2507,I900526,I900491,);
not I_52839 (I900806,I900758);
nand I_52840 (I900503,I900569,I900806);
DFFARX1 I_52841 (I900758,I2507,I900526,I900846,);
not I_52842 (I900854,I900846);
not I_52843 (I900871,I1220491);
not I_52844 (I900888,I1220494);
nor I_52845 (I900905,I900888,I1220485);
nor I_52846 (I900518,I900854,I900905);
nor I_52847 (I900936,I900888,I1220482);
and I_52848 (I900953,I900936,I1220488);
or I_52849 (I900970,I900953,I1220497);
DFFARX1 I_52850 (I900970,I2507,I900526,I900996,);
nor I_52851 (I900506,I900996,I900552);
not I_52852 (I901018,I900996);
and I_52853 (I901035,I901018,I900552);
nor I_52854 (I900500,I900577,I901035);
nand I_52855 (I901066,I901018,I900628);
nor I_52856 (I900494,I900888,I901066);
nand I_52857 (I900497,I901018,I900806);
nand I_52858 (I901111,I900628,I1220494);
nor I_52859 (I900509,I900871,I901111);
not I_52860 (I901172,I2514);
DFFARX1 I_52861 (I701818,I2507,I901172,I901198,);
DFFARX1 I_52862 (I701812,I2507,I901172,I901215,);
not I_52863 (I901223,I901215);
not I_52864 (I901240,I701827);
nor I_52865 (I901257,I901240,I701812);
not I_52866 (I901274,I701821);
nor I_52867 (I901291,I901257,I701830);
nor I_52868 (I901308,I901215,I901291);
DFFARX1 I_52869 (I901308,I2507,I901172,I901158,);
nor I_52870 (I901339,I701830,I701812);
nand I_52871 (I901356,I901339,I701827);
DFFARX1 I_52872 (I901356,I2507,I901172,I901161,);
nor I_52873 (I901387,I901274,I701830);
nand I_52874 (I901404,I901387,I701815);
nor I_52875 (I901421,I901198,I901404);
DFFARX1 I_52876 (I901421,I2507,I901172,I901137,);
not I_52877 (I901452,I901404);
nand I_52878 (I901149,I901215,I901452);
DFFARX1 I_52879 (I901404,I2507,I901172,I901492,);
not I_52880 (I901500,I901492);
not I_52881 (I901517,I701830);
not I_52882 (I901534,I701824);
nor I_52883 (I901551,I901534,I701821);
nor I_52884 (I901164,I901500,I901551);
nor I_52885 (I901582,I901534,I701833);
and I_52886 (I901599,I901582,I701836);
or I_52887 (I901616,I901599,I701815);
DFFARX1 I_52888 (I901616,I2507,I901172,I901642,);
nor I_52889 (I901152,I901642,I901198);
not I_52890 (I901664,I901642);
and I_52891 (I901681,I901664,I901198);
nor I_52892 (I901146,I901223,I901681);
nand I_52893 (I901712,I901664,I901274);
nor I_52894 (I901140,I901534,I901712);
nand I_52895 (I901143,I901664,I901452);
nand I_52896 (I901757,I901274,I701824);
nor I_52897 (I901155,I901517,I901757);
not I_52898 (I901818,I2514);
DFFARX1 I_52899 (I136563,I2507,I901818,I901844,);
DFFARX1 I_52900 (I136566,I2507,I901818,I901861,);
not I_52901 (I901869,I901861);
not I_52902 (I901886,I136551);
nor I_52903 (I901903,I901886,I136545);
not I_52904 (I901920,I136554);
nor I_52905 (I901937,I901903,I136569);
nor I_52906 (I901954,I901861,I901937);
DFFARX1 I_52907 (I901954,I2507,I901818,I901804,);
nor I_52908 (I901985,I136569,I136545);
nand I_52909 (I902002,I901985,I136551);
DFFARX1 I_52910 (I902002,I2507,I901818,I901807,);
nor I_52911 (I902033,I901920,I136569);
nand I_52912 (I902050,I902033,I136572);
nor I_52913 (I902067,I901844,I902050);
DFFARX1 I_52914 (I902067,I2507,I901818,I901783,);
not I_52915 (I902098,I902050);
nand I_52916 (I901795,I901861,I902098);
DFFARX1 I_52917 (I902050,I2507,I901818,I902138,);
not I_52918 (I902146,I902138);
not I_52919 (I902163,I136569);
not I_52920 (I902180,I136548);
nor I_52921 (I902197,I902180,I136554);
nor I_52922 (I901810,I902146,I902197);
nor I_52923 (I902228,I902180,I136557);
and I_52924 (I902245,I902228,I136545);
or I_52925 (I902262,I902245,I136560);
DFFARX1 I_52926 (I902262,I2507,I901818,I902288,);
nor I_52927 (I901798,I902288,I901844);
not I_52928 (I902310,I902288);
and I_52929 (I902327,I902310,I901844);
nor I_52930 (I901792,I901869,I902327);
nand I_52931 (I902358,I902310,I901920);
nor I_52932 (I901786,I902180,I902358);
nand I_52933 (I901789,I902310,I902098);
nand I_52934 (I902403,I901920,I136548);
nor I_52935 (I901801,I902163,I902403);
not I_52936 (I902464,I2514);
DFFARX1 I_52937 (I437077,I2507,I902464,I902490,);
DFFARX1 I_52938 (I437074,I2507,I902464,I902507,);
not I_52939 (I902515,I902507);
not I_52940 (I902532,I437089);
nor I_52941 (I902549,I902532,I437092);
not I_52942 (I902566,I437080);
nor I_52943 (I902583,I902549,I437086);
nor I_52944 (I902600,I902507,I902583);
DFFARX1 I_52945 (I902600,I2507,I902464,I902450,);
nor I_52946 (I902631,I437086,I437092);
nand I_52947 (I902648,I902631,I437089);
DFFARX1 I_52948 (I902648,I2507,I902464,I902453,);
nor I_52949 (I902679,I902566,I437086);
nand I_52950 (I902696,I902679,I437098);
nor I_52951 (I902713,I902490,I902696);
DFFARX1 I_52952 (I902713,I2507,I902464,I902429,);
not I_52953 (I902744,I902696);
nand I_52954 (I902441,I902507,I902744);
DFFARX1 I_52955 (I902696,I2507,I902464,I902784,);
not I_52956 (I902792,I902784);
not I_52957 (I902809,I437086);
not I_52958 (I902826,I437071);
nor I_52959 (I902843,I902826,I437080);
nor I_52960 (I902456,I902792,I902843);
nor I_52961 (I902874,I902826,I437083);
and I_52962 (I902891,I902874,I437071);
or I_52963 (I902908,I902891,I437095);
DFFARX1 I_52964 (I902908,I2507,I902464,I902934,);
nor I_52965 (I902444,I902934,I902490);
not I_52966 (I902956,I902934);
and I_52967 (I902973,I902956,I902490);
nor I_52968 (I902438,I902515,I902973);
nand I_52969 (I903004,I902956,I902566);
nor I_52970 (I902432,I902826,I903004);
nand I_52971 (I902435,I902956,I902744);
nand I_52972 (I903049,I902566,I437071);
nor I_52973 (I902447,I902809,I903049);
not I_52974 (I903110,I2514);
DFFARX1 I_52975 (I616849,I2507,I903110,I903136,);
DFFARX1 I_52976 (I616861,I2507,I903110,I903153,);
not I_52977 (I903161,I903153);
not I_52978 (I903178,I616870);
nor I_52979 (I903195,I903178,I616846);
not I_52980 (I903212,I616864);
nor I_52981 (I903229,I903195,I616858);
nor I_52982 (I903246,I903153,I903229);
DFFARX1 I_52983 (I903246,I2507,I903110,I903096,);
nor I_52984 (I903277,I616858,I616846);
nand I_52985 (I903294,I903277,I616870);
DFFARX1 I_52986 (I903294,I2507,I903110,I903099,);
nor I_52987 (I903325,I903212,I616858);
nand I_52988 (I903342,I903325,I616852);
nor I_52989 (I903359,I903136,I903342);
DFFARX1 I_52990 (I903359,I2507,I903110,I903075,);
not I_52991 (I903390,I903342);
nand I_52992 (I903087,I903153,I903390);
DFFARX1 I_52993 (I903342,I2507,I903110,I903430,);
not I_52994 (I903438,I903430);
not I_52995 (I903455,I616858);
not I_52996 (I903472,I616867);
nor I_52997 (I903489,I903472,I616864);
nor I_52998 (I903102,I903438,I903489);
nor I_52999 (I903520,I903472,I616849);
and I_53000 (I903537,I903520,I616846);
or I_53001 (I903554,I903537,I616855);
DFFARX1 I_53002 (I903554,I2507,I903110,I903580,);
nor I_53003 (I903090,I903580,I903136);
not I_53004 (I903602,I903580);
and I_53005 (I903619,I903602,I903136);
nor I_53006 (I903084,I903161,I903619);
nand I_53007 (I903650,I903602,I903212);
nor I_53008 (I903078,I903472,I903650);
nand I_53009 (I903081,I903602,I903390);
nand I_53010 (I903695,I903212,I616867);
nor I_53011 (I903093,I903455,I903695);
not I_53012 (I903756,I2514);
DFFARX1 I_53013 (I1171676,I2507,I903756,I903782,);
DFFARX1 I_53014 (I1171658,I2507,I903756,I903799,);
not I_53015 (I903807,I903799);
not I_53016 (I903824,I1171667);
nor I_53017 (I903841,I903824,I1171679);
not I_53018 (I903858,I1171661);
nor I_53019 (I903875,I903841,I1171670);
nor I_53020 (I903892,I903799,I903875);
DFFARX1 I_53021 (I903892,I2507,I903756,I903742,);
nor I_53022 (I903923,I1171670,I1171679);
nand I_53023 (I903940,I903923,I1171667);
DFFARX1 I_53024 (I903940,I2507,I903756,I903745,);
nor I_53025 (I903971,I903858,I1171670);
nand I_53026 (I903988,I903971,I1171682);
nor I_53027 (I904005,I903782,I903988);
DFFARX1 I_53028 (I904005,I2507,I903756,I903721,);
not I_53029 (I904036,I903988);
nand I_53030 (I903733,I903799,I904036);
DFFARX1 I_53031 (I903988,I2507,I903756,I904076,);
not I_53032 (I904084,I904076);
not I_53033 (I904101,I1171670);
not I_53034 (I904118,I1171658);
nor I_53035 (I904135,I904118,I1171661);
nor I_53036 (I903748,I904084,I904135);
nor I_53037 (I904166,I904118,I1171664);
and I_53038 (I904183,I904166,I1171673);
or I_53039 (I904200,I904183,I1171661);
DFFARX1 I_53040 (I904200,I2507,I903756,I904226,);
nor I_53041 (I903736,I904226,I903782);
not I_53042 (I904248,I904226);
and I_53043 (I904265,I904248,I903782);
nor I_53044 (I903730,I903807,I904265);
nand I_53045 (I904296,I904248,I903858);
nor I_53046 (I903724,I904118,I904296);
nand I_53047 (I903727,I904248,I904036);
nand I_53048 (I904341,I903858,I1171658);
nor I_53049 (I903739,I904101,I904341);
not I_53050 (I904402,I2514);
DFFARX1 I_53051 (I587371,I2507,I904402,I904428,);
DFFARX1 I_53052 (I587383,I2507,I904402,I904445,);
not I_53053 (I904453,I904445);
not I_53054 (I904470,I587392);
nor I_53055 (I904487,I904470,I587368);
not I_53056 (I904504,I587386);
nor I_53057 (I904521,I904487,I587380);
nor I_53058 (I904538,I904445,I904521);
DFFARX1 I_53059 (I904538,I2507,I904402,I904388,);
nor I_53060 (I904569,I587380,I587368);
nand I_53061 (I904586,I904569,I587392);
DFFARX1 I_53062 (I904586,I2507,I904402,I904391,);
nor I_53063 (I904617,I904504,I587380);
nand I_53064 (I904634,I904617,I587374);
nor I_53065 (I904651,I904428,I904634);
DFFARX1 I_53066 (I904651,I2507,I904402,I904367,);
not I_53067 (I904682,I904634);
nand I_53068 (I904379,I904445,I904682);
DFFARX1 I_53069 (I904634,I2507,I904402,I904722,);
not I_53070 (I904730,I904722);
not I_53071 (I904747,I587380);
not I_53072 (I904764,I587389);
nor I_53073 (I904781,I904764,I587386);
nor I_53074 (I904394,I904730,I904781);
nor I_53075 (I904812,I904764,I587371);
and I_53076 (I904829,I904812,I587368);
or I_53077 (I904846,I904829,I587377);
DFFARX1 I_53078 (I904846,I2507,I904402,I904872,);
nor I_53079 (I904382,I904872,I904428);
not I_53080 (I904894,I904872);
and I_53081 (I904911,I904894,I904428);
nor I_53082 (I904376,I904453,I904911);
nand I_53083 (I904942,I904894,I904504);
nor I_53084 (I904370,I904764,I904942);
nand I_53085 (I904373,I904894,I904682);
nand I_53086 (I904987,I904504,I587389);
nor I_53087 (I904385,I904747,I904987);
not I_53088 (I905048,I2514);
DFFARX1 I_53089 (I222826,I2507,I905048,I905074,);
DFFARX1 I_53090 (I222838,I2507,I905048,I905091,);
not I_53091 (I905099,I905091);
not I_53092 (I905116,I222844);
nor I_53093 (I905133,I905116,I222829);
not I_53094 (I905150,I222820);
nor I_53095 (I905167,I905133,I222841);
nor I_53096 (I905184,I905091,I905167);
DFFARX1 I_53097 (I905184,I2507,I905048,I905034,);
nor I_53098 (I905215,I222841,I222829);
nand I_53099 (I905232,I905215,I222844);
DFFARX1 I_53100 (I905232,I2507,I905048,I905037,);
nor I_53101 (I905263,I905150,I222841);
nand I_53102 (I905280,I905263,I222823);
nor I_53103 (I905297,I905074,I905280);
DFFARX1 I_53104 (I905297,I2507,I905048,I905013,);
not I_53105 (I905328,I905280);
nand I_53106 (I905025,I905091,I905328);
DFFARX1 I_53107 (I905280,I2507,I905048,I905368,);
not I_53108 (I905376,I905368);
not I_53109 (I905393,I222841);
not I_53110 (I905410,I222832);
nor I_53111 (I905427,I905410,I222820);
nor I_53112 (I905040,I905376,I905427);
nor I_53113 (I905458,I905410,I222835);
and I_53114 (I905475,I905458,I222823);
or I_53115 (I905492,I905475,I222820);
DFFARX1 I_53116 (I905492,I2507,I905048,I905518,);
nor I_53117 (I905028,I905518,I905074);
not I_53118 (I905540,I905518);
and I_53119 (I905557,I905540,I905074);
nor I_53120 (I905022,I905099,I905557);
nand I_53121 (I905588,I905540,I905150);
nor I_53122 (I905016,I905410,I905588);
nand I_53123 (I905019,I905540,I905328);
nand I_53124 (I905633,I905150,I222832);
nor I_53125 (I905031,I905393,I905633);
not I_53126 (I905694,I2514);
DFFARX1 I_53127 (I26402,I2507,I905694,I905720,);
DFFARX1 I_53128 (I26408,I2507,I905694,I905737,);
not I_53129 (I905745,I905737);
not I_53130 (I905762,I26402);
nor I_53131 (I905779,I905762,I26414);
not I_53132 (I905796,I26426);
nor I_53133 (I905813,I905779,I26420);
nor I_53134 (I905830,I905737,I905813);
DFFARX1 I_53135 (I905830,I2507,I905694,I905680,);
nor I_53136 (I905861,I26420,I26414);
nand I_53137 (I905878,I905861,I26402);
DFFARX1 I_53138 (I905878,I2507,I905694,I905683,);
nor I_53139 (I905909,I905796,I26420);
nand I_53140 (I905926,I905909,I26405);
nor I_53141 (I905943,I905720,I905926);
DFFARX1 I_53142 (I905943,I2507,I905694,I905659,);
not I_53143 (I905974,I905926);
nand I_53144 (I905671,I905737,I905974);
DFFARX1 I_53145 (I905926,I2507,I905694,I906014,);
not I_53146 (I906022,I906014);
not I_53147 (I906039,I26420);
not I_53148 (I906056,I26405);
nor I_53149 (I906073,I906056,I26426);
nor I_53150 (I905686,I906022,I906073);
nor I_53151 (I906104,I906056,I26423);
and I_53152 (I906121,I906104,I26417);
or I_53153 (I906138,I906121,I26411);
DFFARX1 I_53154 (I906138,I2507,I905694,I906164,);
nor I_53155 (I905674,I906164,I905720);
not I_53156 (I906186,I906164);
and I_53157 (I906203,I906186,I905720);
nor I_53158 (I905668,I905745,I906203);
nand I_53159 (I906234,I906186,I905796);
nor I_53160 (I905662,I906056,I906234);
nand I_53161 (I905665,I906186,I905974);
nand I_53162 (I906279,I905796,I26405);
nor I_53163 (I905677,I906039,I906279);
not I_53164 (I906340,I2514);
DFFARX1 I_53165 (I1102316,I2507,I906340,I906366,);
DFFARX1 I_53166 (I1102298,I2507,I906340,I906383,);
not I_53167 (I906391,I906383);
not I_53168 (I906408,I1102307);
nor I_53169 (I906425,I906408,I1102319);
not I_53170 (I906442,I1102301);
nor I_53171 (I906459,I906425,I1102310);
nor I_53172 (I906476,I906383,I906459);
DFFARX1 I_53173 (I906476,I2507,I906340,I906326,);
nor I_53174 (I906507,I1102310,I1102319);
nand I_53175 (I906524,I906507,I1102307);
DFFARX1 I_53176 (I906524,I2507,I906340,I906329,);
nor I_53177 (I906555,I906442,I1102310);
nand I_53178 (I906572,I906555,I1102322);
nor I_53179 (I906589,I906366,I906572);
DFFARX1 I_53180 (I906589,I2507,I906340,I906305,);
not I_53181 (I906620,I906572);
nand I_53182 (I906317,I906383,I906620);
DFFARX1 I_53183 (I906572,I2507,I906340,I906660,);
not I_53184 (I906668,I906660);
not I_53185 (I906685,I1102310);
not I_53186 (I906702,I1102298);
nor I_53187 (I906719,I906702,I1102301);
nor I_53188 (I906332,I906668,I906719);
nor I_53189 (I906750,I906702,I1102304);
and I_53190 (I906767,I906750,I1102313);
or I_53191 (I906784,I906767,I1102301);
DFFARX1 I_53192 (I906784,I2507,I906340,I906810,);
nor I_53193 (I906320,I906810,I906366);
not I_53194 (I906832,I906810);
and I_53195 (I906849,I906832,I906366);
nor I_53196 (I906314,I906391,I906849);
nand I_53197 (I906880,I906832,I906442);
nor I_53198 (I906308,I906702,I906880);
nand I_53199 (I906311,I906832,I906620);
nand I_53200 (I906925,I906442,I1102298);
nor I_53201 (I906323,I906685,I906925);
not I_53202 (I906986,I2514);
DFFARX1 I_53203 (I101236,I2507,I906986,I907012,);
DFFARX1 I_53204 (I101242,I2507,I906986,I907029,);
not I_53205 (I907037,I907029);
not I_53206 (I907054,I101260);
nor I_53207 (I907071,I907054,I101239);
not I_53208 (I907088,I101245);
nor I_53209 (I907105,I907071,I101251);
nor I_53210 (I907122,I907029,I907105);
DFFARX1 I_53211 (I907122,I2507,I906986,I906972,);
nor I_53212 (I907153,I101251,I101239);
nand I_53213 (I907170,I907153,I101260);
DFFARX1 I_53214 (I907170,I2507,I906986,I906975,);
nor I_53215 (I907201,I907088,I101251);
nand I_53216 (I907218,I907201,I101257);
nor I_53217 (I907235,I907012,I907218);
DFFARX1 I_53218 (I907235,I2507,I906986,I906951,);
not I_53219 (I907266,I907218);
nand I_53220 (I906963,I907029,I907266);
DFFARX1 I_53221 (I907218,I2507,I906986,I907306,);
not I_53222 (I907314,I907306);
not I_53223 (I907331,I101251);
not I_53224 (I907348,I101239);
nor I_53225 (I907365,I907348,I101245);
nor I_53226 (I906978,I907314,I907365);
nor I_53227 (I907396,I907348,I101248);
and I_53228 (I907413,I907396,I101236);
or I_53229 (I907430,I907413,I101254);
DFFARX1 I_53230 (I907430,I2507,I906986,I907456,);
nor I_53231 (I906966,I907456,I907012);
not I_53232 (I907478,I907456);
and I_53233 (I907495,I907478,I907012);
nor I_53234 (I906960,I907037,I907495);
nand I_53235 (I907526,I907478,I907088);
nor I_53236 (I906954,I907348,I907526);
nand I_53237 (I906957,I907478,I907266);
nand I_53238 (I907571,I907088,I101239);
nor I_53239 (I906969,I907331,I907571);
not I_53240 (I907632,I2514);
DFFARX1 I_53241 (I646330,I2507,I907632,I907658,);
DFFARX1 I_53242 (I646324,I2507,I907632,I907675,);
not I_53243 (I907683,I907675);
not I_53244 (I907700,I646339);
nor I_53245 (I907717,I907700,I646324);
not I_53246 (I907734,I646333);
nor I_53247 (I907751,I907717,I646342);
nor I_53248 (I907768,I907675,I907751);
DFFARX1 I_53249 (I907768,I2507,I907632,I907618,);
nor I_53250 (I907799,I646342,I646324);
nand I_53251 (I907816,I907799,I646339);
DFFARX1 I_53252 (I907816,I2507,I907632,I907621,);
nor I_53253 (I907847,I907734,I646342);
nand I_53254 (I907864,I907847,I646327);
nor I_53255 (I907881,I907658,I907864);
DFFARX1 I_53256 (I907881,I2507,I907632,I907597,);
not I_53257 (I907912,I907864);
nand I_53258 (I907609,I907675,I907912);
DFFARX1 I_53259 (I907864,I2507,I907632,I907952,);
not I_53260 (I907960,I907952);
not I_53261 (I907977,I646342);
not I_53262 (I907994,I646336);
nor I_53263 (I908011,I907994,I646333);
nor I_53264 (I907624,I907960,I908011);
nor I_53265 (I908042,I907994,I646345);
and I_53266 (I908059,I908042,I646348);
or I_53267 (I908076,I908059,I646327);
DFFARX1 I_53268 (I908076,I2507,I907632,I908102,);
nor I_53269 (I907612,I908102,I907658);
not I_53270 (I908124,I908102);
and I_53271 (I908141,I908124,I907658);
nor I_53272 (I907606,I907683,I908141);
nand I_53273 (I908172,I908124,I907734);
nor I_53274 (I907600,I907994,I908172);
nand I_53275 (I907603,I908124,I907912);
nand I_53276 (I908217,I907734,I646336);
nor I_53277 (I907615,I907977,I908217);
not I_53278 (I908278,I2514);
DFFARX1 I_53279 (I1066480,I2507,I908278,I908304,);
DFFARX1 I_53280 (I1066462,I2507,I908278,I908321,);
not I_53281 (I908329,I908321);
not I_53282 (I908346,I1066471);
nor I_53283 (I908363,I908346,I1066483);
not I_53284 (I908380,I1066465);
nor I_53285 (I908397,I908363,I1066474);
nor I_53286 (I908414,I908321,I908397);
DFFARX1 I_53287 (I908414,I2507,I908278,I908264,);
nor I_53288 (I908445,I1066474,I1066483);
nand I_53289 (I908462,I908445,I1066471);
DFFARX1 I_53290 (I908462,I2507,I908278,I908267,);
nor I_53291 (I908493,I908380,I1066474);
nand I_53292 (I908510,I908493,I1066486);
nor I_53293 (I908527,I908304,I908510);
DFFARX1 I_53294 (I908527,I2507,I908278,I908243,);
not I_53295 (I908558,I908510);
nand I_53296 (I908255,I908321,I908558);
DFFARX1 I_53297 (I908510,I2507,I908278,I908598,);
not I_53298 (I908606,I908598);
not I_53299 (I908623,I1066474);
not I_53300 (I908640,I1066462);
nor I_53301 (I908657,I908640,I1066465);
nor I_53302 (I908270,I908606,I908657);
nor I_53303 (I908688,I908640,I1066468);
and I_53304 (I908705,I908688,I1066477);
or I_53305 (I908722,I908705,I1066465);
DFFARX1 I_53306 (I908722,I2507,I908278,I908748,);
nor I_53307 (I908258,I908748,I908304);
not I_53308 (I908770,I908748);
and I_53309 (I908787,I908770,I908304);
nor I_53310 (I908252,I908329,I908787);
nand I_53311 (I908818,I908770,I908380);
nor I_53312 (I908246,I908640,I908818);
nand I_53313 (I908249,I908770,I908558);
nand I_53314 (I908863,I908380,I1066462);
nor I_53315 (I908261,I908623,I908863);
not I_53316 (I908924,I2514);
DFFARX1 I_53317 (I255460,I2507,I908924,I908950,);
DFFARX1 I_53318 (I255466,I2507,I908924,I908967,);
not I_53319 (I908975,I908967);
not I_53320 (I908992,I255487);
nor I_53321 (I909009,I908992,I255475);
not I_53322 (I909026,I255484);
nor I_53323 (I909043,I909009,I255469);
nor I_53324 (I909060,I908967,I909043);
DFFARX1 I_53325 (I909060,I2507,I908924,I908910,);
nor I_53326 (I909091,I255469,I255475);
nand I_53327 (I909108,I909091,I255487);
DFFARX1 I_53328 (I909108,I2507,I908924,I908913,);
nor I_53329 (I909139,I909026,I255469);
nand I_53330 (I909156,I909139,I255460);
nor I_53331 (I909173,I908950,I909156);
DFFARX1 I_53332 (I909173,I2507,I908924,I908889,);
not I_53333 (I909204,I909156);
nand I_53334 (I908901,I908967,I909204);
DFFARX1 I_53335 (I909156,I2507,I908924,I909244,);
not I_53336 (I909252,I909244);
not I_53337 (I909269,I255469);
not I_53338 (I909286,I255472);
nor I_53339 (I909303,I909286,I255484);
nor I_53340 (I908916,I909252,I909303);
nor I_53341 (I909334,I909286,I255481);
and I_53342 (I909351,I909334,I255463);
or I_53343 (I909368,I909351,I255478);
DFFARX1 I_53344 (I909368,I2507,I908924,I909394,);
nor I_53345 (I908904,I909394,I908950);
not I_53346 (I909416,I909394);
and I_53347 (I909433,I909416,I908950);
nor I_53348 (I908898,I908975,I909433);
nand I_53349 (I909464,I909416,I909026);
nor I_53350 (I908892,I909286,I909464);
nand I_53351 (I908895,I909416,I909204);
nand I_53352 (I909509,I909026,I255472);
nor I_53353 (I908907,I909269,I909509);
not I_53354 (I909570,I2514);
DFFARX1 I_53355 (I1318997,I2507,I909570,I909596,);
DFFARX1 I_53356 (I1319021,I2507,I909570,I909613,);
not I_53357 (I909621,I909613);
not I_53358 (I909638,I1319003);
nor I_53359 (I909655,I909638,I1319012);
not I_53360 (I909672,I1318997);
nor I_53361 (I909689,I909655,I1319018);
nor I_53362 (I909706,I909613,I909689);
DFFARX1 I_53363 (I909706,I2507,I909570,I909556,);
nor I_53364 (I909737,I1319018,I1319012);
nand I_53365 (I909754,I909737,I1319003);
DFFARX1 I_53366 (I909754,I2507,I909570,I909559,);
nor I_53367 (I909785,I909672,I1319018);
nand I_53368 (I909802,I909785,I1319015);
nor I_53369 (I909819,I909596,I909802);
DFFARX1 I_53370 (I909819,I2507,I909570,I909535,);
not I_53371 (I909850,I909802);
nand I_53372 (I909547,I909613,I909850);
DFFARX1 I_53373 (I909802,I2507,I909570,I909890,);
not I_53374 (I909898,I909890);
not I_53375 (I909915,I1319018);
not I_53376 (I909932,I1319009);
nor I_53377 (I909949,I909932,I1318997);
nor I_53378 (I909562,I909898,I909949);
nor I_53379 (I909980,I909932,I1319000);
and I_53380 (I909997,I909980,I1319024);
or I_53381 (I910014,I909997,I1319006);
DFFARX1 I_53382 (I910014,I2507,I909570,I910040,);
nor I_53383 (I909550,I910040,I909596);
not I_53384 (I910062,I910040);
and I_53385 (I910079,I910062,I909596);
nor I_53386 (I909544,I909621,I910079);
nand I_53387 (I910110,I910062,I909672);
nor I_53388 (I909538,I909932,I910110);
nand I_53389 (I909541,I910062,I909850);
nand I_53390 (I910155,I909672,I1319009);
nor I_53391 (I909553,I909915,I910155);
not I_53392 (I910216,I2514);
DFFARX1 I_53393 (I1023044,I2507,I910216,I910242,);
DFFARX1 I_53394 (I1023047,I2507,I910216,I910259,);
not I_53395 (I910267,I910259);
not I_53396 (I910284,I1023044);
nor I_53397 (I910301,I910284,I1023056);
not I_53398 (I910318,I1023065);
nor I_53399 (I910335,I910301,I1023053);
nor I_53400 (I910352,I910259,I910335);
DFFARX1 I_53401 (I910352,I2507,I910216,I910202,);
nor I_53402 (I910383,I1023053,I1023056);
nand I_53403 (I910400,I910383,I1023044);
DFFARX1 I_53404 (I910400,I2507,I910216,I910205,);
nor I_53405 (I910431,I910318,I1023053);
nand I_53406 (I910448,I910431,I1023059);
nor I_53407 (I910465,I910242,I910448);
DFFARX1 I_53408 (I910465,I2507,I910216,I910181,);
not I_53409 (I910496,I910448);
nand I_53410 (I910193,I910259,I910496);
DFFARX1 I_53411 (I910448,I2507,I910216,I910536,);
not I_53412 (I910544,I910536);
not I_53413 (I910561,I1023053);
not I_53414 (I910578,I1023050);
nor I_53415 (I910595,I910578,I1023065);
nor I_53416 (I910208,I910544,I910595);
nor I_53417 (I910626,I910578,I1023062);
and I_53418 (I910643,I910626,I1023050);
or I_53419 (I910660,I910643,I1023047);
DFFARX1 I_53420 (I910660,I2507,I910216,I910686,);
nor I_53421 (I910196,I910686,I910242);
not I_53422 (I910708,I910686);
and I_53423 (I910725,I910708,I910242);
nor I_53424 (I910190,I910267,I910725);
nand I_53425 (I910756,I910708,I910318);
nor I_53426 (I910184,I910578,I910756);
nand I_53427 (I910187,I910708,I910496);
nand I_53428 (I910801,I910318,I1023050);
nor I_53429 (I910199,I910561,I910801);
not I_53430 (I910862,I2514);
DFFARX1 I_53431 (I613959,I2507,I910862,I910888,);
DFFARX1 I_53432 (I613971,I2507,I910862,I910905,);
not I_53433 (I910913,I910905);
not I_53434 (I910930,I613980);
nor I_53435 (I910947,I910930,I613956);
not I_53436 (I910964,I613974);
nor I_53437 (I910981,I910947,I613968);
nor I_53438 (I910998,I910905,I910981);
DFFARX1 I_53439 (I910998,I2507,I910862,I910848,);
nor I_53440 (I911029,I613968,I613956);
nand I_53441 (I911046,I911029,I613980);
DFFARX1 I_53442 (I911046,I2507,I910862,I910851,);
nor I_53443 (I911077,I910964,I613968);
nand I_53444 (I911094,I911077,I613962);
nor I_53445 (I911111,I910888,I911094);
DFFARX1 I_53446 (I911111,I2507,I910862,I910827,);
not I_53447 (I911142,I911094);
nand I_53448 (I910839,I910905,I911142);
DFFARX1 I_53449 (I911094,I2507,I910862,I911182,);
not I_53450 (I911190,I911182);
not I_53451 (I911207,I613968);
not I_53452 (I911224,I613977);
nor I_53453 (I911241,I911224,I613974);
nor I_53454 (I910854,I911190,I911241);
nor I_53455 (I911272,I911224,I613959);
and I_53456 (I911289,I911272,I613956);
or I_53457 (I911306,I911289,I613965);
DFFARX1 I_53458 (I911306,I2507,I910862,I911332,);
nor I_53459 (I910842,I911332,I910888);
not I_53460 (I911354,I911332);
and I_53461 (I911371,I911354,I910888);
nor I_53462 (I910836,I910913,I911371);
nand I_53463 (I911402,I911354,I910964);
nor I_53464 (I910830,I911224,I911402);
nand I_53465 (I910833,I911354,I911142);
nand I_53466 (I911447,I910964,I613977);
nor I_53467 (I910845,I911207,I911447);
not I_53468 (I911508,I2514);
DFFARX1 I_53469 (I74886,I2507,I911508,I911534,);
DFFARX1 I_53470 (I74892,I2507,I911508,I911551,);
not I_53471 (I911559,I911551);
not I_53472 (I911576,I74910);
nor I_53473 (I911593,I911576,I74889);
not I_53474 (I911610,I74895);
nor I_53475 (I911627,I911593,I74901);
nor I_53476 (I911644,I911551,I911627);
DFFARX1 I_53477 (I911644,I2507,I911508,I911494,);
nor I_53478 (I911675,I74901,I74889);
nand I_53479 (I911692,I911675,I74910);
DFFARX1 I_53480 (I911692,I2507,I911508,I911497,);
nor I_53481 (I911723,I911610,I74901);
nand I_53482 (I911740,I911723,I74907);
nor I_53483 (I911757,I911534,I911740);
DFFARX1 I_53484 (I911757,I2507,I911508,I911473,);
not I_53485 (I911788,I911740);
nand I_53486 (I911485,I911551,I911788);
DFFARX1 I_53487 (I911740,I2507,I911508,I911828,);
not I_53488 (I911836,I911828);
not I_53489 (I911853,I74901);
not I_53490 (I911870,I74889);
nor I_53491 (I911887,I911870,I74895);
nor I_53492 (I911500,I911836,I911887);
nor I_53493 (I911918,I911870,I74898);
and I_53494 (I911935,I911918,I74886);
or I_53495 (I911952,I911935,I74904);
DFFARX1 I_53496 (I911952,I2507,I911508,I911978,);
nor I_53497 (I911488,I911978,I911534);
not I_53498 (I912000,I911978);
and I_53499 (I912017,I912000,I911534);
nor I_53500 (I911482,I911559,I912017);
nand I_53501 (I912048,I912000,I911610);
nor I_53502 (I911476,I911870,I912048);
nand I_53503 (I911479,I912000,I911788);
nand I_53504 (I912093,I911610,I74889);
nor I_53505 (I911491,I911853,I912093);
not I_53506 (I912154,I2514);
DFFARX1 I_53507 (I289715,I2507,I912154,I912180,);
DFFARX1 I_53508 (I289721,I2507,I912154,I912197,);
not I_53509 (I912205,I912197);
not I_53510 (I912222,I289742);
nor I_53511 (I912239,I912222,I289730);
not I_53512 (I912256,I289739);
nor I_53513 (I912273,I912239,I289724);
nor I_53514 (I912290,I912197,I912273);
DFFARX1 I_53515 (I912290,I2507,I912154,I912140,);
nor I_53516 (I912321,I289724,I289730);
nand I_53517 (I912338,I912321,I289742);
DFFARX1 I_53518 (I912338,I2507,I912154,I912143,);
nor I_53519 (I912369,I912256,I289724);
nand I_53520 (I912386,I912369,I289715);
nor I_53521 (I912403,I912180,I912386);
DFFARX1 I_53522 (I912403,I2507,I912154,I912119,);
not I_53523 (I912434,I912386);
nand I_53524 (I912131,I912197,I912434);
DFFARX1 I_53525 (I912386,I2507,I912154,I912474,);
not I_53526 (I912482,I912474);
not I_53527 (I912499,I289724);
not I_53528 (I912516,I289727);
nor I_53529 (I912533,I912516,I289739);
nor I_53530 (I912146,I912482,I912533);
nor I_53531 (I912564,I912516,I289736);
and I_53532 (I912581,I912564,I289718);
or I_53533 (I912598,I912581,I289733);
DFFARX1 I_53534 (I912598,I2507,I912154,I912624,);
nor I_53535 (I912134,I912624,I912180);
not I_53536 (I912646,I912624);
and I_53537 (I912663,I912646,I912180);
nor I_53538 (I912128,I912205,I912663);
nand I_53539 (I912694,I912646,I912256);
nor I_53540 (I912122,I912516,I912694);
nand I_53541 (I912125,I912646,I912434);
nand I_53542 (I912739,I912256,I289727);
nor I_53543 (I912137,I912499,I912739);
not I_53544 (I912800,I2514);
DFFARX1 I_53545 (I108087,I2507,I912800,I912826,);
DFFARX1 I_53546 (I108093,I2507,I912800,I912843,);
not I_53547 (I912851,I912843);
not I_53548 (I912868,I108111);
nor I_53549 (I912885,I912868,I108090);
not I_53550 (I912902,I108096);
nor I_53551 (I912919,I912885,I108102);
nor I_53552 (I912936,I912843,I912919);
DFFARX1 I_53553 (I912936,I2507,I912800,I912786,);
nor I_53554 (I912967,I108102,I108090);
nand I_53555 (I912984,I912967,I108111);
DFFARX1 I_53556 (I912984,I2507,I912800,I912789,);
nor I_53557 (I913015,I912902,I108102);
nand I_53558 (I913032,I913015,I108108);
nor I_53559 (I913049,I912826,I913032);
DFFARX1 I_53560 (I913049,I2507,I912800,I912765,);
not I_53561 (I913080,I913032);
nand I_53562 (I912777,I912843,I913080);
DFFARX1 I_53563 (I913032,I2507,I912800,I913120,);
not I_53564 (I913128,I913120);
not I_53565 (I913145,I108102);
not I_53566 (I913162,I108090);
nor I_53567 (I913179,I913162,I108096);
nor I_53568 (I912792,I913128,I913179);
nor I_53569 (I913210,I913162,I108099);
and I_53570 (I913227,I913210,I108087);
or I_53571 (I913244,I913227,I108105);
DFFARX1 I_53572 (I913244,I2507,I912800,I913270,);
nor I_53573 (I912780,I913270,I912826);
not I_53574 (I913292,I913270);
and I_53575 (I913309,I913292,I912826);
nor I_53576 (I912774,I912851,I913309);
nand I_53577 (I913340,I913292,I912902);
nor I_53578 (I912768,I913162,I913340);
nand I_53579 (I912771,I913292,I913080);
nand I_53580 (I913385,I912902,I108090);
nor I_53581 (I912783,I913145,I913385);
not I_53582 (I913446,I2514);
DFFARX1 I_53583 (I789079,I2507,I913446,I913472,);
DFFARX1 I_53584 (I789076,I2507,I913446,I913489,);
not I_53585 (I913497,I913489);
not I_53586 (I913514,I789076);
nor I_53587 (I913531,I913514,I789079);
not I_53588 (I913548,I789091);
nor I_53589 (I913565,I913531,I789085);
nor I_53590 (I913582,I913489,I913565);
DFFARX1 I_53591 (I913582,I2507,I913446,I913432,);
nor I_53592 (I913613,I789085,I789079);
nand I_53593 (I913630,I913613,I789076);
DFFARX1 I_53594 (I913630,I2507,I913446,I913435,);
nor I_53595 (I913661,I913548,I789085);
nand I_53596 (I913678,I913661,I789073);
nor I_53597 (I913695,I913472,I913678);
DFFARX1 I_53598 (I913695,I2507,I913446,I913411,);
not I_53599 (I913726,I913678);
nand I_53600 (I913423,I913489,I913726);
DFFARX1 I_53601 (I913678,I2507,I913446,I913766,);
not I_53602 (I913774,I913766);
not I_53603 (I913791,I789085);
not I_53604 (I913808,I789082);
nor I_53605 (I913825,I913808,I789091);
nor I_53606 (I913438,I913774,I913825);
nor I_53607 (I913856,I913808,I789088);
and I_53608 (I913873,I913856,I789094);
or I_53609 (I913890,I913873,I789073);
DFFARX1 I_53610 (I913890,I2507,I913446,I913916,);
nor I_53611 (I913426,I913916,I913472);
not I_53612 (I913938,I913916);
and I_53613 (I913955,I913938,I913472);
nor I_53614 (I913420,I913497,I913955);
nand I_53615 (I913986,I913938,I913548);
nor I_53616 (I913414,I913808,I913986);
nand I_53617 (I913417,I913938,I913726);
nand I_53618 (I914031,I913548,I789082);
nor I_53619 (I913429,I913791,I914031);
not I_53620 (I914092,I2514);
DFFARX1 I_53621 (I281283,I2507,I914092,I914118,);
DFFARX1 I_53622 (I281289,I2507,I914092,I914135,);
not I_53623 (I914143,I914135);
not I_53624 (I914160,I281310);
nor I_53625 (I914177,I914160,I281298);
not I_53626 (I914194,I281307);
nor I_53627 (I914211,I914177,I281292);
nor I_53628 (I914228,I914135,I914211);
DFFARX1 I_53629 (I914228,I2507,I914092,I914078,);
nor I_53630 (I914259,I281292,I281298);
nand I_53631 (I914276,I914259,I281310);
DFFARX1 I_53632 (I914276,I2507,I914092,I914081,);
nor I_53633 (I914307,I914194,I281292);
nand I_53634 (I914324,I914307,I281283);
nor I_53635 (I914341,I914118,I914324);
DFFARX1 I_53636 (I914341,I2507,I914092,I914057,);
not I_53637 (I914372,I914324);
nand I_53638 (I914069,I914135,I914372);
DFFARX1 I_53639 (I914324,I2507,I914092,I914412,);
not I_53640 (I914420,I914412);
not I_53641 (I914437,I281292);
not I_53642 (I914454,I281295);
nor I_53643 (I914471,I914454,I281307);
nor I_53644 (I914084,I914420,I914471);
nor I_53645 (I914502,I914454,I281304);
and I_53646 (I914519,I914502,I281286);
or I_53647 (I914536,I914519,I281301);
DFFARX1 I_53648 (I914536,I2507,I914092,I914562,);
nor I_53649 (I914072,I914562,I914118);
not I_53650 (I914584,I914562);
and I_53651 (I914601,I914584,I914118);
nor I_53652 (I914066,I914143,I914601);
nand I_53653 (I914632,I914584,I914194);
nor I_53654 (I914060,I914454,I914632);
nand I_53655 (I914063,I914584,I914372);
nand I_53656 (I914677,I914194,I281295);
nor I_53657 (I914075,I914437,I914677);
not I_53658 (I914738,I2514);
DFFARX1 I_53659 (I50644,I2507,I914738,I914764,);
DFFARX1 I_53660 (I50650,I2507,I914738,I914781,);
not I_53661 (I914789,I914781);
not I_53662 (I914806,I50668);
nor I_53663 (I914823,I914806,I50647);
not I_53664 (I914840,I50653);
nor I_53665 (I914857,I914823,I50659);
nor I_53666 (I914874,I914781,I914857);
DFFARX1 I_53667 (I914874,I2507,I914738,I914724,);
nor I_53668 (I914905,I50659,I50647);
nand I_53669 (I914922,I914905,I50668);
DFFARX1 I_53670 (I914922,I2507,I914738,I914727,);
nor I_53671 (I914953,I914840,I50659);
nand I_53672 (I914970,I914953,I50665);
nor I_53673 (I914987,I914764,I914970);
DFFARX1 I_53674 (I914987,I2507,I914738,I914703,);
not I_53675 (I915018,I914970);
nand I_53676 (I914715,I914781,I915018);
DFFARX1 I_53677 (I914970,I2507,I914738,I915058,);
not I_53678 (I915066,I915058);
not I_53679 (I915083,I50659);
not I_53680 (I915100,I50647);
nor I_53681 (I915117,I915100,I50653);
nor I_53682 (I914730,I915066,I915117);
nor I_53683 (I915148,I915100,I50656);
and I_53684 (I915165,I915148,I50644);
or I_53685 (I915182,I915165,I50662);
DFFARX1 I_53686 (I915182,I2507,I914738,I915208,);
nor I_53687 (I914718,I915208,I914764);
not I_53688 (I915230,I915208);
and I_53689 (I915247,I915230,I914764);
nor I_53690 (I914712,I914789,I915247);
nand I_53691 (I915278,I915230,I914840);
nor I_53692 (I914706,I915100,I915278);
nand I_53693 (I914709,I915230,I915018);
nand I_53694 (I915323,I914840,I50647);
nor I_53695 (I914721,I915083,I915323);
not I_53696 (I915384,I2514);
DFFARX1 I_53697 (I221041,I2507,I915384,I915410,);
DFFARX1 I_53698 (I221053,I2507,I915384,I915427,);
not I_53699 (I915435,I915427);
not I_53700 (I915452,I221059);
nor I_53701 (I915469,I915452,I221044);
not I_53702 (I915486,I221035);
nor I_53703 (I915503,I915469,I221056);
nor I_53704 (I915520,I915427,I915503);
DFFARX1 I_53705 (I915520,I2507,I915384,I915370,);
nor I_53706 (I915551,I221056,I221044);
nand I_53707 (I915568,I915551,I221059);
DFFARX1 I_53708 (I915568,I2507,I915384,I915373,);
nor I_53709 (I915599,I915486,I221056);
nand I_53710 (I915616,I915599,I221038);
nor I_53711 (I915633,I915410,I915616);
DFFARX1 I_53712 (I915633,I2507,I915384,I915349,);
not I_53713 (I915664,I915616);
nand I_53714 (I915361,I915427,I915664);
DFFARX1 I_53715 (I915616,I2507,I915384,I915704,);
not I_53716 (I915712,I915704);
not I_53717 (I915729,I221056);
not I_53718 (I915746,I221047);
nor I_53719 (I915763,I915746,I221035);
nor I_53720 (I915376,I915712,I915763);
nor I_53721 (I915794,I915746,I221050);
and I_53722 (I915811,I915794,I221038);
or I_53723 (I915828,I915811,I221035);
DFFARX1 I_53724 (I915828,I2507,I915384,I915854,);
nor I_53725 (I915364,I915854,I915410);
not I_53726 (I915876,I915854);
and I_53727 (I915893,I915876,I915410);
nor I_53728 (I915358,I915435,I915893);
nand I_53729 (I915924,I915876,I915486);
nor I_53730 (I915352,I915746,I915924);
nand I_53731 (I915355,I915876,I915664);
nand I_53732 (I915969,I915486,I221047);
nor I_53733 (I915367,I915729,I915969);
not I_53734 (I916030,I2514);
DFFARX1 I_53735 (I571187,I2507,I916030,I916056,);
DFFARX1 I_53736 (I571199,I2507,I916030,I916073,);
not I_53737 (I916081,I916073);
not I_53738 (I916098,I571208);
nor I_53739 (I916115,I916098,I571184);
not I_53740 (I916132,I571202);
nor I_53741 (I916149,I916115,I571196);
nor I_53742 (I916166,I916073,I916149);
DFFARX1 I_53743 (I916166,I2507,I916030,I916016,);
nor I_53744 (I916197,I571196,I571184);
nand I_53745 (I916214,I916197,I571208);
DFFARX1 I_53746 (I916214,I2507,I916030,I916019,);
nor I_53747 (I916245,I916132,I571196);
nand I_53748 (I916262,I916245,I571190);
nor I_53749 (I916279,I916056,I916262);
DFFARX1 I_53750 (I916279,I2507,I916030,I915995,);
not I_53751 (I916310,I916262);
nand I_53752 (I916007,I916073,I916310);
DFFARX1 I_53753 (I916262,I2507,I916030,I916350,);
not I_53754 (I916358,I916350);
not I_53755 (I916375,I571196);
not I_53756 (I916392,I571205);
nor I_53757 (I916409,I916392,I571202);
nor I_53758 (I916022,I916358,I916409);
nor I_53759 (I916440,I916392,I571187);
and I_53760 (I916457,I916440,I571184);
or I_53761 (I916474,I916457,I571193);
DFFARX1 I_53762 (I916474,I2507,I916030,I916500,);
nor I_53763 (I916010,I916500,I916056);
not I_53764 (I916522,I916500);
and I_53765 (I916539,I916522,I916056);
nor I_53766 (I916004,I916081,I916539);
nand I_53767 (I916570,I916522,I916132);
nor I_53768 (I915998,I916392,I916570);
nand I_53769 (I916001,I916522,I916310);
nand I_53770 (I916615,I916132,I571205);
nor I_53771 (I916013,I916375,I916615);
not I_53772 (I916676,I2514);
DFFARX1 I_53773 (I739966,I2507,I916676,I916702,);
DFFARX1 I_53774 (I739960,I2507,I916676,I916719,);
not I_53775 (I916727,I916719);
not I_53776 (I916744,I739975);
nor I_53777 (I916761,I916744,I739960);
not I_53778 (I916778,I739969);
nor I_53779 (I916795,I916761,I739978);
nor I_53780 (I916812,I916719,I916795);
DFFARX1 I_53781 (I916812,I2507,I916676,I916662,);
nor I_53782 (I916843,I739978,I739960);
nand I_53783 (I916860,I916843,I739975);
DFFARX1 I_53784 (I916860,I2507,I916676,I916665,);
nor I_53785 (I916891,I916778,I739978);
nand I_53786 (I916908,I916891,I739963);
nor I_53787 (I916925,I916702,I916908);
DFFARX1 I_53788 (I916925,I2507,I916676,I916641,);
not I_53789 (I916956,I916908);
nand I_53790 (I916653,I916719,I916956);
DFFARX1 I_53791 (I916908,I2507,I916676,I916996,);
not I_53792 (I917004,I916996);
not I_53793 (I917021,I739978);
not I_53794 (I917038,I739972);
nor I_53795 (I917055,I917038,I739969);
nor I_53796 (I916668,I917004,I917055);
nor I_53797 (I917086,I917038,I739981);
and I_53798 (I917103,I917086,I739984);
or I_53799 (I917120,I917103,I739963);
DFFARX1 I_53800 (I917120,I2507,I916676,I917146,);
nor I_53801 (I916656,I917146,I916702);
not I_53802 (I917168,I917146);
and I_53803 (I917185,I917168,I916702);
nor I_53804 (I916650,I916727,I917185);
nand I_53805 (I917216,I917168,I916778);
nor I_53806 (I916644,I917038,I917216);
nand I_53807 (I916647,I917168,I916956);
nand I_53808 (I917261,I916778,I739972);
nor I_53809 (I916659,I917021,I917261);
not I_53810 (I917322,I2514);
DFFARX1 I_53811 (I61184,I2507,I917322,I917348,);
DFFARX1 I_53812 (I61190,I2507,I917322,I917365,);
not I_53813 (I917373,I917365);
not I_53814 (I917390,I61208);
nor I_53815 (I917407,I917390,I61187);
not I_53816 (I917424,I61193);
nor I_53817 (I917441,I917407,I61199);
nor I_53818 (I917458,I917365,I917441);
DFFARX1 I_53819 (I917458,I2507,I917322,I917308,);
nor I_53820 (I917489,I61199,I61187);
nand I_53821 (I917506,I917489,I61208);
DFFARX1 I_53822 (I917506,I2507,I917322,I917311,);
nor I_53823 (I917537,I917424,I61199);
nand I_53824 (I917554,I917537,I61205);
nor I_53825 (I917571,I917348,I917554);
DFFARX1 I_53826 (I917571,I2507,I917322,I917287,);
not I_53827 (I917602,I917554);
nand I_53828 (I917299,I917365,I917602);
DFFARX1 I_53829 (I917554,I2507,I917322,I917642,);
not I_53830 (I917650,I917642);
not I_53831 (I917667,I61199);
not I_53832 (I917684,I61187);
nor I_53833 (I917701,I917684,I61193);
nor I_53834 (I917314,I917650,I917701);
nor I_53835 (I917732,I917684,I61196);
and I_53836 (I917749,I917732,I61184);
or I_53837 (I917766,I917749,I61202);
DFFARX1 I_53838 (I917766,I2507,I917322,I917792,);
nor I_53839 (I917302,I917792,I917348);
not I_53840 (I917814,I917792);
and I_53841 (I917831,I917814,I917348);
nor I_53842 (I917296,I917373,I917831);
nand I_53843 (I917862,I917814,I917424);
nor I_53844 (I917290,I917684,I917862);
nand I_53845 (I917293,I917814,I917602);
nand I_53846 (I917907,I917424,I61187);
nor I_53847 (I917305,I917667,I917907);
not I_53848 (I917968,I2514);
DFFARX1 I_53849 (I226991,I2507,I917968,I917994,);
DFFARX1 I_53850 (I227003,I2507,I917968,I918011,);
not I_53851 (I918019,I918011);
not I_53852 (I918036,I227009);
nor I_53853 (I918053,I918036,I226994);
not I_53854 (I918070,I226985);
nor I_53855 (I918087,I918053,I227006);
nor I_53856 (I918104,I918011,I918087);
DFFARX1 I_53857 (I918104,I2507,I917968,I917954,);
nor I_53858 (I918135,I227006,I226994);
nand I_53859 (I918152,I918135,I227009);
DFFARX1 I_53860 (I918152,I2507,I917968,I917957,);
nor I_53861 (I918183,I918070,I227006);
nand I_53862 (I918200,I918183,I226988);
nor I_53863 (I918217,I917994,I918200);
DFFARX1 I_53864 (I918217,I2507,I917968,I917933,);
not I_53865 (I918248,I918200);
nand I_53866 (I917945,I918011,I918248);
DFFARX1 I_53867 (I918200,I2507,I917968,I918288,);
not I_53868 (I918296,I918288);
not I_53869 (I918313,I227006);
not I_53870 (I918330,I226997);
nor I_53871 (I918347,I918330,I226985);
nor I_53872 (I917960,I918296,I918347);
nor I_53873 (I918378,I918330,I227000);
and I_53874 (I918395,I918378,I226988);
or I_53875 (I918412,I918395,I226985);
DFFARX1 I_53876 (I918412,I2507,I917968,I918438,);
nor I_53877 (I917948,I918438,I917994);
not I_53878 (I918460,I918438);
and I_53879 (I918477,I918460,I917994);
nor I_53880 (I917942,I918019,I918477);
nand I_53881 (I918508,I918460,I918070);
nor I_53882 (I917936,I918330,I918508);
nand I_53883 (I917939,I918460,I918248);
nand I_53884 (I918553,I918070,I226997);
nor I_53885 (I917951,I918313,I918553);
not I_53886 (I918614,I2514);
DFFARX1 I_53887 (I427829,I2507,I918614,I918640,);
DFFARX1 I_53888 (I427826,I2507,I918614,I918657,);
not I_53889 (I918665,I918657);
not I_53890 (I918682,I427841);
nor I_53891 (I918699,I918682,I427844);
not I_53892 (I918716,I427832);
nor I_53893 (I918733,I918699,I427838);
nor I_53894 (I918750,I918657,I918733);
DFFARX1 I_53895 (I918750,I2507,I918614,I918600,);
nor I_53896 (I918781,I427838,I427844);
nand I_53897 (I918798,I918781,I427841);
DFFARX1 I_53898 (I918798,I2507,I918614,I918603,);
nor I_53899 (I918829,I918716,I427838);
nand I_53900 (I918846,I918829,I427850);
nor I_53901 (I918863,I918640,I918846);
DFFARX1 I_53902 (I918863,I2507,I918614,I918579,);
not I_53903 (I918894,I918846);
nand I_53904 (I918591,I918657,I918894);
DFFARX1 I_53905 (I918846,I2507,I918614,I918934,);
not I_53906 (I918942,I918934);
not I_53907 (I918959,I427838);
not I_53908 (I918976,I427823);
nor I_53909 (I918993,I918976,I427832);
nor I_53910 (I918606,I918942,I918993);
nor I_53911 (I919024,I918976,I427835);
and I_53912 (I919041,I919024,I427823);
or I_53913 (I919058,I919041,I427847);
DFFARX1 I_53914 (I919058,I2507,I918614,I919084,);
nor I_53915 (I918594,I919084,I918640);
not I_53916 (I919106,I919084);
and I_53917 (I919123,I919106,I918640);
nor I_53918 (I918588,I918665,I919123);
nand I_53919 (I919154,I919106,I918716);
nor I_53920 (I918582,I918976,I919154);
nand I_53921 (I918585,I919106,I918894);
nand I_53922 (I919199,I918716,I427823);
nor I_53923 (I918597,I918959,I919199);
not I_53924 (I919260,I2514);
DFFARX1 I_53925 (I1081508,I2507,I919260,I919286,);
DFFARX1 I_53926 (I1081490,I2507,I919260,I919303,);
not I_53927 (I919311,I919303);
not I_53928 (I919328,I1081499);
nor I_53929 (I919345,I919328,I1081511);
not I_53930 (I919362,I1081493);
nor I_53931 (I919379,I919345,I1081502);
nor I_53932 (I919396,I919303,I919379);
DFFARX1 I_53933 (I919396,I2507,I919260,I919246,);
nor I_53934 (I919427,I1081502,I1081511);
nand I_53935 (I919444,I919427,I1081499);
DFFARX1 I_53936 (I919444,I2507,I919260,I919249,);
nor I_53937 (I919475,I919362,I1081502);
nand I_53938 (I919492,I919475,I1081514);
nor I_53939 (I919509,I919286,I919492);
DFFARX1 I_53940 (I919509,I2507,I919260,I919225,);
not I_53941 (I919540,I919492);
nand I_53942 (I919237,I919303,I919540);
DFFARX1 I_53943 (I919492,I2507,I919260,I919580,);
not I_53944 (I919588,I919580);
not I_53945 (I919605,I1081502);
not I_53946 (I919622,I1081490);
nor I_53947 (I919639,I919622,I1081493);
nor I_53948 (I919252,I919588,I919639);
nor I_53949 (I919670,I919622,I1081496);
and I_53950 (I919687,I919670,I1081505);
or I_53951 (I919704,I919687,I1081493);
DFFARX1 I_53952 (I919704,I2507,I919260,I919730,);
nor I_53953 (I919240,I919730,I919286);
not I_53954 (I919752,I919730);
and I_53955 (I919769,I919752,I919286);
nor I_53956 (I919234,I919311,I919769);
nand I_53957 (I919800,I919752,I919362);
nor I_53958 (I919228,I919622,I919800);
nand I_53959 (I919231,I919752,I919540);
nand I_53960 (I919845,I919362,I1081490);
nor I_53961 (I919243,I919605,I919845);
not I_53962 (I919906,I2514);
DFFARX1 I_53963 (I691992,I2507,I919906,I919932,);
DFFARX1 I_53964 (I691986,I2507,I919906,I919949,);
not I_53965 (I919957,I919949);
not I_53966 (I919974,I692001);
nor I_53967 (I919991,I919974,I691986);
not I_53968 (I920008,I691995);
nor I_53969 (I920025,I919991,I692004);
nor I_53970 (I920042,I919949,I920025);
DFFARX1 I_53971 (I920042,I2507,I919906,I919892,);
nor I_53972 (I920073,I692004,I691986);
nand I_53973 (I920090,I920073,I692001);
DFFARX1 I_53974 (I920090,I2507,I919906,I919895,);
nor I_53975 (I920121,I920008,I692004);
nand I_53976 (I920138,I920121,I691989);
nor I_53977 (I920155,I919932,I920138);
DFFARX1 I_53978 (I920155,I2507,I919906,I919871,);
not I_53979 (I920186,I920138);
nand I_53980 (I919883,I919949,I920186);
DFFARX1 I_53981 (I920138,I2507,I919906,I920226,);
not I_53982 (I920234,I920226);
not I_53983 (I920251,I692004);
not I_53984 (I920268,I691998);
nor I_53985 (I920285,I920268,I691995);
nor I_53986 (I919898,I920234,I920285);
nor I_53987 (I920316,I920268,I692007);
and I_53988 (I920333,I920316,I692010);
or I_53989 (I920350,I920333,I691989);
DFFARX1 I_53990 (I920350,I2507,I919906,I920376,);
nor I_53991 (I919886,I920376,I919932);
not I_53992 (I920398,I920376);
and I_53993 (I920415,I920398,I919932);
nor I_53994 (I919880,I919957,I920415);
nand I_53995 (I920446,I920398,I920008);
nor I_53996 (I919874,I920268,I920446);
nand I_53997 (I919877,I920398,I920186);
nand I_53998 (I920491,I920008,I691998);
nor I_53999 (I919889,I920251,I920491);
not I_54000 (I920552,I2514);
DFFARX1 I_54001 (I717424,I2507,I920552,I920578,);
DFFARX1 I_54002 (I717418,I2507,I920552,I920595,);
not I_54003 (I920603,I920595);
not I_54004 (I920620,I717433);
nor I_54005 (I920637,I920620,I717418);
not I_54006 (I920654,I717427);
nor I_54007 (I920671,I920637,I717436);
nor I_54008 (I920688,I920595,I920671);
DFFARX1 I_54009 (I920688,I2507,I920552,I920538,);
nor I_54010 (I920719,I717436,I717418);
nand I_54011 (I920736,I920719,I717433);
DFFARX1 I_54012 (I920736,I2507,I920552,I920541,);
nor I_54013 (I920767,I920654,I717436);
nand I_54014 (I920784,I920767,I717421);
nor I_54015 (I920801,I920578,I920784);
DFFARX1 I_54016 (I920801,I2507,I920552,I920517,);
not I_54017 (I920832,I920784);
nand I_54018 (I920529,I920595,I920832);
DFFARX1 I_54019 (I920784,I2507,I920552,I920872,);
not I_54020 (I920880,I920872);
not I_54021 (I920897,I717436);
not I_54022 (I920914,I717430);
nor I_54023 (I920931,I920914,I717427);
nor I_54024 (I920544,I920880,I920931);
nor I_54025 (I920962,I920914,I717439);
and I_54026 (I920979,I920962,I717442);
or I_54027 (I920996,I920979,I717421);
DFFARX1 I_54028 (I920996,I2507,I920552,I921022,);
nor I_54029 (I920532,I921022,I920578);
not I_54030 (I921044,I921022);
and I_54031 (I921061,I921044,I920578);
nor I_54032 (I920526,I920603,I921061);
nand I_54033 (I921092,I921044,I920654);
nor I_54034 (I920520,I920914,I921092);
nand I_54035 (I920523,I921044,I920832);
nand I_54036 (I921137,I920654,I717430);
nor I_54037 (I920535,I920897,I921137);
not I_54038 (I921198,I2514);
DFFARX1 I_54039 (I253352,I2507,I921198,I921224,);
DFFARX1 I_54040 (I253358,I2507,I921198,I921241,);
not I_54041 (I921249,I921241);
not I_54042 (I921266,I253379);
nor I_54043 (I921283,I921266,I253367);
not I_54044 (I921300,I253376);
nor I_54045 (I921317,I921283,I253361);
nor I_54046 (I921334,I921241,I921317);
DFFARX1 I_54047 (I921334,I2507,I921198,I921184,);
nor I_54048 (I921365,I253361,I253367);
nand I_54049 (I921382,I921365,I253379);
DFFARX1 I_54050 (I921382,I2507,I921198,I921187,);
nor I_54051 (I921413,I921300,I253361);
nand I_54052 (I921430,I921413,I253352);
nor I_54053 (I921447,I921224,I921430);
DFFARX1 I_54054 (I921447,I2507,I921198,I921163,);
not I_54055 (I921478,I921430);
nand I_54056 (I921175,I921241,I921478);
DFFARX1 I_54057 (I921430,I2507,I921198,I921518,);
not I_54058 (I921526,I921518);
not I_54059 (I921543,I253361);
not I_54060 (I921560,I253364);
nor I_54061 (I921577,I921560,I253376);
nor I_54062 (I921190,I921526,I921577);
nor I_54063 (I921608,I921560,I253373);
and I_54064 (I921625,I921608,I253355);
or I_54065 (I921642,I921625,I253370);
DFFARX1 I_54066 (I921642,I2507,I921198,I921668,);
nor I_54067 (I921178,I921668,I921224);
not I_54068 (I921690,I921668);
and I_54069 (I921707,I921690,I921224);
nor I_54070 (I921172,I921249,I921707);
nand I_54071 (I921738,I921690,I921300);
nor I_54072 (I921166,I921560,I921738);
nand I_54073 (I921169,I921690,I921478);
nand I_54074 (I921783,I921300,I253364);
nor I_54075 (I921181,I921543,I921783);
not I_54076 (I921844,I2514);
DFFARX1 I_54077 (I297093,I2507,I921844,I921870,);
DFFARX1 I_54078 (I297099,I2507,I921844,I921887,);
not I_54079 (I921895,I921887);
not I_54080 (I921912,I297120);
nor I_54081 (I921929,I921912,I297108);
not I_54082 (I921946,I297117);
nor I_54083 (I921963,I921929,I297102);
nor I_54084 (I921980,I921887,I921963);
DFFARX1 I_54085 (I921980,I2507,I921844,I921830,);
nor I_54086 (I922011,I297102,I297108);
nand I_54087 (I922028,I922011,I297120);
DFFARX1 I_54088 (I922028,I2507,I921844,I921833,);
nor I_54089 (I922059,I921946,I297102);
nand I_54090 (I922076,I922059,I297093);
nor I_54091 (I922093,I921870,I922076);
DFFARX1 I_54092 (I922093,I2507,I921844,I921809,);
not I_54093 (I922124,I922076);
nand I_54094 (I921821,I921887,I922124);
DFFARX1 I_54095 (I922076,I2507,I921844,I922164,);
not I_54096 (I922172,I922164);
not I_54097 (I922189,I297102);
not I_54098 (I922206,I297105);
nor I_54099 (I922223,I922206,I297117);
nor I_54100 (I921836,I922172,I922223);
nor I_54101 (I922254,I922206,I297114);
and I_54102 (I922271,I922254,I297096);
or I_54103 (I922288,I922271,I297111);
DFFARX1 I_54104 (I922288,I2507,I921844,I922314,);
nor I_54105 (I921824,I922314,I921870);
not I_54106 (I922336,I922314);
and I_54107 (I922353,I922336,I921870);
nor I_54108 (I921818,I921895,I922353);
nand I_54109 (I922384,I922336,I921946);
nor I_54110 (I921812,I922206,I922384);
nand I_54111 (I921815,I922336,I922124);
nand I_54112 (I922429,I921946,I297105);
nor I_54113 (I921827,I922189,I922429);
not I_54114 (I922490,I2514);
DFFARX1 I_54115 (I1115610,I2507,I922490,I922516,);
DFFARX1 I_54116 (I1115592,I2507,I922490,I922533,);
not I_54117 (I922541,I922533);
not I_54118 (I922558,I1115601);
nor I_54119 (I922575,I922558,I1115613);
not I_54120 (I922592,I1115595);
nor I_54121 (I922609,I922575,I1115604);
nor I_54122 (I922626,I922533,I922609);
DFFARX1 I_54123 (I922626,I2507,I922490,I922476,);
nor I_54124 (I922657,I1115604,I1115613);
nand I_54125 (I922674,I922657,I1115601);
DFFARX1 I_54126 (I922674,I2507,I922490,I922479,);
nor I_54127 (I922705,I922592,I1115604);
nand I_54128 (I922722,I922705,I1115616);
nor I_54129 (I922739,I922516,I922722);
DFFARX1 I_54130 (I922739,I2507,I922490,I922455,);
not I_54131 (I922770,I922722);
nand I_54132 (I922467,I922533,I922770);
DFFARX1 I_54133 (I922722,I2507,I922490,I922810,);
not I_54134 (I922818,I922810);
not I_54135 (I922835,I1115604);
not I_54136 (I922852,I1115592);
nor I_54137 (I922869,I922852,I1115595);
nor I_54138 (I922482,I922818,I922869);
nor I_54139 (I922900,I922852,I1115598);
and I_54140 (I922917,I922900,I1115607);
or I_54141 (I922934,I922917,I1115595);
DFFARX1 I_54142 (I922934,I2507,I922490,I922960,);
nor I_54143 (I922470,I922960,I922516);
not I_54144 (I922982,I922960);
and I_54145 (I922999,I922982,I922516);
nor I_54146 (I922464,I922541,I922999);
nand I_54147 (I923030,I922982,I922592);
nor I_54148 (I922458,I922852,I923030);
nand I_54149 (I922461,I922982,I922770);
nand I_54150 (I923075,I922592,I1115592);
nor I_54151 (I922473,I922835,I923075);
not I_54152 (I923136,I2514);
DFFARX1 I_54153 (I1146244,I2507,I923136,I923162,);
DFFARX1 I_54154 (I1146226,I2507,I923136,I923179,);
not I_54155 (I923187,I923179);
not I_54156 (I923204,I1146235);
nor I_54157 (I923221,I923204,I1146247);
not I_54158 (I923238,I1146229);
nor I_54159 (I923255,I923221,I1146238);
nor I_54160 (I923272,I923179,I923255);
DFFARX1 I_54161 (I923272,I2507,I923136,I923122,);
nor I_54162 (I923303,I1146238,I1146247);
nand I_54163 (I923320,I923303,I1146235);
DFFARX1 I_54164 (I923320,I2507,I923136,I923125,);
nor I_54165 (I923351,I923238,I1146238);
nand I_54166 (I923368,I923351,I1146250);
nor I_54167 (I923385,I923162,I923368);
DFFARX1 I_54168 (I923385,I2507,I923136,I923101,);
not I_54169 (I923416,I923368);
nand I_54170 (I923113,I923179,I923416);
DFFARX1 I_54171 (I923368,I2507,I923136,I923456,);
not I_54172 (I923464,I923456);
not I_54173 (I923481,I1146238);
not I_54174 (I923498,I1146226);
nor I_54175 (I923515,I923498,I1146229);
nor I_54176 (I923128,I923464,I923515);
nor I_54177 (I923546,I923498,I1146232);
and I_54178 (I923563,I923546,I1146241);
or I_54179 (I923580,I923563,I1146229);
DFFARX1 I_54180 (I923580,I2507,I923136,I923606,);
nor I_54181 (I923116,I923606,I923162);
not I_54182 (I923628,I923606);
and I_54183 (I923645,I923628,I923162);
nor I_54184 (I923110,I923187,I923645);
nand I_54185 (I923676,I923628,I923238);
nor I_54186 (I923104,I923498,I923676);
nand I_54187 (I923107,I923628,I923416);
nand I_54188 (I923721,I923238,I1146226);
nor I_54189 (I923119,I923481,I923721);
not I_54190 (I923782,I2514);
DFFARX1 I_54191 (I283391,I2507,I923782,I923808,);
DFFARX1 I_54192 (I283397,I2507,I923782,I923825,);
not I_54193 (I923833,I923825);
not I_54194 (I923850,I283418);
nor I_54195 (I923867,I923850,I283406);
not I_54196 (I923884,I283415);
nor I_54197 (I923901,I923867,I283400);
nor I_54198 (I923918,I923825,I923901);
DFFARX1 I_54199 (I923918,I2507,I923782,I923768,);
nor I_54200 (I923949,I283400,I283406);
nand I_54201 (I923966,I923949,I283418);
DFFARX1 I_54202 (I923966,I2507,I923782,I923771,);
nor I_54203 (I923997,I923884,I283400);
nand I_54204 (I924014,I923997,I283391);
nor I_54205 (I924031,I923808,I924014);
DFFARX1 I_54206 (I924031,I2507,I923782,I923747,);
not I_54207 (I924062,I924014);
nand I_54208 (I923759,I923825,I924062);
DFFARX1 I_54209 (I924014,I2507,I923782,I924102,);
not I_54210 (I924110,I924102);
not I_54211 (I924127,I283400);
not I_54212 (I924144,I283403);
nor I_54213 (I924161,I924144,I283415);
nor I_54214 (I923774,I924110,I924161);
nor I_54215 (I924192,I924144,I283412);
and I_54216 (I924209,I924192,I283394);
or I_54217 (I924226,I924209,I283409);
DFFARX1 I_54218 (I924226,I2507,I923782,I924252,);
nor I_54219 (I923762,I924252,I923808);
not I_54220 (I924274,I924252);
and I_54221 (I924291,I924274,I923808);
nor I_54222 (I923756,I923833,I924291);
nand I_54223 (I924322,I924274,I923884);
nor I_54224 (I923750,I924144,I924322);
nand I_54225 (I923753,I924274,I924062);
nand I_54226 (I924367,I923884,I283403);
nor I_54227 (I923765,I924127,I924367);
not I_54228 (I924428,I2514);
DFFARX1 I_54229 (I174036,I2507,I924428,I924454,);
DFFARX1 I_54230 (I174048,I2507,I924428,I924471,);
not I_54231 (I924479,I924471);
not I_54232 (I924496,I174054);
nor I_54233 (I924513,I924496,I174039);
not I_54234 (I924530,I174030);
nor I_54235 (I924547,I924513,I174051);
nor I_54236 (I924564,I924471,I924547);
DFFARX1 I_54237 (I924564,I2507,I924428,I924414,);
nor I_54238 (I924595,I174051,I174039);
nand I_54239 (I924612,I924595,I174054);
DFFARX1 I_54240 (I924612,I2507,I924428,I924417,);
nor I_54241 (I924643,I924530,I174051);
nand I_54242 (I924660,I924643,I174033);
nor I_54243 (I924677,I924454,I924660);
DFFARX1 I_54244 (I924677,I2507,I924428,I924393,);
not I_54245 (I924708,I924660);
nand I_54246 (I924405,I924471,I924708);
DFFARX1 I_54247 (I924660,I2507,I924428,I924748,);
not I_54248 (I924756,I924748);
not I_54249 (I924773,I174051);
not I_54250 (I924790,I174042);
nor I_54251 (I924807,I924790,I174030);
nor I_54252 (I924420,I924756,I924807);
nor I_54253 (I924838,I924790,I174045);
and I_54254 (I924855,I924838,I174033);
or I_54255 (I924872,I924855,I174030);
DFFARX1 I_54256 (I924872,I2507,I924428,I924898,);
nor I_54257 (I924408,I924898,I924454);
not I_54258 (I924920,I924898);
and I_54259 (I924937,I924920,I924454);
nor I_54260 (I924402,I924479,I924937);
nand I_54261 (I924968,I924920,I924530);
nor I_54262 (I924396,I924790,I924968);
nand I_54263 (I924399,I924920,I924708);
nand I_54264 (I925013,I924530,I174042);
nor I_54265 (I924411,I924773,I925013);
not I_54266 (I925074,I2514);
DFFARX1 I_54267 (I292350,I2507,I925074,I925100,);
DFFARX1 I_54268 (I292356,I2507,I925074,I925117,);
not I_54269 (I925125,I925117);
not I_54270 (I925142,I292377);
nor I_54271 (I925159,I925142,I292365);
not I_54272 (I925176,I292374);
nor I_54273 (I925193,I925159,I292359);
nor I_54274 (I925210,I925117,I925193);
DFFARX1 I_54275 (I925210,I2507,I925074,I925060,);
nor I_54276 (I925241,I292359,I292365);
nand I_54277 (I925258,I925241,I292377);
DFFARX1 I_54278 (I925258,I2507,I925074,I925063,);
nor I_54279 (I925289,I925176,I292359);
nand I_54280 (I925306,I925289,I292350);
nor I_54281 (I925323,I925100,I925306);
DFFARX1 I_54282 (I925323,I2507,I925074,I925039,);
not I_54283 (I925354,I925306);
nand I_54284 (I925051,I925117,I925354);
DFFARX1 I_54285 (I925306,I2507,I925074,I925394,);
not I_54286 (I925402,I925394);
not I_54287 (I925419,I292359);
not I_54288 (I925436,I292362);
nor I_54289 (I925453,I925436,I292374);
nor I_54290 (I925066,I925402,I925453);
nor I_54291 (I925484,I925436,I292371);
and I_54292 (I925501,I925484,I292353);
or I_54293 (I925518,I925501,I292368);
DFFARX1 I_54294 (I925518,I2507,I925074,I925544,);
nor I_54295 (I925054,I925544,I925100);
not I_54296 (I925566,I925544);
and I_54297 (I925583,I925566,I925100);
nor I_54298 (I925048,I925125,I925583);
nand I_54299 (I925614,I925566,I925176);
nor I_54300 (I925042,I925436,I925614);
nand I_54301 (I925045,I925566,I925354);
nand I_54302 (I925659,I925176,I292362);
nor I_54303 (I925057,I925419,I925659);
not I_54304 (I925720,I2514);
DFFARX1 I_54305 (I403893,I2507,I925720,I925746,);
DFFARX1 I_54306 (I403890,I2507,I925720,I925763,);
not I_54307 (I925771,I925763);
not I_54308 (I925788,I403905);
nor I_54309 (I925805,I925788,I403908);
not I_54310 (I925822,I403896);
nor I_54311 (I925839,I925805,I403902);
nor I_54312 (I925856,I925763,I925839);
DFFARX1 I_54313 (I925856,I2507,I925720,I925706,);
nor I_54314 (I925887,I403902,I403908);
nand I_54315 (I925904,I925887,I403905);
DFFARX1 I_54316 (I925904,I2507,I925720,I925709,);
nor I_54317 (I925935,I925822,I403902);
nand I_54318 (I925952,I925935,I403914);
nor I_54319 (I925969,I925746,I925952);
DFFARX1 I_54320 (I925969,I2507,I925720,I925685,);
not I_54321 (I926000,I925952);
nand I_54322 (I925697,I925763,I926000);
DFFARX1 I_54323 (I925952,I2507,I925720,I926040,);
not I_54324 (I926048,I926040);
not I_54325 (I926065,I403902);
not I_54326 (I926082,I403887);
nor I_54327 (I926099,I926082,I403896);
nor I_54328 (I925712,I926048,I926099);
nor I_54329 (I926130,I926082,I403899);
and I_54330 (I926147,I926130,I403887);
or I_54331 (I926164,I926147,I403911);
DFFARX1 I_54332 (I926164,I2507,I925720,I926190,);
nor I_54333 (I925700,I926190,I925746);
not I_54334 (I926212,I926190);
and I_54335 (I926229,I926212,I925746);
nor I_54336 (I925694,I925771,I926229);
nand I_54337 (I926260,I926212,I925822);
nor I_54338 (I925688,I926082,I926260);
nand I_54339 (I925691,I926212,I926000);
nand I_54340 (I926305,I925822,I403887);
nor I_54341 (I925703,I926065,I926305);
not I_54342 (I926366,I2514);
DFFARX1 I_54343 (I130748,I2507,I926366,I926392,);
DFFARX1 I_54344 (I130754,I2507,I926366,I926409,);
not I_54345 (I926417,I926409);
not I_54346 (I926434,I130772);
nor I_54347 (I926451,I926434,I130751);
not I_54348 (I926468,I130757);
nor I_54349 (I926485,I926451,I130763);
nor I_54350 (I926502,I926409,I926485);
DFFARX1 I_54351 (I926502,I2507,I926366,I926352,);
nor I_54352 (I926533,I130763,I130751);
nand I_54353 (I926550,I926533,I130772);
DFFARX1 I_54354 (I926550,I2507,I926366,I926355,);
nor I_54355 (I926581,I926468,I130763);
nand I_54356 (I926598,I926581,I130769);
nor I_54357 (I926615,I926392,I926598);
DFFARX1 I_54358 (I926615,I2507,I926366,I926331,);
not I_54359 (I926646,I926598);
nand I_54360 (I926343,I926409,I926646);
DFFARX1 I_54361 (I926598,I2507,I926366,I926686,);
not I_54362 (I926694,I926686);
not I_54363 (I926711,I130763);
not I_54364 (I926728,I130751);
nor I_54365 (I926745,I926728,I130757);
nor I_54366 (I926358,I926694,I926745);
nor I_54367 (I926776,I926728,I130760);
and I_54368 (I926793,I926776,I130748);
or I_54369 (I926810,I926793,I130766);
DFFARX1 I_54370 (I926810,I2507,I926366,I926836,);
nor I_54371 (I926346,I926836,I926392);
not I_54372 (I926858,I926836);
and I_54373 (I926875,I926858,I926392);
nor I_54374 (I926340,I926417,I926875);
nand I_54375 (I926906,I926858,I926468);
nor I_54376 (I926334,I926728,I926906);
nand I_54377 (I926337,I926858,I926646);
nand I_54378 (I926951,I926468,I130751);
nor I_54379 (I926349,I926711,I926951);
not I_54380 (I927012,I2514);
DFFARX1 I_54381 (I1317212,I2507,I927012,I927038,);
DFFARX1 I_54382 (I1317236,I2507,I927012,I927055,);
not I_54383 (I927063,I927055);
not I_54384 (I927080,I1317218);
nor I_54385 (I927097,I927080,I1317227);
not I_54386 (I927114,I1317212);
nor I_54387 (I927131,I927097,I1317233);
nor I_54388 (I927148,I927055,I927131);
DFFARX1 I_54389 (I927148,I2507,I927012,I926998,);
nor I_54390 (I927179,I1317233,I1317227);
nand I_54391 (I927196,I927179,I1317218);
DFFARX1 I_54392 (I927196,I2507,I927012,I927001,);
nor I_54393 (I927227,I927114,I1317233);
nand I_54394 (I927244,I927227,I1317230);
nor I_54395 (I927261,I927038,I927244);
DFFARX1 I_54396 (I927261,I2507,I927012,I926977,);
not I_54397 (I927292,I927244);
nand I_54398 (I926989,I927055,I927292);
DFFARX1 I_54399 (I927244,I2507,I927012,I927332,);
not I_54400 (I927340,I927332);
not I_54401 (I927357,I1317233);
not I_54402 (I927374,I1317224);
nor I_54403 (I927391,I927374,I1317212);
nor I_54404 (I927004,I927340,I927391);
nor I_54405 (I927422,I927374,I1317215);
and I_54406 (I927439,I927422,I1317239);
or I_54407 (I927456,I927439,I1317221);
DFFARX1 I_54408 (I927456,I2507,I927012,I927482,);
nor I_54409 (I926992,I927482,I927038);
not I_54410 (I927504,I927482);
and I_54411 (I927521,I927504,I927038);
nor I_54412 (I926986,I927063,I927521);
nand I_54413 (I927552,I927504,I927114);
nor I_54414 (I926980,I927374,I927552);
nand I_54415 (I926983,I927504,I927292);
nand I_54416 (I927597,I927114,I1317224);
nor I_54417 (I926995,I927357,I927597);
not I_54418 (I927658,I2514);
DFFARX1 I_54419 (I1219956,I2507,I927658,I927684,);
DFFARX1 I_54420 (I1219962,I2507,I927658,I927701,);
not I_54421 (I927709,I927701);
not I_54422 (I927726,I1219959);
nor I_54423 (I927743,I927726,I1219938);
not I_54424 (I927760,I1219941);
nor I_54425 (I927777,I927743,I1219947);
nor I_54426 (I927794,I927701,I927777);
DFFARX1 I_54427 (I927794,I2507,I927658,I927644,);
nor I_54428 (I927825,I1219947,I1219938);
nand I_54429 (I927842,I927825,I1219959);
DFFARX1 I_54430 (I927842,I2507,I927658,I927647,);
nor I_54431 (I927873,I927760,I1219947);
nand I_54432 (I927890,I927873,I1219941);
nor I_54433 (I927907,I927684,I927890);
DFFARX1 I_54434 (I927907,I2507,I927658,I927623,);
not I_54435 (I927938,I927890);
nand I_54436 (I927635,I927701,I927938);
DFFARX1 I_54437 (I927890,I2507,I927658,I927978,);
not I_54438 (I927986,I927978);
not I_54439 (I928003,I1219947);
not I_54440 (I928020,I1219950);
nor I_54441 (I928037,I928020,I1219941);
nor I_54442 (I927650,I927986,I928037);
nor I_54443 (I928068,I928020,I1219938);
and I_54444 (I928085,I928068,I1219944);
or I_54445 (I928102,I928085,I1219953);
DFFARX1 I_54446 (I928102,I2507,I927658,I928128,);
nor I_54447 (I927638,I928128,I927684);
not I_54448 (I928150,I928128);
and I_54449 (I928167,I928150,I927684);
nor I_54450 (I927632,I927709,I928167);
nand I_54451 (I928198,I928150,I927760);
nor I_54452 (I927626,I928020,I928198);
nand I_54453 (I927629,I928150,I927938);
nand I_54454 (I928243,I927760,I1219950);
nor I_54455 (I927641,I928003,I928243);
not I_54456 (I928304,I2514);
DFFARX1 I_54457 (I823334,I2507,I928304,I928330,);
DFFARX1 I_54458 (I823331,I2507,I928304,I928347,);
not I_54459 (I928355,I928347);
not I_54460 (I928372,I823331);
nor I_54461 (I928389,I928372,I823334);
not I_54462 (I928406,I823346);
nor I_54463 (I928423,I928389,I823340);
nor I_54464 (I928440,I928347,I928423);
DFFARX1 I_54465 (I928440,I2507,I928304,I928290,);
nor I_54466 (I928471,I823340,I823334);
nand I_54467 (I928488,I928471,I823331);
DFFARX1 I_54468 (I928488,I2507,I928304,I928293,);
nor I_54469 (I928519,I928406,I823340);
nand I_54470 (I928536,I928519,I823328);
nor I_54471 (I928553,I928330,I928536);
DFFARX1 I_54472 (I928553,I2507,I928304,I928269,);
not I_54473 (I928584,I928536);
nand I_54474 (I928281,I928347,I928584);
DFFARX1 I_54475 (I928536,I2507,I928304,I928624,);
not I_54476 (I928632,I928624);
not I_54477 (I928649,I823340);
not I_54478 (I928666,I823337);
nor I_54479 (I928683,I928666,I823346);
nor I_54480 (I928296,I928632,I928683);
nor I_54481 (I928714,I928666,I823343);
and I_54482 (I928731,I928714,I823349);
or I_54483 (I928748,I928731,I823328);
DFFARX1 I_54484 (I928748,I2507,I928304,I928774,);
nor I_54485 (I928284,I928774,I928330);
not I_54486 (I928796,I928774);
and I_54487 (I928813,I928796,I928330);
nor I_54488 (I928278,I928355,I928813);
nand I_54489 (I928844,I928796,I928406);
nor I_54490 (I928272,I928666,I928844);
nand I_54491 (I928275,I928796,I928584);
nand I_54492 (I928889,I928406,I823337);
nor I_54493 (I928287,I928649,I928889);
not I_54494 (I928950,I2514);
DFFARX1 I_54495 (I1294645,I2507,I928950,I928976,);
DFFARX1 I_54496 (I1294639,I2507,I928950,I928993,);
not I_54497 (I929001,I928993);
not I_54498 (I929018,I1294648);
nor I_54499 (I929035,I929018,I1294660);
not I_54500 (I929052,I1294642);
nor I_54501 (I929069,I929035,I1294639);
nor I_54502 (I929086,I928993,I929069);
DFFARX1 I_54503 (I929086,I2507,I928950,I928936,);
nor I_54504 (I929117,I1294639,I1294660);
nand I_54505 (I929134,I929117,I1294648);
DFFARX1 I_54506 (I929134,I2507,I928950,I928939,);
nor I_54507 (I929165,I929052,I1294639);
nand I_54508 (I929182,I929165,I1294636);
nor I_54509 (I929199,I928976,I929182);
DFFARX1 I_54510 (I929199,I2507,I928950,I928915,);
not I_54511 (I929230,I929182);
nand I_54512 (I928927,I928993,I929230);
DFFARX1 I_54513 (I929182,I2507,I928950,I929270,);
not I_54514 (I929278,I929270);
not I_54515 (I929295,I1294639);
not I_54516 (I929312,I1294657);
nor I_54517 (I929329,I929312,I1294642);
nor I_54518 (I928942,I929278,I929329);
nor I_54519 (I929360,I929312,I1294651);
and I_54520 (I929377,I929360,I1294636);
or I_54521 (I929394,I929377,I1294654);
DFFARX1 I_54522 (I929394,I2507,I928950,I929420,);
nor I_54523 (I928930,I929420,I928976);
not I_54524 (I929442,I929420);
and I_54525 (I929459,I929442,I928976);
nor I_54526 (I928924,I929001,I929459);
nand I_54527 (I929490,I929442,I929052);
nor I_54528 (I928918,I929312,I929490);
nand I_54529 (I928921,I929442,I929230);
nand I_54530 (I929535,I929052,I1294657);
nor I_54531 (I928933,I929295,I929535);
not I_54532 (I929596,I2514);
DFFARX1 I_54533 (I164516,I2507,I929596,I929622,);
DFFARX1 I_54534 (I164528,I2507,I929596,I929639,);
not I_54535 (I929647,I929639);
not I_54536 (I929664,I164534);
nor I_54537 (I929681,I929664,I164519);
not I_54538 (I929698,I164510);
nor I_54539 (I929715,I929681,I164531);
nor I_54540 (I929732,I929639,I929715);
DFFARX1 I_54541 (I929732,I2507,I929596,I929582,);
nor I_54542 (I929763,I164531,I164519);
nand I_54543 (I929780,I929763,I164534);
DFFARX1 I_54544 (I929780,I2507,I929596,I929585,);
nor I_54545 (I929811,I929698,I164531);
nand I_54546 (I929828,I929811,I164513);
nor I_54547 (I929845,I929622,I929828);
DFFARX1 I_54548 (I929845,I2507,I929596,I929561,);
not I_54549 (I929876,I929828);
nand I_54550 (I929573,I929639,I929876);
DFFARX1 I_54551 (I929828,I2507,I929596,I929916,);
not I_54552 (I929924,I929916);
not I_54553 (I929941,I164531);
not I_54554 (I929958,I164522);
nor I_54555 (I929975,I929958,I164510);
nor I_54556 (I929588,I929924,I929975);
nor I_54557 (I930006,I929958,I164525);
and I_54558 (I930023,I930006,I164513);
or I_54559 (I930040,I930023,I164510);
DFFARX1 I_54560 (I930040,I2507,I929596,I930066,);
nor I_54561 (I929576,I930066,I929622);
not I_54562 (I930088,I930066);
and I_54563 (I930105,I930088,I929622);
nor I_54564 (I929570,I929647,I930105);
nand I_54565 (I930136,I930088,I929698);
nor I_54566 (I929564,I929958,I930136);
nand I_54567 (I929567,I930088,I929876);
nand I_54568 (I930181,I929698,I164522);
nor I_54569 (I929579,I929941,I930181);
not I_54570 (I930242,I2514);
DFFARX1 I_54571 (I165706,I2507,I930242,I930268,);
DFFARX1 I_54572 (I165718,I2507,I930242,I930285,);
not I_54573 (I930293,I930285);
not I_54574 (I930310,I165724);
nor I_54575 (I930327,I930310,I165709);
not I_54576 (I930344,I165700);
nor I_54577 (I930361,I930327,I165721);
nor I_54578 (I930378,I930285,I930361);
DFFARX1 I_54579 (I930378,I2507,I930242,I930228,);
nor I_54580 (I930409,I165721,I165709);
nand I_54581 (I930426,I930409,I165724);
DFFARX1 I_54582 (I930426,I2507,I930242,I930231,);
nor I_54583 (I930457,I930344,I165721);
nand I_54584 (I930474,I930457,I165703);
nor I_54585 (I930491,I930268,I930474);
DFFARX1 I_54586 (I930491,I2507,I930242,I930207,);
not I_54587 (I930522,I930474);
nand I_54588 (I930219,I930285,I930522);
DFFARX1 I_54589 (I930474,I2507,I930242,I930562,);
not I_54590 (I930570,I930562);
not I_54591 (I930587,I165721);
not I_54592 (I930604,I165712);
nor I_54593 (I930621,I930604,I165700);
nor I_54594 (I930234,I930570,I930621);
nor I_54595 (I930652,I930604,I165715);
and I_54596 (I930669,I930652,I165703);
or I_54597 (I930686,I930669,I165700);
DFFARX1 I_54598 (I930686,I2507,I930242,I930712,);
nor I_54599 (I930222,I930712,I930268);
not I_54600 (I930734,I930712);
and I_54601 (I930751,I930734,I930268);
nor I_54602 (I930216,I930293,I930751);
nand I_54603 (I930782,I930734,I930344);
nor I_54604 (I930210,I930604,I930782);
nand I_54605 (I930213,I930734,I930522);
nand I_54606 (I930827,I930344,I165712);
nor I_54607 (I930225,I930587,I930827);
not I_54608 (I930888,I2514);
DFFARX1 I_54609 (I500637,I2507,I930888,I930914,);
DFFARX1 I_54610 (I500649,I2507,I930888,I930931,);
not I_54611 (I930939,I930931);
not I_54612 (I930956,I500634);
nor I_54613 (I930973,I930956,I500652);
not I_54614 (I930990,I500658);
nor I_54615 (I931007,I930973,I500640);
nor I_54616 (I931024,I930931,I931007);
DFFARX1 I_54617 (I931024,I2507,I930888,I930874,);
nor I_54618 (I931055,I500640,I500652);
nand I_54619 (I931072,I931055,I500634);
DFFARX1 I_54620 (I931072,I2507,I930888,I930877,);
nor I_54621 (I931103,I930990,I500640);
nand I_54622 (I931120,I931103,I500643);
nor I_54623 (I931137,I930914,I931120);
DFFARX1 I_54624 (I931137,I2507,I930888,I930853,);
not I_54625 (I931168,I931120);
nand I_54626 (I930865,I930931,I931168);
DFFARX1 I_54627 (I931120,I2507,I930888,I931208,);
not I_54628 (I931216,I931208);
not I_54629 (I931233,I500640);
not I_54630 (I931250,I500646);
nor I_54631 (I931267,I931250,I500658);
nor I_54632 (I930880,I931216,I931267);
nor I_54633 (I931298,I931250,I500655);
and I_54634 (I931315,I931298,I500634);
or I_54635 (I931332,I931315,I500637);
DFFARX1 I_54636 (I931332,I2507,I930888,I931358,);
nor I_54637 (I930868,I931358,I930914);
not I_54638 (I931380,I931358);
and I_54639 (I931397,I931380,I930914);
nor I_54640 (I930862,I930939,I931397);
nand I_54641 (I931428,I931380,I930990);
nor I_54642 (I930856,I931250,I931428);
nand I_54643 (I930859,I931380,I931168);
nand I_54644 (I931473,I930990,I500646);
nor I_54645 (I930871,I931233,I931473);
not I_54646 (I931534,I2514);
DFFARX1 I_54647 (I622051,I2507,I931534,I931560,);
DFFARX1 I_54648 (I622063,I2507,I931534,I931577,);
not I_54649 (I931585,I931577);
not I_54650 (I931602,I622072);
nor I_54651 (I931619,I931602,I622048);
not I_54652 (I931636,I622066);
nor I_54653 (I931653,I931619,I622060);
nor I_54654 (I931670,I931577,I931653);
DFFARX1 I_54655 (I931670,I2507,I931534,I931520,);
nor I_54656 (I931701,I622060,I622048);
nand I_54657 (I931718,I931701,I622072);
DFFARX1 I_54658 (I931718,I2507,I931534,I931523,);
nor I_54659 (I931749,I931636,I622060);
nand I_54660 (I931766,I931749,I622054);
nor I_54661 (I931783,I931560,I931766);
DFFARX1 I_54662 (I931783,I2507,I931534,I931499,);
not I_54663 (I931814,I931766);
nand I_54664 (I931511,I931577,I931814);
DFFARX1 I_54665 (I931766,I2507,I931534,I931854,);
not I_54666 (I931862,I931854);
not I_54667 (I931879,I622060);
not I_54668 (I931896,I622069);
nor I_54669 (I931913,I931896,I622066);
nor I_54670 (I931526,I931862,I931913);
nor I_54671 (I931944,I931896,I622051);
and I_54672 (I931961,I931944,I622048);
or I_54673 (I931978,I931961,I622057);
DFFARX1 I_54674 (I931978,I2507,I931534,I932004,);
nor I_54675 (I931514,I932004,I931560);
not I_54676 (I932026,I932004);
and I_54677 (I932043,I932026,I931560);
nor I_54678 (I931508,I931585,I932043);
nand I_54679 (I932074,I932026,I931636);
nor I_54680 (I931502,I931896,I932074);
nand I_54681 (I931505,I932026,I931814);
nand I_54682 (I932119,I931636,I622069);
nor I_54683 (I931517,I931879,I932119);
not I_54684 (I932180,I2514);
DFFARX1 I_54685 (I1139308,I2507,I932180,I932206,);
DFFARX1 I_54686 (I1139290,I2507,I932180,I932223,);
not I_54687 (I932231,I932223);
not I_54688 (I932248,I1139299);
nor I_54689 (I932265,I932248,I1139311);
not I_54690 (I932282,I1139293);
nor I_54691 (I932299,I932265,I1139302);
nor I_54692 (I932316,I932223,I932299);
DFFARX1 I_54693 (I932316,I2507,I932180,I932166,);
nor I_54694 (I932347,I1139302,I1139311);
nand I_54695 (I932364,I932347,I1139299);
DFFARX1 I_54696 (I932364,I2507,I932180,I932169,);
nor I_54697 (I932395,I932282,I1139302);
nand I_54698 (I932412,I932395,I1139314);
nor I_54699 (I932429,I932206,I932412);
DFFARX1 I_54700 (I932429,I2507,I932180,I932145,);
not I_54701 (I932460,I932412);
nand I_54702 (I932157,I932223,I932460);
DFFARX1 I_54703 (I932412,I2507,I932180,I932500,);
not I_54704 (I932508,I932500);
not I_54705 (I932525,I1139302);
not I_54706 (I932542,I1139290);
nor I_54707 (I932559,I932542,I1139293);
nor I_54708 (I932172,I932508,I932559);
nor I_54709 (I932590,I932542,I1139296);
and I_54710 (I932607,I932590,I1139305);
or I_54711 (I932624,I932607,I1139293);
DFFARX1 I_54712 (I932624,I2507,I932180,I932650,);
nor I_54713 (I932160,I932650,I932206);
not I_54714 (I932672,I932650);
and I_54715 (I932689,I932672,I932206);
nor I_54716 (I932154,I932231,I932689);
nand I_54717 (I932720,I932672,I932282);
nor I_54718 (I932148,I932542,I932720);
nand I_54719 (I932151,I932672,I932460);
nand I_54720 (I932765,I932282,I1139290);
nor I_54721 (I932163,I932525,I932765);
not I_54722 (I932826,I2514);
DFFARX1 I_54723 (I591417,I2507,I932826,I932852,);
DFFARX1 I_54724 (I591429,I2507,I932826,I932869,);
not I_54725 (I932877,I932869);
not I_54726 (I932894,I591438);
nor I_54727 (I932911,I932894,I591414);
not I_54728 (I932928,I591432);
nor I_54729 (I932945,I932911,I591426);
nor I_54730 (I932962,I932869,I932945);
DFFARX1 I_54731 (I932962,I2507,I932826,I932812,);
nor I_54732 (I932993,I591426,I591414);
nand I_54733 (I933010,I932993,I591438);
DFFARX1 I_54734 (I933010,I2507,I932826,I932815,);
nor I_54735 (I933041,I932928,I591426);
nand I_54736 (I933058,I933041,I591420);
nor I_54737 (I933075,I932852,I933058);
DFFARX1 I_54738 (I933075,I2507,I932826,I932791,);
not I_54739 (I933106,I933058);
nand I_54740 (I932803,I932869,I933106);
DFFARX1 I_54741 (I933058,I2507,I932826,I933146,);
not I_54742 (I933154,I933146);
not I_54743 (I933171,I591426);
not I_54744 (I933188,I591435);
nor I_54745 (I933205,I933188,I591432);
nor I_54746 (I932818,I933154,I933205);
nor I_54747 (I933236,I933188,I591417);
and I_54748 (I933253,I933236,I591414);
or I_54749 (I933270,I933253,I591423);
DFFARX1 I_54750 (I933270,I2507,I932826,I933296,);
nor I_54751 (I932806,I933296,I932852);
not I_54752 (I933318,I933296);
and I_54753 (I933335,I933318,I932852);
nor I_54754 (I932800,I932877,I933335);
nand I_54755 (I933366,I933318,I932928);
nor I_54756 (I932794,I933188,I933366);
nand I_54757 (I932797,I933318,I933106);
nand I_54758 (I933411,I932928,I591435);
nor I_54759 (I932809,I933171,I933411);
not I_54760 (I933472,I2514);
DFFARX1 I_54761 (I575811,I2507,I933472,I933498,);
DFFARX1 I_54762 (I575823,I2507,I933472,I933515,);
not I_54763 (I933523,I933515);
not I_54764 (I933540,I575832);
nor I_54765 (I933557,I933540,I575808);
not I_54766 (I933574,I575826);
nor I_54767 (I933591,I933557,I575820);
nor I_54768 (I933608,I933515,I933591);
DFFARX1 I_54769 (I933608,I2507,I933472,I933458,);
nor I_54770 (I933639,I575820,I575808);
nand I_54771 (I933656,I933639,I575832);
DFFARX1 I_54772 (I933656,I2507,I933472,I933461,);
nor I_54773 (I933687,I933574,I575820);
nand I_54774 (I933704,I933687,I575814);
nor I_54775 (I933721,I933498,I933704);
DFFARX1 I_54776 (I933721,I2507,I933472,I933437,);
not I_54777 (I933752,I933704);
nand I_54778 (I933449,I933515,I933752);
DFFARX1 I_54779 (I933704,I2507,I933472,I933792,);
not I_54780 (I933800,I933792);
not I_54781 (I933817,I575820);
not I_54782 (I933834,I575829);
nor I_54783 (I933851,I933834,I575826);
nor I_54784 (I933464,I933800,I933851);
nor I_54785 (I933882,I933834,I575811);
and I_54786 (I933899,I933882,I575808);
or I_54787 (I933916,I933899,I575817);
DFFARX1 I_54788 (I933916,I2507,I933472,I933942,);
nor I_54789 (I933452,I933942,I933498);
not I_54790 (I933964,I933942);
and I_54791 (I933981,I933964,I933498);
nor I_54792 (I933446,I933523,I933981);
nand I_54793 (I934012,I933964,I933574);
nor I_54794 (I933440,I933834,I934012);
nand I_54795 (I933443,I933964,I933752);
nand I_54796 (I934057,I933574,I575829);
nor I_54797 (I933455,I933817,I934057);
not I_54798 (I934118,I2514);
DFFARX1 I_54799 (I1316617,I2507,I934118,I934144,);
DFFARX1 I_54800 (I1316641,I2507,I934118,I934161,);
not I_54801 (I934169,I934161);
not I_54802 (I934186,I1316623);
nor I_54803 (I934203,I934186,I1316632);
not I_54804 (I934220,I1316617);
nor I_54805 (I934237,I934203,I1316638);
nor I_54806 (I934254,I934161,I934237);
DFFARX1 I_54807 (I934254,I2507,I934118,I934104,);
nor I_54808 (I934285,I1316638,I1316632);
nand I_54809 (I934302,I934285,I1316623);
DFFARX1 I_54810 (I934302,I2507,I934118,I934107,);
nor I_54811 (I934333,I934220,I1316638);
nand I_54812 (I934350,I934333,I1316635);
nor I_54813 (I934367,I934144,I934350);
DFFARX1 I_54814 (I934367,I2507,I934118,I934083,);
not I_54815 (I934398,I934350);
nand I_54816 (I934095,I934161,I934398);
DFFARX1 I_54817 (I934350,I2507,I934118,I934438,);
not I_54818 (I934446,I934438);
not I_54819 (I934463,I1316638);
not I_54820 (I934480,I1316629);
nor I_54821 (I934497,I934480,I1316617);
nor I_54822 (I934110,I934446,I934497);
nor I_54823 (I934528,I934480,I1316620);
and I_54824 (I934545,I934528,I1316644);
or I_54825 (I934562,I934545,I1316626);
DFFARX1 I_54826 (I934562,I2507,I934118,I934588,);
nor I_54827 (I934098,I934588,I934144);
not I_54828 (I934610,I934588);
and I_54829 (I934627,I934610,I934144);
nor I_54830 (I934092,I934169,I934627);
nand I_54831 (I934658,I934610,I934220);
nor I_54832 (I934086,I934480,I934658);
nand I_54833 (I934089,I934610,I934398);
nand I_54834 (I934703,I934220,I1316629);
nor I_54835 (I934101,I934463,I934703);
not I_54836 (I934764,I2514);
DFFARX1 I_54837 (I88061,I2507,I934764,I934790,);
DFFARX1 I_54838 (I88067,I2507,I934764,I934807,);
not I_54839 (I934815,I934807);
not I_54840 (I934832,I88085);
nor I_54841 (I934849,I934832,I88064);
not I_54842 (I934866,I88070);
nor I_54843 (I934883,I934849,I88076);
nor I_54844 (I934900,I934807,I934883);
DFFARX1 I_54845 (I934900,I2507,I934764,I934750,);
nor I_54846 (I934931,I88076,I88064);
nand I_54847 (I934948,I934931,I88085);
DFFARX1 I_54848 (I934948,I2507,I934764,I934753,);
nor I_54849 (I934979,I934866,I88076);
nand I_54850 (I934996,I934979,I88082);
nor I_54851 (I935013,I934790,I934996);
DFFARX1 I_54852 (I935013,I2507,I934764,I934729,);
not I_54853 (I935044,I934996);
nand I_54854 (I934741,I934807,I935044);
DFFARX1 I_54855 (I934996,I2507,I934764,I935084,);
not I_54856 (I935092,I935084);
not I_54857 (I935109,I88076);
not I_54858 (I935126,I88064);
nor I_54859 (I935143,I935126,I88070);
nor I_54860 (I934756,I935092,I935143);
nor I_54861 (I935174,I935126,I88073);
and I_54862 (I935191,I935174,I88061);
or I_54863 (I935208,I935191,I88079);
DFFARX1 I_54864 (I935208,I2507,I934764,I935234,);
nor I_54865 (I934744,I935234,I934790);
not I_54866 (I935256,I935234);
and I_54867 (I935273,I935256,I934790);
nor I_54868 (I934738,I934815,I935273);
nand I_54869 (I935304,I935256,I934866);
nor I_54870 (I934732,I935126,I935304);
nand I_54871 (I934735,I935256,I935044);
nand I_54872 (I935349,I934866,I88064);
nor I_54873 (I934747,I935109,I935349);
not I_54874 (I935410,I2514);
DFFARX1 I_54875 (I358225,I2507,I935410,I935436,);
DFFARX1 I_54876 (I358231,I2507,I935410,I935453,);
not I_54877 (I935461,I935453);
not I_54878 (I935478,I358252);
nor I_54879 (I935495,I935478,I358240);
not I_54880 (I935512,I358249);
nor I_54881 (I935529,I935495,I358234);
nor I_54882 (I935546,I935453,I935529);
DFFARX1 I_54883 (I935546,I2507,I935410,I935396,);
nor I_54884 (I935577,I358234,I358240);
nand I_54885 (I935594,I935577,I358252);
DFFARX1 I_54886 (I935594,I2507,I935410,I935399,);
nor I_54887 (I935625,I935512,I358234);
nand I_54888 (I935642,I935625,I358225);
nor I_54889 (I935659,I935436,I935642);
DFFARX1 I_54890 (I935659,I2507,I935410,I935375,);
not I_54891 (I935690,I935642);
nand I_54892 (I935387,I935453,I935690);
DFFARX1 I_54893 (I935642,I2507,I935410,I935730,);
not I_54894 (I935738,I935730);
not I_54895 (I935755,I358234);
not I_54896 (I935772,I358237);
nor I_54897 (I935789,I935772,I358249);
nor I_54898 (I935402,I935738,I935789);
nor I_54899 (I935820,I935772,I358246);
and I_54900 (I935837,I935820,I358228);
or I_54901 (I935854,I935837,I358243);
DFFARX1 I_54902 (I935854,I2507,I935410,I935880,);
nor I_54903 (I935390,I935880,I935436);
not I_54904 (I935902,I935880);
and I_54905 (I935919,I935902,I935436);
nor I_54906 (I935384,I935461,I935919);
nand I_54907 (I935950,I935902,I935512);
nor I_54908 (I935378,I935772,I935950);
nand I_54909 (I935381,I935902,I935690);
nand I_54910 (I935995,I935512,I358237);
nor I_54911 (I935393,I935755,I935995);
not I_54912 (I936056,I2514);
DFFARX1 I_54913 (I83845,I2507,I936056,I936082,);
DFFARX1 I_54914 (I83851,I2507,I936056,I936099,);
not I_54915 (I936107,I936099);
not I_54916 (I936124,I83869);
nor I_54917 (I936141,I936124,I83848);
not I_54918 (I936158,I83854);
nor I_54919 (I936175,I936141,I83860);
nor I_54920 (I936192,I936099,I936175);
DFFARX1 I_54921 (I936192,I2507,I936056,I936042,);
nor I_54922 (I936223,I83860,I83848);
nand I_54923 (I936240,I936223,I83869);
DFFARX1 I_54924 (I936240,I2507,I936056,I936045,);
nor I_54925 (I936271,I936158,I83860);
nand I_54926 (I936288,I936271,I83866);
nor I_54927 (I936305,I936082,I936288);
DFFARX1 I_54928 (I936305,I2507,I936056,I936021,);
not I_54929 (I936336,I936288);
nand I_54930 (I936033,I936099,I936336);
DFFARX1 I_54931 (I936288,I2507,I936056,I936376,);
not I_54932 (I936384,I936376);
not I_54933 (I936401,I83860);
not I_54934 (I936418,I83848);
nor I_54935 (I936435,I936418,I83854);
nor I_54936 (I936048,I936384,I936435);
nor I_54937 (I936466,I936418,I83857);
and I_54938 (I936483,I936466,I83845);
or I_54939 (I936500,I936483,I83863);
DFFARX1 I_54940 (I936500,I2507,I936056,I936526,);
nor I_54941 (I936036,I936526,I936082);
not I_54942 (I936548,I936526);
and I_54943 (I936565,I936548,I936082);
nor I_54944 (I936030,I936107,I936565);
nand I_54945 (I936596,I936548,I936158);
nor I_54946 (I936024,I936418,I936596);
nand I_54947 (I936027,I936548,I936336);
nand I_54948 (I936641,I936158,I83848);
nor I_54949 (I936039,I936401,I936641);
not I_54950 (I936702,I2514);
DFFARX1 I_54951 (I104925,I2507,I936702,I936728,);
DFFARX1 I_54952 (I104931,I2507,I936702,I936745,);
not I_54953 (I936753,I936745);
not I_54954 (I936770,I104949);
nor I_54955 (I936787,I936770,I104928);
not I_54956 (I936804,I104934);
nor I_54957 (I936821,I936787,I104940);
nor I_54958 (I936838,I936745,I936821);
DFFARX1 I_54959 (I936838,I2507,I936702,I936688,);
nor I_54960 (I936869,I104940,I104928);
nand I_54961 (I936886,I936869,I104949);
DFFARX1 I_54962 (I936886,I2507,I936702,I936691,);
nor I_54963 (I936917,I936804,I104940);
nand I_54964 (I936934,I936917,I104946);
nor I_54965 (I936951,I936728,I936934);
DFFARX1 I_54966 (I936951,I2507,I936702,I936667,);
not I_54967 (I936982,I936934);
nand I_54968 (I936679,I936745,I936982);
DFFARX1 I_54969 (I936934,I2507,I936702,I937022,);
not I_54970 (I937030,I937022);
not I_54971 (I937047,I104940);
not I_54972 (I937064,I104928);
nor I_54973 (I937081,I937064,I104934);
nor I_54974 (I936694,I937030,I937081);
nor I_54975 (I937112,I937064,I104937);
and I_54976 (I937129,I937112,I104925);
or I_54977 (I937146,I937129,I104943);
DFFARX1 I_54978 (I937146,I2507,I936702,I937172,);
nor I_54979 (I936682,I937172,I936728);
not I_54980 (I937194,I937172);
and I_54981 (I937211,I937194,I936728);
nor I_54982 (I936676,I936753,I937211);
nand I_54983 (I937242,I937194,I936804);
nor I_54984 (I936670,I937064,I937242);
nand I_54985 (I936673,I937194,I936982);
nand I_54986 (I937287,I936804,I104928);
nor I_54987 (I936685,I937047,I937287);
not I_54988 (I937348,I2514);
DFFARX1 I_54989 (I1214516,I2507,I937348,I937374,);
DFFARX1 I_54990 (I1214522,I2507,I937348,I937391,);
not I_54991 (I937399,I937391);
not I_54992 (I937416,I1214519);
nor I_54993 (I937433,I937416,I1214498);
not I_54994 (I937450,I1214501);
nor I_54995 (I937467,I937433,I1214507);
nor I_54996 (I937484,I937391,I937467);
DFFARX1 I_54997 (I937484,I2507,I937348,I937334,);
nor I_54998 (I937515,I1214507,I1214498);
nand I_54999 (I937532,I937515,I1214519);
DFFARX1 I_55000 (I937532,I2507,I937348,I937337,);
nor I_55001 (I937563,I937450,I1214507);
nand I_55002 (I937580,I937563,I1214501);
nor I_55003 (I937597,I937374,I937580);
DFFARX1 I_55004 (I937597,I2507,I937348,I937313,);
not I_55005 (I937628,I937580);
nand I_55006 (I937325,I937391,I937628);
DFFARX1 I_55007 (I937580,I2507,I937348,I937668,);
not I_55008 (I937676,I937668);
not I_55009 (I937693,I1214507);
not I_55010 (I937710,I1214510);
nor I_55011 (I937727,I937710,I1214501);
nor I_55012 (I937340,I937676,I937727);
nor I_55013 (I937758,I937710,I1214498);
and I_55014 (I937775,I937758,I1214504);
or I_55015 (I937792,I937775,I1214513);
DFFARX1 I_55016 (I937792,I2507,I937348,I937818,);
nor I_55017 (I937328,I937818,I937374);
not I_55018 (I937840,I937818);
and I_55019 (I937857,I937840,I937374);
nor I_55020 (I937322,I937399,I937857);
nand I_55021 (I937888,I937840,I937450);
nor I_55022 (I937316,I937710,I937888);
nand I_55023 (I937319,I937840,I937628);
nand I_55024 (I937933,I937450,I1214510);
nor I_55025 (I937331,I937693,I937933);
not I_55026 (I937994,I2514);
DFFARX1 I_55027 (I41685,I2507,I937994,I938020,);
DFFARX1 I_55028 (I41691,I2507,I937994,I938037,);
not I_55029 (I938045,I938037);
not I_55030 (I938062,I41685);
nor I_55031 (I938079,I938062,I41697);
not I_55032 (I938096,I41709);
nor I_55033 (I938113,I938079,I41703);
nor I_55034 (I938130,I938037,I938113);
DFFARX1 I_55035 (I938130,I2507,I937994,I937980,);
nor I_55036 (I938161,I41703,I41697);
nand I_55037 (I938178,I938161,I41685);
DFFARX1 I_55038 (I938178,I2507,I937994,I937983,);
nor I_55039 (I938209,I938096,I41703);
nand I_55040 (I938226,I938209,I41688);
nor I_55041 (I938243,I938020,I938226);
DFFARX1 I_55042 (I938243,I2507,I937994,I937959,);
not I_55043 (I938274,I938226);
nand I_55044 (I937971,I938037,I938274);
DFFARX1 I_55045 (I938226,I2507,I937994,I938314,);
not I_55046 (I938322,I938314);
not I_55047 (I938339,I41703);
not I_55048 (I938356,I41688);
nor I_55049 (I938373,I938356,I41709);
nor I_55050 (I937986,I938322,I938373);
nor I_55051 (I938404,I938356,I41706);
and I_55052 (I938421,I938404,I41700);
or I_55053 (I938438,I938421,I41694);
DFFARX1 I_55054 (I938438,I2507,I937994,I938464,);
nor I_55055 (I937974,I938464,I938020);
not I_55056 (I938486,I938464);
and I_55057 (I938503,I938486,I938020);
nor I_55058 (I937968,I938045,I938503);
nand I_55059 (I938534,I938486,I938096);
nor I_55060 (I937962,I938356,I938534);
nand I_55061 (I937965,I938486,I938274);
nand I_55062 (I938579,I938096,I41688);
nor I_55063 (I937977,I938339,I938579);
not I_55064 (I938640,I2514);
DFFARX1 I_55065 (I773490,I2507,I938640,I938666,);
DFFARX1 I_55066 (I773484,I2507,I938640,I938683,);
not I_55067 (I938691,I938683);
not I_55068 (I938708,I773499);
nor I_55069 (I938725,I938708,I773484);
not I_55070 (I938742,I773493);
nor I_55071 (I938759,I938725,I773502);
nor I_55072 (I938776,I938683,I938759);
DFFARX1 I_55073 (I938776,I2507,I938640,I938626,);
nor I_55074 (I938807,I773502,I773484);
nand I_55075 (I938824,I938807,I773499);
DFFARX1 I_55076 (I938824,I2507,I938640,I938629,);
nor I_55077 (I938855,I938742,I773502);
nand I_55078 (I938872,I938855,I773487);
nor I_55079 (I938889,I938666,I938872);
DFFARX1 I_55080 (I938889,I2507,I938640,I938605,);
not I_55081 (I938920,I938872);
nand I_55082 (I938617,I938683,I938920);
DFFARX1 I_55083 (I938872,I2507,I938640,I938960,);
not I_55084 (I938968,I938960);
not I_55085 (I938985,I773502);
not I_55086 (I939002,I773496);
nor I_55087 (I939019,I939002,I773493);
nor I_55088 (I938632,I938968,I939019);
nor I_55089 (I939050,I939002,I773505);
and I_55090 (I939067,I939050,I773508);
or I_55091 (I939084,I939067,I773487);
DFFARX1 I_55092 (I939084,I2507,I938640,I939110,);
nor I_55093 (I938620,I939110,I938666);
not I_55094 (I939132,I939110);
and I_55095 (I939149,I939132,I938666);
nor I_55096 (I938614,I938691,I939149);
nand I_55097 (I939180,I939132,I938742);
nor I_55098 (I938608,I939002,I939180);
nand I_55099 (I938611,I939132,I938920);
nand I_55100 (I939225,I938742,I773496);
nor I_55101 (I938623,I938985,I939225);
not I_55102 (I939286,I2514);
DFFARX1 I_55103 (I350320,I2507,I939286,I939312,);
DFFARX1 I_55104 (I350326,I2507,I939286,I939329,);
not I_55105 (I939337,I939329);
not I_55106 (I939354,I350347);
nor I_55107 (I939371,I939354,I350335);
not I_55108 (I939388,I350344);
nor I_55109 (I939405,I939371,I350329);
nor I_55110 (I939422,I939329,I939405);
DFFARX1 I_55111 (I939422,I2507,I939286,I939272,);
nor I_55112 (I939453,I350329,I350335);
nand I_55113 (I939470,I939453,I350347);
DFFARX1 I_55114 (I939470,I2507,I939286,I939275,);
nor I_55115 (I939501,I939388,I350329);
nand I_55116 (I939518,I939501,I350320);
nor I_55117 (I939535,I939312,I939518);
DFFARX1 I_55118 (I939535,I2507,I939286,I939251,);
not I_55119 (I939566,I939518);
nand I_55120 (I939263,I939329,I939566);
DFFARX1 I_55121 (I939518,I2507,I939286,I939606,);
not I_55122 (I939614,I939606);
not I_55123 (I939631,I350329);
not I_55124 (I939648,I350332);
nor I_55125 (I939665,I939648,I350344);
nor I_55126 (I939278,I939614,I939665);
nor I_55127 (I939696,I939648,I350341);
and I_55128 (I939713,I939696,I350323);
or I_55129 (I939730,I939713,I350338);
DFFARX1 I_55130 (I939730,I2507,I939286,I939756,);
nor I_55131 (I939266,I939756,I939312);
not I_55132 (I939778,I939756);
and I_55133 (I939795,I939778,I939312);
nor I_55134 (I939260,I939337,I939795);
nand I_55135 (I939826,I939778,I939388);
nor I_55136 (I939254,I939648,I939826);
nand I_55137 (I939257,I939778,I939566);
nand I_55138 (I939871,I939388,I350332);
nor I_55139 (I939269,I939631,I939871);
not I_55140 (I939932,I2514);
DFFARX1 I_55141 (I665982,I2507,I939932,I939958,);
DFFARX1 I_55142 (I665976,I2507,I939932,I939975,);
not I_55143 (I939983,I939975);
not I_55144 (I940000,I665991);
nor I_55145 (I940017,I940000,I665976);
not I_55146 (I940034,I665985);
nor I_55147 (I940051,I940017,I665994);
nor I_55148 (I940068,I939975,I940051);
DFFARX1 I_55149 (I940068,I2507,I939932,I939918,);
nor I_55150 (I940099,I665994,I665976);
nand I_55151 (I940116,I940099,I665991);
DFFARX1 I_55152 (I940116,I2507,I939932,I939921,);
nor I_55153 (I940147,I940034,I665994);
nand I_55154 (I940164,I940147,I665979);
nor I_55155 (I940181,I939958,I940164);
DFFARX1 I_55156 (I940181,I2507,I939932,I939897,);
not I_55157 (I940212,I940164);
nand I_55158 (I939909,I939975,I940212);
DFFARX1 I_55159 (I940164,I2507,I939932,I940252,);
not I_55160 (I940260,I940252);
not I_55161 (I940277,I665994);
not I_55162 (I940294,I665988);
nor I_55163 (I940311,I940294,I665985);
nor I_55164 (I939924,I940260,I940311);
nor I_55165 (I940342,I940294,I665997);
and I_55166 (I940359,I940342,I666000);
or I_55167 (I940376,I940359,I665979);
DFFARX1 I_55168 (I940376,I2507,I939932,I940402,);
nor I_55169 (I939912,I940402,I939958);
not I_55170 (I940424,I940402);
and I_55171 (I940441,I940424,I939958);
nor I_55172 (I939906,I939983,I940441);
nand I_55173 (I940472,I940424,I940034);
nor I_55174 (I939900,I940294,I940472);
nand I_55175 (I939903,I940424,I940212);
nand I_55176 (I940517,I940034,I665988);
nor I_55177 (I939915,I940277,I940517);
not I_55178 (I940578,I2514);
DFFARX1 I_55179 (I1368977,I2507,I940578,I940604,);
DFFARX1 I_55180 (I1369001,I2507,I940578,I940621,);
not I_55181 (I940629,I940621);
not I_55182 (I940646,I1368983);
nor I_55183 (I940663,I940646,I1368992);
not I_55184 (I940680,I1368977);
nor I_55185 (I940697,I940663,I1368998);
nor I_55186 (I940714,I940621,I940697);
DFFARX1 I_55187 (I940714,I2507,I940578,I940564,);
nor I_55188 (I940745,I1368998,I1368992);
nand I_55189 (I940762,I940745,I1368983);
DFFARX1 I_55190 (I940762,I2507,I940578,I940567,);
nor I_55191 (I940793,I940680,I1368998);
nand I_55192 (I940810,I940793,I1368995);
nor I_55193 (I940827,I940604,I940810);
DFFARX1 I_55194 (I940827,I2507,I940578,I940543,);
not I_55195 (I940858,I940810);
nand I_55196 (I940555,I940621,I940858);
DFFARX1 I_55197 (I940810,I2507,I940578,I940898,);
not I_55198 (I940906,I940898);
not I_55199 (I940923,I1368998);
not I_55200 (I940940,I1368989);
nor I_55201 (I940957,I940940,I1368977);
nor I_55202 (I940570,I940906,I940957);
nor I_55203 (I940988,I940940,I1368980);
and I_55204 (I941005,I940988,I1369004);
or I_55205 (I941022,I941005,I1368986);
DFFARX1 I_55206 (I941022,I2507,I940578,I941048,);
nor I_55207 (I940558,I941048,I940604);
not I_55208 (I941070,I941048);
and I_55209 (I941087,I941070,I940604);
nor I_55210 (I940552,I940629,I941087);
nand I_55211 (I941118,I941070,I940680);
nor I_55212 (I940546,I940940,I941118);
nand I_55213 (I940549,I941070,I940858);
nand I_55214 (I941163,I940680,I1368989);
nor I_55215 (I940561,I940923,I941163);
not I_55216 (I941224,I2514);
DFFARX1 I_55217 (I257568,I2507,I941224,I941250,);
DFFARX1 I_55218 (I257574,I2507,I941224,I941267,);
not I_55219 (I941275,I941267);
not I_55220 (I941292,I257595);
nor I_55221 (I941309,I941292,I257583);
not I_55222 (I941326,I257592);
nor I_55223 (I941343,I941309,I257577);
nor I_55224 (I941360,I941267,I941343);
DFFARX1 I_55225 (I941360,I2507,I941224,I941210,);
nor I_55226 (I941391,I257577,I257583);
nand I_55227 (I941408,I941391,I257595);
DFFARX1 I_55228 (I941408,I2507,I941224,I941213,);
nor I_55229 (I941439,I941326,I257577);
nand I_55230 (I941456,I941439,I257568);
nor I_55231 (I941473,I941250,I941456);
DFFARX1 I_55232 (I941473,I2507,I941224,I941189,);
not I_55233 (I941504,I941456);
nand I_55234 (I941201,I941267,I941504);
DFFARX1 I_55235 (I941456,I2507,I941224,I941544,);
not I_55236 (I941552,I941544);
not I_55237 (I941569,I257577);
not I_55238 (I941586,I257580);
nor I_55239 (I941603,I941586,I257592);
nor I_55240 (I941216,I941552,I941603);
nor I_55241 (I941634,I941586,I257589);
and I_55242 (I941651,I941634,I257571);
or I_55243 (I941668,I941651,I257586);
DFFARX1 I_55244 (I941668,I2507,I941224,I941694,);
nor I_55245 (I941204,I941694,I941250);
not I_55246 (I941716,I941694);
and I_55247 (I941733,I941716,I941250);
nor I_55248 (I941198,I941275,I941733);
nand I_55249 (I941764,I941716,I941326);
nor I_55250 (I941192,I941586,I941764);
nand I_55251 (I941195,I941716,I941504);
nand I_55252 (I941809,I941326,I257580);
nor I_55253 (I941207,I941569,I941809);
not I_55254 (I941870,I2514);
DFFARX1 I_55255 (I793822,I2507,I941870,I941896,);
DFFARX1 I_55256 (I793819,I2507,I941870,I941913,);
not I_55257 (I941921,I941913);
not I_55258 (I941938,I793819);
nor I_55259 (I941955,I941938,I793822);
not I_55260 (I941972,I793834);
nor I_55261 (I941989,I941955,I793828);
nor I_55262 (I942006,I941913,I941989);
DFFARX1 I_55263 (I942006,I2507,I941870,I941856,);
nor I_55264 (I942037,I793828,I793822);
nand I_55265 (I942054,I942037,I793819);
DFFARX1 I_55266 (I942054,I2507,I941870,I941859,);
nor I_55267 (I942085,I941972,I793828);
nand I_55268 (I942102,I942085,I793816);
nor I_55269 (I942119,I941896,I942102);
DFFARX1 I_55270 (I942119,I2507,I941870,I941835,);
not I_55271 (I942150,I942102);
nand I_55272 (I941847,I941913,I942150);
DFFARX1 I_55273 (I942102,I2507,I941870,I942190,);
not I_55274 (I942198,I942190);
not I_55275 (I942215,I793828);
not I_55276 (I942232,I793825);
nor I_55277 (I942249,I942232,I793834);
nor I_55278 (I941862,I942198,I942249);
nor I_55279 (I942280,I942232,I793831);
and I_55280 (I942297,I942280,I793837);
or I_55281 (I942314,I942297,I793816);
DFFARX1 I_55282 (I942314,I2507,I941870,I942340,);
nor I_55283 (I941850,I942340,I941896);
not I_55284 (I942362,I942340);
and I_55285 (I942379,I942362,I941896);
nor I_55286 (I941844,I941921,I942379);
nand I_55287 (I942410,I942362,I941972);
nor I_55288 (I941838,I942232,I942410);
nand I_55289 (I941841,I942362,I942150);
nand I_55290 (I942455,I941972,I793825);
nor I_55291 (I941853,I942215,I942455);
not I_55292 (I942516,I2514);
DFFARX1 I_55293 (I462645,I2507,I942516,I942542,);
DFFARX1 I_55294 (I462642,I2507,I942516,I942559,);
not I_55295 (I942567,I942559);
not I_55296 (I942584,I462657);
nor I_55297 (I942601,I942584,I462660);
not I_55298 (I942618,I462648);
nor I_55299 (I942635,I942601,I462654);
nor I_55300 (I942652,I942559,I942635);
DFFARX1 I_55301 (I942652,I2507,I942516,I942502,);
nor I_55302 (I942683,I462654,I462660);
nand I_55303 (I942700,I942683,I462657);
DFFARX1 I_55304 (I942700,I2507,I942516,I942505,);
nor I_55305 (I942731,I942618,I462654);
nand I_55306 (I942748,I942731,I462666);
nor I_55307 (I942765,I942542,I942748);
DFFARX1 I_55308 (I942765,I2507,I942516,I942481,);
not I_55309 (I942796,I942748);
nand I_55310 (I942493,I942559,I942796);
DFFARX1 I_55311 (I942748,I2507,I942516,I942836,);
not I_55312 (I942844,I942836);
not I_55313 (I942861,I462654);
not I_55314 (I942878,I462639);
nor I_55315 (I942895,I942878,I462648);
nor I_55316 (I942508,I942844,I942895);
nor I_55317 (I942926,I942878,I462651);
and I_55318 (I942943,I942926,I462639);
or I_55319 (I942960,I942943,I462663);
DFFARX1 I_55320 (I942960,I2507,I942516,I942986,);
nor I_55321 (I942496,I942986,I942542);
not I_55322 (I943008,I942986);
and I_55323 (I943025,I943008,I942542);
nor I_55324 (I942490,I942567,I943025);
nand I_55325 (I943056,I943008,I942618);
nor I_55326 (I942484,I942878,I943056);
nand I_55327 (I942487,I943008,I942796);
nand I_55328 (I943101,I942618,I462639);
nor I_55329 (I942499,I942861,I943101);
not I_55330 (I943162,I2514);
DFFARX1 I_55331 (I619161,I2507,I943162,I943188,);
DFFARX1 I_55332 (I619173,I2507,I943162,I943205,);
not I_55333 (I943213,I943205);
not I_55334 (I943230,I619182);
nor I_55335 (I943247,I943230,I619158);
not I_55336 (I943264,I619176);
nor I_55337 (I943281,I943247,I619170);
nor I_55338 (I943298,I943205,I943281);
DFFARX1 I_55339 (I943298,I2507,I943162,I943148,);
nor I_55340 (I943329,I619170,I619158);
nand I_55341 (I943346,I943329,I619182);
DFFARX1 I_55342 (I943346,I2507,I943162,I943151,);
nor I_55343 (I943377,I943264,I619170);
nand I_55344 (I943394,I943377,I619164);
nor I_55345 (I943411,I943188,I943394);
DFFARX1 I_55346 (I943411,I2507,I943162,I943127,);
not I_55347 (I943442,I943394);
nand I_55348 (I943139,I943205,I943442);
DFFARX1 I_55349 (I943394,I2507,I943162,I943482,);
not I_55350 (I943490,I943482);
not I_55351 (I943507,I619170);
not I_55352 (I943524,I619179);
nor I_55353 (I943541,I943524,I619176);
nor I_55354 (I943154,I943490,I943541);
nor I_55355 (I943572,I943524,I619161);
and I_55356 (I943589,I943572,I619158);
or I_55357 (I943606,I943589,I619167);
DFFARX1 I_55358 (I943606,I2507,I943162,I943632,);
nor I_55359 (I943142,I943632,I943188);
not I_55360 (I943654,I943632);
and I_55361 (I943671,I943654,I943188);
nor I_55362 (I943136,I943213,I943671);
nand I_55363 (I943702,I943654,I943264);
nor I_55364 (I943130,I943524,I943702);
nand I_55365 (I943133,I943654,I943442);
nand I_55366 (I943747,I943264,I619179);
nor I_55367 (I943145,I943507,I943747);
not I_55368 (I943808,I2514);
DFFARX1 I_55369 (I796984,I2507,I943808,I943834,);
DFFARX1 I_55370 (I796981,I2507,I943808,I943851,);
not I_55371 (I943859,I943851);
not I_55372 (I943876,I796981);
nor I_55373 (I943893,I943876,I796984);
not I_55374 (I943910,I796996);
nor I_55375 (I943927,I943893,I796990);
nor I_55376 (I943944,I943851,I943927);
DFFARX1 I_55377 (I943944,I2507,I943808,I943794,);
nor I_55378 (I943975,I796990,I796984);
nand I_55379 (I943992,I943975,I796981);
DFFARX1 I_55380 (I943992,I2507,I943808,I943797,);
nor I_55381 (I944023,I943910,I796990);
nand I_55382 (I944040,I944023,I796978);
nor I_55383 (I944057,I943834,I944040);
DFFARX1 I_55384 (I944057,I2507,I943808,I943773,);
not I_55385 (I944088,I944040);
nand I_55386 (I943785,I943851,I944088);
DFFARX1 I_55387 (I944040,I2507,I943808,I944128,);
not I_55388 (I944136,I944128);
not I_55389 (I944153,I796990);
not I_55390 (I944170,I796987);
nor I_55391 (I944187,I944170,I796996);
nor I_55392 (I943800,I944136,I944187);
nor I_55393 (I944218,I944170,I796993);
and I_55394 (I944235,I944218,I796999);
or I_55395 (I944252,I944235,I796978);
DFFARX1 I_55396 (I944252,I2507,I943808,I944278,);
nor I_55397 (I943788,I944278,I943834);
not I_55398 (I944300,I944278);
and I_55399 (I944317,I944300,I943834);
nor I_55400 (I943782,I943859,I944317);
nand I_55401 (I944348,I944300,I943910);
nor I_55402 (I943776,I944170,I944348);
nand I_55403 (I943779,I944300,I944088);
nand I_55404 (I944393,I943910,I796987);
nor I_55405 (I943791,I944153,I944393);
not I_55406 (I944454,I2514);
DFFARX1 I_55407 (I309214,I2507,I944454,I944480,);
DFFARX1 I_55408 (I309220,I2507,I944454,I944497,);
not I_55409 (I944505,I944497);
not I_55410 (I944522,I309241);
nor I_55411 (I944539,I944522,I309229);
not I_55412 (I944556,I309238);
nor I_55413 (I944573,I944539,I309223);
nor I_55414 (I944590,I944497,I944573);
DFFARX1 I_55415 (I944590,I2507,I944454,I944440,);
nor I_55416 (I944621,I309223,I309229);
nand I_55417 (I944638,I944621,I309241);
DFFARX1 I_55418 (I944638,I2507,I944454,I944443,);
nor I_55419 (I944669,I944556,I309223);
nand I_55420 (I944686,I944669,I309214);
nor I_55421 (I944703,I944480,I944686);
DFFARX1 I_55422 (I944703,I2507,I944454,I944419,);
not I_55423 (I944734,I944686);
nand I_55424 (I944431,I944497,I944734);
DFFARX1 I_55425 (I944686,I2507,I944454,I944774,);
not I_55426 (I944782,I944774);
not I_55427 (I944799,I309223);
not I_55428 (I944816,I309226);
nor I_55429 (I944833,I944816,I309238);
nor I_55430 (I944446,I944782,I944833);
nor I_55431 (I944864,I944816,I309235);
and I_55432 (I944881,I944864,I309217);
or I_55433 (I944898,I944881,I309232);
DFFARX1 I_55434 (I944898,I2507,I944454,I944924,);
nor I_55435 (I944434,I944924,I944480);
not I_55436 (I944946,I944924);
and I_55437 (I944963,I944946,I944480);
nor I_55438 (I944428,I944505,I944963);
nand I_55439 (I944994,I944946,I944556);
nor I_55440 (I944422,I944816,I944994);
nand I_55441 (I944425,I944946,I944734);
nand I_55442 (I945039,I944556,I309226);
nor I_55443 (I944437,I944799,I945039);
not I_55444 (I945100,I2514);
DFFARX1 I_55445 (I203786,I2507,I945100,I945126,);
DFFARX1 I_55446 (I203798,I2507,I945100,I945143,);
not I_55447 (I945151,I945143);
not I_55448 (I945168,I203804);
nor I_55449 (I945185,I945168,I203789);
not I_55450 (I945202,I203780);
nor I_55451 (I945219,I945185,I203801);
nor I_55452 (I945236,I945143,I945219);
DFFARX1 I_55453 (I945236,I2507,I945100,I945086,);
nor I_55454 (I945267,I203801,I203789);
nand I_55455 (I945284,I945267,I203804);
DFFARX1 I_55456 (I945284,I2507,I945100,I945089,);
nor I_55457 (I945315,I945202,I203801);
nand I_55458 (I945332,I945315,I203783);
nor I_55459 (I945349,I945126,I945332);
DFFARX1 I_55460 (I945349,I2507,I945100,I945065,);
not I_55461 (I945380,I945332);
nand I_55462 (I945077,I945143,I945380);
DFFARX1 I_55463 (I945332,I2507,I945100,I945420,);
not I_55464 (I945428,I945420);
not I_55465 (I945445,I203801);
not I_55466 (I945462,I203792);
nor I_55467 (I945479,I945462,I203780);
nor I_55468 (I945092,I945428,I945479);
nor I_55469 (I945510,I945462,I203795);
and I_55470 (I945527,I945510,I203783);
or I_55471 (I945544,I945527,I203780);
DFFARX1 I_55472 (I945544,I2507,I945100,I945570,);
nor I_55473 (I945080,I945570,I945126);
not I_55474 (I945592,I945570);
and I_55475 (I945609,I945592,I945126);
nor I_55476 (I945074,I945151,I945609);
nand I_55477 (I945640,I945592,I945202);
nor I_55478 (I945068,I945462,I945640);
nand I_55479 (I945071,I945592,I945380);
nand I_55480 (I945685,I945202,I203792);
nor I_55481 (I945083,I945445,I945685);
not I_55482 (I945746,I2514);
DFFARX1 I_55483 (I387573,I2507,I945746,I945772,);
DFFARX1 I_55484 (I387570,I2507,I945746,I945789,);
not I_55485 (I945797,I945789);
not I_55486 (I945814,I387585);
nor I_55487 (I945831,I945814,I387588);
not I_55488 (I945848,I387576);
nor I_55489 (I945865,I945831,I387582);
nor I_55490 (I945882,I945789,I945865);
DFFARX1 I_55491 (I945882,I2507,I945746,I945732,);
nor I_55492 (I945913,I387582,I387588);
nand I_55493 (I945930,I945913,I387585);
DFFARX1 I_55494 (I945930,I2507,I945746,I945735,);
nor I_55495 (I945961,I945848,I387582);
nand I_55496 (I945978,I945961,I387594);
nor I_55497 (I945995,I945772,I945978);
DFFARX1 I_55498 (I945995,I2507,I945746,I945711,);
not I_55499 (I946026,I945978);
nand I_55500 (I945723,I945789,I946026);
DFFARX1 I_55501 (I945978,I2507,I945746,I946066,);
not I_55502 (I946074,I946066);
not I_55503 (I946091,I387582);
not I_55504 (I946108,I387567);
nor I_55505 (I946125,I946108,I387576);
nor I_55506 (I945738,I946074,I946125);
nor I_55507 (I946156,I946108,I387579);
and I_55508 (I946173,I946156,I387567);
or I_55509 (I946190,I946173,I387591);
DFFARX1 I_55510 (I946190,I2507,I945746,I946216,);
nor I_55511 (I945726,I946216,I945772);
not I_55512 (I946238,I946216);
and I_55513 (I946255,I946238,I945772);
nor I_55514 (I945720,I945797,I946255);
nand I_55515 (I946286,I946238,I945848);
nor I_55516 (I945714,I946108,I946286);
nand I_55517 (I945717,I946238,I946026);
nand I_55518 (I946331,I945848,I387567);
nor I_55519 (I945729,I946091,I946331);
not I_55520 (I946392,I2514);
DFFARX1 I_55521 (I432181,I2507,I946392,I946418,);
DFFARX1 I_55522 (I432178,I2507,I946392,I946435,);
not I_55523 (I946443,I946435);
not I_55524 (I946460,I432193);
nor I_55525 (I946477,I946460,I432196);
not I_55526 (I946494,I432184);
nor I_55527 (I946511,I946477,I432190);
nor I_55528 (I946528,I946435,I946511);
DFFARX1 I_55529 (I946528,I2507,I946392,I946378,);
nor I_55530 (I946559,I432190,I432196);
nand I_55531 (I946576,I946559,I432193);
DFFARX1 I_55532 (I946576,I2507,I946392,I946381,);
nor I_55533 (I946607,I946494,I432190);
nand I_55534 (I946624,I946607,I432202);
nor I_55535 (I946641,I946418,I946624);
DFFARX1 I_55536 (I946641,I2507,I946392,I946357,);
not I_55537 (I946672,I946624);
nand I_55538 (I946369,I946435,I946672);
DFFARX1 I_55539 (I946624,I2507,I946392,I946712,);
not I_55540 (I946720,I946712);
not I_55541 (I946737,I432190);
not I_55542 (I946754,I432175);
nor I_55543 (I946771,I946754,I432184);
nor I_55544 (I946384,I946720,I946771);
nor I_55545 (I946802,I946754,I432187);
and I_55546 (I946819,I946802,I432175);
or I_55547 (I946836,I946819,I432199);
DFFARX1 I_55548 (I946836,I2507,I946392,I946862,);
nor I_55549 (I946372,I946862,I946418);
not I_55550 (I946884,I946862);
and I_55551 (I946901,I946884,I946418);
nor I_55552 (I946366,I946443,I946901);
nand I_55553 (I946932,I946884,I946494);
nor I_55554 (I946360,I946754,I946932);
nand I_55555 (I946363,I946884,I946672);
nand I_55556 (I946977,I946494,I432175);
nor I_55557 (I946375,I946737,I946977);
not I_55558 (I947038,I2514);
DFFARX1 I_55559 (I1276727,I2507,I947038,I947064,);
DFFARX1 I_55560 (I1276721,I2507,I947038,I947081,);
not I_55561 (I947089,I947081);
not I_55562 (I947106,I1276730);
nor I_55563 (I947123,I947106,I1276742);
not I_55564 (I947140,I1276724);
nor I_55565 (I947157,I947123,I1276721);
nor I_55566 (I947174,I947081,I947157);
DFFARX1 I_55567 (I947174,I2507,I947038,I947024,);
nor I_55568 (I947205,I1276721,I1276742);
nand I_55569 (I947222,I947205,I1276730);
DFFARX1 I_55570 (I947222,I2507,I947038,I947027,);
nor I_55571 (I947253,I947140,I1276721);
nand I_55572 (I947270,I947253,I1276718);
nor I_55573 (I947287,I947064,I947270);
DFFARX1 I_55574 (I947287,I2507,I947038,I947003,);
not I_55575 (I947318,I947270);
nand I_55576 (I947015,I947081,I947318);
DFFARX1 I_55577 (I947270,I2507,I947038,I947358,);
not I_55578 (I947366,I947358);
not I_55579 (I947383,I1276721);
not I_55580 (I947400,I1276739);
nor I_55581 (I947417,I947400,I1276724);
nor I_55582 (I947030,I947366,I947417);
nor I_55583 (I947448,I947400,I1276733);
and I_55584 (I947465,I947448,I1276718);
or I_55585 (I947482,I947465,I1276736);
DFFARX1 I_55586 (I947482,I2507,I947038,I947508,);
nor I_55587 (I947018,I947508,I947064);
not I_55588 (I947530,I947508);
and I_55589 (I947547,I947530,I947064);
nor I_55590 (I947012,I947089,I947547);
nand I_55591 (I947578,I947530,I947140);
nor I_55592 (I947006,I947400,I947578);
nand I_55593 (I947009,I947530,I947318);
nand I_55594 (I947623,I947140,I1276739);
nor I_55595 (I947021,I947383,I947623);
not I_55596 (I947684,I2514);
DFFARX1 I_55597 (I73832,I2507,I947684,I947710,);
DFFARX1 I_55598 (I73838,I2507,I947684,I947727,);
not I_55599 (I947735,I947727);
not I_55600 (I947752,I73856);
nor I_55601 (I947769,I947752,I73835);
not I_55602 (I947786,I73841);
nor I_55603 (I947803,I947769,I73847);
nor I_55604 (I947820,I947727,I947803);
DFFARX1 I_55605 (I947820,I2507,I947684,I947670,);
nor I_55606 (I947851,I73847,I73835);
nand I_55607 (I947868,I947851,I73856);
DFFARX1 I_55608 (I947868,I2507,I947684,I947673,);
nor I_55609 (I947899,I947786,I73847);
nand I_55610 (I947916,I947899,I73853);
nor I_55611 (I947933,I947710,I947916);
DFFARX1 I_55612 (I947933,I2507,I947684,I947649,);
not I_55613 (I947964,I947916);
nand I_55614 (I947661,I947727,I947964);
DFFARX1 I_55615 (I947916,I2507,I947684,I948004,);
not I_55616 (I948012,I948004);
not I_55617 (I948029,I73847);
not I_55618 (I948046,I73835);
nor I_55619 (I948063,I948046,I73841);
nor I_55620 (I947676,I948012,I948063);
nor I_55621 (I948094,I948046,I73844);
and I_55622 (I948111,I948094,I73832);
or I_55623 (I948128,I948111,I73850);
DFFARX1 I_55624 (I948128,I2507,I947684,I948154,);
nor I_55625 (I947664,I948154,I947710);
not I_55626 (I948176,I948154);
and I_55627 (I948193,I948176,I947710);
nor I_55628 (I947658,I947735,I948193);
nand I_55629 (I948224,I948176,I947786);
nor I_55630 (I947652,I948046,I948224);
nand I_55631 (I947655,I948176,I947964);
nand I_55632 (I948269,I947786,I73835);
nor I_55633 (I947667,I948029,I948269);
not I_55634 (I948330,I2514);
DFFARX1 I_55635 (I382677,I2507,I948330,I948356,);
DFFARX1 I_55636 (I382674,I2507,I948330,I948373,);
not I_55637 (I948381,I948373);
not I_55638 (I948398,I382689);
nor I_55639 (I948415,I948398,I382692);
not I_55640 (I948432,I382680);
nor I_55641 (I948449,I948415,I382686);
nor I_55642 (I948466,I948373,I948449);
DFFARX1 I_55643 (I948466,I2507,I948330,I948316,);
nor I_55644 (I948497,I382686,I382692);
nand I_55645 (I948514,I948497,I382689);
DFFARX1 I_55646 (I948514,I2507,I948330,I948319,);
nor I_55647 (I948545,I948432,I382686);
nand I_55648 (I948562,I948545,I382698);
nor I_55649 (I948579,I948356,I948562);
DFFARX1 I_55650 (I948579,I2507,I948330,I948295,);
not I_55651 (I948610,I948562);
nand I_55652 (I948307,I948373,I948610);
DFFARX1 I_55653 (I948562,I2507,I948330,I948650,);
not I_55654 (I948658,I948650);
not I_55655 (I948675,I382686);
not I_55656 (I948692,I382671);
nor I_55657 (I948709,I948692,I382680);
nor I_55658 (I948322,I948658,I948709);
nor I_55659 (I948740,I948692,I382683);
and I_55660 (I948757,I948740,I382671);
or I_55661 (I948774,I948757,I382695);
DFFARX1 I_55662 (I948774,I2507,I948330,I948800,);
nor I_55663 (I948310,I948800,I948356);
not I_55664 (I948822,I948800);
and I_55665 (I948839,I948822,I948356);
nor I_55666 (I948304,I948381,I948839);
nand I_55667 (I948870,I948822,I948432);
nor I_55668 (I948298,I948692,I948870);
nand I_55669 (I948301,I948822,I948610);
nand I_55670 (I948915,I948432,I382671);
nor I_55671 (I948313,I948675,I948915);
not I_55672 (I948976,I2514);
DFFARX1 I_55673 (I507777,I2507,I948976,I949002,);
DFFARX1 I_55674 (I507789,I2507,I948976,I949019,);
not I_55675 (I949027,I949019);
not I_55676 (I949044,I507774);
nor I_55677 (I949061,I949044,I507792);
not I_55678 (I949078,I507798);
nor I_55679 (I949095,I949061,I507780);
nor I_55680 (I949112,I949019,I949095);
DFFARX1 I_55681 (I949112,I2507,I948976,I948962,);
nor I_55682 (I949143,I507780,I507792);
nand I_55683 (I949160,I949143,I507774);
DFFARX1 I_55684 (I949160,I2507,I948976,I948965,);
nor I_55685 (I949191,I949078,I507780);
nand I_55686 (I949208,I949191,I507783);
nor I_55687 (I949225,I949002,I949208);
DFFARX1 I_55688 (I949225,I2507,I948976,I948941,);
not I_55689 (I949256,I949208);
nand I_55690 (I948953,I949019,I949256);
DFFARX1 I_55691 (I949208,I2507,I948976,I949296,);
not I_55692 (I949304,I949296);
not I_55693 (I949321,I507780);
not I_55694 (I949338,I507786);
nor I_55695 (I949355,I949338,I507798);
nor I_55696 (I948968,I949304,I949355);
nor I_55697 (I949386,I949338,I507795);
and I_55698 (I949403,I949386,I507774);
or I_55699 (I949420,I949403,I507777);
DFFARX1 I_55700 (I949420,I2507,I948976,I949446,);
nor I_55701 (I948956,I949446,I949002);
not I_55702 (I949468,I949446);
and I_55703 (I949485,I949468,I949002);
nor I_55704 (I948950,I949027,I949485);
nand I_55705 (I949516,I949468,I949078);
nor I_55706 (I948944,I949338,I949516);
nand I_55707 (I948947,I949468,I949256);
nand I_55708 (I949561,I949078,I507786);
nor I_55709 (I948959,I949321,I949561);
not I_55710 (I949622,I2514);
DFFARX1 I_55711 (I1077462,I2507,I949622,I949648,);
DFFARX1 I_55712 (I1077444,I2507,I949622,I949665,);
not I_55713 (I949673,I949665);
not I_55714 (I949690,I1077453);
nor I_55715 (I949707,I949690,I1077465);
not I_55716 (I949724,I1077447);
nor I_55717 (I949741,I949707,I1077456);
nor I_55718 (I949758,I949665,I949741);
DFFARX1 I_55719 (I949758,I2507,I949622,I949608,);
nor I_55720 (I949789,I1077456,I1077465);
nand I_55721 (I949806,I949789,I1077453);
DFFARX1 I_55722 (I949806,I2507,I949622,I949611,);
nor I_55723 (I949837,I949724,I1077456);
nand I_55724 (I949854,I949837,I1077468);
nor I_55725 (I949871,I949648,I949854);
DFFARX1 I_55726 (I949871,I2507,I949622,I949587,);
not I_55727 (I949902,I949854);
nand I_55728 (I949599,I949665,I949902);
DFFARX1 I_55729 (I949854,I2507,I949622,I949942,);
not I_55730 (I949950,I949942);
not I_55731 (I949967,I1077456);
not I_55732 (I949984,I1077444);
nor I_55733 (I950001,I949984,I1077447);
nor I_55734 (I949614,I949950,I950001);
nor I_55735 (I950032,I949984,I1077450);
and I_55736 (I950049,I950032,I1077459);
or I_55737 (I950066,I950049,I1077447);
DFFARX1 I_55738 (I950066,I2507,I949622,I950092,);
nor I_55739 (I949602,I950092,I949648);
not I_55740 (I950114,I950092);
and I_55741 (I950131,I950114,I949648);
nor I_55742 (I949596,I949673,I950131);
nand I_55743 (I950162,I950114,I949724);
nor I_55744 (I949590,I949984,I950162);
nand I_55745 (I949593,I950114,I949902);
nand I_55746 (I950207,I949724,I1077444);
nor I_55747 (I949605,I949967,I950207);
not I_55748 (I950268,I2514);
DFFARX1 I_55749 (I248411,I2507,I950268,I950294,);
DFFARX1 I_55750 (I248423,I2507,I950268,I950311,);
not I_55751 (I950319,I950311);
not I_55752 (I950336,I248429);
nor I_55753 (I950353,I950336,I248414);
not I_55754 (I950370,I248405);
nor I_55755 (I950387,I950353,I248426);
nor I_55756 (I950404,I950311,I950387);
DFFARX1 I_55757 (I950404,I2507,I950268,I950254,);
nor I_55758 (I950435,I248426,I248414);
nand I_55759 (I950452,I950435,I248429);
DFFARX1 I_55760 (I950452,I2507,I950268,I950257,);
nor I_55761 (I950483,I950370,I248426);
nand I_55762 (I950500,I950483,I248408);
nor I_55763 (I950517,I950294,I950500);
DFFARX1 I_55764 (I950517,I2507,I950268,I950233,);
not I_55765 (I950548,I950500);
nand I_55766 (I950245,I950311,I950548);
DFFARX1 I_55767 (I950500,I2507,I950268,I950588,);
not I_55768 (I950596,I950588);
not I_55769 (I950613,I248426);
not I_55770 (I950630,I248417);
nor I_55771 (I950647,I950630,I248405);
nor I_55772 (I950260,I950596,I950647);
nor I_55773 (I950678,I950630,I248420);
and I_55774 (I950695,I950678,I248408);
or I_55775 (I950712,I950695,I248405);
DFFARX1 I_55776 (I950712,I2507,I950268,I950738,);
nor I_55777 (I950248,I950738,I950294);
not I_55778 (I950760,I950738);
and I_55779 (I950777,I950760,I950294);
nor I_55780 (I950242,I950319,I950777);
nand I_55781 (I950808,I950760,I950370);
nor I_55782 (I950236,I950630,I950808);
nand I_55783 (I950239,I950760,I950548);
nand I_55784 (I950853,I950370,I248417);
nor I_55785 (I950251,I950613,I950853);
not I_55786 (I950914,I2514);
DFFARX1 I_55787 (I157376,I2507,I950914,I950940,);
DFFARX1 I_55788 (I157388,I2507,I950914,I950957,);
not I_55789 (I950965,I950957);
not I_55790 (I950982,I157394);
nor I_55791 (I950999,I950982,I157379);
not I_55792 (I951016,I157370);
nor I_55793 (I951033,I950999,I157391);
nor I_55794 (I951050,I950957,I951033);
DFFARX1 I_55795 (I951050,I2507,I950914,I950900,);
nor I_55796 (I951081,I157391,I157379);
nand I_55797 (I951098,I951081,I157394);
DFFARX1 I_55798 (I951098,I2507,I950914,I950903,);
nor I_55799 (I951129,I951016,I157391);
nand I_55800 (I951146,I951129,I157373);
nor I_55801 (I951163,I950940,I951146);
DFFARX1 I_55802 (I951163,I2507,I950914,I950879,);
not I_55803 (I951194,I951146);
nand I_55804 (I950891,I950957,I951194);
DFFARX1 I_55805 (I951146,I2507,I950914,I951234,);
not I_55806 (I951242,I951234);
not I_55807 (I951259,I157391);
not I_55808 (I951276,I157382);
nor I_55809 (I951293,I951276,I157370);
nor I_55810 (I950906,I951242,I951293);
nor I_55811 (I951324,I951276,I157385);
and I_55812 (I951341,I951324,I157373);
or I_55813 (I951358,I951341,I157370);
DFFARX1 I_55814 (I951358,I2507,I950914,I951384,);
nor I_55815 (I950894,I951384,I950940);
not I_55816 (I951406,I951384);
and I_55817 (I951423,I951406,I950940);
nor I_55818 (I950888,I950965,I951423);
nand I_55819 (I951454,I951406,I951016);
nor I_55820 (I950882,I951276,I951454);
nand I_55821 (I950885,I951406,I951194);
nand I_55822 (I951499,I951016,I157382);
nor I_55823 (I950897,I951259,I951499);
not I_55824 (I951560,I2514);
DFFARX1 I_55825 (I1042679,I2507,I951560,I951586,);
DFFARX1 I_55826 (I1042682,I2507,I951560,I951603,);
not I_55827 (I951611,I951603);
not I_55828 (I951628,I1042679);
nor I_55829 (I951645,I951628,I1042691);
not I_55830 (I951662,I1042700);
nor I_55831 (I951679,I951645,I1042688);
nor I_55832 (I951696,I951603,I951679);
DFFARX1 I_55833 (I951696,I2507,I951560,I951546,);
nor I_55834 (I951727,I1042688,I1042691);
nand I_55835 (I951744,I951727,I1042679);
DFFARX1 I_55836 (I951744,I2507,I951560,I951549,);
nor I_55837 (I951775,I951662,I1042688);
nand I_55838 (I951792,I951775,I1042694);
nor I_55839 (I951809,I951586,I951792);
DFFARX1 I_55840 (I951809,I2507,I951560,I951525,);
not I_55841 (I951840,I951792);
nand I_55842 (I951537,I951603,I951840);
DFFARX1 I_55843 (I951792,I2507,I951560,I951880,);
not I_55844 (I951888,I951880);
not I_55845 (I951905,I1042688);
not I_55846 (I951922,I1042685);
nor I_55847 (I951939,I951922,I1042700);
nor I_55848 (I951552,I951888,I951939);
nor I_55849 (I951970,I951922,I1042697);
and I_55850 (I951987,I951970,I1042685);
or I_55851 (I952004,I951987,I1042682);
DFFARX1 I_55852 (I952004,I2507,I951560,I952030,);
nor I_55853 (I951540,I952030,I951586);
not I_55854 (I952052,I952030);
and I_55855 (I952069,I952052,I951586);
nor I_55856 (I951534,I951611,I952069);
nand I_55857 (I952100,I952052,I951662);
nor I_55858 (I951528,I951922,I952100);
nand I_55859 (I951531,I952052,I951840);
nand I_55860 (I952145,I951662,I1042685);
nor I_55861 (I951543,I951905,I952145);
not I_55862 (I952206,I2514);
DFFARX1 I_55863 (I1333277,I2507,I952206,I952232,);
DFFARX1 I_55864 (I1333301,I2507,I952206,I952249,);
not I_55865 (I952257,I952249);
not I_55866 (I952274,I1333283);
nor I_55867 (I952291,I952274,I1333292);
not I_55868 (I952308,I1333277);
nor I_55869 (I952325,I952291,I1333298);
nor I_55870 (I952342,I952249,I952325);
DFFARX1 I_55871 (I952342,I2507,I952206,I952192,);
nor I_55872 (I952373,I1333298,I1333292);
nand I_55873 (I952390,I952373,I1333283);
DFFARX1 I_55874 (I952390,I2507,I952206,I952195,);
nor I_55875 (I952421,I952308,I1333298);
nand I_55876 (I952438,I952421,I1333295);
nor I_55877 (I952455,I952232,I952438);
DFFARX1 I_55878 (I952455,I2507,I952206,I952171,);
not I_55879 (I952486,I952438);
nand I_55880 (I952183,I952249,I952486);
DFFARX1 I_55881 (I952438,I2507,I952206,I952526,);
not I_55882 (I952534,I952526);
not I_55883 (I952551,I1333298);
not I_55884 (I952568,I1333289);
nor I_55885 (I952585,I952568,I1333277);
nor I_55886 (I952198,I952534,I952585);
nor I_55887 (I952616,I952568,I1333280);
and I_55888 (I952633,I952616,I1333304);
or I_55889 (I952650,I952633,I1333286);
DFFARX1 I_55890 (I952650,I2507,I952206,I952676,);
nor I_55891 (I952186,I952676,I952232);
not I_55892 (I952698,I952676);
and I_55893 (I952715,I952698,I952232);
nor I_55894 (I952180,I952257,I952715);
nand I_55895 (I952746,I952698,I952308);
nor I_55896 (I952174,I952568,I952746);
nand I_55897 (I952177,I952698,I952486);
nand I_55898 (I952791,I952308,I1333289);
nor I_55899 (I952189,I952551,I952791);
not I_55900 (I952852,I2514);
DFFARX1 I_55901 (I288661,I2507,I952852,I952878,);
DFFARX1 I_55902 (I288667,I2507,I952852,I952895,);
not I_55903 (I952903,I952895);
not I_55904 (I952920,I288688);
nor I_55905 (I952937,I952920,I288676);
not I_55906 (I952954,I288685);
nor I_55907 (I952971,I952937,I288670);
nor I_55908 (I952988,I952895,I952971);
DFFARX1 I_55909 (I952988,I2507,I952852,I952838,);
nor I_55910 (I953019,I288670,I288676);
nand I_55911 (I953036,I953019,I288688);
DFFARX1 I_55912 (I953036,I2507,I952852,I952841,);
nor I_55913 (I953067,I952954,I288670);
nand I_55914 (I953084,I953067,I288661);
nor I_55915 (I953101,I952878,I953084);
DFFARX1 I_55916 (I953101,I2507,I952852,I952817,);
not I_55917 (I953132,I953084);
nand I_55918 (I952829,I952895,I953132);
DFFARX1 I_55919 (I953084,I2507,I952852,I953172,);
not I_55920 (I953180,I953172);
not I_55921 (I953197,I288670);
not I_55922 (I953214,I288673);
nor I_55923 (I953231,I953214,I288685);
nor I_55924 (I952844,I953180,I953231);
nor I_55925 (I953262,I953214,I288682);
and I_55926 (I953279,I953262,I288664);
or I_55927 (I953296,I953279,I288679);
DFFARX1 I_55928 (I953296,I2507,I952852,I953322,);
nor I_55929 (I952832,I953322,I952878);
not I_55930 (I953344,I953322);
and I_55931 (I953361,I953344,I952878);
nor I_55932 (I952826,I952903,I953361);
nand I_55933 (I953392,I953344,I952954);
nor I_55934 (I952820,I953214,I953392);
nand I_55935 (I952823,I953344,I953132);
nand I_55936 (I953437,I952954,I288673);
nor I_55937 (I952835,I953197,I953437);
not I_55938 (I953498,I2514);
DFFARX1 I_55939 (I80683,I2507,I953498,I953524,);
DFFARX1 I_55940 (I80689,I2507,I953498,I953541,);
not I_55941 (I953549,I953541);
not I_55942 (I953566,I80707);
nor I_55943 (I953583,I953566,I80686);
not I_55944 (I953600,I80692);
nor I_55945 (I953617,I953583,I80698);
nor I_55946 (I953634,I953541,I953617);
DFFARX1 I_55947 (I953634,I2507,I953498,I953484,);
nor I_55948 (I953665,I80698,I80686);
nand I_55949 (I953682,I953665,I80707);
DFFARX1 I_55950 (I953682,I2507,I953498,I953487,);
nor I_55951 (I953713,I953600,I80698);
nand I_55952 (I953730,I953713,I80704);
nor I_55953 (I953747,I953524,I953730);
DFFARX1 I_55954 (I953747,I2507,I953498,I953463,);
not I_55955 (I953778,I953730);
nand I_55956 (I953475,I953541,I953778);
DFFARX1 I_55957 (I953730,I2507,I953498,I953818,);
not I_55958 (I953826,I953818);
not I_55959 (I953843,I80698);
not I_55960 (I953860,I80686);
nor I_55961 (I953877,I953860,I80692);
nor I_55962 (I953490,I953826,I953877);
nor I_55963 (I953908,I953860,I80695);
and I_55964 (I953925,I953908,I80683);
or I_55965 (I953942,I953925,I80701);
DFFARX1 I_55966 (I953942,I2507,I953498,I953968,);
nor I_55967 (I953478,I953968,I953524);
not I_55968 (I953990,I953968);
and I_55969 (I954007,I953990,I953524);
nor I_55970 (I953472,I953549,I954007);
nand I_55971 (I954038,I953990,I953600);
nor I_55972 (I953466,I953860,I954038);
nand I_55973 (I953469,I953990,I953778);
nand I_55974 (I954083,I953600,I80686);
nor I_55975 (I953481,I953843,I954083);
not I_55976 (I954144,I2514);
DFFARX1 I_55977 (I86480,I2507,I954144,I954170,);
DFFARX1 I_55978 (I86486,I2507,I954144,I954187,);
not I_55979 (I954195,I954187);
not I_55980 (I954212,I86504);
nor I_55981 (I954229,I954212,I86483);
not I_55982 (I954246,I86489);
nor I_55983 (I954263,I954229,I86495);
nor I_55984 (I954280,I954187,I954263);
DFFARX1 I_55985 (I954280,I2507,I954144,I954130,);
nor I_55986 (I954311,I86495,I86483);
nand I_55987 (I954328,I954311,I86504);
DFFARX1 I_55988 (I954328,I2507,I954144,I954133,);
nor I_55989 (I954359,I954246,I86495);
nand I_55990 (I954376,I954359,I86501);
nor I_55991 (I954393,I954170,I954376);
DFFARX1 I_55992 (I954393,I2507,I954144,I954109,);
not I_55993 (I954424,I954376);
nand I_55994 (I954121,I954187,I954424);
DFFARX1 I_55995 (I954376,I2507,I954144,I954464,);
not I_55996 (I954472,I954464);
not I_55997 (I954489,I86495);
not I_55998 (I954506,I86483);
nor I_55999 (I954523,I954506,I86489);
nor I_56000 (I954136,I954472,I954523);
nor I_56001 (I954554,I954506,I86492);
and I_56002 (I954571,I954554,I86480);
or I_56003 (I954588,I954571,I86498);
DFFARX1 I_56004 (I954588,I2507,I954144,I954614,);
nor I_56005 (I954124,I954614,I954170);
not I_56006 (I954636,I954614);
and I_56007 (I954653,I954636,I954170);
nor I_56008 (I954118,I954195,I954653);
nand I_56009 (I954684,I954636,I954246);
nor I_56010 (I954112,I954506,I954684);
nand I_56011 (I954115,I954636,I954424);
nand I_56012 (I954729,I954246,I86483);
nor I_56013 (I954127,I954489,I954729);
not I_56014 (I954790,I2514);
DFFARX1 I_56015 (I161541,I2507,I954790,I954816,);
DFFARX1 I_56016 (I161553,I2507,I954790,I954833,);
not I_56017 (I954841,I954833);
not I_56018 (I954858,I161559);
nor I_56019 (I954875,I954858,I161544);
not I_56020 (I954892,I161535);
nor I_56021 (I954909,I954875,I161556);
nor I_56022 (I954926,I954833,I954909);
DFFARX1 I_56023 (I954926,I2507,I954790,I954776,);
nor I_56024 (I954957,I161556,I161544);
nand I_56025 (I954974,I954957,I161559);
DFFARX1 I_56026 (I954974,I2507,I954790,I954779,);
nor I_56027 (I955005,I954892,I161556);
nand I_56028 (I955022,I955005,I161538);
nor I_56029 (I955039,I954816,I955022);
DFFARX1 I_56030 (I955039,I2507,I954790,I954755,);
not I_56031 (I955070,I955022);
nand I_56032 (I954767,I954833,I955070);
DFFARX1 I_56033 (I955022,I2507,I954790,I955110,);
not I_56034 (I955118,I955110);
not I_56035 (I955135,I161556);
not I_56036 (I955152,I161547);
nor I_56037 (I955169,I955152,I161535);
nor I_56038 (I954782,I955118,I955169);
nor I_56039 (I955200,I955152,I161550);
and I_56040 (I955217,I955200,I161538);
or I_56041 (I955234,I955217,I161535);
DFFARX1 I_56042 (I955234,I2507,I954790,I955260,);
nor I_56043 (I954770,I955260,I954816);
not I_56044 (I955282,I955260);
and I_56045 (I955299,I955282,I954816);
nor I_56046 (I954764,I954841,I955299);
nand I_56047 (I955330,I955282,I954892);
nor I_56048 (I954758,I955152,I955330);
nand I_56049 (I954761,I955282,I955070);
nand I_56050 (I955375,I954892,I161547);
nor I_56051 (I954773,I955135,I955375);
not I_56052 (I955436,I2514);
DFFARX1 I_56053 (I1323757,I2507,I955436,I955462,);
DFFARX1 I_56054 (I1323781,I2507,I955436,I955479,);
not I_56055 (I955487,I955479);
not I_56056 (I955504,I1323763);
nor I_56057 (I955521,I955504,I1323772);
not I_56058 (I955538,I1323757);
nor I_56059 (I955555,I955521,I1323778);
nor I_56060 (I955572,I955479,I955555);
DFFARX1 I_56061 (I955572,I2507,I955436,I955422,);
nor I_56062 (I955603,I1323778,I1323772);
nand I_56063 (I955620,I955603,I1323763);
DFFARX1 I_56064 (I955620,I2507,I955436,I955425,);
nor I_56065 (I955651,I955538,I1323778);
nand I_56066 (I955668,I955651,I1323775);
nor I_56067 (I955685,I955462,I955668);
DFFARX1 I_56068 (I955685,I2507,I955436,I955401,);
not I_56069 (I955716,I955668);
nand I_56070 (I955413,I955479,I955716);
DFFARX1 I_56071 (I955668,I2507,I955436,I955756,);
not I_56072 (I955764,I955756);
not I_56073 (I955781,I1323778);
not I_56074 (I955798,I1323769);
nor I_56075 (I955815,I955798,I1323757);
nor I_56076 (I955428,I955764,I955815);
nor I_56077 (I955846,I955798,I1323760);
and I_56078 (I955863,I955846,I1323784);
or I_56079 (I955880,I955863,I1323766);
DFFARX1 I_56080 (I955880,I2507,I955436,I955906,);
nor I_56081 (I955416,I955906,I955462);
not I_56082 (I955928,I955906);
and I_56083 (I955945,I955928,I955462);
nor I_56084 (I955410,I955487,I955945);
nand I_56085 (I955976,I955928,I955538);
nor I_56086 (I955404,I955798,I955976);
nand I_56087 (I955407,I955928,I955716);
nand I_56088 (I956021,I955538,I1323769);
nor I_56089 (I955419,I955781,I956021);
not I_56090 (I956082,I2514);
DFFARX1 I_56091 (I36415,I2507,I956082,I956108,);
DFFARX1 I_56092 (I36421,I2507,I956082,I956125,);
not I_56093 (I956133,I956125);
not I_56094 (I956150,I36415);
nor I_56095 (I956167,I956150,I36427);
not I_56096 (I956184,I36439);
nor I_56097 (I956201,I956167,I36433);
nor I_56098 (I956218,I956125,I956201);
DFFARX1 I_56099 (I956218,I2507,I956082,I956068,);
nor I_56100 (I956249,I36433,I36427);
nand I_56101 (I956266,I956249,I36415);
DFFARX1 I_56102 (I956266,I2507,I956082,I956071,);
nor I_56103 (I956297,I956184,I36433);
nand I_56104 (I956314,I956297,I36418);
nor I_56105 (I956331,I956108,I956314);
DFFARX1 I_56106 (I956331,I2507,I956082,I956047,);
not I_56107 (I956362,I956314);
nand I_56108 (I956059,I956125,I956362);
DFFARX1 I_56109 (I956314,I2507,I956082,I956402,);
not I_56110 (I956410,I956402);
not I_56111 (I956427,I36433);
not I_56112 (I956444,I36418);
nor I_56113 (I956461,I956444,I36439);
nor I_56114 (I956074,I956410,I956461);
nor I_56115 (I956492,I956444,I36436);
and I_56116 (I956509,I956492,I36430);
or I_56117 (I956526,I956509,I36424);
DFFARX1 I_56118 (I956526,I2507,I956082,I956552,);
nor I_56119 (I956062,I956552,I956108);
not I_56120 (I956574,I956552);
and I_56121 (I956591,I956574,I956108);
nor I_56122 (I956056,I956133,I956591);
nand I_56123 (I956622,I956574,I956184);
nor I_56124 (I956050,I956444,I956622);
nand I_56125 (I956053,I956574,I956362);
nand I_56126 (I956667,I956184,I36418);
nor I_56127 (I956065,I956427,I956667);
not I_56128 (I956728,I2514);
DFFARX1 I_56129 (I873399,I2507,I956728,I956754,);
DFFARX1 I_56130 (I873396,I2507,I956728,I956771,);
not I_56131 (I956779,I956771);
not I_56132 (I956796,I873396);
nor I_56133 (I956813,I956796,I873399);
not I_56134 (I956830,I873411);
nor I_56135 (I956847,I956813,I873405);
nor I_56136 (I956864,I956771,I956847);
DFFARX1 I_56137 (I956864,I2507,I956728,I956714,);
nor I_56138 (I956895,I873405,I873399);
nand I_56139 (I956912,I956895,I873396);
DFFARX1 I_56140 (I956912,I2507,I956728,I956717,);
nor I_56141 (I956943,I956830,I873405);
nand I_56142 (I956960,I956943,I873393);
nor I_56143 (I956977,I956754,I956960);
DFFARX1 I_56144 (I956977,I2507,I956728,I956693,);
not I_56145 (I957008,I956960);
nand I_56146 (I956705,I956771,I957008);
DFFARX1 I_56147 (I956960,I2507,I956728,I957048,);
not I_56148 (I957056,I957048);
not I_56149 (I957073,I873405);
not I_56150 (I957090,I873402);
nor I_56151 (I957107,I957090,I873411);
nor I_56152 (I956720,I957056,I957107);
nor I_56153 (I957138,I957090,I873408);
and I_56154 (I957155,I957138,I873414);
or I_56155 (I957172,I957155,I873393);
DFFARX1 I_56156 (I957172,I2507,I956728,I957198,);
nor I_56157 (I956708,I957198,I956754);
not I_56158 (I957220,I957198);
and I_56159 (I957237,I957220,I956754);
nor I_56160 (I956702,I956779,I957237);
nand I_56161 (I957268,I957220,I956830);
nor I_56162 (I956696,I957090,I957268);
nand I_56163 (I956699,I957220,I957008);
nand I_56164 (I957313,I956830,I873402);
nor I_56165 (I956711,I957073,I957313);
not I_56166 (I957374,I2514);
DFFARX1 I_56167 (I107033,I2507,I957374,I957400,);
DFFARX1 I_56168 (I107039,I2507,I957374,I957417,);
not I_56169 (I957425,I957417);
not I_56170 (I957442,I107057);
nor I_56171 (I957459,I957442,I107036);
not I_56172 (I957476,I107042);
nor I_56173 (I957493,I957459,I107048);
nor I_56174 (I957510,I957417,I957493);
DFFARX1 I_56175 (I957510,I2507,I957374,I957360,);
nor I_56176 (I957541,I107048,I107036);
nand I_56177 (I957558,I957541,I107057);
DFFARX1 I_56178 (I957558,I2507,I957374,I957363,);
nor I_56179 (I957589,I957476,I107048);
nand I_56180 (I957606,I957589,I107054);
nor I_56181 (I957623,I957400,I957606);
DFFARX1 I_56182 (I957623,I2507,I957374,I957339,);
not I_56183 (I957654,I957606);
nand I_56184 (I957351,I957417,I957654);
DFFARX1 I_56185 (I957606,I2507,I957374,I957694,);
not I_56186 (I957702,I957694);
not I_56187 (I957719,I107048);
not I_56188 (I957736,I107036);
nor I_56189 (I957753,I957736,I107042);
nor I_56190 (I957366,I957702,I957753);
nor I_56191 (I957784,I957736,I107045);
and I_56192 (I957801,I957784,I107033);
or I_56193 (I957818,I957801,I107051);
DFFARX1 I_56194 (I957818,I2507,I957374,I957844,);
nor I_56195 (I957354,I957844,I957400);
not I_56196 (I957866,I957844);
and I_56197 (I957883,I957866,I957400);
nor I_56198 (I957348,I957425,I957883);
nand I_56199 (I957914,I957866,I957476);
nor I_56200 (I957342,I957736,I957914);
nand I_56201 (I957345,I957866,I957654);
nand I_56202 (I957959,I957476,I107036);
nor I_56203 (I957357,I957719,I957959);
not I_56204 (I958020,I2514);
DFFARX1 I_56205 (I108614,I2507,I958020,I958046,);
DFFARX1 I_56206 (I108620,I2507,I958020,I958063,);
not I_56207 (I958071,I958063);
not I_56208 (I958088,I108638);
nor I_56209 (I958105,I958088,I108617);
not I_56210 (I958122,I108623);
nor I_56211 (I958139,I958105,I108629);
nor I_56212 (I958156,I958063,I958139);
DFFARX1 I_56213 (I958156,I2507,I958020,I958006,);
nor I_56214 (I958187,I108629,I108617);
nand I_56215 (I958204,I958187,I108638);
DFFARX1 I_56216 (I958204,I2507,I958020,I958009,);
nor I_56217 (I958235,I958122,I108629);
nand I_56218 (I958252,I958235,I108635);
nor I_56219 (I958269,I958046,I958252);
DFFARX1 I_56220 (I958269,I2507,I958020,I957985,);
not I_56221 (I958300,I958252);
nand I_56222 (I957997,I958063,I958300);
DFFARX1 I_56223 (I958252,I2507,I958020,I958340,);
not I_56224 (I958348,I958340);
not I_56225 (I958365,I108629);
not I_56226 (I958382,I108617);
nor I_56227 (I958399,I958382,I108623);
nor I_56228 (I958012,I958348,I958399);
nor I_56229 (I958430,I958382,I108626);
and I_56230 (I958447,I958430,I108614);
or I_56231 (I958464,I958447,I108632);
DFFARX1 I_56232 (I958464,I2507,I958020,I958490,);
nor I_56233 (I958000,I958490,I958046);
not I_56234 (I958512,I958490);
and I_56235 (I958529,I958512,I958046);
nor I_56236 (I957994,I958071,I958529);
nand I_56237 (I958560,I958512,I958122);
nor I_56238 (I957988,I958382,I958560);
nand I_56239 (I957991,I958512,I958300);
nand I_56240 (I958605,I958122,I108617);
nor I_56241 (I958003,I958365,I958605);
not I_56242 (I958666,I2514);
DFFARX1 I_56243 (I478965,I2507,I958666,I958692,);
DFFARX1 I_56244 (I478962,I2507,I958666,I958709,);
not I_56245 (I958717,I958709);
not I_56246 (I958734,I478977);
nor I_56247 (I958751,I958734,I478980);
not I_56248 (I958768,I478968);
nor I_56249 (I958785,I958751,I478974);
nor I_56250 (I958802,I958709,I958785);
DFFARX1 I_56251 (I958802,I2507,I958666,I958652,);
nor I_56252 (I958833,I478974,I478980);
nand I_56253 (I958850,I958833,I478977);
DFFARX1 I_56254 (I958850,I2507,I958666,I958655,);
nor I_56255 (I958881,I958768,I478974);
nand I_56256 (I958898,I958881,I478986);
nor I_56257 (I958915,I958692,I958898);
DFFARX1 I_56258 (I958915,I2507,I958666,I958631,);
not I_56259 (I958946,I958898);
nand I_56260 (I958643,I958709,I958946);
DFFARX1 I_56261 (I958898,I2507,I958666,I958986,);
not I_56262 (I958994,I958986);
not I_56263 (I959011,I478974);
not I_56264 (I959028,I478959);
nor I_56265 (I959045,I959028,I478968);
nor I_56266 (I958658,I958994,I959045);
nor I_56267 (I959076,I959028,I478971);
and I_56268 (I959093,I959076,I478959);
or I_56269 (I959110,I959093,I478983);
DFFARX1 I_56270 (I959110,I2507,I958666,I959136,);
nor I_56271 (I958646,I959136,I958692);
not I_56272 (I959158,I959136);
and I_56273 (I959175,I959158,I958692);
nor I_56274 (I958640,I958717,I959175);
nand I_56275 (I959206,I959158,I958768);
nor I_56276 (I958634,I959028,I959206);
nand I_56277 (I958637,I959158,I958946);
nand I_56278 (I959251,I958768,I478959);
nor I_56279 (I958649,I959011,I959251);
not I_56280 (I959312,I2514);
DFFARX1 I_56281 (I677542,I2507,I959312,I959338,);
DFFARX1 I_56282 (I677536,I2507,I959312,I959355,);
not I_56283 (I959363,I959355);
not I_56284 (I959380,I677551);
nor I_56285 (I959397,I959380,I677536);
not I_56286 (I959414,I677545);
nor I_56287 (I959431,I959397,I677554);
nor I_56288 (I959448,I959355,I959431);
DFFARX1 I_56289 (I959448,I2507,I959312,I959298,);
nor I_56290 (I959479,I677554,I677536);
nand I_56291 (I959496,I959479,I677551);
DFFARX1 I_56292 (I959496,I2507,I959312,I959301,);
nor I_56293 (I959527,I959414,I677554);
nand I_56294 (I959544,I959527,I677539);
nor I_56295 (I959561,I959338,I959544);
DFFARX1 I_56296 (I959561,I2507,I959312,I959277,);
not I_56297 (I959592,I959544);
nand I_56298 (I959289,I959355,I959592);
DFFARX1 I_56299 (I959544,I2507,I959312,I959632,);
not I_56300 (I959640,I959632);
not I_56301 (I959657,I677554);
not I_56302 (I959674,I677548);
nor I_56303 (I959691,I959674,I677545);
nor I_56304 (I959304,I959640,I959691);
nor I_56305 (I959722,I959674,I677557);
and I_56306 (I959739,I959722,I677560);
or I_56307 (I959756,I959739,I677539);
DFFARX1 I_56308 (I959756,I2507,I959312,I959782,);
nor I_56309 (I959292,I959782,I959338);
not I_56310 (I959804,I959782);
and I_56311 (I959821,I959804,I959338);
nor I_56312 (I959286,I959363,I959821);
nand I_56313 (I959852,I959804,I959414);
nor I_56314 (I959280,I959674,I959852);
nand I_56315 (I959283,I959804,I959592);
nand I_56316 (I959897,I959414,I677548);
nor I_56317 (I959295,I959657,I959897);
not I_56318 (I959958,I2514);
DFFARX1 I_56319 (I42739,I2507,I959958,I959984,);
DFFARX1 I_56320 (I42745,I2507,I959958,I960001,);
not I_56321 (I960009,I960001);
not I_56322 (I960026,I42739);
nor I_56323 (I960043,I960026,I42751);
not I_56324 (I960060,I42763);
nor I_56325 (I960077,I960043,I42757);
nor I_56326 (I960094,I960001,I960077);
DFFARX1 I_56327 (I960094,I2507,I959958,I959944,);
nor I_56328 (I960125,I42757,I42751);
nand I_56329 (I960142,I960125,I42739);
DFFARX1 I_56330 (I960142,I2507,I959958,I959947,);
nor I_56331 (I960173,I960060,I42757);
nand I_56332 (I960190,I960173,I42742);
nor I_56333 (I960207,I959984,I960190);
DFFARX1 I_56334 (I960207,I2507,I959958,I959923,);
not I_56335 (I960238,I960190);
nand I_56336 (I959935,I960001,I960238);
DFFARX1 I_56337 (I960190,I2507,I959958,I960278,);
not I_56338 (I960286,I960278);
not I_56339 (I960303,I42757);
not I_56340 (I960320,I42742);
nor I_56341 (I960337,I960320,I42763);
nor I_56342 (I959950,I960286,I960337);
nor I_56343 (I960368,I960320,I42760);
and I_56344 (I960385,I960368,I42754);
or I_56345 (I960402,I960385,I42748);
DFFARX1 I_56346 (I960402,I2507,I959958,I960428,);
nor I_56347 (I959938,I960428,I959984);
not I_56348 (I960450,I960428);
and I_56349 (I960467,I960450,I959984);
nor I_56350 (I959932,I960009,I960467);
nand I_56351 (I960498,I960450,I960060);
nor I_56352 (I959926,I960320,I960498);
nand I_56353 (I959929,I960450,I960238);
nand I_56354 (I960543,I960060,I42742);
nor I_56355 (I959941,I960303,I960543);
not I_56356 (I960604,I2514);
DFFARX1 I_56357 (I1376117,I2507,I960604,I960630,);
DFFARX1 I_56358 (I1376141,I2507,I960604,I960647,);
not I_56359 (I960655,I960647);
not I_56360 (I960672,I1376123);
nor I_56361 (I960689,I960672,I1376132);
not I_56362 (I960706,I1376117);
nor I_56363 (I960723,I960689,I1376138);
nor I_56364 (I960740,I960647,I960723);
DFFARX1 I_56365 (I960740,I2507,I960604,I960590,);
nor I_56366 (I960771,I1376138,I1376132);
nand I_56367 (I960788,I960771,I1376123);
DFFARX1 I_56368 (I960788,I2507,I960604,I960593,);
nor I_56369 (I960819,I960706,I1376138);
nand I_56370 (I960836,I960819,I1376135);
nor I_56371 (I960853,I960630,I960836);
DFFARX1 I_56372 (I960853,I2507,I960604,I960569,);
not I_56373 (I960884,I960836);
nand I_56374 (I960581,I960647,I960884);
DFFARX1 I_56375 (I960836,I2507,I960604,I960924,);
not I_56376 (I960932,I960924);
not I_56377 (I960949,I1376138);
not I_56378 (I960966,I1376129);
nor I_56379 (I960983,I960966,I1376117);
nor I_56380 (I960596,I960932,I960983);
nor I_56381 (I961014,I960966,I1376120);
and I_56382 (I961031,I961014,I1376144);
or I_56383 (I961048,I961031,I1376126);
DFFARX1 I_56384 (I961048,I2507,I960604,I961074,);
nor I_56385 (I960584,I961074,I960630);
not I_56386 (I961096,I961074);
and I_56387 (I961113,I961096,I960630);
nor I_56388 (I960578,I960655,I961113);
nand I_56389 (I961144,I961096,I960706);
nor I_56390 (I960572,I960966,I961144);
nand I_56391 (I960575,I961096,I960884);
nand I_56392 (I961189,I960706,I1376129);
nor I_56393 (I960587,I960949,I961189);
not I_56394 (I961250,I2514);
DFFARX1 I_56395 (I232346,I2507,I961250,I961276,);
DFFARX1 I_56396 (I232358,I2507,I961250,I961293,);
not I_56397 (I961301,I961293);
not I_56398 (I961318,I232364);
nor I_56399 (I961335,I961318,I232349);
not I_56400 (I961352,I232340);
nor I_56401 (I961369,I961335,I232361);
nor I_56402 (I961386,I961293,I961369);
DFFARX1 I_56403 (I961386,I2507,I961250,I961236,);
nor I_56404 (I961417,I232361,I232349);
nand I_56405 (I961434,I961417,I232364);
DFFARX1 I_56406 (I961434,I2507,I961250,I961239,);
nor I_56407 (I961465,I961352,I232361);
nand I_56408 (I961482,I961465,I232343);
nor I_56409 (I961499,I961276,I961482);
DFFARX1 I_56410 (I961499,I2507,I961250,I961215,);
not I_56411 (I961530,I961482);
nand I_56412 (I961227,I961293,I961530);
DFFARX1 I_56413 (I961482,I2507,I961250,I961570,);
not I_56414 (I961578,I961570);
not I_56415 (I961595,I232361);
not I_56416 (I961612,I232352);
nor I_56417 (I961629,I961612,I232340);
nor I_56418 (I961242,I961578,I961629);
nor I_56419 (I961660,I961612,I232355);
and I_56420 (I961677,I961660,I232343);
or I_56421 (I961694,I961677,I232340);
DFFARX1 I_56422 (I961694,I2507,I961250,I961720,);
nor I_56423 (I961230,I961720,I961276);
not I_56424 (I961742,I961720);
and I_56425 (I961759,I961742,I961276);
nor I_56426 (I961224,I961301,I961759);
nand I_56427 (I961790,I961742,I961352);
nor I_56428 (I961218,I961612,I961790);
nand I_56429 (I961221,I961742,I961530);
nand I_56430 (I961835,I961352,I232352);
nor I_56431 (I961233,I961595,I961835);
not I_56432 (I961896,I2514);
DFFARX1 I_56433 (I1338037,I2507,I961896,I961922,);
DFFARX1 I_56434 (I1338061,I2507,I961896,I961939,);
not I_56435 (I961947,I961939);
not I_56436 (I961964,I1338043);
nor I_56437 (I961981,I961964,I1338052);
not I_56438 (I961998,I1338037);
nor I_56439 (I962015,I961981,I1338058);
nor I_56440 (I962032,I961939,I962015);
DFFARX1 I_56441 (I962032,I2507,I961896,I961882,);
nor I_56442 (I962063,I1338058,I1338052);
nand I_56443 (I962080,I962063,I1338043);
DFFARX1 I_56444 (I962080,I2507,I961896,I961885,);
nor I_56445 (I962111,I961998,I1338058);
nand I_56446 (I962128,I962111,I1338055);
nor I_56447 (I962145,I961922,I962128);
DFFARX1 I_56448 (I962145,I2507,I961896,I961861,);
not I_56449 (I962176,I962128);
nand I_56450 (I961873,I961939,I962176);
DFFARX1 I_56451 (I962128,I2507,I961896,I962216,);
not I_56452 (I962224,I962216);
not I_56453 (I962241,I1338058);
not I_56454 (I962258,I1338049);
nor I_56455 (I962275,I962258,I1338037);
nor I_56456 (I961888,I962224,I962275);
nor I_56457 (I962306,I962258,I1338040);
and I_56458 (I962323,I962306,I1338064);
or I_56459 (I962340,I962323,I1338046);
DFFARX1 I_56460 (I962340,I2507,I961896,I962366,);
nor I_56461 (I961876,I962366,I961922);
not I_56462 (I962388,I962366);
and I_56463 (I962405,I962388,I961922);
nor I_56464 (I961870,I961947,I962405);
nand I_56465 (I962436,I962388,I961998);
nor I_56466 (I961864,I962258,I962436);
nand I_56467 (I961867,I962388,I962176);
nand I_56468 (I962481,I961998,I1338049);
nor I_56469 (I961879,I962241,I962481);
not I_56470 (I962542,I2514);
DFFARX1 I_56471 (I585637,I2507,I962542,I962568,);
DFFARX1 I_56472 (I585649,I2507,I962542,I962585,);
not I_56473 (I962593,I962585);
not I_56474 (I962610,I585658);
nor I_56475 (I962627,I962610,I585634);
not I_56476 (I962644,I585652);
nor I_56477 (I962661,I962627,I585646);
nor I_56478 (I962678,I962585,I962661);
DFFARX1 I_56479 (I962678,I2507,I962542,I962528,);
nor I_56480 (I962709,I585646,I585634);
nand I_56481 (I962726,I962709,I585658);
DFFARX1 I_56482 (I962726,I2507,I962542,I962531,);
nor I_56483 (I962757,I962644,I585646);
nand I_56484 (I962774,I962757,I585640);
nor I_56485 (I962791,I962568,I962774);
DFFARX1 I_56486 (I962791,I2507,I962542,I962507,);
not I_56487 (I962822,I962774);
nand I_56488 (I962519,I962585,I962822);
DFFARX1 I_56489 (I962774,I2507,I962542,I962862,);
not I_56490 (I962870,I962862);
not I_56491 (I962887,I585646);
not I_56492 (I962904,I585655);
nor I_56493 (I962921,I962904,I585652);
nor I_56494 (I962534,I962870,I962921);
nor I_56495 (I962952,I962904,I585637);
and I_56496 (I962969,I962952,I585634);
or I_56497 (I962986,I962969,I585643);
DFFARX1 I_56498 (I962986,I2507,I962542,I963012,);
nor I_56499 (I962522,I963012,I962568);
not I_56500 (I963034,I963012);
and I_56501 (I963051,I963034,I962568);
nor I_56502 (I962516,I962593,I963051);
nand I_56503 (I963082,I963034,I962644);
nor I_56504 (I962510,I962904,I963082);
nand I_56505 (I962513,I963034,I962822);
nand I_56506 (I963127,I962644,I585655);
nor I_56507 (I962525,I962887,I963127);
not I_56508 (I963188,I2514);
DFFARX1 I_56509 (I353482,I2507,I963188,I963214,);
DFFARX1 I_56510 (I353488,I2507,I963188,I963231,);
not I_56511 (I963239,I963231);
not I_56512 (I963256,I353509);
nor I_56513 (I963273,I963256,I353497);
not I_56514 (I963290,I353506);
nor I_56515 (I963307,I963273,I353491);
nor I_56516 (I963324,I963231,I963307);
DFFARX1 I_56517 (I963324,I2507,I963188,I963174,);
nor I_56518 (I963355,I353491,I353497);
nand I_56519 (I963372,I963355,I353509);
DFFARX1 I_56520 (I963372,I2507,I963188,I963177,);
nor I_56521 (I963403,I963290,I353491);
nand I_56522 (I963420,I963403,I353482);
nor I_56523 (I963437,I963214,I963420);
DFFARX1 I_56524 (I963437,I2507,I963188,I963153,);
not I_56525 (I963468,I963420);
nand I_56526 (I963165,I963231,I963468);
DFFARX1 I_56527 (I963420,I2507,I963188,I963508,);
not I_56528 (I963516,I963508);
not I_56529 (I963533,I353491);
not I_56530 (I963550,I353494);
nor I_56531 (I963567,I963550,I353506);
nor I_56532 (I963180,I963516,I963567);
nor I_56533 (I963598,I963550,I353503);
and I_56534 (I963615,I963598,I353485);
or I_56535 (I963632,I963615,I353500);
DFFARX1 I_56536 (I963632,I2507,I963188,I963658,);
nor I_56537 (I963168,I963658,I963214);
not I_56538 (I963680,I963658);
and I_56539 (I963697,I963680,I963214);
nor I_56540 (I963162,I963239,I963697);
nand I_56541 (I963728,I963680,I963290);
nor I_56542 (I963156,I963550,I963728);
nand I_56543 (I963159,I963680,I963468);
nand I_56544 (I963773,I963290,I353494);
nor I_56545 (I963171,I963533,I963773);
not I_56546 (I963834,I2514);
DFFARX1 I_56547 (I1305361,I2507,I963834,I963860,);
DFFARX1 I_56548 (I1305358,I2507,I963834,I963877,);
not I_56549 (I963885,I963877);
not I_56550 (I963902,I1305355);
nor I_56551 (I963919,I963902,I1305346);
not I_56552 (I963936,I1305367);
nor I_56553 (I963953,I963919,I1305346);
nor I_56554 (I963970,I963877,I963953);
DFFARX1 I_56555 (I963970,I2507,I963834,I963820,);
nor I_56556 (I964001,I1305346,I1305346);
nand I_56557 (I964018,I964001,I1305355);
DFFARX1 I_56558 (I964018,I2507,I963834,I963823,);
nor I_56559 (I964049,I963936,I1305346);
nand I_56560 (I964066,I964049,I1305370);
nor I_56561 (I964083,I963860,I964066);
DFFARX1 I_56562 (I964083,I2507,I963834,I963799,);
not I_56563 (I964114,I964066);
nand I_56564 (I963811,I963877,I964114);
DFFARX1 I_56565 (I964066,I2507,I963834,I964154,);
not I_56566 (I964162,I964154);
not I_56567 (I964179,I1305346);
not I_56568 (I964196,I1305349);
nor I_56569 (I964213,I964196,I1305367);
nor I_56570 (I963826,I964162,I964213);
nor I_56571 (I964244,I964196,I1305352);
and I_56572 (I964261,I964244,I1305373);
or I_56573 (I964278,I964261,I1305364);
DFFARX1 I_56574 (I964278,I2507,I963834,I964304,);
nor I_56575 (I963814,I964304,I963860);
not I_56576 (I964326,I964304);
and I_56577 (I964343,I964326,I963860);
nor I_56578 (I963808,I963885,I964343);
nand I_56579 (I964374,I964326,I963936);
nor I_56580 (I963802,I964196,I964374);
nand I_56581 (I963805,I964326,I964114);
nand I_56582 (I964419,I963936,I1305349);
nor I_56583 (I963817,I964179,I964419);
not I_56584 (I964480,I2514);
DFFARX1 I_56585 (I337145,I2507,I964480,I964506,);
DFFARX1 I_56586 (I337151,I2507,I964480,I964523,);
not I_56587 (I964531,I964523);
not I_56588 (I964548,I337172);
nor I_56589 (I964565,I964548,I337160);
not I_56590 (I964582,I337169);
nor I_56591 (I964599,I964565,I337154);
nor I_56592 (I964616,I964523,I964599);
DFFARX1 I_56593 (I964616,I2507,I964480,I964466,);
nor I_56594 (I964647,I337154,I337160);
nand I_56595 (I964664,I964647,I337172);
DFFARX1 I_56596 (I964664,I2507,I964480,I964469,);
nor I_56597 (I964695,I964582,I337154);
nand I_56598 (I964712,I964695,I337145);
nor I_56599 (I964729,I964506,I964712);
DFFARX1 I_56600 (I964729,I2507,I964480,I964445,);
not I_56601 (I964760,I964712);
nand I_56602 (I964457,I964523,I964760);
DFFARX1 I_56603 (I964712,I2507,I964480,I964800,);
not I_56604 (I964808,I964800);
not I_56605 (I964825,I337154);
not I_56606 (I964842,I337157);
nor I_56607 (I964859,I964842,I337169);
nor I_56608 (I964472,I964808,I964859);
nor I_56609 (I964890,I964842,I337166);
and I_56610 (I964907,I964890,I337148);
or I_56611 (I964924,I964907,I337163);
DFFARX1 I_56612 (I964924,I2507,I964480,I964950,);
nor I_56613 (I964460,I964950,I964506);
not I_56614 (I964972,I964950);
and I_56615 (I964989,I964972,I964506);
nor I_56616 (I964454,I964531,I964989);
nand I_56617 (I965020,I964972,I964582);
nor I_56618 (I964448,I964842,I965020);
nand I_56619 (I964451,I964972,I964760);
nand I_56620 (I965065,I964582,I337157);
nor I_56621 (I964463,I964825,I965065);
not I_56622 (I965126,I2514);
DFFARX1 I_56623 (I370873,I2507,I965126,I965152,);
DFFARX1 I_56624 (I370879,I2507,I965126,I965169,);
not I_56625 (I965177,I965169);
not I_56626 (I965194,I370900);
nor I_56627 (I965211,I965194,I370888);
not I_56628 (I965228,I370897);
nor I_56629 (I965245,I965211,I370882);
nor I_56630 (I965262,I965169,I965245);
DFFARX1 I_56631 (I965262,I2507,I965126,I965112,);
nor I_56632 (I965293,I370882,I370888);
nand I_56633 (I965310,I965293,I370900);
DFFARX1 I_56634 (I965310,I2507,I965126,I965115,);
nor I_56635 (I965341,I965228,I370882);
nand I_56636 (I965358,I965341,I370873);
nor I_56637 (I965375,I965152,I965358);
DFFARX1 I_56638 (I965375,I2507,I965126,I965091,);
not I_56639 (I965406,I965358);
nand I_56640 (I965103,I965169,I965406);
DFFARX1 I_56641 (I965358,I2507,I965126,I965446,);
not I_56642 (I965454,I965446);
not I_56643 (I965471,I370882);
not I_56644 (I965488,I370885);
nor I_56645 (I965505,I965488,I370897);
nor I_56646 (I965118,I965454,I965505);
nor I_56647 (I965536,I965488,I370894);
and I_56648 (I965553,I965536,I370876);
or I_56649 (I965570,I965553,I370891);
DFFARX1 I_56650 (I965570,I2507,I965126,I965596,);
nor I_56651 (I965106,I965596,I965152);
not I_56652 (I965618,I965596);
and I_56653 (I965635,I965618,I965152);
nor I_56654 (I965100,I965177,I965635);
nand I_56655 (I965666,I965618,I965228);
nor I_56656 (I965094,I965488,I965666);
nand I_56657 (I965097,I965618,I965406);
nand I_56658 (I965711,I965228,I370885);
nor I_56659 (I965109,I965471,I965711);
not I_56660 (I965772,I2514);
DFFARX1 I_56661 (I1221044,I2507,I965772,I965798,);
DFFARX1 I_56662 (I1221050,I2507,I965772,I965815,);
not I_56663 (I965823,I965815);
not I_56664 (I965840,I1221047);
nor I_56665 (I965857,I965840,I1221026);
not I_56666 (I965874,I1221029);
nor I_56667 (I965891,I965857,I1221035);
nor I_56668 (I965908,I965815,I965891);
DFFARX1 I_56669 (I965908,I2507,I965772,I965758,);
nor I_56670 (I965939,I1221035,I1221026);
nand I_56671 (I965956,I965939,I1221047);
DFFARX1 I_56672 (I965956,I2507,I965772,I965761,);
nor I_56673 (I965987,I965874,I1221035);
nand I_56674 (I966004,I965987,I1221029);
nor I_56675 (I966021,I965798,I966004);
DFFARX1 I_56676 (I966021,I2507,I965772,I965737,);
not I_56677 (I966052,I966004);
nand I_56678 (I965749,I965815,I966052);
DFFARX1 I_56679 (I966004,I2507,I965772,I966092,);
not I_56680 (I966100,I966092);
not I_56681 (I966117,I1221035);
not I_56682 (I966134,I1221038);
nor I_56683 (I966151,I966134,I1221029);
nor I_56684 (I965764,I966100,I966151);
nor I_56685 (I966182,I966134,I1221026);
and I_56686 (I966199,I966182,I1221032);
or I_56687 (I966216,I966199,I1221041);
DFFARX1 I_56688 (I966216,I2507,I965772,I966242,);
nor I_56689 (I965752,I966242,I965798);
not I_56690 (I966264,I966242);
and I_56691 (I966281,I966264,I965798);
nor I_56692 (I965746,I965823,I966281);
nand I_56693 (I966312,I966264,I965874);
nor I_56694 (I965740,I966134,I966312);
nand I_56695 (I965743,I966264,I966052);
nand I_56696 (I966357,I965874,I1221038);
nor I_56697 (I965755,I966117,I966357);
not I_56698 (I966418,I2514);
DFFARX1 I_56699 (I104398,I2507,I966418,I966444,);
DFFARX1 I_56700 (I104404,I2507,I966418,I966461,);
not I_56701 (I966469,I966461);
not I_56702 (I966486,I104422);
nor I_56703 (I966503,I966486,I104401);
not I_56704 (I966520,I104407);
nor I_56705 (I966537,I966503,I104413);
nor I_56706 (I966554,I966461,I966537);
DFFARX1 I_56707 (I966554,I2507,I966418,I966404,);
nor I_56708 (I966585,I104413,I104401);
nand I_56709 (I966602,I966585,I104422);
DFFARX1 I_56710 (I966602,I2507,I966418,I966407,);
nor I_56711 (I966633,I966520,I104413);
nand I_56712 (I966650,I966633,I104419);
nor I_56713 (I966667,I966444,I966650);
DFFARX1 I_56714 (I966667,I2507,I966418,I966383,);
not I_56715 (I966698,I966650);
nand I_56716 (I966395,I966461,I966698);
DFFARX1 I_56717 (I966650,I2507,I966418,I966738,);
not I_56718 (I966746,I966738);
not I_56719 (I966763,I104413);
not I_56720 (I966780,I104401);
nor I_56721 (I966797,I966780,I104407);
nor I_56722 (I966410,I966746,I966797);
nor I_56723 (I966828,I966780,I104410);
and I_56724 (I966845,I966828,I104398);
or I_56725 (I966862,I966845,I104416);
DFFARX1 I_56726 (I966862,I2507,I966418,I966888,);
nor I_56727 (I966398,I966888,I966444);
not I_56728 (I966910,I966888);
and I_56729 (I966927,I966910,I966444);
nor I_56730 (I966392,I966469,I966927);
nand I_56731 (I966958,I966910,I966520);
nor I_56732 (I966386,I966780,I966958);
nand I_56733 (I966389,I966910,I966698);
nand I_56734 (I967003,I966520,I104401);
nor I_56735 (I966401,I966763,I967003);
not I_56736 (I967064,I2514);
DFFARX1 I_56737 (I100709,I2507,I967064,I967090,);
DFFARX1 I_56738 (I100715,I2507,I967064,I967107,);
not I_56739 (I967115,I967107);
not I_56740 (I967132,I100733);
nor I_56741 (I967149,I967132,I100712);
not I_56742 (I967166,I100718);
nor I_56743 (I967183,I967149,I100724);
nor I_56744 (I967200,I967107,I967183);
DFFARX1 I_56745 (I967200,I2507,I967064,I967050,);
nor I_56746 (I967231,I100724,I100712);
nand I_56747 (I967248,I967231,I100733);
DFFARX1 I_56748 (I967248,I2507,I967064,I967053,);
nor I_56749 (I967279,I967166,I100724);
nand I_56750 (I967296,I967279,I100730);
nor I_56751 (I967313,I967090,I967296);
DFFARX1 I_56752 (I967313,I2507,I967064,I967029,);
not I_56753 (I967344,I967296);
nand I_56754 (I967041,I967107,I967344);
DFFARX1 I_56755 (I967296,I2507,I967064,I967384,);
not I_56756 (I967392,I967384);
not I_56757 (I967409,I100724);
not I_56758 (I967426,I100712);
nor I_56759 (I967443,I967426,I100718);
nor I_56760 (I967056,I967392,I967443);
nor I_56761 (I967474,I967426,I100721);
and I_56762 (I967491,I967474,I100709);
or I_56763 (I967508,I967491,I100727);
DFFARX1 I_56764 (I967508,I2507,I967064,I967534,);
nor I_56765 (I967044,I967534,I967090);
not I_56766 (I967556,I967534);
and I_56767 (I967573,I967556,I967090);
nor I_56768 (I967038,I967115,I967573);
nand I_56769 (I967604,I967556,I967166);
nor I_56770 (I967032,I967426,I967604);
nand I_56771 (I967035,I967556,I967344);
nand I_56772 (I967649,I967166,I100712);
nor I_56773 (I967047,I967409,I967649);
not I_56774 (I967710,I2514);
DFFARX1 I_56775 (I530387,I2507,I967710,I967736,);
DFFARX1 I_56776 (I530399,I2507,I967710,I967753,);
not I_56777 (I967761,I967753);
not I_56778 (I967778,I530384);
nor I_56779 (I967795,I967778,I530402);
not I_56780 (I967812,I530408);
nor I_56781 (I967829,I967795,I530390);
nor I_56782 (I967846,I967753,I967829);
DFFARX1 I_56783 (I967846,I2507,I967710,I967696,);
nor I_56784 (I967877,I530390,I530402);
nand I_56785 (I967894,I967877,I530384);
DFFARX1 I_56786 (I967894,I2507,I967710,I967699,);
nor I_56787 (I967925,I967812,I530390);
nand I_56788 (I967942,I967925,I530393);
nor I_56789 (I967959,I967736,I967942);
DFFARX1 I_56790 (I967959,I2507,I967710,I967675,);
not I_56791 (I967990,I967942);
nand I_56792 (I967687,I967753,I967990);
DFFARX1 I_56793 (I967942,I2507,I967710,I968030,);
not I_56794 (I968038,I968030);
not I_56795 (I968055,I530390);
not I_56796 (I968072,I530396);
nor I_56797 (I968089,I968072,I530408);
nor I_56798 (I967702,I968038,I968089);
nor I_56799 (I968120,I968072,I530405);
and I_56800 (I968137,I968120,I530384);
or I_56801 (I968154,I968137,I530387);
DFFARX1 I_56802 (I968154,I2507,I967710,I968180,);
nor I_56803 (I967690,I968180,I967736);
not I_56804 (I968202,I968180);
and I_56805 (I968219,I968202,I967736);
nor I_56806 (I967684,I967761,I968219);
nand I_56807 (I968250,I968202,I967812);
nor I_56808 (I967678,I968072,I968250);
nand I_56809 (I967681,I968202,I967990);
nand I_56810 (I968295,I967812,I530396);
nor I_56811 (I967693,I968055,I968295);
not I_56812 (I968356,I2514);
DFFARX1 I_56813 (I1203466,I2507,I968356,I968382,);
DFFARX1 I_56814 (I1203448,I2507,I968356,I968399,);
not I_56815 (I968407,I968399);
not I_56816 (I968424,I1203457);
nor I_56817 (I968441,I968424,I1203469);
not I_56818 (I968458,I1203451);
nor I_56819 (I968475,I968441,I1203460);
nor I_56820 (I968492,I968399,I968475);
DFFARX1 I_56821 (I968492,I2507,I968356,I968342,);
nor I_56822 (I968523,I1203460,I1203469);
nand I_56823 (I968540,I968523,I1203457);
DFFARX1 I_56824 (I968540,I2507,I968356,I968345,);
nor I_56825 (I968571,I968458,I1203460);
nand I_56826 (I968588,I968571,I1203472);
nor I_56827 (I968605,I968382,I968588);
DFFARX1 I_56828 (I968605,I2507,I968356,I968321,);
not I_56829 (I968636,I968588);
nand I_56830 (I968333,I968399,I968636);
DFFARX1 I_56831 (I968588,I2507,I968356,I968676,);
not I_56832 (I968684,I968676);
not I_56833 (I968701,I1203460);
not I_56834 (I968718,I1203448);
nor I_56835 (I968735,I968718,I1203451);
nor I_56836 (I968348,I968684,I968735);
nor I_56837 (I968766,I968718,I1203454);
and I_56838 (I968783,I968766,I1203463);
or I_56839 (I968800,I968783,I1203451);
DFFARX1 I_56840 (I968800,I2507,I968356,I968826,);
nor I_56841 (I968336,I968826,I968382);
not I_56842 (I968848,I968826);
and I_56843 (I968865,I968848,I968382);
nor I_56844 (I968330,I968407,I968865);
nand I_56845 (I968896,I968848,I968458);
nor I_56846 (I968324,I968718,I968896);
nand I_56847 (I968327,I968848,I968636);
nand I_56848 (I968941,I968458,I1203448);
nor I_56849 (I968339,I968701,I968941);
not I_56850 (I969002,I2514);
DFFARX1 I_56851 (I767710,I2507,I969002,I969028,);
DFFARX1 I_56852 (I767704,I2507,I969002,I969045,);
not I_56853 (I969053,I969045);
not I_56854 (I969070,I767719);
nor I_56855 (I969087,I969070,I767704);
not I_56856 (I969104,I767713);
nor I_56857 (I969121,I969087,I767722);
nor I_56858 (I969138,I969045,I969121);
DFFARX1 I_56859 (I969138,I2507,I969002,I968988,);
nor I_56860 (I969169,I767722,I767704);
nand I_56861 (I969186,I969169,I767719);
DFFARX1 I_56862 (I969186,I2507,I969002,I968991,);
nor I_56863 (I969217,I969104,I767722);
nand I_56864 (I969234,I969217,I767707);
nor I_56865 (I969251,I969028,I969234);
DFFARX1 I_56866 (I969251,I2507,I969002,I968967,);
not I_56867 (I969282,I969234);
nand I_56868 (I968979,I969045,I969282);
DFFARX1 I_56869 (I969234,I2507,I969002,I969322,);
not I_56870 (I969330,I969322);
not I_56871 (I969347,I767722);
not I_56872 (I969364,I767716);
nor I_56873 (I969381,I969364,I767713);
nor I_56874 (I968994,I969330,I969381);
nor I_56875 (I969412,I969364,I767725);
and I_56876 (I969429,I969412,I767728);
or I_56877 (I969446,I969429,I767707);
DFFARX1 I_56878 (I969446,I2507,I969002,I969472,);
nor I_56879 (I968982,I969472,I969028);
not I_56880 (I969494,I969472);
and I_56881 (I969511,I969494,I969028);
nor I_56882 (I968976,I969053,I969511);
nand I_56883 (I969542,I969494,I969104);
nor I_56884 (I968970,I969364,I969542);
nand I_56885 (I968973,I969494,I969282);
nand I_56886 (I969587,I969104,I767716);
nor I_56887 (I968985,I969347,I969587);
not I_56888 (I969648,I2514);
DFFARX1 I_56889 (I559049,I2507,I969648,I969674,);
DFFARX1 I_56890 (I559061,I2507,I969648,I969691,);
not I_56891 (I969699,I969691);
not I_56892 (I969716,I559070);
nor I_56893 (I969733,I969716,I559046);
not I_56894 (I969750,I559064);
nor I_56895 (I969767,I969733,I559058);
nor I_56896 (I969784,I969691,I969767);
DFFARX1 I_56897 (I969784,I2507,I969648,I969634,);
nor I_56898 (I969815,I559058,I559046);
nand I_56899 (I969832,I969815,I559070);
DFFARX1 I_56900 (I969832,I2507,I969648,I969637,);
nor I_56901 (I969863,I969750,I559058);
nand I_56902 (I969880,I969863,I559052);
nor I_56903 (I969897,I969674,I969880);
DFFARX1 I_56904 (I969897,I2507,I969648,I969613,);
not I_56905 (I969928,I969880);
nand I_56906 (I969625,I969691,I969928);
DFFARX1 I_56907 (I969880,I2507,I969648,I969968,);
not I_56908 (I969976,I969968);
not I_56909 (I969993,I559058);
not I_56910 (I970010,I559067);
nor I_56911 (I970027,I970010,I559064);
nor I_56912 (I969640,I969976,I970027);
nor I_56913 (I970058,I970010,I559049);
and I_56914 (I970075,I970058,I559046);
or I_56915 (I970092,I970075,I559055);
DFFARX1 I_56916 (I970092,I2507,I969648,I970118,);
nor I_56917 (I969628,I970118,I969674);
not I_56918 (I970140,I970118);
and I_56919 (I970157,I970140,I969674);
nor I_56920 (I969622,I969699,I970157);
nand I_56921 (I970188,I970140,I969750);
nor I_56922 (I969616,I970010,I970188);
nand I_56923 (I969619,I970140,I969928);
nand I_56924 (I970233,I969750,I559067);
nor I_56925 (I969631,I969993,I970233);
not I_56926 (I970294,I2514);
DFFARX1 I_56927 (I128640,I2507,I970294,I970320,);
DFFARX1 I_56928 (I128646,I2507,I970294,I970337,);
not I_56929 (I970345,I970337);
not I_56930 (I970362,I128664);
nor I_56931 (I970379,I970362,I128643);
not I_56932 (I970396,I128649);
nor I_56933 (I970413,I970379,I128655);
nor I_56934 (I970430,I970337,I970413);
DFFARX1 I_56935 (I970430,I2507,I970294,I970280,);
nor I_56936 (I970461,I128655,I128643);
nand I_56937 (I970478,I970461,I128664);
DFFARX1 I_56938 (I970478,I2507,I970294,I970283,);
nor I_56939 (I970509,I970396,I128655);
nand I_56940 (I970526,I970509,I128661);
nor I_56941 (I970543,I970320,I970526);
DFFARX1 I_56942 (I970543,I2507,I970294,I970259,);
not I_56943 (I970574,I970526);
nand I_56944 (I970271,I970337,I970574);
DFFARX1 I_56945 (I970526,I2507,I970294,I970614,);
not I_56946 (I970622,I970614);
not I_56947 (I970639,I128655);
not I_56948 (I970656,I128643);
nor I_56949 (I970673,I970656,I128649);
nor I_56950 (I970286,I970622,I970673);
nor I_56951 (I970704,I970656,I128652);
and I_56952 (I970721,I970704,I128640);
or I_56953 (I970738,I970721,I128658);
DFFARX1 I_56954 (I970738,I2507,I970294,I970764,);
nor I_56955 (I970274,I970764,I970320);
not I_56956 (I970786,I970764);
and I_56957 (I970803,I970786,I970320);
nor I_56958 (I970268,I970345,I970803);
nand I_56959 (I970834,I970786,I970396);
nor I_56960 (I970262,I970656,I970834);
nand I_56961 (I970265,I970786,I970574);
nand I_56962 (I970879,I970396,I128643);
nor I_56963 (I970277,I970639,I970879);
not I_56964 (I970940,I2514);
DFFARX1 I_56965 (I876561,I2507,I970940,I970966,);
DFFARX1 I_56966 (I876558,I2507,I970940,I970983,);
not I_56967 (I970991,I970983);
not I_56968 (I971008,I876558);
nor I_56969 (I971025,I971008,I876561);
not I_56970 (I971042,I876573);
nor I_56971 (I971059,I971025,I876567);
nor I_56972 (I971076,I970983,I971059);
DFFARX1 I_56973 (I971076,I2507,I970940,I970926,);
nor I_56974 (I971107,I876567,I876561);
nand I_56975 (I971124,I971107,I876558);
DFFARX1 I_56976 (I971124,I2507,I970940,I970929,);
nor I_56977 (I971155,I971042,I876567);
nand I_56978 (I971172,I971155,I876555);
nor I_56979 (I971189,I970966,I971172);
DFFARX1 I_56980 (I971189,I2507,I970940,I970905,);
not I_56981 (I971220,I971172);
nand I_56982 (I970917,I970983,I971220);
DFFARX1 I_56983 (I971172,I2507,I970940,I971260,);
not I_56984 (I971268,I971260);
not I_56985 (I971285,I876567);
not I_56986 (I971302,I876564);
nor I_56987 (I971319,I971302,I876573);
nor I_56988 (I970932,I971268,I971319);
nor I_56989 (I971350,I971302,I876570);
and I_56990 (I971367,I971350,I876576);
or I_56991 (I971384,I971367,I876555);
DFFARX1 I_56992 (I971384,I2507,I970940,I971410,);
nor I_56993 (I970920,I971410,I970966);
not I_56994 (I971432,I971410);
and I_56995 (I971449,I971432,I970966);
nor I_56996 (I970914,I970991,I971449);
nand I_56997 (I971480,I971432,I971042);
nor I_56998 (I970908,I971302,I971480);
nand I_56999 (I970911,I971432,I971220);
nand I_57000 (I971525,I971042,I876564);
nor I_57001 (I970923,I971285,I971525);
not I_57002 (I971586,I2514);
DFFARX1 I_57003 (I355063,I2507,I971586,I971612,);
DFFARX1 I_57004 (I355069,I2507,I971586,I971629,);
not I_57005 (I971637,I971629);
not I_57006 (I971654,I355090);
nor I_57007 (I971671,I971654,I355078);
not I_57008 (I971688,I355087);
nor I_57009 (I971705,I971671,I355072);
nor I_57010 (I971722,I971629,I971705);
DFFARX1 I_57011 (I971722,I2507,I971586,I971572,);
nor I_57012 (I971753,I355072,I355078);
nand I_57013 (I971770,I971753,I355090);
DFFARX1 I_57014 (I971770,I2507,I971586,I971575,);
nor I_57015 (I971801,I971688,I355072);
nand I_57016 (I971818,I971801,I355063);
nor I_57017 (I971835,I971612,I971818);
DFFARX1 I_57018 (I971835,I2507,I971586,I971551,);
not I_57019 (I971866,I971818);
nand I_57020 (I971563,I971629,I971866);
DFFARX1 I_57021 (I971818,I2507,I971586,I971906,);
not I_57022 (I971914,I971906);
not I_57023 (I971931,I355072);
not I_57024 (I971948,I355075);
nor I_57025 (I971965,I971948,I355087);
nor I_57026 (I971578,I971914,I971965);
nor I_57027 (I971996,I971948,I355084);
and I_57028 (I972013,I971996,I355066);
or I_57029 (I972030,I972013,I355081);
DFFARX1 I_57030 (I972030,I2507,I971586,I972056,);
nor I_57031 (I971566,I972056,I971612);
not I_57032 (I972078,I972056);
and I_57033 (I972095,I972078,I971612);
nor I_57034 (I971560,I971637,I972095);
nand I_57035 (I972126,I972078,I971688);
nor I_57036 (I971554,I971948,I972126);
nand I_57037 (I971557,I972078,I971866);
nand I_57038 (I972171,I971688,I355075);
nor I_57039 (I971569,I971931,I972171);
not I_57040 (I972232,I2514);
DFFARX1 I_57041 (I435989,I2507,I972232,I972258,);
DFFARX1 I_57042 (I435986,I2507,I972232,I972275,);
not I_57043 (I972283,I972275);
not I_57044 (I972300,I436001);
nor I_57045 (I972317,I972300,I436004);
not I_57046 (I972334,I435992);
nor I_57047 (I972351,I972317,I435998);
nor I_57048 (I972368,I972275,I972351);
DFFARX1 I_57049 (I972368,I2507,I972232,I972218,);
nor I_57050 (I972399,I435998,I436004);
nand I_57051 (I972416,I972399,I436001);
DFFARX1 I_57052 (I972416,I2507,I972232,I972221,);
nor I_57053 (I972447,I972334,I435998);
nand I_57054 (I972464,I972447,I436010);
nor I_57055 (I972481,I972258,I972464);
DFFARX1 I_57056 (I972481,I2507,I972232,I972197,);
not I_57057 (I972512,I972464);
nand I_57058 (I972209,I972275,I972512);
DFFARX1 I_57059 (I972464,I2507,I972232,I972552,);
not I_57060 (I972560,I972552);
not I_57061 (I972577,I435998);
not I_57062 (I972594,I435983);
nor I_57063 (I972611,I972594,I435992);
nor I_57064 (I972224,I972560,I972611);
nor I_57065 (I972642,I972594,I435995);
and I_57066 (I972659,I972642,I435983);
or I_57067 (I972676,I972659,I436007);
DFFARX1 I_57068 (I972676,I2507,I972232,I972702,);
nor I_57069 (I972212,I972702,I972258);
not I_57070 (I972724,I972702);
and I_57071 (I972741,I972724,I972258);
nor I_57072 (I972206,I972283,I972741);
nand I_57073 (I972772,I972724,I972334);
nor I_57074 (I972200,I972594,I972772);
nand I_57075 (I972203,I972724,I972512);
nand I_57076 (I972817,I972334,I435983);
nor I_57077 (I972215,I972577,I972817);
not I_57078 (I972878,I2514);
DFFARX1 I_57079 (I806470,I2507,I972878,I972904,);
DFFARX1 I_57080 (I806467,I2507,I972878,I972921,);
not I_57081 (I972929,I972921);
not I_57082 (I972946,I806467);
nor I_57083 (I972963,I972946,I806470);
not I_57084 (I972980,I806482);
nor I_57085 (I972997,I972963,I806476);
nor I_57086 (I973014,I972921,I972997);
DFFARX1 I_57087 (I973014,I2507,I972878,I972864,);
nor I_57088 (I973045,I806476,I806470);
nand I_57089 (I973062,I973045,I806467);
DFFARX1 I_57090 (I973062,I2507,I972878,I972867,);
nor I_57091 (I973093,I972980,I806476);
nand I_57092 (I973110,I973093,I806464);
nor I_57093 (I973127,I972904,I973110);
DFFARX1 I_57094 (I973127,I2507,I972878,I972843,);
not I_57095 (I973158,I973110);
nand I_57096 (I972855,I972921,I973158);
DFFARX1 I_57097 (I973110,I2507,I972878,I973198,);
not I_57098 (I973206,I973198);
not I_57099 (I973223,I806476);
not I_57100 (I973240,I806473);
nor I_57101 (I973257,I973240,I806482);
nor I_57102 (I972870,I973206,I973257);
nor I_57103 (I973288,I973240,I806479);
and I_57104 (I973305,I973288,I806485);
or I_57105 (I973322,I973305,I806464);
DFFARX1 I_57106 (I973322,I2507,I972878,I973348,);
nor I_57107 (I972858,I973348,I972904);
not I_57108 (I973370,I973348);
and I_57109 (I973387,I973370,I972904);
nor I_57110 (I972852,I972929,I973387);
nand I_57111 (I973418,I973370,I972980);
nor I_57112 (I972846,I973240,I973418);
nand I_57113 (I972849,I973370,I973158);
nand I_57114 (I973463,I972980,I806473);
nor I_57115 (I972861,I973223,I973463);
not I_57116 (I973524,I2514);
DFFARX1 I_57117 (I1026410,I2507,I973524,I973550,);
DFFARX1 I_57118 (I1026413,I2507,I973524,I973567,);
not I_57119 (I973575,I973567);
not I_57120 (I973592,I1026410);
nor I_57121 (I973609,I973592,I1026422);
not I_57122 (I973626,I1026431);
nor I_57123 (I973643,I973609,I1026419);
nor I_57124 (I973660,I973567,I973643);
DFFARX1 I_57125 (I973660,I2507,I973524,I973510,);
nor I_57126 (I973691,I1026419,I1026422);
nand I_57127 (I973708,I973691,I1026410);
DFFARX1 I_57128 (I973708,I2507,I973524,I973513,);
nor I_57129 (I973739,I973626,I1026419);
nand I_57130 (I973756,I973739,I1026425);
nor I_57131 (I973773,I973550,I973756);
DFFARX1 I_57132 (I973773,I2507,I973524,I973489,);
not I_57133 (I973804,I973756);
nand I_57134 (I973501,I973567,I973804);
DFFARX1 I_57135 (I973756,I2507,I973524,I973844,);
not I_57136 (I973852,I973844);
not I_57137 (I973869,I1026419);
not I_57138 (I973886,I1026416);
nor I_57139 (I973903,I973886,I1026431);
nor I_57140 (I973516,I973852,I973903);
nor I_57141 (I973934,I973886,I1026428);
and I_57142 (I973951,I973934,I1026416);
or I_57143 (I973968,I973951,I1026413);
DFFARX1 I_57144 (I973968,I2507,I973524,I973994,);
nor I_57145 (I973504,I973994,I973550);
not I_57146 (I974016,I973994);
and I_57147 (I974033,I974016,I973550);
nor I_57148 (I973498,I973575,I974033);
nand I_57149 (I974064,I974016,I973626);
nor I_57150 (I973492,I973886,I974064);
nand I_57151 (I973495,I974016,I973804);
nand I_57152 (I974109,I973626,I1026416);
nor I_57153 (I973507,I973869,I974109);
not I_57154 (I974170,I2514);
DFFARX1 I_57155 (I791714,I2507,I974170,I974196,);
DFFARX1 I_57156 (I791711,I2507,I974170,I974213,);
not I_57157 (I974221,I974213);
not I_57158 (I974238,I791711);
nor I_57159 (I974255,I974238,I791714);
not I_57160 (I974272,I791726);
nor I_57161 (I974289,I974255,I791720);
nor I_57162 (I974306,I974213,I974289);
DFFARX1 I_57163 (I974306,I2507,I974170,I974156,);
nor I_57164 (I974337,I791720,I791714);
nand I_57165 (I974354,I974337,I791711);
DFFARX1 I_57166 (I974354,I2507,I974170,I974159,);
nor I_57167 (I974385,I974272,I791720);
nand I_57168 (I974402,I974385,I791708);
nor I_57169 (I974419,I974196,I974402);
DFFARX1 I_57170 (I974419,I2507,I974170,I974135,);
not I_57171 (I974450,I974402);
nand I_57172 (I974147,I974213,I974450);
DFFARX1 I_57173 (I974402,I2507,I974170,I974490,);
not I_57174 (I974498,I974490);
not I_57175 (I974515,I791720);
not I_57176 (I974532,I791717);
nor I_57177 (I974549,I974532,I791726);
nor I_57178 (I974162,I974498,I974549);
nor I_57179 (I974580,I974532,I791723);
and I_57180 (I974597,I974580,I791729);
or I_57181 (I974614,I974597,I791708);
DFFARX1 I_57182 (I974614,I2507,I974170,I974640,);
nor I_57183 (I974150,I974640,I974196);
not I_57184 (I974662,I974640);
and I_57185 (I974679,I974662,I974196);
nor I_57186 (I974144,I974221,I974679);
nand I_57187 (I974710,I974662,I974272);
nor I_57188 (I974138,I974532,I974710);
nand I_57189 (I974141,I974662,I974450);
nand I_57190 (I974755,I974272,I791717);
nor I_57191 (I974153,I974515,I974755);
not I_57192 (I974816,I2514);
DFFARX1 I_57193 (I469173,I2507,I974816,I974842,);
DFFARX1 I_57194 (I469170,I2507,I974816,I974859,);
not I_57195 (I974867,I974859);
not I_57196 (I974884,I469185);
nor I_57197 (I974901,I974884,I469188);
not I_57198 (I974918,I469176);
nor I_57199 (I974935,I974901,I469182);
nor I_57200 (I974952,I974859,I974935);
DFFARX1 I_57201 (I974952,I2507,I974816,I974802,);
nor I_57202 (I974983,I469182,I469188);
nand I_57203 (I975000,I974983,I469185);
DFFARX1 I_57204 (I975000,I2507,I974816,I974805,);
nor I_57205 (I975031,I974918,I469182);
nand I_57206 (I975048,I975031,I469194);
nor I_57207 (I975065,I974842,I975048);
DFFARX1 I_57208 (I975065,I2507,I974816,I974781,);
not I_57209 (I975096,I975048);
nand I_57210 (I974793,I974859,I975096);
DFFARX1 I_57211 (I975048,I2507,I974816,I975136,);
not I_57212 (I975144,I975136);
not I_57213 (I975161,I469182);
not I_57214 (I975178,I469167);
nor I_57215 (I975195,I975178,I469176);
nor I_57216 (I974808,I975144,I975195);
nor I_57217 (I975226,I975178,I469179);
and I_57218 (I975243,I975226,I469167);
or I_57219 (I975260,I975243,I469191);
DFFARX1 I_57220 (I975260,I2507,I974816,I975286,);
nor I_57221 (I974796,I975286,I974842);
not I_57222 (I975308,I975286);
and I_57223 (I975325,I975308,I974842);
nor I_57224 (I974790,I974867,I975325);
nand I_57225 (I975356,I975308,I974918);
nor I_57226 (I974784,I975178,I975356);
nand I_57227 (I974787,I975308,I975096);
nand I_57228 (I975401,I974918,I469167);
nor I_57229 (I974799,I975161,I975401);
not I_57230 (I975462,I2514);
DFFARX1 I_57231 (I589683,I2507,I975462,I975488,);
DFFARX1 I_57232 (I589695,I2507,I975462,I975505,);
not I_57233 (I975513,I975505);
not I_57234 (I975530,I589704);
nor I_57235 (I975547,I975530,I589680);
not I_57236 (I975564,I589698);
nor I_57237 (I975581,I975547,I589692);
nor I_57238 (I975598,I975505,I975581);
DFFARX1 I_57239 (I975598,I2507,I975462,I975448,);
nor I_57240 (I975629,I589692,I589680);
nand I_57241 (I975646,I975629,I589704);
DFFARX1 I_57242 (I975646,I2507,I975462,I975451,);
nor I_57243 (I975677,I975564,I589692);
nand I_57244 (I975694,I975677,I589686);
nor I_57245 (I975711,I975488,I975694);
DFFARX1 I_57246 (I975711,I2507,I975462,I975427,);
not I_57247 (I975742,I975694);
nand I_57248 (I975439,I975505,I975742);
DFFARX1 I_57249 (I975694,I2507,I975462,I975782,);
not I_57250 (I975790,I975782);
not I_57251 (I975807,I589692);
not I_57252 (I975824,I589701);
nor I_57253 (I975841,I975824,I589698);
nor I_57254 (I975454,I975790,I975841);
nor I_57255 (I975872,I975824,I589683);
and I_57256 (I975889,I975872,I589680);
or I_57257 (I975906,I975889,I589689);
DFFARX1 I_57258 (I975906,I2507,I975462,I975932,);
nor I_57259 (I975442,I975932,I975488);
not I_57260 (I975954,I975932);
and I_57261 (I975971,I975954,I975488);
nor I_57262 (I975436,I975513,I975971);
nand I_57263 (I976002,I975954,I975564);
nor I_57264 (I975430,I975824,I976002);
nand I_57265 (I975433,I975954,I975742);
nand I_57266 (I976047,I975564,I589701);
nor I_57267 (I975445,I975807,I976047);
not I_57268 (I976108,I2514);
DFFARX1 I_57269 (I325551,I2507,I976108,I976134,);
DFFARX1 I_57270 (I325557,I2507,I976108,I976151,);
not I_57271 (I976159,I976151);
not I_57272 (I976176,I325578);
nor I_57273 (I976193,I976176,I325566);
not I_57274 (I976210,I325575);
nor I_57275 (I976227,I976193,I325560);
nor I_57276 (I976244,I976151,I976227);
DFFARX1 I_57277 (I976244,I2507,I976108,I976094,);
nor I_57278 (I976275,I325560,I325566);
nand I_57279 (I976292,I976275,I325578);
DFFARX1 I_57280 (I976292,I2507,I976108,I976097,);
nor I_57281 (I976323,I976210,I325560);
nand I_57282 (I976340,I976323,I325551);
nor I_57283 (I976357,I976134,I976340);
DFFARX1 I_57284 (I976357,I2507,I976108,I976073,);
not I_57285 (I976388,I976340);
nand I_57286 (I976085,I976151,I976388);
DFFARX1 I_57287 (I976340,I2507,I976108,I976428,);
not I_57288 (I976436,I976428);
not I_57289 (I976453,I325560);
not I_57290 (I976470,I325563);
nor I_57291 (I976487,I976470,I325575);
nor I_57292 (I976100,I976436,I976487);
nor I_57293 (I976518,I976470,I325572);
and I_57294 (I976535,I976518,I325554);
or I_57295 (I976552,I976535,I325569);
DFFARX1 I_57296 (I976552,I2507,I976108,I976578,);
nor I_57297 (I976088,I976578,I976134);
not I_57298 (I976600,I976578);
and I_57299 (I976617,I976600,I976134);
nor I_57300 (I976082,I976159,I976617);
nand I_57301 (I976648,I976600,I976210);
nor I_57302 (I976076,I976470,I976648);
nand I_57303 (I976079,I976600,I976388);
nand I_57304 (I976693,I976210,I325563);
nor I_57305 (I976091,I976453,I976693);
not I_57306 (I976754,I2514);
DFFARX1 I_57307 (I286026,I2507,I976754,I976780,);
DFFARX1 I_57308 (I286032,I2507,I976754,I976797,);
not I_57309 (I976805,I976797);
not I_57310 (I976822,I286053);
nor I_57311 (I976839,I976822,I286041);
not I_57312 (I976856,I286050);
nor I_57313 (I976873,I976839,I286035);
nor I_57314 (I976890,I976797,I976873);
DFFARX1 I_57315 (I976890,I2507,I976754,I976740,);
nor I_57316 (I976921,I286035,I286041);
nand I_57317 (I976938,I976921,I286053);
DFFARX1 I_57318 (I976938,I2507,I976754,I976743,);
nor I_57319 (I976969,I976856,I286035);
nand I_57320 (I976986,I976969,I286026);
nor I_57321 (I977003,I976780,I976986);
DFFARX1 I_57322 (I977003,I2507,I976754,I976719,);
not I_57323 (I977034,I976986);
nand I_57324 (I976731,I976797,I977034);
DFFARX1 I_57325 (I976986,I2507,I976754,I977074,);
not I_57326 (I977082,I977074);
not I_57327 (I977099,I286035);
not I_57328 (I977116,I286038);
nor I_57329 (I977133,I977116,I286050);
nor I_57330 (I976746,I977082,I977133);
nor I_57331 (I977164,I977116,I286047);
and I_57332 (I977181,I977164,I286029);
or I_57333 (I977198,I977181,I286044);
DFFARX1 I_57334 (I977198,I2507,I976754,I977224,);
nor I_57335 (I976734,I977224,I976780);
not I_57336 (I977246,I977224);
and I_57337 (I977263,I977246,I976780);
nor I_57338 (I976728,I976805,I977263);
nand I_57339 (I977294,I977246,I976856);
nor I_57340 (I976722,I977116,I977294);
nand I_57341 (I976725,I977246,I977034);
nand I_57342 (I977339,I976856,I286038);
nor I_57343 (I976737,I977099,I977339);
not I_57344 (I977400,I2514);
DFFARX1 I_57345 (I637660,I2507,I977400,I977426,);
DFFARX1 I_57346 (I637654,I2507,I977400,I977443,);
not I_57347 (I977451,I977443);
not I_57348 (I977468,I637669);
nor I_57349 (I977485,I977468,I637654);
not I_57350 (I977502,I637663);
nor I_57351 (I977519,I977485,I637672);
nor I_57352 (I977536,I977443,I977519);
DFFARX1 I_57353 (I977536,I2507,I977400,I977386,);
nor I_57354 (I977567,I637672,I637654);
nand I_57355 (I977584,I977567,I637669);
DFFARX1 I_57356 (I977584,I2507,I977400,I977389,);
nor I_57357 (I977615,I977502,I637672);
nand I_57358 (I977632,I977615,I637657);
nor I_57359 (I977649,I977426,I977632);
DFFARX1 I_57360 (I977649,I2507,I977400,I977365,);
not I_57361 (I977680,I977632);
nand I_57362 (I977377,I977443,I977680);
DFFARX1 I_57363 (I977632,I2507,I977400,I977720,);
not I_57364 (I977728,I977720);
not I_57365 (I977745,I637672);
not I_57366 (I977762,I637666);
nor I_57367 (I977779,I977762,I637663);
nor I_57368 (I977392,I977728,I977779);
nor I_57369 (I977810,I977762,I637675);
and I_57370 (I977827,I977810,I637678);
or I_57371 (I977844,I977827,I637657);
DFFARX1 I_57372 (I977844,I2507,I977400,I977870,);
nor I_57373 (I977380,I977870,I977426);
not I_57374 (I977892,I977870);
and I_57375 (I977909,I977892,I977426);
nor I_57376 (I977374,I977451,I977909);
nand I_57377 (I977940,I977892,I977502);
nor I_57378 (I977368,I977762,I977940);
nand I_57379 (I977371,I977892,I977680);
nand I_57380 (I977985,I977502,I637666);
nor I_57381 (I977383,I977745,I977985);
not I_57382 (I978046,I2514);
DFFARX1 I_57383 (I379957,I2507,I978046,I978072,);
DFFARX1 I_57384 (I379954,I2507,I978046,I978089,);
not I_57385 (I978097,I978089);
not I_57386 (I978114,I379969);
nor I_57387 (I978131,I978114,I379972);
not I_57388 (I978148,I379960);
nor I_57389 (I978165,I978131,I379966);
nor I_57390 (I978182,I978089,I978165);
DFFARX1 I_57391 (I978182,I2507,I978046,I978032,);
nor I_57392 (I978213,I379966,I379972);
nand I_57393 (I978230,I978213,I379969);
DFFARX1 I_57394 (I978230,I2507,I978046,I978035,);
nor I_57395 (I978261,I978148,I379966);
nand I_57396 (I978278,I978261,I379978);
nor I_57397 (I978295,I978072,I978278);
DFFARX1 I_57398 (I978295,I2507,I978046,I978011,);
not I_57399 (I978326,I978278);
nand I_57400 (I978023,I978089,I978326);
DFFARX1 I_57401 (I978278,I2507,I978046,I978366,);
not I_57402 (I978374,I978366);
not I_57403 (I978391,I379966);
not I_57404 (I978408,I379951);
nor I_57405 (I978425,I978408,I379960);
nor I_57406 (I978038,I978374,I978425);
nor I_57407 (I978456,I978408,I379963);
and I_57408 (I978473,I978456,I379951);
or I_57409 (I978490,I978473,I379975);
DFFARX1 I_57410 (I978490,I2507,I978046,I978516,);
nor I_57411 (I978026,I978516,I978072);
not I_57412 (I978538,I978516);
and I_57413 (I978555,I978538,I978072);
nor I_57414 (I978020,I978097,I978555);
nand I_57415 (I978586,I978538,I978148);
nor I_57416 (I978014,I978408,I978586);
nand I_57417 (I978017,I978538,I978326);
nand I_57418 (I978631,I978148,I379951);
nor I_57419 (I978029,I978391,I978631);
not I_57420 (I978692,I2514);
DFFARX1 I_57421 (I1156648,I2507,I978692,I978718,);
DFFARX1 I_57422 (I1156630,I2507,I978692,I978735,);
not I_57423 (I978743,I978735);
not I_57424 (I978760,I1156639);
nor I_57425 (I978777,I978760,I1156651);
not I_57426 (I978794,I1156633);
nor I_57427 (I978811,I978777,I1156642);
nor I_57428 (I978828,I978735,I978811);
DFFARX1 I_57429 (I978828,I2507,I978692,I978678,);
nor I_57430 (I978859,I1156642,I1156651);
nand I_57431 (I978876,I978859,I1156639);
DFFARX1 I_57432 (I978876,I2507,I978692,I978681,);
nor I_57433 (I978907,I978794,I1156642);
nand I_57434 (I978924,I978907,I1156654);
nor I_57435 (I978941,I978718,I978924);
DFFARX1 I_57436 (I978941,I2507,I978692,I978657,);
not I_57437 (I978972,I978924);
nand I_57438 (I978669,I978735,I978972);
DFFARX1 I_57439 (I978924,I2507,I978692,I979012,);
not I_57440 (I979020,I979012);
not I_57441 (I979037,I1156642);
not I_57442 (I979054,I1156630);
nor I_57443 (I979071,I979054,I1156633);
nor I_57444 (I978684,I979020,I979071);
nor I_57445 (I979102,I979054,I1156636);
and I_57446 (I979119,I979102,I1156645);
or I_57447 (I979136,I979119,I1156633);
DFFARX1 I_57448 (I979136,I2507,I978692,I979162,);
nor I_57449 (I978672,I979162,I978718);
not I_57450 (I979184,I979162);
and I_57451 (I979201,I979184,I978718);
nor I_57452 (I978666,I978743,I979201);
nand I_57453 (I979232,I979184,I978794);
nor I_57454 (I978660,I979054,I979232);
nand I_57455 (I978663,I979184,I978972);
nand I_57456 (I979277,I978794,I1156630);
nor I_57457 (I978675,I979037,I979277);
not I_57458 (I979338,I2514);
DFFARX1 I_57459 (I670028,I2507,I979338,I979364,);
DFFARX1 I_57460 (I670022,I2507,I979338,I979381,);
not I_57461 (I979389,I979381);
not I_57462 (I979406,I670037);
nor I_57463 (I979423,I979406,I670022);
not I_57464 (I979440,I670031);
nor I_57465 (I979457,I979423,I670040);
nor I_57466 (I979474,I979381,I979457);
DFFARX1 I_57467 (I979474,I2507,I979338,I979324,);
nor I_57468 (I979505,I670040,I670022);
nand I_57469 (I979522,I979505,I670037);
DFFARX1 I_57470 (I979522,I2507,I979338,I979327,);
nor I_57471 (I979553,I979440,I670040);
nand I_57472 (I979570,I979553,I670025);
nor I_57473 (I979587,I979364,I979570);
DFFARX1 I_57474 (I979587,I2507,I979338,I979303,);
not I_57475 (I979618,I979570);
nand I_57476 (I979315,I979381,I979618);
DFFARX1 I_57477 (I979570,I2507,I979338,I979658,);
not I_57478 (I979666,I979658);
not I_57479 (I979683,I670040);
not I_57480 (I979700,I670034);
nor I_57481 (I979717,I979700,I670031);
nor I_57482 (I979330,I979666,I979717);
nor I_57483 (I979748,I979700,I670043);
and I_57484 (I979765,I979748,I670046);
or I_57485 (I979782,I979765,I670025);
DFFARX1 I_57486 (I979782,I2507,I979338,I979808,);
nor I_57487 (I979318,I979808,I979364);
not I_57488 (I979830,I979808);
and I_57489 (I979847,I979830,I979364);
nor I_57490 (I979312,I979389,I979847);
nand I_57491 (I979878,I979830,I979440);
nor I_57492 (I979306,I979700,I979878);
nand I_57493 (I979309,I979830,I979618);
nand I_57494 (I979923,I979440,I670034);
nor I_57495 (I979321,I979683,I979923);
not I_57496 (I979984,I2514);
DFFARX1 I_57497 (I1388017,I2507,I979984,I980010,);
DFFARX1 I_57498 (I1388041,I2507,I979984,I980027,);
not I_57499 (I980035,I980027);
not I_57500 (I980052,I1388023);
nor I_57501 (I980069,I980052,I1388032);
not I_57502 (I980086,I1388017);
nor I_57503 (I980103,I980069,I1388038);
nor I_57504 (I980120,I980027,I980103);
DFFARX1 I_57505 (I980120,I2507,I979984,I979970,);
nor I_57506 (I980151,I1388038,I1388032);
nand I_57507 (I980168,I980151,I1388023);
DFFARX1 I_57508 (I980168,I2507,I979984,I979973,);
nor I_57509 (I980199,I980086,I1388038);
nand I_57510 (I980216,I980199,I1388035);
nor I_57511 (I980233,I980010,I980216);
DFFARX1 I_57512 (I980233,I2507,I979984,I979949,);
not I_57513 (I980264,I980216);
nand I_57514 (I979961,I980027,I980264);
DFFARX1 I_57515 (I980216,I2507,I979984,I980304,);
not I_57516 (I980312,I980304);
not I_57517 (I980329,I1388038);
not I_57518 (I980346,I1388029);
nor I_57519 (I980363,I980346,I1388017);
nor I_57520 (I979976,I980312,I980363);
nor I_57521 (I980394,I980346,I1388020);
and I_57522 (I980411,I980394,I1388044);
or I_57523 (I980428,I980411,I1388026);
DFFARX1 I_57524 (I980428,I2507,I979984,I980454,);
nor I_57525 (I979964,I980454,I980010);
not I_57526 (I980476,I980454);
and I_57527 (I980493,I980476,I980010);
nor I_57528 (I979958,I980035,I980493);
nand I_57529 (I980524,I980476,I980086);
nor I_57530 (I979952,I980346,I980524);
nand I_57531 (I979955,I980476,I980264);
nand I_57532 (I980569,I980086,I1388029);
nor I_57533 (I979967,I980329,I980569);
not I_57534 (I980630,I2514);
DFFARX1 I_57535 (I32199,I2507,I980630,I980656,);
DFFARX1 I_57536 (I32205,I2507,I980630,I980673,);
not I_57537 (I980681,I980673);
not I_57538 (I980698,I32199);
nor I_57539 (I980715,I980698,I32211);
not I_57540 (I980732,I32223);
nor I_57541 (I980749,I980715,I32217);
nor I_57542 (I980766,I980673,I980749);
DFFARX1 I_57543 (I980766,I2507,I980630,I980616,);
nor I_57544 (I980797,I32217,I32211);
nand I_57545 (I980814,I980797,I32199);
DFFARX1 I_57546 (I980814,I2507,I980630,I980619,);
nor I_57547 (I980845,I980732,I32217);
nand I_57548 (I980862,I980845,I32202);
nor I_57549 (I980879,I980656,I980862);
DFFARX1 I_57550 (I980879,I2507,I980630,I980595,);
not I_57551 (I980910,I980862);
nand I_57552 (I980607,I980673,I980910);
DFFARX1 I_57553 (I980862,I2507,I980630,I980950,);
not I_57554 (I980958,I980950);
not I_57555 (I980975,I32217);
not I_57556 (I980992,I32202);
nor I_57557 (I981009,I980992,I32223);
nor I_57558 (I980622,I980958,I981009);
nor I_57559 (I981040,I980992,I32220);
and I_57560 (I981057,I981040,I32214);
or I_57561 (I981074,I981057,I32208);
DFFARX1 I_57562 (I981074,I2507,I980630,I981100,);
nor I_57563 (I980610,I981100,I980656);
not I_57564 (I981122,I981100);
and I_57565 (I981139,I981122,I980656);
nor I_57566 (I980604,I980681,I981139);
nand I_57567 (I981170,I981122,I980732);
nor I_57568 (I980598,I980992,I981170);
nand I_57569 (I980601,I981122,I980910);
nand I_57570 (I981215,I980732,I32202);
nor I_57571 (I980613,I980975,I981215);
not I_57572 (I981276,I2514);
DFFARX1 I_57573 (I787498,I2507,I981276,I981302,);
DFFARX1 I_57574 (I787495,I2507,I981276,I981319,);
not I_57575 (I981327,I981319);
not I_57576 (I981344,I787495);
nor I_57577 (I981361,I981344,I787498);
not I_57578 (I981378,I787510);
nor I_57579 (I981395,I981361,I787504);
nor I_57580 (I981412,I981319,I981395);
DFFARX1 I_57581 (I981412,I2507,I981276,I981262,);
nor I_57582 (I981443,I787504,I787498);
nand I_57583 (I981460,I981443,I787495);
DFFARX1 I_57584 (I981460,I2507,I981276,I981265,);
nor I_57585 (I981491,I981378,I787504);
nand I_57586 (I981508,I981491,I787492);
nor I_57587 (I981525,I981302,I981508);
DFFARX1 I_57588 (I981525,I2507,I981276,I981241,);
not I_57589 (I981556,I981508);
nand I_57590 (I981253,I981319,I981556);
DFFARX1 I_57591 (I981508,I2507,I981276,I981596,);
not I_57592 (I981604,I981596);
not I_57593 (I981621,I787504);
not I_57594 (I981638,I787501);
nor I_57595 (I981655,I981638,I787510);
nor I_57596 (I981268,I981604,I981655);
nor I_57597 (I981686,I981638,I787507);
and I_57598 (I981703,I981686,I787513);
or I_57599 (I981720,I981703,I787492);
DFFARX1 I_57600 (I981720,I2507,I981276,I981746,);
nor I_57601 (I981256,I981746,I981302);
not I_57602 (I981768,I981746);
and I_57603 (I981785,I981768,I981302);
nor I_57604 (I981250,I981327,I981785);
nand I_57605 (I981816,I981768,I981378);
nor I_57606 (I981244,I981638,I981816);
nand I_57607 (I981247,I981768,I981556);
nand I_57608 (I981861,I981378,I787501);
nor I_57609 (I981259,I981621,I981861);
not I_57610 (I981922,I2514);
DFFARX1 I_57611 (I653844,I2507,I981922,I981948,);
DFFARX1 I_57612 (I653838,I2507,I981922,I981965,);
not I_57613 (I981973,I981965);
not I_57614 (I981990,I653853);
nor I_57615 (I982007,I981990,I653838);
not I_57616 (I982024,I653847);
nor I_57617 (I982041,I982007,I653856);
nor I_57618 (I982058,I981965,I982041);
DFFARX1 I_57619 (I982058,I2507,I981922,I981908,);
nor I_57620 (I982089,I653856,I653838);
nand I_57621 (I982106,I982089,I653853);
DFFARX1 I_57622 (I982106,I2507,I981922,I981911,);
nor I_57623 (I982137,I982024,I653856);
nand I_57624 (I982154,I982137,I653841);
nor I_57625 (I982171,I981948,I982154);
DFFARX1 I_57626 (I982171,I2507,I981922,I981887,);
not I_57627 (I982202,I982154);
nand I_57628 (I981899,I981965,I982202);
DFFARX1 I_57629 (I982154,I2507,I981922,I982242,);
not I_57630 (I982250,I982242);
not I_57631 (I982267,I653856);
not I_57632 (I982284,I653850);
nor I_57633 (I982301,I982284,I653847);
nor I_57634 (I981914,I982250,I982301);
nor I_57635 (I982332,I982284,I653859);
and I_57636 (I982349,I982332,I653862);
or I_57637 (I982366,I982349,I653841);
DFFARX1 I_57638 (I982366,I2507,I981922,I982392,);
nor I_57639 (I981902,I982392,I981948);
not I_57640 (I982414,I982392);
and I_57641 (I982431,I982414,I981948);
nor I_57642 (I981896,I981973,I982431);
nand I_57643 (I982462,I982414,I982024);
nor I_57644 (I981890,I982284,I982462);
nand I_57645 (I981893,I982414,I982202);
nand I_57646 (I982507,I982024,I653850);
nor I_57647 (I981905,I982267,I982507);
not I_57648 (I982568,I2514);
DFFARX1 I_57649 (I32726,I2507,I982568,I982594,);
DFFARX1 I_57650 (I32732,I2507,I982568,I982611,);
not I_57651 (I982619,I982611);
not I_57652 (I982636,I32726);
nor I_57653 (I982653,I982636,I32738);
not I_57654 (I982670,I32750);
nor I_57655 (I982687,I982653,I32744);
nor I_57656 (I982704,I982611,I982687);
DFFARX1 I_57657 (I982704,I2507,I982568,I982554,);
nor I_57658 (I982735,I32744,I32738);
nand I_57659 (I982752,I982735,I32726);
DFFARX1 I_57660 (I982752,I2507,I982568,I982557,);
nor I_57661 (I982783,I982670,I32744);
nand I_57662 (I982800,I982783,I32729);
nor I_57663 (I982817,I982594,I982800);
DFFARX1 I_57664 (I982817,I2507,I982568,I982533,);
not I_57665 (I982848,I982800);
nand I_57666 (I982545,I982611,I982848);
DFFARX1 I_57667 (I982800,I2507,I982568,I982888,);
not I_57668 (I982896,I982888);
not I_57669 (I982913,I32744);
not I_57670 (I982930,I32729);
nor I_57671 (I982947,I982930,I32750);
nor I_57672 (I982560,I982896,I982947);
nor I_57673 (I982978,I982930,I32747);
and I_57674 (I982995,I982978,I32741);
or I_57675 (I983012,I982995,I32735);
DFFARX1 I_57676 (I983012,I2507,I982568,I983038,);
nor I_57677 (I982548,I983038,I982594);
not I_57678 (I983060,I983038);
and I_57679 (I983077,I983060,I982594);
nor I_57680 (I982542,I982619,I983077);
nand I_57681 (I983108,I983060,I982670);
nor I_57682 (I982536,I982930,I983108);
nand I_57683 (I982539,I983060,I982848);
nand I_57684 (I983153,I982670,I32729);
nor I_57685 (I982551,I982913,I983153);
not I_57686 (I983214,I2514);
DFFARX1 I_57687 (I1212340,I2507,I983214,I983240,);
DFFARX1 I_57688 (I1212346,I2507,I983214,I983257,);
not I_57689 (I983265,I983257);
not I_57690 (I983282,I1212343);
nor I_57691 (I983299,I983282,I1212322);
not I_57692 (I983316,I1212325);
nor I_57693 (I983333,I983299,I1212331);
nor I_57694 (I983350,I983257,I983333);
DFFARX1 I_57695 (I983350,I2507,I983214,I983200,);
nor I_57696 (I983381,I1212331,I1212322);
nand I_57697 (I983398,I983381,I1212343);
DFFARX1 I_57698 (I983398,I2507,I983214,I983203,);
nor I_57699 (I983429,I983316,I1212331);
nand I_57700 (I983446,I983429,I1212325);
nor I_57701 (I983463,I983240,I983446);
DFFARX1 I_57702 (I983463,I2507,I983214,I983179,);
not I_57703 (I983494,I983446);
nand I_57704 (I983191,I983257,I983494);
DFFARX1 I_57705 (I983446,I2507,I983214,I983534,);
not I_57706 (I983542,I983534);
not I_57707 (I983559,I1212331);
not I_57708 (I983576,I1212334);
nor I_57709 (I983593,I983576,I1212325);
nor I_57710 (I983206,I983542,I983593);
nor I_57711 (I983624,I983576,I1212322);
and I_57712 (I983641,I983624,I1212328);
or I_57713 (I983658,I983641,I1212337);
DFFARX1 I_57714 (I983658,I2507,I983214,I983684,);
nor I_57715 (I983194,I983684,I983240);
not I_57716 (I983706,I983684);
and I_57717 (I983723,I983706,I983240);
nor I_57718 (I983188,I983265,I983723);
nand I_57719 (I983754,I983706,I983316);
nor I_57720 (I983182,I983576,I983754);
nand I_57721 (I983185,I983706,I983494);
nand I_57722 (I983799,I983316,I1212334);
nor I_57723 (I983197,I983559,I983799);
not I_57724 (I983860,I2514);
DFFARX1 I_57725 (I680432,I2507,I983860,I983886,);
DFFARX1 I_57726 (I680426,I2507,I983860,I983903,);
not I_57727 (I983911,I983903);
not I_57728 (I983928,I680441);
nor I_57729 (I983945,I983928,I680426);
not I_57730 (I983962,I680435);
nor I_57731 (I983979,I983945,I680444);
nor I_57732 (I983996,I983903,I983979);
DFFARX1 I_57733 (I983996,I2507,I983860,I983846,);
nor I_57734 (I984027,I680444,I680426);
nand I_57735 (I984044,I984027,I680441);
DFFARX1 I_57736 (I984044,I2507,I983860,I983849,);
nor I_57737 (I984075,I983962,I680444);
nand I_57738 (I984092,I984075,I680429);
nor I_57739 (I984109,I983886,I984092);
DFFARX1 I_57740 (I984109,I2507,I983860,I983825,);
not I_57741 (I984140,I984092);
nand I_57742 (I983837,I983903,I984140);
DFFARX1 I_57743 (I984092,I2507,I983860,I984180,);
not I_57744 (I984188,I984180);
not I_57745 (I984205,I680444);
not I_57746 (I984222,I680438);
nor I_57747 (I984239,I984222,I680435);
nor I_57748 (I983852,I984188,I984239);
nor I_57749 (I984270,I984222,I680447);
and I_57750 (I984287,I984270,I680450);
or I_57751 (I984304,I984287,I680429);
DFFARX1 I_57752 (I984304,I2507,I983860,I984330,);
nor I_57753 (I983840,I984330,I983886);
not I_57754 (I984352,I984330);
and I_57755 (I984369,I984352,I983886);
nor I_57756 (I983834,I983911,I984369);
nand I_57757 (I984400,I984352,I983962);
nor I_57758 (I983828,I984222,I984400);
nand I_57759 (I983831,I984352,I984140);
nand I_57760 (I984445,I983962,I680438);
nor I_57761 (I983843,I984205,I984445);
not I_57762 (I984506,I2514);
DFFARX1 I_57763 (I788025,I2507,I984506,I984532,);
DFFARX1 I_57764 (I788022,I2507,I984506,I984549,);
not I_57765 (I984557,I984549);
not I_57766 (I984574,I788022);
nor I_57767 (I984591,I984574,I788025);
not I_57768 (I984608,I788037);
nor I_57769 (I984625,I984591,I788031);
nor I_57770 (I984642,I984549,I984625);
DFFARX1 I_57771 (I984642,I2507,I984506,I984492,);
nor I_57772 (I984673,I788031,I788025);
nand I_57773 (I984690,I984673,I788022);
DFFARX1 I_57774 (I984690,I2507,I984506,I984495,);
nor I_57775 (I984721,I984608,I788031);
nand I_57776 (I984738,I984721,I788019);
nor I_57777 (I984755,I984532,I984738);
DFFARX1 I_57778 (I984755,I2507,I984506,I984471,);
not I_57779 (I984786,I984738);
nand I_57780 (I984483,I984549,I984786);
DFFARX1 I_57781 (I984738,I2507,I984506,I984826,);
not I_57782 (I984834,I984826);
not I_57783 (I984851,I788031);
not I_57784 (I984868,I788028);
nor I_57785 (I984885,I984868,I788037);
nor I_57786 (I984498,I984834,I984885);
nor I_57787 (I984916,I984868,I788034);
and I_57788 (I984933,I984916,I788040);
or I_57789 (I984950,I984933,I788019);
DFFARX1 I_57790 (I984950,I2507,I984506,I984976,);
nor I_57791 (I984486,I984976,I984532);
not I_57792 (I984998,I984976);
and I_57793 (I985015,I984998,I984532);
nor I_57794 (I984480,I984557,I985015);
nand I_57795 (I985046,I984998,I984608);
nor I_57796 (I984474,I984868,I985046);
nand I_57797 (I984477,I984998,I984786);
nand I_57798 (I985091,I984608,I788028);
nor I_57799 (I984489,I984851,I985091);
not I_57800 (I985152,I2514);
DFFARX1 I_57801 (I681010,I2507,I985152,I985178,);
DFFARX1 I_57802 (I681004,I2507,I985152,I985195,);
not I_57803 (I985203,I985195);
not I_57804 (I985220,I681019);
nor I_57805 (I985237,I985220,I681004);
not I_57806 (I985254,I681013);
nor I_57807 (I985271,I985237,I681022);
nor I_57808 (I985288,I985195,I985271);
DFFARX1 I_57809 (I985288,I2507,I985152,I985138,);
nor I_57810 (I985319,I681022,I681004);
nand I_57811 (I985336,I985319,I681019);
DFFARX1 I_57812 (I985336,I2507,I985152,I985141,);
nor I_57813 (I985367,I985254,I681022);
nand I_57814 (I985384,I985367,I681007);
nor I_57815 (I985401,I985178,I985384);
DFFARX1 I_57816 (I985401,I2507,I985152,I985117,);
not I_57817 (I985432,I985384);
nand I_57818 (I985129,I985195,I985432);
DFFARX1 I_57819 (I985384,I2507,I985152,I985472,);
not I_57820 (I985480,I985472);
not I_57821 (I985497,I681022);
not I_57822 (I985514,I681016);
nor I_57823 (I985531,I985514,I681013);
nor I_57824 (I985144,I985480,I985531);
nor I_57825 (I985562,I985514,I681025);
and I_57826 (I985579,I985562,I681028);
or I_57827 (I985596,I985579,I681007);
DFFARX1 I_57828 (I985596,I2507,I985152,I985622,);
nor I_57829 (I985132,I985622,I985178);
not I_57830 (I985644,I985622);
and I_57831 (I985661,I985644,I985178);
nor I_57832 (I985126,I985203,I985661);
nand I_57833 (I985692,I985644,I985254);
nor I_57834 (I985120,I985514,I985692);
nand I_57835 (I985123,I985644,I985432);
nand I_57836 (I985737,I985254,I681016);
nor I_57837 (I985135,I985497,I985737);
not I_57838 (I985798,I2514);
DFFARX1 I_57839 (I566563,I2507,I985798,I985824,);
DFFARX1 I_57840 (I566575,I2507,I985798,I985841,);
not I_57841 (I985849,I985841);
not I_57842 (I985866,I566584);
nor I_57843 (I985883,I985866,I566560);
not I_57844 (I985900,I566578);
nor I_57845 (I985917,I985883,I566572);
nor I_57846 (I985934,I985841,I985917);
DFFARX1 I_57847 (I985934,I2507,I985798,I985784,);
nor I_57848 (I985965,I566572,I566560);
nand I_57849 (I985982,I985965,I566584);
DFFARX1 I_57850 (I985982,I2507,I985798,I985787,);
nor I_57851 (I986013,I985900,I566572);
nand I_57852 (I986030,I986013,I566566);
nor I_57853 (I986047,I985824,I986030);
DFFARX1 I_57854 (I986047,I2507,I985798,I985763,);
not I_57855 (I986078,I986030);
nand I_57856 (I985775,I985841,I986078);
DFFARX1 I_57857 (I986030,I2507,I985798,I986118,);
not I_57858 (I986126,I986118);
not I_57859 (I986143,I566572);
not I_57860 (I986160,I566581);
nor I_57861 (I986177,I986160,I566578);
nor I_57862 (I985790,I986126,I986177);
nor I_57863 (I986208,I986160,I566563);
and I_57864 (I986225,I986208,I566560);
or I_57865 (I986242,I986225,I566569);
DFFARX1 I_57866 (I986242,I2507,I985798,I986268,);
nor I_57867 (I985778,I986268,I985824);
not I_57868 (I986290,I986268);
and I_57869 (I986307,I986290,I985824);
nor I_57870 (I985772,I985849,I986307);
nand I_57871 (I986338,I986290,I985900);
nor I_57872 (I985766,I986160,I986338);
nand I_57873 (I985769,I986290,I986078);
nand I_57874 (I986383,I985900,I566581);
nor I_57875 (I985781,I986143,I986383);
not I_57876 (I986444,I2514);
DFFARX1 I_57877 (I1109252,I2507,I986444,I986470,);
DFFARX1 I_57878 (I1109234,I2507,I986444,I986487,);
not I_57879 (I986495,I986487);
not I_57880 (I986512,I1109243);
nor I_57881 (I986529,I986512,I1109255);
not I_57882 (I986546,I1109237);
nor I_57883 (I986563,I986529,I1109246);
nor I_57884 (I986580,I986487,I986563);
DFFARX1 I_57885 (I986580,I2507,I986444,I986430,);
nor I_57886 (I986611,I1109246,I1109255);
nand I_57887 (I986628,I986611,I1109243);
DFFARX1 I_57888 (I986628,I2507,I986444,I986433,);
nor I_57889 (I986659,I986546,I1109246);
nand I_57890 (I986676,I986659,I1109258);
nor I_57891 (I986693,I986470,I986676);
DFFARX1 I_57892 (I986693,I2507,I986444,I986409,);
not I_57893 (I986724,I986676);
nand I_57894 (I986421,I986487,I986724);
DFFARX1 I_57895 (I986676,I2507,I986444,I986764,);
not I_57896 (I986772,I986764);
not I_57897 (I986789,I1109246);
not I_57898 (I986806,I1109234);
nor I_57899 (I986823,I986806,I1109237);
nor I_57900 (I986436,I986772,I986823);
nor I_57901 (I986854,I986806,I1109240);
and I_57902 (I986871,I986854,I1109249);
or I_57903 (I986888,I986871,I1109237);
DFFARX1 I_57904 (I986888,I2507,I986444,I986914,);
nor I_57905 (I986424,I986914,I986470);
not I_57906 (I986936,I986914);
and I_57907 (I986953,I986936,I986470);
nor I_57908 (I986418,I986495,I986953);
nand I_57909 (I986984,I986936,I986546);
nor I_57910 (I986412,I986806,I986984);
nand I_57911 (I986415,I986936,I986724);
nand I_57912 (I987029,I986546,I1109234);
nor I_57913 (I986427,I986789,I987029);
not I_57914 (I987090,I2514);
DFFARX1 I_57915 (I487125,I2507,I987090,I987116,);
DFFARX1 I_57916 (I487122,I2507,I987090,I987133,);
not I_57917 (I987141,I987133);
not I_57918 (I987158,I487137);
nor I_57919 (I987175,I987158,I487140);
not I_57920 (I987192,I487128);
nor I_57921 (I987209,I987175,I487134);
nor I_57922 (I987226,I987133,I987209);
DFFARX1 I_57923 (I987226,I2507,I987090,I987076,);
nor I_57924 (I987257,I487134,I487140);
nand I_57925 (I987274,I987257,I487137);
DFFARX1 I_57926 (I987274,I2507,I987090,I987079,);
nor I_57927 (I987305,I987192,I487134);
nand I_57928 (I987322,I987305,I487146);
nor I_57929 (I987339,I987116,I987322);
DFFARX1 I_57930 (I987339,I2507,I987090,I987055,);
not I_57931 (I987370,I987322);
nand I_57932 (I987067,I987133,I987370);
DFFARX1 I_57933 (I987322,I2507,I987090,I987410,);
not I_57934 (I987418,I987410);
not I_57935 (I987435,I487134);
not I_57936 (I987452,I487119);
nor I_57937 (I987469,I987452,I487128);
nor I_57938 (I987082,I987418,I987469);
nor I_57939 (I987500,I987452,I487131);
and I_57940 (I987517,I987500,I487119);
or I_57941 (I987534,I987517,I487143);
DFFARX1 I_57942 (I987534,I2507,I987090,I987560,);
nor I_57943 (I987070,I987560,I987116);
not I_57944 (I987582,I987560);
and I_57945 (I987599,I987582,I987116);
nor I_57946 (I987064,I987141,I987599);
nand I_57947 (I987630,I987582,I987192);
nor I_57948 (I987058,I987452,I987630);
nand I_57949 (I987061,I987582,I987370);
nand I_57950 (I987675,I987192,I487119);
nor I_57951 (I987073,I987435,I987675);
not I_57952 (I987736,I2514);
DFFARX1 I_57953 (I351374,I2507,I987736,I987762,);
DFFARX1 I_57954 (I351380,I2507,I987736,I987779,);
not I_57955 (I987787,I987779);
not I_57956 (I987804,I351401);
nor I_57957 (I987821,I987804,I351389);
not I_57958 (I987838,I351398);
nor I_57959 (I987855,I987821,I351383);
nor I_57960 (I987872,I987779,I987855);
DFFARX1 I_57961 (I987872,I2507,I987736,I987722,);
nor I_57962 (I987903,I351383,I351389);
nand I_57963 (I987920,I987903,I351401);
DFFARX1 I_57964 (I987920,I2507,I987736,I987725,);
nor I_57965 (I987951,I987838,I351383);
nand I_57966 (I987968,I987951,I351374);
nor I_57967 (I987985,I987762,I987968);
DFFARX1 I_57968 (I987985,I2507,I987736,I987701,);
not I_57969 (I988016,I987968);
nand I_57970 (I987713,I987779,I988016);
DFFARX1 I_57971 (I987968,I2507,I987736,I988056,);
not I_57972 (I988064,I988056);
not I_57973 (I988081,I351383);
not I_57974 (I988098,I351386);
nor I_57975 (I988115,I988098,I351398);
nor I_57976 (I987728,I988064,I988115);
nor I_57977 (I988146,I988098,I351395);
and I_57978 (I988163,I988146,I351377);
or I_57979 (I988180,I988163,I351392);
DFFARX1 I_57980 (I988180,I2507,I987736,I988206,);
nor I_57981 (I987716,I988206,I987762);
not I_57982 (I988228,I988206);
and I_57983 (I988245,I988228,I987762);
nor I_57984 (I987710,I987787,I988245);
nand I_57985 (I988276,I988228,I987838);
nor I_57986 (I987704,I988098,I988276);
nand I_57987 (I987707,I988228,I988016);
nand I_57988 (I988321,I987838,I351386);
nor I_57989 (I987719,I988081,I988321);
not I_57990 (I988382,I2514);
DFFARX1 I_57991 (I68562,I2507,I988382,I988408,);
DFFARX1 I_57992 (I68568,I2507,I988382,I988425,);
not I_57993 (I988433,I988425);
not I_57994 (I988450,I68586);
nor I_57995 (I988467,I988450,I68565);
not I_57996 (I988484,I68571);
nor I_57997 (I988501,I988467,I68577);
nor I_57998 (I988518,I988425,I988501);
DFFARX1 I_57999 (I988518,I2507,I988382,I988368,);
nor I_58000 (I988549,I68577,I68565);
nand I_58001 (I988566,I988549,I68586);
DFFARX1 I_58002 (I988566,I2507,I988382,I988371,);
nor I_58003 (I988597,I988484,I68577);
nand I_58004 (I988614,I988597,I68583);
nor I_58005 (I988631,I988408,I988614);
DFFARX1 I_58006 (I988631,I2507,I988382,I988347,);
not I_58007 (I988662,I988614);
nand I_58008 (I988359,I988425,I988662);
DFFARX1 I_58009 (I988614,I2507,I988382,I988702,);
not I_58010 (I988710,I988702);
not I_58011 (I988727,I68577);
not I_58012 (I988744,I68565);
nor I_58013 (I988761,I988744,I68571);
nor I_58014 (I988374,I988710,I988761);
nor I_58015 (I988792,I988744,I68574);
and I_58016 (I988809,I988792,I68562);
or I_58017 (I988826,I988809,I68580);
DFFARX1 I_58018 (I988826,I2507,I988382,I988852,);
nor I_58019 (I988362,I988852,I988408);
not I_58020 (I988874,I988852);
and I_58021 (I988891,I988874,I988408);
nor I_58022 (I988356,I988433,I988891);
nand I_58023 (I988922,I988874,I988484);
nor I_58024 (I988350,I988744,I988922);
nand I_58025 (I988353,I988874,I988662);
nand I_58026 (I988967,I988484,I68565);
nor I_58027 (I988365,I988727,I988967);
not I_58028 (I989028,I2514);
DFFARX1 I_58029 (I334510,I2507,I989028,I989054,);
DFFARX1 I_58030 (I334516,I2507,I989028,I989071,);
not I_58031 (I989079,I989071);
not I_58032 (I989096,I334537);
nor I_58033 (I989113,I989096,I334525);
not I_58034 (I989130,I334534);
nor I_58035 (I989147,I989113,I334519);
nor I_58036 (I989164,I989071,I989147);
DFFARX1 I_58037 (I989164,I2507,I989028,I989014,);
nor I_58038 (I989195,I334519,I334525);
nand I_58039 (I989212,I989195,I334537);
DFFARX1 I_58040 (I989212,I2507,I989028,I989017,);
nor I_58041 (I989243,I989130,I334519);
nand I_58042 (I989260,I989243,I334510);
nor I_58043 (I989277,I989054,I989260);
DFFARX1 I_58044 (I989277,I2507,I989028,I988993,);
not I_58045 (I989308,I989260);
nand I_58046 (I989005,I989071,I989308);
DFFARX1 I_58047 (I989260,I2507,I989028,I989348,);
not I_58048 (I989356,I989348);
not I_58049 (I989373,I334519);
not I_58050 (I989390,I334522);
nor I_58051 (I989407,I989390,I334534);
nor I_58052 (I989020,I989356,I989407);
nor I_58053 (I989438,I989390,I334531);
and I_58054 (I989455,I989438,I334513);
or I_58055 (I989472,I989455,I334528);
DFFARX1 I_58056 (I989472,I2507,I989028,I989498,);
nor I_58057 (I989008,I989498,I989054);
not I_58058 (I989520,I989498);
and I_58059 (I989537,I989520,I989054);
nor I_58060 (I989002,I989079,I989537);
nand I_58061 (I989568,I989520,I989130);
nor I_58062 (I988996,I989390,I989568);
nand I_58063 (I988999,I989520,I989308);
nand I_58064 (I989613,I989130,I334522);
nor I_58065 (I989011,I989373,I989613);
not I_58066 (I989674,I2514);
DFFARX1 I_58067 (I180581,I2507,I989674,I989700,);
DFFARX1 I_58068 (I180593,I2507,I989674,I989717,);
not I_58069 (I989725,I989717);
not I_58070 (I989742,I180599);
nor I_58071 (I989759,I989742,I180584);
not I_58072 (I989776,I180575);
nor I_58073 (I989793,I989759,I180596);
nor I_58074 (I989810,I989717,I989793);
DFFARX1 I_58075 (I989810,I2507,I989674,I989660,);
nor I_58076 (I989841,I180596,I180584);
nand I_58077 (I989858,I989841,I180599);
DFFARX1 I_58078 (I989858,I2507,I989674,I989663,);
nor I_58079 (I989889,I989776,I180596);
nand I_58080 (I989906,I989889,I180578);
nor I_58081 (I989923,I989700,I989906);
DFFARX1 I_58082 (I989923,I2507,I989674,I989639,);
not I_58083 (I989954,I989906);
nand I_58084 (I989651,I989717,I989954);
DFFARX1 I_58085 (I989906,I2507,I989674,I989994,);
not I_58086 (I990002,I989994);
not I_58087 (I990019,I180596);
not I_58088 (I990036,I180587);
nor I_58089 (I990053,I990036,I180575);
nor I_58090 (I989666,I990002,I990053);
nor I_58091 (I990084,I990036,I180590);
and I_58092 (I990101,I990084,I180578);
or I_58093 (I990118,I990101,I180575);
DFFARX1 I_58094 (I990118,I2507,I989674,I990144,);
nor I_58095 (I989654,I990144,I989700);
not I_58096 (I990166,I990144);
and I_58097 (I990183,I990166,I989700);
nor I_58098 (I989648,I989725,I990183);
nand I_58099 (I990214,I990166,I989776);
nor I_58100 (I989642,I990036,I990214);
nand I_58101 (I989645,I990166,I989954);
nand I_58102 (I990259,I989776,I180587);
nor I_58103 (I989657,I990019,I990259);
not I_58104 (I990320,I2514);
DFFARX1 I_58105 (I330294,I2507,I990320,I990346,);
DFFARX1 I_58106 (I330300,I2507,I990320,I990363,);
not I_58107 (I990371,I990363);
not I_58108 (I990388,I330321);
nor I_58109 (I990405,I990388,I330309);
not I_58110 (I990422,I330318);
nor I_58111 (I990439,I990405,I330303);
nor I_58112 (I990456,I990363,I990439);
DFFARX1 I_58113 (I990456,I2507,I990320,I990306,);
nor I_58114 (I990487,I330303,I330309);
nand I_58115 (I990504,I990487,I330321);
DFFARX1 I_58116 (I990504,I2507,I990320,I990309,);
nor I_58117 (I990535,I990422,I330303);
nand I_58118 (I990552,I990535,I330294);
nor I_58119 (I990569,I990346,I990552);
DFFARX1 I_58120 (I990569,I2507,I990320,I990285,);
not I_58121 (I990600,I990552);
nand I_58122 (I990297,I990363,I990600);
DFFARX1 I_58123 (I990552,I2507,I990320,I990640,);
not I_58124 (I990648,I990640);
not I_58125 (I990665,I330303);
not I_58126 (I990682,I330306);
nor I_58127 (I990699,I990682,I330318);
nor I_58128 (I990312,I990648,I990699);
nor I_58129 (I990730,I990682,I330315);
and I_58130 (I990747,I990730,I330297);
or I_58131 (I990764,I990747,I330312);
DFFARX1 I_58132 (I990764,I2507,I990320,I990790,);
nor I_58133 (I990300,I990790,I990346);
not I_58134 (I990812,I990790);
and I_58135 (I990829,I990812,I990346);
nor I_58136 (I990294,I990371,I990829);
nand I_58137 (I990860,I990812,I990422);
nor I_58138 (I990288,I990682,I990860);
nand I_58139 (I990291,I990812,I990600);
nand I_58140 (I990905,I990422,I330306);
nor I_58141 (I990303,I990665,I990905);
not I_58142 (I990966,I2514);
DFFARX1 I_58143 (I632458,I2507,I990966,I990992,);
DFFARX1 I_58144 (I632452,I2507,I990966,I991009,);
not I_58145 (I991017,I991009);
not I_58146 (I991034,I632467);
nor I_58147 (I991051,I991034,I632452);
not I_58148 (I991068,I632461);
nor I_58149 (I991085,I991051,I632470);
nor I_58150 (I991102,I991009,I991085);
DFFARX1 I_58151 (I991102,I2507,I990966,I990952,);
nor I_58152 (I991133,I632470,I632452);
nand I_58153 (I991150,I991133,I632467);
DFFARX1 I_58154 (I991150,I2507,I990966,I990955,);
nor I_58155 (I991181,I991068,I632470);
nand I_58156 (I991198,I991181,I632455);
nor I_58157 (I991215,I990992,I991198);
DFFARX1 I_58158 (I991215,I2507,I990966,I990931,);
not I_58159 (I991246,I991198);
nand I_58160 (I990943,I991009,I991246);
DFFARX1 I_58161 (I991198,I2507,I990966,I991286,);
not I_58162 (I991294,I991286);
not I_58163 (I991311,I632470);
not I_58164 (I991328,I632464);
nor I_58165 (I991345,I991328,I632461);
nor I_58166 (I990958,I991294,I991345);
nor I_58167 (I991376,I991328,I632473);
and I_58168 (I991393,I991376,I632476);
or I_58169 (I991410,I991393,I632455);
DFFARX1 I_58170 (I991410,I2507,I990966,I991436,);
nor I_58171 (I990946,I991436,I990992);
not I_58172 (I991458,I991436);
and I_58173 (I991475,I991458,I990992);
nor I_58174 (I990940,I991017,I991475);
nand I_58175 (I991506,I991458,I991068);
nor I_58176 (I990934,I991328,I991506);
nand I_58177 (I990937,I991458,I991246);
nand I_58178 (I991551,I991068,I632464);
nor I_58179 (I990949,I991311,I991551);
not I_58180 (I991612,I2514);
DFFARX1 I_58181 (I144893,I2507,I991612,I991638,);
DFFARX1 I_58182 (I144896,I2507,I991612,I991655,);
not I_58183 (I991663,I991655);
not I_58184 (I991680,I144881);
nor I_58185 (I991697,I991680,I144875);
not I_58186 (I991714,I144884);
nor I_58187 (I991731,I991697,I144899);
nor I_58188 (I991748,I991655,I991731);
DFFARX1 I_58189 (I991748,I2507,I991612,I991598,);
nor I_58190 (I991779,I144899,I144875);
nand I_58191 (I991796,I991779,I144881);
DFFARX1 I_58192 (I991796,I2507,I991612,I991601,);
nor I_58193 (I991827,I991714,I144899);
nand I_58194 (I991844,I991827,I144902);
nor I_58195 (I991861,I991638,I991844);
DFFARX1 I_58196 (I991861,I2507,I991612,I991577,);
not I_58197 (I991892,I991844);
nand I_58198 (I991589,I991655,I991892);
DFFARX1 I_58199 (I991844,I2507,I991612,I991932,);
not I_58200 (I991940,I991932);
not I_58201 (I991957,I144899);
not I_58202 (I991974,I144878);
nor I_58203 (I991991,I991974,I144884);
nor I_58204 (I991604,I991940,I991991);
nor I_58205 (I992022,I991974,I144887);
and I_58206 (I992039,I992022,I144875);
or I_58207 (I992056,I992039,I144890);
DFFARX1 I_58208 (I992056,I2507,I991612,I992082,);
nor I_58209 (I991592,I992082,I991638);
not I_58210 (I992104,I992082);
and I_58211 (I992121,I992104,I991638);
nor I_58212 (I991586,I991663,I992121);
nand I_58213 (I992152,I992104,I991714);
nor I_58214 (I991580,I991974,I992152);
nand I_58215 (I991583,I992104,I991892);
nand I_58216 (I992197,I991714,I144878);
nor I_58217 (I991595,I991957,I992197);
not I_58218 (I992258,I2514);
DFFARX1 I_58219 (I122843,I2507,I992258,I992284,);
DFFARX1 I_58220 (I122849,I2507,I992258,I992301,);
not I_58221 (I992309,I992301);
not I_58222 (I992326,I122867);
nor I_58223 (I992343,I992326,I122846);
not I_58224 (I992360,I122852);
nor I_58225 (I992377,I992343,I122858);
nor I_58226 (I992394,I992301,I992377);
DFFARX1 I_58227 (I992394,I2507,I992258,I992244,);
nor I_58228 (I992425,I122858,I122846);
nand I_58229 (I992442,I992425,I122867);
DFFARX1 I_58230 (I992442,I2507,I992258,I992247,);
nor I_58231 (I992473,I992360,I122858);
nand I_58232 (I992490,I992473,I122864);
nor I_58233 (I992507,I992284,I992490);
DFFARX1 I_58234 (I992507,I2507,I992258,I992223,);
not I_58235 (I992538,I992490);
nand I_58236 (I992235,I992301,I992538);
DFFARX1 I_58237 (I992490,I2507,I992258,I992578,);
not I_58238 (I992586,I992578);
not I_58239 (I992603,I122858);
not I_58240 (I992620,I122846);
nor I_58241 (I992637,I992620,I122852);
nor I_58242 (I992250,I992586,I992637);
nor I_58243 (I992668,I992620,I122855);
and I_58244 (I992685,I992668,I122843);
or I_58245 (I992702,I992685,I122861);
DFFARX1 I_58246 (I992702,I2507,I992258,I992728,);
nor I_58247 (I992238,I992728,I992284);
not I_58248 (I992750,I992728);
and I_58249 (I992767,I992750,I992284);
nor I_58250 (I992232,I992309,I992767);
nand I_58251 (I992798,I992750,I992360);
nor I_58252 (I992226,I992620,I992798);
nand I_58253 (I992229,I992750,I992538);
nand I_58254 (I992843,I992360,I122846);
nor I_58255 (I992241,I992603,I992843);
not I_58256 (I992904,I2514);
DFFARX1 I_58257 (I1191906,I2507,I992904,I992930,);
DFFARX1 I_58258 (I1191888,I2507,I992904,I992947,);
not I_58259 (I992955,I992947);
not I_58260 (I992972,I1191897);
nor I_58261 (I992989,I992972,I1191909);
not I_58262 (I993006,I1191891);
nor I_58263 (I993023,I992989,I1191900);
nor I_58264 (I993040,I992947,I993023);
DFFARX1 I_58265 (I993040,I2507,I992904,I992890,);
nor I_58266 (I993071,I1191900,I1191909);
nand I_58267 (I993088,I993071,I1191897);
DFFARX1 I_58268 (I993088,I2507,I992904,I992893,);
nor I_58269 (I993119,I993006,I1191900);
nand I_58270 (I993136,I993119,I1191912);
nor I_58271 (I993153,I992930,I993136);
DFFARX1 I_58272 (I993153,I2507,I992904,I992869,);
not I_58273 (I993184,I993136);
nand I_58274 (I992881,I992947,I993184);
DFFARX1 I_58275 (I993136,I2507,I992904,I993224,);
not I_58276 (I993232,I993224);
not I_58277 (I993249,I1191900);
not I_58278 (I993266,I1191888);
nor I_58279 (I993283,I993266,I1191891);
nor I_58280 (I992896,I993232,I993283);
nor I_58281 (I993314,I993266,I1191894);
and I_58282 (I993331,I993314,I1191903);
or I_58283 (I993348,I993331,I1191891);
DFFARX1 I_58284 (I993348,I2507,I992904,I993374,);
nor I_58285 (I992884,I993374,I992930);
not I_58286 (I993396,I993374);
and I_58287 (I993413,I993396,I992930);
nor I_58288 (I992878,I992955,I993413);
nand I_58289 (I993444,I993396,I993006);
nor I_58290 (I992872,I993266,I993444);
nand I_58291 (I992875,I993396,I993184);
nand I_58292 (I993489,I993006,I1191888);
nor I_58293 (I992887,I993249,I993489);
not I_58294 (I993550,I2514);
DFFARX1 I_58295 (I481141,I2507,I993550,I993576,);
DFFARX1 I_58296 (I481138,I2507,I993550,I993593,);
not I_58297 (I993601,I993593);
not I_58298 (I993618,I481153);
nor I_58299 (I993635,I993618,I481156);
not I_58300 (I993652,I481144);
nor I_58301 (I993669,I993635,I481150);
nor I_58302 (I993686,I993593,I993669);
DFFARX1 I_58303 (I993686,I2507,I993550,I993536,);
nor I_58304 (I993717,I481150,I481156);
nand I_58305 (I993734,I993717,I481153);
DFFARX1 I_58306 (I993734,I2507,I993550,I993539,);
nor I_58307 (I993765,I993652,I481150);
nand I_58308 (I993782,I993765,I481162);
nor I_58309 (I993799,I993576,I993782);
DFFARX1 I_58310 (I993799,I2507,I993550,I993515,);
not I_58311 (I993830,I993782);
nand I_58312 (I993527,I993593,I993830);
DFFARX1 I_58313 (I993782,I2507,I993550,I993870,);
not I_58314 (I993878,I993870);
not I_58315 (I993895,I481150);
not I_58316 (I993912,I481135);
nor I_58317 (I993929,I993912,I481144);
nor I_58318 (I993542,I993878,I993929);
nor I_58319 (I993960,I993912,I481147);
and I_58320 (I993977,I993960,I481135);
or I_58321 (I993994,I993977,I481159);
DFFARX1 I_58322 (I993994,I2507,I993550,I994020,);
nor I_58323 (I993530,I994020,I993576);
not I_58324 (I994042,I994020);
and I_58325 (I994059,I994042,I993576);
nor I_58326 (I993524,I993601,I994059);
nand I_58327 (I994090,I994042,I993652);
nor I_58328 (I993518,I993912,I994090);
nand I_58329 (I993521,I994042,I993830);
nand I_58330 (I994135,I993652,I481135);
nor I_58331 (I993533,I993895,I994135);
not I_58332 (I994196,I2514);
DFFARX1 I_58333 (I543443,I2507,I994196,I994222,);
DFFARX1 I_58334 (I543455,I2507,I994196,I994239,);
not I_58335 (I994247,I994239);
not I_58336 (I994264,I543464);
nor I_58337 (I994281,I994264,I543440);
not I_58338 (I994298,I543458);
nor I_58339 (I994315,I994281,I543452);
nor I_58340 (I994332,I994239,I994315);
DFFARX1 I_58341 (I994332,I2507,I994196,I994182,);
nor I_58342 (I994363,I543452,I543440);
nand I_58343 (I994380,I994363,I543464);
DFFARX1 I_58344 (I994380,I2507,I994196,I994185,);
nor I_58345 (I994411,I994298,I543452);
nand I_58346 (I994428,I994411,I543446);
nor I_58347 (I994445,I994222,I994428);
DFFARX1 I_58348 (I994445,I2507,I994196,I994161,);
not I_58349 (I994476,I994428);
nand I_58350 (I994173,I994239,I994476);
DFFARX1 I_58351 (I994428,I2507,I994196,I994516,);
not I_58352 (I994524,I994516);
not I_58353 (I994541,I543452);
not I_58354 (I994558,I543461);
nor I_58355 (I994575,I994558,I543458);
nor I_58356 (I994188,I994524,I994575);
nor I_58357 (I994606,I994558,I543443);
and I_58358 (I994623,I994606,I543440);
or I_58359 (I994640,I994623,I543449);
DFFARX1 I_58360 (I994640,I2507,I994196,I994666,);
nor I_58361 (I994176,I994666,I994222);
not I_58362 (I994688,I994666);
and I_58363 (I994705,I994688,I994222);
nor I_58364 (I994170,I994247,I994705);
nand I_58365 (I994736,I994688,I994298);
nor I_58366 (I994164,I994558,I994736);
nand I_58367 (I994167,I994688,I994476);
nand I_58368 (I994781,I994298,I543461);
nor I_58369 (I994179,I994541,I994781);
not I_58370 (I994842,I2514);
DFFARX1 I_58371 (I1073994,I2507,I994842,I994868,);
DFFARX1 I_58372 (I1073976,I2507,I994842,I994885,);
not I_58373 (I994893,I994885);
not I_58374 (I994910,I1073985);
nor I_58375 (I994927,I994910,I1073997);
not I_58376 (I994944,I1073979);
nor I_58377 (I994961,I994927,I1073988);
nor I_58378 (I994978,I994885,I994961);
DFFARX1 I_58379 (I994978,I2507,I994842,I994828,);
nor I_58380 (I995009,I1073988,I1073997);
nand I_58381 (I995026,I995009,I1073985);
DFFARX1 I_58382 (I995026,I2507,I994842,I994831,);
nor I_58383 (I995057,I994944,I1073988);
nand I_58384 (I995074,I995057,I1074000);
nor I_58385 (I995091,I994868,I995074);
DFFARX1 I_58386 (I995091,I2507,I994842,I994807,);
not I_58387 (I995122,I995074);
nand I_58388 (I994819,I994885,I995122);
DFFARX1 I_58389 (I995074,I2507,I994842,I995162,);
not I_58390 (I995170,I995162);
not I_58391 (I995187,I1073988);
not I_58392 (I995204,I1073976);
nor I_58393 (I995221,I995204,I1073979);
nor I_58394 (I994834,I995170,I995221);
nor I_58395 (I995252,I995204,I1073982);
and I_58396 (I995269,I995252,I1073991);
or I_58397 (I995286,I995269,I1073979);
DFFARX1 I_58398 (I995286,I2507,I994842,I995312,);
nor I_58399 (I994822,I995312,I994868);
not I_58400 (I995334,I995312);
and I_58401 (I995351,I995334,I994868);
nor I_58402 (I994816,I994893,I995351);
nand I_58403 (I995382,I995334,I994944);
nor I_58404 (I994810,I995204,I995382);
nand I_58405 (I994813,I995334,I995122);
nand I_58406 (I995427,I994944,I1073976);
nor I_58407 (I994825,I995187,I995427);
not I_58408 (I995488,I2514);
DFFARX1 I_58409 (I238296,I2507,I995488,I995514,);
DFFARX1 I_58410 (I238308,I2507,I995488,I995531,);
not I_58411 (I995539,I995531);
not I_58412 (I995556,I238314);
nor I_58413 (I995573,I995556,I238299);
not I_58414 (I995590,I238290);
nor I_58415 (I995607,I995573,I238311);
nor I_58416 (I995624,I995531,I995607);
DFFARX1 I_58417 (I995624,I2507,I995488,I995474,);
nor I_58418 (I995655,I238311,I238299);
nand I_58419 (I995672,I995655,I238314);
DFFARX1 I_58420 (I995672,I2507,I995488,I995477,);
nor I_58421 (I995703,I995590,I238311);
nand I_58422 (I995720,I995703,I238293);
nor I_58423 (I995737,I995514,I995720);
DFFARX1 I_58424 (I995737,I2507,I995488,I995453,);
not I_58425 (I995768,I995720);
nand I_58426 (I995465,I995531,I995768);
DFFARX1 I_58427 (I995720,I2507,I995488,I995808,);
not I_58428 (I995816,I995808);
not I_58429 (I995833,I238311);
not I_58430 (I995850,I238302);
nor I_58431 (I995867,I995850,I238290);
nor I_58432 (I995480,I995816,I995867);
nor I_58433 (I995898,I995850,I238305);
and I_58434 (I995915,I995898,I238293);
or I_58435 (I995932,I995915,I238290);
DFFARX1 I_58436 (I995932,I2507,I995488,I995958,);
nor I_58437 (I995468,I995958,I995514);
not I_58438 (I995980,I995958);
and I_58439 (I995997,I995980,I995514);
nor I_58440 (I995462,I995539,I995997);
nand I_58441 (I996028,I995980,I995590);
nor I_58442 (I995456,I995850,I996028);
nand I_58443 (I995459,I995980,I995768);
nand I_58444 (I996073,I995590,I238302);
nor I_58445 (I995471,I995833,I996073);
not I_58446 (I996134,I2514);
DFFARX1 I_58447 (I469717,I2507,I996134,I996160,);
DFFARX1 I_58448 (I469714,I2507,I996134,I996177,);
not I_58449 (I996185,I996177);
not I_58450 (I996202,I469729);
nor I_58451 (I996219,I996202,I469732);
not I_58452 (I996236,I469720);
nor I_58453 (I996253,I996219,I469726);
nor I_58454 (I996270,I996177,I996253);
DFFARX1 I_58455 (I996270,I2507,I996134,I996120,);
nor I_58456 (I996301,I469726,I469732);
nand I_58457 (I996318,I996301,I469729);
DFFARX1 I_58458 (I996318,I2507,I996134,I996123,);
nor I_58459 (I996349,I996236,I469726);
nand I_58460 (I996366,I996349,I469738);
nor I_58461 (I996383,I996160,I996366);
DFFARX1 I_58462 (I996383,I2507,I996134,I996099,);
not I_58463 (I996414,I996366);
nand I_58464 (I996111,I996177,I996414);
DFFARX1 I_58465 (I996366,I2507,I996134,I996454,);
not I_58466 (I996462,I996454);
not I_58467 (I996479,I469726);
not I_58468 (I996496,I469711);
nor I_58469 (I996513,I996496,I469720);
nor I_58470 (I996126,I996462,I996513);
nor I_58471 (I996544,I996496,I469723);
and I_58472 (I996561,I996544,I469711);
or I_58473 (I996578,I996561,I469735);
DFFARX1 I_58474 (I996578,I2507,I996134,I996604,);
nor I_58475 (I996114,I996604,I996160);
not I_58476 (I996626,I996604);
and I_58477 (I996643,I996626,I996160);
nor I_58478 (I996108,I996185,I996643);
nand I_58479 (I996674,I996626,I996236);
nor I_58480 (I996102,I996496,I996674);
nand I_58481 (I996105,I996626,I996414);
nand I_58482 (I996719,I996236,I469711);
nor I_58483 (I996117,I996479,I996719);
not I_58484 (I996780,I2514);
DFFARX1 I_58485 (I1085554,I2507,I996780,I996806,);
DFFARX1 I_58486 (I1085536,I2507,I996780,I996823,);
not I_58487 (I996831,I996823);
not I_58488 (I996848,I1085545);
nor I_58489 (I996865,I996848,I1085557);
not I_58490 (I996882,I1085539);
nor I_58491 (I996899,I996865,I1085548);
nor I_58492 (I996916,I996823,I996899);
DFFARX1 I_58493 (I996916,I2507,I996780,I996766,);
nor I_58494 (I996947,I1085548,I1085557);
nand I_58495 (I996964,I996947,I1085545);
DFFARX1 I_58496 (I996964,I2507,I996780,I996769,);
nor I_58497 (I996995,I996882,I1085548);
nand I_58498 (I997012,I996995,I1085560);
nor I_58499 (I997029,I996806,I997012);
DFFARX1 I_58500 (I997029,I2507,I996780,I996745,);
not I_58501 (I997060,I997012);
nand I_58502 (I996757,I996823,I997060);
DFFARX1 I_58503 (I997012,I2507,I996780,I997100,);
not I_58504 (I997108,I997100);
not I_58505 (I997125,I1085548);
not I_58506 (I997142,I1085536);
nor I_58507 (I997159,I997142,I1085539);
nor I_58508 (I996772,I997108,I997159);
nor I_58509 (I997190,I997142,I1085542);
and I_58510 (I997207,I997190,I1085551);
or I_58511 (I997224,I997207,I1085539);
DFFARX1 I_58512 (I997224,I2507,I996780,I997250,);
nor I_58513 (I996760,I997250,I996806);
not I_58514 (I997272,I997250);
and I_58515 (I997289,I997272,I996806);
nor I_58516 (I996754,I996831,I997289);
nand I_58517 (I997320,I997272,I996882);
nor I_58518 (I996748,I997142,I997320);
nand I_58519 (I996751,I997272,I997060);
nand I_58520 (I997365,I996882,I1085536);
nor I_58521 (I996763,I997125,I997365);
not I_58522 (I997426,I2514);
DFFARX1 I_58523 (I24294,I2507,I997426,I997452,);
DFFARX1 I_58524 (I24300,I2507,I997426,I997469,);
not I_58525 (I997477,I997469);
not I_58526 (I997494,I24294);
nor I_58527 (I997511,I997494,I24306);
not I_58528 (I997528,I24318);
nor I_58529 (I997545,I997511,I24312);
nor I_58530 (I997562,I997469,I997545);
DFFARX1 I_58531 (I997562,I2507,I997426,I997412,);
nor I_58532 (I997593,I24312,I24306);
nand I_58533 (I997610,I997593,I24294);
DFFARX1 I_58534 (I997610,I2507,I997426,I997415,);
nor I_58535 (I997641,I997528,I24312);
nand I_58536 (I997658,I997641,I24297);
nor I_58537 (I997675,I997452,I997658);
DFFARX1 I_58538 (I997675,I2507,I997426,I997391,);
not I_58539 (I997706,I997658);
nand I_58540 (I997403,I997469,I997706);
DFFARX1 I_58541 (I997658,I2507,I997426,I997746,);
not I_58542 (I997754,I997746);
not I_58543 (I997771,I24312);
not I_58544 (I997788,I24297);
nor I_58545 (I997805,I997788,I24318);
nor I_58546 (I997418,I997754,I997805);
nor I_58547 (I997836,I997788,I24315);
and I_58548 (I997853,I997836,I24309);
or I_58549 (I997870,I997853,I24303);
DFFARX1 I_58550 (I997870,I2507,I997426,I997896,);
nor I_58551 (I997406,I997896,I997452);
not I_58552 (I997918,I997896);
and I_58553 (I997935,I997918,I997452);
nor I_58554 (I997400,I997477,I997935);
nand I_58555 (I997966,I997918,I997528);
nor I_58556 (I997394,I997788,I997966);
nand I_58557 (I997397,I997918,I997706);
nand I_58558 (I998011,I997528,I24297);
nor I_58559 (I997409,I997771,I998011);
not I_58560 (I998072,I2514);
DFFARX1 I_58561 (I1393967,I2507,I998072,I998098,);
DFFARX1 I_58562 (I1393991,I2507,I998072,I998115,);
not I_58563 (I998123,I998115);
not I_58564 (I998140,I1393973);
nor I_58565 (I998157,I998140,I1393982);
not I_58566 (I998174,I1393967);
nor I_58567 (I998191,I998157,I1393988);
nor I_58568 (I998208,I998115,I998191);
DFFARX1 I_58569 (I998208,I2507,I998072,I998058,);
nor I_58570 (I998239,I1393988,I1393982);
nand I_58571 (I998256,I998239,I1393973);
DFFARX1 I_58572 (I998256,I2507,I998072,I998061,);
nor I_58573 (I998287,I998174,I1393988);
nand I_58574 (I998304,I998287,I1393985);
nor I_58575 (I998321,I998098,I998304);
DFFARX1 I_58576 (I998321,I2507,I998072,I998037,);
not I_58577 (I998352,I998304);
nand I_58578 (I998049,I998115,I998352);
DFFARX1 I_58579 (I998304,I2507,I998072,I998392,);
not I_58580 (I998400,I998392);
not I_58581 (I998417,I1393988);
not I_58582 (I998434,I1393979);
nor I_58583 (I998451,I998434,I1393967);
nor I_58584 (I998064,I998400,I998451);
nor I_58585 (I998482,I998434,I1393970);
and I_58586 (I998499,I998482,I1393994);
or I_58587 (I998516,I998499,I1393976);
DFFARX1 I_58588 (I998516,I2507,I998072,I998542,);
nor I_58589 (I998052,I998542,I998098);
not I_58590 (I998564,I998542);
and I_58591 (I998581,I998564,I998098);
nor I_58592 (I998046,I998123,I998581);
nand I_58593 (I998612,I998564,I998174);
nor I_58594 (I998040,I998434,I998612);
nand I_58595 (I998043,I998564,I998352);
nand I_58596 (I998657,I998174,I1393979);
nor I_58597 (I998055,I998417,I998657);
not I_58598 (I998718,I2514);
DFFARX1 I_58599 (I859170,I2507,I998718,I998744,);
DFFARX1 I_58600 (I859167,I2507,I998718,I998761,);
not I_58601 (I998769,I998761);
not I_58602 (I998786,I859167);
nor I_58603 (I998803,I998786,I859170);
not I_58604 (I998820,I859182);
nor I_58605 (I998837,I998803,I859176);
nor I_58606 (I998854,I998761,I998837);
DFFARX1 I_58607 (I998854,I2507,I998718,I998704,);
nor I_58608 (I998885,I859176,I859170);
nand I_58609 (I998902,I998885,I859167);
DFFARX1 I_58610 (I998902,I2507,I998718,I998707,);
nor I_58611 (I998933,I998820,I859176);
nand I_58612 (I998950,I998933,I859164);
nor I_58613 (I998967,I998744,I998950);
DFFARX1 I_58614 (I998967,I2507,I998718,I998683,);
not I_58615 (I998998,I998950);
nand I_58616 (I998695,I998761,I998998);
DFFARX1 I_58617 (I998950,I2507,I998718,I999038,);
not I_58618 (I999046,I999038);
not I_58619 (I999063,I859176);
not I_58620 (I999080,I859173);
nor I_58621 (I999097,I999080,I859182);
nor I_58622 (I998710,I999046,I999097);
nor I_58623 (I999128,I999080,I859179);
and I_58624 (I999145,I999128,I859185);
or I_58625 (I999162,I999145,I859164);
DFFARX1 I_58626 (I999162,I2507,I998718,I999188,);
nor I_58627 (I998698,I999188,I998744);
not I_58628 (I999210,I999188);
and I_58629 (I999227,I999210,I998744);
nor I_58630 (I998692,I998769,I999227);
nand I_58631 (I999258,I999210,I998820);
nor I_58632 (I998686,I999080,I999258);
nand I_58633 (I998689,I999210,I998998);
nand I_58634 (I999303,I998820,I859173);
nor I_58635 (I998701,I999063,I999303);
not I_58636 (I999364,I2514);
DFFARX1 I_58637 (I1175722,I2507,I999364,I999390,);
DFFARX1 I_58638 (I1175704,I2507,I999364,I999407,);
not I_58639 (I999415,I999407);
not I_58640 (I999432,I1175713);
nor I_58641 (I999449,I999432,I1175725);
not I_58642 (I999466,I1175707);
nor I_58643 (I999483,I999449,I1175716);
nor I_58644 (I999500,I999407,I999483);
DFFARX1 I_58645 (I999500,I2507,I999364,I999350,);
nor I_58646 (I999531,I1175716,I1175725);
nand I_58647 (I999548,I999531,I1175713);
DFFARX1 I_58648 (I999548,I2507,I999364,I999353,);
nor I_58649 (I999579,I999466,I1175716);
nand I_58650 (I999596,I999579,I1175728);
nor I_58651 (I999613,I999390,I999596);
DFFARX1 I_58652 (I999613,I2507,I999364,I999329,);
not I_58653 (I999644,I999596);
nand I_58654 (I999341,I999407,I999644);
DFFARX1 I_58655 (I999596,I2507,I999364,I999684,);
not I_58656 (I999692,I999684);
not I_58657 (I999709,I1175716);
not I_58658 (I999726,I1175704);
nor I_58659 (I999743,I999726,I1175707);
nor I_58660 (I999356,I999692,I999743);
nor I_58661 (I999774,I999726,I1175710);
and I_58662 (I999791,I999774,I1175719);
or I_58663 (I999808,I999791,I1175707);
DFFARX1 I_58664 (I999808,I2507,I999364,I999834,);
nor I_58665 (I999344,I999834,I999390);
not I_58666 (I999856,I999834);
and I_58667 (I999873,I999856,I999390);
nor I_58668 (I999338,I999415,I999873);
nand I_58669 (I999904,I999856,I999466);
nor I_58670 (I999332,I999726,I999904);
nand I_58671 (I999335,I999856,I999644);
nand I_58672 (I999949,I999466,I1175704);
nor I_58673 (I999347,I999709,I999949);
not I_58674 (I1000010,I2514);
DFFARX1 I_58675 (I645752,I2507,I1000010,I1000036,);
DFFARX1 I_58676 (I645746,I2507,I1000010,I1000053,);
not I_58677 (I1000061,I1000053);
not I_58678 (I1000078,I645761);
nor I_58679 (I1000095,I1000078,I645746);
not I_58680 (I1000112,I645755);
nor I_58681 (I1000129,I1000095,I645764);
nor I_58682 (I1000146,I1000053,I1000129);
DFFARX1 I_58683 (I1000146,I2507,I1000010,I999996,);
nor I_58684 (I1000177,I645764,I645746);
nand I_58685 (I1000194,I1000177,I645761);
DFFARX1 I_58686 (I1000194,I2507,I1000010,I999999,);
nor I_58687 (I1000225,I1000112,I645764);
nand I_58688 (I1000242,I1000225,I645749);
nor I_58689 (I1000259,I1000036,I1000242);
DFFARX1 I_58690 (I1000259,I2507,I1000010,I999975,);
not I_58691 (I1000290,I1000242);
nand I_58692 (I999987,I1000053,I1000290);
DFFARX1 I_58693 (I1000242,I2507,I1000010,I1000330,);
not I_58694 (I1000338,I1000330);
not I_58695 (I1000355,I645764);
not I_58696 (I1000372,I645758);
nor I_58697 (I1000389,I1000372,I645755);
nor I_58698 (I1000002,I1000338,I1000389);
nor I_58699 (I1000420,I1000372,I645767);
and I_58700 (I1000437,I1000420,I645770);
or I_58701 (I1000454,I1000437,I645749);
DFFARX1 I_58702 (I1000454,I2507,I1000010,I1000480,);
nor I_58703 (I999990,I1000480,I1000036);
not I_58704 (I1000502,I1000480);
and I_58705 (I1000519,I1000502,I1000036);
nor I_58706 (I999984,I1000061,I1000519);
nand I_58707 (I1000550,I1000502,I1000112);
nor I_58708 (I999978,I1000372,I1000550);
nand I_58709 (I999981,I1000502,I1000290);
nand I_58710 (I1000595,I1000112,I645758);
nor I_58711 (I999993,I1000355,I1000595);
not I_58712 (I1000656,I2514);
DFFARX1 I_58713 (I592573,I2507,I1000656,I1000682,);
DFFARX1 I_58714 (I592585,I2507,I1000656,I1000699,);
not I_58715 (I1000707,I1000699);
not I_58716 (I1000724,I592594);
nor I_58717 (I1000741,I1000724,I592570);
not I_58718 (I1000758,I592588);
nor I_58719 (I1000775,I1000741,I592582);
nor I_58720 (I1000792,I1000699,I1000775);
DFFARX1 I_58721 (I1000792,I2507,I1000656,I1000642,);
nor I_58722 (I1000823,I592582,I592570);
nand I_58723 (I1000840,I1000823,I592594);
DFFARX1 I_58724 (I1000840,I2507,I1000656,I1000645,);
nor I_58725 (I1000871,I1000758,I592582);
nand I_58726 (I1000888,I1000871,I592576);
nor I_58727 (I1000905,I1000682,I1000888);
DFFARX1 I_58728 (I1000905,I2507,I1000656,I1000621,);
not I_58729 (I1000936,I1000888);
nand I_58730 (I1000633,I1000699,I1000936);
DFFARX1 I_58731 (I1000888,I2507,I1000656,I1000976,);
not I_58732 (I1000984,I1000976);
not I_58733 (I1001001,I592582);
not I_58734 (I1001018,I592591);
nor I_58735 (I1001035,I1001018,I592588);
nor I_58736 (I1000648,I1000984,I1001035);
nor I_58737 (I1001066,I1001018,I592573);
and I_58738 (I1001083,I1001066,I592570);
or I_58739 (I1001100,I1001083,I592579);
DFFARX1 I_58740 (I1001100,I2507,I1000656,I1001126,);
nor I_58741 (I1000636,I1001126,I1000682);
not I_58742 (I1001148,I1001126);
and I_58743 (I1001165,I1001148,I1000682);
nor I_58744 (I1000630,I1000707,I1001165);
nand I_58745 (I1001196,I1001148,I1000758);
nor I_58746 (I1000624,I1001018,I1001196);
nand I_58747 (I1000627,I1001148,I1000936);
nand I_58748 (I1001241,I1000758,I592591);
nor I_58749 (I1000639,I1001001,I1001241);
not I_58750 (I1001302,I2514);
DFFARX1 I_58751 (I1199420,I2507,I1001302,I1001328,);
DFFARX1 I_58752 (I1199402,I2507,I1001302,I1001345,);
not I_58753 (I1001353,I1001345);
not I_58754 (I1001370,I1199411);
nor I_58755 (I1001387,I1001370,I1199423);
not I_58756 (I1001404,I1199405);
nor I_58757 (I1001421,I1001387,I1199414);
nor I_58758 (I1001438,I1001345,I1001421);
DFFARX1 I_58759 (I1001438,I2507,I1001302,I1001288,);
nor I_58760 (I1001469,I1199414,I1199423);
nand I_58761 (I1001486,I1001469,I1199411);
DFFARX1 I_58762 (I1001486,I2507,I1001302,I1001291,);
nor I_58763 (I1001517,I1001404,I1199414);
nand I_58764 (I1001534,I1001517,I1199426);
nor I_58765 (I1001551,I1001328,I1001534);
DFFARX1 I_58766 (I1001551,I2507,I1001302,I1001267,);
not I_58767 (I1001582,I1001534);
nand I_58768 (I1001279,I1001345,I1001582);
DFFARX1 I_58769 (I1001534,I2507,I1001302,I1001622,);
not I_58770 (I1001630,I1001622);
not I_58771 (I1001647,I1199414);
not I_58772 (I1001664,I1199402);
nor I_58773 (I1001681,I1001664,I1199405);
nor I_58774 (I1001294,I1001630,I1001681);
nor I_58775 (I1001712,I1001664,I1199408);
and I_58776 (I1001729,I1001712,I1199417);
or I_58777 (I1001746,I1001729,I1199405);
DFFARX1 I_58778 (I1001746,I2507,I1001302,I1001772,);
nor I_58779 (I1001282,I1001772,I1001328);
not I_58780 (I1001794,I1001772);
and I_58781 (I1001811,I1001794,I1001328);
nor I_58782 (I1001276,I1001353,I1001811);
nand I_58783 (I1001842,I1001794,I1001404);
nor I_58784 (I1001270,I1001664,I1001842);
nand I_58785 (I1001273,I1001794,I1001582);
nand I_58786 (I1001887,I1001404,I1199402);
nor I_58787 (I1001285,I1001647,I1001887);
not I_58788 (I1001948,I2514);
DFFARX1 I_58789 (I1381472,I2507,I1001948,I1001974,);
DFFARX1 I_58790 (I1381496,I2507,I1001948,I1001991,);
not I_58791 (I1001999,I1001991);
not I_58792 (I1002016,I1381478);
nor I_58793 (I1002033,I1002016,I1381487);
not I_58794 (I1002050,I1381472);
nor I_58795 (I1002067,I1002033,I1381493);
nor I_58796 (I1002084,I1001991,I1002067);
DFFARX1 I_58797 (I1002084,I2507,I1001948,I1001934,);
nor I_58798 (I1002115,I1381493,I1381487);
nand I_58799 (I1002132,I1002115,I1381478);
DFFARX1 I_58800 (I1002132,I2507,I1001948,I1001937,);
nor I_58801 (I1002163,I1002050,I1381493);
nand I_58802 (I1002180,I1002163,I1381490);
nor I_58803 (I1002197,I1001974,I1002180);
DFFARX1 I_58804 (I1002197,I2507,I1001948,I1001913,);
not I_58805 (I1002228,I1002180);
nand I_58806 (I1001925,I1001991,I1002228);
DFFARX1 I_58807 (I1002180,I2507,I1001948,I1002268,);
not I_58808 (I1002276,I1002268);
not I_58809 (I1002293,I1381493);
not I_58810 (I1002310,I1381484);
nor I_58811 (I1002327,I1002310,I1381472);
nor I_58812 (I1001940,I1002276,I1002327);
nor I_58813 (I1002358,I1002310,I1381475);
and I_58814 (I1002375,I1002358,I1381499);
or I_58815 (I1002392,I1002375,I1381481);
DFFARX1 I_58816 (I1002392,I2507,I1001948,I1002418,);
nor I_58817 (I1001928,I1002418,I1001974);
not I_58818 (I1002440,I1002418);
and I_58819 (I1002457,I1002440,I1001974);
nor I_58820 (I1001922,I1001999,I1002457);
nand I_58821 (I1002488,I1002440,I1002050);
nor I_58822 (I1001916,I1002310,I1002488);
nand I_58823 (I1001919,I1002440,I1002228);
nand I_58824 (I1002533,I1002050,I1381484);
nor I_58825 (I1001931,I1002293,I1002533);
not I_58826 (I1002594,I2514);
DFFARX1 I_58827 (I1083820,I2507,I1002594,I1002620,);
DFFARX1 I_58828 (I1083802,I2507,I1002594,I1002637,);
not I_58829 (I1002645,I1002637);
not I_58830 (I1002662,I1083811);
nor I_58831 (I1002679,I1002662,I1083823);
not I_58832 (I1002696,I1083805);
nor I_58833 (I1002713,I1002679,I1083814);
nor I_58834 (I1002730,I1002637,I1002713);
DFFARX1 I_58835 (I1002730,I2507,I1002594,I1002580,);
nor I_58836 (I1002761,I1083814,I1083823);
nand I_58837 (I1002778,I1002761,I1083811);
DFFARX1 I_58838 (I1002778,I2507,I1002594,I1002583,);
nor I_58839 (I1002809,I1002696,I1083814);
nand I_58840 (I1002826,I1002809,I1083826);
nor I_58841 (I1002843,I1002620,I1002826);
DFFARX1 I_58842 (I1002843,I2507,I1002594,I1002559,);
not I_58843 (I1002874,I1002826);
nand I_58844 (I1002571,I1002637,I1002874);
DFFARX1 I_58845 (I1002826,I2507,I1002594,I1002914,);
not I_58846 (I1002922,I1002914);
not I_58847 (I1002939,I1083814);
not I_58848 (I1002956,I1083802);
nor I_58849 (I1002973,I1002956,I1083805);
nor I_58850 (I1002586,I1002922,I1002973);
nor I_58851 (I1003004,I1002956,I1083808);
and I_58852 (I1003021,I1003004,I1083817);
or I_58853 (I1003038,I1003021,I1083805);
DFFARX1 I_58854 (I1003038,I2507,I1002594,I1003064,);
nor I_58855 (I1002574,I1003064,I1002620);
not I_58856 (I1003086,I1003064);
and I_58857 (I1003103,I1003086,I1002620);
nor I_58858 (I1002568,I1002645,I1003103);
nand I_58859 (I1003134,I1003086,I1002696);
nor I_58860 (I1002562,I1002956,I1003134);
nand I_58861 (I1002565,I1003086,I1002874);
nand I_58862 (I1003179,I1002696,I1083802);
nor I_58863 (I1002577,I1002939,I1003179);
not I_58864 (I1003240,I2514);
DFFARX1 I_58865 (I1366597,I2507,I1003240,I1003266,);
DFFARX1 I_58866 (I1366621,I2507,I1003240,I1003283,);
not I_58867 (I1003291,I1003283);
not I_58868 (I1003308,I1366603);
nor I_58869 (I1003325,I1003308,I1366612);
not I_58870 (I1003342,I1366597);
nor I_58871 (I1003359,I1003325,I1366618);
nor I_58872 (I1003376,I1003283,I1003359);
DFFARX1 I_58873 (I1003376,I2507,I1003240,I1003226,);
nor I_58874 (I1003407,I1366618,I1366612);
nand I_58875 (I1003424,I1003407,I1366603);
DFFARX1 I_58876 (I1003424,I2507,I1003240,I1003229,);
nor I_58877 (I1003455,I1003342,I1366618);
nand I_58878 (I1003472,I1003455,I1366615);
nor I_58879 (I1003489,I1003266,I1003472);
DFFARX1 I_58880 (I1003489,I2507,I1003240,I1003205,);
not I_58881 (I1003520,I1003472);
nand I_58882 (I1003217,I1003283,I1003520);
DFFARX1 I_58883 (I1003472,I2507,I1003240,I1003560,);
not I_58884 (I1003568,I1003560);
not I_58885 (I1003585,I1366618);
not I_58886 (I1003602,I1366609);
nor I_58887 (I1003619,I1003602,I1366597);
nor I_58888 (I1003232,I1003568,I1003619);
nor I_58889 (I1003650,I1003602,I1366600);
and I_58890 (I1003667,I1003650,I1366624);
or I_58891 (I1003684,I1003667,I1366606);
DFFARX1 I_58892 (I1003684,I2507,I1003240,I1003710,);
nor I_58893 (I1003220,I1003710,I1003266);
not I_58894 (I1003732,I1003710);
and I_58895 (I1003749,I1003732,I1003266);
nor I_58896 (I1003214,I1003291,I1003749);
nand I_58897 (I1003780,I1003732,I1003342);
nor I_58898 (I1003208,I1003602,I1003780);
nand I_58899 (I1003211,I1003732,I1003520);
nand I_58900 (I1003825,I1003342,I1366609);
nor I_58901 (I1003223,I1003585,I1003825);
not I_58902 (I1003886,I2514);
DFFARX1 I_58903 (I400085,I2507,I1003886,I1003912,);
DFFARX1 I_58904 (I400082,I2507,I1003886,I1003929,);
not I_58905 (I1003937,I1003929);
not I_58906 (I1003954,I400097);
nor I_58907 (I1003971,I1003954,I400100);
not I_58908 (I1003988,I400088);
nor I_58909 (I1004005,I1003971,I400094);
nor I_58910 (I1004022,I1003929,I1004005);
DFFARX1 I_58911 (I1004022,I2507,I1003886,I1003872,);
nor I_58912 (I1004053,I400094,I400100);
nand I_58913 (I1004070,I1004053,I400097);
DFFARX1 I_58914 (I1004070,I2507,I1003886,I1003875,);
nor I_58915 (I1004101,I1003988,I400094);
nand I_58916 (I1004118,I1004101,I400106);
nor I_58917 (I1004135,I1003912,I1004118);
DFFARX1 I_58918 (I1004135,I2507,I1003886,I1003851,);
not I_58919 (I1004166,I1004118);
nand I_58920 (I1003863,I1003929,I1004166);
DFFARX1 I_58921 (I1004118,I2507,I1003886,I1004206,);
not I_58922 (I1004214,I1004206);
not I_58923 (I1004231,I400094);
not I_58924 (I1004248,I400079);
nor I_58925 (I1004265,I1004248,I400088);
nor I_58926 (I1003878,I1004214,I1004265);
nor I_58927 (I1004296,I1004248,I400091);
and I_58928 (I1004313,I1004296,I400079);
or I_58929 (I1004330,I1004313,I400103);
DFFARX1 I_58930 (I1004330,I2507,I1003886,I1004356,);
nor I_58931 (I1003866,I1004356,I1003912);
not I_58932 (I1004378,I1004356);
and I_58933 (I1004395,I1004378,I1003912);
nor I_58934 (I1003860,I1003937,I1004395);
nand I_58935 (I1004426,I1004378,I1003988);
nor I_58936 (I1003854,I1004248,I1004426);
nand I_58937 (I1003857,I1004378,I1004166);
nand I_58938 (I1004471,I1003988,I400079);
nor I_58939 (I1003869,I1004231,I1004471);
not I_58940 (I1004532,I2514);
DFFARX1 I_58941 (I1243348,I2507,I1004532,I1004558,);
DFFARX1 I_58942 (I1243354,I2507,I1004532,I1004575,);
not I_58943 (I1004583,I1004575);
not I_58944 (I1004600,I1243351);
nor I_58945 (I1004617,I1004600,I1243330);
not I_58946 (I1004634,I1243333);
nor I_58947 (I1004651,I1004617,I1243339);
nor I_58948 (I1004668,I1004575,I1004651);
DFFARX1 I_58949 (I1004668,I2507,I1004532,I1004518,);
nor I_58950 (I1004699,I1243339,I1243330);
nand I_58951 (I1004716,I1004699,I1243351);
DFFARX1 I_58952 (I1004716,I2507,I1004532,I1004521,);
nor I_58953 (I1004747,I1004634,I1243339);
nand I_58954 (I1004764,I1004747,I1243333);
nor I_58955 (I1004781,I1004558,I1004764);
DFFARX1 I_58956 (I1004781,I2507,I1004532,I1004497,);
not I_58957 (I1004812,I1004764);
nand I_58958 (I1004509,I1004575,I1004812);
DFFARX1 I_58959 (I1004764,I2507,I1004532,I1004852,);
not I_58960 (I1004860,I1004852);
not I_58961 (I1004877,I1243339);
not I_58962 (I1004894,I1243342);
nor I_58963 (I1004911,I1004894,I1243333);
nor I_58964 (I1004524,I1004860,I1004911);
nor I_58965 (I1004942,I1004894,I1243330);
and I_58966 (I1004959,I1004942,I1243336);
or I_58967 (I1004976,I1004959,I1243345);
DFFARX1 I_58968 (I1004976,I2507,I1004532,I1005002,);
nor I_58969 (I1004512,I1005002,I1004558);
not I_58970 (I1005024,I1005002);
and I_58971 (I1005041,I1005024,I1004558);
nor I_58972 (I1004506,I1004583,I1005041);
nand I_58973 (I1005072,I1005024,I1004634);
nor I_58974 (I1004500,I1004894,I1005072);
nand I_58975 (I1004503,I1005024,I1004812);
nand I_58976 (I1005117,I1004634,I1243342);
nor I_58977 (I1004515,I1004877,I1005117);
not I_58978 (I1005178,I2514);
DFFARX1 I_58979 (I290769,I2507,I1005178,I1005204,);
DFFARX1 I_58980 (I290775,I2507,I1005178,I1005221,);
not I_58981 (I1005229,I1005221);
not I_58982 (I1005246,I290796);
nor I_58983 (I1005263,I1005246,I290784);
not I_58984 (I1005280,I290793);
nor I_58985 (I1005297,I1005263,I290778);
nor I_58986 (I1005314,I1005221,I1005297);
DFFARX1 I_58987 (I1005314,I2507,I1005178,I1005164,);
nor I_58988 (I1005345,I290778,I290784);
nand I_58989 (I1005362,I1005345,I290796);
DFFARX1 I_58990 (I1005362,I2507,I1005178,I1005167,);
nor I_58991 (I1005393,I1005280,I290778);
nand I_58992 (I1005410,I1005393,I290769);
nor I_58993 (I1005427,I1005204,I1005410);
DFFARX1 I_58994 (I1005427,I2507,I1005178,I1005143,);
not I_58995 (I1005458,I1005410);
nand I_58996 (I1005155,I1005221,I1005458);
DFFARX1 I_58997 (I1005410,I2507,I1005178,I1005498,);
not I_58998 (I1005506,I1005498);
not I_58999 (I1005523,I290778);
not I_59000 (I1005540,I290781);
nor I_59001 (I1005557,I1005540,I290793);
nor I_59002 (I1005170,I1005506,I1005557);
nor I_59003 (I1005588,I1005540,I290790);
and I_59004 (I1005605,I1005588,I290772);
or I_59005 (I1005622,I1005605,I290787);
DFFARX1 I_59006 (I1005622,I2507,I1005178,I1005648,);
nor I_59007 (I1005158,I1005648,I1005204);
not I_59008 (I1005670,I1005648);
and I_59009 (I1005687,I1005670,I1005204);
nor I_59010 (I1005152,I1005229,I1005687);
nand I_59011 (I1005718,I1005670,I1005280);
nor I_59012 (I1005146,I1005540,I1005718);
nand I_59013 (I1005149,I1005670,I1005458);
nand I_59014 (I1005763,I1005280,I290781);
nor I_59015 (I1005161,I1005523,I1005763);
not I_59016 (I1005824,I2514);
DFFARX1 I_59017 (I695460,I2507,I1005824,I1005850,);
DFFARX1 I_59018 (I695454,I2507,I1005824,I1005867,);
not I_59019 (I1005875,I1005867);
not I_59020 (I1005892,I695469);
nor I_59021 (I1005909,I1005892,I695454);
not I_59022 (I1005926,I695463);
nor I_59023 (I1005943,I1005909,I695472);
nor I_59024 (I1005960,I1005867,I1005943);
DFFARX1 I_59025 (I1005960,I2507,I1005824,I1005810,);
nor I_59026 (I1005991,I695472,I695454);
nand I_59027 (I1006008,I1005991,I695469);
DFFARX1 I_59028 (I1006008,I2507,I1005824,I1005813,);
nor I_59029 (I1006039,I1005926,I695472);
nand I_59030 (I1006056,I1006039,I695457);
nor I_59031 (I1006073,I1005850,I1006056);
DFFARX1 I_59032 (I1006073,I2507,I1005824,I1005789,);
not I_59033 (I1006104,I1006056);
nand I_59034 (I1005801,I1005867,I1006104);
DFFARX1 I_59035 (I1006056,I2507,I1005824,I1006144,);
not I_59036 (I1006152,I1006144);
not I_59037 (I1006169,I695472);
not I_59038 (I1006186,I695466);
nor I_59039 (I1006203,I1006186,I695463);
nor I_59040 (I1005816,I1006152,I1006203);
nor I_59041 (I1006234,I1006186,I695475);
and I_59042 (I1006251,I1006234,I695478);
or I_59043 (I1006268,I1006251,I695457);
DFFARX1 I_59044 (I1006268,I2507,I1005824,I1006294,);
nor I_59045 (I1005804,I1006294,I1005850);
not I_59046 (I1006316,I1006294);
and I_59047 (I1006333,I1006316,I1005850);
nor I_59048 (I1005798,I1005875,I1006333);
nand I_59049 (I1006364,I1006316,I1005926);
nor I_59050 (I1005792,I1006186,I1006364);
nand I_59051 (I1005795,I1006316,I1006104);
nand I_59052 (I1006409,I1005926,I695466);
nor I_59053 (I1005807,I1006169,I1006409);
not I_59054 (I1006470,I2514);
DFFARX1 I_59055 (I768288,I2507,I1006470,I1006496,);
DFFARX1 I_59056 (I768282,I2507,I1006470,I1006513,);
not I_59057 (I1006521,I1006513);
not I_59058 (I1006538,I768297);
nor I_59059 (I1006555,I1006538,I768282);
not I_59060 (I1006572,I768291);
nor I_59061 (I1006589,I1006555,I768300);
nor I_59062 (I1006606,I1006513,I1006589);
DFFARX1 I_59063 (I1006606,I2507,I1006470,I1006456,);
nor I_59064 (I1006637,I768300,I768282);
nand I_59065 (I1006654,I1006637,I768297);
DFFARX1 I_59066 (I1006654,I2507,I1006470,I1006459,);
nor I_59067 (I1006685,I1006572,I768300);
nand I_59068 (I1006702,I1006685,I768285);
nor I_59069 (I1006719,I1006496,I1006702);
DFFARX1 I_59070 (I1006719,I2507,I1006470,I1006435,);
not I_59071 (I1006750,I1006702);
nand I_59072 (I1006447,I1006513,I1006750);
DFFARX1 I_59073 (I1006702,I2507,I1006470,I1006790,);
not I_59074 (I1006798,I1006790);
not I_59075 (I1006815,I768300);
not I_59076 (I1006832,I768294);
nor I_59077 (I1006849,I1006832,I768291);
nor I_59078 (I1006462,I1006798,I1006849);
nor I_59079 (I1006880,I1006832,I768303);
and I_59080 (I1006897,I1006880,I768306);
or I_59081 (I1006914,I1006897,I768285);
DFFARX1 I_59082 (I1006914,I2507,I1006470,I1006940,);
nor I_59083 (I1006450,I1006940,I1006496);
not I_59084 (I1006962,I1006940);
and I_59085 (I1006979,I1006962,I1006496);
nor I_59086 (I1006444,I1006521,I1006979);
nand I_59087 (I1007010,I1006962,I1006572);
nor I_59088 (I1006438,I1006832,I1007010);
nand I_59089 (I1006441,I1006962,I1006750);
nand I_59090 (I1007055,I1006572,I768294);
nor I_59091 (I1006453,I1006815,I1007055);
not I_59092 (I1007116,I2514);
DFFARX1 I_59093 (I63292,I2507,I1007116,I1007142,);
DFFARX1 I_59094 (I63298,I2507,I1007116,I1007159,);
not I_59095 (I1007167,I1007159);
not I_59096 (I1007184,I63316);
nor I_59097 (I1007201,I1007184,I63295);
not I_59098 (I1007218,I63301);
nor I_59099 (I1007235,I1007201,I63307);
nor I_59100 (I1007252,I1007159,I1007235);
DFFARX1 I_59101 (I1007252,I2507,I1007116,I1007102,);
nor I_59102 (I1007283,I63307,I63295);
nand I_59103 (I1007300,I1007283,I63316);
DFFARX1 I_59104 (I1007300,I2507,I1007116,I1007105,);
nor I_59105 (I1007331,I1007218,I63307);
nand I_59106 (I1007348,I1007331,I63313);
nor I_59107 (I1007365,I1007142,I1007348);
DFFARX1 I_59108 (I1007365,I2507,I1007116,I1007081,);
not I_59109 (I1007396,I1007348);
nand I_59110 (I1007093,I1007159,I1007396);
DFFARX1 I_59111 (I1007348,I2507,I1007116,I1007436,);
not I_59112 (I1007444,I1007436);
not I_59113 (I1007461,I63307);
not I_59114 (I1007478,I63295);
nor I_59115 (I1007495,I1007478,I63301);
nor I_59116 (I1007108,I1007444,I1007495);
nor I_59117 (I1007526,I1007478,I63304);
and I_59118 (I1007543,I1007526,I63292);
or I_59119 (I1007560,I1007543,I63310);
DFFARX1 I_59120 (I1007560,I2507,I1007116,I1007586,);
nor I_59121 (I1007096,I1007586,I1007142);
not I_59122 (I1007608,I1007586);
and I_59123 (I1007625,I1007608,I1007142);
nor I_59124 (I1007090,I1007167,I1007625);
nand I_59125 (I1007656,I1007608,I1007218);
nor I_59126 (I1007084,I1007478,I1007656);
nand I_59127 (I1007087,I1007608,I1007396);
nand I_59128 (I1007701,I1007218,I63295);
nor I_59129 (I1007099,I1007461,I1007701);
not I_59130 (I1007762,I2514);
DFFARX1 I_59131 (I779066,I2507,I1007762,I1007788,);
DFFARX1 I_59132 (I779063,I2507,I1007762,I1007805,);
not I_59133 (I1007813,I1007805);
not I_59134 (I1007830,I779063);
nor I_59135 (I1007847,I1007830,I779066);
not I_59136 (I1007864,I779078);
nor I_59137 (I1007881,I1007847,I779072);
nor I_59138 (I1007898,I1007805,I1007881);
DFFARX1 I_59139 (I1007898,I2507,I1007762,I1007748,);
nor I_59140 (I1007929,I779072,I779066);
nand I_59141 (I1007946,I1007929,I779063);
DFFARX1 I_59142 (I1007946,I2507,I1007762,I1007751,);
nor I_59143 (I1007977,I1007864,I779072);
nand I_59144 (I1007994,I1007977,I779060);
nor I_59145 (I1008011,I1007788,I1007994);
DFFARX1 I_59146 (I1008011,I2507,I1007762,I1007727,);
not I_59147 (I1008042,I1007994);
nand I_59148 (I1007739,I1007805,I1008042);
DFFARX1 I_59149 (I1007994,I2507,I1007762,I1008082,);
not I_59150 (I1008090,I1008082);
not I_59151 (I1008107,I779072);
not I_59152 (I1008124,I779069);
nor I_59153 (I1008141,I1008124,I779078);
nor I_59154 (I1007754,I1008090,I1008141);
nor I_59155 (I1008172,I1008124,I779075);
and I_59156 (I1008189,I1008172,I779081);
or I_59157 (I1008206,I1008189,I779060);
DFFARX1 I_59158 (I1008206,I2507,I1007762,I1008232,);
nor I_59159 (I1007742,I1008232,I1007788);
not I_59160 (I1008254,I1008232);
and I_59161 (I1008271,I1008254,I1007788);
nor I_59162 (I1007736,I1007813,I1008271);
nand I_59163 (I1008302,I1008254,I1007864);
nor I_59164 (I1007730,I1008124,I1008302);
nand I_59165 (I1007733,I1008254,I1008042);
nand I_59166 (I1008347,I1007864,I779069);
nor I_59167 (I1007745,I1008107,I1008347);
not I_59168 (I1008408,I2514);
DFFARX1 I_59169 (I631880,I2507,I1008408,I1008434,);
DFFARX1 I_59170 (I631874,I2507,I1008408,I1008451,);
not I_59171 (I1008459,I1008451);
not I_59172 (I1008476,I631889);
nor I_59173 (I1008493,I1008476,I631874);
not I_59174 (I1008510,I631883);
nor I_59175 (I1008527,I1008493,I631892);
nor I_59176 (I1008544,I1008451,I1008527);
DFFARX1 I_59177 (I1008544,I2507,I1008408,I1008394,);
nor I_59178 (I1008575,I631892,I631874);
nand I_59179 (I1008592,I1008575,I631889);
DFFARX1 I_59180 (I1008592,I2507,I1008408,I1008397,);
nor I_59181 (I1008623,I1008510,I631892);
nand I_59182 (I1008640,I1008623,I631877);
nor I_59183 (I1008657,I1008434,I1008640);
DFFARX1 I_59184 (I1008657,I2507,I1008408,I1008373,);
not I_59185 (I1008688,I1008640);
nand I_59186 (I1008385,I1008451,I1008688);
DFFARX1 I_59187 (I1008640,I2507,I1008408,I1008728,);
not I_59188 (I1008736,I1008728);
not I_59189 (I1008753,I631892);
not I_59190 (I1008770,I631886);
nor I_59191 (I1008787,I1008770,I631883);
nor I_59192 (I1008400,I1008736,I1008787);
nor I_59193 (I1008818,I1008770,I631895);
and I_59194 (I1008835,I1008818,I631898);
or I_59195 (I1008852,I1008835,I631877);
DFFARX1 I_59196 (I1008852,I2507,I1008408,I1008878,);
nor I_59197 (I1008388,I1008878,I1008434);
not I_59198 (I1008900,I1008878);
and I_59199 (I1008917,I1008900,I1008434);
nor I_59200 (I1008382,I1008459,I1008917);
nand I_59201 (I1008948,I1008900,I1008510);
nor I_59202 (I1008376,I1008770,I1008948);
nand I_59203 (I1008379,I1008900,I1008688);
nand I_59204 (I1008993,I1008510,I631886);
nor I_59205 (I1008391,I1008753,I1008993);
not I_59206 (I1009048,I2514);
DFFARX1 I_59207 (I250211,I2507,I1009048,I1009074,);
DFFARX1 I_59208 (I1009074,I2507,I1009048,I1009091,);
not I_59209 (I1009040,I1009091);
not I_59210 (I1009113,I1009074);
DFFARX1 I_59211 (I250208,I2507,I1009048,I1009139,);
nand I_59212 (I1009147,I1009139,I250202);
not I_59213 (I1009164,I250202);
not I_59214 (I1009181,I250199);
nand I_59215 (I1009198,I250193,I250190);
and I_59216 (I1009215,I250193,I250190);
not I_59217 (I1009232,I250205);
nand I_59218 (I1009249,I1009232,I1009181);
nor I_59219 (I1009022,I1009249,I1009147);
nor I_59220 (I1009280,I1009164,I1009249);
nand I_59221 (I1009025,I1009215,I1009280);
not I_59222 (I1009311,I250217);
nor I_59223 (I1009328,I1009311,I250193);
nor I_59224 (I1009345,I1009328,I250205);
nor I_59225 (I1009362,I1009113,I1009345);
DFFARX1 I_59226 (I1009362,I2507,I1009048,I1009034,);
not I_59227 (I1009393,I1009328);
DFFARX1 I_59228 (I1009393,I2507,I1009048,I1009037,);
and I_59229 (I1009031,I1009139,I1009328);
nor I_59230 (I1009438,I1009311,I250214);
and I_59231 (I1009455,I1009438,I250190);
or I_59232 (I1009472,I1009455,I250196);
DFFARX1 I_59233 (I1009472,I2507,I1009048,I1009498,);
nor I_59234 (I1009506,I1009498,I1009232);
DFFARX1 I_59235 (I1009506,I2507,I1009048,I1009019,);
nand I_59236 (I1009537,I1009498,I1009139);
nand I_59237 (I1009554,I1009232,I1009537);
nor I_59238 (I1009028,I1009554,I1009198);
not I_59239 (I1009609,I2514);
DFFARX1 I_59240 (I317667,I2507,I1009609,I1009635,);
DFFARX1 I_59241 (I1009635,I2507,I1009609,I1009652,);
not I_59242 (I1009601,I1009652);
not I_59243 (I1009674,I1009635);
DFFARX1 I_59244 (I317664,I2507,I1009609,I1009700,);
nand I_59245 (I1009708,I1009700,I317658);
not I_59246 (I1009725,I317658);
not I_59247 (I1009742,I317655);
nand I_59248 (I1009759,I317649,I317646);
and I_59249 (I1009776,I317649,I317646);
not I_59250 (I1009793,I317661);
nand I_59251 (I1009810,I1009793,I1009742);
nor I_59252 (I1009583,I1009810,I1009708);
nor I_59253 (I1009841,I1009725,I1009810);
nand I_59254 (I1009586,I1009776,I1009841);
not I_59255 (I1009872,I317673);
nor I_59256 (I1009889,I1009872,I317649);
nor I_59257 (I1009906,I1009889,I317661);
nor I_59258 (I1009923,I1009674,I1009906);
DFFARX1 I_59259 (I1009923,I2507,I1009609,I1009595,);
not I_59260 (I1009954,I1009889);
DFFARX1 I_59261 (I1009954,I2507,I1009609,I1009598,);
and I_59262 (I1009592,I1009700,I1009889);
nor I_59263 (I1009999,I1009872,I317670);
and I_59264 (I1010016,I1009999,I317646);
or I_59265 (I1010033,I1010016,I317652);
DFFARX1 I_59266 (I1010033,I2507,I1009609,I1010059,);
nor I_59267 (I1010067,I1010059,I1009793);
DFFARX1 I_59268 (I1010067,I2507,I1009609,I1009580,);
nand I_59269 (I1010098,I1010059,I1009700);
nand I_59270 (I1010115,I1009793,I1010098);
nor I_59271 (I1009589,I1010115,I1009759);
not I_59272 (I1010170,I2514);
DFFARX1 I_59273 (I299222,I2507,I1010170,I1010196,);
DFFARX1 I_59274 (I1010196,I2507,I1010170,I1010213,);
not I_59275 (I1010162,I1010213);
not I_59276 (I1010235,I1010196);
DFFARX1 I_59277 (I299219,I2507,I1010170,I1010261,);
nand I_59278 (I1010269,I1010261,I299213);
not I_59279 (I1010286,I299213);
not I_59280 (I1010303,I299210);
nand I_59281 (I1010320,I299204,I299201);
and I_59282 (I1010337,I299204,I299201);
not I_59283 (I1010354,I299216);
nand I_59284 (I1010371,I1010354,I1010303);
nor I_59285 (I1010144,I1010371,I1010269);
nor I_59286 (I1010402,I1010286,I1010371);
nand I_59287 (I1010147,I1010337,I1010402);
not I_59288 (I1010433,I299228);
nor I_59289 (I1010450,I1010433,I299204);
nor I_59290 (I1010467,I1010450,I299216);
nor I_59291 (I1010484,I1010235,I1010467);
DFFARX1 I_59292 (I1010484,I2507,I1010170,I1010156,);
not I_59293 (I1010515,I1010450);
DFFARX1 I_59294 (I1010515,I2507,I1010170,I1010159,);
and I_59295 (I1010153,I1010261,I1010450);
nor I_59296 (I1010560,I1010433,I299225);
and I_59297 (I1010577,I1010560,I299201);
or I_59298 (I1010594,I1010577,I299207);
DFFARX1 I_59299 (I1010594,I2507,I1010170,I1010620,);
nor I_59300 (I1010628,I1010620,I1010354);
DFFARX1 I_59301 (I1010628,I2507,I1010170,I1010141,);
nand I_59302 (I1010659,I1010620,I1010261);
nand I_59303 (I1010676,I1010354,I1010659);
nor I_59304 (I1010150,I1010676,I1010320);
not I_59305 (I1010731,I2514);
DFFARX1 I_59306 (I1182655,I2507,I1010731,I1010757,);
DFFARX1 I_59307 (I1010757,I2507,I1010731,I1010774,);
not I_59308 (I1010723,I1010774);
not I_59309 (I1010796,I1010757);
DFFARX1 I_59310 (I1182646,I2507,I1010731,I1010822,);
nand I_59311 (I1010830,I1010822,I1182643);
not I_59312 (I1010847,I1182643);
not I_59313 (I1010864,I1182652);
nand I_59314 (I1010881,I1182661,I1182643);
and I_59315 (I1010898,I1182661,I1182643);
not I_59316 (I1010915,I1182640);
nand I_59317 (I1010932,I1010915,I1010864);
nor I_59318 (I1010705,I1010932,I1010830);
nor I_59319 (I1010963,I1010847,I1010932);
nand I_59320 (I1010708,I1010898,I1010963);
not I_59321 (I1010994,I1182649);
nor I_59322 (I1011011,I1010994,I1182661);
nor I_59323 (I1011028,I1011011,I1182640);
nor I_59324 (I1011045,I1010796,I1011028);
DFFARX1 I_59325 (I1011045,I2507,I1010731,I1010717,);
not I_59326 (I1011076,I1011011);
DFFARX1 I_59327 (I1011076,I2507,I1010731,I1010720,);
and I_59328 (I1010714,I1010822,I1011011);
nor I_59329 (I1011121,I1010994,I1182664);
and I_59330 (I1011138,I1011121,I1182640);
or I_59331 (I1011155,I1011138,I1182658);
DFFARX1 I_59332 (I1011155,I2507,I1010731,I1011181,);
nor I_59333 (I1011189,I1011181,I1010915);
DFFARX1 I_59334 (I1011189,I2507,I1010731,I1010702,);
nand I_59335 (I1011220,I1011181,I1010822);
nand I_59336 (I1011237,I1010915,I1011220);
nor I_59337 (I1010711,I1011237,I1010881);
not I_59338 (I1011292,I2514);
DFFARX1 I_59339 (I244243,I2507,I1011292,I1011318,);
DFFARX1 I_59340 (I1011318,I2507,I1011292,I1011335,);
not I_59341 (I1011284,I1011335);
not I_59342 (I1011357,I1011318);
DFFARX1 I_59343 (I244258,I2507,I1011292,I1011383,);
nand I_59344 (I1011391,I1011383,I244240);
not I_59345 (I1011408,I244240);
not I_59346 (I1011425,I244249);
nand I_59347 (I1011442,I244255,I244246);
and I_59348 (I1011459,I244255,I244246);
not I_59349 (I1011476,I244243);
nand I_59350 (I1011493,I1011476,I1011425);
nor I_59351 (I1011266,I1011493,I1011391);
nor I_59352 (I1011524,I1011408,I1011493);
nand I_59353 (I1011269,I1011459,I1011524);
not I_59354 (I1011555,I244240);
nor I_59355 (I1011572,I1011555,I244255);
nor I_59356 (I1011589,I1011572,I244243);
nor I_59357 (I1011606,I1011357,I1011589);
DFFARX1 I_59358 (I1011606,I2507,I1011292,I1011278,);
not I_59359 (I1011637,I1011572);
DFFARX1 I_59360 (I1011637,I2507,I1011292,I1011281,);
and I_59361 (I1011275,I1011383,I1011572);
nor I_59362 (I1011682,I1011555,I244264);
and I_59363 (I1011699,I1011682,I244261);
or I_59364 (I1011716,I1011699,I244252);
DFFARX1 I_59365 (I1011716,I2507,I1011292,I1011742,);
nor I_59366 (I1011750,I1011742,I1011476);
DFFARX1 I_59367 (I1011750,I2507,I1011292,I1011263,);
nand I_59368 (I1011781,I1011742,I1011383);
nand I_59369 (I1011798,I1011476,I1011781);
nor I_59370 (I1011272,I1011798,I1011442);
not I_59371 (I1011853,I2514);
DFFARX1 I_59372 (I840728,I2507,I1011853,I1011879,);
DFFARX1 I_59373 (I1011879,I2507,I1011853,I1011896,);
not I_59374 (I1011845,I1011896);
not I_59375 (I1011918,I1011879);
DFFARX1 I_59376 (I840725,I2507,I1011853,I1011944,);
nand I_59377 (I1011952,I1011944,I840740);
not I_59378 (I1011969,I840740);
not I_59379 (I1011986,I840737);
nand I_59380 (I1012003,I840734,I840722);
and I_59381 (I1012020,I840734,I840722);
not I_59382 (I1012037,I840719);
nand I_59383 (I1012054,I1012037,I1011986);
nor I_59384 (I1011827,I1012054,I1011952);
nor I_59385 (I1012085,I1011969,I1012054);
nand I_59386 (I1011830,I1012020,I1012085);
not I_59387 (I1012116,I840725);
nor I_59388 (I1012133,I1012116,I840734);
nor I_59389 (I1012150,I1012133,I840719);
nor I_59390 (I1012167,I1011918,I1012150);
DFFARX1 I_59391 (I1012167,I2507,I1011853,I1011839,);
not I_59392 (I1012198,I1012133);
DFFARX1 I_59393 (I1012198,I2507,I1011853,I1011842,);
and I_59394 (I1011836,I1011944,I1012133);
nor I_59395 (I1012243,I1012116,I840731);
and I_59396 (I1012260,I1012243,I840719);
or I_59397 (I1012277,I1012260,I840722);
DFFARX1 I_59398 (I1012277,I2507,I1011853,I1012303,);
nor I_59399 (I1012311,I1012303,I1012037);
DFFARX1 I_59400 (I1012311,I2507,I1011853,I1011824,);
nand I_59401 (I1012342,I1012303,I1011944);
nand I_59402 (I1012359,I1012037,I1012342);
nor I_59403 (I1011833,I1012359,I1012003);
not I_59404 (I1012414,I2514);
DFFARX1 I_59405 (I1292905,I2507,I1012414,I1012440,);
DFFARX1 I_59406 (I1012440,I2507,I1012414,I1012457,);
not I_59407 (I1012406,I1012457);
not I_59408 (I1012479,I1012440);
DFFARX1 I_59409 (I1292902,I2507,I1012414,I1012505,);
nand I_59410 (I1012513,I1012505,I1292908);
not I_59411 (I1012530,I1292908);
not I_59412 (I1012547,I1292917);
nand I_59413 (I1012564,I1292911,I1292905);
and I_59414 (I1012581,I1292911,I1292905);
not I_59415 (I1012598,I1292923);
nand I_59416 (I1012615,I1012598,I1012547);
nor I_59417 (I1012388,I1012615,I1012513);
nor I_59418 (I1012646,I1012530,I1012615);
nand I_59419 (I1012391,I1012581,I1012646);
not I_59420 (I1012677,I1292920);
nor I_59421 (I1012694,I1012677,I1292911);
nor I_59422 (I1012711,I1012694,I1292923);
nor I_59423 (I1012728,I1012479,I1012711);
DFFARX1 I_59424 (I1012728,I2507,I1012414,I1012400,);
not I_59425 (I1012759,I1012694);
DFFARX1 I_59426 (I1012759,I2507,I1012414,I1012403,);
and I_59427 (I1012397,I1012505,I1012694);
nor I_59428 (I1012804,I1012677,I1292914);
and I_59429 (I1012821,I1012804,I1292926);
or I_59430 (I1012838,I1012821,I1292902);
DFFARX1 I_59431 (I1012838,I2507,I1012414,I1012864,);
nor I_59432 (I1012872,I1012864,I1012598);
DFFARX1 I_59433 (I1012872,I2507,I1012414,I1012385,);
nand I_59434 (I1012903,I1012864,I1012505);
nand I_59435 (I1012920,I1012598,I1012903);
nor I_59436 (I1012394,I1012920,I1012564);
not I_59437 (I1012975,I2514);
DFFARX1 I_59438 (I552688,I2507,I1012975,I1013001,);
DFFARX1 I_59439 (I1013001,I2507,I1012975,I1013018,);
not I_59440 (I1012967,I1013018);
not I_59441 (I1013040,I1013001);
DFFARX1 I_59442 (I552703,I2507,I1012975,I1013066,);
nand I_59443 (I1013074,I1013066,I552694);
not I_59444 (I1013091,I552694);
not I_59445 (I1013108,I552700);
nand I_59446 (I1013125,I552697,I552706);
and I_59447 (I1013142,I552697,I552706);
not I_59448 (I1013159,I552691);
nand I_59449 (I1013176,I1013159,I1013108);
nor I_59450 (I1012949,I1013176,I1013074);
nor I_59451 (I1013207,I1013091,I1013176);
nand I_59452 (I1012952,I1013142,I1013207);
not I_59453 (I1013238,I552688);
nor I_59454 (I1013255,I1013238,I552697);
nor I_59455 (I1013272,I1013255,I552691);
nor I_59456 (I1013289,I1013040,I1013272);
DFFARX1 I_59457 (I1013289,I2507,I1012975,I1012961,);
not I_59458 (I1013320,I1013255);
DFFARX1 I_59459 (I1013320,I2507,I1012975,I1012964,);
and I_59460 (I1012958,I1013066,I1013255);
nor I_59461 (I1013365,I1013238,I552712);
and I_59462 (I1013382,I1013365,I552691);
or I_59463 (I1013399,I1013382,I552709);
DFFARX1 I_59464 (I1013399,I2507,I1012975,I1013425,);
nor I_59465 (I1013433,I1013425,I1013159);
DFFARX1 I_59466 (I1013433,I2507,I1012975,I1012946,);
nand I_59467 (I1013464,I1013425,I1013066);
nand I_59468 (I1013481,I1013159,I1013464);
nor I_59469 (I1012955,I1013481,I1013125);
not I_59470 (I1013536,I2514);
DFFARX1 I_59471 (I744587,I2507,I1013536,I1013562,);
DFFARX1 I_59472 (I1013562,I2507,I1013536,I1013579,);
not I_59473 (I1013528,I1013579);
not I_59474 (I1013601,I1013562);
DFFARX1 I_59475 (I744599,I2507,I1013536,I1013627,);
nand I_59476 (I1013635,I1013627,I744608);
not I_59477 (I1013652,I744608);
not I_59478 (I1013669,I744590);
nand I_59479 (I1013686,I744593,I744584);
and I_59480 (I1013703,I744593,I744584);
not I_59481 (I1013720,I744602);
nand I_59482 (I1013737,I1013720,I1013669);
nor I_59483 (I1013510,I1013737,I1013635);
nor I_59484 (I1013768,I1013652,I1013737);
nand I_59485 (I1013513,I1013703,I1013768);
not I_59486 (I1013799,I744605);
nor I_59487 (I1013816,I1013799,I744593);
nor I_59488 (I1013833,I1013816,I744602);
nor I_59489 (I1013850,I1013601,I1013833);
DFFARX1 I_59490 (I1013850,I2507,I1013536,I1013522,);
not I_59491 (I1013881,I1013816);
DFFARX1 I_59492 (I1013881,I2507,I1013536,I1013525,);
and I_59493 (I1013519,I1013627,I1013816);
nor I_59494 (I1013926,I1013799,I744584);
and I_59495 (I1013943,I1013926,I744596);
or I_59496 (I1013960,I1013943,I744587);
DFFARX1 I_59497 (I1013960,I2507,I1013536,I1013986,);
nor I_59498 (I1013994,I1013986,I1013720);
DFFARX1 I_59499 (I1013994,I2507,I1013536,I1013507,);
nand I_59500 (I1014025,I1013986,I1013627);
nand I_59501 (I1014042,I1013720,I1014025);
nor I_59502 (I1013516,I1014042,I1013686);
not I_59503 (I1014097,I2514);
DFFARX1 I_59504 (I979303,I2507,I1014097,I1014123,);
DFFARX1 I_59505 (I1014123,I2507,I1014097,I1014140,);
not I_59506 (I1014089,I1014140);
not I_59507 (I1014162,I1014123);
DFFARX1 I_59508 (I979330,I2507,I1014097,I1014188,);
nand I_59509 (I1014196,I1014188,I979321);
not I_59510 (I1014213,I979321);
not I_59511 (I1014230,I979303);
nand I_59512 (I1014247,I979315,I979318);
and I_59513 (I1014264,I979315,I979318);
not I_59514 (I1014281,I979327);
nand I_59515 (I1014298,I1014281,I1014230);
nor I_59516 (I1014071,I1014298,I1014196);
nor I_59517 (I1014329,I1014213,I1014298);
nand I_59518 (I1014074,I1014264,I1014329);
not I_59519 (I1014360,I979312);
nor I_59520 (I1014377,I1014360,I979315);
nor I_59521 (I1014394,I1014377,I979327);
nor I_59522 (I1014411,I1014162,I1014394);
DFFARX1 I_59523 (I1014411,I2507,I1014097,I1014083,);
not I_59524 (I1014442,I1014377);
DFFARX1 I_59525 (I1014442,I2507,I1014097,I1014086,);
and I_59526 (I1014080,I1014188,I1014377);
nor I_59527 (I1014487,I1014360,I979306);
and I_59528 (I1014504,I1014487,I979309);
or I_59529 (I1014521,I1014504,I979324);
DFFARX1 I_59530 (I1014521,I2507,I1014097,I1014547,);
nor I_59531 (I1014555,I1014547,I1014281);
DFFARX1 I_59532 (I1014555,I2507,I1014097,I1014068,);
nand I_59533 (I1014586,I1014547,I1014188);
nand I_59534 (I1014603,I1014281,I1014586);
nor I_59535 (I1014077,I1014603,I1014247);
not I_59536 (I1014658,I2514);
DFFARX1 I_59537 (I416967,I2507,I1014658,I1014684,);
DFFARX1 I_59538 (I1014684,I2507,I1014658,I1014701,);
not I_59539 (I1014650,I1014701);
not I_59540 (I1014723,I1014684);
DFFARX1 I_59541 (I416955,I2507,I1014658,I1014749,);
nand I_59542 (I1014757,I1014749,I416961);
not I_59543 (I1014774,I416961);
not I_59544 (I1014791,I416958);
nand I_59545 (I1014808,I416946,I416943);
and I_59546 (I1014825,I416946,I416943);
not I_59547 (I1014842,I416970);
nand I_59548 (I1014859,I1014842,I1014791);
nor I_59549 (I1014632,I1014859,I1014757);
nor I_59550 (I1014890,I1014774,I1014859);
nand I_59551 (I1014635,I1014825,I1014890);
not I_59552 (I1014921,I416943);
nor I_59553 (I1014938,I1014921,I416946);
nor I_59554 (I1014955,I1014938,I416970);
nor I_59555 (I1014972,I1014723,I1014955);
DFFARX1 I_59556 (I1014972,I2507,I1014658,I1014644,);
not I_59557 (I1015003,I1014938);
DFFARX1 I_59558 (I1015003,I2507,I1014658,I1014647,);
and I_59559 (I1014641,I1014749,I1014938);
nor I_59560 (I1015048,I1014921,I416952);
and I_59561 (I1015065,I1015048,I416949);
or I_59562 (I1015082,I1015065,I416964);
DFFARX1 I_59563 (I1015082,I2507,I1014658,I1015108,);
nor I_59564 (I1015116,I1015108,I1014842);
DFFARX1 I_59565 (I1015116,I2507,I1014658,I1014629,);
nand I_59566 (I1015147,I1015108,I1014749);
nand I_59567 (I1015164,I1014842,I1015147);
nor I_59568 (I1014638,I1015164,I1014808);
not I_59569 (I1015219,I2514);
DFFARX1 I_59570 (I1308897,I2507,I1015219,I1015245,);
DFFARX1 I_59571 (I1015245,I2507,I1015219,I1015262,);
not I_59572 (I1015211,I1015262);
not I_59573 (I1015284,I1015245);
DFFARX1 I_59574 (I1308891,I2507,I1015219,I1015310,);
nand I_59575 (I1015318,I1015310,I1308882);
not I_59576 (I1015335,I1308882);
not I_59577 (I1015352,I1308909);
nand I_59578 (I1015369,I1308894,I1308903);
and I_59579 (I1015386,I1308894,I1308903);
not I_59580 (I1015403,I1308888);
nand I_59581 (I1015420,I1015403,I1015352);
nor I_59582 (I1015193,I1015420,I1015318);
nor I_59583 (I1015451,I1015335,I1015420);
nand I_59584 (I1015196,I1015386,I1015451);
not I_59585 (I1015482,I1308906);
nor I_59586 (I1015499,I1015482,I1308894);
nor I_59587 (I1015516,I1015499,I1308888);
nor I_59588 (I1015533,I1015284,I1015516);
DFFARX1 I_59589 (I1015533,I2507,I1015219,I1015205,);
not I_59590 (I1015564,I1015499);
DFFARX1 I_59591 (I1015564,I2507,I1015219,I1015208,);
and I_59592 (I1015202,I1015310,I1015499);
nor I_59593 (I1015609,I1015482,I1308900);
and I_59594 (I1015626,I1015609,I1308882);
or I_59595 (I1015643,I1015626,I1308885);
DFFARX1 I_59596 (I1015643,I2507,I1015219,I1015669,);
nor I_59597 (I1015677,I1015669,I1015403);
DFFARX1 I_59598 (I1015677,I2507,I1015219,I1015190,);
nand I_59599 (I1015708,I1015669,I1015310);
nand I_59600 (I1015725,I1015403,I1015708);
nor I_59601 (I1015199,I1015725,I1015369);
not I_59602 (I1015780,I2514);
DFFARX1 I_59603 (I775799,I2507,I1015780,I1015806,);
DFFARX1 I_59604 (I1015806,I2507,I1015780,I1015823,);
not I_59605 (I1015772,I1015823);
not I_59606 (I1015845,I1015806);
DFFARX1 I_59607 (I775811,I2507,I1015780,I1015871,);
nand I_59608 (I1015879,I1015871,I775820);
not I_59609 (I1015896,I775820);
not I_59610 (I1015913,I775802);
nand I_59611 (I1015930,I775805,I775796);
and I_59612 (I1015947,I775805,I775796);
not I_59613 (I1015964,I775814);
nand I_59614 (I1015981,I1015964,I1015913);
nor I_59615 (I1015754,I1015981,I1015879);
nor I_59616 (I1016012,I1015896,I1015981);
nand I_59617 (I1015757,I1015947,I1016012);
not I_59618 (I1016043,I775817);
nor I_59619 (I1016060,I1016043,I775805);
nor I_59620 (I1016077,I1016060,I775814);
nor I_59621 (I1016094,I1015845,I1016077);
DFFARX1 I_59622 (I1016094,I2507,I1015780,I1015766,);
not I_59623 (I1016125,I1016060);
DFFARX1 I_59624 (I1016125,I2507,I1015780,I1015769,);
and I_59625 (I1015763,I1015871,I1016060);
nor I_59626 (I1016170,I1016043,I775796);
and I_59627 (I1016187,I1016170,I775808);
or I_59628 (I1016204,I1016187,I775799);
DFFARX1 I_59629 (I1016204,I2507,I1015780,I1016230,);
nor I_59630 (I1016238,I1016230,I1015964);
DFFARX1 I_59631 (I1016238,I2507,I1015780,I1015751,);
nand I_59632 (I1016269,I1016230,I1015871);
nand I_59633 (I1016286,I1015964,I1016269);
nor I_59634 (I1015760,I1016286,I1015930);
not I_59635 (I1016341,I2514);
DFFARX1 I_59636 (I119166,I2507,I1016341,I1016367,);
DFFARX1 I_59637 (I1016367,I2507,I1016341,I1016384,);
not I_59638 (I1016333,I1016384);
not I_59639 (I1016406,I1016367);
DFFARX1 I_59640 (I119154,I2507,I1016341,I1016432,);
nand I_59641 (I1016440,I1016432,I119169);
not I_59642 (I1016457,I119169);
not I_59643 (I1016474,I119157);
nand I_59644 (I1016491,I119178,I119172);
and I_59645 (I1016508,I119178,I119172);
not I_59646 (I1016525,I119160);
nand I_59647 (I1016542,I1016525,I1016474);
nor I_59648 (I1016315,I1016542,I1016440);
nor I_59649 (I1016573,I1016457,I1016542);
nand I_59650 (I1016318,I1016508,I1016573);
not I_59651 (I1016604,I119163);
nor I_59652 (I1016621,I1016604,I119178);
nor I_59653 (I1016638,I1016621,I119160);
nor I_59654 (I1016655,I1016406,I1016638);
DFFARX1 I_59655 (I1016655,I2507,I1016341,I1016327,);
not I_59656 (I1016686,I1016621);
DFFARX1 I_59657 (I1016686,I2507,I1016341,I1016330,);
and I_59658 (I1016324,I1016432,I1016621);
nor I_59659 (I1016731,I1016604,I119157);
and I_59660 (I1016748,I1016731,I119154);
or I_59661 (I1016765,I1016748,I119175);
DFFARX1 I_59662 (I1016765,I2507,I1016341,I1016791,);
nor I_59663 (I1016799,I1016791,I1016525);
DFFARX1 I_59664 (I1016799,I2507,I1016341,I1016312,);
nand I_59665 (I1016830,I1016791,I1016432);
nand I_59666 (I1016847,I1016525,I1016830);
nor I_59667 (I1016321,I1016847,I1016491);
not I_59668 (I1016902,I2514);
DFFARX1 I_59669 (I927623,I2507,I1016902,I1016928,);
DFFARX1 I_59670 (I1016928,I2507,I1016902,I1016945,);
not I_59671 (I1016894,I1016945);
not I_59672 (I1016967,I1016928);
DFFARX1 I_59673 (I927650,I2507,I1016902,I1016993,);
nand I_59674 (I1017001,I1016993,I927641);
not I_59675 (I1017018,I927641);
not I_59676 (I1017035,I927623);
nand I_59677 (I1017052,I927635,I927638);
and I_59678 (I1017069,I927635,I927638);
not I_59679 (I1017086,I927647);
nand I_59680 (I1017103,I1017086,I1017035);
nor I_59681 (I1016876,I1017103,I1017001);
nor I_59682 (I1017134,I1017018,I1017103);
nand I_59683 (I1016879,I1017069,I1017134);
not I_59684 (I1017165,I927632);
nor I_59685 (I1017182,I1017165,I927635);
nor I_59686 (I1017199,I1017182,I927647);
nor I_59687 (I1017216,I1016967,I1017199);
DFFARX1 I_59688 (I1017216,I2507,I1016902,I1016888,);
not I_59689 (I1017247,I1017182);
DFFARX1 I_59690 (I1017247,I2507,I1016902,I1016891,);
and I_59691 (I1016885,I1016993,I1017182);
nor I_59692 (I1017292,I1017165,I927626);
and I_59693 (I1017309,I1017292,I927629);
or I_59694 (I1017326,I1017309,I927644);
DFFARX1 I_59695 (I1017326,I2507,I1016902,I1017352,);
nor I_59696 (I1017360,I1017352,I1017086);
DFFARX1 I_59697 (I1017360,I2507,I1016902,I1016873,);
nand I_59698 (I1017391,I1017352,I1016993);
nand I_59699 (I1017408,I1017086,I1017391);
nor I_59700 (I1016882,I1017408,I1017052);
not I_59701 (I1017463,I2514);
DFFARX1 I_59702 (I1068789,I2507,I1017463,I1017489,);
DFFARX1 I_59703 (I1017489,I2507,I1017463,I1017506,);
not I_59704 (I1017455,I1017506);
not I_59705 (I1017528,I1017489);
DFFARX1 I_59706 (I1068780,I2507,I1017463,I1017554,);
nand I_59707 (I1017562,I1017554,I1068777);
not I_59708 (I1017579,I1068777);
not I_59709 (I1017596,I1068786);
nand I_59710 (I1017613,I1068795,I1068777);
and I_59711 (I1017630,I1068795,I1068777);
not I_59712 (I1017647,I1068774);
nand I_59713 (I1017664,I1017647,I1017596);
nor I_59714 (I1017437,I1017664,I1017562);
nor I_59715 (I1017695,I1017579,I1017664);
nand I_59716 (I1017440,I1017630,I1017695);
not I_59717 (I1017726,I1068783);
nor I_59718 (I1017743,I1017726,I1068795);
nor I_59719 (I1017760,I1017743,I1068774);
nor I_59720 (I1017777,I1017528,I1017760);
DFFARX1 I_59721 (I1017777,I2507,I1017463,I1017449,);
not I_59722 (I1017808,I1017743);
DFFARX1 I_59723 (I1017808,I2507,I1017463,I1017452,);
and I_59724 (I1017446,I1017554,I1017743);
nor I_59725 (I1017853,I1017726,I1068798);
and I_59726 (I1017870,I1017853,I1068774);
or I_59727 (I1017887,I1017870,I1068792);
DFFARX1 I_59728 (I1017887,I2507,I1017463,I1017913,);
nor I_59729 (I1017921,I1017913,I1017647);
DFFARX1 I_59730 (I1017921,I2507,I1017463,I1017434,);
nand I_59731 (I1017952,I1017913,I1017554);
nand I_59732 (I1017969,I1017647,I1017952);
nor I_59733 (I1017443,I1017969,I1017613);
not I_59734 (I1018024,I2514);
DFFARX1 I_59735 (I513742,I2507,I1018024,I1018050,);
DFFARX1 I_59736 (I1018050,I2507,I1018024,I1018067,);
not I_59737 (I1018016,I1018067);
not I_59738 (I1018089,I1018050);
DFFARX1 I_59739 (I513739,I2507,I1018024,I1018115,);
nand I_59740 (I1018123,I1018115,I513733);
not I_59741 (I1018140,I513733);
not I_59742 (I1018157,I513745);
nand I_59743 (I1018174,I513748,I513727);
and I_59744 (I1018191,I513748,I513727);
not I_59745 (I1018208,I513724);
nand I_59746 (I1018225,I1018208,I1018157);
nor I_59747 (I1017998,I1018225,I1018123);
nor I_59748 (I1018256,I1018140,I1018225);
nand I_59749 (I1018001,I1018191,I1018256);
not I_59750 (I1018287,I513730);
nor I_59751 (I1018304,I1018287,I513748);
nor I_59752 (I1018321,I1018304,I513724);
nor I_59753 (I1018338,I1018089,I1018321);
DFFARX1 I_59754 (I1018338,I2507,I1018024,I1018010,);
not I_59755 (I1018369,I1018304);
DFFARX1 I_59756 (I1018369,I2507,I1018024,I1018013,);
and I_59757 (I1018007,I1018115,I1018304);
nor I_59758 (I1018414,I1018287,I513724);
and I_59759 (I1018431,I1018414,I513736);
or I_59760 (I1018448,I1018431,I513727);
DFFARX1 I_59761 (I1018448,I2507,I1018024,I1018474,);
nor I_59762 (I1018482,I1018474,I1018208);
DFFARX1 I_59763 (I1018482,I2507,I1018024,I1017995,);
nand I_59764 (I1018513,I1018474,I1018115);
nand I_59765 (I1018530,I1018208,I1018513);
nor I_59766 (I1018004,I1018530,I1018174);
not I_59767 (I1018585,I2514);
DFFARX1 I_59768 (I441991,I2507,I1018585,I1018611,);
DFFARX1 I_59769 (I1018611,I2507,I1018585,I1018628,);
not I_59770 (I1018577,I1018628);
not I_59771 (I1018650,I1018611);
DFFARX1 I_59772 (I441979,I2507,I1018585,I1018676,);
nand I_59773 (I1018684,I1018676,I441985);
not I_59774 (I1018701,I441985);
not I_59775 (I1018718,I441982);
nand I_59776 (I1018735,I441970,I441967);
and I_59777 (I1018752,I441970,I441967);
not I_59778 (I1018769,I441994);
nand I_59779 (I1018786,I1018769,I1018718);
nor I_59780 (I1018559,I1018786,I1018684);
nor I_59781 (I1018817,I1018701,I1018786);
nand I_59782 (I1018562,I1018752,I1018817);
not I_59783 (I1018848,I441967);
nor I_59784 (I1018865,I1018848,I441970);
nor I_59785 (I1018882,I1018865,I441994);
nor I_59786 (I1018899,I1018650,I1018882);
DFFARX1 I_59787 (I1018899,I2507,I1018585,I1018571,);
not I_59788 (I1018930,I1018865);
DFFARX1 I_59789 (I1018930,I2507,I1018585,I1018574,);
and I_59790 (I1018568,I1018676,I1018865);
nor I_59791 (I1018975,I1018848,I441976);
and I_59792 (I1018992,I1018975,I441973);
or I_59793 (I1019009,I1018992,I441988);
DFFARX1 I_59794 (I1019009,I2507,I1018585,I1019035,);
nor I_59795 (I1019043,I1019035,I1018769);
DFFARX1 I_59796 (I1019043,I2507,I1018585,I1018556,);
nand I_59797 (I1019074,I1019035,I1018676);
nand I_59798 (I1019091,I1018769,I1019074);
nor I_59799 (I1018565,I1019091,I1018735);
not I_59800 (I1019146,I2514);
DFFARX1 I_59801 (I763661,I2507,I1019146,I1019172,);
DFFARX1 I_59802 (I1019172,I2507,I1019146,I1019189,);
not I_59803 (I1019138,I1019189);
not I_59804 (I1019211,I1019172);
DFFARX1 I_59805 (I763673,I2507,I1019146,I1019237,);
nand I_59806 (I1019245,I1019237,I763682);
not I_59807 (I1019262,I763682);
not I_59808 (I1019279,I763664);
nand I_59809 (I1019296,I763667,I763658);
and I_59810 (I1019313,I763667,I763658);
not I_59811 (I1019330,I763676);
nand I_59812 (I1019347,I1019330,I1019279);
nor I_59813 (I1019120,I1019347,I1019245);
nor I_59814 (I1019378,I1019262,I1019347);
nand I_59815 (I1019123,I1019313,I1019378);
not I_59816 (I1019409,I763679);
nor I_59817 (I1019426,I1019409,I763667);
nor I_59818 (I1019443,I1019426,I763676);
nor I_59819 (I1019460,I1019211,I1019443);
DFFARX1 I_59820 (I1019460,I2507,I1019146,I1019132,);
not I_59821 (I1019491,I1019426);
DFFARX1 I_59822 (I1019491,I2507,I1019146,I1019135,);
and I_59823 (I1019129,I1019237,I1019426);
nor I_59824 (I1019536,I1019409,I763658);
and I_59825 (I1019553,I1019536,I763670);
or I_59826 (I1019570,I1019553,I763661);
DFFARX1 I_59827 (I1019570,I2507,I1019146,I1019596,);
nor I_59828 (I1019604,I1019596,I1019330);
DFFARX1 I_59829 (I1019604,I2507,I1019146,I1019117,);
nand I_59830 (I1019635,I1019596,I1019237);
nand I_59831 (I1019652,I1019330,I1019635);
nor I_59832 (I1019126,I1019652,I1019296);
not I_59833 (I1019707,I2514);
DFFARX1 I_59834 (I1067055,I2507,I1019707,I1019733,);
DFFARX1 I_59835 (I1019733,I2507,I1019707,I1019750,);
not I_59836 (I1019699,I1019750);
not I_59837 (I1019772,I1019733);
DFFARX1 I_59838 (I1067046,I2507,I1019707,I1019798,);
nand I_59839 (I1019806,I1019798,I1067043);
not I_59840 (I1019823,I1067043);
not I_59841 (I1019840,I1067052);
nand I_59842 (I1019857,I1067061,I1067043);
and I_59843 (I1019874,I1067061,I1067043);
not I_59844 (I1019891,I1067040);
nand I_59845 (I1019908,I1019891,I1019840);
nor I_59846 (I1019681,I1019908,I1019806);
nor I_59847 (I1019939,I1019823,I1019908);
nand I_59848 (I1019684,I1019874,I1019939);
not I_59849 (I1019970,I1067049);
nor I_59850 (I1019987,I1019970,I1067061);
nor I_59851 (I1020004,I1019987,I1067040);
nor I_59852 (I1020021,I1019772,I1020004);
DFFARX1 I_59853 (I1020021,I2507,I1019707,I1019693,);
not I_59854 (I1020052,I1019987);
DFFARX1 I_59855 (I1020052,I2507,I1019707,I1019696,);
and I_59856 (I1019690,I1019798,I1019987);
nor I_59857 (I1020097,I1019970,I1067064);
and I_59858 (I1020114,I1020097,I1067040);
or I_59859 (I1020131,I1020114,I1067058);
DFFARX1 I_59860 (I1020131,I2507,I1019707,I1020157,);
nor I_59861 (I1020165,I1020157,I1019891);
DFFARX1 I_59862 (I1020165,I2507,I1019707,I1019678,);
nand I_59863 (I1020196,I1020157,I1019798);
nand I_59864 (I1020213,I1019891,I1020196);
nor I_59865 (I1019687,I1020213,I1019857);
not I_59866 (I1020268,I2514);
DFFARX1 I_59867 (I718577,I2507,I1020268,I1020294,);
DFFARX1 I_59868 (I1020294,I2507,I1020268,I1020311,);
not I_59869 (I1020260,I1020311);
not I_59870 (I1020333,I1020294);
DFFARX1 I_59871 (I718589,I2507,I1020268,I1020359,);
nand I_59872 (I1020367,I1020359,I718598);
not I_59873 (I1020384,I718598);
not I_59874 (I1020401,I718580);
nand I_59875 (I1020418,I718583,I718574);
and I_59876 (I1020435,I718583,I718574);
not I_59877 (I1020452,I718592);
nand I_59878 (I1020469,I1020452,I1020401);
nor I_59879 (I1020242,I1020469,I1020367);
nor I_59880 (I1020500,I1020384,I1020469);
nand I_59881 (I1020245,I1020435,I1020500);
not I_59882 (I1020531,I718595);
nor I_59883 (I1020548,I1020531,I718583);
nor I_59884 (I1020565,I1020548,I718592);
nor I_59885 (I1020582,I1020333,I1020565);
DFFARX1 I_59886 (I1020582,I2507,I1020268,I1020254,);
not I_59887 (I1020613,I1020548);
DFFARX1 I_59888 (I1020613,I2507,I1020268,I1020257,);
and I_59889 (I1020251,I1020359,I1020548);
nor I_59890 (I1020658,I1020531,I718574);
and I_59891 (I1020675,I1020658,I718586);
or I_59892 (I1020692,I1020675,I718577);
DFFARX1 I_59893 (I1020692,I2507,I1020268,I1020718,);
nor I_59894 (I1020726,I1020718,I1020452);
DFFARX1 I_59895 (I1020726,I2507,I1020268,I1020239,);
nand I_59896 (I1020757,I1020718,I1020359);
nand I_59897 (I1020774,I1020452,I1020757);
nor I_59898 (I1020248,I1020774,I1020418);
not I_59899 (I1020829,I2514);
DFFARX1 I_59900 (I908243,I2507,I1020829,I1020855,);
DFFARX1 I_59901 (I1020855,I2507,I1020829,I1020872,);
not I_59902 (I1020821,I1020872);
not I_59903 (I1020894,I1020855);
DFFARX1 I_59904 (I908270,I2507,I1020829,I1020920,);
nand I_59905 (I1020928,I1020920,I908261);
not I_59906 (I1020945,I908261);
not I_59907 (I1020962,I908243);
nand I_59908 (I1020979,I908255,I908258);
and I_59909 (I1020996,I908255,I908258);
not I_59910 (I1021013,I908267);
nand I_59911 (I1021030,I1021013,I1020962);
nor I_59912 (I1020803,I1021030,I1020928);
nor I_59913 (I1021061,I1020945,I1021030);
nand I_59914 (I1020806,I1020996,I1021061);
not I_59915 (I1021092,I908252);
nor I_59916 (I1021109,I1021092,I908255);
nor I_59917 (I1021126,I1021109,I908267);
nor I_59918 (I1021143,I1020894,I1021126);
DFFARX1 I_59919 (I1021143,I2507,I1020829,I1020815,);
not I_59920 (I1021174,I1021109);
DFFARX1 I_59921 (I1021174,I2507,I1020829,I1020818,);
and I_59922 (I1020812,I1020920,I1021109);
nor I_59923 (I1021219,I1021092,I908246);
and I_59924 (I1021236,I1021219,I908249);
or I_59925 (I1021253,I1021236,I908264);
DFFARX1 I_59926 (I1021253,I2507,I1020829,I1021279,);
nor I_59927 (I1021287,I1021279,I1021013);
DFFARX1 I_59928 (I1021287,I2507,I1020829,I1020800,);
nand I_59929 (I1021318,I1021279,I1020920);
nand I_59930 (I1021335,I1021013,I1021318);
nor I_59931 (I1020809,I1021335,I1020979);
not I_59932 (I1021390,I2514);
DFFARX1 I_59933 (I178198,I2507,I1021390,I1021416,);
DFFARX1 I_59934 (I1021416,I2507,I1021390,I1021433,);
not I_59935 (I1021382,I1021433);
not I_59936 (I1021455,I1021416);
DFFARX1 I_59937 (I178213,I2507,I1021390,I1021481,);
nand I_59938 (I1021489,I1021481,I178195);
not I_59939 (I1021506,I178195);
not I_59940 (I1021523,I178204);
nand I_59941 (I1021540,I178210,I178201);
and I_59942 (I1021557,I178210,I178201);
not I_59943 (I1021574,I178198);
nand I_59944 (I1021591,I1021574,I1021523);
nor I_59945 (I1021364,I1021591,I1021489);
nor I_59946 (I1021622,I1021506,I1021591);
nand I_59947 (I1021367,I1021557,I1021622);
not I_59948 (I1021653,I178195);
nor I_59949 (I1021670,I1021653,I178210);
nor I_59950 (I1021687,I1021670,I178198);
nor I_59951 (I1021704,I1021455,I1021687);
DFFARX1 I_59952 (I1021704,I2507,I1021390,I1021376,);
not I_59953 (I1021735,I1021670);
DFFARX1 I_59954 (I1021735,I2507,I1021390,I1021379,);
and I_59955 (I1021373,I1021481,I1021670);
nor I_59956 (I1021780,I1021653,I178219);
and I_59957 (I1021797,I1021780,I178216);
or I_59958 (I1021814,I1021797,I178207);
DFFARX1 I_59959 (I1021814,I2507,I1021390,I1021840,);
nor I_59960 (I1021848,I1021840,I1021574);
DFFARX1 I_59961 (I1021848,I2507,I1021390,I1021361,);
nand I_59962 (I1021879,I1021840,I1021481);
nand I_59963 (I1021896,I1021574,I1021879);
nor I_59964 (I1021370,I1021896,I1021540);
not I_59965 (I1021951,I2514);
DFFARX1 I_59966 (I764239,I2507,I1021951,I1021977,);
DFFARX1 I_59967 (I1021977,I2507,I1021951,I1021994,);
not I_59968 (I1021943,I1021994);
not I_59969 (I1022016,I1021977);
DFFARX1 I_59970 (I764251,I2507,I1021951,I1022042,);
nand I_59971 (I1022050,I1022042,I764260);
not I_59972 (I1022067,I764260);
not I_59973 (I1022084,I764242);
nand I_59974 (I1022101,I764245,I764236);
and I_59975 (I1022118,I764245,I764236);
not I_59976 (I1022135,I764254);
nand I_59977 (I1022152,I1022135,I1022084);
nor I_59978 (I1021925,I1022152,I1022050);
nor I_59979 (I1022183,I1022067,I1022152);
nand I_59980 (I1021928,I1022118,I1022183);
not I_59981 (I1022214,I764257);
nor I_59982 (I1022231,I1022214,I764245);
nor I_59983 (I1022248,I1022231,I764254);
nor I_59984 (I1022265,I1022016,I1022248);
DFFARX1 I_59985 (I1022265,I2507,I1021951,I1021937,);
not I_59986 (I1022296,I1022231);
DFFARX1 I_59987 (I1022296,I2507,I1021951,I1021940,);
and I_59988 (I1021934,I1022042,I1022231);
nor I_59989 (I1022341,I1022214,I764236);
and I_59990 (I1022358,I1022341,I764248);
or I_59991 (I1022375,I1022358,I764239);
DFFARX1 I_59992 (I1022375,I2507,I1021951,I1022401,);
nor I_59993 (I1022409,I1022401,I1022135);
DFFARX1 I_59994 (I1022409,I2507,I1021951,I1021922,);
nand I_59995 (I1022440,I1022401,I1022042);
nand I_59996 (I1022457,I1022135,I1022440);
nor I_59997 (I1021931,I1022457,I1022101);
not I_59998 (I1022512,I2514);
DFFARX1 I_59999 (I1345787,I2507,I1022512,I1022538,);
DFFARX1 I_60000 (I1022538,I2507,I1022512,I1022555,);
not I_60001 (I1022504,I1022555);
not I_60002 (I1022577,I1022538);
DFFARX1 I_60003 (I1345781,I2507,I1022512,I1022603,);
nand I_60004 (I1022611,I1022603,I1345772);
not I_60005 (I1022628,I1345772);
not I_60006 (I1022645,I1345799);
nand I_60007 (I1022662,I1345784,I1345793);
and I_60008 (I1022679,I1345784,I1345793);
not I_60009 (I1022696,I1345778);
nand I_60010 (I1022713,I1022696,I1022645);
nor I_60011 (I1022486,I1022713,I1022611);
nor I_60012 (I1022744,I1022628,I1022713);
nand I_60013 (I1022489,I1022679,I1022744);
not I_60014 (I1022775,I1345796);
nor I_60015 (I1022792,I1022775,I1345784);
nor I_60016 (I1022809,I1022792,I1345778);
nor I_60017 (I1022826,I1022577,I1022809);
DFFARX1 I_60018 (I1022826,I2507,I1022512,I1022498,);
not I_60019 (I1022857,I1022792);
DFFARX1 I_60020 (I1022857,I2507,I1022512,I1022501,);
and I_60021 (I1022495,I1022603,I1022792);
nor I_60022 (I1022902,I1022775,I1345790);
and I_60023 (I1022919,I1022902,I1345772);
or I_60024 (I1022936,I1022919,I1345775);
DFFARX1 I_60025 (I1022936,I2507,I1022512,I1022962,);
nor I_60026 (I1022970,I1022962,I1022696);
DFFARX1 I_60027 (I1022970,I2507,I1022512,I1022483,);
nand I_60028 (I1023001,I1022962,I1022603);
nand I_60029 (I1023018,I1022696,I1023001);
nor I_60030 (I1022492,I1023018,I1022662);
not I_60031 (I1023073,I2514);
DFFARX1 I_60032 (I1222120,I2507,I1023073,I1023099,);
DFFARX1 I_60033 (I1023099,I2507,I1023073,I1023116,);
not I_60034 (I1023065,I1023116);
not I_60035 (I1023138,I1023099);
DFFARX1 I_60036 (I1222126,I2507,I1023073,I1023164,);
nand I_60037 (I1023172,I1023164,I1222135);
not I_60038 (I1023189,I1222135);
not I_60039 (I1023206,I1222114);
nand I_60040 (I1023223,I1222117,I1222117);
and I_60041 (I1023240,I1222117,I1222117);
not I_60042 (I1023257,I1222129);
nand I_60043 (I1023274,I1023257,I1023206);
nor I_60044 (I1023047,I1023274,I1023172);
nor I_60045 (I1023305,I1023189,I1023274);
nand I_60046 (I1023050,I1023240,I1023305);
not I_60047 (I1023336,I1222123);
nor I_60048 (I1023353,I1023336,I1222117);
nor I_60049 (I1023370,I1023353,I1222129);
nor I_60050 (I1023387,I1023138,I1023370);
DFFARX1 I_60051 (I1023387,I2507,I1023073,I1023059,);
not I_60052 (I1023418,I1023353);
DFFARX1 I_60053 (I1023418,I2507,I1023073,I1023062,);
and I_60054 (I1023056,I1023164,I1023353);
nor I_60055 (I1023463,I1023336,I1222138);
and I_60056 (I1023480,I1023463,I1222114);
or I_60057 (I1023497,I1023480,I1222132);
DFFARX1 I_60058 (I1023497,I2507,I1023073,I1023523,);
nor I_60059 (I1023531,I1023523,I1023257);
DFFARX1 I_60060 (I1023531,I2507,I1023073,I1023044,);
nand I_60061 (I1023562,I1023523,I1023164);
nand I_60062 (I1023579,I1023257,I1023562);
nor I_60063 (I1023053,I1023579,I1023223);
not I_60064 (I1023634,I2514);
DFFARX1 I_60065 (I981887,I2507,I1023634,I1023660,);
DFFARX1 I_60066 (I1023660,I2507,I1023634,I1023677,);
not I_60067 (I1023626,I1023677);
not I_60068 (I1023699,I1023660);
DFFARX1 I_60069 (I981914,I2507,I1023634,I1023725,);
nand I_60070 (I1023733,I1023725,I981905);
not I_60071 (I1023750,I981905);
not I_60072 (I1023767,I981887);
nand I_60073 (I1023784,I981899,I981902);
and I_60074 (I1023801,I981899,I981902);
not I_60075 (I1023818,I981911);
nand I_60076 (I1023835,I1023818,I1023767);
nor I_60077 (I1023608,I1023835,I1023733);
nor I_60078 (I1023866,I1023750,I1023835);
nand I_60079 (I1023611,I1023801,I1023866);
not I_60080 (I1023897,I981896);
nor I_60081 (I1023914,I1023897,I981899);
nor I_60082 (I1023931,I1023914,I981911);
nor I_60083 (I1023948,I1023699,I1023931);
DFFARX1 I_60084 (I1023948,I2507,I1023634,I1023620,);
not I_60085 (I1023979,I1023914);
DFFARX1 I_60086 (I1023979,I2507,I1023634,I1023623,);
and I_60087 (I1023617,I1023725,I1023914);
nor I_60088 (I1024024,I1023897,I981890);
and I_60089 (I1024041,I1024024,I981893);
or I_60090 (I1024058,I1024041,I981908);
DFFARX1 I_60091 (I1024058,I2507,I1023634,I1024084,);
nor I_60092 (I1024092,I1024084,I1023818);
DFFARX1 I_60093 (I1024092,I2507,I1023634,I1023605,);
nand I_60094 (I1024123,I1024084,I1023725);
nand I_60095 (I1024140,I1023818,I1024123);
nor I_60096 (I1023614,I1024140,I1023784);
not I_60097 (I1024195,I2514);
DFFARX1 I_60098 (I552110,I2507,I1024195,I1024221,);
DFFARX1 I_60099 (I1024221,I2507,I1024195,I1024238,);
not I_60100 (I1024187,I1024238);
not I_60101 (I1024260,I1024221);
DFFARX1 I_60102 (I552125,I2507,I1024195,I1024286,);
nand I_60103 (I1024294,I1024286,I552116);
not I_60104 (I1024311,I552116);
not I_60105 (I1024328,I552122);
nand I_60106 (I1024345,I552119,I552128);
and I_60107 (I1024362,I552119,I552128);
not I_60108 (I1024379,I552113);
nand I_60109 (I1024396,I1024379,I1024328);
nor I_60110 (I1024169,I1024396,I1024294);
nor I_60111 (I1024427,I1024311,I1024396);
nand I_60112 (I1024172,I1024362,I1024427);
not I_60113 (I1024458,I552110);
nor I_60114 (I1024475,I1024458,I552119);
nor I_60115 (I1024492,I1024475,I552113);
nor I_60116 (I1024509,I1024260,I1024492);
DFFARX1 I_60117 (I1024509,I2507,I1024195,I1024181,);
not I_60118 (I1024540,I1024475);
DFFARX1 I_60119 (I1024540,I2507,I1024195,I1024184,);
and I_60120 (I1024178,I1024286,I1024475);
nor I_60121 (I1024585,I1024458,I552134);
and I_60122 (I1024602,I1024585,I552113);
or I_60123 (I1024619,I1024602,I552131);
DFFARX1 I_60124 (I1024619,I2507,I1024195,I1024645,);
nor I_60125 (I1024653,I1024645,I1024379);
DFFARX1 I_60126 (I1024653,I2507,I1024195,I1024166,);
nand I_60127 (I1024684,I1024645,I1024286);
nand I_60128 (I1024701,I1024379,I1024684);
nor I_60129 (I1024175,I1024701,I1024345);
not I_60130 (I1024756,I2514);
DFFARX1 I_60131 (I317140,I2507,I1024756,I1024782,);
DFFARX1 I_60132 (I1024782,I2507,I1024756,I1024799,);
not I_60133 (I1024748,I1024799);
not I_60134 (I1024821,I1024782);
DFFARX1 I_60135 (I317137,I2507,I1024756,I1024847,);
nand I_60136 (I1024855,I1024847,I317131);
not I_60137 (I1024872,I317131);
not I_60138 (I1024889,I317128);
nand I_60139 (I1024906,I317122,I317119);
and I_60140 (I1024923,I317122,I317119);
not I_60141 (I1024940,I317134);
nand I_60142 (I1024957,I1024940,I1024889);
nor I_60143 (I1024730,I1024957,I1024855);
nor I_60144 (I1024988,I1024872,I1024957);
nand I_60145 (I1024733,I1024923,I1024988);
not I_60146 (I1025019,I317146);
nor I_60147 (I1025036,I1025019,I317122);
nor I_60148 (I1025053,I1025036,I317134);
nor I_60149 (I1025070,I1024821,I1025053);
DFFARX1 I_60150 (I1025070,I2507,I1024756,I1024742,);
not I_60151 (I1025101,I1025036);
DFFARX1 I_60152 (I1025101,I2507,I1024756,I1024745,);
and I_60153 (I1024739,I1024847,I1025036);
nor I_60154 (I1025146,I1025019,I317143);
and I_60155 (I1025163,I1025146,I317119);
or I_60156 (I1025180,I1025163,I317125);
DFFARX1 I_60157 (I1025180,I2507,I1024756,I1025206,);
nor I_60158 (I1025214,I1025206,I1024940);
DFFARX1 I_60159 (I1025214,I2507,I1024756,I1024727,);
nand I_60160 (I1025245,I1025206,I1024847);
nand I_60161 (I1025262,I1024940,I1025245);
nor I_60162 (I1024736,I1025262,I1024906);
not I_60163 (I1025317,I2514);
DFFARX1 I_60164 (I1230280,I2507,I1025317,I1025343,);
DFFARX1 I_60165 (I1025343,I2507,I1025317,I1025360,);
not I_60166 (I1025309,I1025360);
not I_60167 (I1025382,I1025343);
DFFARX1 I_60168 (I1230286,I2507,I1025317,I1025408,);
nand I_60169 (I1025416,I1025408,I1230295);
not I_60170 (I1025433,I1230295);
not I_60171 (I1025450,I1230274);
nand I_60172 (I1025467,I1230277,I1230277);
and I_60173 (I1025484,I1230277,I1230277);
not I_60174 (I1025501,I1230289);
nand I_60175 (I1025518,I1025501,I1025450);
nor I_60176 (I1025291,I1025518,I1025416);
nor I_60177 (I1025549,I1025433,I1025518);
nand I_60178 (I1025294,I1025484,I1025549);
not I_60179 (I1025580,I1230283);
nor I_60180 (I1025597,I1025580,I1230277);
nor I_60181 (I1025614,I1025597,I1230289);
nor I_60182 (I1025631,I1025382,I1025614);
DFFARX1 I_60183 (I1025631,I2507,I1025317,I1025303,);
not I_60184 (I1025662,I1025597);
DFFARX1 I_60185 (I1025662,I2507,I1025317,I1025306,);
and I_60186 (I1025300,I1025408,I1025597);
nor I_60187 (I1025707,I1025580,I1230298);
and I_60188 (I1025724,I1025707,I1230274);
or I_60189 (I1025741,I1025724,I1230292);
DFFARX1 I_60190 (I1025741,I2507,I1025317,I1025767,);
nor I_60191 (I1025775,I1025767,I1025501);
DFFARX1 I_60192 (I1025775,I2507,I1025317,I1025288,);
nand I_60193 (I1025806,I1025767,I1025408);
nand I_60194 (I1025823,I1025501,I1025806);
nor I_60195 (I1025297,I1025823,I1025467);
not I_60196 (I1025878,I2514);
DFFARX1 I_60197 (I697769,I2507,I1025878,I1025904,);
DFFARX1 I_60198 (I1025904,I2507,I1025878,I1025921,);
not I_60199 (I1025870,I1025921);
not I_60200 (I1025943,I1025904);
DFFARX1 I_60201 (I697781,I2507,I1025878,I1025969,);
nand I_60202 (I1025977,I1025969,I697790);
not I_60203 (I1025994,I697790);
not I_60204 (I1026011,I697772);
nand I_60205 (I1026028,I697775,I697766);
and I_60206 (I1026045,I697775,I697766);
not I_60207 (I1026062,I697784);
nand I_60208 (I1026079,I1026062,I1026011);
nor I_60209 (I1025852,I1026079,I1025977);
nor I_60210 (I1026110,I1025994,I1026079);
nand I_60211 (I1025855,I1026045,I1026110);
not I_60212 (I1026141,I697787);
nor I_60213 (I1026158,I1026141,I697775);
nor I_60214 (I1026175,I1026158,I697784);
nor I_60215 (I1026192,I1025943,I1026175);
DFFARX1 I_60216 (I1026192,I2507,I1025878,I1025864,);
not I_60217 (I1026223,I1026158);
DFFARX1 I_60218 (I1026223,I2507,I1025878,I1025867,);
and I_60219 (I1025861,I1025969,I1026158);
nor I_60220 (I1026268,I1026141,I697766);
and I_60221 (I1026285,I1026268,I697778);
or I_60222 (I1026302,I1026285,I697769);
DFFARX1 I_60223 (I1026302,I2507,I1025878,I1026328,);
nor I_60224 (I1026336,I1026328,I1026062);
DFFARX1 I_60225 (I1026336,I2507,I1025878,I1025849,);
nand I_60226 (I1026367,I1026328,I1025969);
nand I_60227 (I1026384,I1026062,I1026367);
nor I_60228 (I1025858,I1026384,I1026028);
not I_60229 (I1026439,I2514);
DFFARX1 I_60230 (I185933,I2507,I1026439,I1026465,);
DFFARX1 I_60231 (I1026465,I2507,I1026439,I1026482,);
not I_60232 (I1026431,I1026482);
not I_60233 (I1026504,I1026465);
DFFARX1 I_60234 (I185948,I2507,I1026439,I1026530,);
nand I_60235 (I1026538,I1026530,I185930);
not I_60236 (I1026555,I185930);
not I_60237 (I1026572,I185939);
nand I_60238 (I1026589,I185945,I185936);
and I_60239 (I1026606,I185945,I185936);
not I_60240 (I1026623,I185933);
nand I_60241 (I1026640,I1026623,I1026572);
nor I_60242 (I1026413,I1026640,I1026538);
nor I_60243 (I1026671,I1026555,I1026640);
nand I_60244 (I1026416,I1026606,I1026671);
not I_60245 (I1026702,I185930);
nor I_60246 (I1026719,I1026702,I185945);
nor I_60247 (I1026736,I1026719,I185933);
nor I_60248 (I1026753,I1026504,I1026736);
DFFARX1 I_60249 (I1026753,I2507,I1026439,I1026425,);
not I_60250 (I1026784,I1026719);
DFFARX1 I_60251 (I1026784,I2507,I1026439,I1026428,);
and I_60252 (I1026422,I1026530,I1026719);
nor I_60253 (I1026829,I1026702,I185954);
and I_60254 (I1026846,I1026829,I185951);
or I_60255 (I1026863,I1026846,I185942);
DFFARX1 I_60256 (I1026863,I2507,I1026439,I1026889,);
nor I_60257 (I1026897,I1026889,I1026623);
DFFARX1 I_60258 (I1026897,I2507,I1026439,I1026410,);
nand I_60259 (I1026928,I1026889,I1026530);
nand I_60260 (I1026945,I1026623,I1026928);
nor I_60261 (I1026419,I1026945,I1026589);
not I_60262 (I1027000,I2514);
DFFARX1 I_60263 (I673493,I2507,I1027000,I1027026,);
DFFARX1 I_60264 (I1027026,I2507,I1027000,I1027043,);
not I_60265 (I1026992,I1027043);
not I_60266 (I1027065,I1027026);
DFFARX1 I_60267 (I673505,I2507,I1027000,I1027091,);
nand I_60268 (I1027099,I1027091,I673514);
not I_60269 (I1027116,I673514);
not I_60270 (I1027133,I673496);
nand I_60271 (I1027150,I673499,I673490);
and I_60272 (I1027167,I673499,I673490);
not I_60273 (I1027184,I673508);
nand I_60274 (I1027201,I1027184,I1027133);
nor I_60275 (I1026974,I1027201,I1027099);
nor I_60276 (I1027232,I1027116,I1027201);
nand I_60277 (I1026977,I1027167,I1027232);
not I_60278 (I1027263,I673511);
nor I_60279 (I1027280,I1027263,I673499);
nor I_60280 (I1027297,I1027280,I673508);
nor I_60281 (I1027314,I1027065,I1027297);
DFFARX1 I_60282 (I1027314,I2507,I1027000,I1026986,);
not I_60283 (I1027345,I1027280);
DFFARX1 I_60284 (I1027345,I2507,I1027000,I1026989,);
and I_60285 (I1026983,I1027091,I1027280);
nor I_60286 (I1027390,I1027263,I673490);
and I_60287 (I1027407,I1027390,I673502);
or I_60288 (I1027424,I1027407,I673493);
DFFARX1 I_60289 (I1027424,I2507,I1027000,I1027450,);
nor I_60290 (I1027458,I1027450,I1027184);
DFFARX1 I_60291 (I1027458,I2507,I1027000,I1026971,);
nand I_60292 (I1027489,I1027450,I1027091);
nand I_60293 (I1027506,I1027184,I1027489);
nor I_60294 (I1026980,I1027506,I1027150);
not I_60295 (I1027561,I2514);
DFFARX1 I_60296 (I149043,I2507,I1027561,I1027587,);
DFFARX1 I_60297 (I1027587,I2507,I1027561,I1027604,);
not I_60298 (I1027553,I1027604);
not I_60299 (I1027626,I1027587);
DFFARX1 I_60300 (I149058,I2507,I1027561,I1027652,);
nand I_60301 (I1027660,I1027652,I149040);
not I_60302 (I1027677,I149040);
not I_60303 (I1027694,I149049);
nand I_60304 (I1027711,I149055,I149046);
and I_60305 (I1027728,I149055,I149046);
not I_60306 (I1027745,I149043);
nand I_60307 (I1027762,I1027745,I1027694);
nor I_60308 (I1027535,I1027762,I1027660);
nor I_60309 (I1027793,I1027677,I1027762);
nand I_60310 (I1027538,I1027728,I1027793);
not I_60311 (I1027824,I149040);
nor I_60312 (I1027841,I1027824,I149055);
nor I_60313 (I1027858,I1027841,I149043);
nor I_60314 (I1027875,I1027626,I1027858);
DFFARX1 I_60315 (I1027875,I2507,I1027561,I1027547,);
not I_60316 (I1027906,I1027841);
DFFARX1 I_60317 (I1027906,I2507,I1027561,I1027550,);
and I_60318 (I1027544,I1027652,I1027841);
nor I_60319 (I1027951,I1027824,I149064);
and I_60320 (I1027968,I1027951,I149061);
or I_60321 (I1027985,I1027968,I149052);
DFFARX1 I_60322 (I1027985,I2507,I1027561,I1028011,);
nor I_60323 (I1028019,I1028011,I1027745);
DFFARX1 I_60324 (I1028019,I2507,I1027561,I1027532,);
nand I_60325 (I1028050,I1028011,I1027652);
nand I_60326 (I1028067,I1027745,I1028050);
nor I_60327 (I1027541,I1028067,I1027711);
not I_60328 (I1028122,I2514);
DFFARX1 I_60329 (I1233544,I2507,I1028122,I1028148,);
DFFARX1 I_60330 (I1028148,I2507,I1028122,I1028165,);
not I_60331 (I1028114,I1028165);
not I_60332 (I1028187,I1028148);
DFFARX1 I_60333 (I1233550,I2507,I1028122,I1028213,);
nand I_60334 (I1028221,I1028213,I1233559);
not I_60335 (I1028238,I1233559);
not I_60336 (I1028255,I1233538);
nand I_60337 (I1028272,I1233541,I1233541);
and I_60338 (I1028289,I1233541,I1233541);
not I_60339 (I1028306,I1233553);
nand I_60340 (I1028323,I1028306,I1028255);
nor I_60341 (I1028096,I1028323,I1028221);
nor I_60342 (I1028354,I1028238,I1028323);
nand I_60343 (I1028099,I1028289,I1028354);
not I_60344 (I1028385,I1233547);
nor I_60345 (I1028402,I1028385,I1233541);
nor I_60346 (I1028419,I1028402,I1233553);
nor I_60347 (I1028436,I1028187,I1028419);
DFFARX1 I_60348 (I1028436,I2507,I1028122,I1028108,);
not I_60349 (I1028467,I1028402);
DFFARX1 I_60350 (I1028467,I2507,I1028122,I1028111,);
and I_60351 (I1028105,I1028213,I1028402);
nor I_60352 (I1028512,I1028385,I1233562);
and I_60353 (I1028529,I1028512,I1233538);
or I_60354 (I1028546,I1028529,I1233556);
DFFARX1 I_60355 (I1028546,I2507,I1028122,I1028572,);
nor I_60356 (I1028580,I1028572,I1028306);
DFFARX1 I_60357 (I1028580,I2507,I1028122,I1028093,);
nand I_60358 (I1028611,I1028572,I1028213);
nand I_60359 (I1028628,I1028306,I1028611);
nor I_60360 (I1028102,I1028628,I1028272);
not I_60361 (I1028683,I2514);
DFFARX1 I_60362 (I538732,I2507,I1028683,I1028709,);
DFFARX1 I_60363 (I1028709,I2507,I1028683,I1028726,);
not I_60364 (I1028675,I1028726);
not I_60365 (I1028748,I1028709);
DFFARX1 I_60366 (I538729,I2507,I1028683,I1028774,);
nand I_60367 (I1028782,I1028774,I538723);
not I_60368 (I1028799,I538723);
not I_60369 (I1028816,I538735);
nand I_60370 (I1028833,I538738,I538717);
and I_60371 (I1028850,I538738,I538717);
not I_60372 (I1028867,I538714);
nand I_60373 (I1028884,I1028867,I1028816);
nor I_60374 (I1028657,I1028884,I1028782);
nor I_60375 (I1028915,I1028799,I1028884);
nand I_60376 (I1028660,I1028850,I1028915);
not I_60377 (I1028946,I538720);
nor I_60378 (I1028963,I1028946,I538738);
nor I_60379 (I1028980,I1028963,I538714);
nor I_60380 (I1028997,I1028748,I1028980);
DFFARX1 I_60381 (I1028997,I2507,I1028683,I1028669,);
not I_60382 (I1029028,I1028963);
DFFARX1 I_60383 (I1029028,I2507,I1028683,I1028672,);
and I_60384 (I1028666,I1028774,I1028963);
nor I_60385 (I1029073,I1028946,I538714);
and I_60386 (I1029090,I1029073,I538726);
or I_60387 (I1029107,I1029090,I538717);
DFFARX1 I_60388 (I1029107,I2507,I1028683,I1029133,);
nor I_60389 (I1029141,I1029133,I1028867);
DFFARX1 I_60390 (I1029141,I2507,I1028683,I1028654,);
nand I_60391 (I1029172,I1029133,I1028774);
nand I_60392 (I1029189,I1028867,I1029172);
nor I_60393 (I1028663,I1029189,I1028833);
not I_60394 (I1029244,I2514);
DFFARX1 I_60395 (I631299,I2507,I1029244,I1029270,);
DFFARX1 I_60396 (I1029270,I2507,I1029244,I1029287,);
not I_60397 (I1029236,I1029287);
not I_60398 (I1029309,I1029270);
DFFARX1 I_60399 (I631311,I2507,I1029244,I1029335,);
nand I_60400 (I1029343,I1029335,I631320);
not I_60401 (I1029360,I631320);
not I_60402 (I1029377,I631302);
nand I_60403 (I1029394,I631305,I631296);
and I_60404 (I1029411,I631305,I631296);
not I_60405 (I1029428,I631314);
nand I_60406 (I1029445,I1029428,I1029377);
nor I_60407 (I1029218,I1029445,I1029343);
nor I_60408 (I1029476,I1029360,I1029445);
nand I_60409 (I1029221,I1029411,I1029476);
not I_60410 (I1029507,I631317);
nor I_60411 (I1029524,I1029507,I631305);
nor I_60412 (I1029541,I1029524,I631314);
nor I_60413 (I1029558,I1029309,I1029541);
DFFARX1 I_60414 (I1029558,I2507,I1029244,I1029230,);
not I_60415 (I1029589,I1029524);
DFFARX1 I_60416 (I1029589,I2507,I1029244,I1029233,);
and I_60417 (I1029227,I1029335,I1029524);
nor I_60418 (I1029634,I1029507,I631296);
and I_60419 (I1029651,I1029634,I631308);
or I_60420 (I1029668,I1029651,I631299);
DFFARX1 I_60421 (I1029668,I2507,I1029244,I1029694,);
nor I_60422 (I1029702,I1029694,I1029428);
DFFARX1 I_60423 (I1029702,I2507,I1029244,I1029215,);
nand I_60424 (I1029733,I1029694,I1029335);
nand I_60425 (I1029750,I1029428,I1029733);
nor I_60426 (I1029224,I1029750,I1029394);
not I_60427 (I1029805,I2514);
DFFARX1 I_60428 (I612800,I2507,I1029805,I1029831,);
DFFARX1 I_60429 (I1029831,I2507,I1029805,I1029848,);
not I_60430 (I1029797,I1029848);
not I_60431 (I1029870,I1029831);
DFFARX1 I_60432 (I612815,I2507,I1029805,I1029896,);
nand I_60433 (I1029904,I1029896,I612806);
not I_60434 (I1029921,I612806);
not I_60435 (I1029938,I612812);
nand I_60436 (I1029955,I612809,I612818);
and I_60437 (I1029972,I612809,I612818);
not I_60438 (I1029989,I612803);
nand I_60439 (I1030006,I1029989,I1029938);
nor I_60440 (I1029779,I1030006,I1029904);
nor I_60441 (I1030037,I1029921,I1030006);
nand I_60442 (I1029782,I1029972,I1030037);
not I_60443 (I1030068,I612800);
nor I_60444 (I1030085,I1030068,I612809);
nor I_60445 (I1030102,I1030085,I612803);
nor I_60446 (I1030119,I1029870,I1030102);
DFFARX1 I_60447 (I1030119,I2507,I1029805,I1029791,);
not I_60448 (I1030150,I1030085);
DFFARX1 I_60449 (I1030150,I2507,I1029805,I1029794,);
and I_60450 (I1029788,I1029896,I1030085);
nor I_60451 (I1030195,I1030068,I612824);
and I_60452 (I1030212,I1030195,I612803);
or I_60453 (I1030229,I1030212,I612821);
DFFARX1 I_60454 (I1030229,I2507,I1029805,I1030255,);
nor I_60455 (I1030263,I1030255,I1029989);
DFFARX1 I_60456 (I1030263,I2507,I1029805,I1029776,);
nand I_60457 (I1030294,I1030255,I1029896);
nand I_60458 (I1030311,I1029989,I1030294);
nor I_60459 (I1029785,I1030311,I1029955);
not I_60460 (I1030366,I2514);
DFFARX1 I_60461 (I758459,I2507,I1030366,I1030392,);
DFFARX1 I_60462 (I1030392,I2507,I1030366,I1030409,);
not I_60463 (I1030358,I1030409);
not I_60464 (I1030431,I1030392);
DFFARX1 I_60465 (I758471,I2507,I1030366,I1030457,);
nand I_60466 (I1030465,I1030457,I758480);
not I_60467 (I1030482,I758480);
not I_60468 (I1030499,I758462);
nand I_60469 (I1030516,I758465,I758456);
and I_60470 (I1030533,I758465,I758456);
not I_60471 (I1030550,I758474);
nand I_60472 (I1030567,I1030550,I1030499);
nor I_60473 (I1030340,I1030567,I1030465);
nor I_60474 (I1030598,I1030482,I1030567);
nand I_60475 (I1030343,I1030533,I1030598);
not I_60476 (I1030629,I758477);
nor I_60477 (I1030646,I1030629,I758465);
nor I_60478 (I1030663,I1030646,I758474);
nor I_60479 (I1030680,I1030431,I1030663);
DFFARX1 I_60480 (I1030680,I2507,I1030366,I1030352,);
not I_60481 (I1030711,I1030646);
DFFARX1 I_60482 (I1030711,I2507,I1030366,I1030355,);
and I_60483 (I1030349,I1030457,I1030646);
nor I_60484 (I1030756,I1030629,I758456);
and I_60485 (I1030773,I1030756,I758468);
or I_60486 (I1030790,I1030773,I758459);
DFFARX1 I_60487 (I1030790,I2507,I1030366,I1030816,);
nor I_60488 (I1030824,I1030816,I1030550);
DFFARX1 I_60489 (I1030824,I2507,I1030366,I1030337,);
nand I_60490 (I1030855,I1030816,I1030457);
nand I_60491 (I1030872,I1030550,I1030855);
nor I_60492 (I1030346,I1030872,I1030516);
not I_60493 (I1030927,I2514);
DFFARX1 I_60494 (I285520,I2507,I1030927,I1030953,);
DFFARX1 I_60495 (I1030953,I2507,I1030927,I1030970,);
not I_60496 (I1030919,I1030970);
not I_60497 (I1030992,I1030953);
DFFARX1 I_60498 (I285517,I2507,I1030927,I1031018,);
nand I_60499 (I1031026,I1031018,I285511);
not I_60500 (I1031043,I285511);
not I_60501 (I1031060,I285508);
nand I_60502 (I1031077,I285502,I285499);
and I_60503 (I1031094,I285502,I285499);
not I_60504 (I1031111,I285514);
nand I_60505 (I1031128,I1031111,I1031060);
nor I_60506 (I1030901,I1031128,I1031026);
nor I_60507 (I1031159,I1031043,I1031128);
nand I_60508 (I1030904,I1031094,I1031159);
not I_60509 (I1031190,I285526);
nor I_60510 (I1031207,I1031190,I285502);
nor I_60511 (I1031224,I1031207,I285514);
nor I_60512 (I1031241,I1030992,I1031224);
DFFARX1 I_60513 (I1031241,I2507,I1030927,I1030913,);
not I_60514 (I1031272,I1031207);
DFFARX1 I_60515 (I1031272,I2507,I1030927,I1030916,);
and I_60516 (I1030910,I1031018,I1031207);
nor I_60517 (I1031317,I1031190,I285523);
and I_60518 (I1031334,I1031317,I285499);
or I_60519 (I1031351,I1031334,I285505);
DFFARX1 I_60520 (I1031351,I2507,I1030927,I1031377,);
nor I_60521 (I1031385,I1031377,I1031111);
DFFARX1 I_60522 (I1031385,I2507,I1030927,I1030898,);
nand I_60523 (I1031416,I1031377,I1031018);
nand I_60524 (I1031433,I1031111,I1031416);
nor I_60525 (I1030907,I1031433,I1031077);
not I_60526 (I1031488,I2514);
DFFARX1 I_60527 (I1181499,I2507,I1031488,I1031514,);
DFFARX1 I_60528 (I1031514,I2507,I1031488,I1031531,);
not I_60529 (I1031480,I1031531);
not I_60530 (I1031553,I1031514);
DFFARX1 I_60531 (I1181490,I2507,I1031488,I1031579,);
nand I_60532 (I1031587,I1031579,I1181487);
not I_60533 (I1031604,I1181487);
not I_60534 (I1031621,I1181496);
nand I_60535 (I1031638,I1181505,I1181487);
and I_60536 (I1031655,I1181505,I1181487);
not I_60537 (I1031672,I1181484);
nand I_60538 (I1031689,I1031672,I1031621);
nor I_60539 (I1031462,I1031689,I1031587);
nor I_60540 (I1031720,I1031604,I1031689);
nand I_60541 (I1031465,I1031655,I1031720);
not I_60542 (I1031751,I1181493);
nor I_60543 (I1031768,I1031751,I1181505);
nor I_60544 (I1031785,I1031768,I1181484);
nor I_60545 (I1031802,I1031553,I1031785);
DFFARX1 I_60546 (I1031802,I2507,I1031488,I1031474,);
not I_60547 (I1031833,I1031768);
DFFARX1 I_60548 (I1031833,I2507,I1031488,I1031477,);
and I_60549 (I1031471,I1031579,I1031768);
nor I_60550 (I1031878,I1031751,I1181508);
and I_60551 (I1031895,I1031878,I1181484);
or I_60552 (I1031912,I1031895,I1181502);
DFFARX1 I_60553 (I1031912,I2507,I1031488,I1031938,);
nor I_60554 (I1031946,I1031938,I1031672);
DFFARX1 I_60555 (I1031946,I2507,I1031488,I1031459,);
nand I_60556 (I1031977,I1031938,I1031579);
nand I_60557 (I1031994,I1031672,I1031977);
nor I_60558 (I1031468,I1031994,I1031638);
not I_60559 (I1032049,I2514);
DFFARX1 I_60560 (I1090753,I2507,I1032049,I1032075,);
DFFARX1 I_60561 (I1032075,I2507,I1032049,I1032092,);
not I_60562 (I1032041,I1032092);
not I_60563 (I1032114,I1032075);
DFFARX1 I_60564 (I1090744,I2507,I1032049,I1032140,);
nand I_60565 (I1032148,I1032140,I1090741);
not I_60566 (I1032165,I1090741);
not I_60567 (I1032182,I1090750);
nand I_60568 (I1032199,I1090759,I1090741);
and I_60569 (I1032216,I1090759,I1090741);
not I_60570 (I1032233,I1090738);
nand I_60571 (I1032250,I1032233,I1032182);
nor I_60572 (I1032023,I1032250,I1032148);
nor I_60573 (I1032281,I1032165,I1032250);
nand I_60574 (I1032026,I1032216,I1032281);
not I_60575 (I1032312,I1090747);
nor I_60576 (I1032329,I1032312,I1090759);
nor I_60577 (I1032346,I1032329,I1090738);
nor I_60578 (I1032363,I1032114,I1032346);
DFFARX1 I_60579 (I1032363,I2507,I1032049,I1032035,);
not I_60580 (I1032394,I1032329);
DFFARX1 I_60581 (I1032394,I2507,I1032049,I1032038,);
and I_60582 (I1032032,I1032140,I1032329);
nor I_60583 (I1032439,I1032312,I1090762);
and I_60584 (I1032456,I1032439,I1090738);
or I_60585 (I1032473,I1032456,I1090756);
DFFARX1 I_60586 (I1032473,I2507,I1032049,I1032499,);
nor I_60587 (I1032507,I1032499,I1032233);
DFFARX1 I_60588 (I1032507,I2507,I1032049,I1032020,);
nand I_60589 (I1032538,I1032499,I1032140);
nand I_60590 (I1032555,I1032233,I1032538);
nor I_60591 (I1032029,I1032555,I1032199);
not I_60592 (I1032610,I2514);
DFFARX1 I_60593 (I133395,I2507,I1032610,I1032636,);
DFFARX1 I_60594 (I1032636,I2507,I1032610,I1032653,);
not I_60595 (I1032602,I1032653);
not I_60596 (I1032675,I1032636);
DFFARX1 I_60597 (I133383,I2507,I1032610,I1032701,);
nand I_60598 (I1032709,I1032701,I133398);
not I_60599 (I1032726,I133398);
not I_60600 (I1032743,I133386);
nand I_60601 (I1032760,I133407,I133401);
and I_60602 (I1032777,I133407,I133401);
not I_60603 (I1032794,I133389);
nand I_60604 (I1032811,I1032794,I1032743);
nor I_60605 (I1032584,I1032811,I1032709);
nor I_60606 (I1032842,I1032726,I1032811);
nand I_60607 (I1032587,I1032777,I1032842);
not I_60608 (I1032873,I133392);
nor I_60609 (I1032890,I1032873,I133407);
nor I_60610 (I1032907,I1032890,I133389);
nor I_60611 (I1032924,I1032675,I1032907);
DFFARX1 I_60612 (I1032924,I2507,I1032610,I1032596,);
not I_60613 (I1032955,I1032890);
DFFARX1 I_60614 (I1032955,I2507,I1032610,I1032599,);
and I_60615 (I1032593,I1032701,I1032890);
nor I_60616 (I1033000,I1032873,I133386);
and I_60617 (I1033017,I1033000,I133383);
or I_60618 (I1033034,I1033017,I133404);
DFFARX1 I_60619 (I1033034,I2507,I1032610,I1033060,);
nor I_60620 (I1033068,I1033060,I1032794);
DFFARX1 I_60621 (I1033068,I2507,I1032610,I1032581,);
nand I_60622 (I1033099,I1033060,I1032701);
nand I_60623 (I1033116,I1032794,I1033099);
nor I_60624 (I1032590,I1033116,I1032760);
not I_60625 (I1033171,I2514);
DFFARX1 I_60626 (I567138,I2507,I1033171,I1033197,);
DFFARX1 I_60627 (I1033197,I2507,I1033171,I1033214,);
not I_60628 (I1033163,I1033214);
not I_60629 (I1033236,I1033197);
DFFARX1 I_60630 (I567153,I2507,I1033171,I1033262,);
nand I_60631 (I1033270,I1033262,I567144);
not I_60632 (I1033287,I567144);
not I_60633 (I1033304,I567150);
nand I_60634 (I1033321,I567147,I567156);
and I_60635 (I1033338,I567147,I567156);
not I_60636 (I1033355,I567141);
nand I_60637 (I1033372,I1033355,I1033304);
nor I_60638 (I1033145,I1033372,I1033270);
nor I_60639 (I1033403,I1033287,I1033372);
nand I_60640 (I1033148,I1033338,I1033403);
not I_60641 (I1033434,I567138);
nor I_60642 (I1033451,I1033434,I567147);
nor I_60643 (I1033468,I1033451,I567141);
nor I_60644 (I1033485,I1033236,I1033468);
DFFARX1 I_60645 (I1033485,I2507,I1033171,I1033157,);
not I_60646 (I1033516,I1033451);
DFFARX1 I_60647 (I1033516,I2507,I1033171,I1033160,);
and I_60648 (I1033154,I1033262,I1033451);
nor I_60649 (I1033561,I1033434,I567162);
and I_60650 (I1033578,I1033561,I567141);
or I_60651 (I1033595,I1033578,I567159);
DFFARX1 I_60652 (I1033595,I2507,I1033171,I1033621,);
nor I_60653 (I1033629,I1033621,I1033355);
DFFARX1 I_60654 (I1033629,I2507,I1033171,I1033142,);
nand I_60655 (I1033660,I1033621,I1033262);
nand I_60656 (I1033677,I1033355,I1033660);
nor I_60657 (I1033151,I1033677,I1033321);
not I_60658 (I1033732,I2514);
DFFARX1 I_60659 (I789609,I2507,I1033732,I1033758,);
DFFARX1 I_60660 (I1033758,I2507,I1033732,I1033775,);
not I_60661 (I1033724,I1033775);
not I_60662 (I1033797,I1033758);
DFFARX1 I_60663 (I789606,I2507,I1033732,I1033823,);
nand I_60664 (I1033831,I1033823,I789621);
not I_60665 (I1033848,I789621);
not I_60666 (I1033865,I789618);
nand I_60667 (I1033882,I789615,I789603);
and I_60668 (I1033899,I789615,I789603);
not I_60669 (I1033916,I789600);
nand I_60670 (I1033933,I1033916,I1033865);
nor I_60671 (I1033706,I1033933,I1033831);
nor I_60672 (I1033964,I1033848,I1033933);
nand I_60673 (I1033709,I1033899,I1033964);
not I_60674 (I1033995,I789606);
nor I_60675 (I1034012,I1033995,I789615);
nor I_60676 (I1034029,I1034012,I789600);
nor I_60677 (I1034046,I1033797,I1034029);
DFFARX1 I_60678 (I1034046,I2507,I1033732,I1033718,);
not I_60679 (I1034077,I1034012);
DFFARX1 I_60680 (I1034077,I2507,I1033732,I1033721,);
and I_60681 (I1033715,I1033823,I1034012);
nor I_60682 (I1034122,I1033995,I789612);
and I_60683 (I1034139,I1034122,I789600);
or I_60684 (I1034156,I1034139,I789603);
DFFARX1 I_60685 (I1034156,I2507,I1033732,I1034182,);
nor I_60686 (I1034190,I1034182,I1033916);
DFFARX1 I_60687 (I1034190,I2507,I1033732,I1033703,);
nand I_60688 (I1034221,I1034182,I1033823);
nand I_60689 (I1034238,I1033916,I1034221);
nor I_60690 (I1033712,I1034238,I1033882);
not I_60691 (I1034293,I2514);
DFFARX1 I_60692 (I246623,I2507,I1034293,I1034319,);
DFFARX1 I_60693 (I1034319,I2507,I1034293,I1034336,);
not I_60694 (I1034285,I1034336);
not I_60695 (I1034358,I1034319);
DFFARX1 I_60696 (I246638,I2507,I1034293,I1034384,);
nand I_60697 (I1034392,I1034384,I246620);
not I_60698 (I1034409,I246620);
not I_60699 (I1034426,I246629);
nand I_60700 (I1034443,I246635,I246626);
and I_60701 (I1034460,I246635,I246626);
not I_60702 (I1034477,I246623);
nand I_60703 (I1034494,I1034477,I1034426);
nor I_60704 (I1034267,I1034494,I1034392);
nor I_60705 (I1034525,I1034409,I1034494);
nand I_60706 (I1034270,I1034460,I1034525);
not I_60707 (I1034556,I246620);
nor I_60708 (I1034573,I1034556,I246635);
nor I_60709 (I1034590,I1034573,I246623);
nor I_60710 (I1034607,I1034358,I1034590);
DFFARX1 I_60711 (I1034607,I2507,I1034293,I1034279,);
not I_60712 (I1034638,I1034573);
DFFARX1 I_60713 (I1034638,I2507,I1034293,I1034282,);
and I_60714 (I1034276,I1034384,I1034573);
nor I_60715 (I1034683,I1034556,I246644);
and I_60716 (I1034700,I1034683,I246641);
or I_60717 (I1034717,I1034700,I246632);
DFFARX1 I_60718 (I1034717,I2507,I1034293,I1034743,);
nor I_60719 (I1034751,I1034743,I1034477);
DFFARX1 I_60720 (I1034751,I2507,I1034293,I1034264,);
nand I_60721 (I1034782,I1034743,I1034384);
nand I_60722 (I1034799,I1034477,I1034782);
nor I_60723 (I1034273,I1034799,I1034443);
not I_60724 (I1034854,I2514);
DFFARX1 I_60725 (I19042,I2507,I1034854,I1034880,);
DFFARX1 I_60726 (I1034880,I2507,I1034854,I1034897,);
not I_60727 (I1034846,I1034897);
not I_60728 (I1034919,I1034880);
DFFARX1 I_60729 (I19027,I2507,I1034854,I1034945,);
nand I_60730 (I1034953,I1034945,I19039);
not I_60731 (I1034970,I19039);
not I_60732 (I1034987,I19045);
nand I_60733 (I1035004,I19033,I19024);
and I_60734 (I1035021,I19033,I19024);
not I_60735 (I1035038,I19030);
nand I_60736 (I1035055,I1035038,I1034987);
nor I_60737 (I1034828,I1035055,I1034953);
nor I_60738 (I1035086,I1034970,I1035055);
nand I_60739 (I1034831,I1035021,I1035086);
not I_60740 (I1035117,I19036);
nor I_60741 (I1035134,I1035117,I19033);
nor I_60742 (I1035151,I1035134,I19030);
nor I_60743 (I1035168,I1034919,I1035151);
DFFARX1 I_60744 (I1035168,I2507,I1034854,I1034840,);
not I_60745 (I1035199,I1035134);
DFFARX1 I_60746 (I1035199,I2507,I1034854,I1034843,);
and I_60747 (I1034837,I1034945,I1035134);
nor I_60748 (I1035244,I1035117,I19024);
and I_60749 (I1035261,I1035244,I19048);
or I_60750 (I1035278,I1035261,I19027);
DFFARX1 I_60751 (I1035278,I2507,I1034854,I1035304,);
nor I_60752 (I1035312,I1035304,I1035038);
DFFARX1 I_60753 (I1035312,I2507,I1034854,I1034825,);
nand I_60754 (I1035343,I1035304,I1034945);
nand I_60755 (I1035360,I1035038,I1035343);
nor I_60756 (I1034834,I1035360,I1035004);
not I_60757 (I1035415,I2514);
DFFARX1 I_60758 (I805946,I2507,I1035415,I1035441,);
DFFARX1 I_60759 (I1035441,I2507,I1035415,I1035458,);
not I_60760 (I1035407,I1035458);
not I_60761 (I1035480,I1035441);
DFFARX1 I_60762 (I805943,I2507,I1035415,I1035506,);
nand I_60763 (I1035514,I1035506,I805958);
not I_60764 (I1035531,I805958);
not I_60765 (I1035548,I805955);
nand I_60766 (I1035565,I805952,I805940);
and I_60767 (I1035582,I805952,I805940);
not I_60768 (I1035599,I805937);
nand I_60769 (I1035616,I1035599,I1035548);
nor I_60770 (I1035389,I1035616,I1035514);
nor I_60771 (I1035647,I1035531,I1035616);
nand I_60772 (I1035392,I1035582,I1035647);
not I_60773 (I1035678,I805943);
nor I_60774 (I1035695,I1035678,I805952);
nor I_60775 (I1035712,I1035695,I805937);
nor I_60776 (I1035729,I1035480,I1035712);
DFFARX1 I_60777 (I1035729,I2507,I1035415,I1035401,);
not I_60778 (I1035760,I1035695);
DFFARX1 I_60779 (I1035760,I2507,I1035415,I1035404,);
and I_60780 (I1035398,I1035506,I1035695);
nor I_60781 (I1035805,I1035678,I805949);
and I_60782 (I1035822,I1035805,I805937);
or I_60783 (I1035839,I1035822,I805940);
DFFARX1 I_60784 (I1035839,I2507,I1035415,I1035865,);
nor I_60785 (I1035873,I1035865,I1035599);
DFFARX1 I_60786 (I1035873,I2507,I1035415,I1035386,);
nand I_60787 (I1035904,I1035865,I1035506);
nand I_60788 (I1035921,I1035599,I1035904);
nor I_60789 (I1035395,I1035921,I1035565);
not I_60790 (I1035976,I2514);
DFFARX1 I_60791 (I457223,I2507,I1035976,I1036002,);
DFFARX1 I_60792 (I1036002,I2507,I1035976,I1036019,);
not I_60793 (I1035968,I1036019);
not I_60794 (I1036041,I1036002);
DFFARX1 I_60795 (I457211,I2507,I1035976,I1036067,);
nand I_60796 (I1036075,I1036067,I457217);
not I_60797 (I1036092,I457217);
not I_60798 (I1036109,I457214);
nand I_60799 (I1036126,I457202,I457199);
and I_60800 (I1036143,I457202,I457199);
not I_60801 (I1036160,I457226);
nand I_60802 (I1036177,I1036160,I1036109);
nor I_60803 (I1035950,I1036177,I1036075);
nor I_60804 (I1036208,I1036092,I1036177);
nand I_60805 (I1035953,I1036143,I1036208);
not I_60806 (I1036239,I457199);
nor I_60807 (I1036256,I1036239,I457202);
nor I_60808 (I1036273,I1036256,I457226);
nor I_60809 (I1036290,I1036041,I1036273);
DFFARX1 I_60810 (I1036290,I2507,I1035976,I1035962,);
not I_60811 (I1036321,I1036256);
DFFARX1 I_60812 (I1036321,I2507,I1035976,I1035965,);
and I_60813 (I1035959,I1036067,I1036256);
nor I_60814 (I1036366,I1036239,I457208);
and I_60815 (I1036383,I1036366,I457205);
or I_60816 (I1036400,I1036383,I457220);
DFFARX1 I_60817 (I1036400,I2507,I1035976,I1036426,);
nor I_60818 (I1036434,I1036426,I1036160);
DFFARX1 I_60819 (I1036434,I2507,I1035976,I1035947,);
nand I_60820 (I1036465,I1036426,I1036067);
nand I_60821 (I1036482,I1036160,I1036465);
nor I_60822 (I1035956,I1036482,I1036126);
not I_60823 (I1036537,I2514);
DFFARX1 I_60824 (I218063,I2507,I1036537,I1036563,);
DFFARX1 I_60825 (I1036563,I2507,I1036537,I1036580,);
not I_60826 (I1036529,I1036580);
not I_60827 (I1036602,I1036563);
DFFARX1 I_60828 (I218078,I2507,I1036537,I1036628,);
nand I_60829 (I1036636,I1036628,I218060);
not I_60830 (I1036653,I218060);
not I_60831 (I1036670,I218069);
nand I_60832 (I1036687,I218075,I218066);
and I_60833 (I1036704,I218075,I218066);
not I_60834 (I1036721,I218063);
nand I_60835 (I1036738,I1036721,I1036670);
nor I_60836 (I1036511,I1036738,I1036636);
nor I_60837 (I1036769,I1036653,I1036738);
nand I_60838 (I1036514,I1036704,I1036769);
not I_60839 (I1036800,I218060);
nor I_60840 (I1036817,I1036800,I218075);
nor I_60841 (I1036834,I1036817,I218063);
nor I_60842 (I1036851,I1036602,I1036834);
DFFARX1 I_60843 (I1036851,I2507,I1036537,I1036523,);
not I_60844 (I1036882,I1036817);
DFFARX1 I_60845 (I1036882,I2507,I1036537,I1036526,);
and I_60846 (I1036520,I1036628,I1036817);
nor I_60847 (I1036927,I1036800,I218084);
and I_60848 (I1036944,I1036927,I218081);
or I_60849 (I1036961,I1036944,I218072);
DFFARX1 I_60850 (I1036961,I2507,I1036537,I1036987,);
nor I_60851 (I1036995,I1036987,I1036721);
DFFARX1 I_60852 (I1036995,I2507,I1036537,I1036508,);
nand I_60853 (I1037026,I1036987,I1036628);
nand I_60854 (I1037043,I1036721,I1037026);
nor I_60855 (I1036517,I1037043,I1036687);
not I_60856 (I1037098,I2514);
DFFARX1 I_60857 (I1195949,I2507,I1037098,I1037124,);
DFFARX1 I_60858 (I1037124,I2507,I1037098,I1037141,);
not I_60859 (I1037090,I1037141);
not I_60860 (I1037163,I1037124);
DFFARX1 I_60861 (I1195940,I2507,I1037098,I1037189,);
nand I_60862 (I1037197,I1037189,I1195937);
not I_60863 (I1037214,I1195937);
not I_60864 (I1037231,I1195946);
nand I_60865 (I1037248,I1195955,I1195937);
and I_60866 (I1037265,I1195955,I1195937);
not I_60867 (I1037282,I1195934);
nand I_60868 (I1037299,I1037282,I1037231);
nor I_60869 (I1037072,I1037299,I1037197);
nor I_60870 (I1037330,I1037214,I1037299);
nand I_60871 (I1037075,I1037265,I1037330);
not I_60872 (I1037361,I1195943);
nor I_60873 (I1037378,I1037361,I1195955);
nor I_60874 (I1037395,I1037378,I1195934);
nor I_60875 (I1037412,I1037163,I1037395);
DFFARX1 I_60876 (I1037412,I2507,I1037098,I1037084,);
not I_60877 (I1037443,I1037378);
DFFARX1 I_60878 (I1037443,I2507,I1037098,I1037087,);
and I_60879 (I1037081,I1037189,I1037378);
nor I_60880 (I1037488,I1037361,I1195958);
and I_60881 (I1037505,I1037488,I1195934);
or I_60882 (I1037522,I1037505,I1195952);
DFFARX1 I_60883 (I1037522,I2507,I1037098,I1037548,);
nor I_60884 (I1037556,I1037548,I1037282);
DFFARX1 I_60885 (I1037556,I2507,I1037098,I1037069,);
nand I_60886 (I1037587,I1037548,I1037189);
nand I_60887 (I1037604,I1037282,I1037587);
nor I_60888 (I1037078,I1037604,I1037248);
not I_60889 (I1037659,I2514);
DFFARX1 I_60890 (I1197683,I2507,I1037659,I1037685,);
DFFARX1 I_60891 (I1037685,I2507,I1037659,I1037702,);
not I_60892 (I1037651,I1037702);
not I_60893 (I1037724,I1037685);
DFFARX1 I_60894 (I1197674,I2507,I1037659,I1037750,);
nand I_60895 (I1037758,I1037750,I1197671);
not I_60896 (I1037775,I1197671);
not I_60897 (I1037792,I1197680);
nand I_60898 (I1037809,I1197689,I1197671);
and I_60899 (I1037826,I1197689,I1197671);
not I_60900 (I1037843,I1197668);
nand I_60901 (I1037860,I1037843,I1037792);
nor I_60902 (I1037633,I1037860,I1037758);
nor I_60903 (I1037891,I1037775,I1037860);
nand I_60904 (I1037636,I1037826,I1037891);
not I_60905 (I1037922,I1197677);
nor I_60906 (I1037939,I1037922,I1197689);
nor I_60907 (I1037956,I1037939,I1197668);
nor I_60908 (I1037973,I1037724,I1037956);
DFFARX1 I_60909 (I1037973,I2507,I1037659,I1037645,);
not I_60910 (I1038004,I1037939);
DFFARX1 I_60911 (I1038004,I2507,I1037659,I1037648,);
and I_60912 (I1037642,I1037750,I1037939);
nor I_60913 (I1038049,I1037922,I1197692);
and I_60914 (I1038066,I1038049,I1197668);
or I_60915 (I1038083,I1038066,I1197686);
DFFARX1 I_60916 (I1038083,I2507,I1037659,I1038109,);
nor I_60917 (I1038117,I1038109,I1037843);
DFFARX1 I_60918 (I1038117,I2507,I1037659,I1037630,);
nand I_60919 (I1038148,I1038109,I1037750);
nand I_60920 (I1038165,I1037843,I1038148);
nor I_60921 (I1037639,I1038165,I1037809);
not I_60922 (I1038220,I2514);
DFFARX1 I_60923 (I290263,I2507,I1038220,I1038246,);
DFFARX1 I_60924 (I1038246,I2507,I1038220,I1038263,);
not I_60925 (I1038212,I1038263);
not I_60926 (I1038285,I1038246);
DFFARX1 I_60927 (I290260,I2507,I1038220,I1038311,);
nand I_60928 (I1038319,I1038311,I290254);
not I_60929 (I1038336,I290254);
not I_60930 (I1038353,I290251);
nand I_60931 (I1038370,I290245,I290242);
and I_60932 (I1038387,I290245,I290242);
not I_60933 (I1038404,I290257);
nand I_60934 (I1038421,I1038404,I1038353);
nor I_60935 (I1038194,I1038421,I1038319);
nor I_60936 (I1038452,I1038336,I1038421);
nand I_60937 (I1038197,I1038387,I1038452);
not I_60938 (I1038483,I290269);
nor I_60939 (I1038500,I1038483,I290245);
nor I_60940 (I1038517,I1038500,I290257);
nor I_60941 (I1038534,I1038285,I1038517);
DFFARX1 I_60942 (I1038534,I2507,I1038220,I1038206,);
not I_60943 (I1038565,I1038500);
DFFARX1 I_60944 (I1038565,I2507,I1038220,I1038209,);
and I_60945 (I1038203,I1038311,I1038500);
nor I_60946 (I1038610,I1038483,I290266);
and I_60947 (I1038627,I1038610,I290242);
or I_60948 (I1038644,I1038627,I290248);
DFFARX1 I_60949 (I1038644,I2507,I1038220,I1038670,);
nor I_60950 (I1038678,I1038670,I1038404);
DFFARX1 I_60951 (I1038678,I2507,I1038220,I1038191,);
nand I_60952 (I1038709,I1038670,I1038311);
nand I_60953 (I1038726,I1038404,I1038709);
nor I_60954 (I1038200,I1038726,I1038370);
not I_60955 (I1038781,I2514);
DFFARX1 I_60956 (I497082,I2507,I1038781,I1038807,);
DFFARX1 I_60957 (I1038807,I2507,I1038781,I1038824,);
not I_60958 (I1038773,I1038824);
not I_60959 (I1038846,I1038807);
DFFARX1 I_60960 (I497079,I2507,I1038781,I1038872,);
nand I_60961 (I1038880,I1038872,I497073);
not I_60962 (I1038897,I497073);
not I_60963 (I1038914,I497085);
nand I_60964 (I1038931,I497088,I497067);
and I_60965 (I1038948,I497088,I497067);
not I_60966 (I1038965,I497064);
nand I_60967 (I1038982,I1038965,I1038914);
nor I_60968 (I1038755,I1038982,I1038880);
nor I_60969 (I1039013,I1038897,I1038982);
nand I_60970 (I1038758,I1038948,I1039013);
not I_60971 (I1039044,I497070);
nor I_60972 (I1039061,I1039044,I497088);
nor I_60973 (I1039078,I1039061,I497064);
nor I_60974 (I1039095,I1038846,I1039078);
DFFARX1 I_60975 (I1039095,I2507,I1038781,I1038767,);
not I_60976 (I1039126,I1039061);
DFFARX1 I_60977 (I1039126,I2507,I1038781,I1038770,);
and I_60978 (I1038764,I1038872,I1039061);
nor I_60979 (I1039171,I1039044,I497064);
and I_60980 (I1039188,I1039171,I497076);
or I_60981 (I1039205,I1039188,I497067);
DFFARX1 I_60982 (I1039205,I2507,I1038781,I1039231,);
nor I_60983 (I1039239,I1039231,I1038965);
DFFARX1 I_60984 (I1039239,I2507,I1038781,I1038752,);
nand I_60985 (I1039270,I1039231,I1038872);
nand I_60986 (I1039287,I1038965,I1039270);
nor I_60987 (I1038761,I1039287,I1038931);
not I_60988 (I1039342,I2514);
DFFARX1 I_60989 (I47500,I2507,I1039342,I1039368,);
DFFARX1 I_60990 (I1039368,I2507,I1039342,I1039385,);
not I_60991 (I1039334,I1039385);
not I_60992 (I1039407,I1039368);
DFFARX1 I_60993 (I47485,I2507,I1039342,I1039433,);
nand I_60994 (I1039441,I1039433,I47497);
not I_60995 (I1039458,I47497);
not I_60996 (I1039475,I47503);
nand I_60997 (I1039492,I47491,I47482);
and I_60998 (I1039509,I47491,I47482);
not I_60999 (I1039526,I47488);
nand I_61000 (I1039543,I1039526,I1039475);
nor I_61001 (I1039316,I1039543,I1039441);
nor I_61002 (I1039574,I1039458,I1039543);
nand I_61003 (I1039319,I1039509,I1039574);
not I_61004 (I1039605,I47494);
nor I_61005 (I1039622,I1039605,I47491);
nor I_61006 (I1039639,I1039622,I47488);
nor I_61007 (I1039656,I1039407,I1039639);
DFFARX1 I_61008 (I1039656,I2507,I1039342,I1039328,);
not I_61009 (I1039687,I1039622);
DFFARX1 I_61010 (I1039687,I2507,I1039342,I1039331,);
and I_61011 (I1039325,I1039433,I1039622);
nor I_61012 (I1039732,I1039605,I47482);
and I_61013 (I1039749,I1039732,I47506);
or I_61014 (I1039766,I1039749,I47485);
DFFARX1 I_61015 (I1039766,I2507,I1039342,I1039792,);
nor I_61016 (I1039800,I1039792,I1039526);
DFFARX1 I_61017 (I1039800,I2507,I1039342,I1039313,);
nand I_61018 (I1039831,I1039792,I1039433);
nand I_61019 (I1039848,I1039526,I1039831);
nor I_61020 (I1039322,I1039848,I1039492);
not I_61021 (I1039903,I2514);
DFFARX1 I_61022 (I737651,I2507,I1039903,I1039929,);
DFFARX1 I_61023 (I1039929,I2507,I1039903,I1039946,);
not I_61024 (I1039895,I1039946);
not I_61025 (I1039968,I1039929);
DFFARX1 I_61026 (I737663,I2507,I1039903,I1039994,);
nand I_61027 (I1040002,I1039994,I737672);
not I_61028 (I1040019,I737672);
not I_61029 (I1040036,I737654);
nand I_61030 (I1040053,I737657,I737648);
and I_61031 (I1040070,I737657,I737648);
not I_61032 (I1040087,I737666);
nand I_61033 (I1040104,I1040087,I1040036);
nor I_61034 (I1039877,I1040104,I1040002);
nor I_61035 (I1040135,I1040019,I1040104);
nand I_61036 (I1039880,I1040070,I1040135);
not I_61037 (I1040166,I737669);
nor I_61038 (I1040183,I1040166,I737657);
nor I_61039 (I1040200,I1040183,I737666);
nor I_61040 (I1040217,I1039968,I1040200);
DFFARX1 I_61041 (I1040217,I2507,I1039903,I1039889,);
not I_61042 (I1040248,I1040183);
DFFARX1 I_61043 (I1040248,I2507,I1039903,I1039892,);
and I_61044 (I1039886,I1039994,I1040183);
nor I_61045 (I1040293,I1040166,I737648);
and I_61046 (I1040310,I1040293,I737660);
or I_61047 (I1040327,I1040310,I737651);
DFFARX1 I_61048 (I1040327,I2507,I1039903,I1040353,);
nor I_61049 (I1040361,I1040353,I1040087);
DFFARX1 I_61050 (I1040361,I2507,I1039903,I1039874,);
nand I_61051 (I1040392,I1040353,I1039994);
nand I_61052 (I1040409,I1040087,I1040392);
nor I_61053 (I1039883,I1040409,I1040053);
not I_61054 (I1040464,I2514);
DFFARX1 I_61055 (I270764,I2507,I1040464,I1040490,);
DFFARX1 I_61056 (I1040490,I2507,I1040464,I1040507,);
not I_61057 (I1040456,I1040507);
not I_61058 (I1040529,I1040490);
DFFARX1 I_61059 (I270761,I2507,I1040464,I1040555,);
nand I_61060 (I1040563,I1040555,I270755);
not I_61061 (I1040580,I270755);
not I_61062 (I1040597,I270752);
nand I_61063 (I1040614,I270746,I270743);
and I_61064 (I1040631,I270746,I270743);
not I_61065 (I1040648,I270758);
nand I_61066 (I1040665,I1040648,I1040597);
nor I_61067 (I1040438,I1040665,I1040563);
nor I_61068 (I1040696,I1040580,I1040665);
nand I_61069 (I1040441,I1040631,I1040696);
not I_61070 (I1040727,I270770);
nor I_61071 (I1040744,I1040727,I270746);
nor I_61072 (I1040761,I1040744,I270758);
nor I_61073 (I1040778,I1040529,I1040761);
DFFARX1 I_61074 (I1040778,I2507,I1040464,I1040450,);
not I_61075 (I1040809,I1040744);
DFFARX1 I_61076 (I1040809,I2507,I1040464,I1040453,);
and I_61077 (I1040447,I1040555,I1040744);
nor I_61078 (I1040854,I1040727,I270767);
and I_61079 (I1040871,I1040854,I270743);
or I_61080 (I1040888,I1040871,I270749);
DFFARX1 I_61081 (I1040888,I2507,I1040464,I1040914,);
nor I_61082 (I1040922,I1040914,I1040648);
DFFARX1 I_61083 (I1040922,I2507,I1040464,I1040435,);
nand I_61084 (I1040953,I1040914,I1040555);
nand I_61085 (I1040970,I1040648,I1040953);
nor I_61086 (I1040444,I1040970,I1040614);
not I_61087 (I1041025,I2514);
DFFARX1 I_61088 (I727247,I2507,I1041025,I1041051,);
DFFARX1 I_61089 (I1041051,I2507,I1041025,I1041068,);
not I_61090 (I1041017,I1041068);
not I_61091 (I1041090,I1041051);
DFFARX1 I_61092 (I727259,I2507,I1041025,I1041116,);
nand I_61093 (I1041124,I1041116,I727268);
not I_61094 (I1041141,I727268);
not I_61095 (I1041158,I727250);
nand I_61096 (I1041175,I727253,I727244);
and I_61097 (I1041192,I727253,I727244);
not I_61098 (I1041209,I727262);
nand I_61099 (I1041226,I1041209,I1041158);
nor I_61100 (I1040999,I1041226,I1041124);
nor I_61101 (I1041257,I1041141,I1041226);
nand I_61102 (I1041002,I1041192,I1041257);
not I_61103 (I1041288,I727265);
nor I_61104 (I1041305,I1041288,I727253);
nor I_61105 (I1041322,I1041305,I727262);
nor I_61106 (I1041339,I1041090,I1041322);
DFFARX1 I_61107 (I1041339,I2507,I1041025,I1041011,);
not I_61108 (I1041370,I1041305);
DFFARX1 I_61109 (I1041370,I2507,I1041025,I1041014,);
and I_61110 (I1041008,I1041116,I1041305);
nor I_61111 (I1041415,I1041288,I727244);
and I_61112 (I1041432,I1041415,I727256);
or I_61113 (I1041449,I1041432,I727247);
DFFARX1 I_61114 (I1041449,I2507,I1041025,I1041475,);
nor I_61115 (I1041483,I1041475,I1041209);
DFFARX1 I_61116 (I1041483,I2507,I1041025,I1040996,);
nand I_61117 (I1041514,I1041475,I1041116);
nand I_61118 (I1041531,I1041209,I1041514);
nor I_61119 (I1041005,I1041531,I1041175);
not I_61120 (I1041586,I2514);
DFFARX1 I_61121 (I1180343,I2507,I1041586,I1041612,);
DFFARX1 I_61122 (I1041612,I2507,I1041586,I1041629,);
not I_61123 (I1041578,I1041629);
not I_61124 (I1041651,I1041612);
DFFARX1 I_61125 (I1180334,I2507,I1041586,I1041677,);
nand I_61126 (I1041685,I1041677,I1180331);
not I_61127 (I1041702,I1180331);
not I_61128 (I1041719,I1180340);
nand I_61129 (I1041736,I1180349,I1180331);
and I_61130 (I1041753,I1180349,I1180331);
not I_61131 (I1041770,I1180328);
nand I_61132 (I1041787,I1041770,I1041719);
nor I_61133 (I1041560,I1041787,I1041685);
nor I_61134 (I1041818,I1041702,I1041787);
nand I_61135 (I1041563,I1041753,I1041818);
not I_61136 (I1041849,I1180337);
nor I_61137 (I1041866,I1041849,I1180349);
nor I_61138 (I1041883,I1041866,I1180328);
nor I_61139 (I1041900,I1041651,I1041883);
DFFARX1 I_61140 (I1041900,I2507,I1041586,I1041572,);
not I_61141 (I1041931,I1041866);
DFFARX1 I_61142 (I1041931,I2507,I1041586,I1041575,);
and I_61143 (I1041569,I1041677,I1041866);
nor I_61144 (I1041976,I1041849,I1180352);
and I_61145 (I1041993,I1041976,I1180328);
or I_61146 (I1042010,I1041993,I1180346);
DFFARX1 I_61147 (I1042010,I2507,I1041586,I1042036,);
nor I_61148 (I1042044,I1042036,I1041770);
DFFARX1 I_61149 (I1042044,I2507,I1041586,I1041557,);
nand I_61150 (I1042075,I1042036,I1041677);
nand I_61151 (I1042092,I1041770,I1042075);
nor I_61152 (I1041566,I1042092,I1041736);
not I_61153 (I1042147,I2514);
DFFARX1 I_61154 (I837566,I2507,I1042147,I1042173,);
DFFARX1 I_61155 (I1042173,I2507,I1042147,I1042190,);
not I_61156 (I1042139,I1042190);
not I_61157 (I1042212,I1042173);
DFFARX1 I_61158 (I837563,I2507,I1042147,I1042238,);
nand I_61159 (I1042246,I1042238,I837578);
not I_61160 (I1042263,I837578);
not I_61161 (I1042280,I837575);
nand I_61162 (I1042297,I837572,I837560);
and I_61163 (I1042314,I837572,I837560);
not I_61164 (I1042331,I837557);
nand I_61165 (I1042348,I1042331,I1042280);
nor I_61166 (I1042121,I1042348,I1042246);
nor I_61167 (I1042379,I1042263,I1042348);
nand I_61168 (I1042124,I1042314,I1042379);
not I_61169 (I1042410,I837563);
nor I_61170 (I1042427,I1042410,I837572);
nor I_61171 (I1042444,I1042427,I837557);
nor I_61172 (I1042461,I1042212,I1042444);
DFFARX1 I_61173 (I1042461,I2507,I1042147,I1042133,);
not I_61174 (I1042492,I1042427);
DFFARX1 I_61175 (I1042492,I2507,I1042147,I1042136,);
and I_61176 (I1042130,I1042238,I1042427);
nor I_61177 (I1042537,I1042410,I837569);
and I_61178 (I1042554,I1042537,I837557);
or I_61179 (I1042571,I1042554,I837560);
DFFARX1 I_61180 (I1042571,I2507,I1042147,I1042597,);
nor I_61181 (I1042605,I1042597,I1042331);
DFFARX1 I_61182 (I1042605,I2507,I1042147,I1042118,);
nand I_61183 (I1042636,I1042597,I1042238);
nand I_61184 (I1042653,I1042331,I1042636);
nor I_61185 (I1042127,I1042653,I1042297);
not I_61186 (I1042708,I2514);
DFFARX1 I_61187 (I827026,I2507,I1042708,I1042734,);
DFFARX1 I_61188 (I1042734,I2507,I1042708,I1042751,);
not I_61189 (I1042700,I1042751);
not I_61190 (I1042773,I1042734);
DFFARX1 I_61191 (I827023,I2507,I1042708,I1042799,);
nand I_61192 (I1042807,I1042799,I827038);
not I_61193 (I1042824,I827038);
not I_61194 (I1042841,I827035);
nand I_61195 (I1042858,I827032,I827020);
and I_61196 (I1042875,I827032,I827020);
not I_61197 (I1042892,I827017);
nand I_61198 (I1042909,I1042892,I1042841);
nor I_61199 (I1042682,I1042909,I1042807);
nor I_61200 (I1042940,I1042824,I1042909);
nand I_61201 (I1042685,I1042875,I1042940);
not I_61202 (I1042971,I827023);
nor I_61203 (I1042988,I1042971,I827032);
nor I_61204 (I1043005,I1042988,I827017);
nor I_61205 (I1043022,I1042773,I1043005);
DFFARX1 I_61206 (I1043022,I2507,I1042708,I1042694,);
not I_61207 (I1043053,I1042988);
DFFARX1 I_61208 (I1043053,I2507,I1042708,I1042697,);
and I_61209 (I1042691,I1042799,I1042988);
nor I_61210 (I1043098,I1042971,I827029);
and I_61211 (I1043115,I1043098,I827017);
or I_61212 (I1043132,I1043115,I827020);
DFFARX1 I_61213 (I1043132,I2507,I1042708,I1043158,);
nor I_61214 (I1043166,I1043158,I1042892);
DFFARX1 I_61215 (I1043166,I2507,I1042708,I1042679,);
nand I_61216 (I1043197,I1043158,I1042799);
nand I_61217 (I1043214,I1042892,I1043197);
nor I_61218 (I1042688,I1043214,I1042858);
not I_61219 (I1043269,I2514);
DFFARX1 I_61220 (I1248232,I2507,I1043269,I1043295,);
DFFARX1 I_61221 (I1043295,I2507,I1043269,I1043312,);
not I_61222 (I1043261,I1043312);
not I_61223 (I1043334,I1043295);
DFFARX1 I_61224 (I1248238,I2507,I1043269,I1043360,);
nand I_61225 (I1043368,I1043360,I1248247);
not I_61226 (I1043385,I1248247);
not I_61227 (I1043402,I1248226);
nand I_61228 (I1043419,I1248229,I1248229);
and I_61229 (I1043436,I1248229,I1248229);
not I_61230 (I1043453,I1248241);
nand I_61231 (I1043470,I1043453,I1043402);
nor I_61232 (I1043243,I1043470,I1043368);
nor I_61233 (I1043501,I1043385,I1043470);
nand I_61234 (I1043246,I1043436,I1043501);
not I_61235 (I1043532,I1248235);
nor I_61236 (I1043549,I1043532,I1248229);
nor I_61237 (I1043566,I1043549,I1248241);
nor I_61238 (I1043583,I1043334,I1043566);
DFFARX1 I_61239 (I1043583,I2507,I1043269,I1043255,);
not I_61240 (I1043614,I1043549);
DFFARX1 I_61241 (I1043614,I2507,I1043269,I1043258,);
and I_61242 (I1043252,I1043360,I1043549);
nor I_61243 (I1043659,I1043532,I1248250);
and I_61244 (I1043676,I1043659,I1248226);
or I_61245 (I1043693,I1043676,I1248244);
DFFARX1 I_61246 (I1043693,I2507,I1043269,I1043719,);
nor I_61247 (I1043727,I1043719,I1043453);
DFFARX1 I_61248 (I1043727,I2507,I1043269,I1043240,);
nand I_61249 (I1043758,I1043719,I1043360);
nand I_61250 (I1043775,I1043453,I1043758);
nor I_61251 (I1043249,I1043775,I1043419);
not I_61252 (I1043830,I2514);
DFFARX1 I_61253 (I10258,I2507,I1043830,I1043856,);
DFFARX1 I_61254 (I1043856,I2507,I1043830,I1043873,);
not I_61255 (I1043822,I1043873);
not I_61256 (I1043895,I1043856);
DFFARX1 I_61257 (I10270,I2507,I1043830,I1043921,);
nand I_61258 (I1043929,I1043921,I10267);
not I_61259 (I1043946,I10267);
not I_61260 (I1043963,I10258);
nand I_61261 (I1043980,I10252,I10252);
and I_61262 (I1043997,I10252,I10252);
not I_61263 (I1044014,I10273);
nand I_61264 (I1044031,I1044014,I1043963);
nor I_61265 (I1043804,I1044031,I1043929);
nor I_61266 (I1044062,I1043946,I1044031);
nand I_61267 (I1043807,I1043997,I1044062);
not I_61268 (I1044093,I10264);
nor I_61269 (I1044110,I1044093,I10252);
nor I_61270 (I1044127,I1044110,I10273);
nor I_61271 (I1044144,I1043895,I1044127);
DFFARX1 I_61272 (I1044144,I2507,I1043830,I1043816,);
not I_61273 (I1044175,I1044110);
DFFARX1 I_61274 (I1044175,I2507,I1043830,I1043819,);
and I_61275 (I1043813,I1043921,I1044110);
nor I_61276 (I1044220,I1044093,I10255);
and I_61277 (I1044237,I1044220,I10255);
or I_61278 (I1044254,I1044237,I10261);
DFFARX1 I_61279 (I1044254,I2507,I1043830,I1044280,);
nor I_61280 (I1044288,I1044280,I1044014);
DFFARX1 I_61281 (I1044288,I2507,I1043830,I1043801,);
nand I_61282 (I1044319,I1044280,I1043921);
nand I_61283 (I1044336,I1044014,I1044319);
nor I_61284 (I1043810,I1044336,I1043980);
not I_61285 (I1044391,I2514);
DFFARX1 I_61286 (I661933,I2507,I1044391,I1044417,);
DFFARX1 I_61287 (I1044417,I2507,I1044391,I1044434,);
not I_61288 (I1044383,I1044434);
not I_61289 (I1044456,I1044417);
DFFARX1 I_61290 (I661945,I2507,I1044391,I1044482,);
nand I_61291 (I1044490,I1044482,I661954);
not I_61292 (I1044507,I661954);
not I_61293 (I1044524,I661936);
nand I_61294 (I1044541,I661939,I661930);
and I_61295 (I1044558,I661939,I661930);
not I_61296 (I1044575,I661948);
nand I_61297 (I1044592,I1044575,I1044524);
nor I_61298 (I1044365,I1044592,I1044490);
nor I_61299 (I1044623,I1044507,I1044592);
nand I_61300 (I1044368,I1044558,I1044623);
not I_61301 (I1044654,I661951);
nor I_61302 (I1044671,I1044654,I661939);
nor I_61303 (I1044688,I1044671,I661948);
nor I_61304 (I1044705,I1044456,I1044688);
DFFARX1 I_61305 (I1044705,I2507,I1044391,I1044377,);
not I_61306 (I1044736,I1044671);
DFFARX1 I_61307 (I1044736,I2507,I1044391,I1044380,);
and I_61308 (I1044374,I1044482,I1044671);
nor I_61309 (I1044781,I1044654,I661930);
and I_61310 (I1044798,I1044781,I661942);
or I_61311 (I1044815,I1044798,I661933);
DFFARX1 I_61312 (I1044815,I2507,I1044391,I1044841,);
nor I_61313 (I1044849,I1044841,I1044575);
DFFARX1 I_61314 (I1044849,I2507,I1044391,I1044362,);
nand I_61315 (I1044880,I1044841,I1044482);
nand I_61316 (I1044897,I1044575,I1044880);
nor I_61317 (I1044371,I1044897,I1044541);
not I_61318 (I1044952,I2514);
DFFARX1 I_61319 (I974781,I2507,I1044952,I1044978,);
DFFARX1 I_61320 (I1044978,I2507,I1044952,I1044995,);
not I_61321 (I1044944,I1044995);
not I_61322 (I1045017,I1044978);
DFFARX1 I_61323 (I974808,I2507,I1044952,I1045043,);
nand I_61324 (I1045051,I1045043,I974799);
not I_61325 (I1045068,I974799);
not I_61326 (I1045085,I974781);
nand I_61327 (I1045102,I974793,I974796);
and I_61328 (I1045119,I974793,I974796);
not I_61329 (I1045136,I974805);
nand I_61330 (I1045153,I1045136,I1045085);
nor I_61331 (I1044926,I1045153,I1045051);
nor I_61332 (I1045184,I1045068,I1045153);
nand I_61333 (I1044929,I1045119,I1045184);
not I_61334 (I1045215,I974790);
nor I_61335 (I1045232,I1045215,I974793);
nor I_61336 (I1045249,I1045232,I974805);
nor I_61337 (I1045266,I1045017,I1045249);
DFFARX1 I_61338 (I1045266,I2507,I1044952,I1044938,);
not I_61339 (I1045297,I1045232);
DFFARX1 I_61340 (I1045297,I2507,I1044952,I1044941,);
and I_61341 (I1044935,I1045043,I1045232);
nor I_61342 (I1045342,I1045215,I974784);
and I_61343 (I1045359,I1045342,I974787);
or I_61344 (I1045376,I1045359,I974802);
DFFARX1 I_61345 (I1045376,I2507,I1044952,I1045402,);
nor I_61346 (I1045410,I1045402,I1045136);
DFFARX1 I_61347 (I1045410,I2507,I1044952,I1044923,);
nand I_61348 (I1045441,I1045402,I1045043);
nand I_61349 (I1045458,I1045136,I1045441);
nor I_61350 (I1044932,I1045458,I1045102);
not I_61351 (I1045513,I2514);
DFFARX1 I_61352 (I114423,I2507,I1045513,I1045539,);
DFFARX1 I_61353 (I1045539,I2507,I1045513,I1045556,);
not I_61354 (I1045505,I1045556);
not I_61355 (I1045578,I1045539);
DFFARX1 I_61356 (I114411,I2507,I1045513,I1045604,);
nand I_61357 (I1045612,I1045604,I114426);
not I_61358 (I1045629,I114426);
not I_61359 (I1045646,I114414);
nand I_61360 (I1045663,I114435,I114429);
and I_61361 (I1045680,I114435,I114429);
not I_61362 (I1045697,I114417);
nand I_61363 (I1045714,I1045697,I1045646);
nor I_61364 (I1045487,I1045714,I1045612);
nor I_61365 (I1045745,I1045629,I1045714);
nand I_61366 (I1045490,I1045680,I1045745);
not I_61367 (I1045776,I114420);
nor I_61368 (I1045793,I1045776,I114435);
nor I_61369 (I1045810,I1045793,I114417);
nor I_61370 (I1045827,I1045578,I1045810);
DFFARX1 I_61371 (I1045827,I2507,I1045513,I1045499,);
not I_61372 (I1045858,I1045793);
DFFARX1 I_61373 (I1045858,I2507,I1045513,I1045502,);
and I_61374 (I1045496,I1045604,I1045793);
nor I_61375 (I1045903,I1045776,I114414);
and I_61376 (I1045920,I1045903,I114411);
or I_61377 (I1045937,I1045920,I114432);
DFFARX1 I_61378 (I1045937,I2507,I1045513,I1045963,);
nor I_61379 (I1045971,I1045963,I1045697);
DFFARX1 I_61380 (I1045971,I2507,I1045513,I1045484,);
nand I_61381 (I1046002,I1045963,I1045604);
nand I_61382 (I1046019,I1045697,I1046002);
nor I_61383 (I1045493,I1046019,I1045663);
not I_61384 (I1046074,I2514);
DFFARX1 I_61385 (I1385057,I2507,I1046074,I1046100,);
DFFARX1 I_61386 (I1046100,I2507,I1046074,I1046117,);
not I_61387 (I1046066,I1046117);
not I_61388 (I1046139,I1046100);
DFFARX1 I_61389 (I1385051,I2507,I1046074,I1046165,);
nand I_61390 (I1046173,I1046165,I1385042);
not I_61391 (I1046190,I1385042);
not I_61392 (I1046207,I1385069);
nand I_61393 (I1046224,I1385054,I1385063);
and I_61394 (I1046241,I1385054,I1385063);
not I_61395 (I1046258,I1385048);
nand I_61396 (I1046275,I1046258,I1046207);
nor I_61397 (I1046048,I1046275,I1046173);
nor I_61398 (I1046306,I1046190,I1046275);
nand I_61399 (I1046051,I1046241,I1046306);
not I_61400 (I1046337,I1385066);
nor I_61401 (I1046354,I1046337,I1385054);
nor I_61402 (I1046371,I1046354,I1385048);
nor I_61403 (I1046388,I1046139,I1046371);
DFFARX1 I_61404 (I1046388,I2507,I1046074,I1046060,);
not I_61405 (I1046419,I1046354);
DFFARX1 I_61406 (I1046419,I2507,I1046074,I1046063,);
and I_61407 (I1046057,I1046165,I1046354);
nor I_61408 (I1046464,I1046337,I1385060);
and I_61409 (I1046481,I1046464,I1385042);
or I_61410 (I1046498,I1046481,I1385045);
DFFARX1 I_61411 (I1046498,I2507,I1046074,I1046524,);
nor I_61412 (I1046532,I1046524,I1046258);
DFFARX1 I_61413 (I1046532,I2507,I1046074,I1046045,);
nand I_61414 (I1046563,I1046524,I1046165);
nand I_61415 (I1046580,I1046258,I1046563);
nor I_61416 (I1046054,I1046580,I1046224);
not I_61417 (I1046635,I2514);
DFFARX1 I_61418 (I699503,I2507,I1046635,I1046661,);
DFFARX1 I_61419 (I1046661,I2507,I1046635,I1046678,);
not I_61420 (I1046627,I1046678);
not I_61421 (I1046700,I1046661);
DFFARX1 I_61422 (I699515,I2507,I1046635,I1046726,);
nand I_61423 (I1046734,I1046726,I699524);
not I_61424 (I1046751,I699524);
not I_61425 (I1046768,I699506);
nand I_61426 (I1046785,I699509,I699500);
and I_61427 (I1046802,I699509,I699500);
not I_61428 (I1046819,I699518);
nand I_61429 (I1046836,I1046819,I1046768);
nor I_61430 (I1046609,I1046836,I1046734);
nor I_61431 (I1046867,I1046751,I1046836);
nand I_61432 (I1046612,I1046802,I1046867);
not I_61433 (I1046898,I699521);
nor I_61434 (I1046915,I1046898,I699509);
nor I_61435 (I1046932,I1046915,I699518);
nor I_61436 (I1046949,I1046700,I1046932);
DFFARX1 I_61437 (I1046949,I2507,I1046635,I1046621,);
not I_61438 (I1046980,I1046915);
DFFARX1 I_61439 (I1046980,I2507,I1046635,I1046624,);
and I_61440 (I1046618,I1046726,I1046915);
nor I_61441 (I1047025,I1046898,I699500);
and I_61442 (I1047042,I1047025,I699512);
or I_61443 (I1047059,I1047042,I699503);
DFFARX1 I_61444 (I1047059,I2507,I1046635,I1047085,);
nor I_61445 (I1047093,I1047085,I1046819);
DFFARX1 I_61446 (I1047093,I2507,I1046635,I1046606,);
nand I_61447 (I1047124,I1047085,I1046726);
nand I_61448 (I1047141,I1046819,I1047124);
nor I_61449 (I1046615,I1047141,I1046785);
not I_61450 (I1047196,I2514);
DFFARX1 I_61451 (I138949,I2507,I1047196,I1047222,);
DFFARX1 I_61452 (I1047222,I2507,I1047196,I1047239,);
not I_61453 (I1047188,I1047239);
not I_61454 (I1047261,I1047222);
DFFARX1 I_61455 (I138931,I2507,I1047196,I1047287,);
nand I_61456 (I1047295,I1047287,I138925);
not I_61457 (I1047312,I138925);
not I_61458 (I1047329,I138928);
nand I_61459 (I1047346,I138943,I138934);
and I_61460 (I1047363,I138943,I138934);
not I_61461 (I1047380,I138946);
nand I_61462 (I1047397,I1047380,I1047329);
nor I_61463 (I1047170,I1047397,I1047295);
nor I_61464 (I1047428,I1047312,I1047397);
nand I_61465 (I1047173,I1047363,I1047428);
not I_61466 (I1047459,I138940);
nor I_61467 (I1047476,I1047459,I138943);
nor I_61468 (I1047493,I1047476,I138946);
nor I_61469 (I1047510,I1047261,I1047493);
DFFARX1 I_61470 (I1047510,I2507,I1047196,I1047182,);
not I_61471 (I1047541,I1047476);
DFFARX1 I_61472 (I1047541,I2507,I1047196,I1047185,);
and I_61473 (I1047179,I1047287,I1047476);
nor I_61474 (I1047586,I1047459,I138952);
and I_61475 (I1047603,I1047586,I138925);
or I_61476 (I1047620,I1047603,I138937);
DFFARX1 I_61477 (I1047620,I2507,I1047196,I1047646,);
nor I_61478 (I1047654,I1047646,I1047380);
DFFARX1 I_61479 (I1047654,I2507,I1047196,I1047167,);
nand I_61480 (I1047685,I1047646,I1047287);
nand I_61481 (I1047702,I1047380,I1047685);
nor I_61482 (I1047176,I1047702,I1047346);
not I_61483 (I1047757,I2514);
DFFARX1 I_61484 (I234128,I2507,I1047757,I1047783,);
DFFARX1 I_61485 (I1047783,I2507,I1047757,I1047800,);
not I_61486 (I1047749,I1047800);
not I_61487 (I1047822,I1047783);
DFFARX1 I_61488 (I234143,I2507,I1047757,I1047848,);
nand I_61489 (I1047856,I1047848,I234125);
not I_61490 (I1047873,I234125);
not I_61491 (I1047890,I234134);
nand I_61492 (I1047907,I234140,I234131);
and I_61493 (I1047924,I234140,I234131);
not I_61494 (I1047941,I234128);
nand I_61495 (I1047958,I1047941,I1047890);
nor I_61496 (I1047731,I1047958,I1047856);
nor I_61497 (I1047989,I1047873,I1047958);
nand I_61498 (I1047734,I1047924,I1047989);
not I_61499 (I1048020,I234125);
nor I_61500 (I1048037,I1048020,I234140);
nor I_61501 (I1048054,I1048037,I234128);
nor I_61502 (I1048071,I1047822,I1048054);
DFFARX1 I_61503 (I1048071,I2507,I1047757,I1047743,);
not I_61504 (I1048102,I1048037);
DFFARX1 I_61505 (I1048102,I2507,I1047757,I1047746,);
and I_61506 (I1047740,I1047848,I1048037);
nor I_61507 (I1048147,I1048020,I234149);
and I_61508 (I1048164,I1048147,I234146);
or I_61509 (I1048181,I1048164,I234137);
DFFARX1 I_61510 (I1048181,I2507,I1047757,I1048207,);
nor I_61511 (I1048215,I1048207,I1047941);
DFFARX1 I_61512 (I1048215,I2507,I1047757,I1047728,);
nand I_61513 (I1048246,I1048207,I1047848);
nand I_61514 (I1048263,I1047941,I1048246);
nor I_61515 (I1047737,I1048263,I1047907);
not I_61516 (I1048318,I2514);
DFFARX1 I_61517 (I437639,I2507,I1048318,I1048344,);
DFFARX1 I_61518 (I1048344,I2507,I1048318,I1048361,);
not I_61519 (I1048310,I1048361);
not I_61520 (I1048383,I1048344);
DFFARX1 I_61521 (I437627,I2507,I1048318,I1048409,);
nand I_61522 (I1048417,I1048409,I437633);
not I_61523 (I1048434,I437633);
not I_61524 (I1048451,I437630);
nand I_61525 (I1048468,I437618,I437615);
and I_61526 (I1048485,I437618,I437615);
not I_61527 (I1048502,I437642);
nand I_61528 (I1048519,I1048502,I1048451);
nor I_61529 (I1048292,I1048519,I1048417);
nor I_61530 (I1048550,I1048434,I1048519);
nand I_61531 (I1048295,I1048485,I1048550);
not I_61532 (I1048581,I437615);
nor I_61533 (I1048598,I1048581,I437618);
nor I_61534 (I1048615,I1048598,I437642);
nor I_61535 (I1048632,I1048383,I1048615);
DFFARX1 I_61536 (I1048632,I2507,I1048318,I1048304,);
not I_61537 (I1048663,I1048598);
DFFARX1 I_61538 (I1048663,I2507,I1048318,I1048307,);
and I_61539 (I1048301,I1048409,I1048598);
nor I_61540 (I1048708,I1048581,I437624);
and I_61541 (I1048725,I1048708,I437621);
or I_61542 (I1048742,I1048725,I437636);
DFFARX1 I_61543 (I1048742,I2507,I1048318,I1048768,);
nor I_61544 (I1048776,I1048768,I1048502);
DFFARX1 I_61545 (I1048776,I2507,I1048318,I1048289,);
nand I_61546 (I1048807,I1048768,I1048409);
nand I_61547 (I1048824,I1048502,I1048807);
nor I_61548 (I1048298,I1048824,I1048468);
not I_61549 (I1048879,I2514);
DFFARX1 I_61550 (I182958,I2507,I1048879,I1048905,);
DFFARX1 I_61551 (I1048905,I2507,I1048879,I1048922,);
not I_61552 (I1048871,I1048922);
not I_61553 (I1048944,I1048905);
DFFARX1 I_61554 (I182973,I2507,I1048879,I1048970,);
nand I_61555 (I1048978,I1048970,I182955);
not I_61556 (I1048995,I182955);
not I_61557 (I1049012,I182964);
nand I_61558 (I1049029,I182970,I182961);
and I_61559 (I1049046,I182970,I182961);
not I_61560 (I1049063,I182958);
nand I_61561 (I1049080,I1049063,I1049012);
nor I_61562 (I1048853,I1049080,I1048978);
nor I_61563 (I1049111,I1048995,I1049080);
nand I_61564 (I1048856,I1049046,I1049111);
not I_61565 (I1049142,I182955);
nor I_61566 (I1049159,I1049142,I182970);
nor I_61567 (I1049176,I1049159,I182958);
nor I_61568 (I1049193,I1048944,I1049176);
DFFARX1 I_61569 (I1049193,I2507,I1048879,I1048865,);
not I_61570 (I1049224,I1049159);
DFFARX1 I_61571 (I1049224,I2507,I1048879,I1048868,);
and I_61572 (I1048862,I1048970,I1049159);
nor I_61573 (I1049269,I1049142,I182979);
and I_61574 (I1049286,I1049269,I182976);
or I_61575 (I1049303,I1049286,I182967);
DFFARX1 I_61576 (I1049303,I2507,I1048879,I1049329,);
nor I_61577 (I1049337,I1049329,I1049063);
DFFARX1 I_61578 (I1049337,I2507,I1048879,I1048850,);
nand I_61579 (I1049368,I1049329,I1048970);
nand I_61580 (I1049385,I1049063,I1049368);
nor I_61581 (I1048859,I1049385,I1049029);
not I_61582 (I1049440,I2514);
DFFARX1 I_61583 (I609332,I2507,I1049440,I1049466,);
DFFARX1 I_61584 (I1049466,I2507,I1049440,I1049483,);
not I_61585 (I1049432,I1049483);
not I_61586 (I1049505,I1049466);
DFFARX1 I_61587 (I609347,I2507,I1049440,I1049531,);
nand I_61588 (I1049539,I1049531,I609338);
not I_61589 (I1049556,I609338);
not I_61590 (I1049573,I609344);
nand I_61591 (I1049590,I609341,I609350);
and I_61592 (I1049607,I609341,I609350);
not I_61593 (I1049624,I609335);
nand I_61594 (I1049641,I1049624,I1049573);
nor I_61595 (I1049414,I1049641,I1049539);
nor I_61596 (I1049672,I1049556,I1049641);
nand I_61597 (I1049417,I1049607,I1049672);
not I_61598 (I1049703,I609332);
nor I_61599 (I1049720,I1049703,I609341);
nor I_61600 (I1049737,I1049720,I609335);
nor I_61601 (I1049754,I1049505,I1049737);
DFFARX1 I_61602 (I1049754,I2507,I1049440,I1049426,);
not I_61603 (I1049785,I1049720);
DFFARX1 I_61604 (I1049785,I2507,I1049440,I1049429,);
and I_61605 (I1049423,I1049531,I1049720);
nor I_61606 (I1049830,I1049703,I609356);
and I_61607 (I1049847,I1049830,I609335);
or I_61608 (I1049864,I1049847,I609353);
DFFARX1 I_61609 (I1049864,I2507,I1049440,I1049890,);
nor I_61610 (I1049898,I1049890,I1049624);
DFFARX1 I_61611 (I1049898,I2507,I1049440,I1049411,);
nand I_61612 (I1049929,I1049890,I1049531);
nand I_61613 (I1049946,I1049624,I1049929);
nor I_61614 (I1049420,I1049946,I1049590);
not I_61615 (I1050001,I2514);
DFFARX1 I_61616 (I407719,I2507,I1050001,I1050027,);
DFFARX1 I_61617 (I1050027,I2507,I1050001,I1050044,);
not I_61618 (I1049993,I1050044);
not I_61619 (I1050066,I1050027);
DFFARX1 I_61620 (I407707,I2507,I1050001,I1050092,);
nand I_61621 (I1050100,I1050092,I407713);
not I_61622 (I1050117,I407713);
not I_61623 (I1050134,I407710);
nand I_61624 (I1050151,I407698,I407695);
and I_61625 (I1050168,I407698,I407695);
not I_61626 (I1050185,I407722);
nand I_61627 (I1050202,I1050185,I1050134);
nor I_61628 (I1049975,I1050202,I1050100);
nor I_61629 (I1050233,I1050117,I1050202);
nand I_61630 (I1049978,I1050168,I1050233);
not I_61631 (I1050264,I407695);
nor I_61632 (I1050281,I1050264,I407698);
nor I_61633 (I1050298,I1050281,I407722);
nor I_61634 (I1050315,I1050066,I1050298);
DFFARX1 I_61635 (I1050315,I2507,I1050001,I1049987,);
not I_61636 (I1050346,I1050281);
DFFARX1 I_61637 (I1050346,I2507,I1050001,I1049990,);
and I_61638 (I1049984,I1050092,I1050281);
nor I_61639 (I1050391,I1050264,I407704);
and I_61640 (I1050408,I1050391,I407701);
or I_61641 (I1050425,I1050408,I407716);
DFFARX1 I_61642 (I1050425,I2507,I1050001,I1050451,);
nor I_61643 (I1050459,I1050451,I1050185);
DFFARX1 I_61644 (I1050459,I2507,I1050001,I1049972,);
nand I_61645 (I1050490,I1050451,I1050092);
nand I_61646 (I1050507,I1050185,I1050490);
nor I_61647 (I1049981,I1050507,I1050151);
not I_61648 (I1050562,I2514);
DFFARX1 I_61649 (I439815,I2507,I1050562,I1050588,);
DFFARX1 I_61650 (I1050588,I2507,I1050562,I1050605,);
not I_61651 (I1050554,I1050605);
not I_61652 (I1050627,I1050588);
DFFARX1 I_61653 (I439803,I2507,I1050562,I1050653,);
nand I_61654 (I1050661,I1050653,I439809);
not I_61655 (I1050678,I439809);
not I_61656 (I1050695,I439806);
nand I_61657 (I1050712,I439794,I439791);
and I_61658 (I1050729,I439794,I439791);
not I_61659 (I1050746,I439818);
nand I_61660 (I1050763,I1050746,I1050695);
nor I_61661 (I1050536,I1050763,I1050661);
nor I_61662 (I1050794,I1050678,I1050763);
nand I_61663 (I1050539,I1050729,I1050794);
not I_61664 (I1050825,I439791);
nor I_61665 (I1050842,I1050825,I439794);
nor I_61666 (I1050859,I1050842,I439818);
nor I_61667 (I1050876,I1050627,I1050859);
DFFARX1 I_61668 (I1050876,I2507,I1050562,I1050548,);
not I_61669 (I1050907,I1050842);
DFFARX1 I_61670 (I1050907,I2507,I1050562,I1050551,);
and I_61671 (I1050545,I1050653,I1050842);
nor I_61672 (I1050952,I1050825,I439800);
and I_61673 (I1050969,I1050952,I439797);
or I_61674 (I1050986,I1050969,I439812);
DFFARX1 I_61675 (I1050986,I2507,I1050562,I1051012,);
nor I_61676 (I1051020,I1051012,I1050746);
DFFARX1 I_61677 (I1051020,I2507,I1050562,I1050533,);
nand I_61678 (I1051051,I1051012,I1050653);
nand I_61679 (I1051068,I1050746,I1051051);
nor I_61680 (I1050542,I1051068,I1050712);
not I_61681 (I1051123,I2514);
DFFARX1 I_61682 (I1075725,I2507,I1051123,I1051149,);
DFFARX1 I_61683 (I1051149,I2507,I1051123,I1051166,);
not I_61684 (I1051115,I1051166);
not I_61685 (I1051188,I1051149);
DFFARX1 I_61686 (I1075716,I2507,I1051123,I1051214,);
nand I_61687 (I1051222,I1051214,I1075713);
not I_61688 (I1051239,I1075713);
not I_61689 (I1051256,I1075722);
nand I_61690 (I1051273,I1075731,I1075713);
and I_61691 (I1051290,I1075731,I1075713);
not I_61692 (I1051307,I1075710);
nand I_61693 (I1051324,I1051307,I1051256);
nor I_61694 (I1051097,I1051324,I1051222);
nor I_61695 (I1051355,I1051239,I1051324);
nand I_61696 (I1051100,I1051290,I1051355);
not I_61697 (I1051386,I1075719);
nor I_61698 (I1051403,I1051386,I1075731);
nor I_61699 (I1051420,I1051403,I1075710);
nor I_61700 (I1051437,I1051188,I1051420);
DFFARX1 I_61701 (I1051437,I2507,I1051123,I1051109,);
not I_61702 (I1051468,I1051403);
DFFARX1 I_61703 (I1051468,I2507,I1051123,I1051112,);
and I_61704 (I1051106,I1051214,I1051403);
nor I_61705 (I1051513,I1051386,I1075734);
and I_61706 (I1051530,I1051513,I1075710);
or I_61707 (I1051547,I1051530,I1075728);
DFFARX1 I_61708 (I1051547,I2507,I1051123,I1051573,);
nor I_61709 (I1051581,I1051573,I1051307);
DFFARX1 I_61710 (I1051581,I2507,I1051123,I1051094,);
nand I_61711 (I1051612,I1051573,I1051214);
nand I_61712 (I1051629,I1051307,I1051612);
nor I_61713 (I1051103,I1051629,I1051273);
not I_61714 (I1051684,I2514);
DFFARX1 I_61715 (I1323177,I2507,I1051684,I1051710,);
DFFARX1 I_61716 (I1051710,I2507,I1051684,I1051727,);
not I_61717 (I1051676,I1051727);
not I_61718 (I1051749,I1051710);
DFFARX1 I_61719 (I1323171,I2507,I1051684,I1051775,);
nand I_61720 (I1051783,I1051775,I1323162);
not I_61721 (I1051800,I1323162);
not I_61722 (I1051817,I1323189);
nand I_61723 (I1051834,I1323174,I1323183);
and I_61724 (I1051851,I1323174,I1323183);
not I_61725 (I1051868,I1323168);
nand I_61726 (I1051885,I1051868,I1051817);
nor I_61727 (I1051658,I1051885,I1051783);
nor I_61728 (I1051916,I1051800,I1051885);
nand I_61729 (I1051661,I1051851,I1051916);
not I_61730 (I1051947,I1323186);
nor I_61731 (I1051964,I1051947,I1323174);
nor I_61732 (I1051981,I1051964,I1323168);
nor I_61733 (I1051998,I1051749,I1051981);
DFFARX1 I_61734 (I1051998,I2507,I1051684,I1051670,);
not I_61735 (I1052029,I1051964);
DFFARX1 I_61736 (I1052029,I2507,I1051684,I1051673,);
and I_61737 (I1051667,I1051775,I1051964);
nor I_61738 (I1052074,I1051947,I1323180);
and I_61739 (I1052091,I1052074,I1323162);
or I_61740 (I1052108,I1052091,I1323165);
DFFARX1 I_61741 (I1052108,I2507,I1051684,I1052134,);
nor I_61742 (I1052142,I1052134,I1051868);
DFFARX1 I_61743 (I1052142,I2507,I1051684,I1051655,);
nand I_61744 (I1052173,I1052134,I1051775);
nand I_61745 (I1052190,I1051868,I1052173);
nor I_61746 (I1051664,I1052190,I1051834);
not I_61747 (I1052245,I2514);
DFFARX1 I_61748 (I1332697,I2507,I1052245,I1052271,);
DFFARX1 I_61749 (I1052271,I2507,I1052245,I1052288,);
not I_61750 (I1052237,I1052288);
not I_61751 (I1052310,I1052271);
DFFARX1 I_61752 (I1332691,I2507,I1052245,I1052336,);
nand I_61753 (I1052344,I1052336,I1332682);
not I_61754 (I1052361,I1332682);
not I_61755 (I1052378,I1332709);
nand I_61756 (I1052395,I1332694,I1332703);
and I_61757 (I1052412,I1332694,I1332703);
not I_61758 (I1052429,I1332688);
nand I_61759 (I1052446,I1052429,I1052378);
nor I_61760 (I1052219,I1052446,I1052344);
nor I_61761 (I1052477,I1052361,I1052446);
nand I_61762 (I1052222,I1052412,I1052477);
not I_61763 (I1052508,I1332706);
nor I_61764 (I1052525,I1052508,I1332694);
nor I_61765 (I1052542,I1052525,I1332688);
nor I_61766 (I1052559,I1052310,I1052542);
DFFARX1 I_61767 (I1052559,I2507,I1052245,I1052231,);
not I_61768 (I1052590,I1052525);
DFFARX1 I_61769 (I1052590,I2507,I1052245,I1052234,);
and I_61770 (I1052228,I1052336,I1052525);
nor I_61771 (I1052635,I1052508,I1332700);
and I_61772 (I1052652,I1052635,I1332682);
or I_61773 (I1052669,I1052652,I1332685);
DFFARX1 I_61774 (I1052669,I2507,I1052245,I1052695,);
nor I_61775 (I1052703,I1052695,I1052429);
DFFARX1 I_61776 (I1052703,I2507,I1052245,I1052216,);
nand I_61777 (I1052734,I1052695,I1052336);
nand I_61778 (I1052751,I1052429,I1052734);
nor I_61779 (I1052225,I1052751,I1052395);
not I_61780 (I1052806,I2514);
DFFARX1 I_61781 (I419687,I2507,I1052806,I1052832,);
DFFARX1 I_61782 (I1052832,I2507,I1052806,I1052849,);
not I_61783 (I1052798,I1052849);
not I_61784 (I1052871,I1052832);
DFFARX1 I_61785 (I419675,I2507,I1052806,I1052897,);
nand I_61786 (I1052905,I1052897,I419681);
not I_61787 (I1052922,I419681);
not I_61788 (I1052939,I419678);
nand I_61789 (I1052956,I419666,I419663);
and I_61790 (I1052973,I419666,I419663);
not I_61791 (I1052990,I419690);
nand I_61792 (I1053007,I1052990,I1052939);
nor I_61793 (I1052780,I1053007,I1052905);
nor I_61794 (I1053038,I1052922,I1053007);
nand I_61795 (I1052783,I1052973,I1053038);
not I_61796 (I1053069,I419663);
nor I_61797 (I1053086,I1053069,I419666);
nor I_61798 (I1053103,I1053086,I419690);
nor I_61799 (I1053120,I1052871,I1053103);
DFFARX1 I_61800 (I1053120,I2507,I1052806,I1052792,);
not I_61801 (I1053151,I1053086);
DFFARX1 I_61802 (I1053151,I2507,I1052806,I1052795,);
and I_61803 (I1052789,I1052897,I1053086);
nor I_61804 (I1053196,I1053069,I419672);
and I_61805 (I1053213,I1053196,I419669);
or I_61806 (I1053230,I1053213,I419684);
DFFARX1 I_61807 (I1053230,I2507,I1052806,I1053256,);
nor I_61808 (I1053264,I1053256,I1052990);
DFFARX1 I_61809 (I1053264,I2507,I1052806,I1052777,);
nand I_61810 (I1053295,I1053256,I1052897);
nand I_61811 (I1053312,I1052990,I1053295);
nor I_61812 (I1052786,I1053312,I1052956);
not I_61813 (I1053367,I2514);
DFFARX1 I_61814 (I1063009,I2507,I1053367,I1053393,);
DFFARX1 I_61815 (I1053393,I2507,I1053367,I1053410,);
not I_61816 (I1053359,I1053410);
not I_61817 (I1053432,I1053393);
DFFARX1 I_61818 (I1063000,I2507,I1053367,I1053458,);
nand I_61819 (I1053466,I1053458,I1062997);
not I_61820 (I1053483,I1062997);
not I_61821 (I1053500,I1063006);
nand I_61822 (I1053517,I1063015,I1062997);
and I_61823 (I1053534,I1063015,I1062997);
not I_61824 (I1053551,I1062994);
nand I_61825 (I1053568,I1053551,I1053500);
nor I_61826 (I1053341,I1053568,I1053466);
nor I_61827 (I1053599,I1053483,I1053568);
nand I_61828 (I1053344,I1053534,I1053599);
not I_61829 (I1053630,I1063003);
nor I_61830 (I1053647,I1053630,I1063015);
nor I_61831 (I1053664,I1053647,I1062994);
nor I_61832 (I1053681,I1053432,I1053664);
DFFARX1 I_61833 (I1053681,I2507,I1053367,I1053353,);
not I_61834 (I1053712,I1053647);
DFFARX1 I_61835 (I1053712,I2507,I1053367,I1053356,);
and I_61836 (I1053350,I1053458,I1053647);
nor I_61837 (I1053757,I1053630,I1063018);
and I_61838 (I1053774,I1053757,I1062994);
or I_61839 (I1053791,I1053774,I1063012);
DFFARX1 I_61840 (I1053791,I2507,I1053367,I1053817,);
nor I_61841 (I1053825,I1053817,I1053551);
DFFARX1 I_61842 (I1053825,I2507,I1053367,I1053338,);
nand I_61843 (I1053856,I1053817,I1053458);
nand I_61844 (I1053873,I1053551,I1053856);
nor I_61845 (I1053347,I1053873,I1053517);
not I_61846 (I1053928,I2514);
DFFARX1 I_61847 (I1210696,I2507,I1053928,I1053954,);
DFFARX1 I_61848 (I1053954,I2507,I1053928,I1053971,);
not I_61849 (I1053920,I1053971);
not I_61850 (I1053993,I1053954);
DFFARX1 I_61851 (I1210702,I2507,I1053928,I1054019,);
nand I_61852 (I1054027,I1054019,I1210711);
not I_61853 (I1054044,I1210711);
not I_61854 (I1054061,I1210690);
nand I_61855 (I1054078,I1210693,I1210693);
and I_61856 (I1054095,I1210693,I1210693);
not I_61857 (I1054112,I1210705);
nand I_61858 (I1054129,I1054112,I1054061);
nor I_61859 (I1053902,I1054129,I1054027);
nor I_61860 (I1054160,I1054044,I1054129);
nand I_61861 (I1053905,I1054095,I1054160);
not I_61862 (I1054191,I1210699);
nor I_61863 (I1054208,I1054191,I1210693);
nor I_61864 (I1054225,I1054208,I1210705);
nor I_61865 (I1054242,I1053993,I1054225);
DFFARX1 I_61866 (I1054242,I2507,I1053928,I1053914,);
not I_61867 (I1054273,I1054208);
DFFARX1 I_61868 (I1054273,I2507,I1053928,I1053917,);
and I_61869 (I1053911,I1054019,I1054208);
nor I_61870 (I1054318,I1054191,I1210714);
and I_61871 (I1054335,I1054318,I1210690);
or I_61872 (I1054352,I1054335,I1210708);
DFFARX1 I_61873 (I1054352,I2507,I1053928,I1054378,);
nor I_61874 (I1054386,I1054378,I1054112);
DFFARX1 I_61875 (I1054386,I2507,I1053928,I1053899,);
nand I_61876 (I1054417,I1054378,I1054019);
nand I_61877 (I1054434,I1054112,I1054417);
nor I_61878 (I1053908,I1054434,I1054078);
not I_61879 (I1054489,I2514);
DFFARX1 I_61880 (I198428,I2507,I1054489,I1054515,);
DFFARX1 I_61881 (I1054515,I2507,I1054489,I1054532,);
not I_61882 (I1054481,I1054532);
not I_61883 (I1054554,I1054515);
DFFARX1 I_61884 (I198443,I2507,I1054489,I1054580,);
nand I_61885 (I1054588,I1054580,I198425);
not I_61886 (I1054605,I198425);
not I_61887 (I1054622,I198434);
nand I_61888 (I1054639,I198440,I198431);
and I_61889 (I1054656,I198440,I198431);
not I_61890 (I1054673,I198428);
nand I_61891 (I1054690,I1054673,I1054622);
nor I_61892 (I1054463,I1054690,I1054588);
nor I_61893 (I1054721,I1054605,I1054690);
nand I_61894 (I1054466,I1054656,I1054721);
not I_61895 (I1054752,I198425);
nor I_61896 (I1054769,I1054752,I198440);
nor I_61897 (I1054786,I1054769,I198428);
nor I_61898 (I1054803,I1054554,I1054786);
DFFARX1 I_61899 (I1054803,I2507,I1054489,I1054475,);
not I_61900 (I1054834,I1054769);
DFFARX1 I_61901 (I1054834,I2507,I1054489,I1054478,);
and I_61902 (I1054472,I1054580,I1054769);
nor I_61903 (I1054879,I1054752,I198449);
and I_61904 (I1054896,I1054879,I198446);
or I_61905 (I1054913,I1054896,I198437);
DFFARX1 I_61906 (I1054913,I2507,I1054489,I1054939,);
nor I_61907 (I1054947,I1054939,I1054673);
DFFARX1 I_61908 (I1054947,I2507,I1054489,I1054460,);
nand I_61909 (I1054978,I1054939,I1054580);
nand I_61910 (I1054995,I1054673,I1054978);
nor I_61911 (I1054469,I1054995,I1054639);
not I_61912 (I1055050,I2514);
DFFARX1 I_61913 (I678117,I2507,I1055050,I1055076,);
DFFARX1 I_61914 (I1055076,I2507,I1055050,I1055093,);
not I_61915 (I1055042,I1055093);
not I_61916 (I1055115,I1055076);
DFFARX1 I_61917 (I678129,I2507,I1055050,I1055141,);
nand I_61918 (I1055149,I1055141,I678138);
not I_61919 (I1055166,I678138);
not I_61920 (I1055183,I678120);
nand I_61921 (I1055200,I678123,I678114);
and I_61922 (I1055217,I678123,I678114);
not I_61923 (I1055234,I678132);
nand I_61924 (I1055251,I1055234,I1055183);
nor I_61925 (I1055024,I1055251,I1055149);
nor I_61926 (I1055282,I1055166,I1055251);
nand I_61927 (I1055027,I1055217,I1055282);
not I_61928 (I1055313,I678135);
nor I_61929 (I1055330,I1055313,I678123);
nor I_61930 (I1055347,I1055330,I678132);
nor I_61931 (I1055364,I1055115,I1055347);
DFFARX1 I_61932 (I1055364,I2507,I1055050,I1055036,);
not I_61933 (I1055395,I1055330);
DFFARX1 I_61934 (I1055395,I2507,I1055050,I1055039,);
and I_61935 (I1055033,I1055141,I1055330);
nor I_61936 (I1055440,I1055313,I678114);
and I_61937 (I1055457,I1055440,I678126);
or I_61938 (I1055474,I1055457,I678117);
DFFARX1 I_61939 (I1055474,I2507,I1055050,I1055500,);
nor I_61940 (I1055508,I1055500,I1055234);
DFFARX1 I_61941 (I1055508,I2507,I1055050,I1055021,);
nand I_61942 (I1055539,I1055500,I1055141);
nand I_61943 (I1055556,I1055234,I1055539);
nor I_61944 (I1055030,I1055556,I1055200);
not I_61945 (I1055611,I2514);
DFFARX1 I_61946 (I646905,I2507,I1055611,I1055637,);
DFFARX1 I_61947 (I1055637,I2507,I1055611,I1055654,);
not I_61948 (I1055603,I1055654);
not I_61949 (I1055676,I1055637);
DFFARX1 I_61950 (I646917,I2507,I1055611,I1055702,);
nand I_61951 (I1055710,I1055702,I646926);
not I_61952 (I1055727,I646926);
not I_61953 (I1055744,I646908);
nand I_61954 (I1055761,I646911,I646902);
and I_61955 (I1055778,I646911,I646902);
not I_61956 (I1055795,I646920);
nand I_61957 (I1055812,I1055795,I1055744);
nor I_61958 (I1055585,I1055812,I1055710);
nor I_61959 (I1055843,I1055727,I1055812);
nand I_61960 (I1055588,I1055778,I1055843);
not I_61961 (I1055874,I646923);
nor I_61962 (I1055891,I1055874,I646911);
nor I_61963 (I1055908,I1055891,I646920);
nor I_61964 (I1055925,I1055676,I1055908);
DFFARX1 I_61965 (I1055925,I2507,I1055611,I1055597,);
not I_61966 (I1055956,I1055891);
DFFARX1 I_61967 (I1055956,I2507,I1055611,I1055600,);
and I_61968 (I1055594,I1055702,I1055891);
nor I_61969 (I1056001,I1055874,I646902);
and I_61970 (I1056018,I1056001,I646914);
or I_61971 (I1056035,I1056018,I646905);
DFFARX1 I_61972 (I1056035,I2507,I1055611,I1056061,);
nor I_61973 (I1056069,I1056061,I1055795);
DFFARX1 I_61974 (I1056069,I2507,I1055611,I1055582,);
nand I_61975 (I1056100,I1056061,I1055702);
nand I_61976 (I1056117,I1055795,I1056100);
nor I_61977 (I1055591,I1056117,I1055761);
not I_61978 (I1056172,I2514);
DFFARX1 I_61979 (I368259,I2507,I1056172,I1056198,);
DFFARX1 I_61980 (I1056198,I2507,I1056172,I1056215,);
not I_61981 (I1056164,I1056215);
not I_61982 (I1056237,I1056198);
DFFARX1 I_61983 (I368256,I2507,I1056172,I1056263,);
nand I_61984 (I1056271,I1056263,I368250);
not I_61985 (I1056288,I368250);
not I_61986 (I1056305,I368247);
nand I_61987 (I1056322,I368241,I368238);
and I_61988 (I1056339,I368241,I368238);
not I_61989 (I1056356,I368253);
nand I_61990 (I1056373,I1056356,I1056305);
nor I_61991 (I1056146,I1056373,I1056271);
nor I_61992 (I1056404,I1056288,I1056373);
nand I_61993 (I1056149,I1056339,I1056404);
not I_61994 (I1056435,I368265);
nor I_61995 (I1056452,I1056435,I368241);
nor I_61996 (I1056469,I1056452,I368253);
nor I_61997 (I1056486,I1056237,I1056469);
DFFARX1 I_61998 (I1056486,I2507,I1056172,I1056158,);
not I_61999 (I1056517,I1056452);
DFFARX1 I_62000 (I1056517,I2507,I1056172,I1056161,);
and I_62001 (I1056155,I1056263,I1056452);
nor I_62002 (I1056562,I1056435,I368262);
and I_62003 (I1056579,I1056562,I368238);
or I_62004 (I1056596,I1056579,I368244);
DFFARX1 I_62005 (I1056596,I2507,I1056172,I1056622,);
nor I_62006 (I1056630,I1056622,I1056356);
DFFARX1 I_62007 (I1056630,I2507,I1056172,I1056143,);
nand I_62008 (I1056661,I1056622,I1056263);
nand I_62009 (I1056678,I1056356,I1056661);
nor I_62010 (I1056152,I1056678,I1056322);
not I_62011 (I1056733,I2514);
DFFARX1 I_62012 (I1137571,I2507,I1056733,I1056759,);
DFFARX1 I_62013 (I1056759,I2507,I1056733,I1056776,);
not I_62014 (I1056725,I1056776);
not I_62015 (I1056798,I1056759);
DFFARX1 I_62016 (I1137562,I2507,I1056733,I1056824,);
nand I_62017 (I1056832,I1056824,I1137559);
not I_62018 (I1056849,I1137559);
not I_62019 (I1056866,I1137568);
nand I_62020 (I1056883,I1137577,I1137559);
and I_62021 (I1056900,I1137577,I1137559);
not I_62022 (I1056917,I1137556);
nand I_62023 (I1056934,I1056917,I1056866);
nor I_62024 (I1056707,I1056934,I1056832);
nor I_62025 (I1056965,I1056849,I1056934);
nand I_62026 (I1056710,I1056900,I1056965);
not I_62027 (I1056996,I1137565);
nor I_62028 (I1057013,I1056996,I1137577);
nor I_62029 (I1057030,I1057013,I1137556);
nor I_62030 (I1057047,I1056798,I1057030);
DFFARX1 I_62031 (I1057047,I2507,I1056733,I1056719,);
not I_62032 (I1057078,I1057013);
DFFARX1 I_62033 (I1057078,I2507,I1056733,I1056722,);
and I_62034 (I1056716,I1056824,I1057013);
nor I_62035 (I1057123,I1056996,I1137580);
and I_62036 (I1057140,I1057123,I1137556);
or I_62037 (I1057157,I1057140,I1137574);
DFFARX1 I_62038 (I1057157,I2507,I1056733,I1057183,);
nor I_62039 (I1057191,I1057183,I1056917);
DFFARX1 I_62040 (I1057191,I2507,I1056733,I1056704,);
nand I_62041 (I1057222,I1057183,I1056824);
nand I_62042 (I1057239,I1056917,I1057222);
nor I_62043 (I1056713,I1057239,I1056883);
not I_62044 (I1057294,I2514);
DFFARX1 I_62045 (I294479,I2507,I1057294,I1057320,);
DFFARX1 I_62046 (I1057320,I2507,I1057294,I1057337,);
not I_62047 (I1057286,I1057337);
not I_62048 (I1057359,I1057320);
DFFARX1 I_62049 (I294476,I2507,I1057294,I1057385,);
nand I_62050 (I1057393,I1057385,I294470);
not I_62051 (I1057410,I294470);
not I_62052 (I1057427,I294467);
nand I_62053 (I1057444,I294461,I294458);
and I_62054 (I1057461,I294461,I294458);
not I_62055 (I1057478,I294473);
nand I_62056 (I1057495,I1057478,I1057427);
nor I_62057 (I1057268,I1057495,I1057393);
nor I_62058 (I1057526,I1057410,I1057495);
nand I_62059 (I1057271,I1057461,I1057526);
not I_62060 (I1057557,I294485);
nor I_62061 (I1057574,I1057557,I294461);
nor I_62062 (I1057591,I1057574,I294473);
nor I_62063 (I1057608,I1057359,I1057591);
DFFARX1 I_62064 (I1057608,I2507,I1057294,I1057280,);
not I_62065 (I1057639,I1057574);
DFFARX1 I_62066 (I1057639,I2507,I1057294,I1057283,);
and I_62067 (I1057277,I1057385,I1057574);
nor I_62068 (I1057684,I1057557,I294482);
and I_62069 (I1057701,I1057684,I294458);
or I_62070 (I1057718,I1057701,I294464);
DFFARX1 I_62071 (I1057718,I2507,I1057294,I1057744,);
nor I_62072 (I1057752,I1057744,I1057478);
DFFARX1 I_62073 (I1057752,I2507,I1057294,I1057265,);
nand I_62074 (I1057783,I1057744,I1057385);
nand I_62075 (I1057800,I1057478,I1057783);
nor I_62076 (I1057274,I1057800,I1057444);
not I_62077 (I1057855,I2514);
DFFARX1 I_62078 (I381063,I2507,I1057855,I1057881,);
DFFARX1 I_62079 (I1057881,I2507,I1057855,I1057898,);
not I_62080 (I1057847,I1057898);
not I_62081 (I1057920,I1057881);
DFFARX1 I_62082 (I381051,I2507,I1057855,I1057946,);
nand I_62083 (I1057954,I1057946,I381057);
not I_62084 (I1057971,I381057);
not I_62085 (I1057988,I381054);
nand I_62086 (I1058005,I381042,I381039);
and I_62087 (I1058022,I381042,I381039);
not I_62088 (I1058039,I381066);
nand I_62089 (I1058056,I1058039,I1057988);
nor I_62090 (I1057829,I1058056,I1057954);
nor I_62091 (I1058087,I1057971,I1058056);
nand I_62092 (I1057832,I1058022,I1058087);
not I_62093 (I1058118,I381039);
nor I_62094 (I1058135,I1058118,I381042);
nor I_62095 (I1058152,I1058135,I381066);
nor I_62096 (I1058169,I1057920,I1058152);
DFFARX1 I_62097 (I1058169,I2507,I1057855,I1057841,);
not I_62098 (I1058200,I1058135);
DFFARX1 I_62099 (I1058200,I2507,I1057855,I1057844,);
and I_62100 (I1057838,I1057946,I1058135);
nor I_62101 (I1058245,I1058118,I381048);
and I_62102 (I1058262,I1058245,I381045);
or I_62103 (I1058279,I1058262,I381060);
DFFARX1 I_62104 (I1058279,I2507,I1057855,I1058305,);
nor I_62105 (I1058313,I1058305,I1058039);
DFFARX1 I_62106 (I1058313,I2507,I1057855,I1057826,);
nand I_62107 (I1058344,I1058305,I1057946);
nand I_62108 (I1058361,I1058039,I1058344);
nor I_62109 (I1057835,I1058361,I1058005);
not I_62110 (I1058416,I2514);
DFFARX1 I_62111 (I845998,I2507,I1058416,I1058442,);
DFFARX1 I_62112 (I1058442,I2507,I1058416,I1058459,);
not I_62113 (I1058408,I1058459);
not I_62114 (I1058481,I1058442);
DFFARX1 I_62115 (I845995,I2507,I1058416,I1058507,);
nand I_62116 (I1058515,I1058507,I846010);
not I_62117 (I1058532,I846010);
not I_62118 (I1058549,I846007);
nand I_62119 (I1058566,I846004,I845992);
and I_62120 (I1058583,I846004,I845992);
not I_62121 (I1058600,I845989);
nand I_62122 (I1058617,I1058600,I1058549);
nor I_62123 (I1058390,I1058617,I1058515);
nor I_62124 (I1058648,I1058532,I1058617);
nand I_62125 (I1058393,I1058583,I1058648);
not I_62126 (I1058679,I845995);
nor I_62127 (I1058696,I1058679,I846004);
nor I_62128 (I1058713,I1058696,I845989);
nor I_62129 (I1058730,I1058481,I1058713);
DFFARX1 I_62130 (I1058730,I2507,I1058416,I1058402,);
not I_62131 (I1058761,I1058696);
DFFARX1 I_62132 (I1058761,I2507,I1058416,I1058405,);
and I_62133 (I1058399,I1058507,I1058696);
nor I_62134 (I1058806,I1058679,I846001);
and I_62135 (I1058823,I1058806,I845989);
or I_62136 (I1058840,I1058823,I845992);
DFFARX1 I_62137 (I1058840,I2507,I1058416,I1058866,);
nor I_62138 (I1058874,I1058866,I1058600);
DFFARX1 I_62139 (I1058874,I2507,I1058416,I1058387,);
nand I_62140 (I1058905,I1058866,I1058507);
nand I_62141 (I1058922,I1058600,I1058905);
nor I_62142 (I1058396,I1058922,I1058566);
not I_62143 (I1058980,I2514);
DFFARX1 I_62144 (I240670,I2507,I1058980,I1059006,);
and I_62145 (I1059014,I1059006,I240673);
DFFARX1 I_62146 (I1059014,I2507,I1058980,I1058963,);
DFFARX1 I_62147 (I240673,I2507,I1058980,I1059054,);
not I_62148 (I1059062,I240688);
not I_62149 (I1059079,I240694);
nand I_62150 (I1059096,I1059079,I1059062);
nor I_62151 (I1058951,I1059054,I1059096);
DFFARX1 I_62152 (I1059096,I2507,I1058980,I1059136,);
not I_62153 (I1058972,I1059136);
not I_62154 (I1059158,I240682);
nand I_62155 (I1059175,I1059079,I1059158);
DFFARX1 I_62156 (I1059175,I2507,I1058980,I1059201,);
not I_62157 (I1059209,I1059201);
not I_62158 (I1059226,I240679);
nand I_62159 (I1059243,I1059226,I240676);
and I_62160 (I1059260,I1059062,I1059243);
nor I_62161 (I1059277,I1059175,I1059260);
DFFARX1 I_62162 (I1059277,I2507,I1058980,I1058948,);
DFFARX1 I_62163 (I1059260,I2507,I1058980,I1058969,);
nor I_62164 (I1059322,I240679,I240670);
nor I_62165 (I1058960,I1059175,I1059322);
or I_62166 (I1059353,I240679,I240670);
nor I_62167 (I1059370,I240685,I240691);
DFFARX1 I_62168 (I1059370,I2507,I1058980,I1059396,);
not I_62169 (I1059404,I1059396);
nor I_62170 (I1058966,I1059404,I1059209);
nand I_62171 (I1059435,I1059404,I1059054);
not I_62172 (I1059452,I240685);
nand I_62173 (I1059469,I1059452,I1059158);
nand I_62174 (I1059486,I1059404,I1059469);
nand I_62175 (I1058957,I1059486,I1059435);
nand I_62176 (I1058954,I1059469,I1059353);
not I_62177 (I1059558,I2514);
DFFARX1 I_62178 (I1032584,I2507,I1059558,I1059584,);
and I_62179 (I1059592,I1059584,I1032581);
DFFARX1 I_62180 (I1059592,I2507,I1059558,I1059541,);
DFFARX1 I_62181 (I1032587,I2507,I1059558,I1059632,);
not I_62182 (I1059640,I1032590);
not I_62183 (I1059657,I1032584);
nand I_62184 (I1059674,I1059657,I1059640);
nor I_62185 (I1059529,I1059632,I1059674);
DFFARX1 I_62186 (I1059674,I2507,I1059558,I1059714,);
not I_62187 (I1059550,I1059714);
not I_62188 (I1059736,I1032599);
nand I_62189 (I1059753,I1059657,I1059736);
DFFARX1 I_62190 (I1059753,I2507,I1059558,I1059779,);
not I_62191 (I1059787,I1059779);
not I_62192 (I1059804,I1032596);
nand I_62193 (I1059821,I1059804,I1032602);
and I_62194 (I1059838,I1059640,I1059821);
nor I_62195 (I1059855,I1059753,I1059838);
DFFARX1 I_62196 (I1059855,I2507,I1059558,I1059526,);
DFFARX1 I_62197 (I1059838,I2507,I1059558,I1059547,);
nor I_62198 (I1059900,I1032596,I1032581);
nor I_62199 (I1059538,I1059753,I1059900);
or I_62200 (I1059931,I1032596,I1032581);
nor I_62201 (I1059948,I1032593,I1032587);
DFFARX1 I_62202 (I1059948,I2507,I1059558,I1059974,);
not I_62203 (I1059982,I1059974);
nor I_62204 (I1059544,I1059982,I1059787);
nand I_62205 (I1060013,I1059982,I1059632);
not I_62206 (I1060030,I1032593);
nand I_62207 (I1060047,I1060030,I1059736);
nand I_62208 (I1060064,I1059982,I1060047);
nand I_62209 (I1059535,I1060064,I1060013);
nand I_62210 (I1059532,I1060047,I1059931);
not I_62211 (I1060136,I2514);
DFFARX1 I_62212 (I822804,I2507,I1060136,I1060162,);
and I_62213 (I1060170,I1060162,I822810);
DFFARX1 I_62214 (I1060170,I2507,I1060136,I1060119,);
DFFARX1 I_62215 (I822816,I2507,I1060136,I1060210,);
not I_62216 (I1060218,I822801);
not I_62217 (I1060235,I822801);
nand I_62218 (I1060252,I1060235,I1060218);
nor I_62219 (I1060107,I1060210,I1060252);
DFFARX1 I_62220 (I1060252,I2507,I1060136,I1060292,);
not I_62221 (I1060128,I1060292);
not I_62222 (I1060314,I822819);
nand I_62223 (I1060331,I1060235,I1060314);
DFFARX1 I_62224 (I1060331,I2507,I1060136,I1060357,);
not I_62225 (I1060365,I1060357);
not I_62226 (I1060382,I822813);
nand I_62227 (I1060399,I1060382,I822804);
and I_62228 (I1060416,I1060218,I1060399);
nor I_62229 (I1060433,I1060331,I1060416);
DFFARX1 I_62230 (I1060433,I2507,I1060136,I1060104,);
DFFARX1 I_62231 (I1060416,I2507,I1060136,I1060125,);
nor I_62232 (I1060478,I822813,I822822);
nor I_62233 (I1060116,I1060331,I1060478);
or I_62234 (I1060509,I822813,I822822);
nor I_62235 (I1060526,I822807,I822807);
DFFARX1 I_62236 (I1060526,I2507,I1060136,I1060552,);
not I_62237 (I1060560,I1060552);
nor I_62238 (I1060122,I1060560,I1060365);
nand I_62239 (I1060591,I1060560,I1060210);
not I_62240 (I1060608,I822807);
nand I_62241 (I1060625,I1060608,I1060314);
nand I_62242 (I1060642,I1060560,I1060625);
nand I_62243 (I1060113,I1060642,I1060591);
nand I_62244 (I1060110,I1060625,I1060509);
not I_62245 (I1060714,I2514);
DFFARX1 I_62246 (I731305,I2507,I1060714,I1060740,);
and I_62247 (I1060748,I1060740,I731293);
DFFARX1 I_62248 (I1060748,I2507,I1060714,I1060697,);
DFFARX1 I_62249 (I731296,I2507,I1060714,I1060788,);
not I_62250 (I1060796,I731290);
not I_62251 (I1060813,I731314);
nand I_62252 (I1060830,I1060813,I1060796);
nor I_62253 (I1060685,I1060788,I1060830);
DFFARX1 I_62254 (I1060830,I2507,I1060714,I1060870,);
not I_62255 (I1060706,I1060870);
not I_62256 (I1060892,I731302);
nand I_62257 (I1060909,I1060813,I1060892);
DFFARX1 I_62258 (I1060909,I2507,I1060714,I1060935,);
not I_62259 (I1060943,I1060935);
not I_62260 (I1060960,I731311);
nand I_62261 (I1060977,I1060960,I731308);
and I_62262 (I1060994,I1060796,I1060977);
nor I_62263 (I1061011,I1060909,I1060994);
DFFARX1 I_62264 (I1061011,I2507,I1060714,I1060682,);
DFFARX1 I_62265 (I1060994,I2507,I1060714,I1060703,);
nor I_62266 (I1061056,I731311,I731299);
nor I_62267 (I1060694,I1060909,I1061056);
or I_62268 (I1061087,I731311,I731299);
nor I_62269 (I1061104,I731290,I731293);
DFFARX1 I_62270 (I1061104,I2507,I1060714,I1061130,);
not I_62271 (I1061138,I1061130);
nor I_62272 (I1060700,I1061138,I1060943);
nand I_62273 (I1061169,I1061138,I1060788);
not I_62274 (I1061186,I731290);
nand I_62275 (I1061203,I1061186,I1060892);
nand I_62276 (I1061220,I1061138,I1061203);
nand I_62277 (I1060691,I1061220,I1061169);
nand I_62278 (I1060688,I1061203,I1061087);
not I_62279 (I1061292,I2514);
DFFARX1 I_62280 (I315038,I2507,I1061292,I1061318,);
and I_62281 (I1061326,I1061318,I315023);
DFFARX1 I_62282 (I1061326,I2507,I1061292,I1061275,);
DFFARX1 I_62283 (I315029,I2507,I1061292,I1061366,);
not I_62284 (I1061374,I315011);
not I_62285 (I1061391,I315032);
nand I_62286 (I1061408,I1061391,I1061374);
nor I_62287 (I1061263,I1061366,I1061408);
DFFARX1 I_62288 (I1061408,I2507,I1061292,I1061448,);
not I_62289 (I1061284,I1061448);
not I_62290 (I1061470,I315035);
nand I_62291 (I1061487,I1061391,I1061470);
DFFARX1 I_62292 (I1061487,I2507,I1061292,I1061513,);
not I_62293 (I1061521,I1061513);
not I_62294 (I1061538,I315026);
nand I_62295 (I1061555,I1061538,I315014);
and I_62296 (I1061572,I1061374,I1061555);
nor I_62297 (I1061589,I1061487,I1061572);
DFFARX1 I_62298 (I1061589,I2507,I1061292,I1061260,);
DFFARX1 I_62299 (I1061572,I2507,I1061292,I1061281,);
nor I_62300 (I1061634,I315026,I315020);
nor I_62301 (I1061272,I1061487,I1061634);
or I_62302 (I1061665,I315026,I315020);
nor I_62303 (I1061682,I315017,I315011);
DFFARX1 I_62304 (I1061682,I2507,I1061292,I1061708,);
not I_62305 (I1061716,I1061708);
nor I_62306 (I1061278,I1061716,I1061521);
nand I_62307 (I1061747,I1061716,I1061366);
not I_62308 (I1061764,I315017);
nand I_62309 (I1061781,I1061764,I1061470);
nand I_62310 (I1061798,I1061716,I1061781);
nand I_62311 (I1061269,I1061798,I1061747);
nand I_62312 (I1061266,I1061781,I1061665);
not I_62313 (I1061870,I2514);
DFFARX1 I_62314 (I85450,I2507,I1061870,I1061896,);
and I_62315 (I1061904,I1061896,I85426);
DFFARX1 I_62316 (I1061904,I2507,I1061870,I1061853,);
DFFARX1 I_62317 (I85444,I2507,I1061870,I1061944,);
not I_62318 (I1061952,I85432);
not I_62319 (I1061969,I85429);
nand I_62320 (I1061986,I1061969,I1061952);
nor I_62321 (I1061841,I1061944,I1061986);
DFFARX1 I_62322 (I1061986,I2507,I1061870,I1062026,);
not I_62323 (I1061862,I1062026);
not I_62324 (I1062048,I85438);
nand I_62325 (I1062065,I1061969,I1062048);
DFFARX1 I_62326 (I1062065,I2507,I1061870,I1062091,);
not I_62327 (I1062099,I1062091);
not I_62328 (I1062116,I85429);
nand I_62329 (I1062133,I1062116,I85447);
and I_62330 (I1062150,I1061952,I1062133);
nor I_62331 (I1062167,I1062065,I1062150);
DFFARX1 I_62332 (I1062167,I2507,I1061870,I1061838,);
DFFARX1 I_62333 (I1062150,I2507,I1061870,I1061859,);
nor I_62334 (I1062212,I85429,I85441);
nor I_62335 (I1061850,I1062065,I1062212);
or I_62336 (I1062243,I85429,I85441);
nor I_62337 (I1062260,I85435,I85426);
DFFARX1 I_62338 (I1062260,I2507,I1061870,I1062286,);
not I_62339 (I1062294,I1062286);
nor I_62340 (I1061856,I1062294,I1062099);
nand I_62341 (I1062325,I1062294,I1061944);
not I_62342 (I1062342,I85435);
nand I_62343 (I1062359,I1062342,I1062048);
nand I_62344 (I1062376,I1062294,I1062359);
nand I_62345 (I1061847,I1062376,I1062325);
nand I_62346 (I1061844,I1062359,I1062243);
not I_62347 (I1062448,I2514);
DFFARX1 I_62348 (I917939,I2507,I1062448,I1062474,);
and I_62349 (I1062482,I1062474,I917933);
DFFARX1 I_62350 (I1062482,I2507,I1062448,I1062431,);
DFFARX1 I_62351 (I917951,I2507,I1062448,I1062522,);
not I_62352 (I1062530,I917942);
not I_62353 (I1062547,I917954);
nand I_62354 (I1062564,I1062547,I1062530);
nor I_62355 (I1062419,I1062522,I1062564);
DFFARX1 I_62356 (I1062564,I2507,I1062448,I1062604,);
not I_62357 (I1062440,I1062604);
not I_62358 (I1062626,I917960);
nand I_62359 (I1062643,I1062547,I1062626);
DFFARX1 I_62360 (I1062643,I2507,I1062448,I1062669,);
not I_62361 (I1062677,I1062669);
not I_62362 (I1062694,I917936);
nand I_62363 (I1062711,I1062694,I917957);
and I_62364 (I1062728,I1062530,I1062711);
nor I_62365 (I1062745,I1062643,I1062728);
DFFARX1 I_62366 (I1062745,I2507,I1062448,I1062416,);
DFFARX1 I_62367 (I1062728,I2507,I1062448,I1062437,);
nor I_62368 (I1062790,I917936,I917948);
nor I_62369 (I1062428,I1062643,I1062790);
or I_62370 (I1062821,I917936,I917948);
nor I_62371 (I1062838,I917933,I917945);
DFFARX1 I_62372 (I1062838,I2507,I1062448,I1062864,);
not I_62373 (I1062872,I1062864);
nor I_62374 (I1062434,I1062872,I1062677);
nand I_62375 (I1062903,I1062872,I1062522);
not I_62376 (I1062920,I917933);
nand I_62377 (I1062937,I1062920,I1062626);
nand I_62378 (I1062954,I1062872,I1062937);
nand I_62379 (I1062425,I1062954,I1062903);
nand I_62380 (I1062422,I1062937,I1062821);
not I_62381 (I1063026,I2514);
DFFARX1 I_62382 (I260757,I2507,I1063026,I1063052,);
and I_62383 (I1063060,I1063052,I260742);
DFFARX1 I_62384 (I1063060,I2507,I1063026,I1063009,);
DFFARX1 I_62385 (I260748,I2507,I1063026,I1063100,);
not I_62386 (I1063108,I260730);
not I_62387 (I1063125,I260751);
nand I_62388 (I1063142,I1063125,I1063108);
nor I_62389 (I1062997,I1063100,I1063142);
DFFARX1 I_62390 (I1063142,I2507,I1063026,I1063182,);
not I_62391 (I1063018,I1063182);
not I_62392 (I1063204,I260754);
nand I_62393 (I1063221,I1063125,I1063204);
DFFARX1 I_62394 (I1063221,I2507,I1063026,I1063247,);
not I_62395 (I1063255,I1063247);
not I_62396 (I1063272,I260745);
nand I_62397 (I1063289,I1063272,I260733);
and I_62398 (I1063306,I1063108,I1063289);
nor I_62399 (I1063323,I1063221,I1063306);
DFFARX1 I_62400 (I1063323,I2507,I1063026,I1062994,);
DFFARX1 I_62401 (I1063306,I2507,I1063026,I1063015,);
nor I_62402 (I1063368,I260745,I260739);
nor I_62403 (I1063006,I1063221,I1063368);
or I_62404 (I1063399,I260745,I260739);
nor I_62405 (I1063416,I260736,I260730);
DFFARX1 I_62406 (I1063416,I2507,I1063026,I1063442,);
not I_62407 (I1063450,I1063442);
nor I_62408 (I1063012,I1063450,I1063255);
nand I_62409 (I1063481,I1063450,I1063100);
not I_62410 (I1063498,I260736);
nand I_62411 (I1063515,I1063498,I1063204);
nand I_62412 (I1063532,I1063450,I1063515);
nand I_62413 (I1063003,I1063532,I1063481);
nand I_62414 (I1063000,I1063515,I1063399);
not I_62415 (I1063604,I2514);
DFFARX1 I_62416 (I765985,I2507,I1063604,I1063630,);
and I_62417 (I1063638,I1063630,I765973);
DFFARX1 I_62418 (I1063638,I2507,I1063604,I1063587,);
DFFARX1 I_62419 (I765976,I2507,I1063604,I1063678,);
not I_62420 (I1063686,I765970);
not I_62421 (I1063703,I765994);
nand I_62422 (I1063720,I1063703,I1063686);
nor I_62423 (I1063575,I1063678,I1063720);
DFFARX1 I_62424 (I1063720,I2507,I1063604,I1063760,);
not I_62425 (I1063596,I1063760);
not I_62426 (I1063782,I765982);
nand I_62427 (I1063799,I1063703,I1063782);
DFFARX1 I_62428 (I1063799,I2507,I1063604,I1063825,);
not I_62429 (I1063833,I1063825);
not I_62430 (I1063850,I765991);
nand I_62431 (I1063867,I1063850,I765988);
and I_62432 (I1063884,I1063686,I1063867);
nor I_62433 (I1063901,I1063799,I1063884);
DFFARX1 I_62434 (I1063901,I2507,I1063604,I1063572,);
DFFARX1 I_62435 (I1063884,I2507,I1063604,I1063593,);
nor I_62436 (I1063946,I765991,I765979);
nor I_62437 (I1063584,I1063799,I1063946);
or I_62438 (I1063977,I765991,I765979);
nor I_62439 (I1063994,I765970,I765973);
DFFARX1 I_62440 (I1063994,I2507,I1063604,I1064020,);
not I_62441 (I1064028,I1064020);
nor I_62442 (I1063590,I1064028,I1063833);
nand I_62443 (I1064059,I1064028,I1063678);
not I_62444 (I1064076,I765970);
nand I_62445 (I1064093,I1064076,I1063782);
nand I_62446 (I1064110,I1064028,I1064093);
nand I_62447 (I1063581,I1064110,I1064059);
nand I_62448 (I1063578,I1064093,I1063977);
not I_62449 (I1064182,I2514);
DFFARX1 I_62450 (I265500,I2507,I1064182,I1064208,);
and I_62451 (I1064216,I1064208,I265485);
DFFARX1 I_62452 (I1064216,I2507,I1064182,I1064165,);
DFFARX1 I_62453 (I265491,I2507,I1064182,I1064256,);
not I_62454 (I1064264,I265473);
not I_62455 (I1064281,I265494);
nand I_62456 (I1064298,I1064281,I1064264);
nor I_62457 (I1064153,I1064256,I1064298);
DFFARX1 I_62458 (I1064298,I2507,I1064182,I1064338,);
not I_62459 (I1064174,I1064338);
not I_62460 (I1064360,I265497);
nand I_62461 (I1064377,I1064281,I1064360);
DFFARX1 I_62462 (I1064377,I2507,I1064182,I1064403,);
not I_62463 (I1064411,I1064403);
not I_62464 (I1064428,I265488);
nand I_62465 (I1064445,I1064428,I265476);
and I_62466 (I1064462,I1064264,I1064445);
nor I_62467 (I1064479,I1064377,I1064462);
DFFARX1 I_62468 (I1064479,I2507,I1064182,I1064150,);
DFFARX1 I_62469 (I1064462,I2507,I1064182,I1064171,);
nor I_62470 (I1064524,I265488,I265482);
nor I_62471 (I1064162,I1064377,I1064524);
or I_62472 (I1064555,I265488,I265482);
nor I_62473 (I1064572,I265479,I265473);
DFFARX1 I_62474 (I1064572,I2507,I1064182,I1064598,);
not I_62475 (I1064606,I1064598);
nor I_62476 (I1064168,I1064606,I1064411);
nand I_62477 (I1064637,I1064606,I1064256);
not I_62478 (I1064654,I265479);
nand I_62479 (I1064671,I1064654,I1064360);
nand I_62480 (I1064688,I1064606,I1064671);
nand I_62481 (I1064159,I1064688,I1064637);
nand I_62482 (I1064156,I1064671,I1064555);
not I_62483 (I1064760,I2514);
DFFARX1 I_62484 (I880247,I2507,I1064760,I1064786,);
and I_62485 (I1064794,I1064786,I880253);
DFFARX1 I_62486 (I1064794,I2507,I1064760,I1064743,);
DFFARX1 I_62487 (I880259,I2507,I1064760,I1064834,);
not I_62488 (I1064842,I880244);
not I_62489 (I1064859,I880244);
nand I_62490 (I1064876,I1064859,I1064842);
nor I_62491 (I1064731,I1064834,I1064876);
DFFARX1 I_62492 (I1064876,I2507,I1064760,I1064916,);
not I_62493 (I1064752,I1064916);
not I_62494 (I1064938,I880262);
nand I_62495 (I1064955,I1064859,I1064938);
DFFARX1 I_62496 (I1064955,I2507,I1064760,I1064981,);
not I_62497 (I1064989,I1064981);
not I_62498 (I1065006,I880256);
nand I_62499 (I1065023,I1065006,I880247);
and I_62500 (I1065040,I1064842,I1065023);
nor I_62501 (I1065057,I1064955,I1065040);
DFFARX1 I_62502 (I1065057,I2507,I1064760,I1064728,);
DFFARX1 I_62503 (I1065040,I2507,I1064760,I1064749,);
nor I_62504 (I1065102,I880256,I880265);
nor I_62505 (I1064740,I1064955,I1065102);
or I_62506 (I1065133,I880256,I880265);
nor I_62507 (I1065150,I880250,I880250);
DFFARX1 I_62508 (I1065150,I2507,I1064760,I1065176,);
not I_62509 (I1065184,I1065176);
nor I_62510 (I1064746,I1065184,I1064989);
nand I_62511 (I1065215,I1065184,I1064834);
not I_62512 (I1065232,I880250);
nand I_62513 (I1065249,I1065232,I1064938);
nand I_62514 (I1065266,I1065184,I1065249);
nand I_62515 (I1064737,I1065266,I1065215);
nand I_62516 (I1064734,I1065249,I1065133);
not I_62517 (I1065338,I2514);
DFFARX1 I_62518 (I418575,I2507,I1065338,I1065364,);
and I_62519 (I1065372,I1065364,I418590);
DFFARX1 I_62520 (I1065372,I2507,I1065338,I1065321,);
DFFARX1 I_62521 (I418593,I2507,I1065338,I1065412,);
not I_62522 (I1065420,I418587);
not I_62523 (I1065437,I418602);
nand I_62524 (I1065454,I1065437,I1065420);
nor I_62525 (I1065309,I1065412,I1065454);
DFFARX1 I_62526 (I1065454,I2507,I1065338,I1065494,);
not I_62527 (I1065330,I1065494);
not I_62528 (I1065516,I418578);
nand I_62529 (I1065533,I1065437,I1065516);
DFFARX1 I_62530 (I1065533,I2507,I1065338,I1065559,);
not I_62531 (I1065567,I1065559);
not I_62532 (I1065584,I418581);
nand I_62533 (I1065601,I1065584,I418575);
and I_62534 (I1065618,I1065420,I1065601);
nor I_62535 (I1065635,I1065533,I1065618);
DFFARX1 I_62536 (I1065635,I2507,I1065338,I1065306,);
DFFARX1 I_62537 (I1065618,I2507,I1065338,I1065327,);
nor I_62538 (I1065680,I418581,I418584);
nor I_62539 (I1065318,I1065533,I1065680);
or I_62540 (I1065711,I418581,I418584);
nor I_62541 (I1065728,I418599,I418596);
DFFARX1 I_62542 (I1065728,I2507,I1065338,I1065754,);
not I_62543 (I1065762,I1065754);
nor I_62544 (I1065324,I1065762,I1065567);
nand I_62545 (I1065793,I1065762,I1065412);
not I_62546 (I1065810,I418599);
nand I_62547 (I1065827,I1065810,I1065516);
nand I_62548 (I1065844,I1065762,I1065827);
nand I_62549 (I1065315,I1065844,I1065793);
nand I_62550 (I1065312,I1065827,I1065711);
not I_62551 (I1065916,I2514);
DFFARX1 I_62552 (I190690,I2507,I1065916,I1065942,);
and I_62553 (I1065950,I1065942,I190693);
DFFARX1 I_62554 (I1065950,I2507,I1065916,I1065899,);
DFFARX1 I_62555 (I190693,I2507,I1065916,I1065990,);
not I_62556 (I1065998,I190708);
not I_62557 (I1066015,I190714);
nand I_62558 (I1066032,I1066015,I1065998);
nor I_62559 (I1065887,I1065990,I1066032);
DFFARX1 I_62560 (I1066032,I2507,I1065916,I1066072,);
not I_62561 (I1065908,I1066072);
not I_62562 (I1066094,I190702);
nand I_62563 (I1066111,I1066015,I1066094);
DFFARX1 I_62564 (I1066111,I2507,I1065916,I1066137,);
not I_62565 (I1066145,I1066137);
not I_62566 (I1066162,I190699);
nand I_62567 (I1066179,I1066162,I190696);
and I_62568 (I1066196,I1065998,I1066179);
nor I_62569 (I1066213,I1066111,I1066196);
DFFARX1 I_62570 (I1066213,I2507,I1065916,I1065884,);
DFFARX1 I_62571 (I1066196,I2507,I1065916,I1065905,);
nor I_62572 (I1066258,I190699,I190690);
nor I_62573 (I1065896,I1066111,I1066258);
or I_62574 (I1066289,I190699,I190690);
nor I_62575 (I1066306,I190705,I190711);
DFFARX1 I_62576 (I1066306,I2507,I1065916,I1066332,);
not I_62577 (I1066340,I1066332);
nor I_62578 (I1065902,I1066340,I1066145);
nand I_62579 (I1066371,I1066340,I1065990);
not I_62580 (I1066388,I190705);
nand I_62581 (I1066405,I1066388,I1066094);
nand I_62582 (I1066422,I1066340,I1066405);
nand I_62583 (I1065893,I1066422,I1066371);
nand I_62584 (I1065890,I1066405,I1066289);
not I_62585 (I1066494,I2514);
DFFARX1 I_62586 (I802251,I2507,I1066494,I1066520,);
and I_62587 (I1066528,I1066520,I802257);
DFFARX1 I_62588 (I1066528,I2507,I1066494,I1066477,);
DFFARX1 I_62589 (I802263,I2507,I1066494,I1066568,);
not I_62590 (I1066576,I802248);
not I_62591 (I1066593,I802248);
nand I_62592 (I1066610,I1066593,I1066576);
nor I_62593 (I1066465,I1066568,I1066610);
DFFARX1 I_62594 (I1066610,I2507,I1066494,I1066650,);
not I_62595 (I1066486,I1066650);
not I_62596 (I1066672,I802266);
nand I_62597 (I1066689,I1066593,I1066672);
DFFARX1 I_62598 (I1066689,I2507,I1066494,I1066715,);
not I_62599 (I1066723,I1066715);
not I_62600 (I1066740,I802260);
nand I_62601 (I1066757,I1066740,I802251);
and I_62602 (I1066774,I1066576,I1066757);
nor I_62603 (I1066791,I1066689,I1066774);
DFFARX1 I_62604 (I1066791,I2507,I1066494,I1066462,);
DFFARX1 I_62605 (I1066774,I2507,I1066494,I1066483,);
nor I_62606 (I1066836,I802260,I802269);
nor I_62607 (I1066474,I1066689,I1066836);
or I_62608 (I1066867,I802260,I802269);
nor I_62609 (I1066884,I802254,I802254);
DFFARX1 I_62610 (I1066884,I2507,I1066494,I1066910,);
not I_62611 (I1066918,I1066910);
nor I_62612 (I1066480,I1066918,I1066723);
nand I_62613 (I1066949,I1066918,I1066568);
not I_62614 (I1066966,I802254);
nand I_62615 (I1066983,I1066966,I1066672);
nand I_62616 (I1067000,I1066918,I1066983);
nand I_62617 (I1066471,I1067000,I1066949);
nand I_62618 (I1066468,I1066983,I1066867);
not I_62619 (I1067072,I2514);
DFFARX1 I_62620 (I207945,I2507,I1067072,I1067098,);
and I_62621 (I1067106,I1067098,I207948);
DFFARX1 I_62622 (I1067106,I2507,I1067072,I1067055,);
DFFARX1 I_62623 (I207948,I2507,I1067072,I1067146,);
not I_62624 (I1067154,I207963);
not I_62625 (I1067171,I207969);
nand I_62626 (I1067188,I1067171,I1067154);
nor I_62627 (I1067043,I1067146,I1067188);
DFFARX1 I_62628 (I1067188,I2507,I1067072,I1067228,);
not I_62629 (I1067064,I1067228);
not I_62630 (I1067250,I207957);
nand I_62631 (I1067267,I1067171,I1067250);
DFFARX1 I_62632 (I1067267,I2507,I1067072,I1067293,);
not I_62633 (I1067301,I1067293);
not I_62634 (I1067318,I207954);
nand I_62635 (I1067335,I1067318,I207951);
and I_62636 (I1067352,I1067154,I1067335);
nor I_62637 (I1067369,I1067267,I1067352);
DFFARX1 I_62638 (I1067369,I2507,I1067072,I1067040,);
DFFARX1 I_62639 (I1067352,I2507,I1067072,I1067061,);
nor I_62640 (I1067414,I207954,I207945);
nor I_62641 (I1067052,I1067267,I1067414);
or I_62642 (I1067445,I207954,I207945);
nor I_62643 (I1067462,I207960,I207966);
DFFARX1 I_62644 (I1067462,I2507,I1067072,I1067488,);
not I_62645 (I1067496,I1067488);
nor I_62646 (I1067058,I1067496,I1067301);
nand I_62647 (I1067527,I1067496,I1067146);
not I_62648 (I1067544,I207960);
nand I_62649 (I1067561,I1067544,I1067250);
nand I_62650 (I1067578,I1067496,I1067561);
nand I_62651 (I1067049,I1067578,I1067527);
nand I_62652 (I1067046,I1067561,I1067445);
not I_62653 (I1067650,I2514);
DFFARX1 I_62654 (I408239,I2507,I1067650,I1067676,);
and I_62655 (I1067684,I1067676,I408254);
DFFARX1 I_62656 (I1067684,I2507,I1067650,I1067633,);
DFFARX1 I_62657 (I408257,I2507,I1067650,I1067724,);
not I_62658 (I1067732,I408251);
not I_62659 (I1067749,I408266);
nand I_62660 (I1067766,I1067749,I1067732);
nor I_62661 (I1067621,I1067724,I1067766);
DFFARX1 I_62662 (I1067766,I2507,I1067650,I1067806,);
not I_62663 (I1067642,I1067806);
not I_62664 (I1067828,I408242);
nand I_62665 (I1067845,I1067749,I1067828);
DFFARX1 I_62666 (I1067845,I2507,I1067650,I1067871,);
not I_62667 (I1067879,I1067871);
not I_62668 (I1067896,I408245);
nand I_62669 (I1067913,I1067896,I408239);
and I_62670 (I1067930,I1067732,I1067913);
nor I_62671 (I1067947,I1067845,I1067930);
DFFARX1 I_62672 (I1067947,I2507,I1067650,I1067618,);
DFFARX1 I_62673 (I1067930,I2507,I1067650,I1067639,);
nor I_62674 (I1067992,I408245,I408248);
nor I_62675 (I1067630,I1067845,I1067992);
or I_62676 (I1068023,I408245,I408248);
nor I_62677 (I1068040,I408263,I408260);
DFFARX1 I_62678 (I1068040,I2507,I1067650,I1068066,);
not I_62679 (I1068074,I1068066);
nor I_62680 (I1067636,I1068074,I1067879);
nand I_62681 (I1068105,I1068074,I1067724);
not I_62682 (I1068122,I408263);
nand I_62683 (I1068139,I1068122,I1067828);
nand I_62684 (I1068156,I1068074,I1068139);
nand I_62685 (I1067627,I1068156,I1068105);
nand I_62686 (I1067624,I1068139,I1068023);
not I_62687 (I1068228,I2514);
DFFARX1 I_62688 (I712809,I2507,I1068228,I1068254,);
and I_62689 (I1068262,I1068254,I712797);
DFFARX1 I_62690 (I1068262,I2507,I1068228,I1068211,);
DFFARX1 I_62691 (I712800,I2507,I1068228,I1068302,);
not I_62692 (I1068310,I712794);
not I_62693 (I1068327,I712818);
nand I_62694 (I1068344,I1068327,I1068310);
nor I_62695 (I1068199,I1068302,I1068344);
DFFARX1 I_62696 (I1068344,I2507,I1068228,I1068384,);
not I_62697 (I1068220,I1068384);
not I_62698 (I1068406,I712806);
nand I_62699 (I1068423,I1068327,I1068406);
DFFARX1 I_62700 (I1068423,I2507,I1068228,I1068449,);
not I_62701 (I1068457,I1068449);
not I_62702 (I1068474,I712815);
nand I_62703 (I1068491,I1068474,I712812);
and I_62704 (I1068508,I1068310,I1068491);
nor I_62705 (I1068525,I1068423,I1068508);
DFFARX1 I_62706 (I1068525,I2507,I1068228,I1068196,);
DFFARX1 I_62707 (I1068508,I2507,I1068228,I1068217,);
nor I_62708 (I1068570,I712815,I712803);
nor I_62709 (I1068208,I1068423,I1068570);
or I_62710 (I1068601,I712815,I712803);
nor I_62711 (I1068618,I712794,I712797);
DFFARX1 I_62712 (I1068618,I2507,I1068228,I1068644,);
not I_62713 (I1068652,I1068644);
nor I_62714 (I1068214,I1068652,I1068457);
nand I_62715 (I1068683,I1068652,I1068302);
not I_62716 (I1068700,I712794);
nand I_62717 (I1068717,I1068700,I1068406);
nand I_62718 (I1068734,I1068652,I1068717);
nand I_62719 (I1068205,I1068734,I1068683);
nand I_62720 (I1068202,I1068717,I1068601);
not I_62721 (I1068806,I2514);
DFFARX1 I_62722 (I356144,I2507,I1068806,I1068832,);
and I_62723 (I1068840,I1068832,I356129);
DFFARX1 I_62724 (I1068840,I2507,I1068806,I1068789,);
DFFARX1 I_62725 (I356135,I2507,I1068806,I1068880,);
not I_62726 (I1068888,I356117);
not I_62727 (I1068905,I356138);
nand I_62728 (I1068922,I1068905,I1068888);
nor I_62729 (I1068777,I1068880,I1068922);
DFFARX1 I_62730 (I1068922,I2507,I1068806,I1068962,);
not I_62731 (I1068798,I1068962);
not I_62732 (I1068984,I356141);
nand I_62733 (I1069001,I1068905,I1068984);
DFFARX1 I_62734 (I1069001,I2507,I1068806,I1069027,);
not I_62735 (I1069035,I1069027);
not I_62736 (I1069052,I356132);
nand I_62737 (I1069069,I1069052,I356120);
and I_62738 (I1069086,I1068888,I1069069);
nor I_62739 (I1069103,I1069001,I1069086);
DFFARX1 I_62740 (I1069103,I2507,I1068806,I1068774,);
DFFARX1 I_62741 (I1069086,I2507,I1068806,I1068795,);
nor I_62742 (I1069148,I356132,I356126);
nor I_62743 (I1068786,I1069001,I1069148);
or I_62744 (I1069179,I356132,I356126);
nor I_62745 (I1069196,I356123,I356117);
DFFARX1 I_62746 (I1069196,I2507,I1068806,I1069222,);
not I_62747 (I1069230,I1069222);
nor I_62748 (I1068792,I1069230,I1069035);
nand I_62749 (I1069261,I1069230,I1068880);
not I_62750 (I1069278,I356123);
nand I_62751 (I1069295,I1069278,I1068984);
nand I_62752 (I1069312,I1069230,I1069295);
nand I_62753 (I1068783,I1069312,I1069261);
nand I_62754 (I1068780,I1069295,I1069179);
not I_62755 (I1069384,I2514);
DFFARX1 I_62756 (I346658,I2507,I1069384,I1069410,);
and I_62757 (I1069418,I1069410,I346643);
DFFARX1 I_62758 (I1069418,I2507,I1069384,I1069367,);
DFFARX1 I_62759 (I346649,I2507,I1069384,I1069458,);
not I_62760 (I1069466,I346631);
not I_62761 (I1069483,I346652);
nand I_62762 (I1069500,I1069483,I1069466);
nor I_62763 (I1069355,I1069458,I1069500);
DFFARX1 I_62764 (I1069500,I2507,I1069384,I1069540,);
not I_62765 (I1069376,I1069540);
not I_62766 (I1069562,I346655);
nand I_62767 (I1069579,I1069483,I1069562);
DFFARX1 I_62768 (I1069579,I2507,I1069384,I1069605,);
not I_62769 (I1069613,I1069605);
not I_62770 (I1069630,I346646);
nand I_62771 (I1069647,I1069630,I346634);
and I_62772 (I1069664,I1069466,I1069647);
nor I_62773 (I1069681,I1069579,I1069664);
DFFARX1 I_62774 (I1069681,I2507,I1069384,I1069352,);
DFFARX1 I_62775 (I1069664,I2507,I1069384,I1069373,);
nor I_62776 (I1069726,I346646,I346640);
nor I_62777 (I1069364,I1069579,I1069726);
or I_62778 (I1069757,I346646,I346640);
nor I_62779 (I1069774,I346637,I346631);
DFFARX1 I_62780 (I1069774,I2507,I1069384,I1069800,);
not I_62781 (I1069808,I1069800);
nor I_62782 (I1069370,I1069808,I1069613);
nand I_62783 (I1069839,I1069808,I1069458);
not I_62784 (I1069856,I346637);
nand I_62785 (I1069873,I1069856,I1069562);
nand I_62786 (I1069890,I1069808,I1069873);
nand I_62787 (I1069361,I1069890,I1069839);
nand I_62788 (I1069358,I1069873,I1069757);
not I_62789 (I1069962,I2514);
DFFARX1 I_62790 (I1228119,I2507,I1069962,I1069988,);
and I_62791 (I1069996,I1069988,I1228113);
DFFARX1 I_62792 (I1069996,I2507,I1069962,I1069945,);
DFFARX1 I_62793 (I1228098,I2507,I1069962,I1070036,);
not I_62794 (I1070044,I1228104);
not I_62795 (I1070061,I1228116);
nand I_62796 (I1070078,I1070061,I1070044);
nor I_62797 (I1069933,I1070036,I1070078);
DFFARX1 I_62798 (I1070078,I2507,I1069962,I1070118,);
not I_62799 (I1069954,I1070118);
not I_62800 (I1070140,I1228098);
nand I_62801 (I1070157,I1070061,I1070140);
DFFARX1 I_62802 (I1070157,I2507,I1069962,I1070183,);
not I_62803 (I1070191,I1070183);
not I_62804 (I1070208,I1228122);
nand I_62805 (I1070225,I1070208,I1228110);
and I_62806 (I1070242,I1070044,I1070225);
nor I_62807 (I1070259,I1070157,I1070242);
DFFARX1 I_62808 (I1070259,I2507,I1069962,I1069930,);
DFFARX1 I_62809 (I1070242,I2507,I1069962,I1069951,);
nor I_62810 (I1070304,I1228122,I1228101);
nor I_62811 (I1069942,I1070157,I1070304);
or I_62812 (I1070335,I1228122,I1228101);
nor I_62813 (I1070352,I1228107,I1228101);
DFFARX1 I_62814 (I1070352,I2507,I1069962,I1070378,);
not I_62815 (I1070386,I1070378);
nor I_62816 (I1069948,I1070386,I1070191);
nand I_62817 (I1070417,I1070386,I1070036);
not I_62818 (I1070434,I1228107);
nand I_62819 (I1070451,I1070434,I1070140);
nand I_62820 (I1070468,I1070386,I1070451);
nand I_62821 (I1069939,I1070468,I1070417);
nand I_62822 (I1069936,I1070451,I1070335);
not I_62823 (I1070540,I2514);
DFFARX1 I_62824 (I828601,I2507,I1070540,I1070566,);
and I_62825 (I1070574,I1070566,I828607);
DFFARX1 I_62826 (I1070574,I2507,I1070540,I1070523,);
DFFARX1 I_62827 (I828613,I2507,I1070540,I1070614,);
not I_62828 (I1070622,I828598);
not I_62829 (I1070639,I828598);
nand I_62830 (I1070656,I1070639,I1070622);
nor I_62831 (I1070511,I1070614,I1070656);
DFFARX1 I_62832 (I1070656,I2507,I1070540,I1070696,);
not I_62833 (I1070532,I1070696);
not I_62834 (I1070718,I828616);
nand I_62835 (I1070735,I1070639,I1070718);
DFFARX1 I_62836 (I1070735,I2507,I1070540,I1070761,);
not I_62837 (I1070769,I1070761);
not I_62838 (I1070786,I828610);
nand I_62839 (I1070803,I1070786,I828601);
and I_62840 (I1070820,I1070622,I1070803);
nor I_62841 (I1070837,I1070735,I1070820);
DFFARX1 I_62842 (I1070837,I2507,I1070540,I1070508,);
DFFARX1 I_62843 (I1070820,I2507,I1070540,I1070529,);
nor I_62844 (I1070882,I828610,I828619);
nor I_62845 (I1070520,I1070735,I1070882);
or I_62846 (I1070913,I828610,I828619);
nor I_62847 (I1070930,I828604,I828604);
DFFARX1 I_62848 (I1070930,I2507,I1070540,I1070956,);
not I_62849 (I1070964,I1070956);
nor I_62850 (I1070526,I1070964,I1070769);
nand I_62851 (I1070995,I1070964,I1070614);
not I_62852 (I1071012,I828604);
nand I_62853 (I1071029,I1071012,I1070718);
nand I_62854 (I1071046,I1070964,I1071029);
nand I_62855 (I1070517,I1071046,I1070995);
nand I_62856 (I1070514,I1071029,I1070913);
not I_62857 (I1071118,I2514);
DFFARX1 I_62858 (I1329139,I2507,I1071118,I1071144,);
and I_62859 (I1071152,I1071144,I1329121);
DFFARX1 I_62860 (I1071152,I2507,I1071118,I1071101,);
DFFARX1 I_62861 (I1329112,I2507,I1071118,I1071192,);
not I_62862 (I1071200,I1329127);
not I_62863 (I1071217,I1329115);
nand I_62864 (I1071234,I1071217,I1071200);
nor I_62865 (I1071089,I1071192,I1071234);
DFFARX1 I_62866 (I1071234,I2507,I1071118,I1071274,);
not I_62867 (I1071110,I1071274);
not I_62868 (I1071296,I1329124);
nand I_62869 (I1071313,I1071217,I1071296);
DFFARX1 I_62870 (I1071313,I2507,I1071118,I1071339,);
not I_62871 (I1071347,I1071339);
not I_62872 (I1071364,I1329133);
nand I_62873 (I1071381,I1071364,I1329112);
and I_62874 (I1071398,I1071200,I1071381);
nor I_62875 (I1071415,I1071313,I1071398);
DFFARX1 I_62876 (I1071415,I2507,I1071118,I1071086,);
DFFARX1 I_62877 (I1071398,I2507,I1071118,I1071107,);
nor I_62878 (I1071460,I1329133,I1329136);
nor I_62879 (I1071098,I1071313,I1071460);
or I_62880 (I1071491,I1329133,I1329136);
nor I_62881 (I1071508,I1329130,I1329118);
DFFARX1 I_62882 (I1071508,I2507,I1071118,I1071534,);
not I_62883 (I1071542,I1071534);
nor I_62884 (I1071104,I1071542,I1071347);
nand I_62885 (I1071573,I1071542,I1071192);
not I_62886 (I1071590,I1329130);
nand I_62887 (I1071607,I1071590,I1071296);
nand I_62888 (I1071624,I1071542,I1071607);
nand I_62889 (I1071095,I1071624,I1071573);
nand I_62890 (I1071092,I1071607,I1071491);
not I_62891 (I1071696,I2514);
DFFARX1 I_62892 (I703561,I2507,I1071696,I1071722,);
and I_62893 (I1071730,I1071722,I703549);
DFFARX1 I_62894 (I1071730,I2507,I1071696,I1071679,);
DFFARX1 I_62895 (I703552,I2507,I1071696,I1071770,);
not I_62896 (I1071778,I703546);
not I_62897 (I1071795,I703570);
nand I_62898 (I1071812,I1071795,I1071778);
nor I_62899 (I1071667,I1071770,I1071812);
DFFARX1 I_62900 (I1071812,I2507,I1071696,I1071852,);
not I_62901 (I1071688,I1071852);
not I_62902 (I1071874,I703558);
nand I_62903 (I1071891,I1071795,I1071874);
DFFARX1 I_62904 (I1071891,I2507,I1071696,I1071917,);
not I_62905 (I1071925,I1071917);
not I_62906 (I1071942,I703567);
nand I_62907 (I1071959,I1071942,I703564);
and I_62908 (I1071976,I1071778,I1071959);
nor I_62909 (I1071993,I1071891,I1071976);
DFFARX1 I_62910 (I1071993,I2507,I1071696,I1071664,);
DFFARX1 I_62911 (I1071976,I2507,I1071696,I1071685,);
nor I_62912 (I1072038,I703567,I703555);
nor I_62913 (I1071676,I1071891,I1072038);
or I_62914 (I1072069,I703567,I703555);
nor I_62915 (I1072086,I703546,I703549);
DFFARX1 I_62916 (I1072086,I2507,I1071696,I1072112,);
not I_62917 (I1072120,I1072112);
nor I_62918 (I1071682,I1072120,I1071925);
nand I_62919 (I1072151,I1072120,I1071770);
not I_62920 (I1072168,I703546);
nand I_62921 (I1072185,I1072168,I1071874);
nand I_62922 (I1072202,I1072120,I1072185);
nand I_62923 (I1071673,I1072202,I1072151);
nand I_62924 (I1071670,I1072185,I1072069);
not I_62925 (I1072274,I2514);
DFFARX1 I_62926 (I141900,I2507,I1072274,I1072300,);
and I_62927 (I1072308,I1072300,I141924);
DFFARX1 I_62928 (I1072308,I2507,I1072274,I1072257,);
DFFARX1 I_62929 (I141900,I2507,I1072274,I1072348,);
not I_62930 (I1072356,I141918);
not I_62931 (I1072373,I141903);
nand I_62932 (I1072390,I1072373,I1072356);
nor I_62933 (I1072245,I1072348,I1072390);
DFFARX1 I_62934 (I1072390,I2507,I1072274,I1072430,);
not I_62935 (I1072266,I1072430);
not I_62936 (I1072452,I141912);
nand I_62937 (I1072469,I1072373,I1072452);
DFFARX1 I_62938 (I1072469,I2507,I1072274,I1072495,);
not I_62939 (I1072503,I1072495);
not I_62940 (I1072520,I141909);
nand I_62941 (I1072537,I1072520,I141906);
and I_62942 (I1072554,I1072356,I1072537);
nor I_62943 (I1072571,I1072469,I1072554);
DFFARX1 I_62944 (I1072571,I2507,I1072274,I1072242,);
DFFARX1 I_62945 (I1072554,I2507,I1072274,I1072263,);
nor I_62946 (I1072616,I141909,I141915);
nor I_62947 (I1072254,I1072469,I1072616);
or I_62948 (I1072647,I141909,I141915);
nor I_62949 (I1072664,I141921,I141927);
DFFARX1 I_62950 (I1072664,I2507,I1072274,I1072690,);
not I_62951 (I1072698,I1072690);
nor I_62952 (I1072260,I1072698,I1072503);
nand I_62953 (I1072729,I1072698,I1072348);
not I_62954 (I1072746,I141921);
nand I_62955 (I1072763,I1072746,I1072452);
nand I_62956 (I1072780,I1072698,I1072763);
nand I_62957 (I1072251,I1072780,I1072729);
nand I_62958 (I1072248,I1072763,I1072647);
not I_62959 (I1072852,I2514);
DFFARX1 I_62960 (I1256512,I2507,I1072852,I1072878,);
and I_62961 (I1072886,I1072878,I1256494);
DFFARX1 I_62962 (I1072886,I2507,I1072852,I1072835,);
DFFARX1 I_62963 (I1256503,I2507,I1072852,I1072926,);
not I_62964 (I1072934,I1256488);
not I_62965 (I1072951,I1256500);
nand I_62966 (I1072968,I1072951,I1072934);
nor I_62967 (I1072823,I1072926,I1072968);
DFFARX1 I_62968 (I1072968,I2507,I1072852,I1073008,);
not I_62969 (I1072844,I1073008);
not I_62970 (I1073030,I1256491);
nand I_62971 (I1073047,I1072951,I1073030);
DFFARX1 I_62972 (I1073047,I2507,I1072852,I1073073,);
not I_62973 (I1073081,I1073073);
not I_62974 (I1073098,I1256488);
nand I_62975 (I1073115,I1073098,I1256491);
and I_62976 (I1073132,I1072934,I1073115);
nor I_62977 (I1073149,I1073047,I1073132);
DFFARX1 I_62978 (I1073149,I2507,I1072852,I1072820,);
DFFARX1 I_62979 (I1073132,I2507,I1072852,I1072841,);
nor I_62980 (I1073194,I1256488,I1256509);
nor I_62981 (I1072832,I1073047,I1073194);
or I_62982 (I1073225,I1256488,I1256509);
nor I_62983 (I1073242,I1256497,I1256506);
DFFARX1 I_62984 (I1073242,I2507,I1072852,I1073268,);
not I_62985 (I1073276,I1073268);
nor I_62986 (I1072838,I1073276,I1073081);
nand I_62987 (I1073307,I1073276,I1072926);
not I_62988 (I1073324,I1256497);
nand I_62989 (I1073341,I1073324,I1073030);
nand I_62990 (I1073358,I1073276,I1073341);
nand I_62991 (I1072829,I1073358,I1073307);
nand I_62992 (I1072826,I1073341,I1073225);
not I_62993 (I1073430,I2514);
DFFARX1 I_62994 (I848100,I2507,I1073430,I1073456,);
and I_62995 (I1073464,I1073456,I848106);
DFFARX1 I_62996 (I1073464,I2507,I1073430,I1073413,);
DFFARX1 I_62997 (I848112,I2507,I1073430,I1073504,);
not I_62998 (I1073512,I848097);
not I_62999 (I1073529,I848097);
nand I_63000 (I1073546,I1073529,I1073512);
nor I_63001 (I1073401,I1073504,I1073546);
DFFARX1 I_63002 (I1073546,I2507,I1073430,I1073586,);
not I_63003 (I1073422,I1073586);
not I_63004 (I1073608,I848115);
nand I_63005 (I1073625,I1073529,I1073608);
DFFARX1 I_63006 (I1073625,I2507,I1073430,I1073651,);
not I_63007 (I1073659,I1073651);
not I_63008 (I1073676,I848109);
nand I_63009 (I1073693,I1073676,I848100);
and I_63010 (I1073710,I1073512,I1073693);
nor I_63011 (I1073727,I1073625,I1073710);
DFFARX1 I_63012 (I1073727,I2507,I1073430,I1073398,);
DFFARX1 I_63013 (I1073710,I2507,I1073430,I1073419,);
nor I_63014 (I1073772,I848109,I848118);
nor I_63015 (I1073410,I1073625,I1073772);
or I_63016 (I1073803,I848109,I848118);
nor I_63017 (I1073820,I848103,I848103);
DFFARX1 I_63018 (I1073820,I2507,I1073430,I1073846,);
not I_63019 (I1073854,I1073846);
nor I_63020 (I1073416,I1073854,I1073659);
nand I_63021 (I1073885,I1073854,I1073504);
not I_63022 (I1073902,I848103);
nand I_63023 (I1073919,I1073902,I1073608);
nand I_63024 (I1073936,I1073854,I1073919);
nand I_63025 (I1073407,I1073936,I1073885);
nand I_63026 (I1073404,I1073919,I1073803);
not I_63027 (I1074008,I2514);
DFFARX1 I_63028 (I1040438,I2507,I1074008,I1074034,);
and I_63029 (I1074042,I1074034,I1040435);
DFFARX1 I_63030 (I1074042,I2507,I1074008,I1073991,);
DFFARX1 I_63031 (I1040441,I2507,I1074008,I1074082,);
not I_63032 (I1074090,I1040444);
not I_63033 (I1074107,I1040438);
nand I_63034 (I1074124,I1074107,I1074090);
nor I_63035 (I1073979,I1074082,I1074124);
DFFARX1 I_63036 (I1074124,I2507,I1074008,I1074164,);
not I_63037 (I1074000,I1074164);
not I_63038 (I1074186,I1040453);
nand I_63039 (I1074203,I1074107,I1074186);
DFFARX1 I_63040 (I1074203,I2507,I1074008,I1074229,);
not I_63041 (I1074237,I1074229);
not I_63042 (I1074254,I1040450);
nand I_63043 (I1074271,I1074254,I1040456);
and I_63044 (I1074288,I1074090,I1074271);
nor I_63045 (I1074305,I1074203,I1074288);
DFFARX1 I_63046 (I1074305,I2507,I1074008,I1073976,);
DFFARX1 I_63047 (I1074288,I2507,I1074008,I1073997,);
nor I_63048 (I1074350,I1040450,I1040435);
nor I_63049 (I1073988,I1074203,I1074350);
or I_63050 (I1074381,I1040450,I1040435);
nor I_63051 (I1074398,I1040447,I1040441);
DFFARX1 I_63052 (I1074398,I2507,I1074008,I1074424,);
not I_63053 (I1074432,I1074424);
nor I_63054 (I1073994,I1074432,I1074237);
nand I_63055 (I1074463,I1074432,I1074082);
not I_63056 (I1074480,I1040447);
nand I_63057 (I1074497,I1074480,I1074186);
nand I_63058 (I1074514,I1074432,I1074497);
nand I_63059 (I1073985,I1074514,I1074463);
nand I_63060 (I1073982,I1074497,I1074381);
not I_63061 (I1074586,I2514);
DFFARX1 I_63062 (I440335,I2507,I1074586,I1074612,);
and I_63063 (I1074620,I1074612,I440350);
DFFARX1 I_63064 (I1074620,I2507,I1074586,I1074569,);
DFFARX1 I_63065 (I440353,I2507,I1074586,I1074660,);
not I_63066 (I1074668,I440347);
not I_63067 (I1074685,I440362);
nand I_63068 (I1074702,I1074685,I1074668);
nor I_63069 (I1074557,I1074660,I1074702);
DFFARX1 I_63070 (I1074702,I2507,I1074586,I1074742,);
not I_63071 (I1074578,I1074742);
not I_63072 (I1074764,I440338);
nand I_63073 (I1074781,I1074685,I1074764);
DFFARX1 I_63074 (I1074781,I2507,I1074586,I1074807,);
not I_63075 (I1074815,I1074807);
not I_63076 (I1074832,I440341);
nand I_63077 (I1074849,I1074832,I440335);
and I_63078 (I1074866,I1074668,I1074849);
nor I_63079 (I1074883,I1074781,I1074866);
DFFARX1 I_63080 (I1074883,I2507,I1074586,I1074554,);
DFFARX1 I_63081 (I1074866,I2507,I1074586,I1074575,);
nor I_63082 (I1074928,I440341,I440344);
nor I_63083 (I1074566,I1074781,I1074928);
or I_63084 (I1074959,I440341,I440344);
nor I_63085 (I1074976,I440359,I440356);
DFFARX1 I_63086 (I1074976,I2507,I1074586,I1075002,);
not I_63087 (I1075010,I1075002);
nor I_63088 (I1074572,I1075010,I1074815);
nand I_63089 (I1075041,I1075010,I1074660);
not I_63090 (I1075058,I440359);
nand I_63091 (I1075075,I1075058,I1074764);
nand I_63092 (I1075092,I1075010,I1075075);
nand I_63093 (I1074563,I1075092,I1075041);
nand I_63094 (I1074560,I1075075,I1074959);
not I_63095 (I1075164,I2514);
DFFARX1 I_63096 (I952823,I2507,I1075164,I1075190,);
and I_63097 (I1075198,I1075190,I952817);
DFFARX1 I_63098 (I1075198,I2507,I1075164,I1075147,);
DFFARX1 I_63099 (I952835,I2507,I1075164,I1075238,);
not I_63100 (I1075246,I952826);
not I_63101 (I1075263,I952838);
nand I_63102 (I1075280,I1075263,I1075246);
nor I_63103 (I1075135,I1075238,I1075280);
DFFARX1 I_63104 (I1075280,I2507,I1075164,I1075320,);
not I_63105 (I1075156,I1075320);
not I_63106 (I1075342,I952844);
nand I_63107 (I1075359,I1075263,I1075342);
DFFARX1 I_63108 (I1075359,I2507,I1075164,I1075385,);
not I_63109 (I1075393,I1075385);
not I_63110 (I1075410,I952820);
nand I_63111 (I1075427,I1075410,I952841);
and I_63112 (I1075444,I1075246,I1075427);
nor I_63113 (I1075461,I1075359,I1075444);
DFFARX1 I_63114 (I1075461,I2507,I1075164,I1075132,);
DFFARX1 I_63115 (I1075444,I2507,I1075164,I1075153,);
nor I_63116 (I1075506,I952820,I952832);
nor I_63117 (I1075144,I1075359,I1075506);
or I_63118 (I1075537,I952820,I952832);
nor I_63119 (I1075554,I952817,I952829);
DFFARX1 I_63120 (I1075554,I2507,I1075164,I1075580,);
not I_63121 (I1075588,I1075580);
nor I_63122 (I1075150,I1075588,I1075393);
nand I_63123 (I1075619,I1075588,I1075238);
not I_63124 (I1075636,I952817);
nand I_63125 (I1075653,I1075636,I1075342);
nand I_63126 (I1075670,I1075588,I1075653);
nand I_63127 (I1075141,I1075670,I1075619);
nand I_63128 (I1075138,I1075653,I1075537);
not I_63129 (I1075742,I2514);
DFFARX1 I_63130 (I1379714,I2507,I1075742,I1075768,);
and I_63131 (I1075776,I1075768,I1379696);
DFFARX1 I_63132 (I1075776,I2507,I1075742,I1075725,);
DFFARX1 I_63133 (I1379687,I2507,I1075742,I1075816,);
not I_63134 (I1075824,I1379702);
not I_63135 (I1075841,I1379690);
nand I_63136 (I1075858,I1075841,I1075824);
nor I_63137 (I1075713,I1075816,I1075858);
DFFARX1 I_63138 (I1075858,I2507,I1075742,I1075898,);
not I_63139 (I1075734,I1075898);
not I_63140 (I1075920,I1379699);
nand I_63141 (I1075937,I1075841,I1075920);
DFFARX1 I_63142 (I1075937,I2507,I1075742,I1075963,);
not I_63143 (I1075971,I1075963);
not I_63144 (I1075988,I1379708);
nand I_63145 (I1076005,I1075988,I1379687);
and I_63146 (I1076022,I1075824,I1076005);
nor I_63147 (I1076039,I1075937,I1076022);
DFFARX1 I_63148 (I1076039,I2507,I1075742,I1075710,);
DFFARX1 I_63149 (I1076022,I2507,I1075742,I1075731,);
nor I_63150 (I1076084,I1379708,I1379711);
nor I_63151 (I1075722,I1075937,I1076084);
or I_63152 (I1076115,I1379708,I1379711);
nor I_63153 (I1076132,I1379705,I1379693);
DFFARX1 I_63154 (I1076132,I2507,I1075742,I1076158,);
not I_63155 (I1076166,I1076158);
nor I_63156 (I1075728,I1076166,I1075971);
nand I_63157 (I1076197,I1076166,I1075816);
not I_63158 (I1076214,I1379705);
nand I_63159 (I1076231,I1076214,I1075920);
nand I_63160 (I1076248,I1076166,I1076231);
nand I_63161 (I1075719,I1076248,I1076197);
nand I_63162 (I1075716,I1076231,I1076115);
not I_63163 (I1076320,I2514);
DFFARX1 I_63164 (I750957,I2507,I1076320,I1076346,);
and I_63165 (I1076354,I1076346,I750945);
DFFARX1 I_63166 (I1076354,I2507,I1076320,I1076303,);
DFFARX1 I_63167 (I750948,I2507,I1076320,I1076394,);
not I_63168 (I1076402,I750942);
not I_63169 (I1076419,I750966);
nand I_63170 (I1076436,I1076419,I1076402);
nor I_63171 (I1076291,I1076394,I1076436);
DFFARX1 I_63172 (I1076436,I2507,I1076320,I1076476,);
not I_63173 (I1076312,I1076476);
not I_63174 (I1076498,I750954);
nand I_63175 (I1076515,I1076419,I1076498);
DFFARX1 I_63176 (I1076515,I2507,I1076320,I1076541,);
not I_63177 (I1076549,I1076541);
not I_63178 (I1076566,I750963);
nand I_63179 (I1076583,I1076566,I750960);
and I_63180 (I1076600,I1076402,I1076583);
nor I_63181 (I1076617,I1076515,I1076600);
DFFARX1 I_63182 (I1076617,I2507,I1076320,I1076288,);
DFFARX1 I_63183 (I1076600,I2507,I1076320,I1076309,);
nor I_63184 (I1076662,I750963,I750951);
nor I_63185 (I1076300,I1076515,I1076662);
or I_63186 (I1076693,I750963,I750951);
nor I_63187 (I1076710,I750942,I750945);
DFFARX1 I_63188 (I1076710,I2507,I1076320,I1076736,);
not I_63189 (I1076744,I1076736);
nor I_63190 (I1076306,I1076744,I1076549);
nand I_63191 (I1076775,I1076744,I1076394);
not I_63192 (I1076792,I750942);
nand I_63193 (I1076809,I1076792,I1076498);
nand I_63194 (I1076826,I1076744,I1076809);
nand I_63195 (I1076297,I1076826,I1076775);
nand I_63196 (I1076294,I1076809,I1076693);
not I_63197 (I1076898,I2514);
DFFARX1 I_63198 (I945071,I2507,I1076898,I1076924,);
and I_63199 (I1076932,I1076924,I945065);
DFFARX1 I_63200 (I1076932,I2507,I1076898,I1076881,);
DFFARX1 I_63201 (I945083,I2507,I1076898,I1076972,);
not I_63202 (I1076980,I945074);
not I_63203 (I1076997,I945086);
nand I_63204 (I1077014,I1076997,I1076980);
nor I_63205 (I1076869,I1076972,I1077014);
DFFARX1 I_63206 (I1077014,I2507,I1076898,I1077054,);
not I_63207 (I1076890,I1077054);
not I_63208 (I1077076,I945092);
nand I_63209 (I1077093,I1076997,I1077076);
DFFARX1 I_63210 (I1077093,I2507,I1076898,I1077119,);
not I_63211 (I1077127,I1077119);
not I_63212 (I1077144,I945068);
nand I_63213 (I1077161,I1077144,I945089);
and I_63214 (I1077178,I1076980,I1077161);
nor I_63215 (I1077195,I1077093,I1077178);
DFFARX1 I_63216 (I1077195,I2507,I1076898,I1076866,);
DFFARX1 I_63217 (I1077178,I2507,I1076898,I1076887,);
nor I_63218 (I1077240,I945068,I945080);
nor I_63219 (I1076878,I1077093,I1077240);
or I_63220 (I1077271,I945068,I945080);
nor I_63221 (I1077288,I945065,I945077);
DFFARX1 I_63222 (I1077288,I2507,I1076898,I1077314,);
not I_63223 (I1077322,I1077314);
nor I_63224 (I1076884,I1077322,I1077127);
nand I_63225 (I1077353,I1077322,I1076972);
not I_63226 (I1077370,I945065);
nand I_63227 (I1077387,I1077370,I1077076);
nand I_63228 (I1077404,I1077322,I1077387);
nand I_63229 (I1076875,I1077404,I1077353);
nand I_63230 (I1076872,I1077387,I1077271);
not I_63231 (I1077476,I2514);
DFFARX1 I_63232 (I535147,I2507,I1077476,I1077502,);
and I_63233 (I1077510,I1077502,I535162);
DFFARX1 I_63234 (I1077510,I2507,I1077476,I1077459,);
DFFARX1 I_63235 (I535153,I2507,I1077476,I1077550,);
not I_63236 (I1077558,I535147);
not I_63237 (I1077575,I535165);
nand I_63238 (I1077592,I1077575,I1077558);
nor I_63239 (I1077447,I1077550,I1077592);
DFFARX1 I_63240 (I1077592,I2507,I1077476,I1077632,);
not I_63241 (I1077468,I1077632);
not I_63242 (I1077654,I535156);
nand I_63243 (I1077671,I1077575,I1077654);
DFFARX1 I_63244 (I1077671,I2507,I1077476,I1077697,);
not I_63245 (I1077705,I1077697);
not I_63246 (I1077722,I535168);
nand I_63247 (I1077739,I1077722,I535144);
and I_63248 (I1077756,I1077558,I1077739);
nor I_63249 (I1077773,I1077671,I1077756);
DFFARX1 I_63250 (I1077773,I2507,I1077476,I1077444,);
DFFARX1 I_63251 (I1077756,I2507,I1077476,I1077465,);
nor I_63252 (I1077818,I535168,I535144);
nor I_63253 (I1077456,I1077671,I1077818);
or I_63254 (I1077849,I535168,I535144);
nor I_63255 (I1077866,I535150,I535159);
DFFARX1 I_63256 (I1077866,I2507,I1077476,I1077892,);
not I_63257 (I1077900,I1077892);
nor I_63258 (I1077462,I1077900,I1077705);
nand I_63259 (I1077931,I1077900,I1077550);
not I_63260 (I1077948,I535150);
nand I_63261 (I1077965,I1077948,I1077654);
nand I_63262 (I1077982,I1077900,I1077965);
nand I_63263 (I1077453,I1077982,I1077931);
nand I_63264 (I1077450,I1077965,I1077849);
not I_63265 (I1078054,I2514);
DFFARX1 I_63266 (I459375,I2507,I1078054,I1078080,);
and I_63267 (I1078088,I1078080,I459390);
DFFARX1 I_63268 (I1078088,I2507,I1078054,I1078037,);
DFFARX1 I_63269 (I459393,I2507,I1078054,I1078128,);
not I_63270 (I1078136,I459387);
not I_63271 (I1078153,I459402);
nand I_63272 (I1078170,I1078153,I1078136);
nor I_63273 (I1078025,I1078128,I1078170);
DFFARX1 I_63274 (I1078170,I2507,I1078054,I1078210,);
not I_63275 (I1078046,I1078210);
not I_63276 (I1078232,I459378);
nand I_63277 (I1078249,I1078153,I1078232);
DFFARX1 I_63278 (I1078249,I2507,I1078054,I1078275,);
not I_63279 (I1078283,I1078275);
not I_63280 (I1078300,I459381);
nand I_63281 (I1078317,I1078300,I459375);
and I_63282 (I1078334,I1078136,I1078317);
nor I_63283 (I1078351,I1078249,I1078334);
DFFARX1 I_63284 (I1078351,I2507,I1078054,I1078022,);
DFFARX1 I_63285 (I1078334,I2507,I1078054,I1078043,);
nor I_63286 (I1078396,I459381,I459384);
nor I_63287 (I1078034,I1078249,I1078396);
or I_63288 (I1078427,I459381,I459384);
nor I_63289 (I1078444,I459399,I459396);
DFFARX1 I_63290 (I1078444,I2507,I1078054,I1078470,);
not I_63291 (I1078478,I1078470);
nor I_63292 (I1078040,I1078478,I1078283);
nand I_63293 (I1078509,I1078478,I1078128);
not I_63294 (I1078526,I459399);
nand I_63295 (I1078543,I1078526,I1078232);
nand I_63296 (I1078560,I1078478,I1078543);
nand I_63297 (I1078031,I1078560,I1078509);
nand I_63298 (I1078028,I1078543,I1078427);
not I_63299 (I1078632,I2514);
DFFARX1 I_63300 (I1257668,I2507,I1078632,I1078658,);
and I_63301 (I1078666,I1078658,I1257650);
DFFARX1 I_63302 (I1078666,I2507,I1078632,I1078615,);
DFFARX1 I_63303 (I1257659,I2507,I1078632,I1078706,);
not I_63304 (I1078714,I1257644);
not I_63305 (I1078731,I1257656);
nand I_63306 (I1078748,I1078731,I1078714);
nor I_63307 (I1078603,I1078706,I1078748);
DFFARX1 I_63308 (I1078748,I2507,I1078632,I1078788,);
not I_63309 (I1078624,I1078788);
not I_63310 (I1078810,I1257647);
nand I_63311 (I1078827,I1078731,I1078810);
DFFARX1 I_63312 (I1078827,I2507,I1078632,I1078853,);
not I_63313 (I1078861,I1078853);
not I_63314 (I1078878,I1257644);
nand I_63315 (I1078895,I1078878,I1257647);
and I_63316 (I1078912,I1078714,I1078895);
nor I_63317 (I1078929,I1078827,I1078912);
DFFARX1 I_63318 (I1078929,I2507,I1078632,I1078600,);
DFFARX1 I_63319 (I1078912,I2507,I1078632,I1078621,);
nor I_63320 (I1078974,I1257644,I1257665);
nor I_63321 (I1078612,I1078827,I1078974);
or I_63322 (I1079005,I1257644,I1257665);
nor I_63323 (I1079022,I1257653,I1257662);
DFFARX1 I_63324 (I1079022,I2507,I1078632,I1079048,);
not I_63325 (I1079056,I1079048);
nor I_63326 (I1078618,I1079056,I1078861);
nand I_63327 (I1079087,I1079056,I1078706);
not I_63328 (I1079104,I1257653);
nand I_63329 (I1079121,I1079104,I1078810);
nand I_63330 (I1079138,I1079056,I1079121);
nand I_63331 (I1078609,I1079138,I1079087);
nand I_63332 (I1078606,I1079121,I1079005);
not I_63333 (I1079210,I2514);
DFFARX1 I_63334 (I420751,I2507,I1079210,I1079236,);
and I_63335 (I1079244,I1079236,I420766);
DFFARX1 I_63336 (I1079244,I2507,I1079210,I1079193,);
DFFARX1 I_63337 (I420769,I2507,I1079210,I1079284,);
not I_63338 (I1079292,I420763);
not I_63339 (I1079309,I420778);
nand I_63340 (I1079326,I1079309,I1079292);
nor I_63341 (I1079181,I1079284,I1079326);
DFFARX1 I_63342 (I1079326,I2507,I1079210,I1079366,);
not I_63343 (I1079202,I1079366);
not I_63344 (I1079388,I420754);
nand I_63345 (I1079405,I1079309,I1079388);
DFFARX1 I_63346 (I1079405,I2507,I1079210,I1079431,);
not I_63347 (I1079439,I1079431);
not I_63348 (I1079456,I420757);
nand I_63349 (I1079473,I1079456,I420751);
and I_63350 (I1079490,I1079292,I1079473);
nor I_63351 (I1079507,I1079405,I1079490);
DFFARX1 I_63352 (I1079507,I2507,I1079210,I1079178,);
DFFARX1 I_63353 (I1079490,I2507,I1079210,I1079199,);
nor I_63354 (I1079552,I420757,I420760);
nor I_63355 (I1079190,I1079405,I1079552);
or I_63356 (I1079583,I420757,I420760);
nor I_63357 (I1079600,I420775,I420772);
DFFARX1 I_63358 (I1079600,I2507,I1079210,I1079626,);
not I_63359 (I1079634,I1079626);
nor I_63360 (I1079196,I1079634,I1079439);
nand I_63361 (I1079665,I1079634,I1079284);
not I_63362 (I1079682,I420775);
nand I_63363 (I1079699,I1079682,I1079388);
nand I_63364 (I1079716,I1079634,I1079699);
nand I_63365 (I1079187,I1079716,I1079665);
nand I_63366 (I1079184,I1079699,I1079583);
not I_63367 (I1079788,I2514);
DFFARX1 I_63368 (I20605,I2507,I1079788,I1079814,);
and I_63369 (I1079822,I1079814,I20608);
DFFARX1 I_63370 (I1079822,I2507,I1079788,I1079771,);
DFFARX1 I_63371 (I20608,I2507,I1079788,I1079862,);
not I_63372 (I1079870,I20611);
not I_63373 (I1079887,I20626);
nand I_63374 (I1079904,I1079887,I1079870);
nor I_63375 (I1079759,I1079862,I1079904);
DFFARX1 I_63376 (I1079904,I2507,I1079788,I1079944,);
not I_63377 (I1079780,I1079944);
not I_63378 (I1079966,I20620);
nand I_63379 (I1079983,I1079887,I1079966);
DFFARX1 I_63380 (I1079983,I2507,I1079788,I1080009,);
not I_63381 (I1080017,I1080009);
not I_63382 (I1080034,I20623);
nand I_63383 (I1080051,I1080034,I20605);
and I_63384 (I1080068,I1079870,I1080051);
nor I_63385 (I1080085,I1079983,I1080068);
DFFARX1 I_63386 (I1080085,I2507,I1079788,I1079756,);
DFFARX1 I_63387 (I1080068,I2507,I1079788,I1079777,);
nor I_63388 (I1080130,I20623,I20617);
nor I_63389 (I1079768,I1079983,I1080130);
or I_63390 (I1080161,I20623,I20617);
nor I_63391 (I1080178,I20614,I20629);
DFFARX1 I_63392 (I1080178,I2507,I1079788,I1080204,);
not I_63393 (I1080212,I1080204);
nor I_63394 (I1079774,I1080212,I1080017);
nand I_63395 (I1080243,I1080212,I1079862);
not I_63396 (I1080260,I20614);
nand I_63397 (I1080277,I1080260,I1079966);
nand I_63398 (I1080294,I1080212,I1080277);
nand I_63399 (I1079765,I1080294,I1080243);
nand I_63400 (I1079762,I1080277,I1080161);
not I_63401 (I1080366,I2514);
DFFARX1 I_63402 (I1342229,I2507,I1080366,I1080392,);
and I_63403 (I1080400,I1080392,I1342211);
DFFARX1 I_63404 (I1080400,I2507,I1080366,I1080349,);
DFFARX1 I_63405 (I1342202,I2507,I1080366,I1080440,);
not I_63406 (I1080448,I1342217);
not I_63407 (I1080465,I1342205);
nand I_63408 (I1080482,I1080465,I1080448);
nor I_63409 (I1080337,I1080440,I1080482);
DFFARX1 I_63410 (I1080482,I2507,I1080366,I1080522,);
not I_63411 (I1080358,I1080522);
not I_63412 (I1080544,I1342214);
nand I_63413 (I1080561,I1080465,I1080544);
DFFARX1 I_63414 (I1080561,I2507,I1080366,I1080587,);
not I_63415 (I1080595,I1080587);
not I_63416 (I1080612,I1342223);
nand I_63417 (I1080629,I1080612,I1342202);
and I_63418 (I1080646,I1080448,I1080629);
nor I_63419 (I1080663,I1080561,I1080646);
DFFARX1 I_63420 (I1080663,I2507,I1080366,I1080334,);
DFFARX1 I_63421 (I1080646,I2507,I1080366,I1080355,);
nor I_63422 (I1080708,I1342223,I1342226);
nor I_63423 (I1080346,I1080561,I1080708);
or I_63424 (I1080739,I1342223,I1342226);
nor I_63425 (I1080756,I1342220,I1342208);
DFFARX1 I_63426 (I1080756,I2507,I1080366,I1080782,);
not I_63427 (I1080790,I1080782);
nor I_63428 (I1080352,I1080790,I1080595);
nand I_63429 (I1080821,I1080790,I1080440);
not I_63430 (I1080838,I1342220);
nand I_63431 (I1080855,I1080838,I1080544);
nand I_63432 (I1080872,I1080790,I1080855);
nand I_63433 (I1080343,I1080872,I1080821);
nand I_63434 (I1080340,I1080855,I1080739);
not I_63435 (I1080944,I2514);
DFFARX1 I_63436 (I756737,I2507,I1080944,I1080970,);
and I_63437 (I1080978,I1080970,I756725);
DFFARX1 I_63438 (I1080978,I2507,I1080944,I1080927,);
DFFARX1 I_63439 (I756728,I2507,I1080944,I1081018,);
not I_63440 (I1081026,I756722);
not I_63441 (I1081043,I756746);
nand I_63442 (I1081060,I1081043,I1081026);
nor I_63443 (I1080915,I1081018,I1081060);
DFFARX1 I_63444 (I1081060,I2507,I1080944,I1081100,);
not I_63445 (I1080936,I1081100);
not I_63446 (I1081122,I756734);
nand I_63447 (I1081139,I1081043,I1081122);
DFFARX1 I_63448 (I1081139,I2507,I1080944,I1081165,);
not I_63449 (I1081173,I1081165);
not I_63450 (I1081190,I756743);
nand I_63451 (I1081207,I1081190,I756740);
and I_63452 (I1081224,I1081026,I1081207);
nor I_63453 (I1081241,I1081139,I1081224);
DFFARX1 I_63454 (I1081241,I2507,I1080944,I1080912,);
DFFARX1 I_63455 (I1081224,I2507,I1080944,I1080933,);
nor I_63456 (I1081286,I756743,I756731);
nor I_63457 (I1080924,I1081139,I1081286);
or I_63458 (I1081317,I756743,I756731);
nor I_63459 (I1081334,I756722,I756725);
DFFARX1 I_63460 (I1081334,I2507,I1080944,I1081360,);
not I_63461 (I1081368,I1081360);
nor I_63462 (I1080930,I1081368,I1081173);
nand I_63463 (I1081399,I1081368,I1081018);
not I_63464 (I1081416,I756722);
nand I_63465 (I1081433,I1081416,I1081122);
nand I_63466 (I1081450,I1081368,I1081433);
nand I_63467 (I1080921,I1081450,I1081399);
nand I_63468 (I1080918,I1081433,I1081317);
not I_63469 (I1081522,I2514);
DFFARX1 I_63470 (I55411,I2507,I1081522,I1081548,);
and I_63471 (I1081556,I1081548,I55387);
DFFARX1 I_63472 (I1081556,I2507,I1081522,I1081505,);
DFFARX1 I_63473 (I55405,I2507,I1081522,I1081596,);
not I_63474 (I1081604,I55393);
not I_63475 (I1081621,I55390);
nand I_63476 (I1081638,I1081621,I1081604);
nor I_63477 (I1081493,I1081596,I1081638);
DFFARX1 I_63478 (I1081638,I2507,I1081522,I1081678,);
not I_63479 (I1081514,I1081678);
not I_63480 (I1081700,I55399);
nand I_63481 (I1081717,I1081621,I1081700);
DFFARX1 I_63482 (I1081717,I2507,I1081522,I1081743,);
not I_63483 (I1081751,I1081743);
not I_63484 (I1081768,I55390);
nand I_63485 (I1081785,I1081768,I55408);
and I_63486 (I1081802,I1081604,I1081785);
nor I_63487 (I1081819,I1081717,I1081802);
DFFARX1 I_63488 (I1081819,I2507,I1081522,I1081490,);
DFFARX1 I_63489 (I1081802,I2507,I1081522,I1081511,);
nor I_63490 (I1081864,I55390,I55402);
nor I_63491 (I1081502,I1081717,I1081864);
or I_63492 (I1081895,I55390,I55402);
nor I_63493 (I1081912,I55396,I55387);
DFFARX1 I_63494 (I1081912,I2507,I1081522,I1081938,);
not I_63495 (I1081946,I1081938);
nor I_63496 (I1081508,I1081946,I1081751);
nand I_63497 (I1081977,I1081946,I1081596);
not I_63498 (I1081994,I55396);
nand I_63499 (I1082011,I1081994,I1081700);
nand I_63500 (I1082028,I1081946,I1082011);
nand I_63501 (I1081499,I1082028,I1081977);
nand I_63502 (I1081496,I1082011,I1081895);
not I_63503 (I1082100,I2514);
DFFARX1 I_63504 (I1276164,I2507,I1082100,I1082126,);
and I_63505 (I1082134,I1082126,I1276146);
DFFARX1 I_63506 (I1082134,I2507,I1082100,I1082083,);
DFFARX1 I_63507 (I1276155,I2507,I1082100,I1082174,);
not I_63508 (I1082182,I1276140);
not I_63509 (I1082199,I1276152);
nand I_63510 (I1082216,I1082199,I1082182);
nor I_63511 (I1082071,I1082174,I1082216);
DFFARX1 I_63512 (I1082216,I2507,I1082100,I1082256,);
not I_63513 (I1082092,I1082256);
not I_63514 (I1082278,I1276143);
nand I_63515 (I1082295,I1082199,I1082278);
DFFARX1 I_63516 (I1082295,I2507,I1082100,I1082321,);
not I_63517 (I1082329,I1082321);
not I_63518 (I1082346,I1276140);
nand I_63519 (I1082363,I1082346,I1276143);
and I_63520 (I1082380,I1082182,I1082363);
nor I_63521 (I1082397,I1082295,I1082380);
DFFARX1 I_63522 (I1082397,I2507,I1082100,I1082068,);
DFFARX1 I_63523 (I1082380,I2507,I1082100,I1082089,);
nor I_63524 (I1082442,I1276140,I1276161);
nor I_63525 (I1082080,I1082295,I1082442);
or I_63526 (I1082473,I1276140,I1276161);
nor I_63527 (I1082490,I1276149,I1276158);
DFFARX1 I_63528 (I1082490,I2507,I1082100,I1082516,);
not I_63529 (I1082524,I1082516);
nor I_63530 (I1082086,I1082524,I1082329);
nand I_63531 (I1082555,I1082524,I1082174);
not I_63532 (I1082572,I1276149);
nand I_63533 (I1082589,I1082572,I1082278);
nand I_63534 (I1082606,I1082524,I1082589);
nand I_63535 (I1082077,I1082606,I1082555);
nand I_63536 (I1082074,I1082589,I1082473);
not I_63537 (I1082678,I2514);
DFFARX1 I_63538 (I278148,I2507,I1082678,I1082704,);
and I_63539 (I1082712,I1082704,I278133);
DFFARX1 I_63540 (I1082712,I2507,I1082678,I1082661,);
DFFARX1 I_63541 (I278139,I2507,I1082678,I1082752,);
not I_63542 (I1082760,I278121);
not I_63543 (I1082777,I278142);
nand I_63544 (I1082794,I1082777,I1082760);
nor I_63545 (I1082649,I1082752,I1082794);
DFFARX1 I_63546 (I1082794,I2507,I1082678,I1082834,);
not I_63547 (I1082670,I1082834);
not I_63548 (I1082856,I278145);
nand I_63549 (I1082873,I1082777,I1082856);
DFFARX1 I_63550 (I1082873,I2507,I1082678,I1082899,);
not I_63551 (I1082907,I1082899);
not I_63552 (I1082924,I278136);
nand I_63553 (I1082941,I1082924,I278124);
and I_63554 (I1082958,I1082760,I1082941);
nor I_63555 (I1082975,I1082873,I1082958);
DFFARX1 I_63556 (I1082975,I2507,I1082678,I1082646,);
DFFARX1 I_63557 (I1082958,I2507,I1082678,I1082667,);
nor I_63558 (I1083020,I278136,I278130);
nor I_63559 (I1082658,I1082873,I1083020);
or I_63560 (I1083051,I278136,I278130);
nor I_63561 (I1083068,I278127,I278121);
DFFARX1 I_63562 (I1083068,I2507,I1082678,I1083094,);
not I_63563 (I1083102,I1083094);
nor I_63564 (I1082664,I1083102,I1082907);
nand I_63565 (I1083133,I1083102,I1082752);
not I_63566 (I1083150,I278127);
nand I_63567 (I1083167,I1083150,I1082856);
nand I_63568 (I1083184,I1083102,I1083167);
nand I_63569 (I1082655,I1083184,I1083133);
nand I_63570 (I1082652,I1083167,I1083051);
not I_63571 (I1083256,I2514);
DFFARX1 I_63572 (I651541,I2507,I1083256,I1083282,);
and I_63573 (I1083290,I1083282,I651529);
DFFARX1 I_63574 (I1083290,I2507,I1083256,I1083239,);
DFFARX1 I_63575 (I651532,I2507,I1083256,I1083330,);
not I_63576 (I1083338,I651526);
not I_63577 (I1083355,I651550);
nand I_63578 (I1083372,I1083355,I1083338);
nor I_63579 (I1083227,I1083330,I1083372);
DFFARX1 I_63580 (I1083372,I2507,I1083256,I1083412,);
not I_63581 (I1083248,I1083412);
not I_63582 (I1083434,I651538);
nand I_63583 (I1083451,I1083355,I1083434);
DFFARX1 I_63584 (I1083451,I2507,I1083256,I1083477,);
not I_63585 (I1083485,I1083477);
not I_63586 (I1083502,I651547);
nand I_63587 (I1083519,I1083502,I651544);
and I_63588 (I1083536,I1083338,I1083519);
nor I_63589 (I1083553,I1083451,I1083536);
DFFARX1 I_63590 (I1083553,I2507,I1083256,I1083224,);
DFFARX1 I_63591 (I1083536,I2507,I1083256,I1083245,);
nor I_63592 (I1083598,I651547,I651535);
nor I_63593 (I1083236,I1083451,I1083598);
or I_63594 (I1083629,I651547,I651535);
nor I_63595 (I1083646,I651526,I651529);
DFFARX1 I_63596 (I1083646,I2507,I1083256,I1083672,);
not I_63597 (I1083680,I1083672);
nor I_63598 (I1083242,I1083680,I1083485);
nand I_63599 (I1083711,I1083680,I1083330);
not I_63600 (I1083728,I651526);
nand I_63601 (I1083745,I1083728,I1083434);
nand I_63602 (I1083762,I1083680,I1083745);
nand I_63603 (I1083233,I1083762,I1083711);
nand I_63604 (I1083230,I1083745,I1083629);
not I_63605 (I1083834,I2514);
DFFARX1 I_63606 (I92301,I2507,I1083834,I1083860,);
and I_63607 (I1083868,I1083860,I92277);
DFFARX1 I_63608 (I1083868,I2507,I1083834,I1083817,);
DFFARX1 I_63609 (I92295,I2507,I1083834,I1083908,);
not I_63610 (I1083916,I92283);
not I_63611 (I1083933,I92280);
nand I_63612 (I1083950,I1083933,I1083916);
nor I_63613 (I1083805,I1083908,I1083950);
DFFARX1 I_63614 (I1083950,I2507,I1083834,I1083990,);
not I_63615 (I1083826,I1083990);
not I_63616 (I1084012,I92289);
nand I_63617 (I1084029,I1083933,I1084012);
DFFARX1 I_63618 (I1084029,I2507,I1083834,I1084055,);
not I_63619 (I1084063,I1084055);
not I_63620 (I1084080,I92280);
nand I_63621 (I1084097,I1084080,I92298);
and I_63622 (I1084114,I1083916,I1084097);
nor I_63623 (I1084131,I1084029,I1084114);
DFFARX1 I_63624 (I1084131,I2507,I1083834,I1083802,);
DFFARX1 I_63625 (I1084114,I2507,I1083834,I1083823,);
nor I_63626 (I1084176,I92280,I92292);
nor I_63627 (I1083814,I1084029,I1084176);
or I_63628 (I1084207,I92280,I92292);
nor I_63629 (I1084224,I92286,I92277);
DFFARX1 I_63630 (I1084224,I2507,I1083834,I1084250,);
not I_63631 (I1084258,I1084250);
nor I_63632 (I1083820,I1084258,I1084063);
nand I_63633 (I1084289,I1084258,I1083908);
not I_63634 (I1084306,I92286);
nand I_63635 (I1084323,I1084306,I1084012);
nand I_63636 (I1084340,I1084258,I1084323);
nand I_63637 (I1083811,I1084340,I1084289);
nand I_63638 (I1083808,I1084323,I1084207);
not I_63639 (I1084412,I2514);
DFFARX1 I_63640 (I1393399,I2507,I1084412,I1084438,);
and I_63641 (I1084446,I1084438,I1393381);
DFFARX1 I_63642 (I1084446,I2507,I1084412,I1084395,);
DFFARX1 I_63643 (I1393372,I2507,I1084412,I1084486,);
not I_63644 (I1084494,I1393387);
not I_63645 (I1084511,I1393375);
nand I_63646 (I1084528,I1084511,I1084494);
nor I_63647 (I1084383,I1084486,I1084528);
DFFARX1 I_63648 (I1084528,I2507,I1084412,I1084568,);
not I_63649 (I1084404,I1084568);
not I_63650 (I1084590,I1393384);
nand I_63651 (I1084607,I1084511,I1084590);
DFFARX1 I_63652 (I1084607,I2507,I1084412,I1084633,);
not I_63653 (I1084641,I1084633);
not I_63654 (I1084658,I1393393);
nand I_63655 (I1084675,I1084658,I1393372);
and I_63656 (I1084692,I1084494,I1084675);
nor I_63657 (I1084709,I1084607,I1084692);
DFFARX1 I_63658 (I1084709,I2507,I1084412,I1084380,);
DFFARX1 I_63659 (I1084692,I2507,I1084412,I1084401,);
nor I_63660 (I1084754,I1393393,I1393396);
nor I_63661 (I1084392,I1084607,I1084754);
or I_63662 (I1084785,I1393393,I1393396);
nor I_63663 (I1084802,I1393390,I1393378);
DFFARX1 I_63664 (I1084802,I2507,I1084412,I1084828,);
not I_63665 (I1084836,I1084828);
nor I_63666 (I1084398,I1084836,I1084641);
nand I_63667 (I1084867,I1084836,I1084486);
not I_63668 (I1084884,I1393390);
nand I_63669 (I1084901,I1084884,I1084590);
nand I_63670 (I1084918,I1084836,I1084901);
nand I_63671 (I1084389,I1084918,I1084867);
nand I_63672 (I1084386,I1084901,I1084785);
not I_63673 (I1084990,I2514);
DFFARX1 I_63674 (I52776,I2507,I1084990,I1085016,);
and I_63675 (I1085024,I1085016,I52752);
DFFARX1 I_63676 (I1085024,I2507,I1084990,I1084973,);
DFFARX1 I_63677 (I52770,I2507,I1084990,I1085064,);
not I_63678 (I1085072,I52758);
not I_63679 (I1085089,I52755);
nand I_63680 (I1085106,I1085089,I1085072);
nor I_63681 (I1084961,I1085064,I1085106);
DFFARX1 I_63682 (I1085106,I2507,I1084990,I1085146,);
not I_63683 (I1084982,I1085146);
not I_63684 (I1085168,I52764);
nand I_63685 (I1085185,I1085089,I1085168);
DFFARX1 I_63686 (I1085185,I2507,I1084990,I1085211,);
not I_63687 (I1085219,I1085211);
not I_63688 (I1085236,I52755);
nand I_63689 (I1085253,I1085236,I52773);
and I_63690 (I1085270,I1085072,I1085253);
nor I_63691 (I1085287,I1085185,I1085270);
DFFARX1 I_63692 (I1085287,I2507,I1084990,I1084958,);
DFFARX1 I_63693 (I1085270,I2507,I1084990,I1084979,);
nor I_63694 (I1085332,I52755,I52767);
nor I_63695 (I1084970,I1085185,I1085332);
or I_63696 (I1085363,I52755,I52767);
nor I_63697 (I1085380,I52761,I52752);
DFFARX1 I_63698 (I1085380,I2507,I1084990,I1085406,);
not I_63699 (I1085414,I1085406);
nor I_63700 (I1084976,I1085414,I1085219);
nand I_63701 (I1085445,I1085414,I1085064);
not I_63702 (I1085462,I52761);
nand I_63703 (I1085479,I1085462,I1085168);
nand I_63704 (I1085496,I1085414,I1085479);
nand I_63705 (I1084967,I1085496,I1085445);
nand I_63706 (I1084964,I1085479,I1085363);
not I_63707 (I1085568,I2514);
DFFARX1 I_63708 (I837033,I2507,I1085568,I1085594,);
and I_63709 (I1085602,I1085594,I837039);
DFFARX1 I_63710 (I1085602,I2507,I1085568,I1085551,);
DFFARX1 I_63711 (I837045,I2507,I1085568,I1085642,);
not I_63712 (I1085650,I837030);
not I_63713 (I1085667,I837030);
nand I_63714 (I1085684,I1085667,I1085650);
nor I_63715 (I1085539,I1085642,I1085684);
DFFARX1 I_63716 (I1085684,I2507,I1085568,I1085724,);
not I_63717 (I1085560,I1085724);
not I_63718 (I1085746,I837048);
nand I_63719 (I1085763,I1085667,I1085746);
DFFARX1 I_63720 (I1085763,I2507,I1085568,I1085789,);
not I_63721 (I1085797,I1085789);
not I_63722 (I1085814,I837042);
nand I_63723 (I1085831,I1085814,I837033);
and I_63724 (I1085848,I1085650,I1085831);
nor I_63725 (I1085865,I1085763,I1085848);
DFFARX1 I_63726 (I1085865,I2507,I1085568,I1085536,);
DFFARX1 I_63727 (I1085848,I2507,I1085568,I1085557,);
nor I_63728 (I1085910,I837042,I837051);
nor I_63729 (I1085548,I1085763,I1085910);
or I_63730 (I1085941,I837042,I837051);
nor I_63731 (I1085958,I837036,I837036);
DFFARX1 I_63732 (I1085958,I2507,I1085568,I1085984,);
not I_63733 (I1085992,I1085984);
nor I_63734 (I1085554,I1085992,I1085797);
nand I_63735 (I1086023,I1085992,I1085642);
not I_63736 (I1086040,I837036);
nand I_63737 (I1086057,I1086040,I1085746);
nand I_63738 (I1086074,I1085992,I1086057);
nand I_63739 (I1085545,I1086074,I1086023);
nand I_63740 (I1085542,I1086057,I1085941);
not I_63741 (I1086146,I2514);
DFFARX1 I_63742 (I1227031,I2507,I1086146,I1086172,);
and I_63743 (I1086180,I1086172,I1227025);
DFFARX1 I_63744 (I1086180,I2507,I1086146,I1086129,);
DFFARX1 I_63745 (I1227010,I2507,I1086146,I1086220,);
not I_63746 (I1086228,I1227016);
not I_63747 (I1086245,I1227028);
nand I_63748 (I1086262,I1086245,I1086228);
nor I_63749 (I1086117,I1086220,I1086262);
DFFARX1 I_63750 (I1086262,I2507,I1086146,I1086302,);
not I_63751 (I1086138,I1086302);
not I_63752 (I1086324,I1227010);
nand I_63753 (I1086341,I1086245,I1086324);
DFFARX1 I_63754 (I1086341,I2507,I1086146,I1086367,);
not I_63755 (I1086375,I1086367);
not I_63756 (I1086392,I1227034);
nand I_63757 (I1086409,I1086392,I1227022);
and I_63758 (I1086426,I1086228,I1086409);
nor I_63759 (I1086443,I1086341,I1086426);
DFFARX1 I_63760 (I1086443,I2507,I1086146,I1086114,);
DFFARX1 I_63761 (I1086426,I2507,I1086146,I1086135,);
nor I_63762 (I1086488,I1227034,I1227013);
nor I_63763 (I1086126,I1086341,I1086488);
or I_63764 (I1086519,I1227034,I1227013);
nor I_63765 (I1086536,I1227019,I1227013);
DFFARX1 I_63766 (I1086536,I2507,I1086146,I1086562,);
not I_63767 (I1086570,I1086562);
nor I_63768 (I1086132,I1086570,I1086375);
nand I_63769 (I1086601,I1086570,I1086220);
not I_63770 (I1086618,I1227019);
nand I_63771 (I1086635,I1086618,I1086324);
nand I_63772 (I1086652,I1086570,I1086635);
nand I_63773 (I1086123,I1086652,I1086601);
nand I_63774 (I1086120,I1086635,I1086519);
not I_63775 (I1086724,I2514);
DFFARX1 I_63776 (I1261714,I2507,I1086724,I1086750,);
and I_63777 (I1086758,I1086750,I1261696);
DFFARX1 I_63778 (I1086758,I2507,I1086724,I1086707,);
DFFARX1 I_63779 (I1261705,I2507,I1086724,I1086798,);
not I_63780 (I1086806,I1261690);
not I_63781 (I1086823,I1261702);
nand I_63782 (I1086840,I1086823,I1086806);
nor I_63783 (I1086695,I1086798,I1086840);
DFFARX1 I_63784 (I1086840,I2507,I1086724,I1086880,);
not I_63785 (I1086716,I1086880);
not I_63786 (I1086902,I1261693);
nand I_63787 (I1086919,I1086823,I1086902);
DFFARX1 I_63788 (I1086919,I2507,I1086724,I1086945,);
not I_63789 (I1086953,I1086945);
not I_63790 (I1086970,I1261690);
nand I_63791 (I1086987,I1086970,I1261693);
and I_63792 (I1087004,I1086806,I1086987);
nor I_63793 (I1087021,I1086919,I1087004);
DFFARX1 I_63794 (I1087021,I2507,I1086724,I1086692,);
DFFARX1 I_63795 (I1087004,I2507,I1086724,I1086713,);
nor I_63796 (I1087066,I1261690,I1261711);
nor I_63797 (I1086704,I1086919,I1087066);
or I_63798 (I1087097,I1261690,I1261711);
nor I_63799 (I1087114,I1261699,I1261708);
DFFARX1 I_63800 (I1087114,I2507,I1086724,I1087140,);
not I_63801 (I1087148,I1087140);
nor I_63802 (I1086710,I1087148,I1086953);
nand I_63803 (I1087179,I1087148,I1086798);
not I_63804 (I1087196,I1261699);
nand I_63805 (I1087213,I1087196,I1086902);
nand I_63806 (I1087230,I1087148,I1087213);
nand I_63807 (I1086701,I1087230,I1087179);
nand I_63808 (I1086698,I1087213,I1087097);
not I_63809 (I1087302,I2514);
DFFARX1 I_63810 (I726681,I2507,I1087302,I1087328,);
and I_63811 (I1087336,I1087328,I726669);
DFFARX1 I_63812 (I1087336,I2507,I1087302,I1087285,);
DFFARX1 I_63813 (I726672,I2507,I1087302,I1087376,);
not I_63814 (I1087384,I726666);
not I_63815 (I1087401,I726690);
nand I_63816 (I1087418,I1087401,I1087384);
nor I_63817 (I1087273,I1087376,I1087418);
DFFARX1 I_63818 (I1087418,I2507,I1087302,I1087458,);
not I_63819 (I1087294,I1087458);
not I_63820 (I1087480,I726678);
nand I_63821 (I1087497,I1087401,I1087480);
DFFARX1 I_63822 (I1087497,I2507,I1087302,I1087523,);
not I_63823 (I1087531,I1087523);
not I_63824 (I1087548,I726687);
nand I_63825 (I1087565,I1087548,I726684);
and I_63826 (I1087582,I1087384,I1087565);
nor I_63827 (I1087599,I1087497,I1087582);
DFFARX1 I_63828 (I1087599,I2507,I1087302,I1087270,);
DFFARX1 I_63829 (I1087582,I2507,I1087302,I1087291,);
nor I_63830 (I1087644,I726687,I726675);
nor I_63831 (I1087282,I1087497,I1087644);
or I_63832 (I1087675,I726687,I726675);
nor I_63833 (I1087692,I726666,I726669);
DFFARX1 I_63834 (I1087692,I2507,I1087302,I1087718,);
not I_63835 (I1087726,I1087718);
nor I_63836 (I1087288,I1087726,I1087531);
nand I_63837 (I1087757,I1087726,I1087376);
not I_63838 (I1087774,I726666);
nand I_63839 (I1087791,I1087774,I1087480);
nand I_63840 (I1087808,I1087726,I1087791);
nand I_63841 (I1087279,I1087808,I1087757);
nand I_63842 (I1087276,I1087791,I1087675);
not I_63843 (I1087880,I2514);
DFFARX1 I_63844 (I1358294,I2507,I1087880,I1087906,);
and I_63845 (I1087914,I1087906,I1358276);
DFFARX1 I_63846 (I1087914,I2507,I1087880,I1087863,);
DFFARX1 I_63847 (I1358267,I2507,I1087880,I1087954,);
not I_63848 (I1087962,I1358282);
not I_63849 (I1087979,I1358270);
nand I_63850 (I1087996,I1087979,I1087962);
nor I_63851 (I1087851,I1087954,I1087996);
DFFARX1 I_63852 (I1087996,I2507,I1087880,I1088036,);
not I_63853 (I1087872,I1088036);
not I_63854 (I1088058,I1358279);
nand I_63855 (I1088075,I1087979,I1088058);
DFFARX1 I_63856 (I1088075,I2507,I1087880,I1088101,);
not I_63857 (I1088109,I1088101);
not I_63858 (I1088126,I1358288);
nand I_63859 (I1088143,I1088126,I1358267);
and I_63860 (I1088160,I1087962,I1088143);
nor I_63861 (I1088177,I1088075,I1088160);
DFFARX1 I_63862 (I1088177,I2507,I1087880,I1087848,);
DFFARX1 I_63863 (I1088160,I2507,I1087880,I1087869,);
nor I_63864 (I1088222,I1358288,I1358291);
nor I_63865 (I1087860,I1088075,I1088222);
or I_63866 (I1088253,I1358288,I1358291);
nor I_63867 (I1088270,I1358285,I1358273);
DFFARX1 I_63868 (I1088270,I2507,I1087880,I1088296,);
not I_63869 (I1088304,I1088296);
nor I_63870 (I1087866,I1088304,I1088109);
nand I_63871 (I1088335,I1088304,I1087954);
not I_63872 (I1088352,I1358285);
nand I_63873 (I1088369,I1088352,I1088058);
nand I_63874 (I1088386,I1088304,I1088369);
nand I_63875 (I1087857,I1088386,I1088335);
nand I_63876 (I1087854,I1088369,I1088253);
not I_63877 (I1088458,I2514);
DFFARX1 I_63878 (I559639,I2507,I1088458,I1088484,);
and I_63879 (I1088492,I1088484,I559627);
DFFARX1 I_63880 (I1088492,I2507,I1088458,I1088441,);
DFFARX1 I_63881 (I559642,I2507,I1088458,I1088532,);
not I_63882 (I1088540,I559633);
not I_63883 (I1088557,I559624);
nand I_63884 (I1088574,I1088557,I1088540);
nor I_63885 (I1088429,I1088532,I1088574);
DFFARX1 I_63886 (I1088574,I2507,I1088458,I1088614,);
not I_63887 (I1088450,I1088614);
not I_63888 (I1088636,I559630);
nand I_63889 (I1088653,I1088557,I1088636);
DFFARX1 I_63890 (I1088653,I2507,I1088458,I1088679,);
not I_63891 (I1088687,I1088679);
not I_63892 (I1088704,I559645);
nand I_63893 (I1088721,I1088704,I559648);
and I_63894 (I1088738,I1088540,I1088721);
nor I_63895 (I1088755,I1088653,I1088738);
DFFARX1 I_63896 (I1088755,I2507,I1088458,I1088426,);
DFFARX1 I_63897 (I1088738,I2507,I1088458,I1088447,);
nor I_63898 (I1088800,I559645,I559624);
nor I_63899 (I1088438,I1088653,I1088800);
or I_63900 (I1088831,I559645,I559624);
nor I_63901 (I1088848,I559636,I559627);
DFFARX1 I_63902 (I1088848,I2507,I1088458,I1088874,);
not I_63903 (I1088882,I1088874);
nor I_63904 (I1088444,I1088882,I1088687);
nand I_63905 (I1088913,I1088882,I1088532);
not I_63906 (I1088930,I559636);
nand I_63907 (I1088947,I1088930,I1088636);
nand I_63908 (I1088964,I1088882,I1088947);
nand I_63909 (I1088435,I1088964,I1088913);
nand I_63910 (I1088432,I1088947,I1088831);
not I_63911 (I1089036,I2514);
DFFARX1 I_63912 (I887577,I2507,I1089036,I1089062,);
and I_63913 (I1089070,I1089062,I887571);
DFFARX1 I_63914 (I1089070,I2507,I1089036,I1089019,);
DFFARX1 I_63915 (I887589,I2507,I1089036,I1089110,);
not I_63916 (I1089118,I887580);
not I_63917 (I1089135,I887592);
nand I_63918 (I1089152,I1089135,I1089118);
nor I_63919 (I1089007,I1089110,I1089152);
DFFARX1 I_63920 (I1089152,I2507,I1089036,I1089192,);
not I_63921 (I1089028,I1089192);
not I_63922 (I1089214,I887598);
nand I_63923 (I1089231,I1089135,I1089214);
DFFARX1 I_63924 (I1089231,I2507,I1089036,I1089257,);
not I_63925 (I1089265,I1089257);
not I_63926 (I1089282,I887574);
nand I_63927 (I1089299,I1089282,I887595);
and I_63928 (I1089316,I1089118,I1089299);
nor I_63929 (I1089333,I1089231,I1089316);
DFFARX1 I_63930 (I1089333,I2507,I1089036,I1089004,);
DFFARX1 I_63931 (I1089316,I2507,I1089036,I1089025,);
nor I_63932 (I1089378,I887574,I887586);
nor I_63933 (I1089016,I1089231,I1089378);
or I_63934 (I1089409,I887574,I887586);
nor I_63935 (I1089426,I887571,I887583);
DFFARX1 I_63936 (I1089426,I2507,I1089036,I1089452,);
not I_63937 (I1089460,I1089452);
nor I_63938 (I1089022,I1089460,I1089265);
nand I_63939 (I1089491,I1089460,I1089110);
not I_63940 (I1089508,I887571);
nand I_63941 (I1089525,I1089508,I1089214);
nand I_63942 (I1089542,I1089460,I1089525);
nand I_63943 (I1089013,I1089542,I1089491);
nand I_63944 (I1089010,I1089525,I1089409);
not I_63945 (I1089614,I2514);
DFFARX1 I_63946 (I675817,I2507,I1089614,I1089640,);
and I_63947 (I1089648,I1089640,I675805);
DFFARX1 I_63948 (I1089648,I2507,I1089614,I1089597,);
DFFARX1 I_63949 (I675808,I2507,I1089614,I1089688,);
not I_63950 (I1089696,I675802);
not I_63951 (I1089713,I675826);
nand I_63952 (I1089730,I1089713,I1089696);
nor I_63953 (I1089585,I1089688,I1089730);
DFFARX1 I_63954 (I1089730,I2507,I1089614,I1089770,);
not I_63955 (I1089606,I1089770);
not I_63956 (I1089792,I675814);
nand I_63957 (I1089809,I1089713,I1089792);
DFFARX1 I_63958 (I1089809,I2507,I1089614,I1089835,);
not I_63959 (I1089843,I1089835);
not I_63960 (I1089860,I675823);
nand I_63961 (I1089877,I1089860,I675820);
and I_63962 (I1089894,I1089696,I1089877);
nor I_63963 (I1089911,I1089809,I1089894);
DFFARX1 I_63964 (I1089911,I2507,I1089614,I1089582,);
DFFARX1 I_63965 (I1089894,I2507,I1089614,I1089603,);
nor I_63966 (I1089956,I675823,I675811);
nor I_63967 (I1089594,I1089809,I1089956);
or I_63968 (I1089987,I675823,I675811);
nor I_63969 (I1090004,I675802,I675805);
DFFARX1 I_63970 (I1090004,I2507,I1089614,I1090030,);
not I_63971 (I1090038,I1090030);
nor I_63972 (I1089600,I1090038,I1089843);
nand I_63973 (I1090069,I1090038,I1089688);
not I_63974 (I1090086,I675802);
nand I_63975 (I1090103,I1090086,I1089792);
nand I_63976 (I1090120,I1090038,I1090103);
nand I_63977 (I1089591,I1090120,I1090069);
nand I_63978 (I1089588,I1090103,I1089987);
not I_63979 (I1090192,I2514);
DFFARX1 I_63980 (I839141,I2507,I1090192,I1090218,);
and I_63981 (I1090226,I1090218,I839147);
DFFARX1 I_63982 (I1090226,I2507,I1090192,I1090175,);
DFFARX1 I_63983 (I839153,I2507,I1090192,I1090266,);
not I_63984 (I1090274,I839138);
not I_63985 (I1090291,I839138);
nand I_63986 (I1090308,I1090291,I1090274);
nor I_63987 (I1090163,I1090266,I1090308);
DFFARX1 I_63988 (I1090308,I2507,I1090192,I1090348,);
not I_63989 (I1090184,I1090348);
not I_63990 (I1090370,I839156);
nand I_63991 (I1090387,I1090291,I1090370);
DFFARX1 I_63992 (I1090387,I2507,I1090192,I1090413,);
not I_63993 (I1090421,I1090413);
not I_63994 (I1090438,I839150);
nand I_63995 (I1090455,I1090438,I839141);
and I_63996 (I1090472,I1090274,I1090455);
nor I_63997 (I1090489,I1090387,I1090472);
DFFARX1 I_63998 (I1090489,I2507,I1090192,I1090160,);
DFFARX1 I_63999 (I1090472,I2507,I1090192,I1090181,);
nor I_64000 (I1090534,I839150,I839159);
nor I_64001 (I1090172,I1090387,I1090534);
or I_64002 (I1090565,I839150,I839159);
nor I_64003 (I1090582,I839144,I839144);
DFFARX1 I_64004 (I1090582,I2507,I1090192,I1090608,);
not I_64005 (I1090616,I1090608);
nor I_64006 (I1090178,I1090616,I1090421);
nand I_64007 (I1090647,I1090616,I1090266);
not I_64008 (I1090664,I839144);
nand I_64009 (I1090681,I1090664,I1090370);
nand I_64010 (I1090698,I1090616,I1090681);
nand I_64011 (I1090169,I1090698,I1090647);
nand I_64012 (I1090166,I1090681,I1090565);
not I_64013 (I1090770,I2514);
DFFARX1 I_64014 (I1240087,I2507,I1090770,I1090796,);
and I_64015 (I1090804,I1090796,I1240081);
DFFARX1 I_64016 (I1090804,I2507,I1090770,I1090753,);
DFFARX1 I_64017 (I1240066,I2507,I1090770,I1090844,);
not I_64018 (I1090852,I1240072);
not I_64019 (I1090869,I1240084);
nand I_64020 (I1090886,I1090869,I1090852);
nor I_64021 (I1090741,I1090844,I1090886);
DFFARX1 I_64022 (I1090886,I2507,I1090770,I1090926,);
not I_64023 (I1090762,I1090926);
not I_64024 (I1090948,I1240066);
nand I_64025 (I1090965,I1090869,I1090948);
DFFARX1 I_64026 (I1090965,I2507,I1090770,I1090991,);
not I_64027 (I1090999,I1090991);
not I_64028 (I1091016,I1240090);
nand I_64029 (I1091033,I1091016,I1240078);
and I_64030 (I1091050,I1090852,I1091033);
nor I_64031 (I1091067,I1090965,I1091050);
DFFARX1 I_64032 (I1091067,I2507,I1090770,I1090738,);
DFFARX1 I_64033 (I1091050,I2507,I1090770,I1090759,);
nor I_64034 (I1091112,I1240090,I1240069);
nor I_64035 (I1090750,I1090965,I1091112);
or I_64036 (I1091143,I1240090,I1240069);
nor I_64037 (I1091160,I1240075,I1240069);
DFFARX1 I_64038 (I1091160,I2507,I1090770,I1091186,);
not I_64039 (I1091194,I1091186);
nor I_64040 (I1090756,I1091194,I1090999);
nand I_64041 (I1091225,I1091194,I1090844);
not I_64042 (I1091242,I1240075);
nand I_64043 (I1091259,I1091242,I1090948);
nand I_64044 (I1091276,I1091194,I1091259);
nand I_64045 (I1090747,I1091276,I1091225);
nand I_64046 (I1090744,I1091259,I1091143);
not I_64047 (I1091348,I2514);
DFFARX1 I_64048 (I347712,I2507,I1091348,I1091374,);
and I_64049 (I1091382,I1091374,I347697);
DFFARX1 I_64050 (I1091382,I2507,I1091348,I1091331,);
DFFARX1 I_64051 (I347703,I2507,I1091348,I1091422,);
not I_64052 (I1091430,I347685);
not I_64053 (I1091447,I347706);
nand I_64054 (I1091464,I1091447,I1091430);
nor I_64055 (I1091319,I1091422,I1091464);
DFFARX1 I_64056 (I1091464,I2507,I1091348,I1091504,);
not I_64057 (I1091340,I1091504);
not I_64058 (I1091526,I347709);
nand I_64059 (I1091543,I1091447,I1091526);
DFFARX1 I_64060 (I1091543,I2507,I1091348,I1091569,);
not I_64061 (I1091577,I1091569);
not I_64062 (I1091594,I347700);
nand I_64063 (I1091611,I1091594,I347688);
and I_64064 (I1091628,I1091430,I1091611);
nor I_64065 (I1091645,I1091543,I1091628);
DFFARX1 I_64066 (I1091645,I2507,I1091348,I1091316,);
DFFARX1 I_64067 (I1091628,I2507,I1091348,I1091337,);
nor I_64068 (I1091690,I347700,I347694);
nor I_64069 (I1091328,I1091543,I1091690);
or I_64070 (I1091721,I347700,I347694);
nor I_64071 (I1091738,I347691,I347685);
DFFARX1 I_64072 (I1091738,I2507,I1091348,I1091764,);
not I_64073 (I1091772,I1091764);
nor I_64074 (I1091334,I1091772,I1091577);
nand I_64075 (I1091803,I1091772,I1091422);
not I_64076 (I1091820,I347691);
nand I_64077 (I1091837,I1091820,I1091526);
nand I_64078 (I1091854,I1091772,I1091837);
nand I_64079 (I1091325,I1091854,I1091803);
nand I_64080 (I1091322,I1091837,I1091721);
not I_64081 (I1091926,I2514);
DFFARX1 I_64082 (I961867,I2507,I1091926,I1091952,);
and I_64083 (I1091960,I1091952,I961861);
DFFARX1 I_64084 (I1091960,I2507,I1091926,I1091909,);
DFFARX1 I_64085 (I961879,I2507,I1091926,I1092000,);
not I_64086 (I1092008,I961870);
not I_64087 (I1092025,I961882);
nand I_64088 (I1092042,I1092025,I1092008);
nor I_64089 (I1091897,I1092000,I1092042);
DFFARX1 I_64090 (I1092042,I2507,I1091926,I1092082,);
not I_64091 (I1091918,I1092082);
not I_64092 (I1092104,I961888);
nand I_64093 (I1092121,I1092025,I1092104);
DFFARX1 I_64094 (I1092121,I2507,I1091926,I1092147,);
not I_64095 (I1092155,I1092147);
not I_64096 (I1092172,I961864);
nand I_64097 (I1092189,I1092172,I961885);
and I_64098 (I1092206,I1092008,I1092189);
nor I_64099 (I1092223,I1092121,I1092206);
DFFARX1 I_64100 (I1092223,I2507,I1091926,I1091894,);
DFFARX1 I_64101 (I1092206,I2507,I1091926,I1091915,);
nor I_64102 (I1092268,I961864,I961876);
nor I_64103 (I1091906,I1092121,I1092268);
or I_64104 (I1092299,I961864,I961876);
nor I_64105 (I1092316,I961861,I961873);
DFFARX1 I_64106 (I1092316,I2507,I1091926,I1092342,);
not I_64107 (I1092350,I1092342);
nor I_64108 (I1091912,I1092350,I1092155);
nand I_64109 (I1092381,I1092350,I1092000);
not I_64110 (I1092398,I961861);
nand I_64111 (I1092415,I1092398,I1092104);
nand I_64112 (I1092432,I1092350,I1092415);
nand I_64113 (I1091903,I1092432,I1092381);
nand I_64114 (I1091900,I1092415,I1092299);
not I_64115 (I1092504,I2514);
DFFARX1 I_64116 (I1310694,I2507,I1092504,I1092530,);
and I_64117 (I1092538,I1092530,I1310676);
DFFARX1 I_64118 (I1092538,I2507,I1092504,I1092487,);
DFFARX1 I_64119 (I1310667,I2507,I1092504,I1092578,);
not I_64120 (I1092586,I1310682);
not I_64121 (I1092603,I1310670);
nand I_64122 (I1092620,I1092603,I1092586);
nor I_64123 (I1092475,I1092578,I1092620);
DFFARX1 I_64124 (I1092620,I2507,I1092504,I1092660,);
not I_64125 (I1092496,I1092660);
not I_64126 (I1092682,I1310679);
nand I_64127 (I1092699,I1092603,I1092682);
DFFARX1 I_64128 (I1092699,I2507,I1092504,I1092725,);
not I_64129 (I1092733,I1092725);
not I_64130 (I1092750,I1310688);
nand I_64131 (I1092767,I1092750,I1310667);
and I_64132 (I1092784,I1092586,I1092767);
nor I_64133 (I1092801,I1092699,I1092784);
DFFARX1 I_64134 (I1092801,I2507,I1092504,I1092472,);
DFFARX1 I_64135 (I1092784,I2507,I1092504,I1092493,);
nor I_64136 (I1092846,I1310688,I1310691);
nor I_64137 (I1092484,I1092699,I1092846);
or I_64138 (I1092877,I1310688,I1310691);
nor I_64139 (I1092894,I1310685,I1310673);
DFFARX1 I_64140 (I1092894,I2507,I1092504,I1092920,);
not I_64141 (I1092928,I1092920);
nor I_64142 (I1092490,I1092928,I1092733);
nand I_64143 (I1092959,I1092928,I1092578);
not I_64144 (I1092976,I1310685);
nand I_64145 (I1092993,I1092976,I1092682);
nand I_64146 (I1093010,I1092928,I1092993);
nand I_64147 (I1092481,I1093010,I1092959);
nand I_64148 (I1092478,I1092993,I1092877);
not I_64149 (I1093082,I2514);
DFFARX1 I_64150 (I1020803,I2507,I1093082,I1093108,);
and I_64151 (I1093116,I1093108,I1020800);
DFFARX1 I_64152 (I1093116,I2507,I1093082,I1093065,);
DFFARX1 I_64153 (I1020806,I2507,I1093082,I1093156,);
not I_64154 (I1093164,I1020809);
not I_64155 (I1093181,I1020803);
nand I_64156 (I1093198,I1093181,I1093164);
nor I_64157 (I1093053,I1093156,I1093198);
DFFARX1 I_64158 (I1093198,I2507,I1093082,I1093238,);
not I_64159 (I1093074,I1093238);
not I_64160 (I1093260,I1020818);
nand I_64161 (I1093277,I1093181,I1093260);
DFFARX1 I_64162 (I1093277,I2507,I1093082,I1093303,);
not I_64163 (I1093311,I1093303);
not I_64164 (I1093328,I1020815);
nand I_64165 (I1093345,I1093328,I1020821);
and I_64166 (I1093362,I1093164,I1093345);
nor I_64167 (I1093379,I1093277,I1093362);
DFFARX1 I_64168 (I1093379,I2507,I1093082,I1093050,);
DFFARX1 I_64169 (I1093362,I2507,I1093082,I1093071,);
nor I_64170 (I1093424,I1020815,I1020800);
nor I_64171 (I1093062,I1093277,I1093424);
or I_64172 (I1093455,I1020815,I1020800);
nor I_64173 (I1093472,I1020812,I1020806);
DFFARX1 I_64174 (I1093472,I2507,I1093082,I1093498,);
not I_64175 (I1093506,I1093498);
nor I_64176 (I1093068,I1093506,I1093311);
nand I_64177 (I1093537,I1093506,I1093156);
not I_64178 (I1093554,I1020812);
nand I_64179 (I1093571,I1093554,I1093260);
nand I_64180 (I1093588,I1093506,I1093571);
nand I_64181 (I1093059,I1093588,I1093537);
nand I_64182 (I1093056,I1093571,I1093455);
not I_64183 (I1093660,I2514);
DFFARX1 I_64184 (I959929,I2507,I1093660,I1093686,);
and I_64185 (I1093694,I1093686,I959923);
DFFARX1 I_64186 (I1093694,I2507,I1093660,I1093643,);
DFFARX1 I_64187 (I959941,I2507,I1093660,I1093734,);
not I_64188 (I1093742,I959932);
not I_64189 (I1093759,I959944);
nand I_64190 (I1093776,I1093759,I1093742);
nor I_64191 (I1093631,I1093734,I1093776);
DFFARX1 I_64192 (I1093776,I2507,I1093660,I1093816,);
not I_64193 (I1093652,I1093816);
not I_64194 (I1093838,I959950);
nand I_64195 (I1093855,I1093759,I1093838);
DFFARX1 I_64196 (I1093855,I2507,I1093660,I1093881,);
not I_64197 (I1093889,I1093881);
not I_64198 (I1093906,I959926);
nand I_64199 (I1093923,I1093906,I959947);
and I_64200 (I1093940,I1093742,I1093923);
nor I_64201 (I1093957,I1093855,I1093940);
DFFARX1 I_64202 (I1093957,I2507,I1093660,I1093628,);
DFFARX1 I_64203 (I1093940,I2507,I1093660,I1093649,);
nor I_64204 (I1094002,I959926,I959938);
nor I_64205 (I1093640,I1093855,I1094002);
or I_64206 (I1094033,I959926,I959938);
nor I_64207 (I1094050,I959923,I959935);
DFFARX1 I_64208 (I1094050,I2507,I1093660,I1094076,);
not I_64209 (I1094084,I1094076);
nor I_64210 (I1093646,I1094084,I1093889);
nand I_64211 (I1094115,I1094084,I1093734);
not I_64212 (I1094132,I959923);
nand I_64213 (I1094149,I1094132,I1093838);
nand I_64214 (I1094166,I1094084,I1094149);
nand I_64215 (I1093637,I1094166,I1094115);
nand I_64216 (I1093634,I1094149,I1094033);
not I_64217 (I1094238,I2514);
DFFARX1 I_64218 (I8482,I2507,I1094238,I1094264,);
and I_64219 (I1094272,I1094264,I8488);
DFFARX1 I_64220 (I1094272,I2507,I1094238,I1094221,);
DFFARX1 I_64221 (I8467,I2507,I1094238,I1094312,);
not I_64222 (I1094320,I8473);
not I_64223 (I1094337,I8479);
nand I_64224 (I1094354,I1094337,I1094320);
nor I_64225 (I1094209,I1094312,I1094354);
DFFARX1 I_64226 (I1094354,I2507,I1094238,I1094394,);
not I_64227 (I1094230,I1094394);
not I_64228 (I1094416,I8470);
nand I_64229 (I1094433,I1094337,I1094416);
DFFARX1 I_64230 (I1094433,I2507,I1094238,I1094459,);
not I_64231 (I1094467,I1094459);
not I_64232 (I1094484,I8485);
nand I_64233 (I1094501,I1094484,I8470);
and I_64234 (I1094518,I1094320,I1094501);
nor I_64235 (I1094535,I1094433,I1094518);
DFFARX1 I_64236 (I1094535,I2507,I1094238,I1094206,);
DFFARX1 I_64237 (I1094518,I2507,I1094238,I1094227,);
nor I_64238 (I1094580,I8485,I8473);
nor I_64239 (I1094218,I1094433,I1094580);
or I_64240 (I1094611,I8485,I8473);
nor I_64241 (I1094628,I8476,I8467);
DFFARX1 I_64242 (I1094628,I2507,I1094238,I1094654,);
not I_64243 (I1094662,I1094654);
nor I_64244 (I1094224,I1094662,I1094467);
nand I_64245 (I1094693,I1094662,I1094312);
not I_64246 (I1094710,I8476);
nand I_64247 (I1094727,I1094710,I1094416);
nand I_64248 (I1094744,I1094662,I1094727);
nand I_64249 (I1094215,I1094744,I1094693);
nand I_64250 (I1094212,I1094727,I1094611);
not I_64251 (I1094816,I2514);
DFFARX1 I_64252 (I269716,I2507,I1094816,I1094842,);
and I_64253 (I1094850,I1094842,I269701);
DFFARX1 I_64254 (I1094850,I2507,I1094816,I1094799,);
DFFARX1 I_64255 (I269707,I2507,I1094816,I1094890,);
not I_64256 (I1094898,I269689);
not I_64257 (I1094915,I269710);
nand I_64258 (I1094932,I1094915,I1094898);
nor I_64259 (I1094787,I1094890,I1094932);
DFFARX1 I_64260 (I1094932,I2507,I1094816,I1094972,);
not I_64261 (I1094808,I1094972);
not I_64262 (I1094994,I269713);
nand I_64263 (I1095011,I1094915,I1094994);
DFFARX1 I_64264 (I1095011,I2507,I1094816,I1095037,);
not I_64265 (I1095045,I1095037);
not I_64266 (I1095062,I269704);
nand I_64267 (I1095079,I1095062,I269692);
and I_64268 (I1095096,I1094898,I1095079);
nor I_64269 (I1095113,I1095011,I1095096);
DFFARX1 I_64270 (I1095113,I2507,I1094816,I1094784,);
DFFARX1 I_64271 (I1095096,I2507,I1094816,I1094805,);
nor I_64272 (I1095158,I269704,I269698);
nor I_64273 (I1094796,I1095011,I1095158);
or I_64274 (I1095189,I269704,I269698);
nor I_64275 (I1095206,I269695,I269689);
DFFARX1 I_64276 (I1095206,I2507,I1094816,I1095232,);
not I_64277 (I1095240,I1095232);
nor I_64278 (I1094802,I1095240,I1095045);
nand I_64279 (I1095271,I1095240,I1094890);
not I_64280 (I1095288,I269695);
nand I_64281 (I1095305,I1095288,I1094994);
nand I_64282 (I1095322,I1095240,I1095305);
nand I_64283 (I1094793,I1095322,I1095271);
nand I_64284 (I1094790,I1095305,I1095189);
not I_64285 (I1095394,I2514);
DFFARX1 I_64286 (I1275008,I2507,I1095394,I1095420,);
and I_64287 (I1095428,I1095420,I1274990);
DFFARX1 I_64288 (I1095428,I2507,I1095394,I1095377,);
DFFARX1 I_64289 (I1274999,I2507,I1095394,I1095468,);
not I_64290 (I1095476,I1274984);
not I_64291 (I1095493,I1274996);
nand I_64292 (I1095510,I1095493,I1095476);
nor I_64293 (I1095365,I1095468,I1095510);
DFFARX1 I_64294 (I1095510,I2507,I1095394,I1095550,);
not I_64295 (I1095386,I1095550);
not I_64296 (I1095572,I1274987);
nand I_64297 (I1095589,I1095493,I1095572);
DFFARX1 I_64298 (I1095589,I2507,I1095394,I1095615,);
not I_64299 (I1095623,I1095615);
not I_64300 (I1095640,I1274984);
nand I_64301 (I1095657,I1095640,I1274987);
and I_64302 (I1095674,I1095476,I1095657);
nor I_64303 (I1095691,I1095589,I1095674);
DFFARX1 I_64304 (I1095691,I2507,I1095394,I1095362,);
DFFARX1 I_64305 (I1095674,I2507,I1095394,I1095383,);
nor I_64306 (I1095736,I1274984,I1275005);
nor I_64307 (I1095374,I1095589,I1095736);
or I_64308 (I1095767,I1274984,I1275005);
nor I_64309 (I1095784,I1274993,I1275002);
DFFARX1 I_64310 (I1095784,I2507,I1095394,I1095810,);
not I_64311 (I1095818,I1095810);
nor I_64312 (I1095380,I1095818,I1095623);
nand I_64313 (I1095849,I1095818,I1095468);
not I_64314 (I1095866,I1274993);
nand I_64315 (I1095883,I1095866,I1095572);
nand I_64316 (I1095900,I1095818,I1095883);
nand I_64317 (I1095371,I1095900,I1095849);
nand I_64318 (I1095368,I1095883,I1095767);
not I_64319 (I1095972,I2514);
DFFARX1 I_64320 (I1233015,I2507,I1095972,I1095998,);
and I_64321 (I1096006,I1095998,I1233009);
DFFARX1 I_64322 (I1096006,I2507,I1095972,I1095955,);
DFFARX1 I_64323 (I1232994,I2507,I1095972,I1096046,);
not I_64324 (I1096054,I1233000);
not I_64325 (I1096071,I1233012);
nand I_64326 (I1096088,I1096071,I1096054);
nor I_64327 (I1095943,I1096046,I1096088);
DFFARX1 I_64328 (I1096088,I2507,I1095972,I1096128,);
not I_64329 (I1095964,I1096128);
not I_64330 (I1096150,I1232994);
nand I_64331 (I1096167,I1096071,I1096150);
DFFARX1 I_64332 (I1096167,I2507,I1095972,I1096193,);
not I_64333 (I1096201,I1096193);
not I_64334 (I1096218,I1233018);
nand I_64335 (I1096235,I1096218,I1233006);
and I_64336 (I1096252,I1096054,I1096235);
nor I_64337 (I1096269,I1096167,I1096252);
DFFARX1 I_64338 (I1096269,I2507,I1095972,I1095940,);
DFFARX1 I_64339 (I1096252,I2507,I1095972,I1095961,);
nor I_64340 (I1096314,I1233018,I1232997);
nor I_64341 (I1095952,I1096167,I1096314);
or I_64342 (I1096345,I1233018,I1232997);
nor I_64343 (I1096362,I1233003,I1232997);
DFFARX1 I_64344 (I1096362,I2507,I1095972,I1096388,);
not I_64345 (I1096396,I1096388);
nor I_64346 (I1095958,I1096396,I1096201);
nand I_64347 (I1096427,I1096396,I1096046);
not I_64348 (I1096444,I1233003);
nand I_64349 (I1096461,I1096444,I1096150);
nand I_64350 (I1096478,I1096396,I1096461);
nand I_64351 (I1095949,I1096478,I1096427);
nand I_64352 (I1095946,I1096461,I1096345);
not I_64353 (I1096550,I2514);
DFFARX1 I_64354 (I202590,I2507,I1096550,I1096576,);
and I_64355 (I1096584,I1096576,I202593);
DFFARX1 I_64356 (I1096584,I2507,I1096550,I1096533,);
DFFARX1 I_64357 (I202593,I2507,I1096550,I1096624,);
not I_64358 (I1096632,I202608);
not I_64359 (I1096649,I202614);
nand I_64360 (I1096666,I1096649,I1096632);
nor I_64361 (I1096521,I1096624,I1096666);
DFFARX1 I_64362 (I1096666,I2507,I1096550,I1096706,);
not I_64363 (I1096542,I1096706);
not I_64364 (I1096728,I202602);
nand I_64365 (I1096745,I1096649,I1096728);
DFFARX1 I_64366 (I1096745,I2507,I1096550,I1096771,);
not I_64367 (I1096779,I1096771);
not I_64368 (I1096796,I202599);
nand I_64369 (I1096813,I1096796,I202596);
and I_64370 (I1096830,I1096632,I1096813);
nor I_64371 (I1096847,I1096745,I1096830);
DFFARX1 I_64372 (I1096847,I2507,I1096550,I1096518,);
DFFARX1 I_64373 (I1096830,I2507,I1096550,I1096539,);
nor I_64374 (I1096892,I202599,I202590);
nor I_64375 (I1096530,I1096745,I1096892);
or I_64376 (I1096923,I202599,I202590);
nor I_64377 (I1096940,I202605,I202611);
DFFARX1 I_64378 (I1096940,I2507,I1096550,I1096966,);
not I_64379 (I1096974,I1096966);
nor I_64380 (I1096536,I1096974,I1096779);
nand I_64381 (I1097005,I1096974,I1096624);
not I_64382 (I1097022,I202605);
nand I_64383 (I1097039,I1097022,I1096728);
nand I_64384 (I1097056,I1096974,I1097039);
nand I_64385 (I1096527,I1097056,I1097005);
nand I_64386 (I1096524,I1097039,I1096923);
not I_64387 (I1097128,I2514);
DFFARX1 I_64388 (I349820,I2507,I1097128,I1097154,);
and I_64389 (I1097162,I1097154,I349805);
DFFARX1 I_64390 (I1097162,I2507,I1097128,I1097111,);
DFFARX1 I_64391 (I349811,I2507,I1097128,I1097202,);
not I_64392 (I1097210,I349793);
not I_64393 (I1097227,I349814);
nand I_64394 (I1097244,I1097227,I1097210);
nor I_64395 (I1097099,I1097202,I1097244);
DFFARX1 I_64396 (I1097244,I2507,I1097128,I1097284,);
not I_64397 (I1097120,I1097284);
not I_64398 (I1097306,I349817);
nand I_64399 (I1097323,I1097227,I1097306);
DFFARX1 I_64400 (I1097323,I2507,I1097128,I1097349,);
not I_64401 (I1097357,I1097349);
not I_64402 (I1097374,I349808);
nand I_64403 (I1097391,I1097374,I349796);
and I_64404 (I1097408,I1097210,I1097391);
nor I_64405 (I1097425,I1097323,I1097408);
DFFARX1 I_64406 (I1097425,I2507,I1097128,I1097096,);
DFFARX1 I_64407 (I1097408,I2507,I1097128,I1097117,);
nor I_64408 (I1097470,I349808,I349802);
nor I_64409 (I1097108,I1097323,I1097470);
or I_64410 (I1097501,I349808,I349802);
nor I_64411 (I1097518,I349799,I349793);
DFFARX1 I_64412 (I1097518,I2507,I1097128,I1097544,);
not I_64413 (I1097552,I1097544);
nor I_64414 (I1097114,I1097552,I1097357);
nand I_64415 (I1097583,I1097552,I1097202);
not I_64416 (I1097600,I349799);
nand I_64417 (I1097617,I1097600,I1097306);
nand I_64418 (I1097634,I1097552,I1097617);
nand I_64419 (I1097105,I1097634,I1097583);
nand I_64420 (I1097102,I1097617,I1097501);
not I_64421 (I1097706,I2514);
DFFARX1 I_64422 (I155585,I2507,I1097706,I1097732,);
and I_64423 (I1097740,I1097732,I155588);
DFFARX1 I_64424 (I1097740,I2507,I1097706,I1097689,);
DFFARX1 I_64425 (I155588,I2507,I1097706,I1097780,);
not I_64426 (I1097788,I155603);
not I_64427 (I1097805,I155609);
nand I_64428 (I1097822,I1097805,I1097788);
nor I_64429 (I1097677,I1097780,I1097822);
DFFARX1 I_64430 (I1097822,I2507,I1097706,I1097862,);
not I_64431 (I1097698,I1097862);
not I_64432 (I1097884,I155597);
nand I_64433 (I1097901,I1097805,I1097884);
DFFARX1 I_64434 (I1097901,I2507,I1097706,I1097927,);
not I_64435 (I1097935,I1097927);
not I_64436 (I1097952,I155594);
nand I_64437 (I1097969,I1097952,I155591);
and I_64438 (I1097986,I1097788,I1097969);
nor I_64439 (I1098003,I1097901,I1097986);
DFFARX1 I_64440 (I1098003,I2507,I1097706,I1097674,);
DFFARX1 I_64441 (I1097986,I2507,I1097706,I1097695,);
nor I_64442 (I1098048,I155594,I155585);
nor I_64443 (I1097686,I1097901,I1098048);
or I_64444 (I1098079,I155594,I155585);
nor I_64445 (I1098096,I155600,I155606);
DFFARX1 I_64446 (I1098096,I2507,I1097706,I1098122,);
not I_64447 (I1098130,I1098122);
nor I_64448 (I1097692,I1098130,I1097935);
nand I_64449 (I1098161,I1098130,I1097780);
not I_64450 (I1098178,I155600);
nand I_64451 (I1098195,I1098178,I1097884);
nand I_64452 (I1098212,I1098130,I1098195);
nand I_64453 (I1097683,I1098212,I1098161);
nand I_64454 (I1097680,I1098195,I1098079);
not I_64455 (I1098284,I2514);
DFFARX1 I_64456 (I516702,I2507,I1098284,I1098310,);
and I_64457 (I1098318,I1098310,I516717);
DFFARX1 I_64458 (I1098318,I2507,I1098284,I1098267,);
DFFARX1 I_64459 (I516708,I2507,I1098284,I1098358,);
not I_64460 (I1098366,I516702);
not I_64461 (I1098383,I516720);
nand I_64462 (I1098400,I1098383,I1098366);
nor I_64463 (I1098255,I1098358,I1098400);
DFFARX1 I_64464 (I1098400,I2507,I1098284,I1098440,);
not I_64465 (I1098276,I1098440);
not I_64466 (I1098462,I516711);
nand I_64467 (I1098479,I1098383,I1098462);
DFFARX1 I_64468 (I1098479,I2507,I1098284,I1098505,);
not I_64469 (I1098513,I1098505);
not I_64470 (I1098530,I516723);
nand I_64471 (I1098547,I1098530,I516699);
and I_64472 (I1098564,I1098366,I1098547);
nor I_64473 (I1098581,I1098479,I1098564);
DFFARX1 I_64474 (I1098581,I2507,I1098284,I1098252,);
DFFARX1 I_64475 (I1098564,I2507,I1098284,I1098273,);
nor I_64476 (I1098626,I516723,I516699);
nor I_64477 (I1098264,I1098479,I1098626);
or I_64478 (I1098657,I516723,I516699);
nor I_64479 (I1098674,I516705,I516714);
DFFARX1 I_64480 (I1098674,I2507,I1098284,I1098700,);
not I_64481 (I1098708,I1098700);
nor I_64482 (I1098270,I1098708,I1098513);
nand I_64483 (I1098739,I1098708,I1098358);
not I_64484 (I1098756,I516705);
nand I_64485 (I1098773,I1098756,I1098462);
nand I_64486 (I1098790,I1098708,I1098773);
nand I_64487 (I1098261,I1098790,I1098739);
nand I_64488 (I1098258,I1098773,I1098657);
not I_64489 (I1098862,I2514);
DFFARX1 I_64490 (I158560,I2507,I1098862,I1098888,);
and I_64491 (I1098896,I1098888,I158563);
DFFARX1 I_64492 (I1098896,I2507,I1098862,I1098845,);
DFFARX1 I_64493 (I158563,I2507,I1098862,I1098936,);
not I_64494 (I1098944,I158578);
not I_64495 (I1098961,I158584);
nand I_64496 (I1098978,I1098961,I1098944);
nor I_64497 (I1098833,I1098936,I1098978);
DFFARX1 I_64498 (I1098978,I2507,I1098862,I1099018,);
not I_64499 (I1098854,I1099018);
not I_64500 (I1099040,I158572);
nand I_64501 (I1099057,I1098961,I1099040);
DFFARX1 I_64502 (I1099057,I2507,I1098862,I1099083,);
not I_64503 (I1099091,I1099083);
not I_64504 (I1099108,I158569);
nand I_64505 (I1099125,I1099108,I158566);
and I_64506 (I1099142,I1098944,I1099125);
nor I_64507 (I1099159,I1099057,I1099142);
DFFARX1 I_64508 (I1099159,I2507,I1098862,I1098830,);
DFFARX1 I_64509 (I1099142,I2507,I1098862,I1098851,);
nor I_64510 (I1099204,I158569,I158560);
nor I_64511 (I1098842,I1099057,I1099204);
or I_64512 (I1099235,I158569,I158560);
nor I_64513 (I1099252,I158575,I158581);
DFFARX1 I_64514 (I1099252,I2507,I1098862,I1099278,);
not I_64515 (I1099286,I1099278);
nor I_64516 (I1098848,I1099286,I1099091);
nand I_64517 (I1099317,I1099286,I1098936);
not I_64518 (I1099334,I158575);
nand I_64519 (I1099351,I1099334,I1099040);
nand I_64520 (I1099368,I1099286,I1099351);
nand I_64521 (I1098839,I1099368,I1099317);
nand I_64522 (I1098836,I1099351,I1099235);
not I_64523 (I1099440,I2514);
DFFARX1 I_64524 (I799089,I2507,I1099440,I1099466,);
and I_64525 (I1099474,I1099466,I799095);
DFFARX1 I_64526 (I1099474,I2507,I1099440,I1099423,);
DFFARX1 I_64527 (I799101,I2507,I1099440,I1099514,);
not I_64528 (I1099522,I799086);
not I_64529 (I1099539,I799086);
nand I_64530 (I1099556,I1099539,I1099522);
nor I_64531 (I1099411,I1099514,I1099556);
DFFARX1 I_64532 (I1099556,I2507,I1099440,I1099596,);
not I_64533 (I1099432,I1099596);
not I_64534 (I1099618,I799104);
nand I_64535 (I1099635,I1099539,I1099618);
DFFARX1 I_64536 (I1099635,I2507,I1099440,I1099661,);
not I_64537 (I1099669,I1099661);
not I_64538 (I1099686,I799098);
nand I_64539 (I1099703,I1099686,I799089);
and I_64540 (I1099720,I1099522,I1099703);
nor I_64541 (I1099737,I1099635,I1099720);
DFFARX1 I_64542 (I1099737,I2507,I1099440,I1099408,);
DFFARX1 I_64543 (I1099720,I2507,I1099440,I1099429,);
nor I_64544 (I1099782,I799098,I799107);
nor I_64545 (I1099420,I1099635,I1099782);
or I_64546 (I1099813,I799098,I799107);
nor I_64547 (I1099830,I799092,I799092);
DFFARX1 I_64548 (I1099830,I2507,I1099440,I1099856,);
not I_64549 (I1099864,I1099856);
nor I_64550 (I1099426,I1099864,I1099669);
nand I_64551 (I1099895,I1099864,I1099514);
not I_64552 (I1099912,I799092);
nand I_64553 (I1099929,I1099912,I1099618);
nand I_64554 (I1099946,I1099864,I1099929);
nand I_64555 (I1099417,I1099946,I1099895);
nand I_64556 (I1099414,I1099929,I1099813);
not I_64557 (I1100018,I2514);
DFFARX1 I_64558 (I902435,I2507,I1100018,I1100044,);
and I_64559 (I1100052,I1100044,I902429);
DFFARX1 I_64560 (I1100052,I2507,I1100018,I1100001,);
DFFARX1 I_64561 (I902447,I2507,I1100018,I1100092,);
not I_64562 (I1100100,I902438);
not I_64563 (I1100117,I902450);
nand I_64564 (I1100134,I1100117,I1100100);
nor I_64565 (I1099989,I1100092,I1100134);
DFFARX1 I_64566 (I1100134,I2507,I1100018,I1100174,);
not I_64567 (I1100010,I1100174);
not I_64568 (I1100196,I902456);
nand I_64569 (I1100213,I1100117,I1100196);
DFFARX1 I_64570 (I1100213,I2507,I1100018,I1100239,);
not I_64571 (I1100247,I1100239);
not I_64572 (I1100264,I902432);
nand I_64573 (I1100281,I1100264,I902453);
and I_64574 (I1100298,I1100100,I1100281);
nor I_64575 (I1100315,I1100213,I1100298);
DFFARX1 I_64576 (I1100315,I2507,I1100018,I1099986,);
DFFARX1 I_64577 (I1100298,I2507,I1100018,I1100007,);
nor I_64578 (I1100360,I902432,I902444);
nor I_64579 (I1099998,I1100213,I1100360);
or I_64580 (I1100391,I902432,I902444);
nor I_64581 (I1100408,I902429,I902441);
DFFARX1 I_64582 (I1100408,I2507,I1100018,I1100434,);
not I_64583 (I1100442,I1100434);
nor I_64584 (I1100004,I1100442,I1100247);
nand I_64585 (I1100473,I1100442,I1100092);
not I_64586 (I1100490,I902429);
nand I_64587 (I1100507,I1100490,I1100196);
nand I_64588 (I1100524,I1100442,I1100507);
nand I_64589 (I1099995,I1100524,I1100473);
nand I_64590 (I1099992,I1100507,I1100391);
not I_64591 (I1100596,I2514);
DFFARX1 I_64592 (I514917,I2507,I1100596,I1100622,);
and I_64593 (I1100630,I1100622,I514932);
DFFARX1 I_64594 (I1100630,I2507,I1100596,I1100579,);
DFFARX1 I_64595 (I514923,I2507,I1100596,I1100670,);
not I_64596 (I1100678,I514917);
not I_64597 (I1100695,I514935);
nand I_64598 (I1100712,I1100695,I1100678);
nor I_64599 (I1100567,I1100670,I1100712);
DFFARX1 I_64600 (I1100712,I2507,I1100596,I1100752,);
not I_64601 (I1100588,I1100752);
not I_64602 (I1100774,I514926);
nand I_64603 (I1100791,I1100695,I1100774);
DFFARX1 I_64604 (I1100791,I2507,I1100596,I1100817,);
not I_64605 (I1100825,I1100817);
not I_64606 (I1100842,I514938);
nand I_64607 (I1100859,I1100842,I514914);
and I_64608 (I1100876,I1100678,I1100859);
nor I_64609 (I1100893,I1100791,I1100876);
DFFARX1 I_64610 (I1100893,I2507,I1100596,I1100564,);
DFFARX1 I_64611 (I1100876,I2507,I1100596,I1100585,);
nor I_64612 (I1100938,I514938,I514914);
nor I_64613 (I1100576,I1100791,I1100938);
or I_64614 (I1100969,I514938,I514914);
nor I_64615 (I1100986,I514920,I514929);
DFFARX1 I_64616 (I1100986,I2507,I1100596,I1101012,);
not I_64617 (I1101020,I1101012);
nor I_64618 (I1100582,I1101020,I1100825);
nand I_64619 (I1101051,I1101020,I1100670);
not I_64620 (I1101068,I514920);
nand I_64621 (I1101085,I1101068,I1100774);
nand I_64622 (I1101102,I1101020,I1101085);
nand I_64623 (I1100573,I1101102,I1101051);
nand I_64624 (I1100570,I1101085,I1100969);
not I_64625 (I1101174,I2514);
DFFARX1 I_64626 (I979955,I2507,I1101174,I1101200,);
and I_64627 (I1101208,I1101200,I979949);
DFFARX1 I_64628 (I1101208,I2507,I1101174,I1101157,);
DFFARX1 I_64629 (I979967,I2507,I1101174,I1101248,);
not I_64630 (I1101256,I979958);
not I_64631 (I1101273,I979970);
nand I_64632 (I1101290,I1101273,I1101256);
nor I_64633 (I1101145,I1101248,I1101290);
DFFARX1 I_64634 (I1101290,I2507,I1101174,I1101330,);
not I_64635 (I1101166,I1101330);
not I_64636 (I1101352,I979976);
nand I_64637 (I1101369,I1101273,I1101352);
DFFARX1 I_64638 (I1101369,I2507,I1101174,I1101395,);
not I_64639 (I1101403,I1101395);
not I_64640 (I1101420,I979952);
nand I_64641 (I1101437,I1101420,I979973);
and I_64642 (I1101454,I1101256,I1101437);
nor I_64643 (I1101471,I1101369,I1101454);
DFFARX1 I_64644 (I1101471,I2507,I1101174,I1101142,);
DFFARX1 I_64645 (I1101454,I2507,I1101174,I1101163,);
nor I_64646 (I1101516,I979952,I979964);
nor I_64647 (I1101154,I1101369,I1101516);
or I_64648 (I1101547,I979952,I979964);
nor I_64649 (I1101564,I979949,I979961);
DFFARX1 I_64650 (I1101564,I2507,I1101174,I1101590,);
not I_64651 (I1101598,I1101590);
nor I_64652 (I1101160,I1101598,I1101403);
nand I_64653 (I1101629,I1101598,I1101248);
not I_64654 (I1101646,I979949);
nand I_64655 (I1101663,I1101646,I1101352);
nand I_64656 (I1101680,I1101598,I1101663);
nand I_64657 (I1101151,I1101680,I1101629);
nand I_64658 (I1101148,I1101663,I1101547);
not I_64659 (I1101752,I2514);
DFFARX1 I_64660 (I429455,I2507,I1101752,I1101778,);
and I_64661 (I1101786,I1101778,I429470);
DFFARX1 I_64662 (I1101786,I2507,I1101752,I1101735,);
DFFARX1 I_64663 (I429473,I2507,I1101752,I1101826,);
not I_64664 (I1101834,I429467);
not I_64665 (I1101851,I429482);
nand I_64666 (I1101868,I1101851,I1101834);
nor I_64667 (I1101723,I1101826,I1101868);
DFFARX1 I_64668 (I1101868,I2507,I1101752,I1101908,);
not I_64669 (I1101744,I1101908);
not I_64670 (I1101930,I429458);
nand I_64671 (I1101947,I1101851,I1101930);
DFFARX1 I_64672 (I1101947,I2507,I1101752,I1101973,);
not I_64673 (I1101981,I1101973);
not I_64674 (I1101998,I429461);
nand I_64675 (I1102015,I1101998,I429455);
and I_64676 (I1102032,I1101834,I1102015);
nor I_64677 (I1102049,I1101947,I1102032);
DFFARX1 I_64678 (I1102049,I2507,I1101752,I1101720,);
DFFARX1 I_64679 (I1102032,I2507,I1101752,I1101741,);
nor I_64680 (I1102094,I429461,I429464);
nor I_64681 (I1101732,I1101947,I1102094);
or I_64682 (I1102125,I429461,I429464);
nor I_64683 (I1102142,I429479,I429476);
DFFARX1 I_64684 (I1102142,I2507,I1101752,I1102168,);
not I_64685 (I1102176,I1102168);
nor I_64686 (I1101738,I1102176,I1101981);
nand I_64687 (I1102207,I1102176,I1101826);
not I_64688 (I1102224,I429479);
nand I_64689 (I1102241,I1102224,I1101930);
nand I_64690 (I1102258,I1102176,I1102241);
nand I_64691 (I1101729,I1102258,I1102207);
nand I_64692 (I1101726,I1102241,I1102125);
not I_64693 (I1102330,I2514);
DFFARX1 I_64694 (I563107,I2507,I1102330,I1102356,);
and I_64695 (I1102364,I1102356,I563095);
DFFARX1 I_64696 (I1102364,I2507,I1102330,I1102313,);
DFFARX1 I_64697 (I563110,I2507,I1102330,I1102404,);
not I_64698 (I1102412,I563101);
not I_64699 (I1102429,I563092);
nand I_64700 (I1102446,I1102429,I1102412);
nor I_64701 (I1102301,I1102404,I1102446);
DFFARX1 I_64702 (I1102446,I2507,I1102330,I1102486,);
not I_64703 (I1102322,I1102486);
not I_64704 (I1102508,I563098);
nand I_64705 (I1102525,I1102429,I1102508);
DFFARX1 I_64706 (I1102525,I2507,I1102330,I1102551,);
not I_64707 (I1102559,I1102551);
not I_64708 (I1102576,I563113);
nand I_64709 (I1102593,I1102576,I563116);
and I_64710 (I1102610,I1102412,I1102593);
nor I_64711 (I1102627,I1102525,I1102610);
DFFARX1 I_64712 (I1102627,I2507,I1102330,I1102298,);
DFFARX1 I_64713 (I1102610,I2507,I1102330,I1102319,);
nor I_64714 (I1102672,I563113,I563092);
nor I_64715 (I1102310,I1102525,I1102672);
or I_64716 (I1102703,I563113,I563092);
nor I_64717 (I1102720,I563104,I563095);
DFFARX1 I_64718 (I1102720,I2507,I1102330,I1102746,);
not I_64719 (I1102754,I1102746);
nor I_64720 (I1102316,I1102754,I1102559);
nand I_64721 (I1102785,I1102754,I1102404);
not I_64722 (I1102802,I563104);
nand I_64723 (I1102819,I1102802,I1102508);
nand I_64724 (I1102836,I1102754,I1102819);
nand I_64725 (I1102307,I1102836,I1102785);
nand I_64726 (I1102304,I1102819,I1102703);
not I_64727 (I1102908,I2514);
DFFARX1 I_64728 (I372481,I2507,I1102908,I1102934,);
and I_64729 (I1102942,I1102934,I372466);
DFFARX1 I_64730 (I1102942,I2507,I1102908,I1102891,);
DFFARX1 I_64731 (I372472,I2507,I1102908,I1102982,);
not I_64732 (I1102990,I372454);
not I_64733 (I1103007,I372475);
nand I_64734 (I1103024,I1103007,I1102990);
nor I_64735 (I1102879,I1102982,I1103024);
DFFARX1 I_64736 (I1103024,I2507,I1102908,I1103064,);
not I_64737 (I1102900,I1103064);
not I_64738 (I1103086,I372478);
nand I_64739 (I1103103,I1103007,I1103086);
DFFARX1 I_64740 (I1103103,I2507,I1102908,I1103129,);
not I_64741 (I1103137,I1103129);
not I_64742 (I1103154,I372469);
nand I_64743 (I1103171,I1103154,I372457);
and I_64744 (I1103188,I1102990,I1103171);
nor I_64745 (I1103205,I1103103,I1103188);
DFFARX1 I_64746 (I1103205,I2507,I1102908,I1102876,);
DFFARX1 I_64747 (I1103188,I2507,I1102908,I1102897,);
nor I_64748 (I1103250,I372469,I372463);
nor I_64749 (I1102888,I1103103,I1103250);
or I_64750 (I1103281,I372469,I372463);
nor I_64751 (I1103298,I372460,I372454);
DFFARX1 I_64752 (I1103298,I2507,I1102908,I1103324,);
not I_64753 (I1103332,I1103324);
nor I_64754 (I1102894,I1103332,I1103137);
nand I_64755 (I1103363,I1103332,I1102982);
not I_64756 (I1103380,I372460);
nand I_64757 (I1103397,I1103380,I1103086);
nand I_64758 (I1103414,I1103332,I1103397);
nand I_64759 (I1102885,I1103414,I1103363);
nand I_64760 (I1102882,I1103397,I1103281);
not I_64761 (I1103486,I2514);
DFFARX1 I_64762 (I869707,I2507,I1103486,I1103512,);
and I_64763 (I1103520,I1103512,I869713);
DFFARX1 I_64764 (I1103520,I2507,I1103486,I1103469,);
DFFARX1 I_64765 (I869719,I2507,I1103486,I1103560,);
not I_64766 (I1103568,I869704);
not I_64767 (I1103585,I869704);
nand I_64768 (I1103602,I1103585,I1103568);
nor I_64769 (I1103457,I1103560,I1103602);
DFFARX1 I_64770 (I1103602,I2507,I1103486,I1103642,);
not I_64771 (I1103478,I1103642);
not I_64772 (I1103664,I869722);
nand I_64773 (I1103681,I1103585,I1103664);
DFFARX1 I_64774 (I1103681,I2507,I1103486,I1103707,);
not I_64775 (I1103715,I1103707);
not I_64776 (I1103732,I869716);
nand I_64777 (I1103749,I1103732,I869707);
and I_64778 (I1103766,I1103568,I1103749);
nor I_64779 (I1103783,I1103681,I1103766);
DFFARX1 I_64780 (I1103783,I2507,I1103486,I1103454,);
DFFARX1 I_64781 (I1103766,I2507,I1103486,I1103475,);
nor I_64782 (I1103828,I869716,I869725);
nor I_64783 (I1103466,I1103681,I1103828);
or I_64784 (I1103859,I869716,I869725);
nor I_64785 (I1103876,I869710,I869710);
DFFARX1 I_64786 (I1103876,I2507,I1103486,I1103902,);
not I_64787 (I1103910,I1103902);
nor I_64788 (I1103472,I1103910,I1103715);
nand I_64789 (I1103941,I1103910,I1103560);
not I_64790 (I1103958,I869710);
nand I_64791 (I1103975,I1103958,I1103664);
nand I_64792 (I1103992,I1103910,I1103975);
nand I_64793 (I1103463,I1103992,I1103941);
nand I_64794 (I1103460,I1103975,I1103859);
not I_64795 (I1104064,I2514);
DFFARX1 I_64796 (I371427,I2507,I1104064,I1104090,);
and I_64797 (I1104098,I1104090,I371412);
DFFARX1 I_64798 (I1104098,I2507,I1104064,I1104047,);
DFFARX1 I_64799 (I371418,I2507,I1104064,I1104138,);
not I_64800 (I1104146,I371400);
not I_64801 (I1104163,I371421);
nand I_64802 (I1104180,I1104163,I1104146);
nor I_64803 (I1104035,I1104138,I1104180);
DFFARX1 I_64804 (I1104180,I2507,I1104064,I1104220,);
not I_64805 (I1104056,I1104220);
not I_64806 (I1104242,I371424);
nand I_64807 (I1104259,I1104163,I1104242);
DFFARX1 I_64808 (I1104259,I2507,I1104064,I1104285,);
not I_64809 (I1104293,I1104285);
not I_64810 (I1104310,I371415);
nand I_64811 (I1104327,I1104310,I371403);
and I_64812 (I1104344,I1104146,I1104327);
nor I_64813 (I1104361,I1104259,I1104344);
DFFARX1 I_64814 (I1104361,I2507,I1104064,I1104032,);
DFFARX1 I_64815 (I1104344,I2507,I1104064,I1104053,);
nor I_64816 (I1104406,I371415,I371409);
nor I_64817 (I1104044,I1104259,I1104406);
or I_64818 (I1104437,I371415,I371409);
nor I_64819 (I1104454,I371406,I371400);
DFFARX1 I_64820 (I1104454,I2507,I1104064,I1104480,);
not I_64821 (I1104488,I1104480);
nor I_64822 (I1104050,I1104488,I1104293);
nand I_64823 (I1104519,I1104488,I1104138);
not I_64824 (I1104536,I371406);
nand I_64825 (I1104553,I1104536,I1104242);
nand I_64826 (I1104570,I1104488,I1104553);
nand I_64827 (I1104041,I1104570,I1104519);
nand I_64828 (I1104038,I1104553,I1104437);
not I_64829 (I1104642,I2514);
DFFARX1 I_64830 (I1291192,I2507,I1104642,I1104668,);
and I_64831 (I1104676,I1104668,I1291174);
DFFARX1 I_64832 (I1104676,I2507,I1104642,I1104625,);
DFFARX1 I_64833 (I1291183,I2507,I1104642,I1104716,);
not I_64834 (I1104724,I1291168);
not I_64835 (I1104741,I1291180);
nand I_64836 (I1104758,I1104741,I1104724);
nor I_64837 (I1104613,I1104716,I1104758);
DFFARX1 I_64838 (I1104758,I2507,I1104642,I1104798,);
not I_64839 (I1104634,I1104798);
not I_64840 (I1104820,I1291171);
nand I_64841 (I1104837,I1104741,I1104820);
DFFARX1 I_64842 (I1104837,I2507,I1104642,I1104863,);
not I_64843 (I1104871,I1104863);
not I_64844 (I1104888,I1291168);
nand I_64845 (I1104905,I1104888,I1291171);
and I_64846 (I1104922,I1104724,I1104905);
nor I_64847 (I1104939,I1104837,I1104922);
DFFARX1 I_64848 (I1104939,I2507,I1104642,I1104610,);
DFFARX1 I_64849 (I1104922,I2507,I1104642,I1104631,);
nor I_64850 (I1104984,I1291168,I1291189);
nor I_64851 (I1104622,I1104837,I1104984);
or I_64852 (I1105015,I1291168,I1291189);
nor I_64853 (I1105032,I1291177,I1291186);
DFFARX1 I_64854 (I1105032,I2507,I1104642,I1105058,);
not I_64855 (I1105066,I1105058);
nor I_64856 (I1104628,I1105066,I1104871);
nand I_64857 (I1105097,I1105066,I1104716);
not I_64858 (I1105114,I1291177);
nand I_64859 (I1105131,I1105114,I1104820);
nand I_64860 (I1105148,I1105066,I1105131);
nand I_64861 (I1104619,I1105148,I1105097);
nand I_64862 (I1104616,I1105131,I1105015);
not I_64863 (I1105220,I2514);
DFFARX1 I_64864 (I34834,I2507,I1105220,I1105246,);
and I_64865 (I1105254,I1105246,I34837);
DFFARX1 I_64866 (I1105254,I2507,I1105220,I1105203,);
DFFARX1 I_64867 (I34837,I2507,I1105220,I1105294,);
not I_64868 (I1105302,I34840);
not I_64869 (I1105319,I34855);
nand I_64870 (I1105336,I1105319,I1105302);
nor I_64871 (I1105191,I1105294,I1105336);
DFFARX1 I_64872 (I1105336,I2507,I1105220,I1105376,);
not I_64873 (I1105212,I1105376);
not I_64874 (I1105398,I34849);
nand I_64875 (I1105415,I1105319,I1105398);
DFFARX1 I_64876 (I1105415,I2507,I1105220,I1105441,);
not I_64877 (I1105449,I1105441);
not I_64878 (I1105466,I34852);
nand I_64879 (I1105483,I1105466,I34834);
and I_64880 (I1105500,I1105302,I1105483);
nor I_64881 (I1105517,I1105415,I1105500);
DFFARX1 I_64882 (I1105517,I2507,I1105220,I1105188,);
DFFARX1 I_64883 (I1105500,I2507,I1105220,I1105209,);
nor I_64884 (I1105562,I34852,I34846);
nor I_64885 (I1105200,I1105415,I1105562);
or I_64886 (I1105593,I34852,I34846);
nor I_64887 (I1105610,I34843,I34858);
DFFARX1 I_64888 (I1105610,I2507,I1105220,I1105636,);
not I_64889 (I1105644,I1105636);
nor I_64890 (I1105206,I1105644,I1105449);
nand I_64891 (I1105675,I1105644,I1105294);
not I_64892 (I1105692,I34843);
nand I_64893 (I1105709,I1105692,I1105398);
nand I_64894 (I1105726,I1105644,I1105709);
nand I_64895 (I1105197,I1105726,I1105675);
nand I_64896 (I1105194,I1105709,I1105593);
not I_64897 (I1105798,I2514);
DFFARX1 I_64898 (I626109,I2507,I1105798,I1105824,);
and I_64899 (I1105832,I1105824,I626097);
DFFARX1 I_64900 (I1105832,I2507,I1105798,I1105781,);
DFFARX1 I_64901 (I626112,I2507,I1105798,I1105872,);
not I_64902 (I1105880,I626103);
not I_64903 (I1105897,I626094);
nand I_64904 (I1105914,I1105897,I1105880);
nor I_64905 (I1105769,I1105872,I1105914);
DFFARX1 I_64906 (I1105914,I2507,I1105798,I1105954,);
not I_64907 (I1105790,I1105954);
not I_64908 (I1105976,I626100);
nand I_64909 (I1105993,I1105897,I1105976);
DFFARX1 I_64910 (I1105993,I2507,I1105798,I1106019,);
not I_64911 (I1106027,I1106019);
not I_64912 (I1106044,I626115);
nand I_64913 (I1106061,I1106044,I626118);
and I_64914 (I1106078,I1105880,I1106061);
nor I_64915 (I1106095,I1105993,I1106078);
DFFARX1 I_64916 (I1106095,I2507,I1105798,I1105766,);
DFFARX1 I_64917 (I1106078,I2507,I1105798,I1105787,);
nor I_64918 (I1106140,I626115,I626094);
nor I_64919 (I1105778,I1105993,I1106140);
or I_64920 (I1106171,I626115,I626094);
nor I_64921 (I1106188,I626106,I626097);
DFFARX1 I_64922 (I1106188,I2507,I1105798,I1106214,);
not I_64923 (I1106222,I1106214);
nor I_64924 (I1105784,I1106222,I1106027);
nand I_64925 (I1106253,I1106222,I1105872);
not I_64926 (I1106270,I626106);
nand I_64927 (I1106287,I1106270,I1105976);
nand I_64928 (I1106304,I1106222,I1106287);
nand I_64929 (I1105775,I1106304,I1106253);
nand I_64930 (I1105772,I1106287,I1106171);
not I_64931 (I1106376,I2514);
DFFARX1 I_64932 (I403343,I2507,I1106376,I1106402,);
and I_64933 (I1106410,I1106402,I403358);
DFFARX1 I_64934 (I1106410,I2507,I1106376,I1106359,);
DFFARX1 I_64935 (I403361,I2507,I1106376,I1106450,);
not I_64936 (I1106458,I403355);
not I_64937 (I1106475,I403370);
nand I_64938 (I1106492,I1106475,I1106458);
nor I_64939 (I1106347,I1106450,I1106492);
DFFARX1 I_64940 (I1106492,I2507,I1106376,I1106532,);
not I_64941 (I1106368,I1106532);
not I_64942 (I1106554,I403346);
nand I_64943 (I1106571,I1106475,I1106554);
DFFARX1 I_64944 (I1106571,I2507,I1106376,I1106597,);
not I_64945 (I1106605,I1106597);
not I_64946 (I1106622,I403349);
nand I_64947 (I1106639,I1106622,I403343);
and I_64948 (I1106656,I1106458,I1106639);
nor I_64949 (I1106673,I1106571,I1106656);
DFFARX1 I_64950 (I1106673,I2507,I1106376,I1106344,);
DFFARX1 I_64951 (I1106656,I2507,I1106376,I1106365,);
nor I_64952 (I1106718,I403349,I403352);
nor I_64953 (I1106356,I1106571,I1106718);
or I_64954 (I1106749,I403349,I403352);
nor I_64955 (I1106766,I403367,I403364);
DFFARX1 I_64956 (I1106766,I2507,I1106376,I1106792,);
not I_64957 (I1106800,I1106792);
nor I_64958 (I1106362,I1106800,I1106605);
nand I_64959 (I1106831,I1106800,I1106450);
not I_64960 (I1106848,I403367);
nand I_64961 (I1106865,I1106848,I1106554);
nand I_64962 (I1106882,I1106800,I1106865);
nand I_64963 (I1106353,I1106882,I1106831);
nand I_64964 (I1106350,I1106865,I1106749);
not I_64965 (I1106954,I2514);
DFFARX1 I_64966 (I660211,I2507,I1106954,I1106980,);
and I_64967 (I1106988,I1106980,I660199);
DFFARX1 I_64968 (I1106988,I2507,I1106954,I1106937,);
DFFARX1 I_64969 (I660202,I2507,I1106954,I1107028,);
not I_64970 (I1107036,I660196);
not I_64971 (I1107053,I660220);
nand I_64972 (I1107070,I1107053,I1107036);
nor I_64973 (I1106925,I1107028,I1107070);
DFFARX1 I_64974 (I1107070,I2507,I1106954,I1107110,);
not I_64975 (I1106946,I1107110);
not I_64976 (I1107132,I660208);
nand I_64977 (I1107149,I1107053,I1107132);
DFFARX1 I_64978 (I1107149,I2507,I1106954,I1107175,);
not I_64979 (I1107183,I1107175);
not I_64980 (I1107200,I660217);
nand I_64981 (I1107217,I1107200,I660214);
and I_64982 (I1107234,I1107036,I1107217);
nor I_64983 (I1107251,I1107149,I1107234);
DFFARX1 I_64984 (I1107251,I2507,I1106954,I1106922,);
DFFARX1 I_64985 (I1107234,I2507,I1106954,I1106943,);
nor I_64986 (I1107296,I660217,I660205);
nor I_64987 (I1106934,I1107149,I1107296);
or I_64988 (I1107327,I660217,I660205);
nor I_64989 (I1107344,I660196,I660199);
DFFARX1 I_64990 (I1107344,I2507,I1106954,I1107370,);
not I_64991 (I1107378,I1107370);
nor I_64992 (I1106940,I1107378,I1107183);
nand I_64993 (I1107409,I1107378,I1107028);
not I_64994 (I1107426,I660196);
nand I_64995 (I1107443,I1107426,I1107132);
nand I_64996 (I1107460,I1107378,I1107443);
nand I_64997 (I1106931,I1107460,I1107409);
nand I_64998 (I1106928,I1107443,I1107327);
not I_64999 (I1107532,I2514);
DFFARX1 I_65000 (I1240631,I2507,I1107532,I1107558,);
and I_65001 (I1107566,I1107558,I1240625);
DFFARX1 I_65002 (I1107566,I2507,I1107532,I1107515,);
DFFARX1 I_65003 (I1240610,I2507,I1107532,I1107606,);
not I_65004 (I1107614,I1240616);
not I_65005 (I1107631,I1240628);
nand I_65006 (I1107648,I1107631,I1107614);
nor I_65007 (I1107503,I1107606,I1107648);
DFFARX1 I_65008 (I1107648,I2507,I1107532,I1107688,);
not I_65009 (I1107524,I1107688);
not I_65010 (I1107710,I1240610);
nand I_65011 (I1107727,I1107631,I1107710);
DFFARX1 I_65012 (I1107727,I2507,I1107532,I1107753,);
not I_65013 (I1107761,I1107753);
not I_65014 (I1107778,I1240634);
nand I_65015 (I1107795,I1107778,I1240622);
and I_65016 (I1107812,I1107614,I1107795);
nor I_65017 (I1107829,I1107727,I1107812);
DFFARX1 I_65018 (I1107829,I2507,I1107532,I1107500,);
DFFARX1 I_65019 (I1107812,I2507,I1107532,I1107521,);
nor I_65020 (I1107874,I1240634,I1240613);
nor I_65021 (I1107512,I1107727,I1107874);
or I_65022 (I1107905,I1240634,I1240613);
nor I_65023 (I1107922,I1240619,I1240613);
DFFARX1 I_65024 (I1107922,I2507,I1107532,I1107948,);
not I_65025 (I1107956,I1107948);
nor I_65026 (I1107518,I1107956,I1107761);
nand I_65027 (I1107987,I1107956,I1107606);
not I_65028 (I1108004,I1240619);
nand I_65029 (I1108021,I1108004,I1107710);
nand I_65030 (I1108038,I1107956,I1108021);
nand I_65031 (I1107509,I1108038,I1107987);
nand I_65032 (I1107506,I1108021,I1107905);
not I_65033 (I1108110,I2514);
DFFARX1 I_65034 (I709341,I2507,I1108110,I1108136,);
and I_65035 (I1108144,I1108136,I709329);
DFFARX1 I_65036 (I1108144,I2507,I1108110,I1108093,);
DFFARX1 I_65037 (I709332,I2507,I1108110,I1108184,);
not I_65038 (I1108192,I709326);
not I_65039 (I1108209,I709350);
nand I_65040 (I1108226,I1108209,I1108192);
nor I_65041 (I1108081,I1108184,I1108226);
DFFARX1 I_65042 (I1108226,I2507,I1108110,I1108266,);
not I_65043 (I1108102,I1108266);
not I_65044 (I1108288,I709338);
nand I_65045 (I1108305,I1108209,I1108288);
DFFARX1 I_65046 (I1108305,I2507,I1108110,I1108331,);
not I_65047 (I1108339,I1108331);
not I_65048 (I1108356,I709347);
nand I_65049 (I1108373,I1108356,I709344);
and I_65050 (I1108390,I1108192,I1108373);
nor I_65051 (I1108407,I1108305,I1108390);
DFFARX1 I_65052 (I1108407,I2507,I1108110,I1108078,);
DFFARX1 I_65053 (I1108390,I2507,I1108110,I1108099,);
nor I_65054 (I1108452,I709347,I709335);
nor I_65055 (I1108090,I1108305,I1108452);
or I_65056 (I1108483,I709347,I709335);
nor I_65057 (I1108500,I709326,I709329);
DFFARX1 I_65058 (I1108500,I2507,I1108110,I1108526,);
not I_65059 (I1108534,I1108526);
nor I_65060 (I1108096,I1108534,I1108339);
nand I_65061 (I1108565,I1108534,I1108184);
not I_65062 (I1108582,I709326);
nand I_65063 (I1108599,I1108582,I1108288);
nand I_65064 (I1108616,I1108534,I1108599);
nand I_65065 (I1108087,I1108616,I1108565);
nand I_65066 (I1108084,I1108599,I1108483);
not I_65067 (I1108688,I2514);
DFFARX1 I_65068 (I950885,I2507,I1108688,I1108714,);
and I_65069 (I1108722,I1108714,I950879);
DFFARX1 I_65070 (I1108722,I2507,I1108688,I1108671,);
DFFARX1 I_65071 (I950897,I2507,I1108688,I1108762,);
not I_65072 (I1108770,I950888);
not I_65073 (I1108787,I950900);
nand I_65074 (I1108804,I1108787,I1108770);
nor I_65075 (I1108659,I1108762,I1108804);
DFFARX1 I_65076 (I1108804,I2507,I1108688,I1108844,);
not I_65077 (I1108680,I1108844);
not I_65078 (I1108866,I950906);
nand I_65079 (I1108883,I1108787,I1108866);
DFFARX1 I_65080 (I1108883,I2507,I1108688,I1108909,);
not I_65081 (I1108917,I1108909);
not I_65082 (I1108934,I950882);
nand I_65083 (I1108951,I1108934,I950903);
and I_65084 (I1108968,I1108770,I1108951);
nor I_65085 (I1108985,I1108883,I1108968);
DFFARX1 I_65086 (I1108985,I2507,I1108688,I1108656,);
DFFARX1 I_65087 (I1108968,I2507,I1108688,I1108677,);
nor I_65088 (I1109030,I950882,I950894);
nor I_65089 (I1108668,I1108883,I1109030);
or I_65090 (I1109061,I950882,I950894);
nor I_65091 (I1109078,I950879,I950891);
DFFARX1 I_65092 (I1109078,I2507,I1108688,I1109104,);
not I_65093 (I1109112,I1109104);
nor I_65094 (I1108674,I1109112,I1108917);
nand I_65095 (I1109143,I1109112,I1108762);
not I_65096 (I1109160,I950879);
nand I_65097 (I1109177,I1109160,I1108866);
nand I_65098 (I1109194,I1109112,I1109177);
nand I_65099 (I1108665,I1109194,I1109143);
nand I_65100 (I1108662,I1109177,I1109061);
not I_65101 (I1109266,I2514);
DFFARX1 I_65102 (I860221,I2507,I1109266,I1109292,);
and I_65103 (I1109300,I1109292,I860227);
DFFARX1 I_65104 (I1109300,I2507,I1109266,I1109249,);
DFFARX1 I_65105 (I860233,I2507,I1109266,I1109340,);
not I_65106 (I1109348,I860218);
not I_65107 (I1109365,I860218);
nand I_65108 (I1109382,I1109365,I1109348);
nor I_65109 (I1109237,I1109340,I1109382);
DFFARX1 I_65110 (I1109382,I2507,I1109266,I1109422,);
not I_65111 (I1109258,I1109422);
not I_65112 (I1109444,I860236);
nand I_65113 (I1109461,I1109365,I1109444);
DFFARX1 I_65114 (I1109461,I2507,I1109266,I1109487,);
not I_65115 (I1109495,I1109487);
not I_65116 (I1109512,I860230);
nand I_65117 (I1109529,I1109512,I860221);
and I_65118 (I1109546,I1109348,I1109529);
nor I_65119 (I1109563,I1109461,I1109546);
DFFARX1 I_65120 (I1109563,I2507,I1109266,I1109234,);
DFFARX1 I_65121 (I1109546,I2507,I1109266,I1109255,);
nor I_65122 (I1109608,I860230,I860239);
nor I_65123 (I1109246,I1109461,I1109608);
or I_65124 (I1109639,I860230,I860239);
nor I_65125 (I1109656,I860224,I860224);
DFFARX1 I_65126 (I1109656,I2507,I1109266,I1109682,);
not I_65127 (I1109690,I1109682);
nor I_65128 (I1109252,I1109690,I1109495);
nand I_65129 (I1109721,I1109690,I1109340);
not I_65130 (I1109738,I860224);
nand I_65131 (I1109755,I1109738,I1109444);
nand I_65132 (I1109772,I1109690,I1109755);
nand I_65133 (I1109243,I1109772,I1109721);
nand I_65134 (I1109240,I1109755,I1109639);
not I_65135 (I1109844,I2514);
DFFARX1 I_65136 (I780644,I2507,I1109844,I1109870,);
and I_65137 (I1109878,I1109870,I780650);
DFFARX1 I_65138 (I1109878,I2507,I1109844,I1109827,);
DFFARX1 I_65139 (I780656,I2507,I1109844,I1109918,);
not I_65140 (I1109926,I780641);
not I_65141 (I1109943,I780641);
nand I_65142 (I1109960,I1109943,I1109926);
nor I_65143 (I1109815,I1109918,I1109960);
DFFARX1 I_65144 (I1109960,I2507,I1109844,I1110000,);
not I_65145 (I1109836,I1110000);
not I_65146 (I1110022,I780659);
nand I_65147 (I1110039,I1109943,I1110022);
DFFARX1 I_65148 (I1110039,I2507,I1109844,I1110065,);
not I_65149 (I1110073,I1110065);
not I_65150 (I1110090,I780653);
nand I_65151 (I1110107,I1110090,I780644);
and I_65152 (I1110124,I1109926,I1110107);
nor I_65153 (I1110141,I1110039,I1110124);
DFFARX1 I_65154 (I1110141,I2507,I1109844,I1109812,);
DFFARX1 I_65155 (I1110124,I2507,I1109844,I1109833,);
nor I_65156 (I1110186,I780653,I780662);
nor I_65157 (I1109824,I1110039,I1110186);
or I_65158 (I1110217,I780653,I780662);
nor I_65159 (I1110234,I780647,I780647);
DFFARX1 I_65160 (I1110234,I2507,I1109844,I1110260,);
not I_65161 (I1110268,I1110260);
nor I_65162 (I1109830,I1110268,I1110073);
nand I_65163 (I1110299,I1110268,I1109918);
not I_65164 (I1110316,I780647);
nand I_65165 (I1110333,I1110316,I1110022);
nand I_65166 (I1110350,I1110268,I1110333);
nand I_65167 (I1109821,I1110350,I1110299);
nand I_65168 (I1109818,I1110333,I1110217);
not I_65169 (I1110422,I2514);
DFFARX1 I_65170 (I1338659,I2507,I1110422,I1110448,);
and I_65171 (I1110456,I1110448,I1338641);
DFFARX1 I_65172 (I1110456,I2507,I1110422,I1110405,);
DFFARX1 I_65173 (I1338632,I2507,I1110422,I1110496,);
not I_65174 (I1110504,I1338647);
not I_65175 (I1110521,I1338635);
nand I_65176 (I1110538,I1110521,I1110504);
nor I_65177 (I1110393,I1110496,I1110538);
DFFARX1 I_65178 (I1110538,I2507,I1110422,I1110578,);
not I_65179 (I1110414,I1110578);
not I_65180 (I1110600,I1338644);
nand I_65181 (I1110617,I1110521,I1110600);
DFFARX1 I_65182 (I1110617,I2507,I1110422,I1110643,);
not I_65183 (I1110651,I1110643);
not I_65184 (I1110668,I1338653);
nand I_65185 (I1110685,I1110668,I1338632);
and I_65186 (I1110702,I1110504,I1110685);
nor I_65187 (I1110719,I1110617,I1110702);
DFFARX1 I_65188 (I1110719,I2507,I1110422,I1110390,);
DFFARX1 I_65189 (I1110702,I2507,I1110422,I1110411,);
nor I_65190 (I1110764,I1338653,I1338656);
nor I_65191 (I1110402,I1110617,I1110764);
or I_65192 (I1110795,I1338653,I1338656);
nor I_65193 (I1110812,I1338650,I1338638);
DFFARX1 I_65194 (I1110812,I2507,I1110422,I1110838,);
not I_65195 (I1110846,I1110838);
nor I_65196 (I1110408,I1110846,I1110651);
nand I_65197 (I1110877,I1110846,I1110496);
not I_65198 (I1110894,I1338650);
nand I_65199 (I1110911,I1110894,I1110600);
nand I_65200 (I1110928,I1110846,I1110911);
nand I_65201 (I1110399,I1110928,I1110877);
nand I_65202 (I1110396,I1110911,I1110795);
not I_65203 (I1111000,I2514);
DFFARX1 I_65204 (I1324974,I2507,I1111000,I1111026,);
and I_65205 (I1111034,I1111026,I1324956);
DFFARX1 I_65206 (I1111034,I2507,I1111000,I1110983,);
DFFARX1 I_65207 (I1324947,I2507,I1111000,I1111074,);
not I_65208 (I1111082,I1324962);
not I_65209 (I1111099,I1324950);
nand I_65210 (I1111116,I1111099,I1111082);
nor I_65211 (I1110971,I1111074,I1111116);
DFFARX1 I_65212 (I1111116,I2507,I1111000,I1111156,);
not I_65213 (I1110992,I1111156);
not I_65214 (I1111178,I1324959);
nand I_65215 (I1111195,I1111099,I1111178);
DFFARX1 I_65216 (I1111195,I2507,I1111000,I1111221,);
not I_65217 (I1111229,I1111221);
not I_65218 (I1111246,I1324968);
nand I_65219 (I1111263,I1111246,I1324947);
and I_65220 (I1111280,I1111082,I1111263);
nor I_65221 (I1111297,I1111195,I1111280);
DFFARX1 I_65222 (I1111297,I2507,I1111000,I1110968,);
DFFARX1 I_65223 (I1111280,I2507,I1111000,I1110989,);
nor I_65224 (I1111342,I1324968,I1324971);
nor I_65225 (I1110980,I1111195,I1111342);
or I_65226 (I1111373,I1324968,I1324971);
nor I_65227 (I1111390,I1324965,I1324953);
DFFARX1 I_65228 (I1111390,I2507,I1111000,I1111416,);
not I_65229 (I1111424,I1111416);
nor I_65230 (I1110986,I1111424,I1111229);
nand I_65231 (I1111455,I1111424,I1111074);
not I_65232 (I1111472,I1324965);
nand I_65233 (I1111489,I1111472,I1111178);
nand I_65234 (I1111506,I1111424,I1111489);
nand I_65235 (I1110977,I1111506,I1111455);
nand I_65236 (I1110974,I1111489,I1111373);
not I_65237 (I1111578,I2514);
DFFARX1 I_65238 (I1236279,I2507,I1111578,I1111604,);
and I_65239 (I1111612,I1111604,I1236273);
DFFARX1 I_65240 (I1111612,I2507,I1111578,I1111561,);
DFFARX1 I_65241 (I1236258,I2507,I1111578,I1111652,);
not I_65242 (I1111660,I1236264);
not I_65243 (I1111677,I1236276);
nand I_65244 (I1111694,I1111677,I1111660);
nor I_65245 (I1111549,I1111652,I1111694);
DFFARX1 I_65246 (I1111694,I2507,I1111578,I1111734,);
not I_65247 (I1111570,I1111734);
not I_65248 (I1111756,I1236258);
nand I_65249 (I1111773,I1111677,I1111756);
DFFARX1 I_65250 (I1111773,I2507,I1111578,I1111799,);
not I_65251 (I1111807,I1111799);
not I_65252 (I1111824,I1236282);
nand I_65253 (I1111841,I1111824,I1236270);
and I_65254 (I1111858,I1111660,I1111841);
nor I_65255 (I1111875,I1111773,I1111858);
DFFARX1 I_65256 (I1111875,I2507,I1111578,I1111546,);
DFFARX1 I_65257 (I1111858,I2507,I1111578,I1111567,);
nor I_65258 (I1111920,I1236282,I1236261);
nor I_65259 (I1111558,I1111773,I1111920);
or I_65260 (I1111951,I1236282,I1236261);
nor I_65261 (I1111968,I1236267,I1236261);
DFFARX1 I_65262 (I1111968,I2507,I1111578,I1111994,);
not I_65263 (I1112002,I1111994);
nor I_65264 (I1111564,I1112002,I1111807);
nand I_65265 (I1112033,I1112002,I1111652);
not I_65266 (I1112050,I1236267);
nand I_65267 (I1112067,I1112050,I1111756);
nand I_65268 (I1112084,I1112002,I1112067);
nand I_65269 (I1111555,I1112084,I1112033);
nand I_65270 (I1111552,I1112067,I1111951);
not I_65271 (I1112156,I2514);
DFFARX1 I_65272 (I84923,I2507,I1112156,I1112182,);
and I_65273 (I1112190,I1112182,I84899);
DFFARX1 I_65274 (I1112190,I2507,I1112156,I1112139,);
DFFARX1 I_65275 (I84917,I2507,I1112156,I1112230,);
not I_65276 (I1112238,I84905);
not I_65277 (I1112255,I84902);
nand I_65278 (I1112272,I1112255,I1112238);
nor I_65279 (I1112127,I1112230,I1112272);
DFFARX1 I_65280 (I1112272,I2507,I1112156,I1112312,);
not I_65281 (I1112148,I1112312);
not I_65282 (I1112334,I84911);
nand I_65283 (I1112351,I1112255,I1112334);
DFFARX1 I_65284 (I1112351,I2507,I1112156,I1112377,);
not I_65285 (I1112385,I1112377);
not I_65286 (I1112402,I84902);
nand I_65287 (I1112419,I1112402,I84920);
and I_65288 (I1112436,I1112238,I1112419);
nor I_65289 (I1112453,I1112351,I1112436);
DFFARX1 I_65290 (I1112453,I2507,I1112156,I1112124,);
DFFARX1 I_65291 (I1112436,I2507,I1112156,I1112145,);
nor I_65292 (I1112498,I84902,I84914);
nor I_65293 (I1112136,I1112351,I1112498);
or I_65294 (I1112529,I84902,I84914);
nor I_65295 (I1112546,I84908,I84899);
DFFARX1 I_65296 (I1112546,I2507,I1112156,I1112572,);
not I_65297 (I1112580,I1112572);
nor I_65298 (I1112142,I1112580,I1112385);
nand I_65299 (I1112611,I1112580,I1112230);
not I_65300 (I1112628,I84908);
nand I_65301 (I1112645,I1112628,I1112334);
nand I_65302 (I1112662,I1112580,I1112645);
nand I_65303 (I1112133,I1112662,I1112611);
nand I_65304 (I1112130,I1112645,I1112529);
not I_65305 (I1112734,I2514);
DFFARX1 I_65306 (I883409,I2507,I1112734,I1112760,);
and I_65307 (I1112768,I1112760,I883415);
DFFARX1 I_65308 (I1112768,I2507,I1112734,I1112717,);
DFFARX1 I_65309 (I883421,I2507,I1112734,I1112808,);
not I_65310 (I1112816,I883406);
not I_65311 (I1112833,I883406);
nand I_65312 (I1112850,I1112833,I1112816);
nor I_65313 (I1112705,I1112808,I1112850);
DFFARX1 I_65314 (I1112850,I2507,I1112734,I1112890,);
not I_65315 (I1112726,I1112890);
not I_65316 (I1112912,I883424);
nand I_65317 (I1112929,I1112833,I1112912);
DFFARX1 I_65318 (I1112929,I2507,I1112734,I1112955,);
not I_65319 (I1112963,I1112955);
not I_65320 (I1112980,I883418);
nand I_65321 (I1112997,I1112980,I883409);
and I_65322 (I1113014,I1112816,I1112997);
nor I_65323 (I1113031,I1112929,I1113014);
DFFARX1 I_65324 (I1113031,I2507,I1112734,I1112702,);
DFFARX1 I_65325 (I1113014,I2507,I1112734,I1112723,);
nor I_65326 (I1113076,I883418,I883427);
nor I_65327 (I1112714,I1112929,I1113076);
or I_65328 (I1113107,I883418,I883427);
nor I_65329 (I1113124,I883412,I883412);
DFFARX1 I_65330 (I1113124,I2507,I1112734,I1113150,);
not I_65331 (I1113158,I1113150);
nor I_65332 (I1112720,I1113158,I1112963);
nand I_65333 (I1113189,I1113158,I1112808);
not I_65334 (I1113206,I883412);
nand I_65335 (I1113223,I1113206,I1112912);
nand I_65336 (I1113240,I1113158,I1113223);
nand I_65337 (I1112711,I1113240,I1113189);
nand I_65338 (I1112708,I1113223,I1113107);
not I_65339 (I1113312,I2514);
DFFARX1 I_65340 (I126556,I2507,I1113312,I1113338,);
and I_65341 (I1113346,I1113338,I126532);
DFFARX1 I_65342 (I1113346,I2507,I1113312,I1113295,);
DFFARX1 I_65343 (I126550,I2507,I1113312,I1113386,);
not I_65344 (I1113394,I126538);
not I_65345 (I1113411,I126535);
nand I_65346 (I1113428,I1113411,I1113394);
nor I_65347 (I1113283,I1113386,I1113428);
DFFARX1 I_65348 (I1113428,I2507,I1113312,I1113468,);
not I_65349 (I1113304,I1113468);
not I_65350 (I1113490,I126544);
nand I_65351 (I1113507,I1113411,I1113490);
DFFARX1 I_65352 (I1113507,I2507,I1113312,I1113533,);
not I_65353 (I1113541,I1113533);
not I_65354 (I1113558,I126535);
nand I_65355 (I1113575,I1113558,I126553);
and I_65356 (I1113592,I1113394,I1113575);
nor I_65357 (I1113609,I1113507,I1113592);
DFFARX1 I_65358 (I1113609,I2507,I1113312,I1113280,);
DFFARX1 I_65359 (I1113592,I2507,I1113312,I1113301,);
nor I_65360 (I1113654,I126535,I126547);
nor I_65361 (I1113292,I1113507,I1113654);
or I_65362 (I1113685,I126535,I126547);
nor I_65363 (I1113702,I126541,I126532);
DFFARX1 I_65364 (I1113702,I2507,I1113312,I1113728,);
not I_65365 (I1113736,I1113728);
nor I_65366 (I1113298,I1113736,I1113541);
nand I_65367 (I1113767,I1113736,I1113386);
not I_65368 (I1113784,I126541);
nand I_65369 (I1113801,I1113784,I1113490);
nand I_65370 (I1113818,I1113736,I1113801);
nand I_65371 (I1113289,I1113818,I1113767);
nand I_65372 (I1113286,I1113801,I1113685);
not I_65373 (I1113890,I2514);
DFFARX1 I_65374 (I1254778,I2507,I1113890,I1113916,);
and I_65375 (I1113924,I1113916,I1254760);
DFFARX1 I_65376 (I1113924,I2507,I1113890,I1113873,);
DFFARX1 I_65377 (I1254769,I2507,I1113890,I1113964,);
not I_65378 (I1113972,I1254754);
not I_65379 (I1113989,I1254766);
nand I_65380 (I1114006,I1113989,I1113972);
nor I_65381 (I1113861,I1113964,I1114006);
DFFARX1 I_65382 (I1114006,I2507,I1113890,I1114046,);
not I_65383 (I1113882,I1114046);
not I_65384 (I1114068,I1254757);
nand I_65385 (I1114085,I1113989,I1114068);
DFFARX1 I_65386 (I1114085,I2507,I1113890,I1114111,);
not I_65387 (I1114119,I1114111);
not I_65388 (I1114136,I1254754);
nand I_65389 (I1114153,I1114136,I1254757);
and I_65390 (I1114170,I1113972,I1114153);
nor I_65391 (I1114187,I1114085,I1114170);
DFFARX1 I_65392 (I1114187,I2507,I1113890,I1113858,);
DFFARX1 I_65393 (I1114170,I2507,I1113890,I1113879,);
nor I_65394 (I1114232,I1254754,I1254775);
nor I_65395 (I1113870,I1114085,I1114232);
or I_65396 (I1114263,I1254754,I1254775);
nor I_65397 (I1114280,I1254763,I1254772);
DFFARX1 I_65398 (I1114280,I2507,I1113890,I1114306,);
not I_65399 (I1114314,I1114306);
nor I_65400 (I1113876,I1114314,I1114119);
nand I_65401 (I1114345,I1114314,I1113964);
not I_65402 (I1114362,I1254763);
nand I_65403 (I1114379,I1114362,I1114068);
nand I_65404 (I1114396,I1114314,I1114379);
nand I_65405 (I1113867,I1114396,I1114345);
nand I_65406 (I1113864,I1114379,I1114263);
not I_65407 (I1114468,I2514);
DFFARX1 I_65408 (I555015,I2507,I1114468,I1114494,);
and I_65409 (I1114502,I1114494,I555003);
DFFARX1 I_65410 (I1114502,I2507,I1114468,I1114451,);
DFFARX1 I_65411 (I555018,I2507,I1114468,I1114542,);
not I_65412 (I1114550,I555009);
not I_65413 (I1114567,I555000);
nand I_65414 (I1114584,I1114567,I1114550);
nor I_65415 (I1114439,I1114542,I1114584);
DFFARX1 I_65416 (I1114584,I2507,I1114468,I1114624,);
not I_65417 (I1114460,I1114624);
not I_65418 (I1114646,I555006);
nand I_65419 (I1114663,I1114567,I1114646);
DFFARX1 I_65420 (I1114663,I2507,I1114468,I1114689,);
not I_65421 (I1114697,I1114689);
not I_65422 (I1114714,I555021);
nand I_65423 (I1114731,I1114714,I555024);
and I_65424 (I1114748,I1114550,I1114731);
nor I_65425 (I1114765,I1114663,I1114748);
DFFARX1 I_65426 (I1114765,I2507,I1114468,I1114436,);
DFFARX1 I_65427 (I1114748,I2507,I1114468,I1114457,);
nor I_65428 (I1114810,I555021,I555000);
nor I_65429 (I1114448,I1114663,I1114810);
or I_65430 (I1114841,I555021,I555000);
nor I_65431 (I1114858,I555012,I555003);
DFFARX1 I_65432 (I1114858,I2507,I1114468,I1114884,);
not I_65433 (I1114892,I1114884);
nor I_65434 (I1114454,I1114892,I1114697);
nand I_65435 (I1114923,I1114892,I1114542);
not I_65436 (I1114940,I555012);
nand I_65437 (I1114957,I1114940,I1114646);
nand I_65438 (I1114974,I1114892,I1114957);
nand I_65439 (I1114445,I1114974,I1114923);
nand I_65440 (I1114442,I1114957,I1114841);
not I_65441 (I1115046,I2514);
DFFARX1 I_65442 (I284472,I2507,I1115046,I1115072,);
and I_65443 (I1115080,I1115072,I284457);
DFFARX1 I_65444 (I1115080,I2507,I1115046,I1115029,);
DFFARX1 I_65445 (I284463,I2507,I1115046,I1115120,);
not I_65446 (I1115128,I284445);
not I_65447 (I1115145,I284466);
nand I_65448 (I1115162,I1115145,I1115128);
nor I_65449 (I1115017,I1115120,I1115162);
DFFARX1 I_65450 (I1115162,I2507,I1115046,I1115202,);
not I_65451 (I1115038,I1115202);
not I_65452 (I1115224,I284469);
nand I_65453 (I1115241,I1115145,I1115224);
DFFARX1 I_65454 (I1115241,I2507,I1115046,I1115267,);
not I_65455 (I1115275,I1115267);
not I_65456 (I1115292,I284460);
nand I_65457 (I1115309,I1115292,I284448);
and I_65458 (I1115326,I1115128,I1115309);
nor I_65459 (I1115343,I1115241,I1115326);
DFFARX1 I_65460 (I1115343,I2507,I1115046,I1115014,);
DFFARX1 I_65461 (I1115326,I2507,I1115046,I1115035,);
nor I_65462 (I1115388,I284460,I284454);
nor I_65463 (I1115026,I1115241,I1115388);
or I_65464 (I1115419,I284460,I284454);
nor I_65465 (I1115436,I284451,I284445);
DFFARX1 I_65466 (I1115436,I2507,I1115046,I1115462,);
not I_65467 (I1115470,I1115462);
nor I_65468 (I1115032,I1115470,I1115275);
nand I_65469 (I1115501,I1115470,I1115120);
not I_65470 (I1115518,I284451);
nand I_65471 (I1115535,I1115518,I1115224);
nand I_65472 (I1115552,I1115470,I1115535);
nand I_65473 (I1115023,I1115552,I1115501);
nand I_65474 (I1115020,I1115535,I1115419);
not I_65475 (I1115624,I2514);
DFFARX1 I_65476 (I727837,I2507,I1115624,I1115650,);
and I_65477 (I1115658,I1115650,I727825);
DFFARX1 I_65478 (I1115658,I2507,I1115624,I1115607,);
DFFARX1 I_65479 (I727828,I2507,I1115624,I1115698,);
not I_65480 (I1115706,I727822);
not I_65481 (I1115723,I727846);
nand I_65482 (I1115740,I1115723,I1115706);
nor I_65483 (I1115595,I1115698,I1115740);
DFFARX1 I_65484 (I1115740,I2507,I1115624,I1115780,);
not I_65485 (I1115616,I1115780);
not I_65486 (I1115802,I727834);
nand I_65487 (I1115819,I1115723,I1115802);
DFFARX1 I_65488 (I1115819,I2507,I1115624,I1115845,);
not I_65489 (I1115853,I1115845);
not I_65490 (I1115870,I727843);
nand I_65491 (I1115887,I1115870,I727840);
and I_65492 (I1115904,I1115706,I1115887);
nor I_65493 (I1115921,I1115819,I1115904);
DFFARX1 I_65494 (I1115921,I2507,I1115624,I1115592,);
DFFARX1 I_65495 (I1115904,I2507,I1115624,I1115613,);
nor I_65496 (I1115966,I727843,I727831);
nor I_65497 (I1115604,I1115819,I1115966);
or I_65498 (I1115997,I727843,I727831);
nor I_65499 (I1116014,I727822,I727825);
DFFARX1 I_65500 (I1116014,I2507,I1115624,I1116040,);
not I_65501 (I1116048,I1116040);
nor I_65502 (I1115610,I1116048,I1115853);
nand I_65503 (I1116079,I1116048,I1115698);
not I_65504 (I1116096,I727822);
nand I_65505 (I1116113,I1116096,I1115802);
nand I_65506 (I1116130,I1116048,I1116113);
nand I_65507 (I1115601,I1116130,I1116079);
nand I_65508 (I1115598,I1116113,I1115997);
not I_65509 (I1116202,I2514);
DFFARX1 I_65510 (I528007,I2507,I1116202,I1116228,);
and I_65511 (I1116236,I1116228,I528022);
DFFARX1 I_65512 (I1116236,I2507,I1116202,I1116185,);
DFFARX1 I_65513 (I528013,I2507,I1116202,I1116276,);
not I_65514 (I1116284,I528007);
not I_65515 (I1116301,I528025);
nand I_65516 (I1116318,I1116301,I1116284);
nor I_65517 (I1116173,I1116276,I1116318);
DFFARX1 I_65518 (I1116318,I2507,I1116202,I1116358,);
not I_65519 (I1116194,I1116358);
not I_65520 (I1116380,I528016);
nand I_65521 (I1116397,I1116301,I1116380);
DFFARX1 I_65522 (I1116397,I2507,I1116202,I1116423,);
not I_65523 (I1116431,I1116423);
not I_65524 (I1116448,I528028);
nand I_65525 (I1116465,I1116448,I528004);
and I_65526 (I1116482,I1116284,I1116465);
nor I_65527 (I1116499,I1116397,I1116482);
DFFARX1 I_65528 (I1116499,I2507,I1116202,I1116170,);
DFFARX1 I_65529 (I1116482,I2507,I1116202,I1116191,);
nor I_65530 (I1116544,I528028,I528004);
nor I_65531 (I1116182,I1116397,I1116544);
or I_65532 (I1116575,I528028,I528004);
nor I_65533 (I1116592,I528010,I528019);
DFFARX1 I_65534 (I1116592,I2507,I1116202,I1116618,);
not I_65535 (I1116626,I1116618);
nor I_65536 (I1116188,I1116626,I1116431);
nand I_65537 (I1116657,I1116626,I1116276);
not I_65538 (I1116674,I528010);
nand I_65539 (I1116691,I1116674,I1116380);
nand I_65540 (I1116708,I1116626,I1116691);
nand I_65541 (I1116179,I1116708,I1116657);
nand I_65542 (I1116176,I1116691,I1116575);
not I_65543 (I1116780,I2514);
DFFARX1 I_65544 (I1034267,I2507,I1116780,I1116806,);
and I_65545 (I1116814,I1116806,I1034264);
DFFARX1 I_65546 (I1116814,I2507,I1116780,I1116763,);
DFFARX1 I_65547 (I1034270,I2507,I1116780,I1116854,);
not I_65548 (I1116862,I1034273);
not I_65549 (I1116879,I1034267);
nand I_65550 (I1116896,I1116879,I1116862);
nor I_65551 (I1116751,I1116854,I1116896);
DFFARX1 I_65552 (I1116896,I2507,I1116780,I1116936,);
not I_65553 (I1116772,I1116936);
not I_65554 (I1116958,I1034282);
nand I_65555 (I1116975,I1116879,I1116958);
DFFARX1 I_65556 (I1116975,I2507,I1116780,I1117001,);
not I_65557 (I1117009,I1117001);
not I_65558 (I1117026,I1034279);
nand I_65559 (I1117043,I1117026,I1034285);
and I_65560 (I1117060,I1116862,I1117043);
nor I_65561 (I1117077,I1116975,I1117060);
DFFARX1 I_65562 (I1117077,I2507,I1116780,I1116748,);
DFFARX1 I_65563 (I1117060,I2507,I1116780,I1116769,);
nor I_65564 (I1117122,I1034279,I1034264);
nor I_65565 (I1116760,I1116975,I1117122);
or I_65566 (I1117153,I1034279,I1034264);
nor I_65567 (I1117170,I1034276,I1034270);
DFFARX1 I_65568 (I1117170,I2507,I1116780,I1117196,);
not I_65569 (I1117204,I1117196);
nor I_65570 (I1116766,I1117204,I1117009);
nand I_65571 (I1117235,I1117204,I1116854);
not I_65572 (I1117252,I1034276);
nand I_65573 (I1117269,I1117252,I1116958);
nand I_65574 (I1117286,I1117204,I1117269);
nand I_65575 (I1116757,I1117286,I1117235);
nand I_65576 (I1116754,I1117269,I1117153);
not I_65577 (I1117358,I2514);
DFFARX1 I_65578 (I64897,I2507,I1117358,I1117384,);
and I_65579 (I1117392,I1117384,I64873);
DFFARX1 I_65580 (I1117392,I2507,I1117358,I1117341,);
DFFARX1 I_65581 (I64891,I2507,I1117358,I1117432,);
not I_65582 (I1117440,I64879);
not I_65583 (I1117457,I64876);
nand I_65584 (I1117474,I1117457,I1117440);
nor I_65585 (I1117329,I1117432,I1117474);
DFFARX1 I_65586 (I1117474,I2507,I1117358,I1117514,);
not I_65587 (I1117350,I1117514);
not I_65588 (I1117536,I64885);
nand I_65589 (I1117553,I1117457,I1117536);
DFFARX1 I_65590 (I1117553,I2507,I1117358,I1117579,);
not I_65591 (I1117587,I1117579);
not I_65592 (I1117604,I64876);
nand I_65593 (I1117621,I1117604,I64894);
and I_65594 (I1117638,I1117440,I1117621);
nor I_65595 (I1117655,I1117553,I1117638);
DFFARX1 I_65596 (I1117655,I2507,I1117358,I1117326,);
DFFARX1 I_65597 (I1117638,I2507,I1117358,I1117347,);
nor I_65598 (I1117700,I64876,I64888);
nor I_65599 (I1117338,I1117553,I1117700);
or I_65600 (I1117731,I64876,I64888);
nor I_65601 (I1117748,I64882,I64873);
DFFARX1 I_65602 (I1117748,I2507,I1117358,I1117774,);
not I_65603 (I1117782,I1117774);
nor I_65604 (I1117344,I1117782,I1117587);
nand I_65605 (I1117813,I1117782,I1117432);
not I_65606 (I1117830,I64882);
nand I_65607 (I1117847,I1117830,I1117536);
nand I_65608 (I1117864,I1117782,I1117847);
nand I_65609 (I1117335,I1117864,I1117813);
nand I_65610 (I1117332,I1117847,I1117731);
not I_65611 (I1117936,I2514);
DFFARX1 I_65612 (I857059,I2507,I1117936,I1117962,);
and I_65613 (I1117970,I1117962,I857065);
DFFARX1 I_65614 (I1117970,I2507,I1117936,I1117919,);
DFFARX1 I_65615 (I857071,I2507,I1117936,I1118010,);
not I_65616 (I1118018,I857056);
not I_65617 (I1118035,I857056);
nand I_65618 (I1118052,I1118035,I1118018);
nor I_65619 (I1117907,I1118010,I1118052);
DFFARX1 I_65620 (I1118052,I2507,I1117936,I1118092,);
not I_65621 (I1117928,I1118092);
not I_65622 (I1118114,I857074);
nand I_65623 (I1118131,I1118035,I1118114);
DFFARX1 I_65624 (I1118131,I2507,I1117936,I1118157,);
not I_65625 (I1118165,I1118157);
not I_65626 (I1118182,I857068);
nand I_65627 (I1118199,I1118182,I857059);
and I_65628 (I1118216,I1118018,I1118199);
nor I_65629 (I1118233,I1118131,I1118216);
DFFARX1 I_65630 (I1118233,I2507,I1117936,I1117904,);
DFFARX1 I_65631 (I1118216,I2507,I1117936,I1117925,);
nor I_65632 (I1118278,I857068,I857077);
nor I_65633 (I1117916,I1118131,I1118278);
or I_65634 (I1118309,I857068,I857077);
nor I_65635 (I1118326,I857062,I857062);
DFFARX1 I_65636 (I1118326,I2507,I1117936,I1118352,);
not I_65637 (I1118360,I1118352);
nor I_65638 (I1117922,I1118360,I1118165);
nand I_65639 (I1118391,I1118360,I1118010);
not I_65640 (I1118408,I857062);
nand I_65641 (I1118425,I1118408,I1118114);
nand I_65642 (I1118442,I1118360,I1118425);
nand I_65643 (I1117913,I1118442,I1118391);
nand I_65644 (I1117910,I1118425,I1118309);
not I_65645 (I1118514,I2514);
DFFARX1 I_65646 (I992875,I2507,I1118514,I1118540,);
and I_65647 (I1118548,I1118540,I992869);
DFFARX1 I_65648 (I1118548,I2507,I1118514,I1118497,);
DFFARX1 I_65649 (I992887,I2507,I1118514,I1118588,);
not I_65650 (I1118596,I992878);
not I_65651 (I1118613,I992890);
nand I_65652 (I1118630,I1118613,I1118596);
nor I_65653 (I1118485,I1118588,I1118630);
DFFARX1 I_65654 (I1118630,I2507,I1118514,I1118670,);
not I_65655 (I1118506,I1118670);
not I_65656 (I1118692,I992896);
nand I_65657 (I1118709,I1118613,I1118692);
DFFARX1 I_65658 (I1118709,I2507,I1118514,I1118735,);
not I_65659 (I1118743,I1118735);
not I_65660 (I1118760,I992872);
nand I_65661 (I1118777,I1118760,I992893);
and I_65662 (I1118794,I1118596,I1118777);
nor I_65663 (I1118811,I1118709,I1118794);
DFFARX1 I_65664 (I1118811,I2507,I1118514,I1118482,);
DFFARX1 I_65665 (I1118794,I2507,I1118514,I1118503,);
nor I_65666 (I1118856,I992872,I992884);
nor I_65667 (I1118494,I1118709,I1118856);
or I_65668 (I1118887,I992872,I992884);
nor I_65669 (I1118904,I992869,I992881);
DFFARX1 I_65670 (I1118904,I2507,I1118514,I1118930,);
not I_65671 (I1118938,I1118930);
nor I_65672 (I1118500,I1118938,I1118743);
nand I_65673 (I1118969,I1118938,I1118588);
not I_65674 (I1118986,I992869);
nand I_65675 (I1119003,I1118986,I1118692);
nand I_65676 (I1119020,I1118938,I1119003);
nand I_65677 (I1118491,I1119020,I1118969);
nand I_65678 (I1118488,I1119003,I1118887);
not I_65679 (I1119092,I2514);
DFFARX1 I_65680 (I574089,I2507,I1119092,I1119118,);
and I_65681 (I1119126,I1119118,I574077);
DFFARX1 I_65682 (I1119126,I2507,I1119092,I1119075,);
DFFARX1 I_65683 (I574092,I2507,I1119092,I1119166,);
not I_65684 (I1119174,I574083);
not I_65685 (I1119191,I574074);
nand I_65686 (I1119208,I1119191,I1119174);
nor I_65687 (I1119063,I1119166,I1119208);
DFFARX1 I_65688 (I1119208,I2507,I1119092,I1119248,);
not I_65689 (I1119084,I1119248);
not I_65690 (I1119270,I574080);
nand I_65691 (I1119287,I1119191,I1119270);
DFFARX1 I_65692 (I1119287,I2507,I1119092,I1119313,);
not I_65693 (I1119321,I1119313);
not I_65694 (I1119338,I574095);
nand I_65695 (I1119355,I1119338,I574098);
and I_65696 (I1119372,I1119174,I1119355);
nor I_65697 (I1119389,I1119287,I1119372);
DFFARX1 I_65698 (I1119389,I2507,I1119092,I1119060,);
DFFARX1 I_65699 (I1119372,I2507,I1119092,I1119081,);
nor I_65700 (I1119434,I574095,I574074);
nor I_65701 (I1119072,I1119287,I1119434);
or I_65702 (I1119465,I574095,I574074);
nor I_65703 (I1119482,I574086,I574077);
DFFARX1 I_65704 (I1119482,I2507,I1119092,I1119508,);
not I_65705 (I1119516,I1119508);
nor I_65706 (I1119078,I1119516,I1119321);
nand I_65707 (I1119547,I1119516,I1119166);
not I_65708 (I1119564,I574086);
nand I_65709 (I1119581,I1119564,I1119270);
nand I_65710 (I1119598,I1119516,I1119581);
nand I_65711 (I1119069,I1119598,I1119547);
nand I_65712 (I1119066,I1119581,I1119465);
not I_65713 (I1119670,I2514);
DFFARX1 I_65714 (I830182,I2507,I1119670,I1119696,);
and I_65715 (I1119704,I1119696,I830188);
DFFARX1 I_65716 (I1119704,I2507,I1119670,I1119653,);
DFFARX1 I_65717 (I830194,I2507,I1119670,I1119744,);
not I_65718 (I1119752,I830179);
not I_65719 (I1119769,I830179);
nand I_65720 (I1119786,I1119769,I1119752);
nor I_65721 (I1119641,I1119744,I1119786);
DFFARX1 I_65722 (I1119786,I2507,I1119670,I1119826,);
not I_65723 (I1119662,I1119826);
not I_65724 (I1119848,I830197);
nand I_65725 (I1119865,I1119769,I1119848);
DFFARX1 I_65726 (I1119865,I2507,I1119670,I1119891,);
not I_65727 (I1119899,I1119891);
not I_65728 (I1119916,I830191);
nand I_65729 (I1119933,I1119916,I830182);
and I_65730 (I1119950,I1119752,I1119933);
nor I_65731 (I1119967,I1119865,I1119950);
DFFARX1 I_65732 (I1119967,I2507,I1119670,I1119638,);
DFFARX1 I_65733 (I1119950,I2507,I1119670,I1119659,);
nor I_65734 (I1120012,I830191,I830200);
nor I_65735 (I1119650,I1119865,I1120012);
or I_65736 (I1120043,I830191,I830200);
nor I_65737 (I1120060,I830185,I830185);
DFFARX1 I_65738 (I1120060,I2507,I1119670,I1120086,);
not I_65739 (I1120094,I1120086);
nor I_65740 (I1119656,I1120094,I1119899);
nand I_65741 (I1120125,I1120094,I1119744);
not I_65742 (I1120142,I830185);
nand I_65743 (I1120159,I1120142,I1119848);
nand I_65744 (I1120176,I1120094,I1120159);
nand I_65745 (I1119647,I1120176,I1120125);
nand I_65746 (I1119644,I1120159,I1120043);
not I_65747 (I1120248,I2514);
DFFARX1 I_65748 (I238885,I2507,I1120248,I1120274,);
and I_65749 (I1120282,I1120274,I238888);
DFFARX1 I_65750 (I1120282,I2507,I1120248,I1120231,);
DFFARX1 I_65751 (I238888,I2507,I1120248,I1120322,);
not I_65752 (I1120330,I238903);
not I_65753 (I1120347,I238909);
nand I_65754 (I1120364,I1120347,I1120330);
nor I_65755 (I1120219,I1120322,I1120364);
DFFARX1 I_65756 (I1120364,I2507,I1120248,I1120404,);
not I_65757 (I1120240,I1120404);
not I_65758 (I1120426,I238897);
nand I_65759 (I1120443,I1120347,I1120426);
DFFARX1 I_65760 (I1120443,I2507,I1120248,I1120469,);
not I_65761 (I1120477,I1120469);
not I_65762 (I1120494,I238894);
nand I_65763 (I1120511,I1120494,I238891);
and I_65764 (I1120528,I1120330,I1120511);
nor I_65765 (I1120545,I1120443,I1120528);
DFFARX1 I_65766 (I1120545,I2507,I1120248,I1120216,);
DFFARX1 I_65767 (I1120528,I2507,I1120248,I1120237,);
nor I_65768 (I1120590,I238894,I238885);
nor I_65769 (I1120228,I1120443,I1120590);
or I_65770 (I1120621,I238894,I238885);
nor I_65771 (I1120638,I238900,I238906);
DFFARX1 I_65772 (I1120638,I2507,I1120248,I1120664,);
not I_65773 (I1120672,I1120664);
nor I_65774 (I1120234,I1120672,I1120477);
nand I_65775 (I1120703,I1120672,I1120322);
not I_65776 (I1120720,I238900);
nand I_65777 (I1120737,I1120720,I1120426);
nand I_65778 (I1120754,I1120672,I1120737);
nand I_65779 (I1120225,I1120754,I1120703);
nand I_65780 (I1120222,I1120737,I1120621);
not I_65781 (I1120826,I2514);
DFFARX1 I_65782 (I1355914,I2507,I1120826,I1120852,);
and I_65783 (I1120860,I1120852,I1355896);
DFFARX1 I_65784 (I1120860,I2507,I1120826,I1120809,);
DFFARX1 I_65785 (I1355887,I2507,I1120826,I1120900,);
not I_65786 (I1120908,I1355902);
not I_65787 (I1120925,I1355890);
nand I_65788 (I1120942,I1120925,I1120908);
nor I_65789 (I1120797,I1120900,I1120942);
DFFARX1 I_65790 (I1120942,I2507,I1120826,I1120982,);
not I_65791 (I1120818,I1120982);
not I_65792 (I1121004,I1355899);
nand I_65793 (I1121021,I1120925,I1121004);
DFFARX1 I_65794 (I1121021,I2507,I1120826,I1121047,);
not I_65795 (I1121055,I1121047);
not I_65796 (I1121072,I1355908);
nand I_65797 (I1121089,I1121072,I1355887);
and I_65798 (I1121106,I1120908,I1121089);
nor I_65799 (I1121123,I1121021,I1121106);
DFFARX1 I_65800 (I1121123,I2507,I1120826,I1120794,);
DFFARX1 I_65801 (I1121106,I2507,I1120826,I1120815,);
nor I_65802 (I1121168,I1355908,I1355911);
nor I_65803 (I1120806,I1121021,I1121168);
or I_65804 (I1121199,I1355908,I1355911);
nor I_65805 (I1121216,I1355905,I1355893);
DFFARX1 I_65806 (I1121216,I2507,I1120826,I1121242,);
not I_65807 (I1121250,I1121242);
nor I_65808 (I1120812,I1121250,I1121055);
nand I_65809 (I1121281,I1121250,I1120900);
not I_65810 (I1121298,I1355905);
nand I_65811 (I1121315,I1121298,I1121004);
nand I_65812 (I1121332,I1121250,I1121315);
nand I_65813 (I1120803,I1121332,I1121281);
nand I_65814 (I1120800,I1121315,I1121199);
not I_65815 (I1121404,I2514);
DFFARX1 I_65816 (I110746,I2507,I1121404,I1121430,);
and I_65817 (I1121438,I1121430,I110722);
DFFARX1 I_65818 (I1121438,I2507,I1121404,I1121387,);
DFFARX1 I_65819 (I110740,I2507,I1121404,I1121478,);
not I_65820 (I1121486,I110728);
not I_65821 (I1121503,I110725);
nand I_65822 (I1121520,I1121503,I1121486);
nor I_65823 (I1121375,I1121478,I1121520);
DFFARX1 I_65824 (I1121520,I2507,I1121404,I1121560,);
not I_65825 (I1121396,I1121560);
not I_65826 (I1121582,I110734);
nand I_65827 (I1121599,I1121503,I1121582);
DFFARX1 I_65828 (I1121599,I2507,I1121404,I1121625,);
not I_65829 (I1121633,I1121625);
not I_65830 (I1121650,I110725);
nand I_65831 (I1121667,I1121650,I110743);
and I_65832 (I1121684,I1121486,I1121667);
nor I_65833 (I1121701,I1121599,I1121684);
DFFARX1 I_65834 (I1121701,I2507,I1121404,I1121372,);
DFFARX1 I_65835 (I1121684,I2507,I1121404,I1121393,);
nor I_65836 (I1121746,I110725,I110737);
nor I_65837 (I1121384,I1121599,I1121746);
or I_65838 (I1121777,I110725,I110737);
nor I_65839 (I1121794,I110731,I110722);
DFFARX1 I_65840 (I1121794,I2507,I1121404,I1121820,);
not I_65841 (I1121828,I1121820);
nor I_65842 (I1121390,I1121828,I1121633);
nand I_65843 (I1121859,I1121828,I1121478);
not I_65844 (I1121876,I110731);
nand I_65845 (I1121893,I1121876,I1121582);
nand I_65846 (I1121910,I1121828,I1121893);
nand I_65847 (I1121381,I1121910,I1121859);
nand I_65848 (I1121378,I1121893,I1121777);
not I_65849 (I1121982,I2514);
DFFARX1 I_65850 (I998689,I2507,I1121982,I1122008,);
and I_65851 (I1122016,I1122008,I998683);
DFFARX1 I_65852 (I1122016,I2507,I1121982,I1121965,);
DFFARX1 I_65853 (I998701,I2507,I1121982,I1122056,);
not I_65854 (I1122064,I998692);
not I_65855 (I1122081,I998704);
nand I_65856 (I1122098,I1122081,I1122064);
nor I_65857 (I1121953,I1122056,I1122098);
DFFARX1 I_65858 (I1122098,I2507,I1121982,I1122138,);
not I_65859 (I1121974,I1122138);
not I_65860 (I1122160,I998710);
nand I_65861 (I1122177,I1122081,I1122160);
DFFARX1 I_65862 (I1122177,I2507,I1121982,I1122203,);
not I_65863 (I1122211,I1122203);
not I_65864 (I1122228,I998686);
nand I_65865 (I1122245,I1122228,I998707);
and I_65866 (I1122262,I1122064,I1122245);
nor I_65867 (I1122279,I1122177,I1122262);
DFFARX1 I_65868 (I1122279,I2507,I1121982,I1121950,);
DFFARX1 I_65869 (I1122262,I2507,I1121982,I1121971,);
nor I_65870 (I1122324,I998686,I998698);
nor I_65871 (I1121962,I1122177,I1122324);
or I_65872 (I1122355,I998686,I998698);
nor I_65873 (I1122372,I998683,I998695);
DFFARX1 I_65874 (I1122372,I2507,I1121982,I1122398,);
not I_65875 (I1122406,I1122398);
nor I_65876 (I1121968,I1122406,I1122211);
nand I_65877 (I1122437,I1122406,I1122056);
not I_65878 (I1122454,I998683);
nand I_65879 (I1122471,I1122454,I1122160);
nand I_65880 (I1122488,I1122406,I1122471);
nand I_65881 (I1121959,I1122488,I1122437);
nand I_65882 (I1121956,I1122471,I1122355);
not I_65883 (I1122560,I2514);
DFFARX1 I_65884 (I1394589,I2507,I1122560,I1122586,);
and I_65885 (I1122594,I1122586,I1394571);
DFFARX1 I_65886 (I1122594,I2507,I1122560,I1122543,);
DFFARX1 I_65887 (I1394562,I2507,I1122560,I1122634,);
not I_65888 (I1122642,I1394577);
not I_65889 (I1122659,I1394565);
nand I_65890 (I1122676,I1122659,I1122642);
nor I_65891 (I1122531,I1122634,I1122676);
DFFARX1 I_65892 (I1122676,I2507,I1122560,I1122716,);
not I_65893 (I1122552,I1122716);
not I_65894 (I1122738,I1394574);
nand I_65895 (I1122755,I1122659,I1122738);
DFFARX1 I_65896 (I1122755,I2507,I1122560,I1122781,);
not I_65897 (I1122789,I1122781);
not I_65898 (I1122806,I1394583);
nand I_65899 (I1122823,I1122806,I1394562);
and I_65900 (I1122840,I1122642,I1122823);
nor I_65901 (I1122857,I1122755,I1122840);
DFFARX1 I_65902 (I1122857,I2507,I1122560,I1122528,);
DFFARX1 I_65903 (I1122840,I2507,I1122560,I1122549,);
nor I_65904 (I1122902,I1394583,I1394586);
nor I_65905 (I1122540,I1122755,I1122902);
or I_65906 (I1122933,I1394583,I1394586);
nor I_65907 (I1122950,I1394580,I1394568);
DFFARX1 I_65908 (I1122950,I2507,I1122560,I1122976,);
not I_65909 (I1122984,I1122976);
nor I_65910 (I1122546,I1122984,I1122789);
nand I_65911 (I1123015,I1122984,I1122634);
not I_65912 (I1123032,I1394580);
nand I_65913 (I1123049,I1123032,I1122738);
nand I_65914 (I1123066,I1122984,I1123049);
nand I_65915 (I1122537,I1123066,I1123015);
nand I_65916 (I1122534,I1123049,I1122933);
not I_65917 (I1123138,I2514);
DFFARX1 I_65918 (I622641,I2507,I1123138,I1123164,);
and I_65919 (I1123172,I1123164,I622629);
DFFARX1 I_65920 (I1123172,I2507,I1123138,I1123121,);
DFFARX1 I_65921 (I622644,I2507,I1123138,I1123212,);
not I_65922 (I1123220,I622635);
not I_65923 (I1123237,I622626);
nand I_65924 (I1123254,I1123237,I1123220);
nor I_65925 (I1123109,I1123212,I1123254);
DFFARX1 I_65926 (I1123254,I2507,I1123138,I1123294,);
not I_65927 (I1123130,I1123294);
not I_65928 (I1123316,I622632);
nand I_65929 (I1123333,I1123237,I1123316);
DFFARX1 I_65930 (I1123333,I2507,I1123138,I1123359,);
not I_65931 (I1123367,I1123359);
not I_65932 (I1123384,I622647);
nand I_65933 (I1123401,I1123384,I622650);
and I_65934 (I1123418,I1123220,I1123401);
nor I_65935 (I1123435,I1123333,I1123418);
DFFARX1 I_65936 (I1123435,I2507,I1123138,I1123106,);
DFFARX1 I_65937 (I1123418,I2507,I1123138,I1123127,);
nor I_65938 (I1123480,I622647,I622626);
nor I_65939 (I1123118,I1123333,I1123480);
or I_65940 (I1123511,I622647,I622626);
nor I_65941 (I1123528,I622638,I622629);
DFFARX1 I_65942 (I1123528,I2507,I1123138,I1123554,);
not I_65943 (I1123562,I1123554);
nor I_65944 (I1123124,I1123562,I1123367);
nand I_65945 (I1123593,I1123562,I1123212);
not I_65946 (I1123610,I622638);
nand I_65947 (I1123627,I1123610,I1123316);
nand I_65948 (I1123644,I1123562,I1123627);
nand I_65949 (I1123115,I1123644,I1123593);
nand I_65950 (I1123112,I1123627,I1123511);
not I_65951 (I1123716,I2514);
DFFARX1 I_65952 (I169865,I2507,I1123716,I1123742,);
and I_65953 (I1123750,I1123742,I169868);
DFFARX1 I_65954 (I1123750,I2507,I1123716,I1123699,);
DFFARX1 I_65955 (I169868,I2507,I1123716,I1123790,);
not I_65956 (I1123798,I169883);
not I_65957 (I1123815,I169889);
nand I_65958 (I1123832,I1123815,I1123798);
nor I_65959 (I1123687,I1123790,I1123832);
DFFARX1 I_65960 (I1123832,I2507,I1123716,I1123872,);
not I_65961 (I1123708,I1123872);
not I_65962 (I1123894,I169877);
nand I_65963 (I1123911,I1123815,I1123894);
DFFARX1 I_65964 (I1123911,I2507,I1123716,I1123937,);
not I_65965 (I1123945,I1123937);
not I_65966 (I1123962,I169874);
nand I_65967 (I1123979,I1123962,I169871);
and I_65968 (I1123996,I1123798,I1123979);
nor I_65969 (I1124013,I1123911,I1123996);
DFFARX1 I_65970 (I1124013,I2507,I1123716,I1123684,);
DFFARX1 I_65971 (I1123996,I2507,I1123716,I1123705,);
nor I_65972 (I1124058,I169874,I169865);
nor I_65973 (I1123696,I1123911,I1124058);
or I_65974 (I1124089,I169874,I169865);
nor I_65975 (I1124106,I169880,I169886);
DFFARX1 I_65976 (I1124106,I2507,I1123716,I1124132,);
not I_65977 (I1124140,I1124132);
nor I_65978 (I1123702,I1124140,I1123945);
nand I_65979 (I1124171,I1124140,I1123790);
not I_65980 (I1124188,I169880);
nand I_65981 (I1124205,I1124188,I1123894);
nand I_65982 (I1124222,I1124140,I1124205);
nand I_65983 (I1123693,I1124222,I1124171);
nand I_65984 (I1123690,I1124205,I1124089);
not I_65985 (I1124294,I2514);
DFFARX1 I_65986 (I133934,I2507,I1124294,I1124320,);
and I_65987 (I1124328,I1124320,I133910);
DFFARX1 I_65988 (I1124328,I2507,I1124294,I1124277,);
DFFARX1 I_65989 (I133928,I2507,I1124294,I1124368,);
not I_65990 (I1124376,I133916);
not I_65991 (I1124393,I133913);
nand I_65992 (I1124410,I1124393,I1124376);
nor I_65993 (I1124265,I1124368,I1124410);
DFFARX1 I_65994 (I1124410,I2507,I1124294,I1124450,);
not I_65995 (I1124286,I1124450);
not I_65996 (I1124472,I133922);
nand I_65997 (I1124489,I1124393,I1124472);
DFFARX1 I_65998 (I1124489,I2507,I1124294,I1124515,);
not I_65999 (I1124523,I1124515);
not I_66000 (I1124540,I133913);
nand I_66001 (I1124557,I1124540,I133931);
and I_66002 (I1124574,I1124376,I1124557);
nor I_66003 (I1124591,I1124489,I1124574);
DFFARX1 I_66004 (I1124591,I2507,I1124294,I1124262,);
DFFARX1 I_66005 (I1124574,I2507,I1124294,I1124283,);
nor I_66006 (I1124636,I133913,I133925);
nor I_66007 (I1124274,I1124489,I1124636);
or I_66008 (I1124667,I133913,I133925);
nor I_66009 (I1124684,I133919,I133910);
DFFARX1 I_66010 (I1124684,I2507,I1124294,I1124710,);
not I_66011 (I1124718,I1124710);
nor I_66012 (I1124280,I1124718,I1124523);
nand I_66013 (I1124749,I1124718,I1124368);
not I_66014 (I1124766,I133919);
nand I_66015 (I1124783,I1124766,I1124472);
nand I_66016 (I1124800,I1124718,I1124783);
nand I_66017 (I1124271,I1124800,I1124749);
nand I_66018 (I1124268,I1124783,I1124667);
not I_66019 (I1124872,I2514);
DFFARX1 I_66020 (I541692,I2507,I1124872,I1124898,);
and I_66021 (I1124906,I1124898,I541707);
DFFARX1 I_66022 (I1124906,I2507,I1124872,I1124855,);
DFFARX1 I_66023 (I541698,I2507,I1124872,I1124946,);
not I_66024 (I1124954,I541692);
not I_66025 (I1124971,I541710);
nand I_66026 (I1124988,I1124971,I1124954);
nor I_66027 (I1124843,I1124946,I1124988);
DFFARX1 I_66028 (I1124988,I2507,I1124872,I1125028,);
not I_66029 (I1124864,I1125028);
not I_66030 (I1125050,I541701);
nand I_66031 (I1125067,I1124971,I1125050);
DFFARX1 I_66032 (I1125067,I2507,I1124872,I1125093,);
not I_66033 (I1125101,I1125093);
not I_66034 (I1125118,I541713);
nand I_66035 (I1125135,I1125118,I541689);
and I_66036 (I1125152,I1124954,I1125135);
nor I_66037 (I1125169,I1125067,I1125152);
DFFARX1 I_66038 (I1125169,I2507,I1124872,I1124840,);
DFFARX1 I_66039 (I1125152,I2507,I1124872,I1124861,);
nor I_66040 (I1125214,I541713,I541689);
nor I_66041 (I1124852,I1125067,I1125214);
or I_66042 (I1125245,I541713,I541689);
nor I_66043 (I1125262,I541695,I541704);
DFFARX1 I_66044 (I1125262,I2507,I1124872,I1125288,);
not I_66045 (I1125296,I1125288);
nor I_66046 (I1124858,I1125296,I1125101);
nand I_66047 (I1125327,I1125296,I1124946);
not I_66048 (I1125344,I541695);
nand I_66049 (I1125361,I1125344,I1125050);
nand I_66050 (I1125378,I1125296,I1125361);
nand I_66051 (I1124849,I1125378,I1125327);
nand I_66052 (I1124846,I1125361,I1125245);
not I_66053 (I1125450,I2514);
DFFARX1 I_66054 (I423471,I2507,I1125450,I1125476,);
and I_66055 (I1125484,I1125476,I423486);
DFFARX1 I_66056 (I1125484,I2507,I1125450,I1125433,);
DFFARX1 I_66057 (I423489,I2507,I1125450,I1125524,);
not I_66058 (I1125532,I423483);
not I_66059 (I1125549,I423498);
nand I_66060 (I1125566,I1125549,I1125532);
nor I_66061 (I1125421,I1125524,I1125566);
DFFARX1 I_66062 (I1125566,I2507,I1125450,I1125606,);
not I_66063 (I1125442,I1125606);
not I_66064 (I1125628,I423474);
nand I_66065 (I1125645,I1125549,I1125628);
DFFARX1 I_66066 (I1125645,I2507,I1125450,I1125671,);
not I_66067 (I1125679,I1125671);
not I_66068 (I1125696,I423477);
nand I_66069 (I1125713,I1125696,I423471);
and I_66070 (I1125730,I1125532,I1125713);
nor I_66071 (I1125747,I1125645,I1125730);
DFFARX1 I_66072 (I1125747,I2507,I1125450,I1125418,);
DFFARX1 I_66073 (I1125730,I2507,I1125450,I1125439,);
nor I_66074 (I1125792,I423477,I423480);
nor I_66075 (I1125430,I1125645,I1125792);
or I_66076 (I1125823,I423477,I423480);
nor I_66077 (I1125840,I423495,I423492);
DFFARX1 I_66078 (I1125840,I2507,I1125450,I1125866,);
not I_66079 (I1125874,I1125866);
nor I_66080 (I1125436,I1125874,I1125679);
nand I_66081 (I1125905,I1125874,I1125524);
not I_66082 (I1125922,I423495);
nand I_66083 (I1125939,I1125922,I1125628);
nand I_66084 (I1125956,I1125874,I1125939);
nand I_66085 (I1125427,I1125956,I1125905);
nand I_66086 (I1125424,I1125939,I1125823);
not I_66087 (I1126028,I2514);
DFFARX1 I_66088 (I331375,I2507,I1126028,I1126054,);
and I_66089 (I1126062,I1126054,I331360);
DFFARX1 I_66090 (I1126062,I2507,I1126028,I1126011,);
DFFARX1 I_66091 (I331366,I2507,I1126028,I1126102,);
not I_66092 (I1126110,I331348);
not I_66093 (I1126127,I331369);
nand I_66094 (I1126144,I1126127,I1126110);
nor I_66095 (I1125999,I1126102,I1126144);
DFFARX1 I_66096 (I1126144,I2507,I1126028,I1126184,);
not I_66097 (I1126020,I1126184);
not I_66098 (I1126206,I331372);
nand I_66099 (I1126223,I1126127,I1126206);
DFFARX1 I_66100 (I1126223,I2507,I1126028,I1126249,);
not I_66101 (I1126257,I1126249);
not I_66102 (I1126274,I331363);
nand I_66103 (I1126291,I1126274,I331351);
and I_66104 (I1126308,I1126110,I1126291);
nor I_66105 (I1126325,I1126223,I1126308);
DFFARX1 I_66106 (I1126325,I2507,I1126028,I1125996,);
DFFARX1 I_66107 (I1126308,I2507,I1126028,I1126017,);
nor I_66108 (I1126370,I331363,I331357);
nor I_66109 (I1126008,I1126223,I1126370);
or I_66110 (I1126401,I331363,I331357);
nor I_66111 (I1126418,I331354,I331348);
DFFARX1 I_66112 (I1126418,I2507,I1126028,I1126444,);
not I_66113 (I1126452,I1126444);
nor I_66114 (I1126014,I1126452,I1126257);
nand I_66115 (I1126483,I1126452,I1126102);
not I_66116 (I1126500,I331354);
nand I_66117 (I1126517,I1126500,I1126206);
nand I_66118 (I1126534,I1126452,I1126517);
nand I_66119 (I1126005,I1126534,I1126483);
nand I_66120 (I1126002,I1126517,I1126401);
not I_66121 (I1126606,I2514);
DFFARX1 I_66122 (I500042,I2507,I1126606,I1126632,);
and I_66123 (I1126640,I1126632,I500057);
DFFARX1 I_66124 (I1126640,I2507,I1126606,I1126589,);
DFFARX1 I_66125 (I500048,I2507,I1126606,I1126680,);
not I_66126 (I1126688,I500042);
not I_66127 (I1126705,I500060);
nand I_66128 (I1126722,I1126705,I1126688);
nor I_66129 (I1126577,I1126680,I1126722);
DFFARX1 I_66130 (I1126722,I2507,I1126606,I1126762,);
not I_66131 (I1126598,I1126762);
not I_66132 (I1126784,I500051);
nand I_66133 (I1126801,I1126705,I1126784);
DFFARX1 I_66134 (I1126801,I2507,I1126606,I1126827,);
not I_66135 (I1126835,I1126827);
not I_66136 (I1126852,I500063);
nand I_66137 (I1126869,I1126852,I500039);
and I_66138 (I1126886,I1126688,I1126869);
nor I_66139 (I1126903,I1126801,I1126886);
DFFARX1 I_66140 (I1126903,I2507,I1126606,I1126574,);
DFFARX1 I_66141 (I1126886,I2507,I1126606,I1126595,);
nor I_66142 (I1126948,I500063,I500039);
nor I_66143 (I1126586,I1126801,I1126948);
or I_66144 (I1126979,I500063,I500039);
nor I_66145 (I1126996,I500045,I500054);
DFFARX1 I_66146 (I1126996,I2507,I1126606,I1127022,);
not I_66147 (I1127030,I1127022);
nor I_66148 (I1126592,I1127030,I1126835);
nand I_66149 (I1127061,I1127030,I1126680);
not I_66150 (I1127078,I500045);
nand I_66151 (I1127095,I1127078,I1126784);
nand I_66152 (I1127112,I1127030,I1127095);
nand I_66153 (I1126583,I1127112,I1127061);
nand I_66154 (I1126580,I1127095,I1126979);
not I_66155 (I1127184,I2514);
DFFARX1 I_66156 (I738241,I2507,I1127184,I1127210,);
and I_66157 (I1127218,I1127210,I738229);
DFFARX1 I_66158 (I1127218,I2507,I1127184,I1127167,);
DFFARX1 I_66159 (I738232,I2507,I1127184,I1127258,);
not I_66160 (I1127266,I738226);
not I_66161 (I1127283,I738250);
nand I_66162 (I1127300,I1127283,I1127266);
nor I_66163 (I1127155,I1127258,I1127300);
DFFARX1 I_66164 (I1127300,I2507,I1127184,I1127340,);
not I_66165 (I1127176,I1127340);
not I_66166 (I1127362,I738238);
nand I_66167 (I1127379,I1127283,I1127362);
DFFARX1 I_66168 (I1127379,I2507,I1127184,I1127405,);
not I_66169 (I1127413,I1127405);
not I_66170 (I1127430,I738247);
nand I_66171 (I1127447,I1127430,I738244);
and I_66172 (I1127464,I1127266,I1127447);
nor I_66173 (I1127481,I1127379,I1127464);
DFFARX1 I_66174 (I1127481,I2507,I1127184,I1127152,);
DFFARX1 I_66175 (I1127464,I2507,I1127184,I1127173,);
nor I_66176 (I1127526,I738247,I738235);
nor I_66177 (I1127164,I1127379,I1127526);
or I_66178 (I1127557,I738247,I738235);
nor I_66179 (I1127574,I738226,I738229);
DFFARX1 I_66180 (I1127574,I2507,I1127184,I1127600,);
not I_66181 (I1127608,I1127600);
nor I_66182 (I1127170,I1127608,I1127413);
nand I_66183 (I1127639,I1127608,I1127258);
not I_66184 (I1127656,I738226);
nand I_66185 (I1127673,I1127656,I1127362);
nand I_66186 (I1127690,I1127608,I1127673);
nand I_66187 (I1127161,I1127690,I1127639);
nand I_66188 (I1127158,I1127673,I1127557);
not I_66189 (I1127762,I2514);
DFFARX1 I_66190 (I1377334,I2507,I1127762,I1127788,);
and I_66191 (I1127796,I1127788,I1377316);
DFFARX1 I_66192 (I1127796,I2507,I1127762,I1127745,);
DFFARX1 I_66193 (I1377307,I2507,I1127762,I1127836,);
not I_66194 (I1127844,I1377322);
not I_66195 (I1127861,I1377310);
nand I_66196 (I1127878,I1127861,I1127844);
nor I_66197 (I1127733,I1127836,I1127878);
DFFARX1 I_66198 (I1127878,I2507,I1127762,I1127918,);
not I_66199 (I1127754,I1127918);
not I_66200 (I1127940,I1377319);
nand I_66201 (I1127957,I1127861,I1127940);
DFFARX1 I_66202 (I1127957,I2507,I1127762,I1127983,);
not I_66203 (I1127991,I1127983);
not I_66204 (I1128008,I1377328);
nand I_66205 (I1128025,I1128008,I1377307);
and I_66206 (I1128042,I1127844,I1128025);
nor I_66207 (I1128059,I1127957,I1128042);
DFFARX1 I_66208 (I1128059,I2507,I1127762,I1127730,);
DFFARX1 I_66209 (I1128042,I2507,I1127762,I1127751,);
nor I_66210 (I1128104,I1377328,I1377331);
nor I_66211 (I1127742,I1127957,I1128104);
or I_66212 (I1128135,I1377328,I1377331);
nor I_66213 (I1128152,I1377325,I1377313);
DFFARX1 I_66214 (I1128152,I2507,I1127762,I1128178,);
not I_66215 (I1128186,I1128178);
nor I_66216 (I1127748,I1128186,I1127991);
nand I_66217 (I1128217,I1128186,I1127836);
not I_66218 (I1128234,I1377325);
nand I_66219 (I1128251,I1128234,I1127940);
nand I_66220 (I1128268,I1128186,I1128251);
nand I_66221 (I1127739,I1128268,I1128217);
nand I_66222 (I1127736,I1128251,I1128135);
not I_66223 (I1128340,I2514);
DFFARX1 I_66224 (I188905,I2507,I1128340,I1128366,);
and I_66225 (I1128374,I1128366,I188908);
DFFARX1 I_66226 (I1128374,I2507,I1128340,I1128323,);
DFFARX1 I_66227 (I188908,I2507,I1128340,I1128414,);
not I_66228 (I1128422,I188923);
not I_66229 (I1128439,I188929);
nand I_66230 (I1128456,I1128439,I1128422);
nor I_66231 (I1128311,I1128414,I1128456);
DFFARX1 I_66232 (I1128456,I2507,I1128340,I1128496,);
not I_66233 (I1128332,I1128496);
not I_66234 (I1128518,I188917);
nand I_66235 (I1128535,I1128439,I1128518);
DFFARX1 I_66236 (I1128535,I2507,I1128340,I1128561,);
not I_66237 (I1128569,I1128561);
not I_66238 (I1128586,I188914);
nand I_66239 (I1128603,I1128586,I188911);
and I_66240 (I1128620,I1128422,I1128603);
nor I_66241 (I1128637,I1128535,I1128620);
DFFARX1 I_66242 (I1128637,I2507,I1128340,I1128308,);
DFFARX1 I_66243 (I1128620,I2507,I1128340,I1128329,);
nor I_66244 (I1128682,I188914,I188905);
nor I_66245 (I1128320,I1128535,I1128682);
or I_66246 (I1128713,I188914,I188905);
nor I_66247 (I1128730,I188920,I188926);
DFFARX1 I_66248 (I1128730,I2507,I1128340,I1128756,);
not I_66249 (I1128764,I1128756);
nor I_66250 (I1128326,I1128764,I1128569);
nand I_66251 (I1128795,I1128764,I1128414);
not I_66252 (I1128812,I188920);
nand I_66253 (I1128829,I1128812,I1128518);
nand I_66254 (I1128846,I1128764,I1128829);
nand I_66255 (I1128317,I1128846,I1128795);
nand I_66256 (I1128314,I1128829,I1128713);
not I_66257 (I1128918,I2514);
DFFARX1 I_66258 (I1364839,I2507,I1128918,I1128944,);
and I_66259 (I1128952,I1128944,I1364821);
DFFARX1 I_66260 (I1128952,I2507,I1128918,I1128901,);
DFFARX1 I_66261 (I1364812,I2507,I1128918,I1128992,);
not I_66262 (I1129000,I1364827);
not I_66263 (I1129017,I1364815);
nand I_66264 (I1129034,I1129017,I1129000);
nor I_66265 (I1128889,I1128992,I1129034);
DFFARX1 I_66266 (I1129034,I2507,I1128918,I1129074,);
not I_66267 (I1128910,I1129074);
not I_66268 (I1129096,I1364824);
nand I_66269 (I1129113,I1129017,I1129096);
DFFARX1 I_66270 (I1129113,I2507,I1128918,I1129139,);
not I_66271 (I1129147,I1129139);
not I_66272 (I1129164,I1364833);
nand I_66273 (I1129181,I1129164,I1364812);
and I_66274 (I1129198,I1129000,I1129181);
nor I_66275 (I1129215,I1129113,I1129198);
DFFARX1 I_66276 (I1129215,I2507,I1128918,I1128886,);
DFFARX1 I_66277 (I1129198,I2507,I1128918,I1128907,);
nor I_66278 (I1129260,I1364833,I1364836);
nor I_66279 (I1128898,I1129113,I1129260);
or I_66280 (I1129291,I1364833,I1364836);
nor I_66281 (I1129308,I1364830,I1364818);
DFFARX1 I_66282 (I1129308,I2507,I1128918,I1129334,);
not I_66283 (I1129342,I1129334);
nor I_66284 (I1128904,I1129342,I1129147);
nand I_66285 (I1129373,I1129342,I1128992);
not I_66286 (I1129390,I1364830);
nand I_66287 (I1129407,I1129390,I1129096);
nand I_66288 (I1129424,I1129342,I1129407);
nand I_66289 (I1128895,I1129424,I1129373);
nand I_66290 (I1128892,I1129407,I1129291);
not I_66291 (I1129496,I2514);
DFFARX1 I_66292 (I733039,I2507,I1129496,I1129522,);
and I_66293 (I1129530,I1129522,I733027);
DFFARX1 I_66294 (I1129530,I2507,I1129496,I1129479,);
DFFARX1 I_66295 (I733030,I2507,I1129496,I1129570,);
not I_66296 (I1129578,I733024);
not I_66297 (I1129595,I733048);
nand I_66298 (I1129612,I1129595,I1129578);
nor I_66299 (I1129467,I1129570,I1129612);
DFFARX1 I_66300 (I1129612,I2507,I1129496,I1129652,);
not I_66301 (I1129488,I1129652);
not I_66302 (I1129674,I733036);
nand I_66303 (I1129691,I1129595,I1129674);
DFFARX1 I_66304 (I1129691,I2507,I1129496,I1129717,);
not I_66305 (I1129725,I1129717);
not I_66306 (I1129742,I733045);
nand I_66307 (I1129759,I1129742,I733042);
and I_66308 (I1129776,I1129578,I1129759);
nor I_66309 (I1129793,I1129691,I1129776);
DFFARX1 I_66310 (I1129793,I2507,I1129496,I1129464,);
DFFARX1 I_66311 (I1129776,I2507,I1129496,I1129485,);
nor I_66312 (I1129838,I733045,I733033);
nor I_66313 (I1129476,I1129691,I1129838);
or I_66314 (I1129869,I733045,I733033);
nor I_66315 (I1129886,I733024,I733027);
DFFARX1 I_66316 (I1129886,I2507,I1129496,I1129912,);
not I_66317 (I1129920,I1129912);
nor I_66318 (I1129482,I1129920,I1129725);
nand I_66319 (I1129951,I1129920,I1129570);
not I_66320 (I1129968,I733024);
nand I_66321 (I1129985,I1129968,I1129674);
nand I_66322 (I1130002,I1129920,I1129985);
nand I_66323 (I1129473,I1130002,I1129951);
nand I_66324 (I1129470,I1129985,I1129869);
not I_66325 (I1130074,I2514);
DFFARX1 I_66326 (I888223,I2507,I1130074,I1130100,);
and I_66327 (I1130108,I1130100,I888217);
DFFARX1 I_66328 (I1130108,I2507,I1130074,I1130057,);
DFFARX1 I_66329 (I888235,I2507,I1130074,I1130148,);
not I_66330 (I1130156,I888226);
not I_66331 (I1130173,I888238);
nand I_66332 (I1130190,I1130173,I1130156);
nor I_66333 (I1130045,I1130148,I1130190);
DFFARX1 I_66334 (I1130190,I2507,I1130074,I1130230,);
not I_66335 (I1130066,I1130230);
not I_66336 (I1130252,I888244);
nand I_66337 (I1130269,I1130173,I1130252);
DFFARX1 I_66338 (I1130269,I2507,I1130074,I1130295,);
not I_66339 (I1130303,I1130295);
not I_66340 (I1130320,I888220);
nand I_66341 (I1130337,I1130320,I888241);
and I_66342 (I1130354,I1130156,I1130337);
nor I_66343 (I1130371,I1130269,I1130354);
DFFARX1 I_66344 (I1130371,I2507,I1130074,I1130042,);
DFFARX1 I_66345 (I1130354,I2507,I1130074,I1130063,);
nor I_66346 (I1130416,I888220,I888232);
nor I_66347 (I1130054,I1130269,I1130416);
or I_66348 (I1130447,I888220,I888232);
nor I_66349 (I1130464,I888217,I888229);
DFFARX1 I_66350 (I1130464,I2507,I1130074,I1130490,);
not I_66351 (I1130498,I1130490);
nor I_66352 (I1130060,I1130498,I1130303);
nand I_66353 (I1130529,I1130498,I1130148);
not I_66354 (I1130546,I888217);
nand I_66355 (I1130563,I1130546,I1130252);
nand I_66356 (I1130580,I1130498,I1130563);
nand I_66357 (I1130051,I1130580,I1130529);
nand I_66358 (I1130048,I1130563,I1130447);
not I_66359 (I1130652,I2514);
DFFARX1 I_66360 (I34307,I2507,I1130652,I1130678,);
and I_66361 (I1130686,I1130678,I34310);
DFFARX1 I_66362 (I1130686,I2507,I1130652,I1130635,);
DFFARX1 I_66363 (I34310,I2507,I1130652,I1130726,);
not I_66364 (I1130734,I34313);
not I_66365 (I1130751,I34328);
nand I_66366 (I1130768,I1130751,I1130734);
nor I_66367 (I1130623,I1130726,I1130768);
DFFARX1 I_66368 (I1130768,I2507,I1130652,I1130808,);
not I_66369 (I1130644,I1130808);
not I_66370 (I1130830,I34322);
nand I_66371 (I1130847,I1130751,I1130830);
DFFARX1 I_66372 (I1130847,I2507,I1130652,I1130873,);
not I_66373 (I1130881,I1130873);
not I_66374 (I1130898,I34325);
nand I_66375 (I1130915,I1130898,I34307);
and I_66376 (I1130932,I1130734,I1130915);
nor I_66377 (I1130949,I1130847,I1130932);
DFFARX1 I_66378 (I1130949,I2507,I1130652,I1130620,);
DFFARX1 I_66379 (I1130932,I2507,I1130652,I1130641,);
nor I_66380 (I1130994,I34325,I34319);
nor I_66381 (I1130632,I1130847,I1130994);
or I_66382 (I1131025,I34325,I34319);
nor I_66383 (I1131042,I34316,I34331);
DFFARX1 I_66384 (I1131042,I2507,I1130652,I1131068,);
not I_66385 (I1131076,I1131068);
nor I_66386 (I1130638,I1131076,I1130881);
nand I_66387 (I1131107,I1131076,I1130726);
not I_66388 (I1131124,I34316);
nand I_66389 (I1131141,I1131124,I1130830);
nand I_66390 (I1131158,I1131076,I1131141);
nand I_66391 (I1130629,I1131158,I1131107);
nand I_66392 (I1130626,I1131141,I1131025);
not I_66393 (I1131230,I2514);
DFFARX1 I_66394 (I1259402,I2507,I1131230,I1131256,);
and I_66395 (I1131264,I1131256,I1259384);
DFFARX1 I_66396 (I1131264,I2507,I1131230,I1131213,);
DFFARX1 I_66397 (I1259393,I2507,I1131230,I1131304,);
not I_66398 (I1131312,I1259378);
not I_66399 (I1131329,I1259390);
nand I_66400 (I1131346,I1131329,I1131312);
nor I_66401 (I1131201,I1131304,I1131346);
DFFARX1 I_66402 (I1131346,I2507,I1131230,I1131386,);
not I_66403 (I1131222,I1131386);
not I_66404 (I1131408,I1259381);
nand I_66405 (I1131425,I1131329,I1131408);
DFFARX1 I_66406 (I1131425,I2507,I1131230,I1131451,);
not I_66407 (I1131459,I1131451);
not I_66408 (I1131476,I1259378);
nand I_66409 (I1131493,I1131476,I1259381);
and I_66410 (I1131510,I1131312,I1131493);
nor I_66411 (I1131527,I1131425,I1131510);
DFFARX1 I_66412 (I1131527,I2507,I1131230,I1131198,);
DFFARX1 I_66413 (I1131510,I2507,I1131230,I1131219,);
nor I_66414 (I1131572,I1259378,I1259399);
nor I_66415 (I1131210,I1131425,I1131572);
or I_66416 (I1131603,I1259378,I1259399);
nor I_66417 (I1131620,I1259387,I1259396);
DFFARX1 I_66418 (I1131620,I2507,I1131230,I1131646,);
not I_66419 (I1131654,I1131646);
nor I_66420 (I1131216,I1131654,I1131459);
nand I_66421 (I1131685,I1131654,I1131304);
not I_66422 (I1131702,I1259387);
nand I_66423 (I1131719,I1131702,I1131408);
nand I_66424 (I1131736,I1131654,I1131719);
nand I_66425 (I1131207,I1131736,I1131685);
nand I_66426 (I1131204,I1131719,I1131603);
not I_66427 (I1131808,I2514);
DFFARX1 I_66428 (I251271,I2507,I1131808,I1131834,);
and I_66429 (I1131842,I1131834,I251256);
DFFARX1 I_66430 (I1131842,I2507,I1131808,I1131791,);
DFFARX1 I_66431 (I251262,I2507,I1131808,I1131882,);
not I_66432 (I1131890,I251244);
not I_66433 (I1131907,I251265);
nand I_66434 (I1131924,I1131907,I1131890);
nor I_66435 (I1131779,I1131882,I1131924);
DFFARX1 I_66436 (I1131924,I2507,I1131808,I1131964,);
not I_66437 (I1131800,I1131964);
not I_66438 (I1131986,I251268);
nand I_66439 (I1132003,I1131907,I1131986);
DFFARX1 I_66440 (I1132003,I2507,I1131808,I1132029,);
not I_66441 (I1132037,I1132029);
not I_66442 (I1132054,I251259);
nand I_66443 (I1132071,I1132054,I251247);
and I_66444 (I1132088,I1131890,I1132071);
nor I_66445 (I1132105,I1132003,I1132088);
DFFARX1 I_66446 (I1132105,I2507,I1131808,I1131776,);
DFFARX1 I_66447 (I1132088,I2507,I1131808,I1131797,);
nor I_66448 (I1132150,I251259,I251253);
nor I_66449 (I1131788,I1132003,I1132150);
or I_66450 (I1132181,I251259,I251253);
nor I_66451 (I1132198,I251250,I251244);
DFFARX1 I_66452 (I1132198,I2507,I1131808,I1132224,);
not I_66453 (I1132232,I1132224);
nor I_66454 (I1131794,I1132232,I1132037);
nand I_66455 (I1132263,I1132232,I1131882);
not I_66456 (I1132280,I251250);
nand I_66457 (I1132297,I1132280,I1131986);
nand I_66458 (I1132314,I1132232,I1132297);
nand I_66459 (I1131785,I1132314,I1132263);
nand I_66460 (I1131782,I1132297,I1132181);
not I_66461 (I1132386,I2514);
DFFARX1 I_66462 (I171055,I2507,I1132386,I1132412,);
and I_66463 (I1132420,I1132412,I171058);
DFFARX1 I_66464 (I1132420,I2507,I1132386,I1132369,);
DFFARX1 I_66465 (I171058,I2507,I1132386,I1132460,);
not I_66466 (I1132468,I171073);
not I_66467 (I1132485,I171079);
nand I_66468 (I1132502,I1132485,I1132468);
nor I_66469 (I1132357,I1132460,I1132502);
DFFARX1 I_66470 (I1132502,I2507,I1132386,I1132542,);
not I_66471 (I1132378,I1132542);
not I_66472 (I1132564,I171067);
nand I_66473 (I1132581,I1132485,I1132564);
DFFARX1 I_66474 (I1132581,I2507,I1132386,I1132607,);
not I_66475 (I1132615,I1132607);
not I_66476 (I1132632,I171064);
nand I_66477 (I1132649,I1132632,I171061);
and I_66478 (I1132666,I1132468,I1132649);
nor I_66479 (I1132683,I1132581,I1132666);
DFFARX1 I_66480 (I1132683,I2507,I1132386,I1132354,);
DFFARX1 I_66481 (I1132666,I2507,I1132386,I1132375,);
nor I_66482 (I1132728,I171064,I171055);
nor I_66483 (I1132366,I1132581,I1132728);
or I_66484 (I1132759,I171064,I171055);
nor I_66485 (I1132776,I171070,I171076);
DFFARX1 I_66486 (I1132776,I2507,I1132386,I1132802,);
not I_66487 (I1132810,I1132802);
nor I_66488 (I1132372,I1132810,I1132615);
nand I_66489 (I1132841,I1132810,I1132460);
not I_66490 (I1132858,I171070);
nand I_66491 (I1132875,I1132858,I1132564);
nand I_66492 (I1132892,I1132810,I1132875);
nand I_66493 (I1132363,I1132892,I1132841);
nand I_66494 (I1132360,I1132875,I1132759);
not I_66495 (I1132964,I2514);
DFFARX1 I_66496 (I817534,I2507,I1132964,I1132990,);
and I_66497 (I1132998,I1132990,I817540);
DFFARX1 I_66498 (I1132998,I2507,I1132964,I1132947,);
DFFARX1 I_66499 (I817546,I2507,I1132964,I1133038,);
not I_66500 (I1133046,I817531);
not I_66501 (I1133063,I817531);
nand I_66502 (I1133080,I1133063,I1133046);
nor I_66503 (I1132935,I1133038,I1133080);
DFFARX1 I_66504 (I1133080,I2507,I1132964,I1133120,);
not I_66505 (I1132956,I1133120);
not I_66506 (I1133142,I817549);
nand I_66507 (I1133159,I1133063,I1133142);
DFFARX1 I_66508 (I1133159,I2507,I1132964,I1133185,);
not I_66509 (I1133193,I1133185);
not I_66510 (I1133210,I817543);
nand I_66511 (I1133227,I1133210,I817534);
and I_66512 (I1133244,I1133046,I1133227);
nor I_66513 (I1133261,I1133159,I1133244);
DFFARX1 I_66514 (I1133261,I2507,I1132964,I1132932,);
DFFARX1 I_66515 (I1133244,I2507,I1132964,I1132953,);
nor I_66516 (I1133306,I817543,I817552);
nor I_66517 (I1132944,I1133159,I1133306);
or I_66518 (I1133337,I817543,I817552);
nor I_66519 (I1133354,I817537,I817537);
DFFARX1 I_66520 (I1133354,I2507,I1132964,I1133380,);
not I_66521 (I1133388,I1133380);
nor I_66522 (I1132950,I1133388,I1133193);
nand I_66523 (I1133419,I1133388,I1133038);
not I_66524 (I1133436,I817537);
nand I_66525 (I1133453,I1133436,I1133142);
nand I_66526 (I1133470,I1133388,I1133453);
nand I_66527 (I1132941,I1133470,I1133419);
nand I_66528 (I1132938,I1133453,I1133337);
not I_66529 (I1133542,I2514);
DFFARX1 I_66530 (I329267,I2507,I1133542,I1133568,);
and I_66531 (I1133576,I1133568,I329252);
DFFARX1 I_66532 (I1133576,I2507,I1133542,I1133525,);
DFFARX1 I_66533 (I329258,I2507,I1133542,I1133616,);
not I_66534 (I1133624,I329240);
not I_66535 (I1133641,I329261);
nand I_66536 (I1133658,I1133641,I1133624);
nor I_66537 (I1133513,I1133616,I1133658);
DFFARX1 I_66538 (I1133658,I2507,I1133542,I1133698,);
not I_66539 (I1133534,I1133698);
not I_66540 (I1133720,I329264);
nand I_66541 (I1133737,I1133641,I1133720);
DFFARX1 I_66542 (I1133737,I2507,I1133542,I1133763,);
not I_66543 (I1133771,I1133763);
not I_66544 (I1133788,I329255);
nand I_66545 (I1133805,I1133788,I329243);
and I_66546 (I1133822,I1133624,I1133805);
nor I_66547 (I1133839,I1133737,I1133822);
DFFARX1 I_66548 (I1133839,I2507,I1133542,I1133510,);
DFFARX1 I_66549 (I1133822,I2507,I1133542,I1133531,);
nor I_66550 (I1133884,I329255,I329249);
nor I_66551 (I1133522,I1133737,I1133884);
or I_66552 (I1133915,I329255,I329249);
nor I_66553 (I1133932,I329246,I329240);
DFFARX1 I_66554 (I1133932,I2507,I1133542,I1133958,);
not I_66555 (I1133966,I1133958);
nor I_66556 (I1133528,I1133966,I1133771);
nand I_66557 (I1133997,I1133966,I1133616);
not I_66558 (I1134014,I329246);
nand I_66559 (I1134031,I1134014,I1133720);
nand I_66560 (I1134048,I1133966,I1134031);
nand I_66561 (I1133519,I1134048,I1133997);
nand I_66562 (I1133516,I1134031,I1133915);
not I_66563 (I1134120,I2514);
DFFARX1 I_66564 (I247810,I2507,I1134120,I1134146,);
and I_66565 (I1134154,I1134146,I247813);
DFFARX1 I_66566 (I1134154,I2507,I1134120,I1134103,);
DFFARX1 I_66567 (I247813,I2507,I1134120,I1134194,);
not I_66568 (I1134202,I247828);
not I_66569 (I1134219,I247834);
nand I_66570 (I1134236,I1134219,I1134202);
nor I_66571 (I1134091,I1134194,I1134236);
DFFARX1 I_66572 (I1134236,I2507,I1134120,I1134276,);
not I_66573 (I1134112,I1134276);
not I_66574 (I1134298,I247822);
nand I_66575 (I1134315,I1134219,I1134298);
DFFARX1 I_66576 (I1134315,I2507,I1134120,I1134341,);
not I_66577 (I1134349,I1134341);
not I_66578 (I1134366,I247819);
nand I_66579 (I1134383,I1134366,I247816);
and I_66580 (I1134400,I1134202,I1134383);
nor I_66581 (I1134417,I1134315,I1134400);
DFFARX1 I_66582 (I1134417,I2507,I1134120,I1134088,);
DFFARX1 I_66583 (I1134400,I2507,I1134120,I1134109,);
nor I_66584 (I1134462,I247819,I247810);
nor I_66585 (I1134100,I1134315,I1134462);
or I_66586 (I1134493,I247819,I247810);
nor I_66587 (I1134510,I247825,I247831);
DFFARX1 I_66588 (I1134510,I2507,I1134120,I1134536,);
not I_66589 (I1134544,I1134536);
nor I_66590 (I1134106,I1134544,I1134349);
nand I_66591 (I1134575,I1134544,I1134194);
not I_66592 (I1134592,I247825);
nand I_66593 (I1134609,I1134592,I1134298);
nand I_66594 (I1134626,I1134544,I1134609);
nand I_66595 (I1134097,I1134626,I1134575);
nand I_66596 (I1134094,I1134609,I1134493);
not I_66597 (I1134698,I2514);
DFFARX1 I_66598 (I1266338,I2507,I1134698,I1134724,);
and I_66599 (I1134732,I1134724,I1266320);
DFFARX1 I_66600 (I1134732,I2507,I1134698,I1134681,);
DFFARX1 I_66601 (I1266329,I2507,I1134698,I1134772,);
not I_66602 (I1134780,I1266314);
not I_66603 (I1134797,I1266326);
nand I_66604 (I1134814,I1134797,I1134780);
nor I_66605 (I1134669,I1134772,I1134814);
DFFARX1 I_66606 (I1134814,I2507,I1134698,I1134854,);
not I_66607 (I1134690,I1134854);
not I_66608 (I1134876,I1266317);
nand I_66609 (I1134893,I1134797,I1134876);
DFFARX1 I_66610 (I1134893,I2507,I1134698,I1134919,);
not I_66611 (I1134927,I1134919);
not I_66612 (I1134944,I1266314);
nand I_66613 (I1134961,I1134944,I1266317);
and I_66614 (I1134978,I1134780,I1134961);
nor I_66615 (I1134995,I1134893,I1134978);
DFFARX1 I_66616 (I1134995,I2507,I1134698,I1134666,);
DFFARX1 I_66617 (I1134978,I2507,I1134698,I1134687,);
nor I_66618 (I1135040,I1266314,I1266335);
nor I_66619 (I1134678,I1134893,I1135040);
or I_66620 (I1135071,I1266314,I1266335);
nor I_66621 (I1135088,I1266323,I1266332);
DFFARX1 I_66622 (I1135088,I2507,I1134698,I1135114,);
not I_66623 (I1135122,I1135114);
nor I_66624 (I1134684,I1135122,I1134927);
nand I_66625 (I1135153,I1135122,I1134772);
not I_66626 (I1135170,I1266323);
nand I_66627 (I1135187,I1135170,I1134876);
nand I_66628 (I1135204,I1135122,I1135187);
nand I_66629 (I1134675,I1135204,I1135153);
nand I_66630 (I1134672,I1135187,I1135071);
not I_66631 (I1135276,I2514);
DFFARX1 I_66632 (I243645,I2507,I1135276,I1135302,);
and I_66633 (I1135310,I1135302,I243648);
DFFARX1 I_66634 (I1135310,I2507,I1135276,I1135259,);
DFFARX1 I_66635 (I243648,I2507,I1135276,I1135350,);
not I_66636 (I1135358,I243663);
not I_66637 (I1135375,I243669);
nand I_66638 (I1135392,I1135375,I1135358);
nor I_66639 (I1135247,I1135350,I1135392);
DFFARX1 I_66640 (I1135392,I2507,I1135276,I1135432,);
not I_66641 (I1135268,I1135432);
not I_66642 (I1135454,I243657);
nand I_66643 (I1135471,I1135375,I1135454);
DFFARX1 I_66644 (I1135471,I2507,I1135276,I1135497,);
not I_66645 (I1135505,I1135497);
not I_66646 (I1135522,I243654);
nand I_66647 (I1135539,I1135522,I243651);
and I_66648 (I1135556,I1135358,I1135539);
nor I_66649 (I1135573,I1135471,I1135556);
DFFARX1 I_66650 (I1135573,I2507,I1135276,I1135244,);
DFFARX1 I_66651 (I1135556,I2507,I1135276,I1135265,);
nor I_66652 (I1135618,I243654,I243645);
nor I_66653 (I1135256,I1135471,I1135618);
or I_66654 (I1135649,I243654,I243645);
nor I_66655 (I1135666,I243660,I243666);
DFFARX1 I_66656 (I1135666,I2507,I1135276,I1135692,);
not I_66657 (I1135700,I1135692);
nor I_66658 (I1135262,I1135700,I1135505);
nand I_66659 (I1135731,I1135700,I1135350);
not I_66660 (I1135748,I243660);
nand I_66661 (I1135765,I1135748,I1135454);
nand I_66662 (I1135782,I1135700,I1135765);
nand I_66663 (I1135253,I1135782,I1135731);
nand I_66664 (I1135250,I1135765,I1135649);
not I_66665 (I1135854,I2514);
DFFARX1 I_66666 (I474063,I2507,I1135854,I1135880,);
and I_66667 (I1135888,I1135880,I474078);
DFFARX1 I_66668 (I1135888,I2507,I1135854,I1135837,);
DFFARX1 I_66669 (I474081,I2507,I1135854,I1135928,);
not I_66670 (I1135936,I474075);
not I_66671 (I1135953,I474090);
nand I_66672 (I1135970,I1135953,I1135936);
nor I_66673 (I1135825,I1135928,I1135970);
DFFARX1 I_66674 (I1135970,I2507,I1135854,I1136010,);
not I_66675 (I1135846,I1136010);
not I_66676 (I1136032,I474066);
nand I_66677 (I1136049,I1135953,I1136032);
DFFARX1 I_66678 (I1136049,I2507,I1135854,I1136075,);
not I_66679 (I1136083,I1136075);
not I_66680 (I1136100,I474069);
nand I_66681 (I1136117,I1136100,I474063);
and I_66682 (I1136134,I1135936,I1136117);
nor I_66683 (I1136151,I1136049,I1136134);
DFFARX1 I_66684 (I1136151,I2507,I1135854,I1135822,);
DFFARX1 I_66685 (I1136134,I2507,I1135854,I1135843,);
nor I_66686 (I1136196,I474069,I474072);
nor I_66687 (I1135834,I1136049,I1136196);
or I_66688 (I1136227,I474069,I474072);
nor I_66689 (I1136244,I474087,I474084);
DFFARX1 I_66690 (I1136244,I2507,I1135854,I1136270,);
not I_66691 (I1136278,I1136270);
nor I_66692 (I1135840,I1136278,I1136083);
nand I_66693 (I1136309,I1136278,I1135928);
not I_66694 (I1136326,I474087);
nand I_66695 (I1136343,I1136326,I1136032);
nand I_66696 (I1136360,I1136278,I1136343);
nand I_66697 (I1135831,I1136360,I1136309);
nand I_66698 (I1135828,I1136343,I1136227);
not I_66699 (I1136432,I2514);
DFFARX1 I_66700 (I177005,I2507,I1136432,I1136458,);
and I_66701 (I1136466,I1136458,I177008);
DFFARX1 I_66702 (I1136466,I2507,I1136432,I1136415,);
DFFARX1 I_66703 (I177008,I2507,I1136432,I1136506,);
not I_66704 (I1136514,I177023);
not I_66705 (I1136531,I177029);
nand I_66706 (I1136548,I1136531,I1136514);
nor I_66707 (I1136403,I1136506,I1136548);
DFFARX1 I_66708 (I1136548,I2507,I1136432,I1136588,);
not I_66709 (I1136424,I1136588);
not I_66710 (I1136610,I177017);
nand I_66711 (I1136627,I1136531,I1136610);
DFFARX1 I_66712 (I1136627,I2507,I1136432,I1136653,);
not I_66713 (I1136661,I1136653);
not I_66714 (I1136678,I177014);
nand I_66715 (I1136695,I1136678,I177011);
and I_66716 (I1136712,I1136514,I1136695);
nor I_66717 (I1136729,I1136627,I1136712);
DFFARX1 I_66718 (I1136729,I2507,I1136432,I1136400,);
DFFARX1 I_66719 (I1136712,I2507,I1136432,I1136421,);
nor I_66720 (I1136774,I177014,I177005);
nor I_66721 (I1136412,I1136627,I1136774);
or I_66722 (I1136805,I177014,I177005);
nor I_66723 (I1136822,I177020,I177026);
DFFARX1 I_66724 (I1136822,I2507,I1136432,I1136848,);
not I_66725 (I1136856,I1136848);
nor I_66726 (I1136418,I1136856,I1136661);
nand I_66727 (I1136887,I1136856,I1136506);
not I_66728 (I1136904,I177020);
nand I_66729 (I1136921,I1136904,I1136610);
nand I_66730 (I1136938,I1136856,I1136921);
nand I_66731 (I1136409,I1136938,I1136887);
nand I_66732 (I1136406,I1136921,I1136805);
not I_66733 (I1137010,I2514);
DFFARX1 I_66734 (I431087,I2507,I1137010,I1137036,);
and I_66735 (I1137044,I1137036,I431102);
DFFARX1 I_66736 (I1137044,I2507,I1137010,I1136993,);
DFFARX1 I_66737 (I431105,I2507,I1137010,I1137084,);
not I_66738 (I1137092,I431099);
not I_66739 (I1137109,I431114);
nand I_66740 (I1137126,I1137109,I1137092);
nor I_66741 (I1136981,I1137084,I1137126);
DFFARX1 I_66742 (I1137126,I2507,I1137010,I1137166,);
not I_66743 (I1137002,I1137166);
not I_66744 (I1137188,I431090);
nand I_66745 (I1137205,I1137109,I1137188);
DFFARX1 I_66746 (I1137205,I2507,I1137010,I1137231,);
not I_66747 (I1137239,I1137231);
not I_66748 (I1137256,I431093);
nand I_66749 (I1137273,I1137256,I431087);
and I_66750 (I1137290,I1137092,I1137273);
nor I_66751 (I1137307,I1137205,I1137290);
DFFARX1 I_66752 (I1137307,I2507,I1137010,I1136978,);
DFFARX1 I_66753 (I1137290,I2507,I1137010,I1136999,);
nor I_66754 (I1137352,I431093,I431096);
nor I_66755 (I1136990,I1137205,I1137352);
or I_66756 (I1137383,I431093,I431096);
nor I_66757 (I1137400,I431111,I431108);
DFFARX1 I_66758 (I1137400,I2507,I1137010,I1137426,);
not I_66759 (I1137434,I1137426);
nor I_66760 (I1136996,I1137434,I1137239);
nand I_66761 (I1137465,I1137434,I1137084);
not I_66762 (I1137482,I431111);
nand I_66763 (I1137499,I1137482,I1137188);
nand I_66764 (I1137516,I1137434,I1137499);
nand I_66765 (I1136987,I1137516,I1137465);
nand I_66766 (I1136984,I1137499,I1137383);
not I_66767 (I1137588,I2514);
DFFARX1 I_66768 (I1034828,I2507,I1137588,I1137614,);
and I_66769 (I1137622,I1137614,I1034825);
DFFARX1 I_66770 (I1137622,I2507,I1137588,I1137571,);
DFFARX1 I_66771 (I1034831,I2507,I1137588,I1137662,);
not I_66772 (I1137670,I1034834);
not I_66773 (I1137687,I1034828);
nand I_66774 (I1137704,I1137687,I1137670);
nor I_66775 (I1137559,I1137662,I1137704);
DFFARX1 I_66776 (I1137704,I2507,I1137588,I1137744,);
not I_66777 (I1137580,I1137744);
not I_66778 (I1137766,I1034843);
nand I_66779 (I1137783,I1137687,I1137766);
DFFARX1 I_66780 (I1137783,I2507,I1137588,I1137809,);
not I_66781 (I1137817,I1137809);
not I_66782 (I1137834,I1034840);
nand I_66783 (I1137851,I1137834,I1034846);
and I_66784 (I1137868,I1137670,I1137851);
nor I_66785 (I1137885,I1137783,I1137868);
DFFARX1 I_66786 (I1137885,I2507,I1137588,I1137556,);
DFFARX1 I_66787 (I1137868,I2507,I1137588,I1137577,);
nor I_66788 (I1137930,I1034840,I1034825);
nor I_66789 (I1137568,I1137783,I1137930);
or I_66790 (I1137961,I1034840,I1034825);
nor I_66791 (I1137978,I1034837,I1034831);
DFFARX1 I_66792 (I1137978,I2507,I1137588,I1138004,);
not I_66793 (I1138012,I1138004);
nor I_66794 (I1137574,I1138012,I1137817);
nand I_66795 (I1138043,I1138012,I1137662);
not I_66796 (I1138060,I1034837);
nand I_66797 (I1138077,I1138060,I1137766);
nand I_66798 (I1138094,I1138012,I1138077);
nand I_66799 (I1137565,I1138094,I1138043);
nand I_66800 (I1137562,I1138077,I1137961);
not I_66801 (I1138166,I2514);
DFFARX1 I_66802 (I154990,I2507,I1138166,I1138192,);
and I_66803 (I1138200,I1138192,I154993);
DFFARX1 I_66804 (I1138200,I2507,I1138166,I1138149,);
DFFARX1 I_66805 (I154993,I2507,I1138166,I1138240,);
not I_66806 (I1138248,I155008);
not I_66807 (I1138265,I155014);
nand I_66808 (I1138282,I1138265,I1138248);
nor I_66809 (I1138137,I1138240,I1138282);
DFFARX1 I_66810 (I1138282,I2507,I1138166,I1138322,);
not I_66811 (I1138158,I1138322);
not I_66812 (I1138344,I155002);
nand I_66813 (I1138361,I1138265,I1138344);
DFFARX1 I_66814 (I1138361,I2507,I1138166,I1138387,);
not I_66815 (I1138395,I1138387);
not I_66816 (I1138412,I154999);
nand I_66817 (I1138429,I1138412,I154996);
and I_66818 (I1138446,I1138248,I1138429);
nor I_66819 (I1138463,I1138361,I1138446);
DFFARX1 I_66820 (I1138463,I2507,I1138166,I1138134,);
DFFARX1 I_66821 (I1138446,I2507,I1138166,I1138155,);
nor I_66822 (I1138508,I154999,I154990);
nor I_66823 (I1138146,I1138361,I1138508);
or I_66824 (I1138539,I154999,I154990);
nor I_66825 (I1138556,I155005,I155011);
DFFARX1 I_66826 (I1138556,I2507,I1138166,I1138582,);
not I_66827 (I1138590,I1138582);
nor I_66828 (I1138152,I1138590,I1138395);
nand I_66829 (I1138621,I1138590,I1138240);
not I_66830 (I1138638,I155005);
nand I_66831 (I1138655,I1138638,I1138344);
nand I_66832 (I1138672,I1138590,I1138655);
nand I_66833 (I1138143,I1138672,I1138621);
nand I_66834 (I1138140,I1138655,I1138539);
not I_66835 (I1138744,I2514);
DFFARX1 I_66836 (I51722,I2507,I1138744,I1138770,);
and I_66837 (I1138778,I1138770,I51698);
DFFARX1 I_66838 (I1138778,I2507,I1138744,I1138727,);
DFFARX1 I_66839 (I51716,I2507,I1138744,I1138818,);
not I_66840 (I1138826,I51704);
not I_66841 (I1138843,I51701);
nand I_66842 (I1138860,I1138843,I1138826);
nor I_66843 (I1138715,I1138818,I1138860);
DFFARX1 I_66844 (I1138860,I2507,I1138744,I1138900,);
not I_66845 (I1138736,I1138900);
not I_66846 (I1138922,I51710);
nand I_66847 (I1138939,I1138843,I1138922);
DFFARX1 I_66848 (I1138939,I2507,I1138744,I1138965,);
not I_66849 (I1138973,I1138965);
not I_66850 (I1138990,I51701);
nand I_66851 (I1139007,I1138990,I51719);
and I_66852 (I1139024,I1138826,I1139007);
nor I_66853 (I1139041,I1138939,I1139024);
DFFARX1 I_66854 (I1139041,I2507,I1138744,I1138712,);
DFFARX1 I_66855 (I1139024,I2507,I1138744,I1138733,);
nor I_66856 (I1139086,I51701,I51713);
nor I_66857 (I1138724,I1138939,I1139086);
or I_66858 (I1139117,I51701,I51713);
nor I_66859 (I1139134,I51707,I51698);
DFFARX1 I_66860 (I1139134,I2507,I1138744,I1139160,);
not I_66861 (I1139168,I1139160);
nor I_66862 (I1138730,I1139168,I1138973);
nand I_66863 (I1139199,I1139168,I1138818);
not I_66864 (I1139216,I51707);
nand I_66865 (I1139233,I1139216,I1138922);
nand I_66866 (I1139250,I1139168,I1139233);
nand I_66867 (I1138721,I1139250,I1139199);
nand I_66868 (I1138718,I1139233,I1139117);
not I_66869 (I1139322,I2514);
DFFARX1 I_66870 (I185335,I2507,I1139322,I1139348,);
and I_66871 (I1139356,I1139348,I185338);
DFFARX1 I_66872 (I1139356,I2507,I1139322,I1139305,);
DFFARX1 I_66873 (I185338,I2507,I1139322,I1139396,);
not I_66874 (I1139404,I185353);
not I_66875 (I1139421,I185359);
nand I_66876 (I1139438,I1139421,I1139404);
nor I_66877 (I1139293,I1139396,I1139438);
DFFARX1 I_66878 (I1139438,I2507,I1139322,I1139478,);
not I_66879 (I1139314,I1139478);
not I_66880 (I1139500,I185347);
nand I_66881 (I1139517,I1139421,I1139500);
DFFARX1 I_66882 (I1139517,I2507,I1139322,I1139543,);
not I_66883 (I1139551,I1139543);
not I_66884 (I1139568,I185344);
nand I_66885 (I1139585,I1139568,I185341);
and I_66886 (I1139602,I1139404,I1139585);
nor I_66887 (I1139619,I1139517,I1139602);
DFFARX1 I_66888 (I1139619,I2507,I1139322,I1139290,);
DFFARX1 I_66889 (I1139602,I2507,I1139322,I1139311,);
nor I_66890 (I1139664,I185344,I185335);
nor I_66891 (I1139302,I1139517,I1139664);
or I_66892 (I1139695,I185344,I185335);
nor I_66893 (I1139712,I185350,I185356);
DFFARX1 I_66894 (I1139712,I2507,I1139322,I1139738,);
not I_66895 (I1139746,I1139738);
nor I_66896 (I1139308,I1139746,I1139551);
nand I_66897 (I1139777,I1139746,I1139396);
not I_66898 (I1139794,I185350);
nand I_66899 (I1139811,I1139794,I1139500);
nand I_66900 (I1139828,I1139746,I1139811);
nand I_66901 (I1139299,I1139828,I1139777);
nand I_66902 (I1139296,I1139811,I1139695);
not I_66903 (I1139900,I2514);
DFFARX1 I_66904 (I785914,I2507,I1139900,I1139926,);
and I_66905 (I1139934,I1139926,I785920);
DFFARX1 I_66906 (I1139934,I2507,I1139900,I1139883,);
DFFARX1 I_66907 (I785926,I2507,I1139900,I1139974,);
not I_66908 (I1139982,I785911);
not I_66909 (I1139999,I785911);
nand I_66910 (I1140016,I1139999,I1139982);
nor I_66911 (I1139871,I1139974,I1140016);
DFFARX1 I_66912 (I1140016,I2507,I1139900,I1140056,);
not I_66913 (I1139892,I1140056);
not I_66914 (I1140078,I785929);
nand I_66915 (I1140095,I1139999,I1140078);
DFFARX1 I_66916 (I1140095,I2507,I1139900,I1140121,);
not I_66917 (I1140129,I1140121);
not I_66918 (I1140146,I785923);
nand I_66919 (I1140163,I1140146,I785914);
and I_66920 (I1140180,I1139982,I1140163);
nor I_66921 (I1140197,I1140095,I1140180);
DFFARX1 I_66922 (I1140197,I2507,I1139900,I1139868,);
DFFARX1 I_66923 (I1140180,I2507,I1139900,I1139889,);
nor I_66924 (I1140242,I785923,I785932);
nor I_66925 (I1139880,I1140095,I1140242);
or I_66926 (I1140273,I785923,I785932);
nor I_66927 (I1140290,I785917,I785917);
DFFARX1 I_66928 (I1140290,I2507,I1139900,I1140316,);
not I_66929 (I1140324,I1140316);
nor I_66930 (I1139886,I1140324,I1140129);
nand I_66931 (I1140355,I1140324,I1139974);
not I_66932 (I1140372,I785917);
nand I_66933 (I1140389,I1140372,I1140078);
nand I_66934 (I1140406,I1140324,I1140389);
nand I_66935 (I1139877,I1140406,I1140355);
nand I_66936 (I1139874,I1140389,I1140273);
not I_66937 (I1140478,I2514);
DFFARX1 I_66938 (I129191,I2507,I1140478,I1140504,);
and I_66939 (I1140512,I1140504,I129167);
DFFARX1 I_66940 (I1140512,I2507,I1140478,I1140461,);
DFFARX1 I_66941 (I129185,I2507,I1140478,I1140552,);
not I_66942 (I1140560,I129173);
not I_66943 (I1140577,I129170);
nand I_66944 (I1140594,I1140577,I1140560);
nor I_66945 (I1140449,I1140552,I1140594);
DFFARX1 I_66946 (I1140594,I2507,I1140478,I1140634,);
not I_66947 (I1140470,I1140634);
not I_66948 (I1140656,I129179);
nand I_66949 (I1140673,I1140577,I1140656);
DFFARX1 I_66950 (I1140673,I2507,I1140478,I1140699,);
not I_66951 (I1140707,I1140699);
not I_66952 (I1140724,I129170);
nand I_66953 (I1140741,I1140724,I129188);
and I_66954 (I1140758,I1140560,I1140741);
nor I_66955 (I1140775,I1140673,I1140758);
DFFARX1 I_66956 (I1140775,I2507,I1140478,I1140446,);
DFFARX1 I_66957 (I1140758,I2507,I1140478,I1140467,);
nor I_66958 (I1140820,I129170,I129182);
nor I_66959 (I1140458,I1140673,I1140820);
or I_66960 (I1140851,I129170,I129182);
nor I_66961 (I1140868,I129176,I129167);
DFFARX1 I_66962 (I1140868,I2507,I1140478,I1140894,);
not I_66963 (I1140902,I1140894);
nor I_66964 (I1140464,I1140902,I1140707);
nand I_66965 (I1140933,I1140902,I1140552);
not I_66966 (I1140950,I129176);
nand I_66967 (I1140967,I1140950,I1140656);
nand I_66968 (I1140984,I1140902,I1140967);
nand I_66969 (I1140455,I1140984,I1140933);
nand I_66970 (I1140452,I1140967,I1140851);
not I_66971 (I1141056,I2514);
DFFARX1 I_66972 (I401167,I2507,I1141056,I1141082,);
and I_66973 (I1141090,I1141082,I401182);
DFFARX1 I_66974 (I1141090,I2507,I1141056,I1141039,);
DFFARX1 I_66975 (I401185,I2507,I1141056,I1141130,);
not I_66976 (I1141138,I401179);
not I_66977 (I1141155,I401194);
nand I_66978 (I1141172,I1141155,I1141138);
nor I_66979 (I1141027,I1141130,I1141172);
DFFARX1 I_66980 (I1141172,I2507,I1141056,I1141212,);
not I_66981 (I1141048,I1141212);
not I_66982 (I1141234,I401170);
nand I_66983 (I1141251,I1141155,I1141234);
DFFARX1 I_66984 (I1141251,I2507,I1141056,I1141277,);
not I_66985 (I1141285,I1141277);
not I_66986 (I1141302,I401173);
nand I_66987 (I1141319,I1141302,I401167);
and I_66988 (I1141336,I1141138,I1141319);
nor I_66989 (I1141353,I1141251,I1141336);
DFFARX1 I_66990 (I1141353,I2507,I1141056,I1141024,);
DFFARX1 I_66991 (I1141336,I2507,I1141056,I1141045,);
nor I_66992 (I1141398,I401173,I401176);
nor I_66993 (I1141036,I1141251,I1141398);
or I_66994 (I1141429,I401173,I401176);
nor I_66995 (I1141446,I401191,I401188);
DFFARX1 I_66996 (I1141446,I2507,I1141056,I1141472,);
not I_66997 (I1141480,I1141472);
nor I_66998 (I1141042,I1141480,I1141285);
nand I_66999 (I1141511,I1141480,I1141130);
not I_67000 (I1141528,I401191);
nand I_67001 (I1141545,I1141528,I1141234);
nand I_67002 (I1141562,I1141480,I1141545);
nand I_67003 (I1141033,I1141562,I1141511);
nand I_67004 (I1141030,I1141545,I1141429);
not I_67005 (I1141634,I2514);
DFFARX1 I_67006 (I763095,I2507,I1141634,I1141660,);
and I_67007 (I1141668,I1141660,I763083);
DFFARX1 I_67008 (I1141668,I2507,I1141634,I1141617,);
DFFARX1 I_67009 (I763086,I2507,I1141634,I1141708,);
not I_67010 (I1141716,I763080);
not I_67011 (I1141733,I763104);
nand I_67012 (I1141750,I1141733,I1141716);
nor I_67013 (I1141605,I1141708,I1141750);
DFFARX1 I_67014 (I1141750,I2507,I1141634,I1141790,);
not I_67015 (I1141626,I1141790);
not I_67016 (I1141812,I763092);
nand I_67017 (I1141829,I1141733,I1141812);
DFFARX1 I_67018 (I1141829,I2507,I1141634,I1141855,);
not I_67019 (I1141863,I1141855);
not I_67020 (I1141880,I763101);
nand I_67021 (I1141897,I1141880,I763098);
and I_67022 (I1141914,I1141716,I1141897);
nor I_67023 (I1141931,I1141829,I1141914);
DFFARX1 I_67024 (I1141931,I2507,I1141634,I1141602,);
DFFARX1 I_67025 (I1141914,I2507,I1141634,I1141623,);
nor I_67026 (I1141976,I763101,I763089);
nor I_67027 (I1141614,I1141829,I1141976);
or I_67028 (I1142007,I763101,I763089);
nor I_67029 (I1142024,I763080,I763083);
DFFARX1 I_67030 (I1142024,I2507,I1141634,I1142050,);
not I_67031 (I1142058,I1142050);
nor I_67032 (I1141620,I1142058,I1141863);
nand I_67033 (I1142089,I1142058,I1141708);
not I_67034 (I1142106,I763080);
nand I_67035 (I1142123,I1142106,I1141812);
nand I_67036 (I1142140,I1142058,I1142123);
nand I_67037 (I1141611,I1142140,I1142089);
nand I_67038 (I1141608,I1142123,I1142007);
not I_67039 (I1142212,I2514);
DFFARX1 I_67040 (I156775,I2507,I1142212,I1142238,);
and I_67041 (I1142246,I1142238,I156778);
DFFARX1 I_67042 (I1142246,I2507,I1142212,I1142195,);
DFFARX1 I_67043 (I156778,I2507,I1142212,I1142286,);
not I_67044 (I1142294,I156793);
not I_67045 (I1142311,I156799);
nand I_67046 (I1142328,I1142311,I1142294);
nor I_67047 (I1142183,I1142286,I1142328);
DFFARX1 I_67048 (I1142328,I2507,I1142212,I1142368,);
not I_67049 (I1142204,I1142368);
not I_67050 (I1142390,I156787);
nand I_67051 (I1142407,I1142311,I1142390);
DFFARX1 I_67052 (I1142407,I2507,I1142212,I1142433,);
not I_67053 (I1142441,I1142433);
not I_67054 (I1142458,I156784);
nand I_67055 (I1142475,I1142458,I156781);
and I_67056 (I1142492,I1142294,I1142475);
nor I_67057 (I1142509,I1142407,I1142492);
DFFARX1 I_67058 (I1142509,I2507,I1142212,I1142180,);
DFFARX1 I_67059 (I1142492,I2507,I1142212,I1142201,);
nor I_67060 (I1142554,I156784,I156775);
nor I_67061 (I1142192,I1142407,I1142554);
or I_67062 (I1142585,I156784,I156775);
nor I_67063 (I1142602,I156790,I156796);
DFFARX1 I_67064 (I1142602,I2507,I1142212,I1142628,);
not I_67065 (I1142636,I1142628);
nor I_67066 (I1142198,I1142636,I1142441);
nand I_67067 (I1142667,I1142636,I1142286);
not I_67068 (I1142684,I156790);
nand I_67069 (I1142701,I1142684,I1142390);
nand I_67070 (I1142718,I1142636,I1142701);
nand I_67071 (I1142189,I1142718,I1142667);
nand I_67072 (I1142186,I1142701,I1142585);
not I_67073 (I1142790,I2514);
DFFARX1 I_67074 (I608191,I2507,I1142790,I1142816,);
and I_67075 (I1142824,I1142816,I608179);
DFFARX1 I_67076 (I1142824,I2507,I1142790,I1142773,);
DFFARX1 I_67077 (I608194,I2507,I1142790,I1142864,);
not I_67078 (I1142872,I608185);
not I_67079 (I1142889,I608176);
nand I_67080 (I1142906,I1142889,I1142872);
nor I_67081 (I1142761,I1142864,I1142906);
DFFARX1 I_67082 (I1142906,I2507,I1142790,I1142946,);
not I_67083 (I1142782,I1142946);
not I_67084 (I1142968,I608182);
nand I_67085 (I1142985,I1142889,I1142968);
DFFARX1 I_67086 (I1142985,I2507,I1142790,I1143011,);
not I_67087 (I1143019,I1143011);
not I_67088 (I1143036,I608197);
nand I_67089 (I1143053,I1143036,I608200);
and I_67090 (I1143070,I1142872,I1143053);
nor I_67091 (I1143087,I1142985,I1143070);
DFFARX1 I_67092 (I1143087,I2507,I1142790,I1142758,);
DFFARX1 I_67093 (I1143070,I2507,I1142790,I1142779,);
nor I_67094 (I1143132,I608197,I608176);
nor I_67095 (I1142770,I1142985,I1143132);
or I_67096 (I1143163,I608197,I608176);
nor I_67097 (I1143180,I608188,I608179);
DFFARX1 I_67098 (I1143180,I2507,I1142790,I1143206,);
not I_67099 (I1143214,I1143206);
nor I_67100 (I1142776,I1143214,I1143019);
nand I_67101 (I1143245,I1143214,I1142864);
not I_67102 (I1143262,I608188);
nand I_67103 (I1143279,I1143262,I1142968);
nand I_67104 (I1143296,I1143214,I1143279);
nand I_67105 (I1142767,I1143296,I1143245);
nand I_67106 (I1142764,I1143279,I1143163);
not I_67107 (I1143368,I2514);
DFFARX1 I_67108 (I126029,I2507,I1143368,I1143394,);
and I_67109 (I1143402,I1143394,I126005);
DFFARX1 I_67110 (I1143402,I2507,I1143368,I1143351,);
DFFARX1 I_67111 (I126023,I2507,I1143368,I1143442,);
not I_67112 (I1143450,I126011);
not I_67113 (I1143467,I126008);
nand I_67114 (I1143484,I1143467,I1143450);
nor I_67115 (I1143339,I1143442,I1143484);
DFFARX1 I_67116 (I1143484,I2507,I1143368,I1143524,);
not I_67117 (I1143360,I1143524);
not I_67118 (I1143546,I126017);
nand I_67119 (I1143563,I1143467,I1143546);
DFFARX1 I_67120 (I1143563,I2507,I1143368,I1143589,);
not I_67121 (I1143597,I1143589);
not I_67122 (I1143614,I126008);
nand I_67123 (I1143631,I1143614,I126026);
and I_67124 (I1143648,I1143450,I1143631);
nor I_67125 (I1143665,I1143563,I1143648);
DFFARX1 I_67126 (I1143665,I2507,I1143368,I1143336,);
DFFARX1 I_67127 (I1143648,I2507,I1143368,I1143357,);
nor I_67128 (I1143710,I126008,I126020);
nor I_67129 (I1143348,I1143563,I1143710);
or I_67130 (I1143741,I126008,I126020);
nor I_67131 (I1143758,I126014,I126005);
DFFARX1 I_67132 (I1143758,I2507,I1143368,I1143784,);
not I_67133 (I1143792,I1143784);
nor I_67134 (I1143354,I1143792,I1143597);
nand I_67135 (I1143823,I1143792,I1143442);
not I_67136 (I1143840,I126014);
nand I_67137 (I1143857,I1143840,I1143546);
nand I_67138 (I1143874,I1143792,I1143857);
nand I_67139 (I1143345,I1143874,I1143823);
nand I_67140 (I1143342,I1143857,I1143741);
not I_67141 (I1143946,I2514);
DFFARX1 I_67142 (I70694,I2507,I1143946,I1143972,);
and I_67143 (I1143980,I1143972,I70670);
DFFARX1 I_67144 (I1143980,I2507,I1143946,I1143929,);
DFFARX1 I_67145 (I70688,I2507,I1143946,I1144020,);
not I_67146 (I1144028,I70676);
not I_67147 (I1144045,I70673);
nand I_67148 (I1144062,I1144045,I1144028);
nor I_67149 (I1143917,I1144020,I1144062);
DFFARX1 I_67150 (I1144062,I2507,I1143946,I1144102,);
not I_67151 (I1143938,I1144102);
not I_67152 (I1144124,I70682);
nand I_67153 (I1144141,I1144045,I1144124);
DFFARX1 I_67154 (I1144141,I2507,I1143946,I1144167,);
not I_67155 (I1144175,I1144167);
not I_67156 (I1144192,I70673);
nand I_67157 (I1144209,I1144192,I70691);
and I_67158 (I1144226,I1144028,I1144209);
nor I_67159 (I1144243,I1144141,I1144226);
DFFARX1 I_67160 (I1144243,I2507,I1143946,I1143914,);
DFFARX1 I_67161 (I1144226,I2507,I1143946,I1143935,);
nor I_67162 (I1144288,I70673,I70685);
nor I_67163 (I1143926,I1144141,I1144288);
or I_67164 (I1144319,I70673,I70685);
nor I_67165 (I1144336,I70679,I70670);
DFFARX1 I_67166 (I1144336,I2507,I1143946,I1144362,);
not I_67167 (I1144370,I1144362);
nor I_67168 (I1143932,I1144370,I1144175);
nand I_67169 (I1144401,I1144370,I1144020);
not I_67170 (I1144418,I70679);
nand I_67171 (I1144435,I1144418,I1144124);
nand I_67172 (I1144452,I1144370,I1144435);
nand I_67173 (I1143923,I1144452,I1144401);
nand I_67174 (I1143920,I1144435,I1144319);
not I_67175 (I1144524,I2514);
DFFARX1 I_67176 (I270243,I2507,I1144524,I1144550,);
and I_67177 (I1144558,I1144550,I270228);
DFFARX1 I_67178 (I1144558,I2507,I1144524,I1144507,);
DFFARX1 I_67179 (I270234,I2507,I1144524,I1144598,);
not I_67180 (I1144606,I270216);
not I_67181 (I1144623,I270237);
nand I_67182 (I1144640,I1144623,I1144606);
nor I_67183 (I1144495,I1144598,I1144640);
DFFARX1 I_67184 (I1144640,I2507,I1144524,I1144680,);
not I_67185 (I1144516,I1144680);
not I_67186 (I1144702,I270240);
nand I_67187 (I1144719,I1144623,I1144702);
DFFARX1 I_67188 (I1144719,I2507,I1144524,I1144745,);
not I_67189 (I1144753,I1144745);
not I_67190 (I1144770,I270231);
nand I_67191 (I1144787,I1144770,I270219);
and I_67192 (I1144804,I1144606,I1144787);
nor I_67193 (I1144821,I1144719,I1144804);
DFFARX1 I_67194 (I1144821,I2507,I1144524,I1144492,);
DFFARX1 I_67195 (I1144804,I2507,I1144524,I1144513,);
nor I_67196 (I1144866,I270231,I270225);
nor I_67197 (I1144504,I1144719,I1144866);
or I_67198 (I1144897,I270231,I270225);
nor I_67199 (I1144914,I270222,I270216);
DFFARX1 I_67200 (I1144914,I2507,I1144524,I1144940,);
not I_67201 (I1144948,I1144940);
nor I_67202 (I1144510,I1144948,I1144753);
nand I_67203 (I1144979,I1144948,I1144598);
not I_67204 (I1144996,I270222);
nand I_67205 (I1145013,I1144996,I1144702);
nand I_67206 (I1145030,I1144948,I1145013);
nand I_67207 (I1144501,I1145030,I1144979);
nand I_67208 (I1144498,I1145013,I1144897);
not I_67209 (I1145102,I2514);
DFFARX1 I_67210 (I1224311,I2507,I1145102,I1145128,);
and I_67211 (I1145136,I1145128,I1224305);
DFFARX1 I_67212 (I1145136,I2507,I1145102,I1145085,);
DFFARX1 I_67213 (I1224290,I2507,I1145102,I1145176,);
not I_67214 (I1145184,I1224296);
not I_67215 (I1145201,I1224308);
nand I_67216 (I1145218,I1145201,I1145184);
nor I_67217 (I1145073,I1145176,I1145218);
DFFARX1 I_67218 (I1145218,I2507,I1145102,I1145258,);
not I_67219 (I1145094,I1145258);
not I_67220 (I1145280,I1224290);
nand I_67221 (I1145297,I1145201,I1145280);
DFFARX1 I_67222 (I1145297,I2507,I1145102,I1145323,);
not I_67223 (I1145331,I1145323);
not I_67224 (I1145348,I1224314);
nand I_67225 (I1145365,I1145348,I1224302);
and I_67226 (I1145382,I1145184,I1145365);
nor I_67227 (I1145399,I1145297,I1145382);
DFFARX1 I_67228 (I1145399,I2507,I1145102,I1145070,);
DFFARX1 I_67229 (I1145382,I2507,I1145102,I1145091,);
nor I_67230 (I1145444,I1224314,I1224293);
nor I_67231 (I1145082,I1145297,I1145444);
or I_67232 (I1145475,I1224314,I1224293);
nor I_67233 (I1145492,I1224299,I1224293);
DFFARX1 I_67234 (I1145492,I2507,I1145102,I1145518,);
not I_67235 (I1145526,I1145518);
nor I_67236 (I1145088,I1145526,I1145331);
nand I_67237 (I1145557,I1145526,I1145176);
not I_67238 (I1145574,I1224299);
nand I_67239 (I1145591,I1145574,I1145280);
nand I_67240 (I1145608,I1145526,I1145591);
nand I_67241 (I1145079,I1145608,I1145557);
nand I_67242 (I1145076,I1145591,I1145475);
not I_67243 (I1145680,I2514);
DFFARX1 I_67244 (I770031,I2507,I1145680,I1145706,);
and I_67245 (I1145714,I1145706,I770019);
DFFARX1 I_67246 (I1145714,I2507,I1145680,I1145663,);
DFFARX1 I_67247 (I770022,I2507,I1145680,I1145754,);
not I_67248 (I1145762,I770016);
not I_67249 (I1145779,I770040);
nand I_67250 (I1145796,I1145779,I1145762);
nor I_67251 (I1145651,I1145754,I1145796);
DFFARX1 I_67252 (I1145796,I2507,I1145680,I1145836,);
not I_67253 (I1145672,I1145836);
not I_67254 (I1145858,I770028);
nand I_67255 (I1145875,I1145779,I1145858);
DFFARX1 I_67256 (I1145875,I2507,I1145680,I1145901,);
not I_67257 (I1145909,I1145901);
not I_67258 (I1145926,I770037);
nand I_67259 (I1145943,I1145926,I770034);
and I_67260 (I1145960,I1145762,I1145943);
nor I_67261 (I1145977,I1145875,I1145960);
DFFARX1 I_67262 (I1145977,I2507,I1145680,I1145648,);
DFFARX1 I_67263 (I1145960,I2507,I1145680,I1145669,);
nor I_67264 (I1146022,I770037,I770025);
nor I_67265 (I1145660,I1145875,I1146022);
or I_67266 (I1146053,I770037,I770025);
nor I_67267 (I1146070,I770016,I770019);
DFFARX1 I_67268 (I1146070,I2507,I1145680,I1146096,);
not I_67269 (I1146104,I1146096);
nor I_67270 (I1145666,I1146104,I1145909);
nand I_67271 (I1146135,I1146104,I1145754);
not I_67272 (I1146152,I770016);
nand I_67273 (I1146169,I1146152,I1145858);
nand I_67274 (I1146186,I1146104,I1146169);
nand I_67275 (I1145657,I1146186,I1146135);
nand I_67276 (I1145654,I1146169,I1146053);
not I_67277 (I1146258,I2514);
DFFARX1 I_67278 (I345604,I2507,I1146258,I1146284,);
and I_67279 (I1146292,I1146284,I345589);
DFFARX1 I_67280 (I1146292,I2507,I1146258,I1146241,);
DFFARX1 I_67281 (I345595,I2507,I1146258,I1146332,);
not I_67282 (I1146340,I345577);
not I_67283 (I1146357,I345598);
nand I_67284 (I1146374,I1146357,I1146340);
nor I_67285 (I1146229,I1146332,I1146374);
DFFARX1 I_67286 (I1146374,I2507,I1146258,I1146414,);
not I_67287 (I1146250,I1146414);
not I_67288 (I1146436,I345601);
nand I_67289 (I1146453,I1146357,I1146436);
DFFARX1 I_67290 (I1146453,I2507,I1146258,I1146479,);
not I_67291 (I1146487,I1146479);
not I_67292 (I1146504,I345592);
nand I_67293 (I1146521,I1146504,I345580);
and I_67294 (I1146538,I1146340,I1146521);
nor I_67295 (I1146555,I1146453,I1146538);
DFFARX1 I_67296 (I1146555,I2507,I1146258,I1146226,);
DFFARX1 I_67297 (I1146538,I2507,I1146258,I1146247,);
nor I_67298 (I1146600,I345592,I345586);
nor I_67299 (I1146238,I1146453,I1146600);
or I_67300 (I1146631,I345592,I345586);
nor I_67301 (I1146648,I345583,I345577);
DFFARX1 I_67302 (I1146648,I2507,I1146258,I1146674,);
not I_67303 (I1146682,I1146674);
nor I_67304 (I1146244,I1146682,I1146487);
nand I_67305 (I1146713,I1146682,I1146332);
not I_67306 (I1146730,I345583);
nand I_67307 (I1146747,I1146730,I1146436);
nand I_67308 (I1146764,I1146682,I1146747);
nand I_67309 (I1146235,I1146764,I1146713);
nand I_67310 (I1146232,I1146747,I1146631);
not I_67311 (I1146836,I2514);
DFFARX1 I_67312 (I153205,I2507,I1146836,I1146862,);
and I_67313 (I1146870,I1146862,I153208);
DFFARX1 I_67314 (I1146870,I2507,I1146836,I1146819,);
DFFARX1 I_67315 (I153208,I2507,I1146836,I1146910,);
not I_67316 (I1146918,I153223);
not I_67317 (I1146935,I153229);
nand I_67318 (I1146952,I1146935,I1146918);
nor I_67319 (I1146807,I1146910,I1146952);
DFFARX1 I_67320 (I1146952,I2507,I1146836,I1146992,);
not I_67321 (I1146828,I1146992);
not I_67322 (I1147014,I153217);
nand I_67323 (I1147031,I1146935,I1147014);
DFFARX1 I_67324 (I1147031,I2507,I1146836,I1147057,);
not I_67325 (I1147065,I1147057);
not I_67326 (I1147082,I153214);
nand I_67327 (I1147099,I1147082,I153211);
and I_67328 (I1147116,I1146918,I1147099);
nor I_67329 (I1147133,I1147031,I1147116);
DFFARX1 I_67330 (I1147133,I2507,I1146836,I1146804,);
DFFARX1 I_67331 (I1147116,I2507,I1146836,I1146825,);
nor I_67332 (I1147178,I153214,I153205);
nor I_67333 (I1146816,I1147031,I1147178);
or I_67334 (I1147209,I153214,I153205);
nor I_67335 (I1147226,I153220,I153226);
DFFARX1 I_67336 (I1147226,I2507,I1146836,I1147252,);
not I_67337 (I1147260,I1147252);
nor I_67338 (I1146822,I1147260,I1147065);
nand I_67339 (I1147291,I1147260,I1146910);
not I_67340 (I1147308,I153220);
nand I_67341 (I1147325,I1147308,I1147014);
nand I_67342 (I1147342,I1147260,I1147325);
nand I_67343 (I1146813,I1147342,I1147291);
nand I_67344 (I1146810,I1147325,I1147209);
not I_67345 (I1147414,I2514);
DFFARX1 I_67346 (I748067,I2507,I1147414,I1147440,);
and I_67347 (I1147448,I1147440,I748055);
DFFARX1 I_67348 (I1147448,I2507,I1147414,I1147397,);
DFFARX1 I_67349 (I748058,I2507,I1147414,I1147488,);
not I_67350 (I1147496,I748052);
not I_67351 (I1147513,I748076);
nand I_67352 (I1147530,I1147513,I1147496);
nor I_67353 (I1147385,I1147488,I1147530);
DFFARX1 I_67354 (I1147530,I2507,I1147414,I1147570,);
not I_67355 (I1147406,I1147570);
not I_67356 (I1147592,I748064);
nand I_67357 (I1147609,I1147513,I1147592);
DFFARX1 I_67358 (I1147609,I2507,I1147414,I1147635,);
not I_67359 (I1147643,I1147635);
not I_67360 (I1147660,I748073);
nand I_67361 (I1147677,I1147660,I748070);
and I_67362 (I1147694,I1147496,I1147677);
nor I_67363 (I1147711,I1147609,I1147694);
DFFARX1 I_67364 (I1147711,I2507,I1147414,I1147382,);
DFFARX1 I_67365 (I1147694,I2507,I1147414,I1147403,);
nor I_67366 (I1147756,I748073,I748061);
nor I_67367 (I1147394,I1147609,I1147756);
or I_67368 (I1147787,I748073,I748061);
nor I_67369 (I1147804,I748052,I748055);
DFFARX1 I_67370 (I1147804,I2507,I1147414,I1147830,);
not I_67371 (I1147838,I1147830);
nor I_67372 (I1147400,I1147838,I1147643);
nand I_67373 (I1147869,I1147838,I1147488);
not I_67374 (I1147886,I748052);
nand I_67375 (I1147903,I1147886,I1147592);
nand I_67376 (I1147920,I1147838,I1147903);
nand I_67377 (I1147391,I1147920,I1147869);
nand I_67378 (I1147388,I1147903,I1147787);
not I_67379 (I1147992,I2514);
DFFARX1 I_67380 (I1046609,I2507,I1147992,I1148018,);
and I_67381 (I1148026,I1148018,I1046606);
DFFARX1 I_67382 (I1148026,I2507,I1147992,I1147975,);
DFFARX1 I_67383 (I1046612,I2507,I1147992,I1148066,);
not I_67384 (I1148074,I1046615);
not I_67385 (I1148091,I1046609);
nand I_67386 (I1148108,I1148091,I1148074);
nor I_67387 (I1147963,I1148066,I1148108);
DFFARX1 I_67388 (I1148108,I2507,I1147992,I1148148,);
not I_67389 (I1147984,I1148148);
not I_67390 (I1148170,I1046624);
nand I_67391 (I1148187,I1148091,I1148170);
DFFARX1 I_67392 (I1148187,I2507,I1147992,I1148213,);
not I_67393 (I1148221,I1148213);
not I_67394 (I1148238,I1046621);
nand I_67395 (I1148255,I1148238,I1046627);
and I_67396 (I1148272,I1148074,I1148255);
nor I_67397 (I1148289,I1148187,I1148272);
DFFARX1 I_67398 (I1148289,I2507,I1147992,I1147960,);
DFFARX1 I_67399 (I1148272,I2507,I1147992,I1147981,);
nor I_67400 (I1148334,I1046621,I1046606);
nor I_67401 (I1147972,I1148187,I1148334);
or I_67402 (I1148365,I1046621,I1046606);
nor I_67403 (I1148382,I1046618,I1046612);
DFFARX1 I_67404 (I1148382,I2507,I1147992,I1148408,);
not I_67405 (I1148416,I1148408);
nor I_67406 (I1147978,I1148416,I1148221);
nand I_67407 (I1148447,I1148416,I1148066);
not I_67408 (I1148464,I1046618);
nand I_67409 (I1148481,I1148464,I1148170);
nand I_67410 (I1148498,I1148416,I1148481);
nand I_67411 (I1147969,I1148498,I1148447);
nand I_67412 (I1147966,I1148481,I1148365);
not I_67413 (I1148570,I2514);
DFFARX1 I_67414 (I174625,I2507,I1148570,I1148596,);
and I_67415 (I1148604,I1148596,I174628);
DFFARX1 I_67416 (I1148604,I2507,I1148570,I1148553,);
DFFARX1 I_67417 (I174628,I2507,I1148570,I1148644,);
not I_67418 (I1148652,I174643);
not I_67419 (I1148669,I174649);
nand I_67420 (I1148686,I1148669,I1148652);
nor I_67421 (I1148541,I1148644,I1148686);
DFFARX1 I_67422 (I1148686,I2507,I1148570,I1148726,);
not I_67423 (I1148562,I1148726);
not I_67424 (I1148748,I174637);
nand I_67425 (I1148765,I1148669,I1148748);
DFFARX1 I_67426 (I1148765,I2507,I1148570,I1148791,);
not I_67427 (I1148799,I1148791);
not I_67428 (I1148816,I174634);
nand I_67429 (I1148833,I1148816,I174631);
and I_67430 (I1148850,I1148652,I1148833);
nor I_67431 (I1148867,I1148765,I1148850);
DFFARX1 I_67432 (I1148867,I2507,I1148570,I1148538,);
DFFARX1 I_67433 (I1148850,I2507,I1148570,I1148559,);
nor I_67434 (I1148912,I174634,I174625);
nor I_67435 (I1148550,I1148765,I1148912);
or I_67436 (I1148943,I174634,I174625);
nor I_67437 (I1148960,I174640,I174646);
DFFARX1 I_67438 (I1148960,I2507,I1148570,I1148986,);
not I_67439 (I1148994,I1148986);
nor I_67440 (I1148556,I1148994,I1148799);
nand I_67441 (I1149025,I1148994,I1148644);
not I_67442 (I1149042,I174640);
nand I_67443 (I1149059,I1149042,I1148748);
nand I_67444 (I1149076,I1148994,I1149059);
nand I_67445 (I1148547,I1149076,I1149025);
nand I_67446 (I1148544,I1149059,I1148943);
not I_67447 (I1149148,I2514);
DFFARX1 I_67448 (I544611,I2507,I1149148,I1149174,);
and I_67449 (I1149182,I1149174,I544599);
DFFARX1 I_67450 (I1149182,I2507,I1149148,I1149131,);
DFFARX1 I_67451 (I544614,I2507,I1149148,I1149222,);
not I_67452 (I1149230,I544605);
not I_67453 (I1149247,I544596);
nand I_67454 (I1149264,I1149247,I1149230);
nor I_67455 (I1149119,I1149222,I1149264);
DFFARX1 I_67456 (I1149264,I2507,I1149148,I1149304,);
not I_67457 (I1149140,I1149304);
not I_67458 (I1149326,I544602);
nand I_67459 (I1149343,I1149247,I1149326);
DFFARX1 I_67460 (I1149343,I2507,I1149148,I1149369,);
not I_67461 (I1149377,I1149369);
not I_67462 (I1149394,I544617);
nand I_67463 (I1149411,I1149394,I544620);
and I_67464 (I1149428,I1149230,I1149411);
nor I_67465 (I1149445,I1149343,I1149428);
DFFARX1 I_67466 (I1149445,I2507,I1149148,I1149116,);
DFFARX1 I_67467 (I1149428,I2507,I1149148,I1149137,);
nor I_67468 (I1149490,I544617,I544596);
nor I_67469 (I1149128,I1149343,I1149490);
or I_67470 (I1149521,I544617,I544596);
nor I_67471 (I1149538,I544608,I544599);
DFFARX1 I_67472 (I1149538,I2507,I1149148,I1149564,);
not I_67473 (I1149572,I1149564);
nor I_67474 (I1149134,I1149572,I1149377);
nand I_67475 (I1149603,I1149572,I1149222);
not I_67476 (I1149620,I544608);
nand I_67477 (I1149637,I1149620,I1149326);
nand I_67478 (I1149654,I1149572,I1149637);
nand I_67479 (I1149125,I1149654,I1149603);
nand I_67480 (I1149122,I1149637,I1149521);
not I_67481 (I1149726,I2514);
DFFARX1 I_67482 (I661367,I2507,I1149726,I1149752,);
and I_67483 (I1149760,I1149752,I661355);
DFFARX1 I_67484 (I1149760,I2507,I1149726,I1149709,);
DFFARX1 I_67485 (I661358,I2507,I1149726,I1149800,);
not I_67486 (I1149808,I661352);
not I_67487 (I1149825,I661376);
nand I_67488 (I1149842,I1149825,I1149808);
nor I_67489 (I1149697,I1149800,I1149842);
DFFARX1 I_67490 (I1149842,I2507,I1149726,I1149882,);
not I_67491 (I1149718,I1149882);
not I_67492 (I1149904,I661364);
nand I_67493 (I1149921,I1149825,I1149904);
DFFARX1 I_67494 (I1149921,I2507,I1149726,I1149947,);
not I_67495 (I1149955,I1149947);
not I_67496 (I1149972,I661373);
nand I_67497 (I1149989,I1149972,I661370);
and I_67498 (I1150006,I1149808,I1149989);
nor I_67499 (I1150023,I1149921,I1150006);
DFFARX1 I_67500 (I1150023,I2507,I1149726,I1149694,);
DFFARX1 I_67501 (I1150006,I2507,I1149726,I1149715,);
nor I_67502 (I1150068,I661373,I661361);
nor I_67503 (I1149706,I1149921,I1150068);
or I_67504 (I1150099,I661373,I661361);
nor I_67505 (I1150116,I661352,I661355);
DFFARX1 I_67506 (I1150116,I2507,I1149726,I1150142,);
not I_67507 (I1150150,I1150142);
nor I_67508 (I1149712,I1150150,I1149955);
nand I_67509 (I1150181,I1150150,I1149800);
not I_67510 (I1150198,I661352);
nand I_67511 (I1150215,I1150198,I1149904);
nand I_67512 (I1150232,I1150150,I1150215);
nand I_67513 (I1149703,I1150232,I1150181);
nand I_67514 (I1149700,I1150215,I1150099);
not I_67515 (I1150304,I2514);
DFFARX1 I_67516 (I540502,I2507,I1150304,I1150330,);
and I_67517 (I1150338,I1150330,I540517);
DFFARX1 I_67518 (I1150338,I2507,I1150304,I1150287,);
DFFARX1 I_67519 (I540508,I2507,I1150304,I1150378,);
not I_67520 (I1150386,I540502);
not I_67521 (I1150403,I540520);
nand I_67522 (I1150420,I1150403,I1150386);
nor I_67523 (I1150275,I1150378,I1150420);
DFFARX1 I_67524 (I1150420,I2507,I1150304,I1150460,);
not I_67525 (I1150296,I1150460);
not I_67526 (I1150482,I540511);
nand I_67527 (I1150499,I1150403,I1150482);
DFFARX1 I_67528 (I1150499,I2507,I1150304,I1150525,);
not I_67529 (I1150533,I1150525);
not I_67530 (I1150550,I540523);
nand I_67531 (I1150567,I1150550,I540499);
and I_67532 (I1150584,I1150386,I1150567);
nor I_67533 (I1150601,I1150499,I1150584);
DFFARX1 I_67534 (I1150601,I2507,I1150304,I1150272,);
DFFARX1 I_67535 (I1150584,I2507,I1150304,I1150293,);
nor I_67536 (I1150646,I540523,I540499);
nor I_67537 (I1150284,I1150499,I1150646);
or I_67538 (I1150677,I540523,I540499);
nor I_67539 (I1150694,I540505,I540514);
DFFARX1 I_67540 (I1150694,I2507,I1150304,I1150720,);
not I_67541 (I1150728,I1150720);
nor I_67542 (I1150290,I1150728,I1150533);
nand I_67543 (I1150759,I1150728,I1150378);
not I_67544 (I1150776,I540505);
nand I_67545 (I1150793,I1150776,I1150482);
nand I_67546 (I1150810,I1150728,I1150793);
nand I_67547 (I1150281,I1150810,I1150759);
nand I_67548 (I1150278,I1150793,I1150677);
not I_67549 (I1150882,I2514);
DFFARX1 I_67550 (I56465,I2507,I1150882,I1150908,);
and I_67551 (I1150916,I1150908,I56441);
DFFARX1 I_67552 (I1150916,I2507,I1150882,I1150865,);
DFFARX1 I_67553 (I56459,I2507,I1150882,I1150956,);
not I_67554 (I1150964,I56447);
not I_67555 (I1150981,I56444);
nand I_67556 (I1150998,I1150981,I1150964);
nor I_67557 (I1150853,I1150956,I1150998);
DFFARX1 I_67558 (I1150998,I2507,I1150882,I1151038,);
not I_67559 (I1150874,I1151038);
not I_67560 (I1151060,I56453);
nand I_67561 (I1151077,I1150981,I1151060);
DFFARX1 I_67562 (I1151077,I2507,I1150882,I1151103,);
not I_67563 (I1151111,I1151103);
not I_67564 (I1151128,I56444);
nand I_67565 (I1151145,I1151128,I56462);
and I_67566 (I1151162,I1150964,I1151145);
nor I_67567 (I1151179,I1151077,I1151162);
DFFARX1 I_67568 (I1151179,I2507,I1150882,I1150850,);
DFFARX1 I_67569 (I1151162,I2507,I1150882,I1150871,);
nor I_67570 (I1151224,I56444,I56456);
nor I_67571 (I1150862,I1151077,I1151224);
or I_67572 (I1151255,I56444,I56456);
nor I_67573 (I1151272,I56450,I56441);
DFFARX1 I_67574 (I1151272,I2507,I1150882,I1151298,);
not I_67575 (I1151306,I1151298);
nor I_67576 (I1150868,I1151306,I1151111);
nand I_67577 (I1151337,I1151306,I1150956);
not I_67578 (I1151354,I56450);
nand I_67579 (I1151371,I1151354,I1151060);
nand I_67580 (I1151388,I1151306,I1151371);
nand I_67581 (I1150859,I1151388,I1151337);
nand I_67582 (I1150856,I1151371,I1151255);
not I_67583 (I1151460,I2514);
DFFARX1 I_67584 (I657899,I2507,I1151460,I1151486,);
and I_67585 (I1151494,I1151486,I657887);
DFFARX1 I_67586 (I1151494,I2507,I1151460,I1151443,);
DFFARX1 I_67587 (I657890,I2507,I1151460,I1151534,);
not I_67588 (I1151542,I657884);
not I_67589 (I1151559,I657908);
nand I_67590 (I1151576,I1151559,I1151542);
nor I_67591 (I1151431,I1151534,I1151576);
DFFARX1 I_67592 (I1151576,I2507,I1151460,I1151616,);
not I_67593 (I1151452,I1151616);
not I_67594 (I1151638,I657896);
nand I_67595 (I1151655,I1151559,I1151638);
DFFARX1 I_67596 (I1151655,I2507,I1151460,I1151681,);
not I_67597 (I1151689,I1151681);
not I_67598 (I1151706,I657905);
nand I_67599 (I1151723,I1151706,I657902);
and I_67600 (I1151740,I1151542,I1151723);
nor I_67601 (I1151757,I1151655,I1151740);
DFFARX1 I_67602 (I1151757,I2507,I1151460,I1151428,);
DFFARX1 I_67603 (I1151740,I2507,I1151460,I1151449,);
nor I_67604 (I1151802,I657905,I657893);
nor I_67605 (I1151440,I1151655,I1151802);
or I_67606 (I1151833,I657905,I657893);
nor I_67607 (I1151850,I657884,I657887);
DFFARX1 I_67608 (I1151850,I2507,I1151460,I1151876,);
not I_67609 (I1151884,I1151876);
nor I_67610 (I1151446,I1151884,I1151689);
nand I_67611 (I1151915,I1151884,I1151534);
not I_67612 (I1151932,I657884);
nand I_67613 (I1151949,I1151932,I1151638);
nand I_67614 (I1151966,I1151884,I1151949);
nand I_67615 (I1151437,I1151966,I1151915);
nand I_67616 (I1151434,I1151949,I1151833);
not I_67617 (I1152038,I2514);
DFFARX1 I_67618 (I259703,I2507,I1152038,I1152064,);
and I_67619 (I1152072,I1152064,I259688);
DFFARX1 I_67620 (I1152072,I2507,I1152038,I1152021,);
DFFARX1 I_67621 (I259694,I2507,I1152038,I1152112,);
not I_67622 (I1152120,I259676);
not I_67623 (I1152137,I259697);
nand I_67624 (I1152154,I1152137,I1152120);
nor I_67625 (I1152009,I1152112,I1152154);
DFFARX1 I_67626 (I1152154,I2507,I1152038,I1152194,);
not I_67627 (I1152030,I1152194);
not I_67628 (I1152216,I259700);
nand I_67629 (I1152233,I1152137,I1152216);
DFFARX1 I_67630 (I1152233,I2507,I1152038,I1152259,);
not I_67631 (I1152267,I1152259);
not I_67632 (I1152284,I259691);
nand I_67633 (I1152301,I1152284,I259679);
and I_67634 (I1152318,I1152120,I1152301);
nor I_67635 (I1152335,I1152233,I1152318);
DFFARX1 I_67636 (I1152335,I2507,I1152038,I1152006,);
DFFARX1 I_67637 (I1152318,I2507,I1152038,I1152027,);
nor I_67638 (I1152380,I259691,I259685);
nor I_67639 (I1152018,I1152233,I1152380);
or I_67640 (I1152411,I259691,I259685);
nor I_67641 (I1152428,I259682,I259676);
DFFARX1 I_67642 (I1152428,I2507,I1152038,I1152454,);
not I_67643 (I1152462,I1152454);
nor I_67644 (I1152024,I1152462,I1152267);
nand I_67645 (I1152493,I1152462,I1152112);
not I_67646 (I1152510,I259682);
nand I_67647 (I1152527,I1152510,I1152216);
nand I_67648 (I1152544,I1152462,I1152527);
nand I_67649 (I1152015,I1152544,I1152493);
nand I_67650 (I1152012,I1152527,I1152411);
not I_67651 (I1152616,I2514);
DFFARX1 I_67652 (I519082,I2507,I1152616,I1152642,);
and I_67653 (I1152650,I1152642,I519097);
DFFARX1 I_67654 (I1152650,I2507,I1152616,I1152599,);
DFFARX1 I_67655 (I519088,I2507,I1152616,I1152690,);
not I_67656 (I1152698,I519082);
not I_67657 (I1152715,I519100);
nand I_67658 (I1152732,I1152715,I1152698);
nor I_67659 (I1152587,I1152690,I1152732);
DFFARX1 I_67660 (I1152732,I2507,I1152616,I1152772,);
not I_67661 (I1152608,I1152772);
not I_67662 (I1152794,I519091);
nand I_67663 (I1152811,I1152715,I1152794);
DFFARX1 I_67664 (I1152811,I2507,I1152616,I1152837,);
not I_67665 (I1152845,I1152837);
not I_67666 (I1152862,I519103);
nand I_67667 (I1152879,I1152862,I519079);
and I_67668 (I1152896,I1152698,I1152879);
nor I_67669 (I1152913,I1152811,I1152896);
DFFARX1 I_67670 (I1152913,I2507,I1152616,I1152584,);
DFFARX1 I_67671 (I1152896,I2507,I1152616,I1152605,);
nor I_67672 (I1152958,I519103,I519079);
nor I_67673 (I1152596,I1152811,I1152958);
or I_67674 (I1152989,I519103,I519079);
nor I_67675 (I1153006,I519085,I519094);
DFFARX1 I_67676 (I1153006,I2507,I1152616,I1153032,);
not I_67677 (I1153040,I1153032);
nor I_67678 (I1152602,I1153040,I1152845);
nand I_67679 (I1153071,I1153040,I1152690);
not I_67680 (I1153088,I519085);
nand I_67681 (I1153105,I1153088,I1152794);
nand I_67682 (I1153122,I1153040,I1153105);
nand I_67683 (I1152593,I1153122,I1153071);
nand I_67684 (I1152590,I1153105,I1152989);
not I_67685 (I1153194,I2514);
DFFARX1 I_67686 (I1218871,I2507,I1153194,I1153220,);
and I_67687 (I1153228,I1153220,I1218865);
DFFARX1 I_67688 (I1153228,I2507,I1153194,I1153177,);
DFFARX1 I_67689 (I1218850,I2507,I1153194,I1153268,);
not I_67690 (I1153276,I1218856);
not I_67691 (I1153293,I1218868);
nand I_67692 (I1153310,I1153293,I1153276);
nor I_67693 (I1153165,I1153268,I1153310);
DFFARX1 I_67694 (I1153310,I2507,I1153194,I1153350,);
not I_67695 (I1153186,I1153350);
not I_67696 (I1153372,I1218850);
nand I_67697 (I1153389,I1153293,I1153372);
DFFARX1 I_67698 (I1153389,I2507,I1153194,I1153415,);
not I_67699 (I1153423,I1153415);
not I_67700 (I1153440,I1218874);
nand I_67701 (I1153457,I1153440,I1218862);
and I_67702 (I1153474,I1153276,I1153457);
nor I_67703 (I1153491,I1153389,I1153474);
DFFARX1 I_67704 (I1153491,I2507,I1153194,I1153162,);
DFFARX1 I_67705 (I1153474,I2507,I1153194,I1153183,);
nor I_67706 (I1153536,I1218874,I1218853);
nor I_67707 (I1153174,I1153389,I1153536);
or I_67708 (I1153567,I1218874,I1218853);
nor I_67709 (I1153584,I1218859,I1218853);
DFFARX1 I_67710 (I1153584,I2507,I1153194,I1153610,);
not I_67711 (I1153618,I1153610);
nor I_67712 (I1153180,I1153618,I1153423);
nand I_67713 (I1153649,I1153618,I1153268);
not I_67714 (I1153666,I1218859);
nand I_67715 (I1153683,I1153666,I1153372);
nand I_67716 (I1153700,I1153618,I1153683);
nand I_67717 (I1153171,I1153700,I1153649);
nand I_67718 (I1153168,I1153683,I1153567);
not I_67719 (I1153772,I2514);
DFFARX1 I_67720 (I795400,I2507,I1153772,I1153798,);
and I_67721 (I1153806,I1153798,I795406);
DFFARX1 I_67722 (I1153806,I2507,I1153772,I1153755,);
DFFARX1 I_67723 (I795412,I2507,I1153772,I1153846,);
not I_67724 (I1153854,I795397);
not I_67725 (I1153871,I795397);
nand I_67726 (I1153888,I1153871,I1153854);
nor I_67727 (I1153743,I1153846,I1153888);
DFFARX1 I_67728 (I1153888,I2507,I1153772,I1153928,);
not I_67729 (I1153764,I1153928);
not I_67730 (I1153950,I795415);
nand I_67731 (I1153967,I1153871,I1153950);
DFFARX1 I_67732 (I1153967,I2507,I1153772,I1153993,);
not I_67733 (I1154001,I1153993);
not I_67734 (I1154018,I795409);
nand I_67735 (I1154035,I1154018,I795400);
and I_67736 (I1154052,I1153854,I1154035);
nor I_67737 (I1154069,I1153967,I1154052);
DFFARX1 I_67738 (I1154069,I2507,I1153772,I1153740,);
DFFARX1 I_67739 (I1154052,I2507,I1153772,I1153761,);
nor I_67740 (I1154114,I795409,I795418);
nor I_67741 (I1153752,I1153967,I1154114);
or I_67742 (I1154145,I795409,I795418);
nor I_67743 (I1154162,I795403,I795403);
DFFARX1 I_67744 (I1154162,I2507,I1153772,I1154188,);
not I_67745 (I1154196,I1154188);
nor I_67746 (I1153758,I1154196,I1154001);
nand I_67747 (I1154227,I1154196,I1153846);
not I_67748 (I1154244,I795403);
nand I_67749 (I1154261,I1154244,I1153950);
nand I_67750 (I1154278,I1154196,I1154261);
nand I_67751 (I1153749,I1154278,I1154227);
nand I_67752 (I1153746,I1154261,I1154145);
not I_67753 (I1154350,I2514);
DFFARX1 I_67754 (I341388,I2507,I1154350,I1154376,);
and I_67755 (I1154384,I1154376,I341373);
DFFARX1 I_67756 (I1154384,I2507,I1154350,I1154333,);
DFFARX1 I_67757 (I341379,I2507,I1154350,I1154424,);
not I_67758 (I1154432,I341361);
not I_67759 (I1154449,I341382);
nand I_67760 (I1154466,I1154449,I1154432);
nor I_67761 (I1154321,I1154424,I1154466);
DFFARX1 I_67762 (I1154466,I2507,I1154350,I1154506,);
not I_67763 (I1154342,I1154506);
not I_67764 (I1154528,I341385);
nand I_67765 (I1154545,I1154449,I1154528);
DFFARX1 I_67766 (I1154545,I2507,I1154350,I1154571,);
not I_67767 (I1154579,I1154571);
not I_67768 (I1154596,I341376);
nand I_67769 (I1154613,I1154596,I341364);
and I_67770 (I1154630,I1154432,I1154613);
nor I_67771 (I1154647,I1154545,I1154630);
DFFARX1 I_67772 (I1154647,I2507,I1154350,I1154318,);
DFFARX1 I_67773 (I1154630,I2507,I1154350,I1154339,);
nor I_67774 (I1154692,I341376,I341370);
nor I_67775 (I1154330,I1154545,I1154692);
or I_67776 (I1154723,I341376,I341370);
nor I_67777 (I1154740,I341367,I341361);
DFFARX1 I_67778 (I1154740,I2507,I1154350,I1154766,);
not I_67779 (I1154774,I1154766);
nor I_67780 (I1154336,I1154774,I1154579);
nand I_67781 (I1154805,I1154774,I1154424);
not I_67782 (I1154822,I341367);
nand I_67783 (I1154839,I1154822,I1154528);
nand I_67784 (I1154856,I1154774,I1154839);
nand I_67785 (I1154327,I1154856,I1154805);
nand I_67786 (I1154324,I1154839,I1154723);
not I_67787 (I1154928,I2514);
DFFARX1 I_67788 (I1346989,I2507,I1154928,I1154954,);
and I_67789 (I1154962,I1154954,I1346971);
DFFARX1 I_67790 (I1154962,I2507,I1154928,I1154911,);
DFFARX1 I_67791 (I1346962,I2507,I1154928,I1155002,);
not I_67792 (I1155010,I1346977);
not I_67793 (I1155027,I1346965);
nand I_67794 (I1155044,I1155027,I1155010);
nor I_67795 (I1154899,I1155002,I1155044);
DFFARX1 I_67796 (I1155044,I2507,I1154928,I1155084,);
not I_67797 (I1154920,I1155084);
not I_67798 (I1155106,I1346974);
nand I_67799 (I1155123,I1155027,I1155106);
DFFARX1 I_67800 (I1155123,I2507,I1154928,I1155149,);
not I_67801 (I1155157,I1155149);
not I_67802 (I1155174,I1346983);
nand I_67803 (I1155191,I1155174,I1346962);
and I_67804 (I1155208,I1155010,I1155191);
nor I_67805 (I1155225,I1155123,I1155208);
DFFARX1 I_67806 (I1155225,I2507,I1154928,I1154896,);
DFFARX1 I_67807 (I1155208,I2507,I1154928,I1154917,);
nor I_67808 (I1155270,I1346983,I1346986);
nor I_67809 (I1154908,I1155123,I1155270);
or I_67810 (I1155301,I1346983,I1346986);
nor I_67811 (I1155318,I1346980,I1346968);
DFFARX1 I_67812 (I1155318,I2507,I1154928,I1155344,);
not I_67813 (I1155352,I1155344);
nor I_67814 (I1154914,I1155352,I1155157);
nand I_67815 (I1155383,I1155352,I1155002);
not I_67816 (I1155400,I1346980);
nand I_67817 (I1155417,I1155400,I1155106);
nand I_67818 (I1155434,I1155352,I1155417);
nand I_67819 (I1154905,I1155434,I1155383);
nand I_67820 (I1154902,I1155417,I1155301);
not I_67821 (I1155506,I2514);
DFFARX1 I_67822 (I827547,I2507,I1155506,I1155532,);
and I_67823 (I1155540,I1155532,I827553);
DFFARX1 I_67824 (I1155540,I2507,I1155506,I1155489,);
DFFARX1 I_67825 (I827559,I2507,I1155506,I1155580,);
not I_67826 (I1155588,I827544);
not I_67827 (I1155605,I827544);
nand I_67828 (I1155622,I1155605,I1155588);
nor I_67829 (I1155477,I1155580,I1155622);
DFFARX1 I_67830 (I1155622,I2507,I1155506,I1155662,);
not I_67831 (I1155498,I1155662);
not I_67832 (I1155684,I827562);
nand I_67833 (I1155701,I1155605,I1155684);
DFFARX1 I_67834 (I1155701,I2507,I1155506,I1155727,);
not I_67835 (I1155735,I1155727);
not I_67836 (I1155752,I827556);
nand I_67837 (I1155769,I1155752,I827547);
and I_67838 (I1155786,I1155588,I1155769);
nor I_67839 (I1155803,I1155701,I1155786);
DFFARX1 I_67840 (I1155803,I2507,I1155506,I1155474,);
DFFARX1 I_67841 (I1155786,I2507,I1155506,I1155495,);
nor I_67842 (I1155848,I827556,I827565);
nor I_67843 (I1155486,I1155701,I1155848);
or I_67844 (I1155879,I827556,I827565);
nor I_67845 (I1155896,I827550,I827550);
DFFARX1 I_67846 (I1155896,I2507,I1155506,I1155922,);
not I_67847 (I1155930,I1155922);
nor I_67848 (I1155492,I1155930,I1155735);
nand I_67849 (I1155961,I1155930,I1155580);
not I_67850 (I1155978,I827550);
nand I_67851 (I1155995,I1155978,I1155684);
nand I_67852 (I1156012,I1155930,I1155995);
nand I_67853 (I1155483,I1156012,I1155961);
nand I_67854 (I1155480,I1155995,I1155879);
not I_67855 (I1156084,I2514);
DFFARX1 I_67856 (I1052780,I2507,I1156084,I1156110,);
and I_67857 (I1156118,I1156110,I1052777);
DFFARX1 I_67858 (I1156118,I2507,I1156084,I1156067,);
DFFARX1 I_67859 (I1052783,I2507,I1156084,I1156158,);
not I_67860 (I1156166,I1052786);
not I_67861 (I1156183,I1052780);
nand I_67862 (I1156200,I1156183,I1156166);
nor I_67863 (I1156055,I1156158,I1156200);
DFFARX1 I_67864 (I1156200,I2507,I1156084,I1156240,);
not I_67865 (I1156076,I1156240);
not I_67866 (I1156262,I1052795);
nand I_67867 (I1156279,I1156183,I1156262);
DFFARX1 I_67868 (I1156279,I2507,I1156084,I1156305,);
not I_67869 (I1156313,I1156305);
not I_67870 (I1156330,I1052792);
nand I_67871 (I1156347,I1156330,I1052798);
and I_67872 (I1156364,I1156166,I1156347);
nor I_67873 (I1156381,I1156279,I1156364);
DFFARX1 I_67874 (I1156381,I2507,I1156084,I1156052,);
DFFARX1 I_67875 (I1156364,I2507,I1156084,I1156073,);
nor I_67876 (I1156426,I1052792,I1052777);
nor I_67877 (I1156064,I1156279,I1156426);
or I_67878 (I1156457,I1052792,I1052777);
nor I_67879 (I1156474,I1052789,I1052783);
DFFARX1 I_67880 (I1156474,I2507,I1156084,I1156500,);
not I_67881 (I1156508,I1156500);
nor I_67882 (I1156070,I1156508,I1156313);
nand I_67883 (I1156539,I1156508,I1156158);
not I_67884 (I1156556,I1052789);
nand I_67885 (I1156573,I1156556,I1156262);
nand I_67886 (I1156590,I1156508,I1156573);
nand I_67887 (I1156061,I1156590,I1156539);
nand I_67888 (I1156058,I1156573,I1156457);
not I_67889 (I1156662,I2514);
DFFARX1 I_67890 (I399535,I2507,I1156662,I1156688,);
and I_67891 (I1156696,I1156688,I399550);
DFFARX1 I_67892 (I1156696,I2507,I1156662,I1156645,);
DFFARX1 I_67893 (I399553,I2507,I1156662,I1156736,);
not I_67894 (I1156744,I399547);
not I_67895 (I1156761,I399562);
nand I_67896 (I1156778,I1156761,I1156744);
nor I_67897 (I1156633,I1156736,I1156778);
DFFARX1 I_67898 (I1156778,I2507,I1156662,I1156818,);
not I_67899 (I1156654,I1156818);
not I_67900 (I1156840,I399538);
nand I_67901 (I1156857,I1156761,I1156840);
DFFARX1 I_67902 (I1156857,I2507,I1156662,I1156883,);
not I_67903 (I1156891,I1156883);
not I_67904 (I1156908,I399541);
nand I_67905 (I1156925,I1156908,I399535);
and I_67906 (I1156942,I1156744,I1156925);
nor I_67907 (I1156959,I1156857,I1156942);
DFFARX1 I_67908 (I1156959,I2507,I1156662,I1156630,);
DFFARX1 I_67909 (I1156942,I2507,I1156662,I1156651,);
nor I_67910 (I1157004,I399541,I399544);
nor I_67911 (I1156642,I1156857,I1157004);
or I_67912 (I1157035,I399541,I399544);
nor I_67913 (I1157052,I399559,I399556);
DFFARX1 I_67914 (I1157052,I2507,I1156662,I1157078,);
not I_67915 (I1157086,I1157078);
nor I_67916 (I1156648,I1157086,I1156891);
nand I_67917 (I1157117,I1157086,I1156736);
not I_67918 (I1157134,I399559);
nand I_67919 (I1157151,I1157134,I1156840);
nand I_67920 (I1157168,I1157086,I1157151);
nand I_67921 (I1156639,I1157168,I1157117);
nand I_67922 (I1156636,I1157151,I1157035);
not I_67923 (I1157240,I2514);
DFFARX1 I_67924 (I99679,I2507,I1157240,I1157266,);
and I_67925 (I1157274,I1157266,I99655);
DFFARX1 I_67926 (I1157274,I2507,I1157240,I1157223,);
DFFARX1 I_67927 (I99673,I2507,I1157240,I1157314,);
not I_67928 (I1157322,I99661);
not I_67929 (I1157339,I99658);
nand I_67930 (I1157356,I1157339,I1157322);
nor I_67931 (I1157211,I1157314,I1157356);
DFFARX1 I_67932 (I1157356,I2507,I1157240,I1157396,);
not I_67933 (I1157232,I1157396);
not I_67934 (I1157418,I99667);
nand I_67935 (I1157435,I1157339,I1157418);
DFFARX1 I_67936 (I1157435,I2507,I1157240,I1157461,);
not I_67937 (I1157469,I1157461);
not I_67938 (I1157486,I99658);
nand I_67939 (I1157503,I1157486,I99676);
and I_67940 (I1157520,I1157322,I1157503);
nor I_67941 (I1157537,I1157435,I1157520);
DFFARX1 I_67942 (I1157537,I2507,I1157240,I1157208,);
DFFARX1 I_67943 (I1157520,I2507,I1157240,I1157229,);
nor I_67944 (I1157582,I99658,I99670);
nor I_67945 (I1157220,I1157435,I1157582);
or I_67946 (I1157613,I99658,I99670);
nor I_67947 (I1157630,I99664,I99655);
DFFARX1 I_67948 (I1157630,I2507,I1157240,I1157656,);
not I_67949 (I1157664,I1157656);
nor I_67950 (I1157226,I1157664,I1157469);
nand I_67951 (I1157695,I1157664,I1157314);
not I_67952 (I1157712,I99664);
nand I_67953 (I1157729,I1157712,I1157418);
nand I_67954 (I1157746,I1157664,I1157729);
nand I_67955 (I1157217,I1157746,I1157695);
nand I_67956 (I1157214,I1157729,I1157613);
not I_67957 (I1157818,I2514);
DFFARX1 I_67958 (I477871,I2507,I1157818,I1157844,);
and I_67959 (I1157852,I1157844,I477886);
DFFARX1 I_67960 (I1157852,I2507,I1157818,I1157801,);
DFFARX1 I_67961 (I477889,I2507,I1157818,I1157892,);
not I_67962 (I1157900,I477883);
not I_67963 (I1157917,I477898);
nand I_67964 (I1157934,I1157917,I1157900);
nor I_67965 (I1157789,I1157892,I1157934);
DFFARX1 I_67966 (I1157934,I2507,I1157818,I1157974,);
not I_67967 (I1157810,I1157974);
not I_67968 (I1157996,I477874);
nand I_67969 (I1158013,I1157917,I1157996);
DFFARX1 I_67970 (I1158013,I2507,I1157818,I1158039,);
not I_67971 (I1158047,I1158039);
not I_67972 (I1158064,I477877);
nand I_67973 (I1158081,I1158064,I477871);
and I_67974 (I1158098,I1157900,I1158081);
nor I_67975 (I1158115,I1158013,I1158098);
DFFARX1 I_67976 (I1158115,I2507,I1157818,I1157786,);
DFFARX1 I_67977 (I1158098,I2507,I1157818,I1157807,);
nor I_67978 (I1158160,I477877,I477880);
nor I_67979 (I1157798,I1158013,I1158160);
or I_67980 (I1158191,I477877,I477880);
nor I_67981 (I1158208,I477895,I477892);
DFFARX1 I_67982 (I1158208,I2507,I1157818,I1158234,);
not I_67983 (I1158242,I1158234);
nor I_67984 (I1157804,I1158242,I1158047);
nand I_67985 (I1158273,I1158242,I1157892);
not I_67986 (I1158290,I477895);
nand I_67987 (I1158307,I1158290,I1157996);
nand I_67988 (I1158324,I1158242,I1158307);
nand I_67989 (I1157795,I1158324,I1158273);
nand I_67990 (I1157792,I1158307,I1158191);
not I_67991 (I1158396,I2514);
DFFARX1 I_67992 (I1248791,I2507,I1158396,I1158422,);
and I_67993 (I1158430,I1158422,I1248785);
DFFARX1 I_67994 (I1158430,I2507,I1158396,I1158379,);
DFFARX1 I_67995 (I1248770,I2507,I1158396,I1158470,);
not I_67996 (I1158478,I1248776);
not I_67997 (I1158495,I1248788);
nand I_67998 (I1158512,I1158495,I1158478);
nor I_67999 (I1158367,I1158470,I1158512);
DFFARX1 I_68000 (I1158512,I2507,I1158396,I1158552,);
not I_68001 (I1158388,I1158552);
not I_68002 (I1158574,I1248770);
nand I_68003 (I1158591,I1158495,I1158574);
DFFARX1 I_68004 (I1158591,I2507,I1158396,I1158617,);
not I_68005 (I1158625,I1158617);
not I_68006 (I1158642,I1248794);
nand I_68007 (I1158659,I1158642,I1248782);
and I_68008 (I1158676,I1158478,I1158659);
nor I_68009 (I1158693,I1158591,I1158676);
DFFARX1 I_68010 (I1158693,I2507,I1158396,I1158364,);
DFFARX1 I_68011 (I1158676,I2507,I1158396,I1158385,);
nor I_68012 (I1158738,I1248794,I1248773);
nor I_68013 (I1158376,I1158591,I1158738);
or I_68014 (I1158769,I1248794,I1248773);
nor I_68015 (I1158786,I1248779,I1248773);
DFFARX1 I_68016 (I1158786,I2507,I1158396,I1158812,);
not I_68017 (I1158820,I1158812);
nor I_68018 (I1158382,I1158820,I1158625);
nand I_68019 (I1158851,I1158820,I1158470);
not I_68020 (I1158868,I1248779);
nand I_68021 (I1158885,I1158868,I1158574);
nand I_68022 (I1158902,I1158820,I1158885);
nand I_68023 (I1158373,I1158902,I1158851);
nand I_68024 (I1158370,I1158885,I1158769);
not I_68025 (I1158974,I2514);
DFFARX1 I_68026 (I813845,I2507,I1158974,I1159000,);
and I_68027 (I1159008,I1159000,I813851);
DFFARX1 I_68028 (I1159008,I2507,I1158974,I1158957,);
DFFARX1 I_68029 (I813857,I2507,I1158974,I1159048,);
not I_68030 (I1159056,I813842);
not I_68031 (I1159073,I813842);
nand I_68032 (I1159090,I1159073,I1159056);
nor I_68033 (I1158945,I1159048,I1159090);
DFFARX1 I_68034 (I1159090,I2507,I1158974,I1159130,);
not I_68035 (I1158966,I1159130);
not I_68036 (I1159152,I813860);
nand I_68037 (I1159169,I1159073,I1159152);
DFFARX1 I_68038 (I1159169,I2507,I1158974,I1159195,);
not I_68039 (I1159203,I1159195);
not I_68040 (I1159220,I813854);
nand I_68041 (I1159237,I1159220,I813845);
and I_68042 (I1159254,I1159056,I1159237);
nor I_68043 (I1159271,I1159169,I1159254);
DFFARX1 I_68044 (I1159271,I2507,I1158974,I1158942,);
DFFARX1 I_68045 (I1159254,I2507,I1158974,I1158963,);
nor I_68046 (I1159316,I813854,I813863);
nor I_68047 (I1158954,I1159169,I1159316);
or I_68048 (I1159347,I813854,I813863);
nor I_68049 (I1159364,I813848,I813848);
DFFARX1 I_68050 (I1159364,I2507,I1158974,I1159390,);
not I_68051 (I1159398,I1159390);
nor I_68052 (I1158960,I1159398,I1159203);
nand I_68053 (I1159429,I1159398,I1159048);
not I_68054 (I1159446,I813848);
nand I_68055 (I1159463,I1159446,I1159152);
nand I_68056 (I1159480,I1159398,I1159463);
nand I_68057 (I1158951,I1159480,I1159429);
nand I_68058 (I1158948,I1159463,I1159347);
not I_68059 (I1159552,I2514);
DFFARX1 I_68060 (I809629,I2507,I1159552,I1159578,);
and I_68061 (I1159586,I1159578,I809635);
DFFARX1 I_68062 (I1159586,I2507,I1159552,I1159535,);
DFFARX1 I_68063 (I809641,I2507,I1159552,I1159626,);
not I_68064 (I1159634,I809626);
not I_68065 (I1159651,I809626);
nand I_68066 (I1159668,I1159651,I1159634);
nor I_68067 (I1159523,I1159626,I1159668);
DFFARX1 I_68068 (I1159668,I2507,I1159552,I1159708,);
not I_68069 (I1159544,I1159708);
not I_68070 (I1159730,I809644);
nand I_68071 (I1159747,I1159651,I1159730);
DFFARX1 I_68072 (I1159747,I2507,I1159552,I1159773,);
not I_68073 (I1159781,I1159773);
not I_68074 (I1159798,I809638);
nand I_68075 (I1159815,I1159798,I809629);
and I_68076 (I1159832,I1159634,I1159815);
nor I_68077 (I1159849,I1159747,I1159832);
DFFARX1 I_68078 (I1159849,I2507,I1159552,I1159520,);
DFFARX1 I_68079 (I1159832,I2507,I1159552,I1159541,);
nor I_68080 (I1159894,I809638,I809647);
nor I_68081 (I1159532,I1159747,I1159894);
or I_68082 (I1159925,I809638,I809647);
nor I_68083 (I1159942,I809632,I809632);
DFFARX1 I_68084 (I1159942,I2507,I1159552,I1159968,);
not I_68085 (I1159976,I1159968);
nor I_68086 (I1159538,I1159976,I1159781);
nand I_68087 (I1160007,I1159976,I1159626);
not I_68088 (I1160024,I809632);
nand I_68089 (I1160041,I1160024,I1159730);
nand I_68090 (I1160058,I1159976,I1160041);
nand I_68091 (I1159529,I1160058,I1160007);
nand I_68092 (I1159526,I1160041,I1159925);
not I_68093 (I1160130,I2514);
DFFARX1 I_68094 (I455567,I2507,I1160130,I1160156,);
and I_68095 (I1160164,I1160156,I455582);
DFFARX1 I_68096 (I1160164,I2507,I1160130,I1160113,);
DFFARX1 I_68097 (I455585,I2507,I1160130,I1160204,);
not I_68098 (I1160212,I455579);
not I_68099 (I1160229,I455594);
nand I_68100 (I1160246,I1160229,I1160212);
nor I_68101 (I1160101,I1160204,I1160246);
DFFARX1 I_68102 (I1160246,I2507,I1160130,I1160286,);
not I_68103 (I1160122,I1160286);
not I_68104 (I1160308,I455570);
nand I_68105 (I1160325,I1160229,I1160308);
DFFARX1 I_68106 (I1160325,I2507,I1160130,I1160351,);
not I_68107 (I1160359,I1160351);
not I_68108 (I1160376,I455573);
nand I_68109 (I1160393,I1160376,I455567);
and I_68110 (I1160410,I1160212,I1160393);
nor I_68111 (I1160427,I1160325,I1160410);
DFFARX1 I_68112 (I1160427,I2507,I1160130,I1160098,);
DFFARX1 I_68113 (I1160410,I2507,I1160130,I1160119,);
nor I_68114 (I1160472,I455573,I455576);
nor I_68115 (I1160110,I1160325,I1160472);
or I_68116 (I1160503,I455573,I455576);
nor I_68117 (I1160520,I455591,I455588);
DFFARX1 I_68118 (I1160520,I2507,I1160130,I1160546,);
not I_68119 (I1160554,I1160546);
nor I_68120 (I1160116,I1160554,I1160359);
nand I_68121 (I1160585,I1160554,I1160204);
not I_68122 (I1160602,I455591);
nand I_68123 (I1160619,I1160602,I1160308);
nand I_68124 (I1160636,I1160554,I1160619);
nand I_68125 (I1160107,I1160636,I1160585);
nand I_68126 (I1160104,I1160619,I1160503);
not I_68127 (I1160708,I2514);
DFFARX1 I_68128 (I857586,I2507,I1160708,I1160734,);
and I_68129 (I1160742,I1160734,I857592);
DFFARX1 I_68130 (I1160742,I2507,I1160708,I1160691,);
DFFARX1 I_68131 (I857598,I2507,I1160708,I1160782,);
not I_68132 (I1160790,I857583);
not I_68133 (I1160807,I857583);
nand I_68134 (I1160824,I1160807,I1160790);
nor I_68135 (I1160679,I1160782,I1160824);
DFFARX1 I_68136 (I1160824,I2507,I1160708,I1160864,);
not I_68137 (I1160700,I1160864);
not I_68138 (I1160886,I857601);
nand I_68139 (I1160903,I1160807,I1160886);
DFFARX1 I_68140 (I1160903,I2507,I1160708,I1160929,);
not I_68141 (I1160937,I1160929);
not I_68142 (I1160954,I857595);
nand I_68143 (I1160971,I1160954,I857586);
and I_68144 (I1160988,I1160790,I1160971);
nor I_68145 (I1161005,I1160903,I1160988);
DFFARX1 I_68146 (I1161005,I2507,I1160708,I1160676,);
DFFARX1 I_68147 (I1160988,I2507,I1160708,I1160697,);
nor I_68148 (I1161050,I857595,I857604);
nor I_68149 (I1160688,I1160903,I1161050);
or I_68150 (I1161081,I857595,I857604);
nor I_68151 (I1161098,I857589,I857589);
DFFARX1 I_68152 (I1161098,I2507,I1160708,I1161124,);
not I_68153 (I1161132,I1161124);
nor I_68154 (I1160694,I1161132,I1160937);
nand I_68155 (I1161163,I1161132,I1160782);
not I_68156 (I1161180,I857589);
nand I_68157 (I1161197,I1161180,I1160886);
nand I_68158 (I1161214,I1161132,I1161197);
nand I_68159 (I1160685,I1161214,I1161163);
nand I_68160 (I1160682,I1161197,I1161081);
not I_68161 (I1161286,I2514);
DFFARX1 I_68162 (I481679,I2507,I1161286,I1161312,);
and I_68163 (I1161320,I1161312,I481694);
DFFARX1 I_68164 (I1161320,I2507,I1161286,I1161269,);
DFFARX1 I_68165 (I481697,I2507,I1161286,I1161360,);
not I_68166 (I1161368,I481691);
not I_68167 (I1161385,I481706);
nand I_68168 (I1161402,I1161385,I1161368);
nor I_68169 (I1161257,I1161360,I1161402);
DFFARX1 I_68170 (I1161402,I2507,I1161286,I1161442,);
not I_68171 (I1161278,I1161442);
not I_68172 (I1161464,I481682);
nand I_68173 (I1161481,I1161385,I1161464);
DFFARX1 I_68174 (I1161481,I2507,I1161286,I1161507,);
not I_68175 (I1161515,I1161507);
not I_68176 (I1161532,I481685);
nand I_68177 (I1161549,I1161532,I481679);
and I_68178 (I1161566,I1161368,I1161549);
nor I_68179 (I1161583,I1161481,I1161566);
DFFARX1 I_68180 (I1161583,I2507,I1161286,I1161254,);
DFFARX1 I_68181 (I1161566,I2507,I1161286,I1161275,);
nor I_68182 (I1161628,I481685,I481688);
nor I_68183 (I1161266,I1161481,I1161628);
or I_68184 (I1161659,I481685,I481688);
nor I_68185 (I1161676,I481703,I481700);
DFFARX1 I_68186 (I1161676,I2507,I1161286,I1161702,);
not I_68187 (I1161710,I1161702);
nor I_68188 (I1161272,I1161710,I1161515);
nand I_68189 (I1161741,I1161710,I1161360);
not I_68190 (I1161758,I481703);
nand I_68191 (I1161775,I1161758,I1161464);
nand I_68192 (I1161792,I1161710,I1161775);
nand I_68193 (I1161263,I1161792,I1161741);
nand I_68194 (I1161260,I1161775,I1161659);
not I_68195 (I1161864,I2514);
DFFARX1 I_68196 (I815426,I2507,I1161864,I1161890,);
and I_68197 (I1161898,I1161890,I815432);
DFFARX1 I_68198 (I1161898,I2507,I1161864,I1161847,);
DFFARX1 I_68199 (I815438,I2507,I1161864,I1161938,);
not I_68200 (I1161946,I815423);
not I_68201 (I1161963,I815423);
nand I_68202 (I1161980,I1161963,I1161946);
nor I_68203 (I1161835,I1161938,I1161980);
DFFARX1 I_68204 (I1161980,I2507,I1161864,I1162020,);
not I_68205 (I1161856,I1162020);
not I_68206 (I1162042,I815441);
nand I_68207 (I1162059,I1161963,I1162042);
DFFARX1 I_68208 (I1162059,I2507,I1161864,I1162085,);
not I_68209 (I1162093,I1162085);
not I_68210 (I1162110,I815435);
nand I_68211 (I1162127,I1162110,I815426);
and I_68212 (I1162144,I1161946,I1162127);
nor I_68213 (I1162161,I1162059,I1162144);
DFFARX1 I_68214 (I1162161,I2507,I1161864,I1161832,);
DFFARX1 I_68215 (I1162144,I2507,I1161864,I1161853,);
nor I_68216 (I1162206,I815435,I815444);
nor I_68217 (I1161844,I1162059,I1162206);
or I_68218 (I1162237,I815435,I815444);
nor I_68219 (I1162254,I815429,I815429);
DFFARX1 I_68220 (I1162254,I2507,I1161864,I1162280,);
not I_68221 (I1162288,I1162280);
nor I_68222 (I1161850,I1162288,I1162093);
nand I_68223 (I1162319,I1162288,I1161938);
not I_68224 (I1162336,I815429);
nand I_68225 (I1162353,I1162336,I1162042);
nand I_68226 (I1162370,I1162288,I1162353);
nand I_68227 (I1161841,I1162370,I1162319);
nand I_68228 (I1161838,I1162353,I1162237);
not I_68229 (I1162442,I2514);
DFFARX1 I_68230 (I741709,I2507,I1162442,I1162468,);
and I_68231 (I1162476,I1162468,I741697);
DFFARX1 I_68232 (I1162476,I2507,I1162442,I1162425,);
DFFARX1 I_68233 (I741700,I2507,I1162442,I1162516,);
not I_68234 (I1162524,I741694);
not I_68235 (I1162541,I741718);
nand I_68236 (I1162558,I1162541,I1162524);
nor I_68237 (I1162413,I1162516,I1162558);
DFFARX1 I_68238 (I1162558,I2507,I1162442,I1162598,);
not I_68239 (I1162434,I1162598);
not I_68240 (I1162620,I741706);
nand I_68241 (I1162637,I1162541,I1162620);
DFFARX1 I_68242 (I1162637,I2507,I1162442,I1162663,);
not I_68243 (I1162671,I1162663);
not I_68244 (I1162688,I741715);
nand I_68245 (I1162705,I1162688,I741712);
and I_68246 (I1162722,I1162524,I1162705);
nor I_68247 (I1162739,I1162637,I1162722);
DFFARX1 I_68248 (I1162739,I2507,I1162442,I1162410,);
DFFARX1 I_68249 (I1162722,I2507,I1162442,I1162431,);
nor I_68250 (I1162784,I741715,I741703);
nor I_68251 (I1162422,I1162637,I1162784);
or I_68252 (I1162815,I741715,I741703);
nor I_68253 (I1162832,I741694,I741697);
DFFARX1 I_68254 (I1162832,I2507,I1162442,I1162858,);
not I_68255 (I1162866,I1162858);
nor I_68256 (I1162428,I1162866,I1162671);
nand I_68257 (I1162897,I1162866,I1162516);
not I_68258 (I1162914,I741694);
nand I_68259 (I1162931,I1162914,I1162620);
nand I_68260 (I1162948,I1162866,I1162931);
nand I_68261 (I1162419,I1162948,I1162897);
nand I_68262 (I1162416,I1162931,I1162815);
not I_68263 (I1163020,I2514);
DFFARX1 I_68264 (I386479,I2507,I1163020,I1163046,);
and I_68265 (I1163054,I1163046,I386494);
DFFARX1 I_68266 (I1163054,I2507,I1163020,I1163003,);
DFFARX1 I_68267 (I386497,I2507,I1163020,I1163094,);
not I_68268 (I1163102,I386491);
not I_68269 (I1163119,I386506);
nand I_68270 (I1163136,I1163119,I1163102);
nor I_68271 (I1162991,I1163094,I1163136);
DFFARX1 I_68272 (I1163136,I2507,I1163020,I1163176,);
not I_68273 (I1163012,I1163176);
not I_68274 (I1163198,I386482);
nand I_68275 (I1163215,I1163119,I1163198);
DFFARX1 I_68276 (I1163215,I2507,I1163020,I1163241,);
not I_68277 (I1163249,I1163241);
not I_68278 (I1163266,I386485);
nand I_68279 (I1163283,I1163266,I386479);
and I_68280 (I1163300,I1163102,I1163283);
nor I_68281 (I1163317,I1163215,I1163300);
DFFARX1 I_68282 (I1163317,I2507,I1163020,I1162988,);
DFFARX1 I_68283 (I1163300,I2507,I1163020,I1163009,);
nor I_68284 (I1163362,I386485,I386488);
nor I_68285 (I1163000,I1163215,I1163362);
or I_68286 (I1163393,I386485,I386488);
nor I_68287 (I1163410,I386503,I386500);
DFFARX1 I_68288 (I1163410,I2507,I1163020,I1163436,);
not I_68289 (I1163444,I1163436);
nor I_68290 (I1163006,I1163444,I1163249);
nand I_68291 (I1163475,I1163444,I1163094);
not I_68292 (I1163492,I386503);
nand I_68293 (I1163509,I1163492,I1163198);
nand I_68294 (I1163526,I1163444,I1163509);
nand I_68295 (I1162997,I1163526,I1163475);
nand I_68296 (I1162994,I1163509,I1163393);
not I_68297 (I1163598,I2514);
DFFARX1 I_68298 (I1232471,I2507,I1163598,I1163624,);
and I_68299 (I1163632,I1163624,I1232465);
DFFARX1 I_68300 (I1163632,I2507,I1163598,I1163581,);
DFFARX1 I_68301 (I1232450,I2507,I1163598,I1163672,);
not I_68302 (I1163680,I1232456);
not I_68303 (I1163697,I1232468);
nand I_68304 (I1163714,I1163697,I1163680);
nor I_68305 (I1163569,I1163672,I1163714);
DFFARX1 I_68306 (I1163714,I2507,I1163598,I1163754,);
not I_68307 (I1163590,I1163754);
not I_68308 (I1163776,I1232450);
nand I_68309 (I1163793,I1163697,I1163776);
DFFARX1 I_68310 (I1163793,I2507,I1163598,I1163819,);
not I_68311 (I1163827,I1163819);
not I_68312 (I1163844,I1232474);
nand I_68313 (I1163861,I1163844,I1232462);
and I_68314 (I1163878,I1163680,I1163861);
nor I_68315 (I1163895,I1163793,I1163878);
DFFARX1 I_68316 (I1163895,I2507,I1163598,I1163566,);
DFFARX1 I_68317 (I1163878,I2507,I1163598,I1163587,);
nor I_68318 (I1163940,I1232474,I1232453);
nor I_68319 (I1163578,I1163793,I1163940);
or I_68320 (I1163971,I1232474,I1232453);
nor I_68321 (I1163988,I1232459,I1232453);
DFFARX1 I_68322 (I1163988,I2507,I1163598,I1164014,);
not I_68323 (I1164022,I1164014);
nor I_68324 (I1163584,I1164022,I1163827);
nand I_68325 (I1164053,I1164022,I1163672);
not I_68326 (I1164070,I1232459);
nand I_68327 (I1164087,I1164070,I1163776);
nand I_68328 (I1164104,I1164022,I1164087);
nand I_68329 (I1163575,I1164104,I1164053);
nand I_68330 (I1163572,I1164087,I1163971);
not I_68331 (I1164176,I2514);
DFFARX1 I_68332 (I825966,I2507,I1164176,I1164202,);
and I_68333 (I1164210,I1164202,I825972);
DFFARX1 I_68334 (I1164210,I2507,I1164176,I1164159,);
DFFARX1 I_68335 (I825978,I2507,I1164176,I1164250,);
not I_68336 (I1164258,I825963);
not I_68337 (I1164275,I825963);
nand I_68338 (I1164292,I1164275,I1164258);
nor I_68339 (I1164147,I1164250,I1164292);
DFFARX1 I_68340 (I1164292,I2507,I1164176,I1164332,);
not I_68341 (I1164168,I1164332);
not I_68342 (I1164354,I825981);
nand I_68343 (I1164371,I1164275,I1164354);
DFFARX1 I_68344 (I1164371,I2507,I1164176,I1164397,);
not I_68345 (I1164405,I1164397);
not I_68346 (I1164422,I825975);
nand I_68347 (I1164439,I1164422,I825966);
and I_68348 (I1164456,I1164258,I1164439);
nor I_68349 (I1164473,I1164371,I1164456);
DFFARX1 I_68350 (I1164473,I2507,I1164176,I1164144,);
DFFARX1 I_68351 (I1164456,I2507,I1164176,I1164165,);
nor I_68352 (I1164518,I825975,I825984);
nor I_68353 (I1164156,I1164371,I1164518);
or I_68354 (I1164549,I825975,I825984);
nor I_68355 (I1164566,I825969,I825969);
DFFARX1 I_68356 (I1164566,I2507,I1164176,I1164592,);
not I_68357 (I1164600,I1164592);
nor I_68358 (I1164162,I1164600,I1164405);
nand I_68359 (I1164631,I1164600,I1164250);
not I_68360 (I1164648,I825969);
nand I_68361 (I1164665,I1164648,I1164354);
nand I_68362 (I1164682,I1164600,I1164665);
nand I_68363 (I1164153,I1164682,I1164631);
nand I_68364 (I1164150,I1164665,I1164549);
not I_68365 (I1164754,I2514);
DFFARX1 I_68366 (I1299736,I2507,I1164754,I1164780,);
and I_68367 (I1164788,I1164780,I1299763);
DFFARX1 I_68368 (I1164788,I2507,I1164754,I1164737,);
DFFARX1 I_68369 (I1299745,I2507,I1164754,I1164828,);
not I_68370 (I1164836,I1299754);
not I_68371 (I1164853,I1299757);
nand I_68372 (I1164870,I1164853,I1164836);
nor I_68373 (I1164725,I1164828,I1164870);
DFFARX1 I_68374 (I1164870,I2507,I1164754,I1164910,);
not I_68375 (I1164746,I1164910);
not I_68376 (I1164932,I1299751);
nand I_68377 (I1164949,I1164853,I1164932);
DFFARX1 I_68378 (I1164949,I2507,I1164754,I1164975,);
not I_68379 (I1164983,I1164975);
not I_68380 (I1165000,I1299739);
nand I_68381 (I1165017,I1165000,I1299742);
and I_68382 (I1165034,I1164836,I1165017);
nor I_68383 (I1165051,I1164949,I1165034);
DFFARX1 I_68384 (I1165051,I2507,I1164754,I1164722,);
DFFARX1 I_68385 (I1165034,I2507,I1164754,I1164743,);
nor I_68386 (I1165096,I1299739,I1299760);
nor I_68387 (I1164734,I1164949,I1165096);
or I_68388 (I1165127,I1299739,I1299760);
nor I_68389 (I1165144,I1299748,I1299736);
DFFARX1 I_68390 (I1165144,I2507,I1164754,I1165170,);
not I_68391 (I1165178,I1165170);
nor I_68392 (I1164740,I1165178,I1164983);
nand I_68393 (I1165209,I1165178,I1164828);
not I_68394 (I1165226,I1299748);
nand I_68395 (I1165243,I1165226,I1164932);
nand I_68396 (I1165260,I1165178,I1165243);
nand I_68397 (I1164731,I1165260,I1165209);
nand I_68398 (I1164728,I1165243,I1165127);
not I_68399 (I1165332,I2514);
DFFARX1 I_68400 (I821750,I2507,I1165332,I1165358,);
and I_68401 (I1165366,I1165358,I821756);
DFFARX1 I_68402 (I1165366,I2507,I1165332,I1165315,);
DFFARX1 I_68403 (I821762,I2507,I1165332,I1165406,);
not I_68404 (I1165414,I821747);
not I_68405 (I1165431,I821747);
nand I_68406 (I1165448,I1165431,I1165414);
nor I_68407 (I1165303,I1165406,I1165448);
DFFARX1 I_68408 (I1165448,I2507,I1165332,I1165488,);
not I_68409 (I1165324,I1165488);
not I_68410 (I1165510,I821765);
nand I_68411 (I1165527,I1165431,I1165510);
DFFARX1 I_68412 (I1165527,I2507,I1165332,I1165553,);
not I_68413 (I1165561,I1165553);
not I_68414 (I1165578,I821759);
nand I_68415 (I1165595,I1165578,I821750);
and I_68416 (I1165612,I1165414,I1165595);
nor I_68417 (I1165629,I1165527,I1165612);
DFFARX1 I_68418 (I1165629,I2507,I1165332,I1165300,);
DFFARX1 I_68419 (I1165612,I2507,I1165332,I1165321,);
nor I_68420 (I1165674,I821759,I821768);
nor I_68421 (I1165312,I1165527,I1165674);
or I_68422 (I1165705,I821759,I821768);
nor I_68423 (I1165722,I821753,I821753);
DFFARX1 I_68424 (I1165722,I2507,I1165332,I1165748,);
not I_68425 (I1165756,I1165748);
nor I_68426 (I1165318,I1165756,I1165561);
nand I_68427 (I1165787,I1165756,I1165406);
not I_68428 (I1165804,I821753);
nand I_68429 (I1165821,I1165804,I1165510);
nand I_68430 (I1165838,I1165756,I1165821);
nand I_68431 (I1165309,I1165838,I1165787);
nand I_68432 (I1165306,I1165821,I1165705);
not I_68433 (I1165910,I2514);
DFFARX1 I_68434 (I420207,I2507,I1165910,I1165936,);
and I_68435 (I1165944,I1165936,I420222);
DFFARX1 I_68436 (I1165944,I2507,I1165910,I1165893,);
DFFARX1 I_68437 (I420225,I2507,I1165910,I1165984,);
not I_68438 (I1165992,I420219);
not I_68439 (I1166009,I420234);
nand I_68440 (I1166026,I1166009,I1165992);
nor I_68441 (I1165881,I1165984,I1166026);
DFFARX1 I_68442 (I1166026,I2507,I1165910,I1166066,);
not I_68443 (I1165902,I1166066);
not I_68444 (I1166088,I420210);
nand I_68445 (I1166105,I1166009,I1166088);
DFFARX1 I_68446 (I1166105,I2507,I1165910,I1166131,);
not I_68447 (I1166139,I1166131);
not I_68448 (I1166156,I420213);
nand I_68449 (I1166173,I1166156,I420207);
and I_68450 (I1166190,I1165992,I1166173);
nor I_68451 (I1166207,I1166105,I1166190);
DFFARX1 I_68452 (I1166207,I2507,I1165910,I1165878,);
DFFARX1 I_68453 (I1166190,I2507,I1165910,I1165899,);
nor I_68454 (I1166252,I420213,I420216);
nor I_68455 (I1165890,I1166105,I1166252);
or I_68456 (I1166283,I420213,I420216);
nor I_68457 (I1166300,I420231,I420228);
DFFARX1 I_68458 (I1166300,I2507,I1165910,I1166326,);
not I_68459 (I1166334,I1166326);
nor I_68460 (I1165896,I1166334,I1166139);
nand I_68461 (I1166365,I1166334,I1165984);
not I_68462 (I1166382,I420231);
nand I_68463 (I1166399,I1166382,I1166088);
nand I_68464 (I1166416,I1166334,I1166399);
nand I_68465 (I1165887,I1166416,I1166365);
nand I_68466 (I1165884,I1166399,I1166283);
not I_68467 (I1166488,I2514);
DFFARX1 I_68468 (I593741,I2507,I1166488,I1166514,);
and I_68469 (I1166522,I1166514,I593729);
DFFARX1 I_68470 (I1166522,I2507,I1166488,I1166471,);
DFFARX1 I_68471 (I593744,I2507,I1166488,I1166562,);
not I_68472 (I1166570,I593735);
not I_68473 (I1166587,I593726);
nand I_68474 (I1166604,I1166587,I1166570);
nor I_68475 (I1166459,I1166562,I1166604);
DFFARX1 I_68476 (I1166604,I2507,I1166488,I1166644,);
not I_68477 (I1166480,I1166644);
not I_68478 (I1166666,I593732);
nand I_68479 (I1166683,I1166587,I1166666);
DFFARX1 I_68480 (I1166683,I2507,I1166488,I1166709,);
not I_68481 (I1166717,I1166709);
not I_68482 (I1166734,I593747);
nand I_68483 (I1166751,I1166734,I593750);
and I_68484 (I1166768,I1166570,I1166751);
nor I_68485 (I1166785,I1166683,I1166768);
DFFARX1 I_68486 (I1166785,I2507,I1166488,I1166456,);
DFFARX1 I_68487 (I1166768,I2507,I1166488,I1166477,);
nor I_68488 (I1166830,I593747,I593726);
nor I_68489 (I1166468,I1166683,I1166830);
or I_68490 (I1166861,I593747,I593726);
nor I_68491 (I1166878,I593738,I593729);
DFFARX1 I_68492 (I1166878,I2507,I1166488,I1166904,);
not I_68493 (I1166912,I1166904);
nor I_68494 (I1166474,I1166912,I1166717);
nand I_68495 (I1166943,I1166912,I1166562);
not I_68496 (I1166960,I593738);
nand I_68497 (I1166977,I1166960,I1166666);
nand I_68498 (I1166994,I1166912,I1166977);
nand I_68499 (I1166465,I1166994,I1166943);
nand I_68500 (I1166462,I1166977,I1166861);
not I_68501 (I1167066,I2514);
DFFARX1 I_68502 (I719745,I2507,I1167066,I1167092,);
and I_68503 (I1167100,I1167092,I719733);
DFFARX1 I_68504 (I1167100,I2507,I1167066,I1167049,);
DFFARX1 I_68505 (I719736,I2507,I1167066,I1167140,);
not I_68506 (I1167148,I719730);
not I_68507 (I1167165,I719754);
nand I_68508 (I1167182,I1167165,I1167148);
nor I_68509 (I1167037,I1167140,I1167182);
DFFARX1 I_68510 (I1167182,I2507,I1167066,I1167222,);
not I_68511 (I1167058,I1167222);
not I_68512 (I1167244,I719742);
nand I_68513 (I1167261,I1167165,I1167244);
DFFARX1 I_68514 (I1167261,I2507,I1167066,I1167287,);
not I_68515 (I1167295,I1167287);
not I_68516 (I1167312,I719751);
nand I_68517 (I1167329,I1167312,I719748);
and I_68518 (I1167346,I1167148,I1167329);
nor I_68519 (I1167363,I1167261,I1167346);
DFFARX1 I_68520 (I1167363,I2507,I1167066,I1167034,);
DFFARX1 I_68521 (I1167346,I2507,I1167066,I1167055,);
nor I_68522 (I1167408,I719751,I719739);
nor I_68523 (I1167046,I1167261,I1167408);
or I_68524 (I1167439,I719751,I719739);
nor I_68525 (I1167456,I719730,I719733);
DFFARX1 I_68526 (I1167456,I2507,I1167066,I1167482,);
not I_68527 (I1167490,I1167482);
nor I_68528 (I1167052,I1167490,I1167295);
nand I_68529 (I1167521,I1167490,I1167140);
not I_68530 (I1167538,I719730);
nand I_68531 (I1167555,I1167538,I1167244);
nand I_68532 (I1167572,I1167490,I1167555);
nand I_68533 (I1167043,I1167572,I1167521);
nand I_68534 (I1167040,I1167555,I1167439);
not I_68535 (I1167644,I2514);
DFFARX1 I_68536 (I534552,I2507,I1167644,I1167670,);
and I_68537 (I1167678,I1167670,I534567);
DFFARX1 I_68538 (I1167678,I2507,I1167644,I1167627,);
DFFARX1 I_68539 (I534558,I2507,I1167644,I1167718,);
not I_68540 (I1167726,I534552);
not I_68541 (I1167743,I534570);
nand I_68542 (I1167760,I1167743,I1167726);
nor I_68543 (I1167615,I1167718,I1167760);
DFFARX1 I_68544 (I1167760,I2507,I1167644,I1167800,);
not I_68545 (I1167636,I1167800);
not I_68546 (I1167822,I534561);
nand I_68547 (I1167839,I1167743,I1167822);
DFFARX1 I_68548 (I1167839,I2507,I1167644,I1167865,);
not I_68549 (I1167873,I1167865);
not I_68550 (I1167890,I534573);
nand I_68551 (I1167907,I1167890,I534549);
and I_68552 (I1167924,I1167726,I1167907);
nor I_68553 (I1167941,I1167839,I1167924);
DFFARX1 I_68554 (I1167941,I2507,I1167644,I1167612,);
DFFARX1 I_68555 (I1167924,I2507,I1167644,I1167633,);
nor I_68556 (I1167986,I534573,I534549);
nor I_68557 (I1167624,I1167839,I1167986);
or I_68558 (I1168017,I534573,I534549);
nor I_68559 (I1168034,I534555,I534564);
DFFARX1 I_68560 (I1168034,I2507,I1167644,I1168060,);
not I_68561 (I1168068,I1168060);
nor I_68562 (I1167630,I1168068,I1167873);
nand I_68563 (I1168099,I1168068,I1167718);
not I_68564 (I1168116,I534555);
nand I_68565 (I1168133,I1168116,I1167822);
nand I_68566 (I1168150,I1168068,I1168133);
nand I_68567 (I1167621,I1168150,I1168099);
nand I_68568 (I1167618,I1168133,I1168017);
not I_68569 (I1168222,I2514);
DFFARX1 I_68570 (I277094,I2507,I1168222,I1168248,);
and I_68571 (I1168256,I1168248,I277079);
DFFARX1 I_68572 (I1168256,I2507,I1168222,I1168205,);
DFFARX1 I_68573 (I277085,I2507,I1168222,I1168296,);
not I_68574 (I1168304,I277067);
not I_68575 (I1168321,I277088);
nand I_68576 (I1168338,I1168321,I1168304);
nor I_68577 (I1168193,I1168296,I1168338);
DFFARX1 I_68578 (I1168338,I2507,I1168222,I1168378,);
not I_68579 (I1168214,I1168378);
not I_68580 (I1168400,I277091);
nand I_68581 (I1168417,I1168321,I1168400);
DFFARX1 I_68582 (I1168417,I2507,I1168222,I1168443,);
not I_68583 (I1168451,I1168443);
not I_68584 (I1168468,I277082);
nand I_68585 (I1168485,I1168468,I277070);
and I_68586 (I1168502,I1168304,I1168485);
nor I_68587 (I1168519,I1168417,I1168502);
DFFARX1 I_68588 (I1168519,I2507,I1168222,I1168190,);
DFFARX1 I_68589 (I1168502,I2507,I1168222,I1168211,);
nor I_68590 (I1168564,I277082,I277076);
nor I_68591 (I1168202,I1168417,I1168564);
or I_68592 (I1168595,I277082,I277076);
nor I_68593 (I1168612,I277073,I277067);
DFFARX1 I_68594 (I1168612,I2507,I1168222,I1168638,);
not I_68595 (I1168646,I1168638);
nor I_68596 (I1168208,I1168646,I1168451);
nand I_68597 (I1168677,I1168646,I1168296);
not I_68598 (I1168694,I277073);
nand I_68599 (I1168711,I1168694,I1168400);
nand I_68600 (I1168728,I1168646,I1168711);
nand I_68601 (I1168199,I1168728,I1168677);
nand I_68602 (I1168196,I1168711,I1168595);
not I_68603 (I1168800,I2514);
DFFARX1 I_68604 (I134988,I2507,I1168800,I1168826,);
and I_68605 (I1168834,I1168826,I134964);
DFFARX1 I_68606 (I1168834,I2507,I1168800,I1168783,);
DFFARX1 I_68607 (I134982,I2507,I1168800,I1168874,);
not I_68608 (I1168882,I134970);
not I_68609 (I1168899,I134967);
nand I_68610 (I1168916,I1168899,I1168882);
nor I_68611 (I1168771,I1168874,I1168916);
DFFARX1 I_68612 (I1168916,I2507,I1168800,I1168956,);
not I_68613 (I1168792,I1168956);
not I_68614 (I1168978,I134976);
nand I_68615 (I1168995,I1168899,I1168978);
DFFARX1 I_68616 (I1168995,I2507,I1168800,I1169021,);
not I_68617 (I1169029,I1169021);
not I_68618 (I1169046,I134967);
nand I_68619 (I1169063,I1169046,I134985);
and I_68620 (I1169080,I1168882,I1169063);
nor I_68621 (I1169097,I1168995,I1169080);
DFFARX1 I_68622 (I1169097,I2507,I1168800,I1168768,);
DFFARX1 I_68623 (I1169080,I2507,I1168800,I1168789,);
nor I_68624 (I1169142,I134967,I134979);
nor I_68625 (I1168780,I1168995,I1169142);
or I_68626 (I1169173,I134967,I134979);
nor I_68627 (I1169190,I134973,I134964);
DFFARX1 I_68628 (I1169190,I2507,I1168800,I1169216,);
not I_68629 (I1169224,I1169216);
nor I_68630 (I1168786,I1169224,I1169029);
nand I_68631 (I1169255,I1169224,I1168874);
not I_68632 (I1169272,I134973);
nand I_68633 (I1169289,I1169272,I1168978);
nand I_68634 (I1169306,I1169224,I1169289);
nand I_68635 (I1168777,I1169306,I1169255);
nand I_68636 (I1168774,I1169289,I1169173);
not I_68637 (I1169378,I2514);
DFFARX1 I_68638 (I384847,I2507,I1169378,I1169404,);
and I_68639 (I1169412,I1169404,I384862);
DFFARX1 I_68640 (I1169412,I2507,I1169378,I1169361,);
DFFARX1 I_68641 (I384865,I2507,I1169378,I1169452,);
not I_68642 (I1169460,I384859);
not I_68643 (I1169477,I384874);
nand I_68644 (I1169494,I1169477,I1169460);
nor I_68645 (I1169349,I1169452,I1169494);
DFFARX1 I_68646 (I1169494,I2507,I1169378,I1169534,);
not I_68647 (I1169370,I1169534);
not I_68648 (I1169556,I384850);
nand I_68649 (I1169573,I1169477,I1169556);
DFFARX1 I_68650 (I1169573,I2507,I1169378,I1169599,);
not I_68651 (I1169607,I1169599);
not I_68652 (I1169624,I384853);
nand I_68653 (I1169641,I1169624,I384847);
and I_68654 (I1169658,I1169460,I1169641);
nor I_68655 (I1169675,I1169573,I1169658);
DFFARX1 I_68656 (I1169675,I2507,I1169378,I1169346,);
DFFARX1 I_68657 (I1169658,I2507,I1169378,I1169367,);
nor I_68658 (I1169720,I384853,I384856);
nor I_68659 (I1169358,I1169573,I1169720);
or I_68660 (I1169751,I384853,I384856);
nor I_68661 (I1169768,I384871,I384868);
DFFARX1 I_68662 (I1169768,I2507,I1169378,I1169794,);
not I_68663 (I1169802,I1169794);
nor I_68664 (I1169364,I1169802,I1169607);
nand I_68665 (I1169833,I1169802,I1169452);
not I_68666 (I1169850,I384871);
nand I_68667 (I1169867,I1169850,I1169556);
nand I_68668 (I1169884,I1169802,I1169867);
nand I_68669 (I1169355,I1169884,I1169833);
nand I_68670 (I1169352,I1169867,I1169751);
not I_68671 (I1169956,I2514);
DFFARX1 I_68672 (I478415,I2507,I1169956,I1169982,);
and I_68673 (I1169990,I1169982,I478430);
DFFARX1 I_68674 (I1169990,I2507,I1169956,I1169939,);
DFFARX1 I_68675 (I478433,I2507,I1169956,I1170030,);
not I_68676 (I1170038,I478427);
not I_68677 (I1170055,I478442);
nand I_68678 (I1170072,I1170055,I1170038);
nor I_68679 (I1169927,I1170030,I1170072);
DFFARX1 I_68680 (I1170072,I2507,I1169956,I1170112,);
not I_68681 (I1169948,I1170112);
not I_68682 (I1170134,I478418);
nand I_68683 (I1170151,I1170055,I1170134);
DFFARX1 I_68684 (I1170151,I2507,I1169956,I1170177,);
not I_68685 (I1170185,I1170177);
not I_68686 (I1170202,I478421);
nand I_68687 (I1170219,I1170202,I478415);
and I_68688 (I1170236,I1170038,I1170219);
nor I_68689 (I1170253,I1170151,I1170236);
DFFARX1 I_68690 (I1170253,I2507,I1169956,I1169924,);
DFFARX1 I_68691 (I1170236,I2507,I1169956,I1169945,);
nor I_68692 (I1170298,I478421,I478424);
nor I_68693 (I1169936,I1170151,I1170298);
or I_68694 (I1170329,I478421,I478424);
nor I_68695 (I1170346,I478439,I478436);
DFFARX1 I_68696 (I1170346,I2507,I1169956,I1170372,);
not I_68697 (I1170380,I1170372);
nor I_68698 (I1169942,I1170380,I1170185);
nand I_68699 (I1170411,I1170380,I1170030);
not I_68700 (I1170428,I478439);
nand I_68701 (I1170445,I1170428,I1170134);
nand I_68702 (I1170462,I1170380,I1170445);
nand I_68703 (I1169933,I1170462,I1170411);
nand I_68704 (I1169930,I1170445,I1170329);
not I_68705 (I1170534,I2514);
DFFARX1 I_68706 (I659633,I2507,I1170534,I1170560,);
and I_68707 (I1170568,I1170560,I659621);
DFFARX1 I_68708 (I1170568,I2507,I1170534,I1170517,);
DFFARX1 I_68709 (I659624,I2507,I1170534,I1170608,);
not I_68710 (I1170616,I659618);
not I_68711 (I1170633,I659642);
nand I_68712 (I1170650,I1170633,I1170616);
nor I_68713 (I1170505,I1170608,I1170650);
DFFARX1 I_68714 (I1170650,I2507,I1170534,I1170690,);
not I_68715 (I1170526,I1170690);
not I_68716 (I1170712,I659630);
nand I_68717 (I1170729,I1170633,I1170712);
DFFARX1 I_68718 (I1170729,I2507,I1170534,I1170755,);
not I_68719 (I1170763,I1170755);
not I_68720 (I1170780,I659639);
nand I_68721 (I1170797,I1170780,I659636);
and I_68722 (I1170814,I1170616,I1170797);
nor I_68723 (I1170831,I1170729,I1170814);
DFFARX1 I_68724 (I1170831,I2507,I1170534,I1170502,);
DFFARX1 I_68725 (I1170814,I2507,I1170534,I1170523,);
nor I_68726 (I1170876,I659639,I659627);
nor I_68727 (I1170514,I1170729,I1170876);
or I_68728 (I1170907,I659639,I659627);
nor I_68729 (I1170924,I659618,I659621);
DFFARX1 I_68730 (I1170924,I2507,I1170534,I1170950,);
not I_68731 (I1170958,I1170950);
nor I_68732 (I1170520,I1170958,I1170763);
nand I_68733 (I1170989,I1170958,I1170608);
not I_68734 (I1171006,I659618);
nand I_68735 (I1171023,I1171006,I1170712);
nand I_68736 (I1171040,I1170958,I1171023);
nand I_68737 (I1170511,I1171040,I1170989);
nand I_68738 (I1170508,I1171023,I1170907);
not I_68739 (I1171112,I2514);
DFFARX1 I_68740 (I810683,I2507,I1171112,I1171138,);
and I_68741 (I1171146,I1171138,I810689);
DFFARX1 I_68742 (I1171146,I2507,I1171112,I1171095,);
DFFARX1 I_68743 (I810695,I2507,I1171112,I1171186,);
not I_68744 (I1171194,I810680);
not I_68745 (I1171211,I810680);
nand I_68746 (I1171228,I1171211,I1171194);
nor I_68747 (I1171083,I1171186,I1171228);
DFFARX1 I_68748 (I1171228,I2507,I1171112,I1171268,);
not I_68749 (I1171104,I1171268);
not I_68750 (I1171290,I810698);
nand I_68751 (I1171307,I1171211,I1171290);
DFFARX1 I_68752 (I1171307,I2507,I1171112,I1171333,);
not I_68753 (I1171341,I1171333);
not I_68754 (I1171358,I810692);
nand I_68755 (I1171375,I1171358,I810683);
and I_68756 (I1171392,I1171194,I1171375);
nor I_68757 (I1171409,I1171307,I1171392);
DFFARX1 I_68758 (I1171409,I2507,I1171112,I1171080,);
DFFARX1 I_68759 (I1171392,I2507,I1171112,I1171101,);
nor I_68760 (I1171454,I810692,I810701);
nor I_68761 (I1171092,I1171307,I1171454);
or I_68762 (I1171485,I810692,I810701);
nor I_68763 (I1171502,I810686,I810686);
DFFARX1 I_68764 (I1171502,I2507,I1171112,I1171528,);
not I_68765 (I1171536,I1171528);
nor I_68766 (I1171098,I1171536,I1171341);
nand I_68767 (I1171567,I1171536,I1171186);
not I_68768 (I1171584,I810686);
nand I_68769 (I1171601,I1171584,I1171290);
nand I_68770 (I1171618,I1171536,I1171601);
nand I_68771 (I1171089,I1171618,I1171567);
nand I_68772 (I1171086,I1171601,I1171485);
not I_68773 (I1171690,I2514);
DFFARX1 I_68774 (I730727,I2507,I1171690,I1171716,);
and I_68775 (I1171724,I1171716,I730715);
DFFARX1 I_68776 (I1171724,I2507,I1171690,I1171673,);
DFFARX1 I_68777 (I730718,I2507,I1171690,I1171764,);
not I_68778 (I1171772,I730712);
not I_68779 (I1171789,I730736);
nand I_68780 (I1171806,I1171789,I1171772);
nor I_68781 (I1171661,I1171764,I1171806);
DFFARX1 I_68782 (I1171806,I2507,I1171690,I1171846,);
not I_68783 (I1171682,I1171846);
not I_68784 (I1171868,I730724);
nand I_68785 (I1171885,I1171789,I1171868);
DFFARX1 I_68786 (I1171885,I2507,I1171690,I1171911,);
not I_68787 (I1171919,I1171911);
not I_68788 (I1171936,I730733);
nand I_68789 (I1171953,I1171936,I730730);
and I_68790 (I1171970,I1171772,I1171953);
nor I_68791 (I1171987,I1171885,I1171970);
DFFARX1 I_68792 (I1171987,I2507,I1171690,I1171658,);
DFFARX1 I_68793 (I1171970,I2507,I1171690,I1171679,);
nor I_68794 (I1172032,I730733,I730721);
nor I_68795 (I1171670,I1171885,I1172032);
or I_68796 (I1172063,I730733,I730721);
nor I_68797 (I1172080,I730712,I730715);
DFFARX1 I_68798 (I1172080,I2507,I1171690,I1172106,);
not I_68799 (I1172114,I1172106);
nor I_68800 (I1171676,I1172114,I1171919);
nand I_68801 (I1172145,I1172114,I1171764);
not I_68802 (I1172162,I730712);
nand I_68803 (I1172179,I1172162,I1171868);
nand I_68804 (I1172196,I1172114,I1172179);
nand I_68805 (I1171667,I1172196,I1172145);
nand I_68806 (I1171664,I1172179,I1172063);
not I_68807 (I1172268,I2514);
DFFARX1 I_68808 (I1344014,I2507,I1172268,I1172294,);
and I_68809 (I1172302,I1172294,I1343996);
DFFARX1 I_68810 (I1172302,I2507,I1172268,I1172251,);
DFFARX1 I_68811 (I1343987,I2507,I1172268,I1172342,);
not I_68812 (I1172350,I1344002);
not I_68813 (I1172367,I1343990);
nand I_68814 (I1172384,I1172367,I1172350);
nor I_68815 (I1172239,I1172342,I1172384);
DFFARX1 I_68816 (I1172384,I2507,I1172268,I1172424,);
not I_68817 (I1172260,I1172424);
not I_68818 (I1172446,I1343999);
nand I_68819 (I1172463,I1172367,I1172446);
DFFARX1 I_68820 (I1172463,I2507,I1172268,I1172489,);
not I_68821 (I1172497,I1172489);
not I_68822 (I1172514,I1344008);
nand I_68823 (I1172531,I1172514,I1343987);
and I_68824 (I1172548,I1172350,I1172531);
nor I_68825 (I1172565,I1172463,I1172548);
DFFARX1 I_68826 (I1172565,I2507,I1172268,I1172236,);
DFFARX1 I_68827 (I1172548,I2507,I1172268,I1172257,);
nor I_68828 (I1172610,I1344008,I1344011);
nor I_68829 (I1172248,I1172463,I1172610);
or I_68830 (I1172641,I1344008,I1344011);
nor I_68831 (I1172658,I1344005,I1343993);
DFFARX1 I_68832 (I1172658,I2507,I1172268,I1172684,);
not I_68833 (I1172692,I1172684);
nor I_68834 (I1172254,I1172692,I1172497);
nand I_68835 (I1172723,I1172692,I1172342);
not I_68836 (I1172740,I1344005);
nand I_68837 (I1172757,I1172740,I1172446);
nand I_68838 (I1172774,I1172692,I1172757);
nand I_68839 (I1172245,I1172774,I1172723);
nand I_68840 (I1172242,I1172757,I1172641);
not I_68841 (I1172846,I2514);
DFFARX1 I_68842 (I240075,I2507,I1172846,I1172872,);
and I_68843 (I1172880,I1172872,I240078);
DFFARX1 I_68844 (I1172880,I2507,I1172846,I1172829,);
DFFARX1 I_68845 (I240078,I2507,I1172846,I1172920,);
not I_68846 (I1172928,I240093);
not I_68847 (I1172945,I240099);
nand I_68848 (I1172962,I1172945,I1172928);
nor I_68849 (I1172817,I1172920,I1172962);
DFFARX1 I_68850 (I1172962,I2507,I1172846,I1173002,);
not I_68851 (I1172838,I1173002);
not I_68852 (I1173024,I240087);
nand I_68853 (I1173041,I1172945,I1173024);
DFFARX1 I_68854 (I1173041,I2507,I1172846,I1173067,);
not I_68855 (I1173075,I1173067);
not I_68856 (I1173092,I240084);
nand I_68857 (I1173109,I1173092,I240081);
and I_68858 (I1173126,I1172928,I1173109);
nor I_68859 (I1173143,I1173041,I1173126);
DFFARX1 I_68860 (I1173143,I2507,I1172846,I1172814,);
DFFARX1 I_68861 (I1173126,I2507,I1172846,I1172835,);
nor I_68862 (I1173188,I240084,I240075);
nor I_68863 (I1172826,I1173041,I1173188);
or I_68864 (I1173219,I240084,I240075);
nor I_68865 (I1173236,I240090,I240096);
DFFARX1 I_68866 (I1173236,I2507,I1172846,I1173262,);
not I_68867 (I1173270,I1173262);
nor I_68868 (I1172832,I1173270,I1173075);
nand I_68869 (I1173301,I1173270,I1172920);
not I_68870 (I1173318,I240090);
nand I_68871 (I1173335,I1173318,I1173024);
nand I_68872 (I1173352,I1173270,I1173335);
nand I_68873 (I1172823,I1173352,I1173301);
nand I_68874 (I1172820,I1173335,I1173219);
not I_68875 (I1173424,I2514);
DFFARX1 I_68876 (I694313,I2507,I1173424,I1173450,);
and I_68877 (I1173458,I1173450,I694301);
DFFARX1 I_68878 (I1173458,I2507,I1173424,I1173407,);
DFFARX1 I_68879 (I694304,I2507,I1173424,I1173498,);
not I_68880 (I1173506,I694298);
not I_68881 (I1173523,I694322);
nand I_68882 (I1173540,I1173523,I1173506);
nor I_68883 (I1173395,I1173498,I1173540);
DFFARX1 I_68884 (I1173540,I2507,I1173424,I1173580,);
not I_68885 (I1173416,I1173580);
not I_68886 (I1173602,I694310);
nand I_68887 (I1173619,I1173523,I1173602);
DFFARX1 I_68888 (I1173619,I2507,I1173424,I1173645,);
not I_68889 (I1173653,I1173645);
not I_68890 (I1173670,I694319);
nand I_68891 (I1173687,I1173670,I694316);
and I_68892 (I1173704,I1173506,I1173687);
nor I_68893 (I1173721,I1173619,I1173704);
DFFARX1 I_68894 (I1173721,I2507,I1173424,I1173392,);
DFFARX1 I_68895 (I1173704,I2507,I1173424,I1173413,);
nor I_68896 (I1173766,I694319,I694307);
nor I_68897 (I1173404,I1173619,I1173766);
or I_68898 (I1173797,I694319,I694307);
nor I_68899 (I1173814,I694298,I694301);
DFFARX1 I_68900 (I1173814,I2507,I1173424,I1173840,);
not I_68901 (I1173848,I1173840);
nor I_68902 (I1173410,I1173848,I1173653);
nand I_68903 (I1173879,I1173848,I1173498);
not I_68904 (I1173896,I694298);
nand I_68905 (I1173913,I1173896,I1173602);
nand I_68906 (I1173930,I1173848,I1173913);
nand I_68907 (I1173401,I1173930,I1173879);
nand I_68908 (I1173398,I1173913,I1173797);
not I_68909 (I1174002,I2514);
DFFARX1 I_68910 (I572355,I2507,I1174002,I1174028,);
and I_68911 (I1174036,I1174028,I572343);
DFFARX1 I_68912 (I1174036,I2507,I1174002,I1173985,);
DFFARX1 I_68913 (I572358,I2507,I1174002,I1174076,);
not I_68914 (I1174084,I572349);
not I_68915 (I1174101,I572340);
nand I_68916 (I1174118,I1174101,I1174084);
nor I_68917 (I1173973,I1174076,I1174118);
DFFARX1 I_68918 (I1174118,I2507,I1174002,I1174158,);
not I_68919 (I1173994,I1174158);
not I_68920 (I1174180,I572346);
nand I_68921 (I1174197,I1174101,I1174180);
DFFARX1 I_68922 (I1174197,I2507,I1174002,I1174223,);
not I_68923 (I1174231,I1174223);
not I_68924 (I1174248,I572361);
nand I_68925 (I1174265,I1174248,I572364);
and I_68926 (I1174282,I1174084,I1174265);
nor I_68927 (I1174299,I1174197,I1174282);
DFFARX1 I_68928 (I1174299,I2507,I1174002,I1173970,);
DFFARX1 I_68929 (I1174282,I2507,I1174002,I1173991,);
nor I_68930 (I1174344,I572361,I572340);
nor I_68931 (I1173982,I1174197,I1174344);
or I_68932 (I1174375,I572361,I572340);
nor I_68933 (I1174392,I572352,I572343);
DFFARX1 I_68934 (I1174392,I2507,I1174002,I1174418,);
not I_68935 (I1174426,I1174418);
nor I_68936 (I1173988,I1174426,I1174231);
nand I_68937 (I1174457,I1174426,I1174076);
not I_68938 (I1174474,I572352);
nand I_68939 (I1174491,I1174474,I1174180);
nand I_68940 (I1174508,I1174426,I1174491);
nand I_68941 (I1173979,I1174508,I1174457);
nand I_68942 (I1173976,I1174491,I1174375);
not I_68943 (I1174580,I2514);
DFFARX1 I_68944 (I1252055,I2507,I1174580,I1174606,);
and I_68945 (I1174614,I1174606,I1252049);
DFFARX1 I_68946 (I1174614,I2507,I1174580,I1174563,);
DFFARX1 I_68947 (I1252034,I2507,I1174580,I1174654,);
not I_68948 (I1174662,I1252040);
not I_68949 (I1174679,I1252052);
nand I_68950 (I1174696,I1174679,I1174662);
nor I_68951 (I1174551,I1174654,I1174696);
DFFARX1 I_68952 (I1174696,I2507,I1174580,I1174736,);
not I_68953 (I1174572,I1174736);
not I_68954 (I1174758,I1252034);
nand I_68955 (I1174775,I1174679,I1174758);
DFFARX1 I_68956 (I1174775,I2507,I1174580,I1174801,);
not I_68957 (I1174809,I1174801);
not I_68958 (I1174826,I1252058);
nand I_68959 (I1174843,I1174826,I1252046);
and I_68960 (I1174860,I1174662,I1174843);
nor I_68961 (I1174877,I1174775,I1174860);
DFFARX1 I_68962 (I1174877,I2507,I1174580,I1174548,);
DFFARX1 I_68963 (I1174860,I2507,I1174580,I1174569,);
nor I_68964 (I1174922,I1252058,I1252037);
nor I_68965 (I1174560,I1174775,I1174922);
or I_68966 (I1174953,I1252058,I1252037);
nor I_68967 (I1174970,I1252043,I1252037);
DFFARX1 I_68968 (I1174970,I2507,I1174580,I1174996,);
not I_68969 (I1175004,I1174996);
nor I_68970 (I1174566,I1175004,I1174809);
nand I_68971 (I1175035,I1175004,I1174654);
not I_68972 (I1175052,I1252043);
nand I_68973 (I1175069,I1175052,I1174758);
nand I_68974 (I1175086,I1175004,I1175069);
nand I_68975 (I1174557,I1175086,I1175035);
nand I_68976 (I1174554,I1175069,I1174953);
not I_68977 (I1175158,I2514);
DFFARX1 I_68978 (I477327,I2507,I1175158,I1175184,);
and I_68979 (I1175192,I1175184,I477342);
DFFARX1 I_68980 (I1175192,I2507,I1175158,I1175141,);
DFFARX1 I_68981 (I477345,I2507,I1175158,I1175232,);
not I_68982 (I1175240,I477339);
not I_68983 (I1175257,I477354);
nand I_68984 (I1175274,I1175257,I1175240);
nor I_68985 (I1175129,I1175232,I1175274);
DFFARX1 I_68986 (I1175274,I2507,I1175158,I1175314,);
not I_68987 (I1175150,I1175314);
not I_68988 (I1175336,I477330);
nand I_68989 (I1175353,I1175257,I1175336);
DFFARX1 I_68990 (I1175353,I2507,I1175158,I1175379,);
not I_68991 (I1175387,I1175379);
not I_68992 (I1175404,I477333);
nand I_68993 (I1175421,I1175404,I477327);
and I_68994 (I1175438,I1175240,I1175421);
nor I_68995 (I1175455,I1175353,I1175438);
DFFARX1 I_68996 (I1175455,I2507,I1175158,I1175126,);
DFFARX1 I_68997 (I1175438,I2507,I1175158,I1175147,);
nor I_68998 (I1175500,I477333,I477336);
nor I_68999 (I1175138,I1175353,I1175500);
or I_69000 (I1175531,I477333,I477336);
nor I_69001 (I1175548,I477351,I477348);
DFFARX1 I_69002 (I1175548,I2507,I1175158,I1175574,);
not I_69003 (I1175582,I1175574);
nor I_69004 (I1175144,I1175582,I1175387);
nand I_69005 (I1175613,I1175582,I1175232);
not I_69006 (I1175630,I477351);
nand I_69007 (I1175647,I1175630,I1175336);
nand I_69008 (I1175664,I1175582,I1175647);
nand I_69009 (I1175135,I1175664,I1175613);
nand I_69010 (I1175132,I1175647,I1175531);
not I_69011 (I1175736,I2514);
DFFARX1 I_69012 (I1025852,I2507,I1175736,I1175762,);
and I_69013 (I1175770,I1175762,I1025849);
DFFARX1 I_69014 (I1175770,I2507,I1175736,I1175719,);
DFFARX1 I_69015 (I1025855,I2507,I1175736,I1175810,);
not I_69016 (I1175818,I1025858);
not I_69017 (I1175835,I1025852);
nand I_69018 (I1175852,I1175835,I1175818);
nor I_69019 (I1175707,I1175810,I1175852);
DFFARX1 I_69020 (I1175852,I2507,I1175736,I1175892,);
not I_69021 (I1175728,I1175892);
not I_69022 (I1175914,I1025867);
nand I_69023 (I1175931,I1175835,I1175914);
DFFARX1 I_69024 (I1175931,I2507,I1175736,I1175957,);
not I_69025 (I1175965,I1175957);
not I_69026 (I1175982,I1025864);
nand I_69027 (I1175999,I1175982,I1025870);
and I_69028 (I1176016,I1175818,I1175999);
nor I_69029 (I1176033,I1175931,I1176016);
DFFARX1 I_69030 (I1176033,I2507,I1175736,I1175704,);
DFFARX1 I_69031 (I1176016,I2507,I1175736,I1175725,);
nor I_69032 (I1176078,I1025864,I1025849);
nor I_69033 (I1175716,I1175931,I1176078);
or I_69034 (I1176109,I1025864,I1025849);
nor I_69035 (I1176126,I1025861,I1025855);
DFFARX1 I_69036 (I1176126,I2507,I1175736,I1176152,);
not I_69037 (I1176160,I1176152);
nor I_69038 (I1175722,I1176160,I1175965);
nand I_69039 (I1176191,I1176160,I1175810);
not I_69040 (I1176208,I1025861);
nand I_69041 (I1176225,I1176208,I1175914);
nand I_69042 (I1176242,I1176160,I1176225);
nand I_69043 (I1175713,I1176242,I1176191);
nand I_69044 (I1175710,I1176225,I1176109);
not I_69045 (I1176314,I2514);
DFFARX1 I_69046 (I700093,I2507,I1176314,I1176340,);
and I_69047 (I1176348,I1176340,I700081);
DFFARX1 I_69048 (I1176348,I2507,I1176314,I1176297,);
DFFARX1 I_69049 (I700084,I2507,I1176314,I1176388,);
not I_69050 (I1176396,I700078);
not I_69051 (I1176413,I700102);
nand I_69052 (I1176430,I1176413,I1176396);
nor I_69053 (I1176285,I1176388,I1176430);
DFFARX1 I_69054 (I1176430,I2507,I1176314,I1176470,);
not I_69055 (I1176306,I1176470);
not I_69056 (I1176492,I700090);
nand I_69057 (I1176509,I1176413,I1176492);
DFFARX1 I_69058 (I1176509,I2507,I1176314,I1176535,);
not I_69059 (I1176543,I1176535);
not I_69060 (I1176560,I700099);
nand I_69061 (I1176577,I1176560,I700096);
and I_69062 (I1176594,I1176396,I1176577);
nor I_69063 (I1176611,I1176509,I1176594);
DFFARX1 I_69064 (I1176611,I2507,I1176314,I1176282,);
DFFARX1 I_69065 (I1176594,I2507,I1176314,I1176303,);
nor I_69066 (I1176656,I700099,I700087);
nor I_69067 (I1176294,I1176509,I1176656);
or I_69068 (I1176687,I700099,I700087);
nor I_69069 (I1176704,I700078,I700081);
DFFARX1 I_69070 (I1176704,I2507,I1176314,I1176730,);
not I_69071 (I1176738,I1176730);
nor I_69072 (I1176300,I1176738,I1176543);
nand I_69073 (I1176769,I1176738,I1176388);
not I_69074 (I1176786,I700078);
nand I_69075 (I1176803,I1176786,I1176492);
nand I_69076 (I1176820,I1176738,I1176803);
nand I_69077 (I1176291,I1176820,I1176769);
nand I_69078 (I1176288,I1176803,I1176687);
not I_69079 (I1176892,I2514);
DFFARX1 I_69080 (I1011266,I2507,I1176892,I1176918,);
and I_69081 (I1176926,I1176918,I1011263);
DFFARX1 I_69082 (I1176926,I2507,I1176892,I1176875,);
DFFARX1 I_69083 (I1011269,I2507,I1176892,I1176966,);
not I_69084 (I1176974,I1011272);
not I_69085 (I1176991,I1011266);
nand I_69086 (I1177008,I1176991,I1176974);
nor I_69087 (I1176863,I1176966,I1177008);
DFFARX1 I_69088 (I1177008,I2507,I1176892,I1177048,);
not I_69089 (I1176884,I1177048);
not I_69090 (I1177070,I1011281);
nand I_69091 (I1177087,I1176991,I1177070);
DFFARX1 I_69092 (I1177087,I2507,I1176892,I1177113,);
not I_69093 (I1177121,I1177113);
not I_69094 (I1177138,I1011278);
nand I_69095 (I1177155,I1177138,I1011284);
and I_69096 (I1177172,I1176974,I1177155);
nor I_69097 (I1177189,I1177087,I1177172);
DFFARX1 I_69098 (I1177189,I2507,I1176892,I1176860,);
DFFARX1 I_69099 (I1177172,I2507,I1176892,I1176881,);
nor I_69100 (I1177234,I1011278,I1011263);
nor I_69101 (I1176872,I1177087,I1177234);
or I_69102 (I1177265,I1011278,I1011263);
nor I_69103 (I1177282,I1011275,I1011269);
DFFARX1 I_69104 (I1177282,I2507,I1176892,I1177308,);
not I_69105 (I1177316,I1177308);
nor I_69106 (I1176878,I1177316,I1177121);
nand I_69107 (I1177347,I1177316,I1176966);
not I_69108 (I1177364,I1011275);
nand I_69109 (I1177381,I1177364,I1177070);
nand I_69110 (I1177398,I1177316,I1177381);
nand I_69111 (I1176869,I1177398,I1177347);
nand I_69112 (I1176866,I1177381,I1177265);
not I_69113 (I1177470,I2514);
DFFARX1 I_69114 (I506587,I2507,I1177470,I1177496,);
and I_69115 (I1177504,I1177496,I506602);
DFFARX1 I_69116 (I1177504,I2507,I1177470,I1177453,);
DFFARX1 I_69117 (I506593,I2507,I1177470,I1177544,);
not I_69118 (I1177552,I506587);
not I_69119 (I1177569,I506605);
nand I_69120 (I1177586,I1177569,I1177552);
nor I_69121 (I1177441,I1177544,I1177586);
DFFARX1 I_69122 (I1177586,I2507,I1177470,I1177626,);
not I_69123 (I1177462,I1177626);
not I_69124 (I1177648,I506596);
nand I_69125 (I1177665,I1177569,I1177648);
DFFARX1 I_69126 (I1177665,I2507,I1177470,I1177691,);
not I_69127 (I1177699,I1177691);
not I_69128 (I1177716,I506608);
nand I_69129 (I1177733,I1177716,I506584);
and I_69130 (I1177750,I1177552,I1177733);
nor I_69131 (I1177767,I1177665,I1177750);
DFFARX1 I_69132 (I1177767,I2507,I1177470,I1177438,);
DFFARX1 I_69133 (I1177750,I2507,I1177470,I1177459,);
nor I_69134 (I1177812,I506608,I506584);
nor I_69135 (I1177450,I1177665,I1177812);
or I_69136 (I1177843,I506608,I506584);
nor I_69137 (I1177860,I506590,I506599);
DFFARX1 I_69138 (I1177860,I2507,I1177470,I1177886,);
not I_69139 (I1177894,I1177886);
nor I_69140 (I1177456,I1177894,I1177699);
nand I_69141 (I1177925,I1177894,I1177544);
not I_69142 (I1177942,I506590);
nand I_69143 (I1177959,I1177942,I1177648);
nand I_69144 (I1177976,I1177894,I1177959);
nand I_69145 (I1177447,I1177976,I1177925);
nand I_69146 (I1177444,I1177959,I1177843);
not I_69147 (I1178048,I2514);
DFFARX1 I_69148 (I1012388,I2507,I1178048,I1178074,);
and I_69149 (I1178082,I1178074,I1012385);
DFFARX1 I_69150 (I1178082,I2507,I1178048,I1178031,);
DFFARX1 I_69151 (I1012391,I2507,I1178048,I1178122,);
not I_69152 (I1178130,I1012394);
not I_69153 (I1178147,I1012388);
nand I_69154 (I1178164,I1178147,I1178130);
nor I_69155 (I1178019,I1178122,I1178164);
DFFARX1 I_69156 (I1178164,I2507,I1178048,I1178204,);
not I_69157 (I1178040,I1178204);
not I_69158 (I1178226,I1012403);
nand I_69159 (I1178243,I1178147,I1178226);
DFFARX1 I_69160 (I1178243,I2507,I1178048,I1178269,);
not I_69161 (I1178277,I1178269);
not I_69162 (I1178294,I1012400);
nand I_69163 (I1178311,I1178294,I1012406);
and I_69164 (I1178328,I1178130,I1178311);
nor I_69165 (I1178345,I1178243,I1178328);
DFFARX1 I_69166 (I1178345,I2507,I1178048,I1178016,);
DFFARX1 I_69167 (I1178328,I2507,I1178048,I1178037,);
nor I_69168 (I1178390,I1012400,I1012385);
nor I_69169 (I1178028,I1178243,I1178390);
or I_69170 (I1178421,I1012400,I1012385);
nor I_69171 (I1178438,I1012397,I1012391);
DFFARX1 I_69172 (I1178438,I2507,I1178048,I1178464,);
not I_69173 (I1178472,I1178464);
nor I_69174 (I1178034,I1178472,I1178277);
nand I_69175 (I1178503,I1178472,I1178122);
not I_69176 (I1178520,I1012397);
nand I_69177 (I1178537,I1178520,I1178226);
nand I_69178 (I1178554,I1178472,I1178537);
nand I_69179 (I1178025,I1178554,I1178503);
nand I_69180 (I1178022,I1178537,I1178421);
not I_69181 (I1178626,I2514);
DFFARX1 I_69182 (I550391,I2507,I1178626,I1178652,);
and I_69183 (I1178660,I1178652,I550379);
DFFARX1 I_69184 (I1178660,I2507,I1178626,I1178609,);
DFFARX1 I_69185 (I550394,I2507,I1178626,I1178700,);
not I_69186 (I1178708,I550385);
not I_69187 (I1178725,I550376);
nand I_69188 (I1178742,I1178725,I1178708);
nor I_69189 (I1178597,I1178700,I1178742);
DFFARX1 I_69190 (I1178742,I2507,I1178626,I1178782,);
not I_69191 (I1178618,I1178782);
not I_69192 (I1178804,I550382);
nand I_69193 (I1178821,I1178725,I1178804);
DFFARX1 I_69194 (I1178821,I2507,I1178626,I1178847,);
not I_69195 (I1178855,I1178847);
not I_69196 (I1178872,I550397);
nand I_69197 (I1178889,I1178872,I550400);
and I_69198 (I1178906,I1178708,I1178889);
nor I_69199 (I1178923,I1178821,I1178906);
DFFARX1 I_69200 (I1178923,I2507,I1178626,I1178594,);
DFFARX1 I_69201 (I1178906,I2507,I1178626,I1178615,);
nor I_69202 (I1178968,I550397,I550376);
nor I_69203 (I1178606,I1178821,I1178968);
or I_69204 (I1178999,I550397,I550376);
nor I_69205 (I1179016,I550388,I550379);
DFFARX1 I_69206 (I1179016,I2507,I1178626,I1179042,);
not I_69207 (I1179050,I1179042);
nor I_69208 (I1178612,I1179050,I1178855);
nand I_69209 (I1179081,I1179050,I1178700);
not I_69210 (I1179098,I550388);
nand I_69211 (I1179115,I1179098,I1178804);
nand I_69212 (I1179132,I1179050,I1179115);
nand I_69213 (I1178603,I1179132,I1179081);
nand I_69214 (I1178600,I1179115,I1178999);
not I_69215 (I1179204,I2514);
DFFARX1 I_69216 (I742287,I2507,I1179204,I1179230,);
and I_69217 (I1179238,I1179230,I742275);
DFFARX1 I_69218 (I1179238,I2507,I1179204,I1179187,);
DFFARX1 I_69219 (I742278,I2507,I1179204,I1179278,);
not I_69220 (I1179286,I742272);
not I_69221 (I1179303,I742296);
nand I_69222 (I1179320,I1179303,I1179286);
nor I_69223 (I1179175,I1179278,I1179320);
DFFARX1 I_69224 (I1179320,I2507,I1179204,I1179360,);
not I_69225 (I1179196,I1179360);
not I_69226 (I1179382,I742284);
nand I_69227 (I1179399,I1179303,I1179382);
DFFARX1 I_69228 (I1179399,I2507,I1179204,I1179425,);
not I_69229 (I1179433,I1179425);
not I_69230 (I1179450,I742293);
nand I_69231 (I1179467,I1179450,I742290);
and I_69232 (I1179484,I1179286,I1179467);
nor I_69233 (I1179501,I1179399,I1179484);
DFFARX1 I_69234 (I1179501,I2507,I1179204,I1179172,);
DFFARX1 I_69235 (I1179484,I2507,I1179204,I1179193,);
nor I_69236 (I1179546,I742293,I742281);
nor I_69237 (I1179184,I1179399,I1179546);
or I_69238 (I1179577,I742293,I742281);
nor I_69239 (I1179594,I742272,I742275);
DFFARX1 I_69240 (I1179594,I2507,I1179204,I1179620,);
not I_69241 (I1179628,I1179620);
nor I_69242 (I1179190,I1179628,I1179433);
nand I_69243 (I1179659,I1179628,I1179278);
not I_69244 (I1179676,I742272);
nand I_69245 (I1179693,I1179676,I1179382);
nand I_69246 (I1179710,I1179628,I1179693);
nand I_69247 (I1179181,I1179710,I1179659);
nand I_69248 (I1179178,I1179693,I1179577);
not I_69249 (I1179782,I2514);
DFFARX1 I_69250 (I988353,I2507,I1179782,I1179808,);
and I_69251 (I1179816,I1179808,I988347);
DFFARX1 I_69252 (I1179816,I2507,I1179782,I1179765,);
DFFARX1 I_69253 (I988365,I2507,I1179782,I1179856,);
not I_69254 (I1179864,I988356);
not I_69255 (I1179881,I988368);
nand I_69256 (I1179898,I1179881,I1179864);
nor I_69257 (I1179753,I1179856,I1179898);
DFFARX1 I_69258 (I1179898,I2507,I1179782,I1179938,);
not I_69259 (I1179774,I1179938);
not I_69260 (I1179960,I988374);
nand I_69261 (I1179977,I1179881,I1179960);
DFFARX1 I_69262 (I1179977,I2507,I1179782,I1180003,);
not I_69263 (I1180011,I1180003);
not I_69264 (I1180028,I988350);
nand I_69265 (I1180045,I1180028,I988371);
and I_69266 (I1180062,I1179864,I1180045);
nor I_69267 (I1180079,I1179977,I1180062);
DFFARX1 I_69268 (I1180079,I2507,I1179782,I1179750,);
DFFARX1 I_69269 (I1180062,I2507,I1179782,I1179771,);
nor I_69270 (I1180124,I988350,I988362);
nor I_69271 (I1179762,I1179977,I1180124);
or I_69272 (I1180155,I988350,I988362);
nor I_69273 (I1180172,I988347,I988359);
DFFARX1 I_69274 (I1180172,I2507,I1179782,I1180198,);
not I_69275 (I1180206,I1180198);
nor I_69276 (I1179768,I1180206,I1180011);
nand I_69277 (I1180237,I1180206,I1179856);
not I_69278 (I1180254,I988347);
nand I_69279 (I1180271,I1180254,I1179960);
nand I_69280 (I1180288,I1180206,I1180271);
nand I_69281 (I1179759,I1180288,I1180237);
nand I_69282 (I1179756,I1180271,I1180155);
not I_69283 (I1180360,I2514);
DFFARX1 I_69284 (I882355,I2507,I1180360,I1180386,);
and I_69285 (I1180394,I1180386,I882361);
DFFARX1 I_69286 (I1180394,I2507,I1180360,I1180343,);
DFFARX1 I_69287 (I882367,I2507,I1180360,I1180434,);
not I_69288 (I1180442,I882352);
not I_69289 (I1180459,I882352);
nand I_69290 (I1180476,I1180459,I1180442);
nor I_69291 (I1180331,I1180434,I1180476);
DFFARX1 I_69292 (I1180476,I2507,I1180360,I1180516,);
not I_69293 (I1180352,I1180516);
not I_69294 (I1180538,I882370);
nand I_69295 (I1180555,I1180459,I1180538);
DFFARX1 I_69296 (I1180555,I2507,I1180360,I1180581,);
not I_69297 (I1180589,I1180581);
not I_69298 (I1180606,I882364);
nand I_69299 (I1180623,I1180606,I882355);
and I_69300 (I1180640,I1180442,I1180623);
nor I_69301 (I1180657,I1180555,I1180640);
DFFARX1 I_69302 (I1180657,I2507,I1180360,I1180328,);
DFFARX1 I_69303 (I1180640,I2507,I1180360,I1180349,);
nor I_69304 (I1180702,I882364,I882373);
nor I_69305 (I1180340,I1180555,I1180702);
or I_69306 (I1180733,I882364,I882373);
nor I_69307 (I1180750,I882358,I882358);
DFFARX1 I_69308 (I1180750,I2507,I1180360,I1180776,);
not I_69309 (I1180784,I1180776);
nor I_69310 (I1180346,I1180784,I1180589);
nand I_69311 (I1180815,I1180784,I1180434);
not I_69312 (I1180832,I882358);
nand I_69313 (I1180849,I1180832,I1180538);
nand I_69314 (I1180866,I1180784,I1180849);
nand I_69315 (I1180337,I1180866,I1180815);
nand I_69316 (I1180334,I1180849,I1180733);
not I_69317 (I1180938,I2514);
DFFARX1 I_69318 (I3722,I2507,I1180938,I1180964,);
and I_69319 (I1180972,I1180964,I3728);
DFFARX1 I_69320 (I1180972,I2507,I1180938,I1180921,);
DFFARX1 I_69321 (I3707,I2507,I1180938,I1181012,);
not I_69322 (I1181020,I3713);
not I_69323 (I1181037,I3719);
nand I_69324 (I1181054,I1181037,I1181020);
nor I_69325 (I1180909,I1181012,I1181054);
DFFARX1 I_69326 (I1181054,I2507,I1180938,I1181094,);
not I_69327 (I1180930,I1181094);
not I_69328 (I1181116,I3710);
nand I_69329 (I1181133,I1181037,I1181116);
DFFARX1 I_69330 (I1181133,I2507,I1180938,I1181159,);
not I_69331 (I1181167,I1181159);
not I_69332 (I1181184,I3725);
nand I_69333 (I1181201,I1181184,I3710);
and I_69334 (I1181218,I1181020,I1181201);
nor I_69335 (I1181235,I1181133,I1181218);
DFFARX1 I_69336 (I1181235,I2507,I1180938,I1180906,);
DFFARX1 I_69337 (I1181218,I2507,I1180938,I1180927,);
nor I_69338 (I1181280,I3725,I3713);
nor I_69339 (I1180918,I1181133,I1181280);
or I_69340 (I1181311,I3725,I3713);
nor I_69341 (I1181328,I3716,I3707);
DFFARX1 I_69342 (I1181328,I2507,I1180938,I1181354,);
not I_69343 (I1181362,I1181354);
nor I_69344 (I1180924,I1181362,I1181167);
nand I_69345 (I1181393,I1181362,I1181012);
not I_69346 (I1181410,I3716);
nand I_69347 (I1181427,I1181410,I1181116);
nand I_69348 (I1181444,I1181362,I1181427);
nand I_69349 (I1180915,I1181444,I1181393);
nand I_69350 (I1180912,I1181427,I1181311);
not I_69351 (I1181516,I2514);
DFFARX1 I_69352 (I821223,I2507,I1181516,I1181542,);
and I_69353 (I1181550,I1181542,I821229);
DFFARX1 I_69354 (I1181550,I2507,I1181516,I1181499,);
DFFARX1 I_69355 (I821235,I2507,I1181516,I1181590,);
not I_69356 (I1181598,I821220);
not I_69357 (I1181615,I821220);
nand I_69358 (I1181632,I1181615,I1181598);
nor I_69359 (I1181487,I1181590,I1181632);
DFFARX1 I_69360 (I1181632,I2507,I1181516,I1181672,);
not I_69361 (I1181508,I1181672);
not I_69362 (I1181694,I821238);
nand I_69363 (I1181711,I1181615,I1181694);
DFFARX1 I_69364 (I1181711,I2507,I1181516,I1181737,);
not I_69365 (I1181745,I1181737);
not I_69366 (I1181762,I821232);
nand I_69367 (I1181779,I1181762,I821223);
and I_69368 (I1181796,I1181598,I1181779);
nor I_69369 (I1181813,I1181711,I1181796);
DFFARX1 I_69370 (I1181813,I2507,I1181516,I1181484,);
DFFARX1 I_69371 (I1181796,I2507,I1181516,I1181505,);
nor I_69372 (I1181858,I821232,I821241);
nor I_69373 (I1181496,I1181711,I1181858);
or I_69374 (I1181889,I821232,I821241);
nor I_69375 (I1181906,I821226,I821226);
DFFARX1 I_69376 (I1181906,I2507,I1181516,I1181932,);
not I_69377 (I1181940,I1181932);
nor I_69378 (I1181502,I1181940,I1181745);
nand I_69379 (I1181971,I1181940,I1181590);
not I_69380 (I1181988,I821226);
nand I_69381 (I1182005,I1181988,I1181694);
nand I_69382 (I1182022,I1181940,I1182005);
nand I_69383 (I1181493,I1182022,I1181971);
nand I_69384 (I1181490,I1182005,I1181889);
not I_69385 (I1182094,I2514);
DFFARX1 I_69386 (I989645,I2507,I1182094,I1182120,);
and I_69387 (I1182128,I1182120,I989639);
DFFARX1 I_69388 (I1182128,I2507,I1182094,I1182077,);
DFFARX1 I_69389 (I989657,I2507,I1182094,I1182168,);
not I_69390 (I1182176,I989648);
not I_69391 (I1182193,I989660);
nand I_69392 (I1182210,I1182193,I1182176);
nor I_69393 (I1182065,I1182168,I1182210);
DFFARX1 I_69394 (I1182210,I2507,I1182094,I1182250,);
not I_69395 (I1182086,I1182250);
not I_69396 (I1182272,I989666);
nand I_69397 (I1182289,I1182193,I1182272);
DFFARX1 I_69398 (I1182289,I2507,I1182094,I1182315,);
not I_69399 (I1182323,I1182315);
not I_69400 (I1182340,I989642);
nand I_69401 (I1182357,I1182340,I989663);
and I_69402 (I1182374,I1182176,I1182357);
nor I_69403 (I1182391,I1182289,I1182374);
DFFARX1 I_69404 (I1182391,I2507,I1182094,I1182062,);
DFFARX1 I_69405 (I1182374,I2507,I1182094,I1182083,);
nor I_69406 (I1182436,I989642,I989654);
nor I_69407 (I1182074,I1182289,I1182436);
or I_69408 (I1182467,I989642,I989654);
nor I_69409 (I1182484,I989639,I989651);
DFFARX1 I_69410 (I1182484,I2507,I1182094,I1182510,);
not I_69411 (I1182518,I1182510);
nor I_69412 (I1182080,I1182518,I1182323);
nand I_69413 (I1182549,I1182518,I1182168);
not I_69414 (I1182566,I989639);
nand I_69415 (I1182583,I1182566,I1182272);
nand I_69416 (I1182600,I1182518,I1182583);
nand I_69417 (I1182071,I1182600,I1182549);
nand I_69418 (I1182068,I1182583,I1182467);
not I_69419 (I1182672,I2514);
DFFARX1 I_69420 (I114962,I2507,I1182672,I1182698,);
and I_69421 (I1182706,I1182698,I114938);
DFFARX1 I_69422 (I1182706,I2507,I1182672,I1182655,);
DFFARX1 I_69423 (I114956,I2507,I1182672,I1182746,);
not I_69424 (I1182754,I114944);
not I_69425 (I1182771,I114941);
nand I_69426 (I1182788,I1182771,I1182754);
nor I_69427 (I1182643,I1182746,I1182788);
DFFARX1 I_69428 (I1182788,I2507,I1182672,I1182828,);
not I_69429 (I1182664,I1182828);
not I_69430 (I1182850,I114950);
nand I_69431 (I1182867,I1182771,I1182850);
DFFARX1 I_69432 (I1182867,I2507,I1182672,I1182893,);
not I_69433 (I1182901,I1182893);
not I_69434 (I1182918,I114941);
nand I_69435 (I1182935,I1182918,I114959);
and I_69436 (I1182952,I1182754,I1182935);
nor I_69437 (I1182969,I1182867,I1182952);
DFFARX1 I_69438 (I1182969,I2507,I1182672,I1182640,);
DFFARX1 I_69439 (I1182952,I2507,I1182672,I1182661,);
nor I_69440 (I1183014,I114941,I114953);
nor I_69441 (I1182652,I1182867,I1183014);
or I_69442 (I1183045,I114941,I114953);
nor I_69443 (I1183062,I114947,I114938);
DFFARX1 I_69444 (I1183062,I2507,I1182672,I1183088,);
not I_69445 (I1183096,I1183088);
nor I_69446 (I1182658,I1183096,I1182901);
nand I_69447 (I1183127,I1183096,I1182746);
not I_69448 (I1183144,I114947);
nand I_69449 (I1183161,I1183144,I1182850);
nand I_69450 (I1183178,I1183096,I1183161);
nand I_69451 (I1182649,I1183178,I1183127);
nand I_69452 (I1182646,I1183161,I1183045);
not I_69453 (I1183250,I2514);
DFFARX1 I_69454 (I322943,I2507,I1183250,I1183276,);
and I_69455 (I1183284,I1183276,I322928);
DFFARX1 I_69456 (I1183284,I2507,I1183250,I1183233,);
DFFARX1 I_69457 (I322934,I2507,I1183250,I1183324,);
not I_69458 (I1183332,I322916);
not I_69459 (I1183349,I322937);
nand I_69460 (I1183366,I1183349,I1183332);
nor I_69461 (I1183221,I1183324,I1183366);
DFFARX1 I_69462 (I1183366,I2507,I1183250,I1183406,);
not I_69463 (I1183242,I1183406);
not I_69464 (I1183428,I322940);
nand I_69465 (I1183445,I1183349,I1183428);
DFFARX1 I_69466 (I1183445,I2507,I1183250,I1183471,);
not I_69467 (I1183479,I1183471);
not I_69468 (I1183496,I322931);
nand I_69469 (I1183513,I1183496,I322919);
and I_69470 (I1183530,I1183332,I1183513);
nor I_69471 (I1183547,I1183445,I1183530);
DFFARX1 I_69472 (I1183547,I2507,I1183250,I1183218,);
DFFARX1 I_69473 (I1183530,I2507,I1183250,I1183239,);
nor I_69474 (I1183592,I322931,I322925);
nor I_69475 (I1183230,I1183445,I1183592);
or I_69476 (I1183623,I322931,I322925);
nor I_69477 (I1183640,I322922,I322916);
DFFARX1 I_69478 (I1183640,I2507,I1183250,I1183666,);
not I_69479 (I1183674,I1183666);
nor I_69480 (I1183236,I1183674,I1183479);
nand I_69481 (I1183705,I1183674,I1183324);
not I_69482 (I1183722,I322922);
nand I_69483 (I1183739,I1183722,I1183428);
nand I_69484 (I1183756,I1183674,I1183739);
nand I_69485 (I1183227,I1183756,I1183705);
nand I_69486 (I1183224,I1183739,I1183623);
not I_69487 (I1183828,I2514);
DFFARX1 I_69488 (I448495,I2507,I1183828,I1183854,);
and I_69489 (I1183862,I1183854,I448510);
DFFARX1 I_69490 (I1183862,I2507,I1183828,I1183811,);
DFFARX1 I_69491 (I448513,I2507,I1183828,I1183902,);
not I_69492 (I1183910,I448507);
not I_69493 (I1183927,I448522);
nand I_69494 (I1183944,I1183927,I1183910);
nor I_69495 (I1183799,I1183902,I1183944);
DFFARX1 I_69496 (I1183944,I2507,I1183828,I1183984,);
not I_69497 (I1183820,I1183984);
not I_69498 (I1184006,I448498);
nand I_69499 (I1184023,I1183927,I1184006);
DFFARX1 I_69500 (I1184023,I2507,I1183828,I1184049,);
not I_69501 (I1184057,I1184049);
not I_69502 (I1184074,I448501);
nand I_69503 (I1184091,I1184074,I448495);
and I_69504 (I1184108,I1183910,I1184091);
nor I_69505 (I1184125,I1184023,I1184108);
DFFARX1 I_69506 (I1184125,I2507,I1183828,I1183796,);
DFFARX1 I_69507 (I1184108,I2507,I1183828,I1183817,);
nor I_69508 (I1184170,I448501,I448504);
nor I_69509 (I1183808,I1184023,I1184170);
or I_69510 (I1184201,I448501,I448504);
nor I_69511 (I1184218,I448519,I448516);
DFFARX1 I_69512 (I1184218,I2507,I1183828,I1184244,);
not I_69513 (I1184252,I1184244);
nor I_69514 (I1183814,I1184252,I1184057);
nand I_69515 (I1184283,I1184252,I1183902);
not I_69516 (I1184300,I448519);
nand I_69517 (I1184317,I1184300,I1184006);
nand I_69518 (I1184334,I1184252,I1184317);
nand I_69519 (I1183805,I1184334,I1184283);
nand I_69520 (I1183802,I1184317,I1184201);
not I_69521 (I1184406,I2514);
DFFARX1 I_69522 (I688533,I2507,I1184406,I1184432,);
and I_69523 (I1184440,I1184432,I688521);
DFFARX1 I_69524 (I1184440,I2507,I1184406,I1184389,);
DFFARX1 I_69525 (I688524,I2507,I1184406,I1184480,);
not I_69526 (I1184488,I688518);
not I_69527 (I1184505,I688542);
nand I_69528 (I1184522,I1184505,I1184488);
nor I_69529 (I1184377,I1184480,I1184522);
DFFARX1 I_69530 (I1184522,I2507,I1184406,I1184562,);
not I_69531 (I1184398,I1184562);
not I_69532 (I1184584,I688530);
nand I_69533 (I1184601,I1184505,I1184584);
DFFARX1 I_69534 (I1184601,I2507,I1184406,I1184627,);
not I_69535 (I1184635,I1184627);
not I_69536 (I1184652,I688539);
nand I_69537 (I1184669,I1184652,I688536);
and I_69538 (I1184686,I1184488,I1184669);
nor I_69539 (I1184703,I1184601,I1184686);
DFFARX1 I_69540 (I1184703,I2507,I1184406,I1184374,);
DFFARX1 I_69541 (I1184686,I2507,I1184406,I1184395,);
nor I_69542 (I1184748,I688539,I688527);
nor I_69543 (I1184386,I1184601,I1184748);
or I_69544 (I1184779,I688539,I688527);
nor I_69545 (I1184796,I688518,I688521);
DFFARX1 I_69546 (I1184796,I2507,I1184406,I1184822,);
not I_69547 (I1184830,I1184822);
nor I_69548 (I1184392,I1184830,I1184635);
nand I_69549 (I1184861,I1184830,I1184480);
not I_69550 (I1184878,I688518);
nand I_69551 (I1184895,I1184878,I1184584);
nand I_69552 (I1184912,I1184830,I1184895);
nand I_69553 (I1184383,I1184912,I1184861);
nand I_69554 (I1184380,I1184895,I1184779);
not I_69555 (I1184984,I2514);
DFFARX1 I_69556 (I658477,I2507,I1184984,I1185010,);
and I_69557 (I1185018,I1185010,I658465);
DFFARX1 I_69558 (I1185018,I2507,I1184984,I1184967,);
DFFARX1 I_69559 (I658468,I2507,I1184984,I1185058,);
not I_69560 (I1185066,I658462);
not I_69561 (I1185083,I658486);
nand I_69562 (I1185100,I1185083,I1185066);
nor I_69563 (I1184955,I1185058,I1185100);
DFFARX1 I_69564 (I1185100,I2507,I1184984,I1185140,);
not I_69565 (I1184976,I1185140);
not I_69566 (I1185162,I658474);
nand I_69567 (I1185179,I1185083,I1185162);
DFFARX1 I_69568 (I1185179,I2507,I1184984,I1185205,);
not I_69569 (I1185213,I1185205);
not I_69570 (I1185230,I658483);
nand I_69571 (I1185247,I1185230,I658480);
and I_69572 (I1185264,I1185066,I1185247);
nor I_69573 (I1185281,I1185179,I1185264);
DFFARX1 I_69574 (I1185281,I2507,I1184984,I1184952,);
DFFARX1 I_69575 (I1185264,I2507,I1184984,I1184973,);
nor I_69576 (I1185326,I658483,I658471);
nor I_69577 (I1184964,I1185179,I1185326);
or I_69578 (I1185357,I658483,I658471);
nor I_69579 (I1185374,I658462,I658465);
DFFARX1 I_69580 (I1185374,I2507,I1184984,I1185400,);
not I_69581 (I1185408,I1185400);
nor I_69582 (I1184970,I1185408,I1185213);
nand I_69583 (I1185439,I1185408,I1185058);
not I_69584 (I1185456,I658462);
nand I_69585 (I1185473,I1185456,I1185162);
nand I_69586 (I1185490,I1185408,I1185473);
nand I_69587 (I1184961,I1185490,I1185439);
nand I_69588 (I1184958,I1185473,I1185357);
not I_69589 (I1185562,I2514);
DFFARX1 I_69590 (I598943,I2507,I1185562,I1185588,);
and I_69591 (I1185596,I1185588,I598931);
DFFARX1 I_69592 (I1185596,I2507,I1185562,I1185545,);
DFFARX1 I_69593 (I598946,I2507,I1185562,I1185636,);
not I_69594 (I1185644,I598937);
not I_69595 (I1185661,I598928);
nand I_69596 (I1185678,I1185661,I1185644);
nor I_69597 (I1185533,I1185636,I1185678);
DFFARX1 I_69598 (I1185678,I2507,I1185562,I1185718,);
not I_69599 (I1185554,I1185718);
not I_69600 (I1185740,I598934);
nand I_69601 (I1185757,I1185661,I1185740);
DFFARX1 I_69602 (I1185757,I2507,I1185562,I1185783,);
not I_69603 (I1185791,I1185783);
not I_69604 (I1185808,I598949);
nand I_69605 (I1185825,I1185808,I598952);
and I_69606 (I1185842,I1185644,I1185825);
nor I_69607 (I1185859,I1185757,I1185842);
DFFARX1 I_69608 (I1185859,I2507,I1185562,I1185530,);
DFFARX1 I_69609 (I1185842,I2507,I1185562,I1185551,);
nor I_69610 (I1185904,I598949,I598928);
nor I_69611 (I1185542,I1185757,I1185904);
or I_69612 (I1185935,I598949,I598928);
nor I_69613 (I1185952,I598940,I598931);
DFFARX1 I_69614 (I1185952,I2507,I1185562,I1185978,);
not I_69615 (I1185986,I1185978);
nor I_69616 (I1185548,I1185986,I1185791);
nand I_69617 (I1186017,I1185986,I1185636);
not I_69618 (I1186034,I598940);
nand I_69619 (I1186051,I1186034,I1185740);
nand I_69620 (I1186068,I1185986,I1186051);
nand I_69621 (I1185539,I1186068,I1186017);
nand I_69622 (I1185536,I1186051,I1185935);
not I_69623 (I1186140,I2514);
DFFARX1 I_69624 (I95463,I2507,I1186140,I1186166,);
and I_69625 (I1186174,I1186166,I95439);
DFFARX1 I_69626 (I1186174,I2507,I1186140,I1186123,);
DFFARX1 I_69627 (I95457,I2507,I1186140,I1186214,);
not I_69628 (I1186222,I95445);
not I_69629 (I1186239,I95442);
nand I_69630 (I1186256,I1186239,I1186222);
nor I_69631 (I1186111,I1186214,I1186256);
DFFARX1 I_69632 (I1186256,I2507,I1186140,I1186296,);
not I_69633 (I1186132,I1186296);
not I_69634 (I1186318,I95451);
nand I_69635 (I1186335,I1186239,I1186318);
DFFARX1 I_69636 (I1186335,I2507,I1186140,I1186361,);
not I_69637 (I1186369,I1186361);
not I_69638 (I1186386,I95442);
nand I_69639 (I1186403,I1186386,I95460);
and I_69640 (I1186420,I1186222,I1186403);
nor I_69641 (I1186437,I1186335,I1186420);
DFFARX1 I_69642 (I1186437,I2507,I1186140,I1186108,);
DFFARX1 I_69643 (I1186420,I2507,I1186140,I1186129,);
nor I_69644 (I1186482,I95442,I95454);
nor I_69645 (I1186120,I1186335,I1186482);
or I_69646 (I1186513,I95442,I95454);
nor I_69647 (I1186530,I95448,I95439);
DFFARX1 I_69648 (I1186530,I2507,I1186140,I1186556,);
not I_69649 (I1186564,I1186556);
nor I_69650 (I1186126,I1186564,I1186369);
nand I_69651 (I1186595,I1186564,I1186214);
not I_69652 (I1186612,I95448);
nand I_69653 (I1186629,I1186612,I1186318);
nand I_69654 (I1186646,I1186564,I1186629);
nand I_69655 (I1186117,I1186646,I1186595);
nand I_69656 (I1186114,I1186629,I1186513);
not I_69657 (I1186718,I2514);
DFFARX1 I_69658 (I1307719,I2507,I1186718,I1186744,);
and I_69659 (I1186752,I1186744,I1307701);
DFFARX1 I_69660 (I1186752,I2507,I1186718,I1186701,);
DFFARX1 I_69661 (I1307692,I2507,I1186718,I1186792,);
not I_69662 (I1186800,I1307707);
not I_69663 (I1186817,I1307695);
nand I_69664 (I1186834,I1186817,I1186800);
nor I_69665 (I1186689,I1186792,I1186834);
DFFARX1 I_69666 (I1186834,I2507,I1186718,I1186874,);
not I_69667 (I1186710,I1186874);
not I_69668 (I1186896,I1307704);
nand I_69669 (I1186913,I1186817,I1186896);
DFFARX1 I_69670 (I1186913,I2507,I1186718,I1186939,);
not I_69671 (I1186947,I1186939);
not I_69672 (I1186964,I1307713);
nand I_69673 (I1186981,I1186964,I1307692);
and I_69674 (I1186998,I1186800,I1186981);
nor I_69675 (I1187015,I1186913,I1186998);
DFFARX1 I_69676 (I1187015,I2507,I1186718,I1186686,);
DFFARX1 I_69677 (I1186998,I2507,I1186718,I1186707,);
nor I_69678 (I1187060,I1307713,I1307716);
nor I_69679 (I1186698,I1186913,I1187060);
or I_69680 (I1187091,I1307713,I1307716);
nor I_69681 (I1187108,I1307710,I1307698);
DFFARX1 I_69682 (I1187108,I2507,I1186718,I1187134,);
not I_69683 (I1187142,I1187134);
nor I_69684 (I1186704,I1187142,I1186947);
nand I_69685 (I1187173,I1187142,I1186792);
not I_69686 (I1187190,I1307710);
nand I_69687 (I1187207,I1187190,I1186896);
nand I_69688 (I1187224,I1187142,I1187207);
nand I_69689 (I1186695,I1187224,I1187173);
nand I_69690 (I1186692,I1187207,I1187091);
not I_69691 (I1187296,I2514);
DFFARX1 I_69692 (I882882,I2507,I1187296,I1187322,);
and I_69693 (I1187330,I1187322,I882888);
DFFARX1 I_69694 (I1187330,I2507,I1187296,I1187279,);
DFFARX1 I_69695 (I882894,I2507,I1187296,I1187370,);
not I_69696 (I1187378,I882879);
not I_69697 (I1187395,I882879);
nand I_69698 (I1187412,I1187395,I1187378);
nor I_69699 (I1187267,I1187370,I1187412);
DFFARX1 I_69700 (I1187412,I2507,I1187296,I1187452,);
not I_69701 (I1187288,I1187452);
not I_69702 (I1187474,I882897);
nand I_69703 (I1187491,I1187395,I1187474);
DFFARX1 I_69704 (I1187491,I2507,I1187296,I1187517,);
not I_69705 (I1187525,I1187517);
not I_69706 (I1187542,I882891);
nand I_69707 (I1187559,I1187542,I882882);
and I_69708 (I1187576,I1187378,I1187559);
nor I_69709 (I1187593,I1187491,I1187576);
DFFARX1 I_69710 (I1187593,I2507,I1187296,I1187264,);
DFFARX1 I_69711 (I1187576,I2507,I1187296,I1187285,);
nor I_69712 (I1187638,I882891,I882900);
nor I_69713 (I1187276,I1187491,I1187638);
or I_69714 (I1187669,I882891,I882900);
nor I_69715 (I1187686,I882885,I882885);
DFFARX1 I_69716 (I1187686,I2507,I1187296,I1187712,);
not I_69717 (I1187720,I1187712);
nor I_69718 (I1187282,I1187720,I1187525);
nand I_69719 (I1187751,I1187720,I1187370);
not I_69720 (I1187768,I882885);
nand I_69721 (I1187785,I1187768,I1187474);
nand I_69722 (I1187802,I1187720,I1187785);
nand I_69723 (I1187273,I1187802,I1187751);
nand I_69724 (I1187270,I1187785,I1187669);
not I_69725 (I1187874,I2514);
DFFARX1 I_69726 (I123394,I2507,I1187874,I1187900,);
and I_69727 (I1187908,I1187900,I123370);
DFFARX1 I_69728 (I1187908,I2507,I1187874,I1187857,);
DFFARX1 I_69729 (I123388,I2507,I1187874,I1187948,);
not I_69730 (I1187956,I123376);
not I_69731 (I1187973,I123373);
nand I_69732 (I1187990,I1187973,I1187956);
nor I_69733 (I1187845,I1187948,I1187990);
DFFARX1 I_69734 (I1187990,I2507,I1187874,I1188030,);
not I_69735 (I1187866,I1188030);
not I_69736 (I1188052,I123382);
nand I_69737 (I1188069,I1187973,I1188052);
DFFARX1 I_69738 (I1188069,I2507,I1187874,I1188095,);
not I_69739 (I1188103,I1188095);
not I_69740 (I1188120,I123373);
nand I_69741 (I1188137,I1188120,I123391);
and I_69742 (I1188154,I1187956,I1188137);
nor I_69743 (I1188171,I1188069,I1188154);
DFFARX1 I_69744 (I1188171,I2507,I1187874,I1187842,);
DFFARX1 I_69745 (I1188154,I2507,I1187874,I1187863,);
nor I_69746 (I1188216,I123373,I123385);
nor I_69747 (I1187854,I1188069,I1188216);
or I_69748 (I1188247,I123373,I123385);
nor I_69749 (I1188264,I123379,I123370);
DFFARX1 I_69750 (I1188264,I2507,I1187874,I1188290,);
not I_69751 (I1188298,I1188290);
nor I_69752 (I1187860,I1188298,I1188103);
nand I_69753 (I1188329,I1188298,I1187948);
not I_69754 (I1188346,I123379);
nand I_69755 (I1188363,I1188346,I1188052);
nand I_69756 (I1188380,I1188298,I1188363);
nand I_69757 (I1187851,I1188380,I1188329);
nand I_69758 (I1187848,I1188363,I1188247);
not I_69759 (I1188452,I2514);
DFFARX1 I_69760 (I1235191,I2507,I1188452,I1188478,);
and I_69761 (I1188486,I1188478,I1235185);
DFFARX1 I_69762 (I1188486,I2507,I1188452,I1188435,);
DFFARX1 I_69763 (I1235170,I2507,I1188452,I1188526,);
not I_69764 (I1188534,I1235176);
not I_69765 (I1188551,I1235188);
nand I_69766 (I1188568,I1188551,I1188534);
nor I_69767 (I1188423,I1188526,I1188568);
DFFARX1 I_69768 (I1188568,I2507,I1188452,I1188608,);
not I_69769 (I1188444,I1188608);
not I_69770 (I1188630,I1235170);
nand I_69771 (I1188647,I1188551,I1188630);
DFFARX1 I_69772 (I1188647,I2507,I1188452,I1188673,);
not I_69773 (I1188681,I1188673);
not I_69774 (I1188698,I1235194);
nand I_69775 (I1188715,I1188698,I1235182);
and I_69776 (I1188732,I1188534,I1188715);
nor I_69777 (I1188749,I1188647,I1188732);
DFFARX1 I_69778 (I1188749,I2507,I1188452,I1188420,);
DFFARX1 I_69779 (I1188732,I2507,I1188452,I1188441,);
nor I_69780 (I1188794,I1235194,I1235173);
nor I_69781 (I1188432,I1188647,I1188794);
or I_69782 (I1188825,I1235194,I1235173);
nor I_69783 (I1188842,I1235179,I1235173);
DFFARX1 I_69784 (I1188842,I2507,I1188452,I1188868,);
not I_69785 (I1188876,I1188868);
nor I_69786 (I1188438,I1188876,I1188681);
nand I_69787 (I1188907,I1188876,I1188526);
not I_69788 (I1188924,I1235179);
nand I_69789 (I1188941,I1188924,I1188630);
nand I_69790 (I1188958,I1188876,I1188941);
nand I_69791 (I1188429,I1188958,I1188907);
nand I_69792 (I1188426,I1188941,I1188825);
not I_69793 (I1189030,I2514);
DFFARX1 I_69794 (I516107,I2507,I1189030,I1189056,);
and I_69795 (I1189064,I1189056,I516122);
DFFARX1 I_69796 (I1189064,I2507,I1189030,I1189013,);
DFFARX1 I_69797 (I516113,I2507,I1189030,I1189104,);
not I_69798 (I1189112,I516107);
not I_69799 (I1189129,I516125);
nand I_69800 (I1189146,I1189129,I1189112);
nor I_69801 (I1189001,I1189104,I1189146);
DFFARX1 I_69802 (I1189146,I2507,I1189030,I1189186,);
not I_69803 (I1189022,I1189186);
not I_69804 (I1189208,I516116);
nand I_69805 (I1189225,I1189129,I1189208);
DFFARX1 I_69806 (I1189225,I2507,I1189030,I1189251,);
not I_69807 (I1189259,I1189251);
not I_69808 (I1189276,I516128);
nand I_69809 (I1189293,I1189276,I516104);
and I_69810 (I1189310,I1189112,I1189293);
nor I_69811 (I1189327,I1189225,I1189310);
DFFARX1 I_69812 (I1189327,I2507,I1189030,I1188998,);
DFFARX1 I_69813 (I1189310,I2507,I1189030,I1189019,);
nor I_69814 (I1189372,I516128,I516104);
nor I_69815 (I1189010,I1189225,I1189372);
or I_69816 (I1189403,I516128,I516104);
nor I_69817 (I1189420,I516110,I516119);
DFFARX1 I_69818 (I1189420,I2507,I1189030,I1189446,);
not I_69819 (I1189454,I1189446);
nor I_69820 (I1189016,I1189454,I1189259);
nand I_69821 (I1189485,I1189454,I1189104);
not I_69822 (I1189502,I516110);
nand I_69823 (I1189519,I1189502,I1189208);
nand I_69824 (I1189536,I1189454,I1189519);
nand I_69825 (I1189007,I1189536,I1189485);
nand I_69826 (I1189004,I1189519,I1189403);
not I_69827 (I1189608,I2514);
DFFARX1 I_69828 (I987061,I2507,I1189608,I1189634,);
and I_69829 (I1189642,I1189634,I987055);
DFFARX1 I_69830 (I1189642,I2507,I1189608,I1189591,);
DFFARX1 I_69831 (I987073,I2507,I1189608,I1189682,);
not I_69832 (I1189690,I987064);
not I_69833 (I1189707,I987076);
nand I_69834 (I1189724,I1189707,I1189690);
nor I_69835 (I1189579,I1189682,I1189724);
DFFARX1 I_69836 (I1189724,I2507,I1189608,I1189764,);
not I_69837 (I1189600,I1189764);
not I_69838 (I1189786,I987082);
nand I_69839 (I1189803,I1189707,I1189786);
DFFARX1 I_69840 (I1189803,I2507,I1189608,I1189829,);
not I_69841 (I1189837,I1189829);
not I_69842 (I1189854,I987058);
nand I_69843 (I1189871,I1189854,I987079);
and I_69844 (I1189888,I1189690,I1189871);
nor I_69845 (I1189905,I1189803,I1189888);
DFFARX1 I_69846 (I1189905,I2507,I1189608,I1189576,);
DFFARX1 I_69847 (I1189888,I2507,I1189608,I1189597,);
nor I_69848 (I1189950,I987058,I987070);
nor I_69849 (I1189588,I1189803,I1189950);
or I_69850 (I1189981,I987058,I987070);
nor I_69851 (I1189998,I987055,I987067);
DFFARX1 I_69852 (I1189998,I2507,I1189608,I1190024,);
not I_69853 (I1190032,I1190024);
nor I_69854 (I1189594,I1190032,I1189837);
nand I_69855 (I1190063,I1190032,I1189682);
not I_69856 (I1190080,I987055);
nand I_69857 (I1190097,I1190080,I1189786);
nand I_69858 (I1190114,I1190032,I1190097);
nand I_69859 (I1189585,I1190114,I1190063);
nand I_69860 (I1189582,I1190097,I1189981);
not I_69861 (I1190186,I2514);
DFFARX1 I_69862 (I586227,I2507,I1190186,I1190212,);
and I_69863 (I1190220,I1190212,I586215);
DFFARX1 I_69864 (I1190220,I2507,I1190186,I1190169,);
DFFARX1 I_69865 (I586230,I2507,I1190186,I1190260,);
not I_69866 (I1190268,I586221);
not I_69867 (I1190285,I586212);
nand I_69868 (I1190302,I1190285,I1190268);
nor I_69869 (I1190157,I1190260,I1190302);
DFFARX1 I_69870 (I1190302,I2507,I1190186,I1190342,);
not I_69871 (I1190178,I1190342);
not I_69872 (I1190364,I586218);
nand I_69873 (I1190381,I1190285,I1190364);
DFFARX1 I_69874 (I1190381,I2507,I1190186,I1190407,);
not I_69875 (I1190415,I1190407);
not I_69876 (I1190432,I586233);
nand I_69877 (I1190449,I1190432,I586236);
and I_69878 (I1190466,I1190268,I1190449);
nor I_69879 (I1190483,I1190381,I1190466);
DFFARX1 I_69880 (I1190483,I2507,I1190186,I1190154,);
DFFARX1 I_69881 (I1190466,I2507,I1190186,I1190175,);
nor I_69882 (I1190528,I586233,I586212);
nor I_69883 (I1190166,I1190381,I1190528);
or I_69884 (I1190559,I586233,I586212);
nor I_69885 (I1190576,I586224,I586215);
DFFARX1 I_69886 (I1190576,I2507,I1190186,I1190602,);
not I_69887 (I1190610,I1190602);
nor I_69888 (I1190172,I1190610,I1190415);
nand I_69889 (I1190641,I1190610,I1190260);
not I_69890 (I1190658,I586224);
nand I_69891 (I1190675,I1190658,I1190364);
nand I_69892 (I1190692,I1190610,I1190675);
nand I_69893 (I1190163,I1190692,I1190641);
nand I_69894 (I1190160,I1190675,I1190559);
not I_69895 (I1190764,I2514);
DFFARX1 I_69896 (I630155,I2507,I1190764,I1190790,);
and I_69897 (I1190798,I1190790,I630143);
DFFARX1 I_69898 (I1190798,I2507,I1190764,I1190747,);
DFFARX1 I_69899 (I630146,I2507,I1190764,I1190838,);
not I_69900 (I1190846,I630140);
not I_69901 (I1190863,I630164);
nand I_69902 (I1190880,I1190863,I1190846);
nor I_69903 (I1190735,I1190838,I1190880);
DFFARX1 I_69904 (I1190880,I2507,I1190764,I1190920,);
not I_69905 (I1190756,I1190920);
not I_69906 (I1190942,I630152);
nand I_69907 (I1190959,I1190863,I1190942);
DFFARX1 I_69908 (I1190959,I2507,I1190764,I1190985,);
not I_69909 (I1190993,I1190985);
not I_69910 (I1191010,I630161);
nand I_69911 (I1191027,I1191010,I630158);
and I_69912 (I1191044,I1190846,I1191027);
nor I_69913 (I1191061,I1190959,I1191044);
DFFARX1 I_69914 (I1191061,I2507,I1190764,I1190732,);
DFFARX1 I_69915 (I1191044,I2507,I1190764,I1190753,);
nor I_69916 (I1191106,I630161,I630149);
nor I_69917 (I1190744,I1190959,I1191106);
or I_69918 (I1191137,I630161,I630149);
nor I_69919 (I1191154,I630140,I630143);
DFFARX1 I_69920 (I1191154,I2507,I1190764,I1191180,);
not I_69921 (I1191188,I1191180);
nor I_69922 (I1190750,I1191188,I1190993);
nand I_69923 (I1191219,I1191188,I1190838);
not I_69924 (I1191236,I630140);
nand I_69925 (I1191253,I1191236,I1190942);
nand I_69926 (I1191270,I1191188,I1191253);
nand I_69927 (I1190741,I1191270,I1191219);
nand I_69928 (I1190738,I1191253,I1191137);
not I_69929 (I1191342,I2514);
DFFARX1 I_69930 (I1247159,I2507,I1191342,I1191368,);
and I_69931 (I1191376,I1191368,I1247153);
DFFARX1 I_69932 (I1191376,I2507,I1191342,I1191325,);
DFFARX1 I_69933 (I1247138,I2507,I1191342,I1191416,);
not I_69934 (I1191424,I1247144);
not I_69935 (I1191441,I1247156);
nand I_69936 (I1191458,I1191441,I1191424);
nor I_69937 (I1191313,I1191416,I1191458);
DFFARX1 I_69938 (I1191458,I2507,I1191342,I1191498,);
not I_69939 (I1191334,I1191498);
not I_69940 (I1191520,I1247138);
nand I_69941 (I1191537,I1191441,I1191520);
DFFARX1 I_69942 (I1191537,I2507,I1191342,I1191563,);
not I_69943 (I1191571,I1191563);
not I_69944 (I1191588,I1247162);
nand I_69945 (I1191605,I1191588,I1247150);
and I_69946 (I1191622,I1191424,I1191605);
nor I_69947 (I1191639,I1191537,I1191622);
DFFARX1 I_69948 (I1191639,I2507,I1191342,I1191310,);
DFFARX1 I_69949 (I1191622,I2507,I1191342,I1191331,);
nor I_69950 (I1191684,I1247162,I1247141);
nor I_69951 (I1191322,I1191537,I1191684);
or I_69952 (I1191715,I1247162,I1247141);
nor I_69953 (I1191732,I1247147,I1247141);
DFFARX1 I_69954 (I1191732,I2507,I1191342,I1191758,);
not I_69955 (I1191766,I1191758);
nor I_69956 (I1191328,I1191766,I1191571);
nand I_69957 (I1191797,I1191766,I1191416);
not I_69958 (I1191814,I1247147);
nand I_69959 (I1191831,I1191814,I1191520);
nand I_69960 (I1191848,I1191766,I1191831);
nand I_69961 (I1191319,I1191848,I1191797);
nand I_69962 (I1191316,I1191831,I1191715);
not I_69963 (I1191920,I2514);
DFFARX1 I_69964 (I362468,I2507,I1191920,I1191946,);
and I_69965 (I1191954,I1191946,I362453);
DFFARX1 I_69966 (I1191954,I2507,I1191920,I1191903,);
DFFARX1 I_69967 (I362459,I2507,I1191920,I1191994,);
not I_69968 (I1192002,I362441);
not I_69969 (I1192019,I362462);
nand I_69970 (I1192036,I1192019,I1192002);
nor I_69971 (I1191891,I1191994,I1192036);
DFFARX1 I_69972 (I1192036,I2507,I1191920,I1192076,);
not I_69973 (I1191912,I1192076);
not I_69974 (I1192098,I362465);
nand I_69975 (I1192115,I1192019,I1192098);
DFFARX1 I_69976 (I1192115,I2507,I1191920,I1192141,);
not I_69977 (I1192149,I1192141);
not I_69978 (I1192166,I362456);
nand I_69979 (I1192183,I1192166,I362444);
and I_69980 (I1192200,I1192002,I1192183);
nor I_69981 (I1192217,I1192115,I1192200);
DFFARX1 I_69982 (I1192217,I2507,I1191920,I1191888,);
DFFARX1 I_69983 (I1192200,I2507,I1191920,I1191909,);
nor I_69984 (I1192262,I362456,I362450);
nor I_69985 (I1191900,I1192115,I1192262);
or I_69986 (I1192293,I362456,I362450);
nor I_69987 (I1192310,I362447,I362441);
DFFARX1 I_69988 (I1192310,I2507,I1191920,I1192336,);
not I_69989 (I1192344,I1192336);
nor I_69990 (I1191906,I1192344,I1192149);
nand I_69991 (I1192375,I1192344,I1191994);
not I_69992 (I1192392,I362447);
nand I_69993 (I1192409,I1192392,I1192098);
nand I_69994 (I1192426,I1192344,I1192409);
nand I_69995 (I1191897,I1192426,I1192375);
nand I_69996 (I1191894,I1192409,I1192293);
not I_69997 (I1192498,I2514);
DFFARX1 I_69998 (I777482,I2507,I1192498,I1192524,);
and I_69999 (I1192532,I1192524,I777488);
DFFARX1 I_70000 (I1192532,I2507,I1192498,I1192481,);
DFFARX1 I_70001 (I777494,I2507,I1192498,I1192572,);
not I_70002 (I1192580,I777479);
not I_70003 (I1192597,I777479);
nand I_70004 (I1192614,I1192597,I1192580);
nor I_70005 (I1192469,I1192572,I1192614);
DFFARX1 I_70006 (I1192614,I2507,I1192498,I1192654,);
not I_70007 (I1192490,I1192654);
not I_70008 (I1192676,I777497);
nand I_70009 (I1192693,I1192597,I1192676);
DFFARX1 I_70010 (I1192693,I2507,I1192498,I1192719,);
not I_70011 (I1192727,I1192719);
not I_70012 (I1192744,I777491);
nand I_70013 (I1192761,I1192744,I777482);
and I_70014 (I1192778,I1192580,I1192761);
nor I_70015 (I1192795,I1192693,I1192778);
DFFARX1 I_70016 (I1192795,I2507,I1192498,I1192466,);
DFFARX1 I_70017 (I1192778,I2507,I1192498,I1192487,);
nor I_70018 (I1192840,I777491,I777500);
nor I_70019 (I1192478,I1192693,I1192840);
or I_70020 (I1192871,I777491,I777500);
nor I_70021 (I1192888,I777485,I777485);
DFFARX1 I_70022 (I1192888,I2507,I1192498,I1192914,);
not I_70023 (I1192922,I1192914);
nor I_70024 (I1192484,I1192922,I1192727);
nand I_70025 (I1192953,I1192922,I1192572);
not I_70026 (I1192970,I777485);
nand I_70027 (I1192987,I1192970,I1192676);
nand I_70028 (I1193004,I1192922,I1192987);
nand I_70029 (I1192475,I1193004,I1192953);
nand I_70030 (I1192472,I1192987,I1192871);
not I_70031 (I1193076,I2514);
DFFARX1 I_70032 (I314511,I2507,I1193076,I1193102,);
and I_70033 (I1193110,I1193102,I314496);
DFFARX1 I_70034 (I1193110,I2507,I1193076,I1193059,);
DFFARX1 I_70035 (I314502,I2507,I1193076,I1193150,);
not I_70036 (I1193158,I314484);
not I_70037 (I1193175,I314505);
nand I_70038 (I1193192,I1193175,I1193158);
nor I_70039 (I1193047,I1193150,I1193192);
DFFARX1 I_70040 (I1193192,I2507,I1193076,I1193232,);
not I_70041 (I1193068,I1193232);
not I_70042 (I1193254,I314508);
nand I_70043 (I1193271,I1193175,I1193254);
DFFARX1 I_70044 (I1193271,I2507,I1193076,I1193297,);
not I_70045 (I1193305,I1193297);
not I_70046 (I1193322,I314499);
nand I_70047 (I1193339,I1193322,I314487);
and I_70048 (I1193356,I1193158,I1193339);
nor I_70049 (I1193373,I1193271,I1193356);
DFFARX1 I_70050 (I1193373,I2507,I1193076,I1193044,);
DFFARX1 I_70051 (I1193356,I2507,I1193076,I1193065,);
nor I_70052 (I1193418,I314499,I314493);
nor I_70053 (I1193056,I1193271,I1193418);
or I_70054 (I1193449,I314499,I314493);
nor I_70055 (I1193466,I314490,I314484);
DFFARX1 I_70056 (I1193466,I2507,I1193076,I1193492,);
not I_70057 (I1193500,I1193492);
nor I_70058 (I1193062,I1193500,I1193305);
nand I_70059 (I1193531,I1193500,I1193150);
not I_70060 (I1193548,I314490);
nand I_70061 (I1193565,I1193548,I1193254);
nand I_70062 (I1193582,I1193500,I1193565);
nand I_70063 (I1193053,I1193582,I1193531);
nand I_70064 (I1193050,I1193565,I1193449);
not I_70065 (I1193654,I2514);
DFFARX1 I_70066 (I497662,I2507,I1193654,I1193680,);
and I_70067 (I1193688,I1193680,I497677);
DFFARX1 I_70068 (I1193688,I2507,I1193654,I1193637,);
DFFARX1 I_70069 (I497668,I2507,I1193654,I1193728,);
not I_70070 (I1193736,I497662);
not I_70071 (I1193753,I497680);
nand I_70072 (I1193770,I1193753,I1193736);
nor I_70073 (I1193625,I1193728,I1193770);
DFFARX1 I_70074 (I1193770,I2507,I1193654,I1193810,);
not I_70075 (I1193646,I1193810);
not I_70076 (I1193832,I497671);
nand I_70077 (I1193849,I1193753,I1193832);
DFFARX1 I_70078 (I1193849,I2507,I1193654,I1193875,);
not I_70079 (I1193883,I1193875);
not I_70080 (I1193900,I497683);
nand I_70081 (I1193917,I1193900,I497659);
and I_70082 (I1193934,I1193736,I1193917);
nor I_70083 (I1193951,I1193849,I1193934);
DFFARX1 I_70084 (I1193951,I2507,I1193654,I1193622,);
DFFARX1 I_70085 (I1193934,I2507,I1193654,I1193643,);
nor I_70086 (I1193996,I497683,I497659);
nor I_70087 (I1193634,I1193849,I1193996);
or I_70088 (I1194027,I497683,I497659);
nor I_70089 (I1194044,I497665,I497674);
DFFARX1 I_70090 (I1194044,I2507,I1193654,I1194070,);
not I_70091 (I1194078,I1194070);
nor I_70092 (I1193640,I1194078,I1193883);
nand I_70093 (I1194109,I1194078,I1193728);
not I_70094 (I1194126,I497665);
nand I_70095 (I1194143,I1194126,I1193832);
nand I_70096 (I1194160,I1194078,I1194143);
nand I_70097 (I1193631,I1194160,I1194109);
nand I_70098 (I1193628,I1194143,I1194027);
not I_70099 (I1194232,I2514);
DFFARX1 I_70100 (I159155,I2507,I1194232,I1194258,);
and I_70101 (I1194266,I1194258,I159158);
DFFARX1 I_70102 (I1194266,I2507,I1194232,I1194215,);
DFFARX1 I_70103 (I159158,I2507,I1194232,I1194306,);
not I_70104 (I1194314,I159173);
not I_70105 (I1194331,I159179);
nand I_70106 (I1194348,I1194331,I1194314);
nor I_70107 (I1194203,I1194306,I1194348);
DFFARX1 I_70108 (I1194348,I2507,I1194232,I1194388,);
not I_70109 (I1194224,I1194388);
not I_70110 (I1194410,I159167);
nand I_70111 (I1194427,I1194331,I1194410);
DFFARX1 I_70112 (I1194427,I2507,I1194232,I1194453,);
not I_70113 (I1194461,I1194453);
not I_70114 (I1194478,I159164);
nand I_70115 (I1194495,I1194478,I159161);
and I_70116 (I1194512,I1194314,I1194495);
nor I_70117 (I1194529,I1194427,I1194512);
DFFARX1 I_70118 (I1194529,I2507,I1194232,I1194200,);
DFFARX1 I_70119 (I1194512,I2507,I1194232,I1194221,);
nor I_70120 (I1194574,I159164,I159155);
nor I_70121 (I1194212,I1194427,I1194574);
or I_70122 (I1194605,I159164,I159155);
nor I_70123 (I1194622,I159170,I159176);
DFFARX1 I_70124 (I1194622,I2507,I1194232,I1194648,);
not I_70125 (I1194656,I1194648);
nor I_70126 (I1194218,I1194656,I1194461);
nand I_70127 (I1194687,I1194656,I1194306);
not I_70128 (I1194704,I159170);
nand I_70129 (I1194721,I1194704,I1194410);
nand I_70130 (I1194738,I1194656,I1194721);
nand I_70131 (I1194209,I1194738,I1194687);
nand I_70132 (I1194206,I1194721,I1194605);
not I_70133 (I1194810,I2514);
DFFARX1 I_70134 (I659055,I2507,I1194810,I1194836,);
and I_70135 (I1194844,I1194836,I659043);
DFFARX1 I_70136 (I1194844,I2507,I1194810,I1194793,);
DFFARX1 I_70137 (I659046,I2507,I1194810,I1194884,);
not I_70138 (I1194892,I659040);
not I_70139 (I1194909,I659064);
nand I_70140 (I1194926,I1194909,I1194892);
nor I_70141 (I1194781,I1194884,I1194926);
DFFARX1 I_70142 (I1194926,I2507,I1194810,I1194966,);
not I_70143 (I1194802,I1194966);
not I_70144 (I1194988,I659052);
nand I_70145 (I1195005,I1194909,I1194988);
DFFARX1 I_70146 (I1195005,I2507,I1194810,I1195031,);
not I_70147 (I1195039,I1195031);
not I_70148 (I1195056,I659061);
nand I_70149 (I1195073,I1195056,I659058);
and I_70150 (I1195090,I1194892,I1195073);
nor I_70151 (I1195107,I1195005,I1195090);
DFFARX1 I_70152 (I1195107,I2507,I1194810,I1194778,);
DFFARX1 I_70153 (I1195090,I2507,I1194810,I1194799,);
nor I_70154 (I1195152,I659061,I659049);
nor I_70155 (I1194790,I1195005,I1195152);
or I_70156 (I1195183,I659061,I659049);
nor I_70157 (I1195200,I659040,I659043);
DFFARX1 I_70158 (I1195200,I2507,I1194810,I1195226,);
not I_70159 (I1195234,I1195226);
nor I_70160 (I1194796,I1195234,I1195039);
nand I_70161 (I1195265,I1195234,I1194884);
not I_70162 (I1195282,I659040);
nand I_70163 (I1195299,I1195282,I1194988);
nand I_70164 (I1195316,I1195234,I1195299);
nand I_70165 (I1194787,I1195316,I1195265);
nand I_70166 (I1194784,I1195299,I1195183);
not I_70167 (I1195388,I2514);
DFFARX1 I_70168 (I1277898,I2507,I1195388,I1195414,);
and I_70169 (I1195422,I1195414,I1277880);
DFFARX1 I_70170 (I1195422,I2507,I1195388,I1195371,);
DFFARX1 I_70171 (I1277889,I2507,I1195388,I1195462,);
not I_70172 (I1195470,I1277874);
not I_70173 (I1195487,I1277886);
nand I_70174 (I1195504,I1195487,I1195470);
nor I_70175 (I1195359,I1195462,I1195504);
DFFARX1 I_70176 (I1195504,I2507,I1195388,I1195544,);
not I_70177 (I1195380,I1195544);
not I_70178 (I1195566,I1277877);
nand I_70179 (I1195583,I1195487,I1195566);
DFFARX1 I_70180 (I1195583,I2507,I1195388,I1195609,);
not I_70181 (I1195617,I1195609);
not I_70182 (I1195634,I1277874);
nand I_70183 (I1195651,I1195634,I1277877);
and I_70184 (I1195668,I1195470,I1195651);
nor I_70185 (I1195685,I1195583,I1195668);
DFFARX1 I_70186 (I1195685,I2507,I1195388,I1195356,);
DFFARX1 I_70187 (I1195668,I2507,I1195388,I1195377,);
nor I_70188 (I1195730,I1277874,I1277895);
nor I_70189 (I1195368,I1195583,I1195730);
or I_70190 (I1195761,I1277874,I1277895);
nor I_70191 (I1195778,I1277883,I1277892);
DFFARX1 I_70192 (I1195778,I2507,I1195388,I1195804,);
not I_70193 (I1195812,I1195804);
nor I_70194 (I1195374,I1195812,I1195617);
nand I_70195 (I1195843,I1195812,I1195462);
not I_70196 (I1195860,I1277883);
nand I_70197 (I1195877,I1195860,I1195566);
nand I_70198 (I1195894,I1195812,I1195877);
nand I_70199 (I1195365,I1195894,I1195843);
nand I_70200 (I1195362,I1195877,I1195761);
not I_70201 (I1195966,I2514);
DFFARX1 I_70202 (I318200,I2507,I1195966,I1195992,);
and I_70203 (I1196000,I1195992,I318185);
DFFARX1 I_70204 (I1196000,I2507,I1195966,I1195949,);
DFFARX1 I_70205 (I318191,I2507,I1195966,I1196040,);
not I_70206 (I1196048,I318173);
not I_70207 (I1196065,I318194);
nand I_70208 (I1196082,I1196065,I1196048);
nor I_70209 (I1195937,I1196040,I1196082);
DFFARX1 I_70210 (I1196082,I2507,I1195966,I1196122,);
not I_70211 (I1195958,I1196122);
not I_70212 (I1196144,I318197);
nand I_70213 (I1196161,I1196065,I1196144);
DFFARX1 I_70214 (I1196161,I2507,I1195966,I1196187,);
not I_70215 (I1196195,I1196187);
not I_70216 (I1196212,I318188);
nand I_70217 (I1196229,I1196212,I318176);
and I_70218 (I1196246,I1196048,I1196229);
nor I_70219 (I1196263,I1196161,I1196246);
DFFARX1 I_70220 (I1196263,I2507,I1195966,I1195934,);
DFFARX1 I_70221 (I1196246,I2507,I1195966,I1195955,);
nor I_70222 (I1196308,I318188,I318182);
nor I_70223 (I1195946,I1196161,I1196308);
or I_70224 (I1196339,I318188,I318182);
nor I_70225 (I1196356,I318179,I318173);
DFFARX1 I_70226 (I1196356,I2507,I1195966,I1196382,);
not I_70227 (I1196390,I1196382);
nor I_70228 (I1195952,I1196390,I1196195);
nand I_70229 (I1196421,I1196390,I1196040);
not I_70230 (I1196438,I318179);
nand I_70231 (I1196455,I1196438,I1196144);
nand I_70232 (I1196472,I1196390,I1196455);
nand I_70233 (I1195943,I1196472,I1196421);
nand I_70234 (I1195940,I1196455,I1196339);
not I_70235 (I1196544,I2514);
DFFARX1 I_70236 (I118651,I2507,I1196544,I1196570,);
and I_70237 (I1196578,I1196570,I118627);
DFFARX1 I_70238 (I1196578,I2507,I1196544,I1196527,);
DFFARX1 I_70239 (I118645,I2507,I1196544,I1196618,);
not I_70240 (I1196626,I118633);
not I_70241 (I1196643,I118630);
nand I_70242 (I1196660,I1196643,I1196626);
nor I_70243 (I1196515,I1196618,I1196660);
DFFARX1 I_70244 (I1196660,I2507,I1196544,I1196700,);
not I_70245 (I1196536,I1196700);
not I_70246 (I1196722,I118639);
nand I_70247 (I1196739,I1196643,I1196722);
DFFARX1 I_70248 (I1196739,I2507,I1196544,I1196765,);
not I_70249 (I1196773,I1196765);
not I_70250 (I1196790,I118630);
nand I_70251 (I1196807,I1196790,I118648);
and I_70252 (I1196824,I1196626,I1196807);
nor I_70253 (I1196841,I1196739,I1196824);
DFFARX1 I_70254 (I1196841,I2507,I1196544,I1196512,);
DFFARX1 I_70255 (I1196824,I2507,I1196544,I1196533,);
nor I_70256 (I1196886,I118630,I118642);
nor I_70257 (I1196524,I1196739,I1196886);
or I_70258 (I1196917,I118630,I118642);
nor I_70259 (I1196934,I118636,I118627);
DFFARX1 I_70260 (I1196934,I2507,I1196544,I1196960,);
not I_70261 (I1196968,I1196960);
nor I_70262 (I1196530,I1196968,I1196773);
nand I_70263 (I1196999,I1196968,I1196618);
not I_70264 (I1197016,I118636);
nand I_70265 (I1197033,I1197016,I1196722);
nand I_70266 (I1197050,I1196968,I1197033);
nand I_70267 (I1196521,I1197050,I1196999);
nand I_70268 (I1196518,I1197033,I1196917);
not I_70269 (I1197122,I2514);
DFFARX1 I_70270 (I55938,I2507,I1197122,I1197148,);
and I_70271 (I1197156,I1197148,I55914);
DFFARX1 I_70272 (I1197156,I2507,I1197122,I1197105,);
DFFARX1 I_70273 (I55932,I2507,I1197122,I1197196,);
not I_70274 (I1197204,I55920);
not I_70275 (I1197221,I55917);
nand I_70276 (I1197238,I1197221,I1197204);
nor I_70277 (I1197093,I1197196,I1197238);
DFFARX1 I_70278 (I1197238,I2507,I1197122,I1197278,);
not I_70279 (I1197114,I1197278);
not I_70280 (I1197300,I55926);
nand I_70281 (I1197317,I1197221,I1197300);
DFFARX1 I_70282 (I1197317,I2507,I1197122,I1197343,);
not I_70283 (I1197351,I1197343);
not I_70284 (I1197368,I55917);
nand I_70285 (I1197385,I1197368,I55935);
and I_70286 (I1197402,I1197204,I1197385);
nor I_70287 (I1197419,I1197317,I1197402);
DFFARX1 I_70288 (I1197419,I2507,I1197122,I1197090,);
DFFARX1 I_70289 (I1197402,I2507,I1197122,I1197111,);
nor I_70290 (I1197464,I55917,I55929);
nor I_70291 (I1197102,I1197317,I1197464);
or I_70292 (I1197495,I55917,I55929);
nor I_70293 (I1197512,I55923,I55914);
DFFARX1 I_70294 (I1197512,I2507,I1197122,I1197538,);
not I_70295 (I1197546,I1197538);
nor I_70296 (I1197108,I1197546,I1197351);
nand I_70297 (I1197577,I1197546,I1197196);
not I_70298 (I1197594,I55923);
nand I_70299 (I1197611,I1197594,I1197300);
nand I_70300 (I1197628,I1197546,I1197611);
nand I_70301 (I1197099,I1197628,I1197577);
nand I_70302 (I1197096,I1197611,I1197495);
not I_70303 (I1197700,I2514);
DFFARX1 I_70304 (I756159,I2507,I1197700,I1197726,);
and I_70305 (I1197734,I1197726,I756147);
DFFARX1 I_70306 (I1197734,I2507,I1197700,I1197683,);
DFFARX1 I_70307 (I756150,I2507,I1197700,I1197774,);
not I_70308 (I1197782,I756144);
not I_70309 (I1197799,I756168);
nand I_70310 (I1197816,I1197799,I1197782);
nor I_70311 (I1197671,I1197774,I1197816);
DFFARX1 I_70312 (I1197816,I2507,I1197700,I1197856,);
not I_70313 (I1197692,I1197856);
not I_70314 (I1197878,I756156);
nand I_70315 (I1197895,I1197799,I1197878);
DFFARX1 I_70316 (I1197895,I2507,I1197700,I1197921,);
not I_70317 (I1197929,I1197921);
not I_70318 (I1197946,I756165);
nand I_70319 (I1197963,I1197946,I756162);
and I_70320 (I1197980,I1197782,I1197963);
nor I_70321 (I1197997,I1197895,I1197980);
DFFARX1 I_70322 (I1197997,I2507,I1197700,I1197668,);
DFFARX1 I_70323 (I1197980,I2507,I1197700,I1197689,);
nor I_70324 (I1198042,I756165,I756153);
nor I_70325 (I1197680,I1197895,I1198042);
or I_70326 (I1198073,I756165,I756153);
nor I_70327 (I1198090,I756144,I756147);
DFFARX1 I_70328 (I1198090,I2507,I1197700,I1198116,);
not I_70329 (I1198124,I1198116);
nor I_70330 (I1197686,I1198124,I1197929);
nand I_70331 (I1198155,I1198124,I1197774);
not I_70332 (I1198172,I756144);
nand I_70333 (I1198189,I1198172,I1197878);
nand I_70334 (I1198206,I1198124,I1198189);
nand I_70335 (I1197677,I1198206,I1198155);
nand I_70336 (I1197674,I1198189,I1198073);
not I_70337 (I1198278,I2514);
DFFARX1 I_70338 (I1250423,I2507,I1198278,I1198304,);
and I_70339 (I1198312,I1198304,I1250417);
DFFARX1 I_70340 (I1198312,I2507,I1198278,I1198261,);
DFFARX1 I_70341 (I1250402,I2507,I1198278,I1198352,);
not I_70342 (I1198360,I1250408);
not I_70343 (I1198377,I1250420);
nand I_70344 (I1198394,I1198377,I1198360);
nor I_70345 (I1198249,I1198352,I1198394);
DFFARX1 I_70346 (I1198394,I2507,I1198278,I1198434,);
not I_70347 (I1198270,I1198434);
not I_70348 (I1198456,I1250402);
nand I_70349 (I1198473,I1198377,I1198456);
DFFARX1 I_70350 (I1198473,I2507,I1198278,I1198499,);
not I_70351 (I1198507,I1198499);
not I_70352 (I1198524,I1250426);
nand I_70353 (I1198541,I1198524,I1250414);
and I_70354 (I1198558,I1198360,I1198541);
nor I_70355 (I1198575,I1198473,I1198558);
DFFARX1 I_70356 (I1198575,I2507,I1198278,I1198246,);
DFFARX1 I_70357 (I1198558,I2507,I1198278,I1198267,);
nor I_70358 (I1198620,I1250426,I1250405);
nor I_70359 (I1198258,I1198473,I1198620);
or I_70360 (I1198651,I1250426,I1250405);
nor I_70361 (I1198668,I1250411,I1250405);
DFFARX1 I_70362 (I1198668,I2507,I1198278,I1198694,);
not I_70363 (I1198702,I1198694);
nor I_70364 (I1198264,I1198702,I1198507);
nand I_70365 (I1198733,I1198702,I1198352);
not I_70366 (I1198750,I1250411);
nand I_70367 (I1198767,I1198750,I1198456);
nand I_70368 (I1198784,I1198702,I1198767);
nand I_70369 (I1198255,I1198784,I1198733);
nand I_70370 (I1198252,I1198767,I1198651);
not I_70371 (I1198856,I2514);
DFFARX1 I_70372 (I137735,I2507,I1198856,I1198882,);
and I_70373 (I1198890,I1198882,I137759);
DFFARX1 I_70374 (I1198890,I2507,I1198856,I1198839,);
DFFARX1 I_70375 (I137735,I2507,I1198856,I1198930,);
not I_70376 (I1198938,I137753);
not I_70377 (I1198955,I137738);
nand I_70378 (I1198972,I1198955,I1198938);
nor I_70379 (I1198827,I1198930,I1198972);
DFFARX1 I_70380 (I1198972,I2507,I1198856,I1199012,);
not I_70381 (I1198848,I1199012);
not I_70382 (I1199034,I137747);
nand I_70383 (I1199051,I1198955,I1199034);
DFFARX1 I_70384 (I1199051,I2507,I1198856,I1199077,);
not I_70385 (I1199085,I1199077);
not I_70386 (I1199102,I137744);
nand I_70387 (I1199119,I1199102,I137741);
and I_70388 (I1199136,I1198938,I1199119);
nor I_70389 (I1199153,I1199051,I1199136);
DFFARX1 I_70390 (I1199153,I2507,I1198856,I1198824,);
DFFARX1 I_70391 (I1199136,I2507,I1198856,I1198845,);
nor I_70392 (I1199198,I137744,I137750);
nor I_70393 (I1198836,I1199051,I1199198);
or I_70394 (I1199229,I137744,I137750);
nor I_70395 (I1199246,I137756,I137762);
DFFARX1 I_70396 (I1199246,I2507,I1198856,I1199272,);
not I_70397 (I1199280,I1199272);
nor I_70398 (I1198842,I1199280,I1199085);
nand I_70399 (I1199311,I1199280,I1198930);
not I_70400 (I1199328,I137756);
nand I_70401 (I1199345,I1199328,I1199034);
nand I_70402 (I1199362,I1199280,I1199345);
nand I_70403 (I1198833,I1199362,I1199311);
nand I_70404 (I1198830,I1199345,I1199229);
not I_70405 (I1199434,I2514);
DFFARX1 I_70406 (I13754,I2507,I1199434,I1199460,);
and I_70407 (I1199468,I1199460,I13757);
DFFARX1 I_70408 (I1199468,I2507,I1199434,I1199417,);
DFFARX1 I_70409 (I13757,I2507,I1199434,I1199508,);
not I_70410 (I1199516,I13760);
not I_70411 (I1199533,I13775);
nand I_70412 (I1199550,I1199533,I1199516);
nor I_70413 (I1199405,I1199508,I1199550);
DFFARX1 I_70414 (I1199550,I2507,I1199434,I1199590,);
not I_70415 (I1199426,I1199590);
not I_70416 (I1199612,I13769);
nand I_70417 (I1199629,I1199533,I1199612);
DFFARX1 I_70418 (I1199629,I2507,I1199434,I1199655,);
not I_70419 (I1199663,I1199655);
not I_70420 (I1199680,I13772);
nand I_70421 (I1199697,I1199680,I13754);
and I_70422 (I1199714,I1199516,I1199697);
nor I_70423 (I1199731,I1199629,I1199714);
DFFARX1 I_70424 (I1199731,I2507,I1199434,I1199402,);
DFFARX1 I_70425 (I1199714,I2507,I1199434,I1199423,);
nor I_70426 (I1199776,I13772,I13766);
nor I_70427 (I1199414,I1199629,I1199776);
or I_70428 (I1199807,I13772,I13766);
nor I_70429 (I1199824,I13763,I13778);
DFFARX1 I_70430 (I1199824,I2507,I1199434,I1199850,);
not I_70431 (I1199858,I1199850);
nor I_70432 (I1199420,I1199858,I1199663);
nand I_70433 (I1199889,I1199858,I1199508);
not I_70434 (I1199906,I13763);
nand I_70435 (I1199923,I1199906,I1199612);
nand I_70436 (I1199940,I1199858,I1199923);
nand I_70437 (I1199411,I1199940,I1199889);
nand I_70438 (I1199408,I1199923,I1199807);
not I_70439 (I1200012,I2514);
DFFARX1 I_70440 (I1346394,I2507,I1200012,I1200038,);
and I_70441 (I1200046,I1200038,I1346376);
DFFARX1 I_70442 (I1200046,I2507,I1200012,I1199995,);
DFFARX1 I_70443 (I1346367,I2507,I1200012,I1200086,);
not I_70444 (I1200094,I1346382);
not I_70445 (I1200111,I1346370);
nand I_70446 (I1200128,I1200111,I1200094);
nor I_70447 (I1199983,I1200086,I1200128);
DFFARX1 I_70448 (I1200128,I2507,I1200012,I1200168,);
not I_70449 (I1200004,I1200168);
not I_70450 (I1200190,I1346379);
nand I_70451 (I1200207,I1200111,I1200190);
DFFARX1 I_70452 (I1200207,I2507,I1200012,I1200233,);
not I_70453 (I1200241,I1200233);
not I_70454 (I1200258,I1346388);
nand I_70455 (I1200275,I1200258,I1346367);
and I_70456 (I1200292,I1200094,I1200275);
nor I_70457 (I1200309,I1200207,I1200292);
DFFARX1 I_70458 (I1200309,I2507,I1200012,I1199980,);
DFFARX1 I_70459 (I1200292,I2507,I1200012,I1200001,);
nor I_70460 (I1200354,I1346388,I1346391);
nor I_70461 (I1199992,I1200207,I1200354);
or I_70462 (I1200385,I1346388,I1346391);
nor I_70463 (I1200402,I1346385,I1346373);
DFFARX1 I_70464 (I1200402,I2507,I1200012,I1200428,);
not I_70465 (I1200436,I1200428);
nor I_70466 (I1199998,I1200436,I1200241);
nand I_70467 (I1200467,I1200436,I1200086);
not I_70468 (I1200484,I1346385);
nand I_70469 (I1200501,I1200484,I1200190);
nand I_70470 (I1200518,I1200436,I1200501);
nand I_70471 (I1199989,I1200518,I1200467);
nand I_70472 (I1199986,I1200501,I1200385);
not I_70473 (I1200590,I2514);
DFFARX1 I_70474 (I438703,I2507,I1200590,I1200616,);
and I_70475 (I1200624,I1200616,I438718);
DFFARX1 I_70476 (I1200624,I2507,I1200590,I1200573,);
DFFARX1 I_70477 (I438721,I2507,I1200590,I1200664,);
not I_70478 (I1200672,I438715);
not I_70479 (I1200689,I438730);
nand I_70480 (I1200706,I1200689,I1200672);
nor I_70481 (I1200561,I1200664,I1200706);
DFFARX1 I_70482 (I1200706,I2507,I1200590,I1200746,);
not I_70483 (I1200582,I1200746);
not I_70484 (I1200768,I438706);
nand I_70485 (I1200785,I1200689,I1200768);
DFFARX1 I_70486 (I1200785,I2507,I1200590,I1200811,);
not I_70487 (I1200819,I1200811);
not I_70488 (I1200836,I438709);
nand I_70489 (I1200853,I1200836,I438703);
and I_70490 (I1200870,I1200672,I1200853);
nor I_70491 (I1200887,I1200785,I1200870);
DFFARX1 I_70492 (I1200887,I2507,I1200590,I1200558,);
DFFARX1 I_70493 (I1200870,I2507,I1200590,I1200579,);
nor I_70494 (I1200932,I438709,I438712);
nor I_70495 (I1200570,I1200785,I1200932);
or I_70496 (I1200963,I438709,I438712);
nor I_70497 (I1200980,I438727,I438724);
DFFARX1 I_70498 (I1200980,I2507,I1200590,I1201006,);
not I_70499 (I1201014,I1201006);
nor I_70500 (I1200576,I1201014,I1200819);
nand I_70501 (I1201045,I1201014,I1200664);
not I_70502 (I1201062,I438727);
nand I_70503 (I1201079,I1201062,I1200768);
nand I_70504 (I1201096,I1201014,I1201079);
nand I_70505 (I1200567,I1201096,I1201045);
nand I_70506 (I1200564,I1201079,I1200963);
not I_70507 (I1201168,I2514);
DFFARX1 I_70508 (I1210167,I2507,I1201168,I1201194,);
and I_70509 (I1201202,I1201194,I1210161);
DFFARX1 I_70510 (I1201202,I2507,I1201168,I1201151,);
DFFARX1 I_70511 (I1210146,I2507,I1201168,I1201242,);
not I_70512 (I1201250,I1210152);
not I_70513 (I1201267,I1210164);
nand I_70514 (I1201284,I1201267,I1201250);
nor I_70515 (I1201139,I1201242,I1201284);
DFFARX1 I_70516 (I1201284,I2507,I1201168,I1201324,);
not I_70517 (I1201160,I1201324);
not I_70518 (I1201346,I1210146);
nand I_70519 (I1201363,I1201267,I1201346);
DFFARX1 I_70520 (I1201363,I2507,I1201168,I1201389,);
not I_70521 (I1201397,I1201389);
not I_70522 (I1201414,I1210170);
nand I_70523 (I1201431,I1201414,I1210158);
and I_70524 (I1201448,I1201250,I1201431);
nor I_70525 (I1201465,I1201363,I1201448);
DFFARX1 I_70526 (I1201465,I2507,I1201168,I1201136,);
DFFARX1 I_70527 (I1201448,I2507,I1201168,I1201157,);
nor I_70528 (I1201510,I1210170,I1210149);
nor I_70529 (I1201148,I1201363,I1201510);
or I_70530 (I1201541,I1210170,I1210149);
nor I_70531 (I1201558,I1210155,I1210149);
DFFARX1 I_70532 (I1201558,I2507,I1201168,I1201584,);
not I_70533 (I1201592,I1201584);
nor I_70534 (I1201154,I1201592,I1201397);
nand I_70535 (I1201623,I1201592,I1201242);
not I_70536 (I1201640,I1210155);
nand I_70537 (I1201657,I1201640,I1201346);
nand I_70538 (I1201674,I1201592,I1201657);
nand I_70539 (I1201145,I1201674,I1201623);
nand I_70540 (I1201142,I1201657,I1201541);
not I_70541 (I1201746,I2514);
DFFARX1 I_70542 (I491471,I2507,I1201746,I1201772,);
and I_70543 (I1201780,I1201772,I491486);
DFFARX1 I_70544 (I1201780,I2507,I1201746,I1201729,);
DFFARX1 I_70545 (I491489,I2507,I1201746,I1201820,);
not I_70546 (I1201828,I491483);
not I_70547 (I1201845,I491498);
nand I_70548 (I1201862,I1201845,I1201828);
nor I_70549 (I1201717,I1201820,I1201862);
DFFARX1 I_70550 (I1201862,I2507,I1201746,I1201902,);
not I_70551 (I1201738,I1201902);
not I_70552 (I1201924,I491474);
nand I_70553 (I1201941,I1201845,I1201924);
DFFARX1 I_70554 (I1201941,I2507,I1201746,I1201967,);
not I_70555 (I1201975,I1201967);
not I_70556 (I1201992,I491477);
nand I_70557 (I1202009,I1201992,I491471);
and I_70558 (I1202026,I1201828,I1202009);
nor I_70559 (I1202043,I1201941,I1202026);
DFFARX1 I_70560 (I1202043,I2507,I1201746,I1201714,);
DFFARX1 I_70561 (I1202026,I2507,I1201746,I1201735,);
nor I_70562 (I1202088,I491477,I491480);
nor I_70563 (I1201726,I1201941,I1202088);
or I_70564 (I1202119,I491477,I491480);
nor I_70565 (I1202136,I491495,I491492);
DFFARX1 I_70566 (I1202136,I2507,I1201746,I1202162,);
not I_70567 (I1202170,I1202162);
nor I_70568 (I1201732,I1202170,I1201975);
nand I_70569 (I1202201,I1202170,I1201820);
not I_70570 (I1202218,I491495);
nand I_70571 (I1202235,I1202218,I1201924);
nand I_70572 (I1202252,I1202170,I1202235);
nand I_70573 (I1201723,I1202252,I1202201);
nand I_70574 (I1201720,I1202235,I1202119);
not I_70575 (I1202324,I2514);
DFFARX1 I_70576 (I730149,I2507,I1202324,I1202350,);
and I_70577 (I1202358,I1202350,I730137);
DFFARX1 I_70578 (I1202358,I2507,I1202324,I1202307,);
DFFARX1 I_70579 (I730140,I2507,I1202324,I1202398,);
not I_70580 (I1202406,I730134);
not I_70581 (I1202423,I730158);
nand I_70582 (I1202440,I1202423,I1202406);
nor I_70583 (I1202295,I1202398,I1202440);
DFFARX1 I_70584 (I1202440,I2507,I1202324,I1202480,);
not I_70585 (I1202316,I1202480);
not I_70586 (I1202502,I730146);
nand I_70587 (I1202519,I1202423,I1202502);
DFFARX1 I_70588 (I1202519,I2507,I1202324,I1202545,);
not I_70589 (I1202553,I1202545);
not I_70590 (I1202570,I730155);
nand I_70591 (I1202587,I1202570,I730152);
and I_70592 (I1202604,I1202406,I1202587);
nor I_70593 (I1202621,I1202519,I1202604);
DFFARX1 I_70594 (I1202621,I2507,I1202324,I1202292,);
DFFARX1 I_70595 (I1202604,I2507,I1202324,I1202313,);
nor I_70596 (I1202666,I730155,I730143);
nor I_70597 (I1202304,I1202519,I1202666);
or I_70598 (I1202697,I730155,I730143);
nor I_70599 (I1202714,I730134,I730137);
DFFARX1 I_70600 (I1202714,I2507,I1202324,I1202740,);
not I_70601 (I1202748,I1202740);
nor I_70602 (I1202310,I1202748,I1202553);
nand I_70603 (I1202779,I1202748,I1202398);
not I_70604 (I1202796,I730134);
nand I_70605 (I1202813,I1202796,I1202502);
nand I_70606 (I1202830,I1202748,I1202813);
nand I_70607 (I1202301,I1202830,I1202779);
nand I_70608 (I1202298,I1202813,I1202697);
not I_70609 (I1202902,I2514);
DFFARX1 I_70610 (I330848,I2507,I1202902,I1202928,);
and I_70611 (I1202936,I1202928,I330833);
DFFARX1 I_70612 (I1202936,I2507,I1202902,I1202885,);
DFFARX1 I_70613 (I330839,I2507,I1202902,I1202976,);
not I_70614 (I1202984,I330821);
not I_70615 (I1203001,I330842);
nand I_70616 (I1203018,I1203001,I1202984);
nor I_70617 (I1202873,I1202976,I1203018);
DFFARX1 I_70618 (I1203018,I2507,I1202902,I1203058,);
not I_70619 (I1202894,I1203058);
not I_70620 (I1203080,I330845);
nand I_70621 (I1203097,I1203001,I1203080);
DFFARX1 I_70622 (I1203097,I2507,I1202902,I1203123,);
not I_70623 (I1203131,I1203123);
not I_70624 (I1203148,I330836);
nand I_70625 (I1203165,I1203148,I330824);
and I_70626 (I1203182,I1202984,I1203165);
nor I_70627 (I1203199,I1203097,I1203182);
DFFARX1 I_70628 (I1203199,I2507,I1202902,I1202870,);
DFFARX1 I_70629 (I1203182,I2507,I1202902,I1202891,);
nor I_70630 (I1203244,I330836,I330830);
nor I_70631 (I1202882,I1203097,I1203244);
or I_70632 (I1203275,I330836,I330830);
nor I_70633 (I1203292,I330827,I330821);
DFFARX1 I_70634 (I1203292,I2507,I1202902,I1203318,);
not I_70635 (I1203326,I1203318);
nor I_70636 (I1202888,I1203326,I1203131);
nand I_70637 (I1203357,I1203326,I1202976);
not I_70638 (I1203374,I330827);
nand I_70639 (I1203391,I1203374,I1203080);
nand I_70640 (I1203408,I1203326,I1203391);
nand I_70641 (I1202879,I1203408,I1203357);
nand I_70642 (I1202876,I1203391,I1203275);
not I_70643 (I1203480,I2514);
DFFARX1 I_70644 (I892745,I2507,I1203480,I1203506,);
and I_70645 (I1203514,I1203506,I892739);
DFFARX1 I_70646 (I1203514,I2507,I1203480,I1203463,);
DFFARX1 I_70647 (I892757,I2507,I1203480,I1203554,);
not I_70648 (I1203562,I892748);
not I_70649 (I1203579,I892760);
nand I_70650 (I1203596,I1203579,I1203562);
nor I_70651 (I1203451,I1203554,I1203596);
DFFARX1 I_70652 (I1203596,I2507,I1203480,I1203636,);
not I_70653 (I1203472,I1203636);
not I_70654 (I1203658,I892766);
nand I_70655 (I1203675,I1203579,I1203658);
DFFARX1 I_70656 (I1203675,I2507,I1203480,I1203701,);
not I_70657 (I1203709,I1203701);
not I_70658 (I1203726,I892742);
nand I_70659 (I1203743,I1203726,I892763);
and I_70660 (I1203760,I1203562,I1203743);
nor I_70661 (I1203777,I1203675,I1203760);
DFFARX1 I_70662 (I1203777,I2507,I1203480,I1203448,);
DFFARX1 I_70663 (I1203760,I2507,I1203480,I1203469,);
nor I_70664 (I1203822,I892742,I892754);
nor I_70665 (I1203460,I1203675,I1203822);
or I_70666 (I1203853,I892742,I892754);
nor I_70667 (I1203870,I892739,I892751);
DFFARX1 I_70668 (I1203870,I2507,I1203480,I1203896,);
not I_70669 (I1203904,I1203896);
nor I_70670 (I1203466,I1203904,I1203709);
nand I_70671 (I1203935,I1203904,I1203554);
not I_70672 (I1203952,I892739);
nand I_70673 (I1203969,I1203952,I1203658);
nand I_70674 (I1203986,I1203904,I1203969);
nand I_70675 (I1203457,I1203986,I1203935);
nand I_70676 (I1203454,I1203969,I1203853);
not I_70677 (I1204058,I2514);
DFFARX1 I_70678 (I64370,I2507,I1204058,I1204084,);
and I_70679 (I1204092,I1204084,I64346);
DFFARX1 I_70680 (I1204092,I2507,I1204058,I1204041,);
DFFARX1 I_70681 (I64364,I2507,I1204058,I1204132,);
not I_70682 (I1204140,I64352);
not I_70683 (I1204157,I64349);
nand I_70684 (I1204174,I1204157,I1204140);
nor I_70685 (I1204029,I1204132,I1204174);
DFFARX1 I_70686 (I1204174,I2507,I1204058,I1204214,);
not I_70687 (I1204050,I1204214);
not I_70688 (I1204236,I64358);
nand I_70689 (I1204253,I1204157,I1204236);
DFFARX1 I_70690 (I1204253,I2507,I1204058,I1204279,);
not I_70691 (I1204287,I1204279);
not I_70692 (I1204304,I64349);
nand I_70693 (I1204321,I1204304,I64367);
and I_70694 (I1204338,I1204140,I1204321);
nor I_70695 (I1204355,I1204253,I1204338);
DFFARX1 I_70696 (I1204355,I2507,I1204058,I1204026,);
DFFARX1 I_70697 (I1204338,I2507,I1204058,I1204047,);
nor I_70698 (I1204400,I64349,I64361);
nor I_70699 (I1204038,I1204253,I1204400);
or I_70700 (I1204431,I64349,I64361);
nor I_70701 (I1204448,I64355,I64346);
DFFARX1 I_70702 (I1204448,I2507,I1204058,I1204474,);
not I_70703 (I1204482,I1204474);
nor I_70704 (I1204044,I1204482,I1204287);
nand I_70705 (I1204513,I1204482,I1204132);
not I_70706 (I1204530,I64355);
nand I_70707 (I1204547,I1204530,I1204236);
nand I_70708 (I1204564,I1204482,I1204547);
nand I_70709 (I1204035,I1204564,I1204513);
nand I_70710 (I1204032,I1204547,I1204431);
not I_70711 (I1204636,I2514);
DFFARX1 I_70712 (I840195,I2507,I1204636,I1204662,);
and I_70713 (I1204670,I1204662,I840201);
DFFARX1 I_70714 (I1204670,I2507,I1204636,I1204619,);
DFFARX1 I_70715 (I840207,I2507,I1204636,I1204710,);
not I_70716 (I1204718,I840192);
not I_70717 (I1204735,I840192);
nand I_70718 (I1204752,I1204735,I1204718);
nor I_70719 (I1204607,I1204710,I1204752);
DFFARX1 I_70720 (I1204752,I2507,I1204636,I1204792,);
not I_70721 (I1204628,I1204792);
not I_70722 (I1204814,I840210);
nand I_70723 (I1204831,I1204735,I1204814);
DFFARX1 I_70724 (I1204831,I2507,I1204636,I1204857,);
not I_70725 (I1204865,I1204857);
not I_70726 (I1204882,I840204);
nand I_70727 (I1204899,I1204882,I840195);
and I_70728 (I1204916,I1204718,I1204899);
nor I_70729 (I1204933,I1204831,I1204916);
DFFARX1 I_70730 (I1204933,I2507,I1204636,I1204604,);
DFFARX1 I_70731 (I1204916,I2507,I1204636,I1204625,);
nor I_70732 (I1204978,I840204,I840213);
nor I_70733 (I1204616,I1204831,I1204978);
or I_70734 (I1205009,I840204,I840213);
nor I_70735 (I1205026,I840198,I840198);
DFFARX1 I_70736 (I1205026,I2507,I1204636,I1205052,);
not I_70737 (I1205060,I1205052);
nor I_70738 (I1204622,I1205060,I1204865);
nand I_70739 (I1205091,I1205060,I1204710);
not I_70740 (I1205108,I840198);
nand I_70741 (I1205125,I1205108,I1204814);
nand I_70742 (I1205142,I1205060,I1205125);
nand I_70743 (I1204613,I1205142,I1205091);
nand I_70744 (I1204610,I1205125,I1205009);
not I_70745 (I1205214,I2514);
DFFARX1 I_70746 (I1253143,I2507,I1205214,I1205240,);
and I_70747 (I1205248,I1205240,I1253137);
DFFARX1 I_70748 (I1205248,I2507,I1205214,I1205197,);
DFFARX1 I_70749 (I1253122,I2507,I1205214,I1205288,);
not I_70750 (I1205296,I1253128);
not I_70751 (I1205313,I1253140);
nand I_70752 (I1205330,I1205313,I1205296);
nor I_70753 (I1205185,I1205288,I1205330);
DFFARX1 I_70754 (I1205330,I2507,I1205214,I1205370,);
not I_70755 (I1205206,I1205370);
not I_70756 (I1205392,I1253122);
nand I_70757 (I1205409,I1205313,I1205392);
DFFARX1 I_70758 (I1205409,I2507,I1205214,I1205435,);
not I_70759 (I1205443,I1205435);
not I_70760 (I1205460,I1253146);
nand I_70761 (I1205477,I1205460,I1253134);
and I_70762 (I1205494,I1205296,I1205477);
nor I_70763 (I1205511,I1205409,I1205494);
DFFARX1 I_70764 (I1205511,I2507,I1205214,I1205182,);
DFFARX1 I_70765 (I1205494,I2507,I1205214,I1205203,);
nor I_70766 (I1205556,I1253146,I1253125);
nor I_70767 (I1205194,I1205409,I1205556);
or I_70768 (I1205587,I1253146,I1253125);
nor I_70769 (I1205604,I1253131,I1253125);
DFFARX1 I_70770 (I1205604,I2507,I1205214,I1205630,);
not I_70771 (I1205638,I1205630);
nor I_70772 (I1205200,I1205638,I1205443);
nand I_70773 (I1205669,I1205638,I1205288);
not I_70774 (I1205686,I1253131);
nand I_70775 (I1205703,I1205686,I1205392);
nand I_70776 (I1205720,I1205638,I1205703);
nand I_70777 (I1205191,I1205720,I1205669);
nand I_70778 (I1205188,I1205703,I1205587);
not I_70779 (I1205792,I2514);
DFFARX1 I_70780 (I398447,I2507,I1205792,I1205818,);
and I_70781 (I1205826,I1205818,I398462);
DFFARX1 I_70782 (I1205826,I2507,I1205792,I1205775,);
DFFARX1 I_70783 (I398465,I2507,I1205792,I1205866,);
not I_70784 (I1205874,I398459);
not I_70785 (I1205891,I398474);
nand I_70786 (I1205908,I1205891,I1205874);
nor I_70787 (I1205763,I1205866,I1205908);
DFFARX1 I_70788 (I1205908,I2507,I1205792,I1205948,);
not I_70789 (I1205784,I1205948);
not I_70790 (I1205970,I398450);
nand I_70791 (I1205987,I1205891,I1205970);
DFFARX1 I_70792 (I1205987,I2507,I1205792,I1206013,);
not I_70793 (I1206021,I1206013);
not I_70794 (I1206038,I398453);
nand I_70795 (I1206055,I1206038,I398447);
and I_70796 (I1206072,I1205874,I1206055);
nor I_70797 (I1206089,I1205987,I1206072);
DFFARX1 I_70798 (I1206089,I2507,I1205792,I1205760,);
DFFARX1 I_70799 (I1206072,I2507,I1205792,I1205781,);
nor I_70800 (I1206134,I398453,I398456);
nor I_70801 (I1205772,I1205987,I1206134);
or I_70802 (I1206165,I398453,I398456);
nor I_70803 (I1206182,I398471,I398468);
DFFARX1 I_70804 (I1206182,I2507,I1205792,I1206208,);
not I_70805 (I1206216,I1206208);
nor I_70806 (I1205778,I1206216,I1206021);
nand I_70807 (I1206247,I1206216,I1205866);
not I_70808 (I1206264,I398471);
nand I_70809 (I1206281,I1206264,I1205970);
nand I_70810 (I1206298,I1206216,I1206281);
nand I_70811 (I1205769,I1206298,I1206247);
nand I_70812 (I1205766,I1206281,I1206165);
not I_70813 (I1206370,I2514);
DFFARX1 I_70814 (I889509,I2507,I1206370,I1206396,);
nand I_70815 (I1206404,I1206396,I889509);
DFFARX1 I_70816 (I889521,I2507,I1206370,I1206430,);
DFFARX1 I_70817 (I1206430,I2507,I1206370,I1206447,);
not I_70818 (I1206362,I1206447);
not I_70819 (I1206469,I889515);
nor I_70820 (I1206486,I889515,I889536);
not I_70821 (I1206503,I889524);
nand I_70822 (I1206520,I1206469,I1206503);
nor I_70823 (I1206537,I889524,I889515);
and I_70824 (I1206341,I1206537,I1206404);
not I_70825 (I1206568,I889518);
nand I_70826 (I1206585,I1206568,I889533);
nor I_70827 (I1206602,I889518,I889527);
not I_70828 (I1206619,I1206602);
nand I_70829 (I1206344,I1206486,I1206619);
DFFARX1 I_70830 (I1206602,I2507,I1206370,I1206359,);
nor I_70831 (I1206664,I889530,I889524);
nor I_70832 (I1206681,I1206664,I889536);
and I_70833 (I1206698,I1206681,I1206585);
DFFARX1 I_70834 (I1206698,I2507,I1206370,I1206356,);
nor I_70835 (I1206353,I1206664,I1206520);
or I_70836 (I1206350,I1206602,I1206664);
nor I_70837 (I1206757,I889530,I889512);
DFFARX1 I_70838 (I1206757,I2507,I1206370,I1206783,);
not I_70839 (I1206791,I1206783);
nand I_70840 (I1206808,I1206791,I1206469);
nor I_70841 (I1206825,I1206808,I889536);
DFFARX1 I_70842 (I1206825,I2507,I1206370,I1206338,);
nor I_70843 (I1206856,I1206791,I1206520);
nor I_70844 (I1206347,I1206664,I1206856);
not I_70845 (I1206914,I2514);
DFFARX1 I_70846 (I1316049,I2507,I1206914,I1206940,);
nand I_70847 (I1206948,I1206940,I1316034);
DFFARX1 I_70848 (I1316028,I2507,I1206914,I1206974,);
DFFARX1 I_70849 (I1206974,I2507,I1206914,I1206991,);
not I_70850 (I1206906,I1206991);
not I_70851 (I1207013,I1316022);
nor I_70852 (I1207030,I1316022,I1316043);
not I_70853 (I1207047,I1316031);
nand I_70854 (I1207064,I1207013,I1207047);
nor I_70855 (I1207081,I1316031,I1316022);
and I_70856 (I1206885,I1207081,I1206948);
not I_70857 (I1207112,I1316040);
nand I_70858 (I1207129,I1207112,I1316046);
nor I_70859 (I1207146,I1316040,I1316037);
not I_70860 (I1207163,I1207146);
nand I_70861 (I1206888,I1207030,I1207163);
DFFARX1 I_70862 (I1207146,I2507,I1206914,I1206903,);
nor I_70863 (I1207208,I1316025,I1316031);
nor I_70864 (I1207225,I1207208,I1316043);
and I_70865 (I1207242,I1207225,I1207129);
DFFARX1 I_70866 (I1207242,I2507,I1206914,I1206900,);
nor I_70867 (I1206897,I1207208,I1207064);
or I_70868 (I1206894,I1207146,I1207208);
nor I_70869 (I1207301,I1316025,I1316022);
DFFARX1 I_70870 (I1207301,I2507,I1206914,I1207327,);
not I_70871 (I1207335,I1207327);
nand I_70872 (I1207352,I1207335,I1207013);
nor I_70873 (I1207369,I1207352,I1316043);
DFFARX1 I_70874 (I1207369,I2507,I1206914,I1206882,);
nor I_70875 (I1207400,I1207335,I1207064);
nor I_70876 (I1206891,I1207208,I1207400);
not I_70877 (I1207458,I2514);
DFFARX1 I_70878 (I29046,I2507,I1207458,I1207484,);
nand I_70879 (I1207492,I1207484,I29040);
DFFARX1 I_70880 (I29061,I2507,I1207458,I1207518,);
DFFARX1 I_70881 (I1207518,I2507,I1207458,I1207535,);
not I_70882 (I1207450,I1207535);
not I_70883 (I1207557,I29049);
nor I_70884 (I1207574,I29049,I29058);
not I_70885 (I1207591,I29037);
nand I_70886 (I1207608,I1207557,I1207591);
nor I_70887 (I1207625,I29037,I29049);
and I_70888 (I1207429,I1207625,I1207492);
not I_70889 (I1207656,I29055);
nand I_70890 (I1207673,I1207656,I29043);
nor I_70891 (I1207690,I29055,I29037);
not I_70892 (I1207707,I1207690);
nand I_70893 (I1207432,I1207574,I1207707);
DFFARX1 I_70894 (I1207690,I2507,I1207458,I1207447,);
nor I_70895 (I1207752,I29040,I29037);
nor I_70896 (I1207769,I1207752,I29058);
and I_70897 (I1207786,I1207769,I1207673);
DFFARX1 I_70898 (I1207786,I2507,I1207458,I1207444,);
nor I_70899 (I1207441,I1207752,I1207608);
or I_70900 (I1207438,I1207690,I1207752);
nor I_70901 (I1207845,I29040,I29052);
DFFARX1 I_70902 (I1207845,I2507,I1207458,I1207871,);
not I_70903 (I1207879,I1207871);
nand I_70904 (I1207896,I1207879,I1207557);
nor I_70905 (I1207913,I1207896,I29058);
DFFARX1 I_70906 (I1207913,I2507,I1207458,I1207426,);
nor I_70907 (I1207944,I1207879,I1207608);
nor I_70908 (I1207435,I1207752,I1207944);
not I_70909 (I1208002,I2514);
DFFARX1 I_70910 (I1369599,I2507,I1208002,I1208028,);
nand I_70911 (I1208036,I1208028,I1369584);
DFFARX1 I_70912 (I1369578,I2507,I1208002,I1208062,);
DFFARX1 I_70913 (I1208062,I2507,I1208002,I1208079,);
not I_70914 (I1207994,I1208079);
not I_70915 (I1208101,I1369572);
nor I_70916 (I1208118,I1369572,I1369593);
not I_70917 (I1208135,I1369581);
nand I_70918 (I1208152,I1208101,I1208135);
nor I_70919 (I1208169,I1369581,I1369572);
and I_70920 (I1207973,I1208169,I1208036);
not I_70921 (I1208200,I1369590);
nand I_70922 (I1208217,I1208200,I1369596);
nor I_70923 (I1208234,I1369590,I1369587);
not I_70924 (I1208251,I1208234);
nand I_70925 (I1207976,I1208118,I1208251);
DFFARX1 I_70926 (I1208234,I2507,I1208002,I1207991,);
nor I_70927 (I1208296,I1369575,I1369581);
nor I_70928 (I1208313,I1208296,I1369593);
and I_70929 (I1208330,I1208313,I1208217);
DFFARX1 I_70930 (I1208330,I2507,I1208002,I1207988,);
nor I_70931 (I1207985,I1208296,I1208152);
or I_70932 (I1207982,I1208234,I1208296);
nor I_70933 (I1208389,I1369575,I1369572);
DFFARX1 I_70934 (I1208389,I2507,I1208002,I1208415,);
not I_70935 (I1208423,I1208415);
nand I_70936 (I1208440,I1208423,I1208101);
nor I_70937 (I1208457,I1208440,I1369593);
DFFARX1 I_70938 (I1208457,I2507,I1208002,I1207970,);
nor I_70939 (I1208488,I1208423,I1208152);
nor I_70940 (I1207979,I1208296,I1208488);
not I_70941 (I1208546,I2514);
DFFARX1 I_70942 (I1154920,I2507,I1208546,I1208572,);
nand I_70943 (I1208580,I1208572,I1154899);
DFFARX1 I_70944 (I1154896,I2507,I1208546,I1208606,);
DFFARX1 I_70945 (I1208606,I2507,I1208546,I1208623,);
not I_70946 (I1208538,I1208623);
not I_70947 (I1208645,I1154908);
nor I_70948 (I1208662,I1154908,I1154917);
not I_70949 (I1208679,I1154905);
nand I_70950 (I1208696,I1208645,I1208679);
nor I_70951 (I1208713,I1154905,I1154908);
and I_70952 (I1208517,I1208713,I1208580);
not I_70953 (I1208744,I1154914);
nand I_70954 (I1208761,I1208744,I1154911);
nor I_70955 (I1208778,I1154914,I1154896);
not I_70956 (I1208795,I1208778);
nand I_70957 (I1208520,I1208662,I1208795);
DFFARX1 I_70958 (I1208778,I2507,I1208546,I1208535,);
nor I_70959 (I1208840,I1154899,I1154905);
nor I_70960 (I1208857,I1208840,I1154917);
and I_70961 (I1208874,I1208857,I1208761);
DFFARX1 I_70962 (I1208874,I2507,I1208546,I1208532,);
nor I_70963 (I1208529,I1208840,I1208696);
or I_70964 (I1208526,I1208778,I1208840);
nor I_70965 (I1208933,I1154899,I1154902);
DFFARX1 I_70966 (I1208933,I2507,I1208546,I1208959,);
not I_70967 (I1208967,I1208959);
nand I_70968 (I1208984,I1208967,I1208645);
nor I_70969 (I1209001,I1208984,I1154917);
DFFARX1 I_70970 (I1209001,I2507,I1208546,I1208514,);
nor I_70971 (I1209032,I1208967,I1208696);
nor I_70972 (I1208523,I1208840,I1209032);
not I_70973 (I1209090,I2514);
DFFARX1 I_70974 (I39059,I2507,I1209090,I1209116,);
nand I_70975 (I1209124,I1209116,I39053);
DFFARX1 I_70976 (I39074,I2507,I1209090,I1209150,);
DFFARX1 I_70977 (I1209150,I2507,I1209090,I1209167,);
not I_70978 (I1209082,I1209167);
not I_70979 (I1209189,I39062);
nor I_70980 (I1209206,I39062,I39071);
not I_70981 (I1209223,I39050);
nand I_70982 (I1209240,I1209189,I1209223);
nor I_70983 (I1209257,I39050,I39062);
and I_70984 (I1209061,I1209257,I1209124);
not I_70985 (I1209288,I39068);
nand I_70986 (I1209305,I1209288,I39056);
nor I_70987 (I1209322,I39068,I39050);
not I_70988 (I1209339,I1209322);
nand I_70989 (I1209064,I1209206,I1209339);
DFFARX1 I_70990 (I1209322,I2507,I1209090,I1209079,);
nor I_70991 (I1209384,I39053,I39050);
nor I_70992 (I1209401,I1209384,I39071);
and I_70993 (I1209418,I1209401,I1209305);
DFFARX1 I_70994 (I1209418,I2507,I1209090,I1209076,);
nor I_70995 (I1209073,I1209384,I1209240);
or I_70996 (I1209070,I1209322,I1209384);
nor I_70997 (I1209477,I39053,I39065);
DFFARX1 I_70998 (I1209477,I2507,I1209090,I1209503,);
not I_70999 (I1209511,I1209503);
nand I_71000 (I1209528,I1209511,I1209189);
nor I_71001 (I1209545,I1209528,I39071);
DFFARX1 I_71002 (I1209545,I2507,I1209090,I1209058,);
nor I_71003 (I1209576,I1209511,I1209240);
nor I_71004 (I1209067,I1209384,I1209576);
not I_71005 (I1209634,I2514);
DFFARX1 I_71006 (I613399,I2507,I1209634,I1209660,);
nand I_71007 (I1209668,I1209660,I613387);
DFFARX1 I_71008 (I613393,I2507,I1209634,I1209694,);
DFFARX1 I_71009 (I1209694,I2507,I1209634,I1209711,);
not I_71010 (I1209626,I1209711);
not I_71011 (I1209733,I613378);
nor I_71012 (I1209750,I613378,I613390);
not I_71013 (I1209767,I613381);
nand I_71014 (I1209784,I1209733,I1209767);
nor I_71015 (I1209801,I613381,I613378);
and I_71016 (I1209605,I1209801,I1209668);
not I_71017 (I1209832,I613396);
nand I_71018 (I1209849,I1209832,I613378);
nor I_71019 (I1209866,I613396,I613402);
not I_71020 (I1209883,I1209866);
nand I_71021 (I1209608,I1209750,I1209883);
DFFARX1 I_71022 (I1209866,I2507,I1209634,I1209623,);
nor I_71023 (I1209928,I613384,I613381);
nor I_71024 (I1209945,I1209928,I613390);
and I_71025 (I1209962,I1209945,I1209849);
DFFARX1 I_71026 (I1209962,I2507,I1209634,I1209620,);
nor I_71027 (I1209617,I1209928,I1209784);
or I_71028 (I1209614,I1209866,I1209928);
nor I_71029 (I1210021,I613384,I613381);
DFFARX1 I_71030 (I1210021,I2507,I1209634,I1210047,);
not I_71031 (I1210055,I1210047);
nand I_71032 (I1210072,I1210055,I1209733);
nor I_71033 (I1210089,I1210072,I613390);
DFFARX1 I_71034 (I1210089,I2507,I1209634,I1209602,);
nor I_71035 (I1210120,I1210055,I1209784);
nor I_71036 (I1209611,I1209928,I1210120);
not I_71037 (I1210178,I2514);
DFFARX1 I_71038 (I113905,I2507,I1210178,I1210204,);
nand I_71039 (I1210212,I1210204,I113887);
DFFARX1 I_71040 (I113884,I2507,I1210178,I1210238,);
DFFARX1 I_71041 (I1210238,I2507,I1210178,I1210255,);
not I_71042 (I1210170,I1210255);
not I_71043 (I1210277,I113902);
nor I_71044 (I1210294,I113902,I113896);
not I_71045 (I1210311,I113884);
nand I_71046 (I1210328,I1210277,I1210311);
nor I_71047 (I1210345,I113884,I113902);
and I_71048 (I1210149,I1210345,I1210212);
not I_71049 (I1210376,I113893);
nand I_71050 (I1210393,I1210376,I113899);
nor I_71051 (I1210410,I113893,I113887);
not I_71052 (I1210427,I1210410);
nand I_71053 (I1210152,I1210294,I1210427);
DFFARX1 I_71054 (I1210410,I2507,I1210178,I1210167,);
nor I_71055 (I1210472,I113890,I113884);
nor I_71056 (I1210489,I1210472,I113896);
and I_71057 (I1210506,I1210489,I1210393);
DFFARX1 I_71058 (I1210506,I2507,I1210178,I1210164,);
nor I_71059 (I1210161,I1210472,I1210328);
or I_71060 (I1210158,I1210410,I1210472);
nor I_71061 (I1210565,I113890,I113908);
DFFARX1 I_71062 (I1210565,I2507,I1210178,I1210591,);
not I_71063 (I1210599,I1210591);
nand I_71064 (I1210616,I1210599,I1210277);
nor I_71065 (I1210633,I1210616,I113896);
DFFARX1 I_71066 (I1210633,I2507,I1210178,I1210146,);
nor I_71067 (I1210664,I1210599,I1210328);
nor I_71068 (I1210155,I1210472,I1210664);
not I_71069 (I1210722,I2514);
DFFARX1 I_71070 (I207359,I2507,I1210722,I1210748,);
nand I_71071 (I1210756,I1210748,I207374);
DFFARX1 I_71072 (I207371,I2507,I1210722,I1210782,);
DFFARX1 I_71073 (I1210782,I2507,I1210722,I1210799,);
not I_71074 (I1210714,I1210799);
not I_71075 (I1210821,I207350);
nor I_71076 (I1210838,I207350,I207356);
not I_71077 (I1210855,I207362);
nand I_71078 (I1210872,I1210821,I1210855);
nor I_71079 (I1210889,I207362,I207350);
and I_71080 (I1210693,I1210889,I1210756);
not I_71081 (I1210920,I207368);
nand I_71082 (I1210937,I1210920,I207350);
nor I_71083 (I1210954,I207368,I207353);
not I_71084 (I1210971,I1210954);
nand I_71085 (I1210696,I1210838,I1210971);
DFFARX1 I_71086 (I1210954,I2507,I1210722,I1210711,);
nor I_71087 (I1211016,I207353,I207362);
nor I_71088 (I1211033,I1211016,I207356);
and I_71089 (I1211050,I1211033,I1210937);
DFFARX1 I_71090 (I1211050,I2507,I1210722,I1210708,);
nor I_71091 (I1210705,I1211016,I1210872);
or I_71092 (I1210702,I1210954,I1211016);
nor I_71093 (I1211109,I207353,I207365);
DFFARX1 I_71094 (I1211109,I2507,I1210722,I1211135,);
not I_71095 (I1211143,I1211135);
nand I_71096 (I1211160,I1211143,I1210821);
nor I_71097 (I1211177,I1211160,I207356);
DFFARX1 I_71098 (I1211177,I2507,I1210722,I1210690,);
nor I_71099 (I1211208,I1211143,I1210872);
nor I_71100 (I1210699,I1211016,I1211208);
not I_71101 (I1211266,I2514);
DFFARX1 I_71102 (I262323,I2507,I1211266,I1211292,);
nand I_71103 (I1211300,I1211292,I262326);
DFFARX1 I_71104 (I262320,I2507,I1211266,I1211326,);
DFFARX1 I_71105 (I1211326,I2507,I1211266,I1211343,);
not I_71106 (I1211258,I1211343);
not I_71107 (I1211365,I262329);
nor I_71108 (I1211382,I262329,I262314);
not I_71109 (I1211399,I262338);
nand I_71110 (I1211416,I1211365,I1211399);
nor I_71111 (I1211433,I262338,I262329);
and I_71112 (I1211237,I1211433,I1211300);
not I_71113 (I1211464,I262317);
nand I_71114 (I1211481,I1211464,I262335);
nor I_71115 (I1211498,I262317,I262311);
not I_71116 (I1211515,I1211498);
nand I_71117 (I1211240,I1211382,I1211515);
DFFARX1 I_71118 (I1211498,I2507,I1211266,I1211255,);
nor I_71119 (I1211560,I262332,I262338);
nor I_71120 (I1211577,I1211560,I262314);
and I_71121 (I1211594,I1211577,I1211481);
DFFARX1 I_71122 (I1211594,I2507,I1211266,I1211252,);
nor I_71123 (I1211249,I1211560,I1211416);
or I_71124 (I1211246,I1211498,I1211560);
nor I_71125 (I1211653,I262332,I262311);
DFFARX1 I_71126 (I1211653,I2507,I1211266,I1211679,);
not I_71127 (I1211687,I1211679);
nand I_71128 (I1211704,I1211687,I1211365);
nor I_71129 (I1211721,I1211704,I262314);
DFFARX1 I_71130 (I1211721,I2507,I1211266,I1211234,);
nor I_71131 (I1211752,I1211687,I1211416);
nor I_71132 (I1211243,I1211560,I1211752);
not I_71133 (I1211810,I2514);
DFFARX1 I_71134 (I690255,I2507,I1211810,I1211836,);
nand I_71135 (I1211844,I1211836,I690270);
DFFARX1 I_71136 (I690264,I2507,I1211810,I1211870,);
DFFARX1 I_71137 (I1211870,I2507,I1211810,I1211887,);
not I_71138 (I1211802,I1211887);
not I_71139 (I1211909,I690267);
nor I_71140 (I1211926,I690267,I690273);
not I_71141 (I1211943,I690255);
nand I_71142 (I1211960,I1211909,I1211943);
nor I_71143 (I1211977,I690255,I690267);
and I_71144 (I1211781,I1211977,I1211844);
not I_71145 (I1212008,I690252);
nand I_71146 (I1212025,I1212008,I690258);
nor I_71147 (I1212042,I690252,I690252);
not I_71148 (I1212059,I1212042);
nand I_71149 (I1211784,I1211926,I1212059);
DFFARX1 I_71150 (I1212042,I2507,I1211810,I1211799,);
nor I_71151 (I1212104,I690261,I690255);
nor I_71152 (I1212121,I1212104,I690273);
and I_71153 (I1212138,I1212121,I1212025);
DFFARX1 I_71154 (I1212138,I2507,I1211810,I1211796,);
nor I_71155 (I1211793,I1212104,I1211960);
or I_71156 (I1211790,I1212042,I1212104);
nor I_71157 (I1212197,I690261,I690276);
DFFARX1 I_71158 (I1212197,I2507,I1211810,I1212223,);
not I_71159 (I1212231,I1212223);
nand I_71160 (I1212248,I1212231,I1211909);
nor I_71161 (I1212265,I1212248,I690273);
DFFARX1 I_71162 (I1212265,I2507,I1211810,I1211778,);
nor I_71163 (I1212296,I1212231,I1211960);
nor I_71164 (I1211787,I1212104,I1212296);
not I_71165 (I1212354,I2514);
DFFARX1 I_71166 (I772331,I2507,I1212354,I1212380,);
nand I_71167 (I1212388,I1212380,I772346);
DFFARX1 I_71168 (I772340,I2507,I1212354,I1212414,);
DFFARX1 I_71169 (I1212414,I2507,I1212354,I1212431,);
not I_71170 (I1212346,I1212431);
not I_71171 (I1212453,I772343);
nor I_71172 (I1212470,I772343,I772349);
not I_71173 (I1212487,I772331);
nand I_71174 (I1212504,I1212453,I1212487);
nor I_71175 (I1212521,I772331,I772343);
and I_71176 (I1212325,I1212521,I1212388);
not I_71177 (I1212552,I772328);
nand I_71178 (I1212569,I1212552,I772334);
nor I_71179 (I1212586,I772328,I772328);
not I_71180 (I1212603,I1212586);
nand I_71181 (I1212328,I1212470,I1212603);
DFFARX1 I_71182 (I1212586,I2507,I1212354,I1212343,);
nor I_71183 (I1212648,I772337,I772331);
nor I_71184 (I1212665,I1212648,I772349);
and I_71185 (I1212682,I1212665,I1212569);
DFFARX1 I_71186 (I1212682,I2507,I1212354,I1212340,);
nor I_71187 (I1212337,I1212648,I1212504);
or I_71188 (I1212334,I1212586,I1212648);
nor I_71189 (I1212741,I772337,I772352);
DFFARX1 I_71190 (I1212741,I2507,I1212354,I1212767,);
not I_71191 (I1212775,I1212767);
nand I_71192 (I1212792,I1212775,I1212453);
nor I_71193 (I1212809,I1212792,I772349);
DFFARX1 I_71194 (I1212809,I2507,I1212354,I1212322,);
nor I_71195 (I1212840,I1212775,I1212504);
nor I_71196 (I1212331,I1212648,I1212840);
not I_71197 (I1212898,I2514);
DFFARX1 I_71198 (I700659,I2507,I1212898,I1212924,);
nand I_71199 (I1212932,I1212924,I700674);
DFFARX1 I_71200 (I700668,I2507,I1212898,I1212958,);
DFFARX1 I_71201 (I1212958,I2507,I1212898,I1212975,);
not I_71202 (I1212890,I1212975);
not I_71203 (I1212997,I700671);
nor I_71204 (I1213014,I700671,I700677);
not I_71205 (I1213031,I700659);
nand I_71206 (I1213048,I1212997,I1213031);
nor I_71207 (I1213065,I700659,I700671);
and I_71208 (I1212869,I1213065,I1212932);
not I_71209 (I1213096,I700656);
nand I_71210 (I1213113,I1213096,I700662);
nor I_71211 (I1213130,I700656,I700656);
not I_71212 (I1213147,I1213130);
nand I_71213 (I1212872,I1213014,I1213147);
DFFARX1 I_71214 (I1213130,I2507,I1212898,I1212887,);
nor I_71215 (I1213192,I700665,I700659);
nor I_71216 (I1213209,I1213192,I700677);
and I_71217 (I1213226,I1213209,I1213113);
DFFARX1 I_71218 (I1213226,I2507,I1212898,I1212884,);
nor I_71219 (I1212881,I1213192,I1213048);
or I_71220 (I1212878,I1213130,I1213192);
nor I_71221 (I1213285,I700665,I700680);
DFFARX1 I_71222 (I1213285,I2507,I1212898,I1213311,);
not I_71223 (I1213319,I1213311);
nand I_71224 (I1213336,I1213319,I1212997);
nor I_71225 (I1213353,I1213336,I700677);
DFFARX1 I_71226 (I1213353,I2507,I1212898,I1212866,);
nor I_71227 (I1213384,I1213319,I1213048);
nor I_71228 (I1212875,I1213192,I1213384);
not I_71229 (I1213442,I2514);
DFFARX1 I_71230 (I640547,I2507,I1213442,I1213468,);
nand I_71231 (I1213476,I1213468,I640562);
DFFARX1 I_71232 (I640556,I2507,I1213442,I1213502,);
DFFARX1 I_71233 (I1213502,I2507,I1213442,I1213519,);
not I_71234 (I1213434,I1213519);
not I_71235 (I1213541,I640559);
nor I_71236 (I1213558,I640559,I640565);
not I_71237 (I1213575,I640547);
nand I_71238 (I1213592,I1213541,I1213575);
nor I_71239 (I1213609,I640547,I640559);
and I_71240 (I1213413,I1213609,I1213476);
not I_71241 (I1213640,I640544);
nand I_71242 (I1213657,I1213640,I640550);
nor I_71243 (I1213674,I640544,I640544);
not I_71244 (I1213691,I1213674);
nand I_71245 (I1213416,I1213558,I1213691);
DFFARX1 I_71246 (I1213674,I2507,I1213442,I1213431,);
nor I_71247 (I1213736,I640553,I640547);
nor I_71248 (I1213753,I1213736,I640565);
and I_71249 (I1213770,I1213753,I1213657);
DFFARX1 I_71250 (I1213770,I2507,I1213442,I1213428,);
nor I_71251 (I1213425,I1213736,I1213592);
or I_71252 (I1213422,I1213674,I1213736);
nor I_71253 (I1213829,I640553,I640568);
DFFARX1 I_71254 (I1213829,I2507,I1213442,I1213855,);
not I_71255 (I1213863,I1213855);
nand I_71256 (I1213880,I1213863,I1213541);
nor I_71257 (I1213897,I1213880,I640565);
DFFARX1 I_71258 (I1213897,I2507,I1213442,I1213410,);
nor I_71259 (I1213928,I1213863,I1213592);
nor I_71260 (I1213419,I1213736,I1213928);
not I_71261 (I1213986,I2514);
DFFARX1 I_71262 (I1352344,I2507,I1213986,I1214012,);
nand I_71263 (I1214020,I1214012,I1352329);
DFFARX1 I_71264 (I1352323,I2507,I1213986,I1214046,);
DFFARX1 I_71265 (I1214046,I2507,I1213986,I1214063,);
not I_71266 (I1213978,I1214063);
not I_71267 (I1214085,I1352317);
nor I_71268 (I1214102,I1352317,I1352338);
not I_71269 (I1214119,I1352326);
nand I_71270 (I1214136,I1214085,I1214119);
nor I_71271 (I1214153,I1352326,I1352317);
and I_71272 (I1213957,I1214153,I1214020);
not I_71273 (I1214184,I1352335);
nand I_71274 (I1214201,I1214184,I1352341);
nor I_71275 (I1214218,I1352335,I1352332);
not I_71276 (I1214235,I1214218);
nand I_71277 (I1213960,I1214102,I1214235);
DFFARX1 I_71278 (I1214218,I2507,I1213986,I1213975,);
nor I_71279 (I1214280,I1352320,I1352326);
nor I_71280 (I1214297,I1214280,I1352338);
and I_71281 (I1214314,I1214297,I1214201);
DFFARX1 I_71282 (I1214314,I2507,I1213986,I1213972,);
nor I_71283 (I1213969,I1214280,I1214136);
or I_71284 (I1213966,I1214218,I1214280);
nor I_71285 (I1214373,I1352320,I1352317);
DFFARX1 I_71286 (I1214373,I2507,I1213986,I1214399,);
not I_71287 (I1214407,I1214399);
nand I_71288 (I1214424,I1214407,I1214085);
nor I_71289 (I1214441,I1214424,I1352338);
DFFARX1 I_71290 (I1214441,I2507,I1213986,I1213954,);
nor I_71291 (I1214472,I1214407,I1214136);
nor I_71292 (I1213963,I1214280,I1214472);
not I_71293 (I1214530,I2514);
DFFARX1 I_71294 (I368777,I2507,I1214530,I1214556,);
nand I_71295 (I1214564,I1214556,I368780);
DFFARX1 I_71296 (I368774,I2507,I1214530,I1214590,);
DFFARX1 I_71297 (I1214590,I2507,I1214530,I1214607,);
not I_71298 (I1214522,I1214607);
not I_71299 (I1214629,I368783);
nor I_71300 (I1214646,I368783,I368768);
not I_71301 (I1214663,I368792);
nand I_71302 (I1214680,I1214629,I1214663);
nor I_71303 (I1214697,I368792,I368783);
and I_71304 (I1214501,I1214697,I1214564);
not I_71305 (I1214728,I368771);
nand I_71306 (I1214745,I1214728,I368789);
nor I_71307 (I1214762,I368771,I368765);
not I_71308 (I1214779,I1214762);
nand I_71309 (I1214504,I1214646,I1214779);
DFFARX1 I_71310 (I1214762,I2507,I1214530,I1214519,);
nor I_71311 (I1214824,I368786,I368792);
nor I_71312 (I1214841,I1214824,I368768);
and I_71313 (I1214858,I1214841,I1214745);
DFFARX1 I_71314 (I1214858,I2507,I1214530,I1214516,);
nor I_71315 (I1214513,I1214824,I1214680);
or I_71316 (I1214510,I1214762,I1214824);
nor I_71317 (I1214917,I368786,I368765);
DFFARX1 I_71318 (I1214917,I2507,I1214530,I1214943,);
not I_71319 (I1214951,I1214943);
nand I_71320 (I1214968,I1214951,I1214629);
nor I_71321 (I1214985,I1214968,I368768);
DFFARX1 I_71322 (I1214985,I2507,I1214530,I1214498,);
nor I_71323 (I1215016,I1214951,I1214680);
nor I_71324 (I1214507,I1214824,I1215016);
not I_71325 (I1215074,I2514);
DFFARX1 I_71326 (I528599,I2507,I1215074,I1215100,);
nand I_71327 (I1215108,I1215100,I528623);
DFFARX1 I_71328 (I528602,I2507,I1215074,I1215134,);
DFFARX1 I_71329 (I1215134,I2507,I1215074,I1215151,);
not I_71330 (I1215066,I1215151);
not I_71331 (I1215173,I528605);
nor I_71332 (I1215190,I528605,I528620);
not I_71333 (I1215207,I528611);
nand I_71334 (I1215224,I1215173,I1215207);
nor I_71335 (I1215241,I528611,I528605);
and I_71336 (I1215045,I1215241,I1215108);
not I_71337 (I1215272,I528608);
nand I_71338 (I1215289,I1215272,I528602);
nor I_71339 (I1215306,I528608,I528617);
not I_71340 (I1215323,I1215306);
nand I_71341 (I1215048,I1215190,I1215323);
DFFARX1 I_71342 (I1215306,I2507,I1215074,I1215063,);
nor I_71343 (I1215368,I528614,I528611);
nor I_71344 (I1215385,I1215368,I528620);
and I_71345 (I1215402,I1215385,I1215289);
DFFARX1 I_71346 (I1215402,I2507,I1215074,I1215060,);
nor I_71347 (I1215057,I1215368,I1215224);
or I_71348 (I1215054,I1215306,I1215368);
nor I_71349 (I1215461,I528614,I528599);
DFFARX1 I_71350 (I1215461,I2507,I1215074,I1215487,);
not I_71351 (I1215495,I1215487);
nand I_71352 (I1215512,I1215495,I1215173);
nor I_71353 (I1215529,I1215512,I528620);
DFFARX1 I_71354 (I1215529,I2507,I1215074,I1215042,);
nor I_71355 (I1215560,I1215495,I1215224);
nor I_71356 (I1215051,I1215368,I1215560);
not I_71357 (I1215618,I2514);
DFFARX1 I_71358 (I668291,I2507,I1215618,I1215644,);
nand I_71359 (I1215652,I1215644,I668306);
DFFARX1 I_71360 (I668300,I2507,I1215618,I1215678,);
DFFARX1 I_71361 (I1215678,I2507,I1215618,I1215695,);
not I_71362 (I1215610,I1215695);
not I_71363 (I1215717,I668303);
nor I_71364 (I1215734,I668303,I668309);
not I_71365 (I1215751,I668291);
nand I_71366 (I1215768,I1215717,I1215751);
nor I_71367 (I1215785,I668291,I668303);
and I_71368 (I1215589,I1215785,I1215652);
not I_71369 (I1215816,I668288);
nand I_71370 (I1215833,I1215816,I668294);
nor I_71371 (I1215850,I668288,I668288);
not I_71372 (I1215867,I1215850);
nand I_71373 (I1215592,I1215734,I1215867);
DFFARX1 I_71374 (I1215850,I2507,I1215618,I1215607,);
nor I_71375 (I1215912,I668297,I668291);
nor I_71376 (I1215929,I1215912,I668309);
and I_71377 (I1215946,I1215929,I1215833);
DFFARX1 I_71378 (I1215946,I2507,I1215618,I1215604,);
nor I_71379 (I1215601,I1215912,I1215768);
or I_71380 (I1215598,I1215850,I1215912);
nor I_71381 (I1216005,I668297,I668312);
DFFARX1 I_71382 (I1216005,I2507,I1215618,I1216031,);
not I_71383 (I1216039,I1216031);
nand I_71384 (I1216056,I1216039,I1215717);
nor I_71385 (I1216073,I1216056,I668309);
DFFARX1 I_71386 (I1216073,I2507,I1215618,I1215586,);
nor I_71387 (I1216104,I1216039,I1215768);
nor I_71388 (I1215595,I1215912,I1216104);
not I_71389 (I1216162,I2514);
DFFARX1 I_71390 (I896615,I2507,I1216162,I1216188,);
nand I_71391 (I1216196,I1216188,I896615);
DFFARX1 I_71392 (I896627,I2507,I1216162,I1216222,);
DFFARX1 I_71393 (I1216222,I2507,I1216162,I1216239,);
not I_71394 (I1216154,I1216239);
not I_71395 (I1216261,I896621);
nor I_71396 (I1216278,I896621,I896642);
not I_71397 (I1216295,I896630);
nand I_71398 (I1216312,I1216261,I1216295);
nor I_71399 (I1216329,I896630,I896621);
and I_71400 (I1216133,I1216329,I1216196);
not I_71401 (I1216360,I896624);
nand I_71402 (I1216377,I1216360,I896639);
nor I_71403 (I1216394,I896624,I896633);
not I_71404 (I1216411,I1216394);
nand I_71405 (I1216136,I1216278,I1216411);
DFFARX1 I_71406 (I1216394,I2507,I1216162,I1216151,);
nor I_71407 (I1216456,I896636,I896630);
nor I_71408 (I1216473,I1216456,I896642);
and I_71409 (I1216490,I1216473,I1216377);
DFFARX1 I_71410 (I1216490,I2507,I1216162,I1216148,);
nor I_71411 (I1216145,I1216456,I1216312);
or I_71412 (I1216142,I1216394,I1216456);
nor I_71413 (I1216549,I896636,I896618);
DFFARX1 I_71414 (I1216549,I2507,I1216162,I1216575,);
not I_71415 (I1216583,I1216575);
nand I_71416 (I1216600,I1216583,I1216261);
nor I_71417 (I1216617,I1216600,I896642);
DFFARX1 I_71418 (I1216617,I2507,I1216162,I1216130,);
nor I_71419 (I1216648,I1216583,I1216312);
nor I_71420 (I1216139,I1216456,I1216648);
not I_71421 (I1216706,I2514);
DFFARX1 I_71422 (I868129,I2507,I1216706,I1216732,);
nand I_71423 (I1216740,I1216732,I868123);
DFFARX1 I_71424 (I868126,I2507,I1216706,I1216766,);
DFFARX1 I_71425 (I1216766,I2507,I1216706,I1216783,);
not I_71426 (I1216698,I1216783);
not I_71427 (I1216805,I868132);
nor I_71428 (I1216822,I868132,I868126);
not I_71429 (I1216839,I868135);
nand I_71430 (I1216856,I1216805,I1216839);
nor I_71431 (I1216873,I868135,I868132);
and I_71432 (I1216677,I1216873,I1216740);
not I_71433 (I1216904,I868144);
nand I_71434 (I1216921,I1216904,I868138);
nor I_71435 (I1216938,I868144,I868141);
not I_71436 (I1216955,I1216938);
nand I_71437 (I1216680,I1216822,I1216955);
DFFARX1 I_71438 (I1216938,I2507,I1216706,I1216695,);
nor I_71439 (I1217000,I868123,I868135);
nor I_71440 (I1217017,I1217000,I868126);
and I_71441 (I1217034,I1217017,I1216921);
DFFARX1 I_71442 (I1217034,I2507,I1216706,I1216692,);
nor I_71443 (I1216689,I1217000,I1216856);
or I_71444 (I1216686,I1216938,I1217000);
nor I_71445 (I1217093,I868123,I868129);
DFFARX1 I_71446 (I1217093,I2507,I1216706,I1217119,);
not I_71447 (I1217127,I1217119);
nand I_71448 (I1217144,I1217127,I1216805);
nor I_71449 (I1217161,I1217144,I868126);
DFFARX1 I_71450 (I1217161,I2507,I1216706,I1216674,);
nor I_71451 (I1217192,I1217127,I1216856);
nor I_71452 (I1216683,I1217000,I1217192);
not I_71453 (I1217250,I2514);
DFFARX1 I_71454 (I206764,I2507,I1217250,I1217276,);
nand I_71455 (I1217284,I1217276,I206779);
DFFARX1 I_71456 (I206776,I2507,I1217250,I1217310,);
DFFARX1 I_71457 (I1217310,I2507,I1217250,I1217327,);
not I_71458 (I1217242,I1217327);
not I_71459 (I1217349,I206755);
nor I_71460 (I1217366,I206755,I206761);
not I_71461 (I1217383,I206767);
nand I_71462 (I1217400,I1217349,I1217383);
nor I_71463 (I1217417,I206767,I206755);
and I_71464 (I1217221,I1217417,I1217284);
not I_71465 (I1217448,I206773);
nand I_71466 (I1217465,I1217448,I206755);
nor I_71467 (I1217482,I206773,I206758);
not I_71468 (I1217499,I1217482);
nand I_71469 (I1217224,I1217366,I1217499);
DFFARX1 I_71470 (I1217482,I2507,I1217250,I1217239,);
nor I_71471 (I1217544,I206758,I206767);
nor I_71472 (I1217561,I1217544,I206761);
and I_71473 (I1217578,I1217561,I1217465);
DFFARX1 I_71474 (I1217578,I2507,I1217250,I1217236,);
nor I_71475 (I1217233,I1217544,I1217400);
or I_71476 (I1217230,I1217482,I1217544);
nor I_71477 (I1217637,I206758,I206770);
DFFARX1 I_71478 (I1217637,I2507,I1217250,I1217663,);
not I_71479 (I1217671,I1217663);
nand I_71480 (I1217688,I1217671,I1217349);
nor I_71481 (I1217705,I1217688,I206761);
DFFARX1 I_71482 (I1217705,I2507,I1217250,I1217218,);
nor I_71483 (I1217736,I1217671,I1217400);
nor I_71484 (I1217227,I1217544,I1217736);
not I_71485 (I1217794,I2514);
DFFARX1 I_71486 (I1294067,I2507,I1217794,I1217820,);
nand I_71487 (I1217828,I1217820,I1294076);
DFFARX1 I_71488 (I1294079,I2507,I1217794,I1217854,);
DFFARX1 I_71489 (I1217854,I2507,I1217794,I1217871,);
not I_71490 (I1217786,I1217871);
not I_71491 (I1217893,I1294073);
nor I_71492 (I1217910,I1294073,I1294070);
not I_71493 (I1217927,I1294064);
nand I_71494 (I1217944,I1217893,I1217927);
nor I_71495 (I1217961,I1294064,I1294073);
and I_71496 (I1217765,I1217961,I1217828);
not I_71497 (I1217992,I1294061);
nand I_71498 (I1218009,I1217992,I1294058);
nor I_71499 (I1218026,I1294061,I1294058);
not I_71500 (I1218043,I1218026);
nand I_71501 (I1217768,I1217910,I1218043);
DFFARX1 I_71502 (I1218026,I2507,I1217794,I1217783,);
nor I_71503 (I1218088,I1294061,I1294064);
nor I_71504 (I1218105,I1218088,I1294070);
and I_71505 (I1218122,I1218105,I1218009);
DFFARX1 I_71506 (I1218122,I2507,I1217794,I1217780,);
nor I_71507 (I1217777,I1218088,I1217944);
or I_71508 (I1217774,I1218026,I1218088);
nor I_71509 (I1218181,I1294061,I1294082);
DFFARX1 I_71510 (I1218181,I2507,I1217794,I1218207,);
not I_71511 (I1218215,I1218207);
nand I_71512 (I1218232,I1218215,I1217893);
nor I_71513 (I1218249,I1218232,I1294070);
DFFARX1 I_71514 (I1218249,I2507,I1217794,I1217762,);
nor I_71515 (I1218280,I1218215,I1217944);
nor I_71516 (I1217771,I1218088,I1218280);
not I_71517 (I1218338,I2514);
DFFARX1 I_71518 (I1305934,I2507,I1218338,I1218364,);
nand I_71519 (I1218372,I1218364,I1305919);
DFFARX1 I_71520 (I1305913,I2507,I1218338,I1218398,);
DFFARX1 I_71521 (I1218398,I2507,I1218338,I1218415,);
not I_71522 (I1218330,I1218415);
not I_71523 (I1218437,I1305907);
nor I_71524 (I1218454,I1305907,I1305928);
not I_71525 (I1218471,I1305916);
nand I_71526 (I1218488,I1218437,I1218471);
nor I_71527 (I1218505,I1305916,I1305907);
and I_71528 (I1218309,I1218505,I1218372);
not I_71529 (I1218536,I1305925);
nand I_71530 (I1218553,I1218536,I1305931);
nor I_71531 (I1218570,I1305925,I1305922);
not I_71532 (I1218587,I1218570);
nand I_71533 (I1218312,I1218454,I1218587);
DFFARX1 I_71534 (I1218570,I2507,I1218338,I1218327,);
nor I_71535 (I1218632,I1305910,I1305916);
nor I_71536 (I1218649,I1218632,I1305928);
and I_71537 (I1218666,I1218649,I1218553);
DFFARX1 I_71538 (I1218666,I2507,I1218338,I1218324,);
nor I_71539 (I1218321,I1218632,I1218488);
or I_71540 (I1218318,I1218570,I1218632);
nor I_71541 (I1218725,I1305910,I1305907);
DFFARX1 I_71542 (I1218725,I2507,I1218338,I1218751,);
not I_71543 (I1218759,I1218751);
nand I_71544 (I1218776,I1218759,I1218437);
nor I_71545 (I1218793,I1218776,I1305928);
DFFARX1 I_71546 (I1218793,I2507,I1218338,I1218306,);
nor I_71547 (I1218824,I1218759,I1218488);
nor I_71548 (I1218315,I1218632,I1218824);
not I_71549 (I1218882,I2514);
DFFARX1 I_71550 (I338211,I2507,I1218882,I1218908,);
nand I_71551 (I1218916,I1218908,I338214);
DFFARX1 I_71552 (I338208,I2507,I1218882,I1218942,);
DFFARX1 I_71553 (I1218942,I2507,I1218882,I1218959,);
not I_71554 (I1218874,I1218959);
not I_71555 (I1218981,I338217);
nor I_71556 (I1218998,I338217,I338202);
not I_71557 (I1219015,I338226);
nand I_71558 (I1219032,I1218981,I1219015);
nor I_71559 (I1219049,I338226,I338217);
and I_71560 (I1218853,I1219049,I1218916);
not I_71561 (I1219080,I338205);
nand I_71562 (I1219097,I1219080,I338223);
nor I_71563 (I1219114,I338205,I338199);
not I_71564 (I1219131,I1219114);
nand I_71565 (I1218856,I1218998,I1219131);
DFFARX1 I_71566 (I1219114,I2507,I1218882,I1218871,);
nor I_71567 (I1219176,I338220,I338226);
nor I_71568 (I1219193,I1219176,I338202);
and I_71569 (I1219210,I1219193,I1219097);
DFFARX1 I_71570 (I1219210,I2507,I1218882,I1218868,);
nor I_71571 (I1218865,I1219176,I1219032);
or I_71572 (I1218862,I1219114,I1219176);
nor I_71573 (I1219269,I338220,I338199);
DFFARX1 I_71574 (I1219269,I2507,I1218882,I1219295,);
not I_71575 (I1219303,I1219295);
nand I_71576 (I1219320,I1219303,I1218981);
nor I_71577 (I1219337,I1219320,I338202);
DFFARX1 I_71578 (I1219337,I2507,I1218882,I1218850,);
nor I_71579 (I1219368,I1219303,I1219032);
nor I_71580 (I1218859,I1219176,I1219368);
not I_71581 (I1219426,I2514);
DFFARX1 I_71582 (I333468,I2507,I1219426,I1219452,);
nand I_71583 (I1219460,I1219452,I333471);
DFFARX1 I_71584 (I333465,I2507,I1219426,I1219486,);
DFFARX1 I_71585 (I1219486,I2507,I1219426,I1219503,);
not I_71586 (I1219418,I1219503);
not I_71587 (I1219525,I333474);
nor I_71588 (I1219542,I333474,I333459);
not I_71589 (I1219559,I333483);
nand I_71590 (I1219576,I1219525,I1219559);
nor I_71591 (I1219593,I333483,I333474);
and I_71592 (I1219397,I1219593,I1219460);
not I_71593 (I1219624,I333462);
nand I_71594 (I1219641,I1219624,I333480);
nor I_71595 (I1219658,I333462,I333456);
not I_71596 (I1219675,I1219658);
nand I_71597 (I1219400,I1219542,I1219675);
DFFARX1 I_71598 (I1219658,I2507,I1219426,I1219415,);
nor I_71599 (I1219720,I333477,I333483);
nor I_71600 (I1219737,I1219720,I333459);
and I_71601 (I1219754,I1219737,I1219641);
DFFARX1 I_71602 (I1219754,I2507,I1219426,I1219412,);
nor I_71603 (I1219409,I1219720,I1219576);
or I_71604 (I1219406,I1219658,I1219720);
nor I_71605 (I1219813,I333477,I333456);
DFFARX1 I_71606 (I1219813,I2507,I1219426,I1219839,);
not I_71607 (I1219847,I1219839);
nand I_71608 (I1219864,I1219847,I1219525);
nor I_71609 (I1219881,I1219864,I333459);
DFFARX1 I_71610 (I1219881,I2507,I1219426,I1219394,);
nor I_71611 (I1219912,I1219847,I1219576);
nor I_71612 (I1219403,I1219720,I1219912);
not I_71613 (I1219970,I2514);
DFFARX1 I_71614 (I733605,I2507,I1219970,I1219996,);
nand I_71615 (I1220004,I1219996,I733620);
DFFARX1 I_71616 (I733614,I2507,I1219970,I1220030,);
DFFARX1 I_71617 (I1220030,I2507,I1219970,I1220047,);
not I_71618 (I1219962,I1220047);
not I_71619 (I1220069,I733617);
nor I_71620 (I1220086,I733617,I733623);
not I_71621 (I1220103,I733605);
nand I_71622 (I1220120,I1220069,I1220103);
nor I_71623 (I1220137,I733605,I733617);
and I_71624 (I1219941,I1220137,I1220004);
not I_71625 (I1220168,I733602);
nand I_71626 (I1220185,I1220168,I733608);
nor I_71627 (I1220202,I733602,I733602);
not I_71628 (I1220219,I1220202);
nand I_71629 (I1219944,I1220086,I1220219);
DFFARX1 I_71630 (I1220202,I2507,I1219970,I1219959,);
nor I_71631 (I1220264,I733611,I733605);
nor I_71632 (I1220281,I1220264,I733623);
and I_71633 (I1220298,I1220281,I1220185);
DFFARX1 I_71634 (I1220298,I2507,I1219970,I1219956,);
nor I_71635 (I1219953,I1220264,I1220120);
or I_71636 (I1219950,I1220202,I1220264);
nor I_71637 (I1220357,I733611,I733626);
DFFARX1 I_71638 (I1220357,I2507,I1219970,I1220383,);
not I_71639 (I1220391,I1220383);
nand I_71640 (I1220408,I1220391,I1220069);
nor I_71641 (I1220425,I1220408,I733623);
DFFARX1 I_71642 (I1220425,I2507,I1219970,I1219938,);
nor I_71643 (I1220456,I1220391,I1220120);
nor I_71644 (I1219947,I1220264,I1220456);
not I_71645 (I1220514,I2514);
DFFARX1 I_71646 (I1270369,I2507,I1220514,I1220540,);
nand I_71647 (I1220548,I1220540,I1270378);
DFFARX1 I_71648 (I1270381,I2507,I1220514,I1220574,);
DFFARX1 I_71649 (I1220574,I2507,I1220514,I1220591,);
not I_71650 (I1220506,I1220591);
not I_71651 (I1220613,I1270375);
nor I_71652 (I1220630,I1270375,I1270372);
not I_71653 (I1220647,I1270366);
nand I_71654 (I1220664,I1220613,I1220647);
nor I_71655 (I1220681,I1270366,I1270375);
and I_71656 (I1220485,I1220681,I1220548);
not I_71657 (I1220712,I1270363);
nand I_71658 (I1220729,I1220712,I1270360);
nor I_71659 (I1220746,I1270363,I1270360);
not I_71660 (I1220763,I1220746);
nand I_71661 (I1220488,I1220630,I1220763);
DFFARX1 I_71662 (I1220746,I2507,I1220514,I1220503,);
nor I_71663 (I1220808,I1270363,I1270366);
nor I_71664 (I1220825,I1220808,I1270372);
and I_71665 (I1220842,I1220825,I1220729);
DFFARX1 I_71666 (I1220842,I2507,I1220514,I1220500,);
nor I_71667 (I1220497,I1220808,I1220664);
or I_71668 (I1220494,I1220746,I1220808);
nor I_71669 (I1220901,I1270363,I1270384);
DFFARX1 I_71670 (I1220901,I2507,I1220514,I1220927,);
not I_71671 (I1220935,I1220927);
nand I_71672 (I1220952,I1220935,I1220613);
nor I_71673 (I1220969,I1220952,I1270372);
DFFARX1 I_71674 (I1220969,I2507,I1220514,I1220482,);
nor I_71675 (I1221000,I1220935,I1220664);
nor I_71676 (I1220491,I1220808,I1221000);
not I_71677 (I1221058,I2514);
DFFARX1 I_71678 (I1094230,I2507,I1221058,I1221084,);
nand I_71679 (I1221092,I1221084,I1094209);
DFFARX1 I_71680 (I1094206,I2507,I1221058,I1221118,);
DFFARX1 I_71681 (I1221118,I2507,I1221058,I1221135,);
not I_71682 (I1221050,I1221135);
not I_71683 (I1221157,I1094218);
nor I_71684 (I1221174,I1094218,I1094227);
not I_71685 (I1221191,I1094215);
nand I_71686 (I1221208,I1221157,I1221191);
nor I_71687 (I1221225,I1094215,I1094218);
and I_71688 (I1221029,I1221225,I1221092);
not I_71689 (I1221256,I1094224);
nand I_71690 (I1221273,I1221256,I1094221);
nor I_71691 (I1221290,I1094224,I1094206);
not I_71692 (I1221307,I1221290);
nand I_71693 (I1221032,I1221174,I1221307);
DFFARX1 I_71694 (I1221290,I2507,I1221058,I1221047,);
nor I_71695 (I1221352,I1094209,I1094215);
nor I_71696 (I1221369,I1221352,I1094227);
and I_71697 (I1221386,I1221369,I1221273);
DFFARX1 I_71698 (I1221386,I2507,I1221058,I1221044,);
nor I_71699 (I1221041,I1221352,I1221208);
or I_71700 (I1221038,I1221290,I1221352);
nor I_71701 (I1221445,I1094209,I1094212);
DFFARX1 I_71702 (I1221445,I2507,I1221058,I1221471,);
not I_71703 (I1221479,I1221471);
nand I_71704 (I1221496,I1221479,I1221157);
nor I_71705 (I1221513,I1221496,I1094227);
DFFARX1 I_71706 (I1221513,I2507,I1221058,I1221026,);
nor I_71707 (I1221544,I1221479,I1221208);
nor I_71708 (I1221035,I1221352,I1221544);
not I_71709 (I1221602,I2514);
DFFARX1 I_71710 (I1046063,I2507,I1221602,I1221628,);
nand I_71711 (I1221636,I1221628,I1046051);
DFFARX1 I_71712 (I1046045,I2507,I1221602,I1221662,);
DFFARX1 I_71713 (I1221662,I2507,I1221602,I1221679,);
not I_71714 (I1221594,I1221679);
not I_71715 (I1221701,I1046045);
nor I_71716 (I1221718,I1046045,I1046057);
not I_71717 (I1221735,I1046054);
nand I_71718 (I1221752,I1221701,I1221735);
nor I_71719 (I1221769,I1046054,I1046045);
and I_71720 (I1221573,I1221769,I1221636);
not I_71721 (I1221800,I1046048);
nand I_71722 (I1221817,I1221800,I1046060);
nor I_71723 (I1221834,I1046048,I1046066);
not I_71724 (I1221851,I1221834);
nand I_71725 (I1221576,I1221718,I1221851);
DFFARX1 I_71726 (I1221834,I2507,I1221602,I1221591,);
nor I_71727 (I1221896,I1046051,I1046054);
nor I_71728 (I1221913,I1221896,I1046057);
and I_71729 (I1221930,I1221913,I1221817);
DFFARX1 I_71730 (I1221930,I2507,I1221602,I1221588,);
nor I_71731 (I1221585,I1221896,I1221752);
or I_71732 (I1221582,I1221834,I1221896);
nor I_71733 (I1221989,I1046051,I1046048);
DFFARX1 I_71734 (I1221989,I2507,I1221602,I1222015,);
not I_71735 (I1222023,I1222015);
nand I_71736 (I1222040,I1222023,I1221701);
nor I_71737 (I1222057,I1222040,I1046057);
DFFARX1 I_71738 (I1222057,I2507,I1221602,I1221570,);
nor I_71739 (I1222088,I1222023,I1221752);
nor I_71740 (I1221579,I1221896,I1222088);
not I_71741 (I1222146,I2514);
DFFARX1 I_71742 (I340846,I2507,I1222146,I1222172,);
nand I_71743 (I1222180,I1222172,I340849);
DFFARX1 I_71744 (I340843,I2507,I1222146,I1222206,);
DFFARX1 I_71745 (I1222206,I2507,I1222146,I1222223,);
not I_71746 (I1222138,I1222223);
not I_71747 (I1222245,I340852);
nor I_71748 (I1222262,I340852,I340837);
not I_71749 (I1222279,I340861);
nand I_71750 (I1222296,I1222245,I1222279);
nor I_71751 (I1222313,I340861,I340852);
and I_71752 (I1222117,I1222313,I1222180);
not I_71753 (I1222344,I340840);
nand I_71754 (I1222361,I1222344,I340858);
nor I_71755 (I1222378,I340840,I340834);
not I_71756 (I1222395,I1222378);
nand I_71757 (I1222120,I1222262,I1222395);
DFFARX1 I_71758 (I1222378,I2507,I1222146,I1222135,);
nor I_71759 (I1222440,I340855,I340861);
nor I_71760 (I1222457,I1222440,I340837);
and I_71761 (I1222474,I1222457,I1222361);
DFFARX1 I_71762 (I1222474,I2507,I1222146,I1222132,);
nor I_71763 (I1222129,I1222440,I1222296);
or I_71764 (I1222126,I1222378,I1222440);
nor I_71765 (I1222533,I340855,I340834);
DFFARX1 I_71766 (I1222533,I2507,I1222146,I1222559,);
not I_71767 (I1222567,I1222559);
nand I_71768 (I1222584,I1222567,I1222245);
nor I_71769 (I1222601,I1222584,I340837);
DFFARX1 I_71770 (I1222601,I2507,I1222146,I1222114,);
nor I_71771 (I1222632,I1222567,I1222296);
nor I_71772 (I1222123,I1222440,I1222632);
not I_71773 (I1222690,I2514);
DFFARX1 I_71774 (I723201,I2507,I1222690,I1222716,);
nand I_71775 (I1222724,I1222716,I723216);
DFFARX1 I_71776 (I723210,I2507,I1222690,I1222750,);
DFFARX1 I_71777 (I1222750,I2507,I1222690,I1222767,);
not I_71778 (I1222682,I1222767);
not I_71779 (I1222789,I723213);
nor I_71780 (I1222806,I723213,I723219);
not I_71781 (I1222823,I723201);
nand I_71782 (I1222840,I1222789,I1222823);
nor I_71783 (I1222857,I723201,I723213);
and I_71784 (I1222661,I1222857,I1222724);
not I_71785 (I1222888,I723198);
nand I_71786 (I1222905,I1222888,I723204);
nor I_71787 (I1222922,I723198,I723198);
not I_71788 (I1222939,I1222922);
nand I_71789 (I1222664,I1222806,I1222939);
DFFARX1 I_71790 (I1222922,I2507,I1222690,I1222679,);
nor I_71791 (I1222984,I723207,I723201);
nor I_71792 (I1223001,I1222984,I723219);
and I_71793 (I1223018,I1223001,I1222905);
DFFARX1 I_71794 (I1223018,I2507,I1222690,I1222676,);
nor I_71795 (I1222673,I1222984,I1222840);
or I_71796 (I1222670,I1222922,I1222984);
nor I_71797 (I1223077,I723207,I723222);
DFFARX1 I_71798 (I1223077,I2507,I1222690,I1223103,);
not I_71799 (I1223111,I1223103);
nand I_71800 (I1223128,I1223111,I1222789);
nor I_71801 (I1223145,I1223128,I723219);
DFFARX1 I_71802 (I1223145,I2507,I1222690,I1222658,);
nor I_71803 (I1223176,I1223111,I1222840);
nor I_71804 (I1222667,I1222984,I1223176);
not I_71805 (I1223234,I2514);
DFFARX1 I_71806 (I374047,I2507,I1223234,I1223260,);
nand I_71807 (I1223268,I1223260,I374050);
DFFARX1 I_71808 (I374044,I2507,I1223234,I1223294,);
DFFARX1 I_71809 (I1223294,I2507,I1223234,I1223311,);
not I_71810 (I1223226,I1223311);
not I_71811 (I1223333,I374053);
nor I_71812 (I1223350,I374053,I374038);
not I_71813 (I1223367,I374062);
nand I_71814 (I1223384,I1223333,I1223367);
nor I_71815 (I1223401,I374062,I374053);
and I_71816 (I1223205,I1223401,I1223268);
not I_71817 (I1223432,I374041);
nand I_71818 (I1223449,I1223432,I374059);
nor I_71819 (I1223466,I374041,I374035);
not I_71820 (I1223483,I1223466);
nand I_71821 (I1223208,I1223350,I1223483);
DFFARX1 I_71822 (I1223466,I2507,I1223234,I1223223,);
nor I_71823 (I1223528,I374056,I374062);
nor I_71824 (I1223545,I1223528,I374038);
and I_71825 (I1223562,I1223545,I1223449);
DFFARX1 I_71826 (I1223562,I2507,I1223234,I1223220,);
nor I_71827 (I1223217,I1223528,I1223384);
or I_71828 (I1223214,I1223466,I1223528);
nor I_71829 (I1223621,I374056,I374035);
DFFARX1 I_71830 (I1223621,I2507,I1223234,I1223647,);
not I_71831 (I1223655,I1223647);
nand I_71832 (I1223672,I1223655,I1223333);
nor I_71833 (I1223689,I1223672,I374038);
DFFARX1 I_71834 (I1223689,I2507,I1223234,I1223202,);
nor I_71835 (I1223720,I1223655,I1223384);
nor I_71836 (I1223211,I1223528,I1223720);
not I_71837 (I1223778,I2514);
DFFARX1 I_71838 (I645171,I2507,I1223778,I1223804,);
nand I_71839 (I1223812,I1223804,I645186);
DFFARX1 I_71840 (I645180,I2507,I1223778,I1223838,);
DFFARX1 I_71841 (I1223838,I2507,I1223778,I1223855,);
not I_71842 (I1223770,I1223855);
not I_71843 (I1223877,I645183);
nor I_71844 (I1223894,I645183,I645189);
not I_71845 (I1223911,I645171);
nand I_71846 (I1223928,I1223877,I1223911);
nor I_71847 (I1223945,I645171,I645183);
and I_71848 (I1223749,I1223945,I1223812);
not I_71849 (I1223976,I645168);
nand I_71850 (I1223993,I1223976,I645174);
nor I_71851 (I1224010,I645168,I645168);
not I_71852 (I1224027,I1224010);
nand I_71853 (I1223752,I1223894,I1224027);
DFFARX1 I_71854 (I1224010,I2507,I1223778,I1223767,);
nor I_71855 (I1224072,I645177,I645171);
nor I_71856 (I1224089,I1224072,I645189);
and I_71857 (I1224106,I1224089,I1223993);
DFFARX1 I_71858 (I1224106,I2507,I1223778,I1223764,);
nor I_71859 (I1223761,I1224072,I1223928);
or I_71860 (I1223758,I1224010,I1224072);
nor I_71861 (I1224165,I645177,I645192);
DFFARX1 I_71862 (I1224165,I2507,I1223778,I1224191,);
not I_71863 (I1224199,I1224191);
nand I_71864 (I1224216,I1224199,I1223877);
nor I_71865 (I1224233,I1224216,I645189);
DFFARX1 I_71866 (I1224233,I2507,I1223778,I1223746,);
nor I_71867 (I1224264,I1224199,I1223928);
nor I_71868 (I1223755,I1224072,I1224264);
not I_71869 (I1224322,I2514);
DFFARX1 I_71870 (I68056,I2507,I1224322,I1224348,);
nand I_71871 (I1224356,I1224348,I68038);
DFFARX1 I_71872 (I68035,I2507,I1224322,I1224382,);
DFFARX1 I_71873 (I1224382,I2507,I1224322,I1224399,);
not I_71874 (I1224314,I1224399);
not I_71875 (I1224421,I68053);
nor I_71876 (I1224438,I68053,I68047);
not I_71877 (I1224455,I68035);
nand I_71878 (I1224472,I1224421,I1224455);
nor I_71879 (I1224489,I68035,I68053);
and I_71880 (I1224293,I1224489,I1224356);
not I_71881 (I1224520,I68044);
nand I_71882 (I1224537,I1224520,I68050);
nor I_71883 (I1224554,I68044,I68038);
not I_71884 (I1224571,I1224554);
nand I_71885 (I1224296,I1224438,I1224571);
DFFARX1 I_71886 (I1224554,I2507,I1224322,I1224311,);
nor I_71887 (I1224616,I68041,I68035);
nor I_71888 (I1224633,I1224616,I68047);
and I_71889 (I1224650,I1224633,I1224537);
DFFARX1 I_71890 (I1224650,I2507,I1224322,I1224308,);
nor I_71891 (I1224305,I1224616,I1224472);
or I_71892 (I1224302,I1224554,I1224616);
nor I_71893 (I1224709,I68041,I68059);
DFFARX1 I_71894 (I1224709,I2507,I1224322,I1224735,);
not I_71895 (I1224743,I1224735);
nand I_71896 (I1224760,I1224743,I1224421);
nor I_71897 (I1224777,I1224760,I68047);
DFFARX1 I_71898 (I1224777,I2507,I1224322,I1224290,);
nor I_71899 (I1224808,I1224743,I1224472);
nor I_71900 (I1224299,I1224616,I1224808);
not I_71901 (I1224866,I2514);
DFFARX1 I_71902 (I216284,I2507,I1224866,I1224892,);
nand I_71903 (I1224900,I1224892,I216299);
DFFARX1 I_71904 (I216296,I2507,I1224866,I1224926,);
DFFARX1 I_71905 (I1224926,I2507,I1224866,I1224943,);
not I_71906 (I1224858,I1224943);
not I_71907 (I1224965,I216275);
nor I_71908 (I1224982,I216275,I216281);
not I_71909 (I1224999,I216287);
nand I_71910 (I1225016,I1224965,I1224999);
nor I_71911 (I1225033,I216287,I216275);
and I_71912 (I1224837,I1225033,I1224900);
not I_71913 (I1225064,I216293);
nand I_71914 (I1225081,I1225064,I216275);
nor I_71915 (I1225098,I216293,I216278);
not I_71916 (I1225115,I1225098);
nand I_71917 (I1224840,I1224982,I1225115);
DFFARX1 I_71918 (I1225098,I2507,I1224866,I1224855,);
nor I_71919 (I1225160,I216278,I216287);
nor I_71920 (I1225177,I1225160,I216281);
and I_71921 (I1225194,I1225177,I1225081);
DFFARX1 I_71922 (I1225194,I2507,I1224866,I1224852,);
nor I_71923 (I1224849,I1225160,I1225016);
or I_71924 (I1224846,I1225098,I1225160);
nor I_71925 (I1225253,I216278,I216290);
DFFARX1 I_71926 (I1225253,I2507,I1224866,I1225279,);
not I_71927 (I1225287,I1225279);
nand I_71928 (I1225304,I1225287,I1224965);
nor I_71929 (I1225321,I1225304,I216281);
DFFARX1 I_71930 (I1225321,I2507,I1224866,I1224834,);
nor I_71931 (I1225352,I1225287,I1225016);
nor I_71932 (I1224843,I1225160,I1225352);
not I_71933 (I1225410,I2514);
DFFARX1 I_71934 (I820699,I2507,I1225410,I1225436,);
nand I_71935 (I1225444,I1225436,I820693);
DFFARX1 I_71936 (I820696,I2507,I1225410,I1225470,);
DFFARX1 I_71937 (I1225470,I2507,I1225410,I1225487,);
not I_71938 (I1225402,I1225487);
not I_71939 (I1225509,I820702);
nor I_71940 (I1225526,I820702,I820696);
not I_71941 (I1225543,I820705);
nand I_71942 (I1225560,I1225509,I1225543);
nor I_71943 (I1225577,I820705,I820702);
and I_71944 (I1225381,I1225577,I1225444);
not I_71945 (I1225608,I820714);
nand I_71946 (I1225625,I1225608,I820708);
nor I_71947 (I1225642,I820714,I820711);
not I_71948 (I1225659,I1225642);
nand I_71949 (I1225384,I1225526,I1225659);
DFFARX1 I_71950 (I1225642,I2507,I1225410,I1225399,);
nor I_71951 (I1225704,I820693,I820705);
nor I_71952 (I1225721,I1225704,I820696);
and I_71953 (I1225738,I1225721,I1225625);
DFFARX1 I_71954 (I1225738,I2507,I1225410,I1225396,);
nor I_71955 (I1225393,I1225704,I1225560);
or I_71956 (I1225390,I1225642,I1225704);
nor I_71957 (I1225797,I820693,I820699);
DFFARX1 I_71958 (I1225797,I2507,I1225410,I1225823,);
not I_71959 (I1225831,I1225823);
nand I_71960 (I1225848,I1225831,I1225509);
nor I_71961 (I1225865,I1225848,I820696);
DFFARX1 I_71962 (I1225865,I2507,I1225410,I1225378,);
nor I_71963 (I1225896,I1225831,I1225560);
nor I_71964 (I1225387,I1225704,I1225896);
not I_71965 (I1225954,I2514);
DFFARX1 I_71966 (I698925,I2507,I1225954,I1225980,);
nand I_71967 (I1225988,I1225980,I698940);
DFFARX1 I_71968 (I698934,I2507,I1225954,I1226014,);
DFFARX1 I_71969 (I1226014,I2507,I1225954,I1226031,);
not I_71970 (I1225946,I1226031);
not I_71971 (I1226053,I698937);
nor I_71972 (I1226070,I698937,I698943);
not I_71973 (I1226087,I698925);
nand I_71974 (I1226104,I1226053,I1226087);
nor I_71975 (I1226121,I698925,I698937);
and I_71976 (I1225925,I1226121,I1225988);
not I_71977 (I1226152,I698922);
nand I_71978 (I1226169,I1226152,I698928);
nor I_71979 (I1226186,I698922,I698922);
not I_71980 (I1226203,I1226186);
nand I_71981 (I1225928,I1226070,I1226203);
DFFARX1 I_71982 (I1226186,I2507,I1225954,I1225943,);
nor I_71983 (I1226248,I698931,I698925);
nor I_71984 (I1226265,I1226248,I698943);
and I_71985 (I1226282,I1226265,I1226169);
DFFARX1 I_71986 (I1226282,I2507,I1225954,I1225940,);
nor I_71987 (I1225937,I1226248,I1226104);
or I_71988 (I1225934,I1226186,I1226248);
nor I_71989 (I1226341,I698931,I698946);
DFFARX1 I_71990 (I1226341,I2507,I1225954,I1226367,);
not I_71991 (I1226375,I1226367);
nand I_71992 (I1226392,I1226375,I1226053);
nor I_71993 (I1226409,I1226392,I698943);
DFFARX1 I_71994 (I1226409,I2507,I1225954,I1225922,);
nor I_71995 (I1226440,I1226375,I1226104);
nor I_71996 (I1225931,I1226248,I1226440);
not I_71997 (I1226498,I2514);
DFFARX1 I_71998 (I1186132,I2507,I1226498,I1226524,);
nand I_71999 (I1226532,I1226524,I1186111);
DFFARX1 I_72000 (I1186108,I2507,I1226498,I1226558,);
DFFARX1 I_72001 (I1226558,I2507,I1226498,I1226575,);
not I_72002 (I1226490,I1226575);
not I_72003 (I1226597,I1186120);
nor I_72004 (I1226614,I1186120,I1186129);
not I_72005 (I1226631,I1186117);
nand I_72006 (I1226648,I1226597,I1226631);
nor I_72007 (I1226665,I1186117,I1186120);
and I_72008 (I1226469,I1226665,I1226532);
not I_72009 (I1226696,I1186126);
nand I_72010 (I1226713,I1226696,I1186123);
nor I_72011 (I1226730,I1186126,I1186108);
not I_72012 (I1226747,I1226730);
nand I_72013 (I1226472,I1226614,I1226747);
DFFARX1 I_72014 (I1226730,I2507,I1226498,I1226487,);
nor I_72015 (I1226792,I1186111,I1186117);
nor I_72016 (I1226809,I1226792,I1186129);
and I_72017 (I1226826,I1226809,I1226713);
DFFARX1 I_72018 (I1226826,I2507,I1226498,I1226484,);
nor I_72019 (I1226481,I1226792,I1226648);
or I_72020 (I1226478,I1226730,I1226792);
nor I_72021 (I1226885,I1186111,I1186114);
DFFARX1 I_72022 (I1226885,I2507,I1226498,I1226911,);
not I_72023 (I1226919,I1226911);
nand I_72024 (I1226936,I1226919,I1226597);
nor I_72025 (I1226953,I1226936,I1186129);
DFFARX1 I_72026 (I1226953,I2507,I1226498,I1226466,);
nor I_72027 (I1226984,I1226919,I1226648);
nor I_72028 (I1226475,I1226792,I1226984);
not I_72029 (I1227042,I2514);
DFFARX1 I_72030 (I555599,I2507,I1227042,I1227068,);
nand I_72031 (I1227076,I1227068,I555587);
DFFARX1 I_72032 (I555593,I2507,I1227042,I1227102,);
DFFARX1 I_72033 (I1227102,I2507,I1227042,I1227119,);
not I_72034 (I1227034,I1227119);
not I_72035 (I1227141,I555578);
nor I_72036 (I1227158,I555578,I555590);
not I_72037 (I1227175,I555581);
nand I_72038 (I1227192,I1227141,I1227175);
nor I_72039 (I1227209,I555581,I555578);
and I_72040 (I1227013,I1227209,I1227076);
not I_72041 (I1227240,I555596);
nand I_72042 (I1227257,I1227240,I555578);
nor I_72043 (I1227274,I555596,I555602);
not I_72044 (I1227291,I1227274);
nand I_72045 (I1227016,I1227158,I1227291);
DFFARX1 I_72046 (I1227274,I2507,I1227042,I1227031,);
nor I_72047 (I1227336,I555584,I555581);
nor I_72048 (I1227353,I1227336,I555590);
and I_72049 (I1227370,I1227353,I1227257);
DFFARX1 I_72050 (I1227370,I2507,I1227042,I1227028,);
nor I_72051 (I1227025,I1227336,I1227192);
or I_72052 (I1227022,I1227274,I1227336);
nor I_72053 (I1227429,I555584,I555581);
DFFARX1 I_72054 (I1227429,I2507,I1227042,I1227455,);
not I_72055 (I1227463,I1227455);
nand I_72056 (I1227480,I1227463,I1227141);
nor I_72057 (I1227497,I1227480,I555590);
DFFARX1 I_72058 (I1227497,I2507,I1227042,I1227010,);
nor I_72059 (I1227528,I1227463,I1227192);
nor I_72060 (I1227019,I1227336,I1227528);
not I_72061 (I1227586,I2514);
DFFARX1 I_72062 (I1140470,I2507,I1227586,I1227612,);
nand I_72063 (I1227620,I1227612,I1140449);
DFFARX1 I_72064 (I1140446,I2507,I1227586,I1227646,);
DFFARX1 I_72065 (I1227646,I2507,I1227586,I1227663,);
not I_72066 (I1227578,I1227663);
not I_72067 (I1227685,I1140458);
nor I_72068 (I1227702,I1140458,I1140467);
not I_72069 (I1227719,I1140455);
nand I_72070 (I1227736,I1227685,I1227719);
nor I_72071 (I1227753,I1140455,I1140458);
and I_72072 (I1227557,I1227753,I1227620);
not I_72073 (I1227784,I1140464);
nand I_72074 (I1227801,I1227784,I1140461);
nor I_72075 (I1227818,I1140464,I1140446);
not I_72076 (I1227835,I1227818);
nand I_72077 (I1227560,I1227702,I1227835);
DFFARX1 I_72078 (I1227818,I2507,I1227586,I1227575,);
nor I_72079 (I1227880,I1140449,I1140455);
nor I_72080 (I1227897,I1227880,I1140467);
and I_72081 (I1227914,I1227897,I1227801);
DFFARX1 I_72082 (I1227914,I2507,I1227586,I1227572,);
nor I_72083 (I1227569,I1227880,I1227736);
or I_72084 (I1227566,I1227818,I1227880);
nor I_72085 (I1227973,I1140449,I1140452);
DFFARX1 I_72086 (I1227973,I2507,I1227586,I1227999,);
not I_72087 (I1228007,I1227999);
nand I_72088 (I1228024,I1228007,I1227685);
nor I_72089 (I1228041,I1228024,I1140467);
DFFARX1 I_72090 (I1228041,I2507,I1227586,I1227554,);
nor I_72091 (I1228072,I1228007,I1227736);
nor I_72092 (I1227563,I1227880,I1228072);
not I_72093 (I1228130,I2514);
DFFARX1 I_72094 (I2108,I2507,I1228130,I1228156,);
nand I_72095 (I1228164,I1228156,I2068);
DFFARX1 I_72096 (I1428,I2507,I1228130,I1228190,);
DFFARX1 I_72097 (I1228190,I2507,I1228130,I1228207,);
not I_72098 (I1228122,I1228207);
not I_72099 (I1228229,I1828);
nor I_72100 (I1228246,I1828,I1548);
not I_72101 (I1228263,I2388);
nand I_72102 (I1228280,I1228229,I1228263);
nor I_72103 (I1228297,I2388,I1828);
and I_72104 (I1228101,I1228297,I1228164);
not I_72105 (I1228328,I1692);
nand I_72106 (I1228345,I1228328,I2100);
nor I_72107 (I1228362,I1692,I1516);
not I_72108 (I1228379,I1228362);
nand I_72109 (I1228104,I1228246,I1228379);
DFFARX1 I_72110 (I1228362,I2507,I1228130,I1228119,);
nor I_72111 (I1228424,I1484,I2388);
nor I_72112 (I1228441,I1228424,I1548);
and I_72113 (I1228458,I1228441,I1228345);
DFFARX1 I_72114 (I1228458,I2507,I1228130,I1228116,);
nor I_72115 (I1228113,I1228424,I1228280);
or I_72116 (I1228110,I1228362,I1228424);
nor I_72117 (I1228517,I1484,I1540);
DFFARX1 I_72118 (I1228517,I2507,I1228130,I1228543,);
not I_72119 (I1228551,I1228543);
nand I_72120 (I1228568,I1228551,I1228229);
nor I_72121 (I1228585,I1228568,I1548);
DFFARX1 I_72122 (I1228585,I2507,I1228130,I1228098,);
nor I_72123 (I1228616,I1228551,I1228280);
nor I_72124 (I1228107,I1228424,I1228616);
not I_72125 (I1228674,I2514);
DFFARX1 I_72126 (I588545,I2507,I1228674,I1228700,);
nand I_72127 (I1228708,I1228700,I588533);
DFFARX1 I_72128 (I588539,I2507,I1228674,I1228734,);
DFFARX1 I_72129 (I1228734,I2507,I1228674,I1228751,);
not I_72130 (I1228666,I1228751);
not I_72131 (I1228773,I588524);
nor I_72132 (I1228790,I588524,I588536);
not I_72133 (I1228807,I588527);
nand I_72134 (I1228824,I1228773,I1228807);
nor I_72135 (I1228841,I588527,I588524);
and I_72136 (I1228645,I1228841,I1228708);
not I_72137 (I1228872,I588542);
nand I_72138 (I1228889,I1228872,I588524);
nor I_72139 (I1228906,I588542,I588548);
not I_72140 (I1228923,I1228906);
nand I_72141 (I1228648,I1228790,I1228923);
DFFARX1 I_72142 (I1228906,I2507,I1228674,I1228663,);
nor I_72143 (I1228968,I588530,I588527);
nor I_72144 (I1228985,I1228968,I588536);
and I_72145 (I1229002,I1228985,I1228889);
DFFARX1 I_72146 (I1229002,I2507,I1228674,I1228660,);
nor I_72147 (I1228657,I1228968,I1228824);
or I_72148 (I1228654,I1228906,I1228968);
nor I_72149 (I1229061,I588530,I588527);
DFFARX1 I_72150 (I1229061,I2507,I1228674,I1229087,);
not I_72151 (I1229095,I1229087);
nand I_72152 (I1229112,I1229095,I1228773);
nor I_72153 (I1229129,I1229112,I588536);
DFFARX1 I_72154 (I1229129,I2507,I1228674,I1228642,);
nor I_72155 (I1229160,I1229095,I1228824);
nor I_72156 (I1228651,I1228968,I1229160);
not I_72157 (I1229218,I2514);
DFFARX1 I_72158 (I467559,I2507,I1229218,I1229244,);
nand I_72159 (I1229252,I1229244,I467556);
DFFARX1 I_72160 (I467535,I2507,I1229218,I1229278,);
DFFARX1 I_72161 (I1229278,I2507,I1229218,I1229295,);
not I_72162 (I1229210,I1229295);
not I_72163 (I1229317,I467550);
nor I_72164 (I1229334,I467550,I467553);
not I_72165 (I1229351,I467544);
nand I_72166 (I1229368,I1229317,I1229351);
nor I_72167 (I1229385,I467544,I467550);
and I_72168 (I1229189,I1229385,I1229252);
not I_72169 (I1229416,I467541);
nand I_72170 (I1229433,I1229416,I467562);
nor I_72171 (I1229450,I467541,I467538);
not I_72172 (I1229467,I1229450);
nand I_72173 (I1229192,I1229334,I1229467);
DFFARX1 I_72174 (I1229450,I2507,I1229218,I1229207,);
nor I_72175 (I1229512,I467547,I467544);
nor I_72176 (I1229529,I1229512,I467553);
and I_72177 (I1229546,I1229529,I1229433);
DFFARX1 I_72178 (I1229546,I2507,I1229218,I1229204,);
nor I_72179 (I1229201,I1229512,I1229368);
or I_72180 (I1229198,I1229450,I1229512);
nor I_72181 (I1229605,I467547,I467535);
DFFARX1 I_72182 (I1229605,I2507,I1229218,I1229631,);
not I_72183 (I1229639,I1229631);
nand I_72184 (I1229656,I1229639,I1229317);
nor I_72185 (I1229673,I1229656,I467553);
DFFARX1 I_72186 (I1229673,I2507,I1229218,I1229186,);
nor I_72187 (I1229704,I1229639,I1229368);
nor I_72188 (I1229195,I1229512,I1229704);
not I_72189 (I1229762,I2514);
DFFARX1 I_72190 (I11451,I2507,I1229762,I1229788,);
nand I_72191 (I1229796,I1229788,I11463);
DFFARX1 I_72192 (I11460,I2507,I1229762,I1229822,);
DFFARX1 I_72193 (I1229822,I2507,I1229762,I1229839,);
not I_72194 (I1229754,I1229839);
not I_72195 (I1229861,I11448);
nor I_72196 (I1229878,I11448,I11448);
not I_72197 (I1229895,I11442);
nand I_72198 (I1229912,I1229861,I1229895);
nor I_72199 (I1229929,I11442,I11448);
and I_72200 (I1229733,I1229929,I1229796);
not I_72201 (I1229960,I11445);
nand I_72202 (I1229977,I1229960,I11445);
nor I_72203 (I1229994,I11445,I11454);
not I_72204 (I1230011,I1229994);
nand I_72205 (I1229736,I1229878,I1230011);
DFFARX1 I_72206 (I1229994,I2507,I1229762,I1229751,);
nor I_72207 (I1230056,I11442,I11442);
nor I_72208 (I1230073,I1230056,I11448);
and I_72209 (I1230090,I1230073,I1229977);
DFFARX1 I_72210 (I1230090,I2507,I1229762,I1229748,);
nor I_72211 (I1229745,I1230056,I1229912);
or I_72212 (I1229742,I1229994,I1230056);
nor I_72213 (I1230149,I11442,I11457);
DFFARX1 I_72214 (I1230149,I2507,I1229762,I1230175,);
not I_72215 (I1230183,I1230175);
nand I_72216 (I1230200,I1230183,I1229861);
nor I_72217 (I1230217,I1230200,I11448);
DFFARX1 I_72218 (I1230217,I2507,I1229762,I1229730,);
nor I_72219 (I1230248,I1230183,I1229912);
nor I_72220 (I1229739,I1230056,I1230248);
not I_72221 (I1230306,I2514);
DFFARX1 I_72222 (I1180930,I2507,I1230306,I1230332,);
nand I_72223 (I1230340,I1230332,I1180909);
DFFARX1 I_72224 (I1180906,I2507,I1230306,I1230366,);
DFFARX1 I_72225 (I1230366,I2507,I1230306,I1230383,);
not I_72226 (I1230298,I1230383);
not I_72227 (I1230405,I1180918);
nor I_72228 (I1230422,I1180918,I1180927);
not I_72229 (I1230439,I1180915);
nand I_72230 (I1230456,I1230405,I1230439);
nor I_72231 (I1230473,I1180915,I1180918);
and I_72232 (I1230277,I1230473,I1230340);
not I_72233 (I1230504,I1180924);
nand I_72234 (I1230521,I1230504,I1180921);
nor I_72235 (I1230538,I1180924,I1180906);
not I_72236 (I1230555,I1230538);
nand I_72237 (I1230280,I1230422,I1230555);
DFFARX1 I_72238 (I1230538,I2507,I1230306,I1230295,);
nor I_72239 (I1230600,I1180909,I1180915);
nor I_72240 (I1230617,I1230600,I1180927);
and I_72241 (I1230634,I1230617,I1230521);
DFFARX1 I_72242 (I1230634,I2507,I1230306,I1230292,);
nor I_72243 (I1230289,I1230600,I1230456);
or I_72244 (I1230286,I1230538,I1230600);
nor I_72245 (I1230693,I1180909,I1180912);
DFFARX1 I_72246 (I1230693,I2507,I1230306,I1230719,);
not I_72247 (I1230727,I1230719);
nand I_72248 (I1230744,I1230727,I1230405);
nor I_72249 (I1230761,I1230744,I1180927);
DFFARX1 I_72250 (I1230761,I2507,I1230306,I1230274,);
nor I_72251 (I1230792,I1230727,I1230456);
nor I_72252 (I1230283,I1230600,I1230792);
not I_72253 (I1230850,I2514);
DFFARX1 I_72254 (I426215,I2507,I1230850,I1230876,);
nand I_72255 (I1230884,I1230876,I426212);
DFFARX1 I_72256 (I426191,I2507,I1230850,I1230910,);
DFFARX1 I_72257 (I1230910,I2507,I1230850,I1230927,);
not I_72258 (I1230842,I1230927);
not I_72259 (I1230949,I426206);
nor I_72260 (I1230966,I426206,I426209);
not I_72261 (I1230983,I426200);
nand I_72262 (I1231000,I1230949,I1230983);
nor I_72263 (I1231017,I426200,I426206);
and I_72264 (I1230821,I1231017,I1230884);
not I_72265 (I1231048,I426197);
nand I_72266 (I1231065,I1231048,I426218);
nor I_72267 (I1231082,I426197,I426194);
not I_72268 (I1231099,I1231082);
nand I_72269 (I1230824,I1230966,I1231099);
DFFARX1 I_72270 (I1231082,I2507,I1230850,I1230839,);
nor I_72271 (I1231144,I426203,I426200);
nor I_72272 (I1231161,I1231144,I426209);
and I_72273 (I1231178,I1231161,I1231065);
DFFARX1 I_72274 (I1231178,I2507,I1230850,I1230836,);
nor I_72275 (I1230833,I1231144,I1231000);
or I_72276 (I1230830,I1231082,I1231144);
nor I_72277 (I1231237,I426203,I426191);
DFFARX1 I_72278 (I1231237,I2507,I1230850,I1231263,);
not I_72279 (I1231271,I1231263);
nand I_72280 (I1231288,I1231271,I1230949);
nor I_72281 (I1231305,I1231288,I426209);
DFFARX1 I_72282 (I1231305,I2507,I1230850,I1230818,);
nor I_72283 (I1231336,I1231271,I1231000);
nor I_72284 (I1230827,I1231144,I1231336);
not I_72285 (I1231394,I2514);
DFFARX1 I_72286 (I199624,I2507,I1231394,I1231420,);
nand I_72287 (I1231428,I1231420,I199639);
DFFARX1 I_72288 (I199636,I2507,I1231394,I1231454,);
DFFARX1 I_72289 (I1231454,I2507,I1231394,I1231471,);
not I_72290 (I1231386,I1231471);
not I_72291 (I1231493,I199615);
nor I_72292 (I1231510,I199615,I199621);
not I_72293 (I1231527,I199627);
nand I_72294 (I1231544,I1231493,I1231527);
nor I_72295 (I1231561,I199627,I199615);
and I_72296 (I1231365,I1231561,I1231428);
not I_72297 (I1231592,I199633);
nand I_72298 (I1231609,I1231592,I199615);
nor I_72299 (I1231626,I199633,I199618);
not I_72300 (I1231643,I1231626);
nand I_72301 (I1231368,I1231510,I1231643);
DFFARX1 I_72302 (I1231626,I2507,I1231394,I1231383,);
nor I_72303 (I1231688,I199618,I199627);
nor I_72304 (I1231705,I1231688,I199621);
and I_72305 (I1231722,I1231705,I1231609);
DFFARX1 I_72306 (I1231722,I2507,I1231394,I1231380,);
nor I_72307 (I1231377,I1231688,I1231544);
or I_72308 (I1231374,I1231626,I1231688);
nor I_72309 (I1231781,I199618,I199630);
DFFARX1 I_72310 (I1231781,I2507,I1231394,I1231807,);
not I_72311 (I1231815,I1231807);
nand I_72312 (I1231832,I1231815,I1231493);
nor I_72313 (I1231849,I1231832,I199621);
DFFARX1 I_72314 (I1231849,I2507,I1231394,I1231362,);
nor I_72315 (I1231880,I1231815,I1231544);
nor I_72316 (I1231371,I1231688,I1231880);
not I_72317 (I1231938,I2514);
DFFARX1 I_72318 (I1196536,I2507,I1231938,I1231964,);
nand I_72319 (I1231972,I1231964,I1196515);
DFFARX1 I_72320 (I1196512,I2507,I1231938,I1231998,);
DFFARX1 I_72321 (I1231998,I2507,I1231938,I1232015,);
not I_72322 (I1231930,I1232015);
not I_72323 (I1232037,I1196524);
nor I_72324 (I1232054,I1196524,I1196533);
not I_72325 (I1232071,I1196521);
nand I_72326 (I1232088,I1232037,I1232071);
nor I_72327 (I1232105,I1196521,I1196524);
and I_72328 (I1231909,I1232105,I1231972);
not I_72329 (I1232136,I1196530);
nand I_72330 (I1232153,I1232136,I1196527);
nor I_72331 (I1232170,I1196530,I1196512);
not I_72332 (I1232187,I1232170);
nand I_72333 (I1231912,I1232054,I1232187);
DFFARX1 I_72334 (I1232170,I2507,I1231938,I1231927,);
nor I_72335 (I1232232,I1196515,I1196521);
nor I_72336 (I1232249,I1232232,I1196533);
and I_72337 (I1232266,I1232249,I1232153);
DFFARX1 I_72338 (I1232266,I2507,I1231938,I1231924,);
nor I_72339 (I1231921,I1232232,I1232088);
or I_72340 (I1231918,I1232170,I1232232);
nor I_72341 (I1232325,I1196515,I1196518);
DFFARX1 I_72342 (I1232325,I2507,I1231938,I1232351,);
not I_72343 (I1232359,I1232351);
nand I_72344 (I1232376,I1232359,I1232037);
nor I_72345 (I1232393,I1232376,I1196533);
DFFARX1 I_72346 (I1232393,I2507,I1231938,I1231906,);
nor I_72347 (I1232424,I1232359,I1232088);
nor I_72348 (I1231915,I1232232,I1232424);
not I_72349 (I1232482,I2514);
DFFARX1 I_72350 (I772909,I2507,I1232482,I1232508,);
nand I_72351 (I1232516,I1232508,I772924);
DFFARX1 I_72352 (I772918,I2507,I1232482,I1232542,);
DFFARX1 I_72353 (I1232542,I2507,I1232482,I1232559,);
not I_72354 (I1232474,I1232559);
not I_72355 (I1232581,I772921);
nor I_72356 (I1232598,I772921,I772927);
not I_72357 (I1232615,I772909);
nand I_72358 (I1232632,I1232581,I1232615);
nor I_72359 (I1232649,I772909,I772921);
and I_72360 (I1232453,I1232649,I1232516);
not I_72361 (I1232680,I772906);
nand I_72362 (I1232697,I1232680,I772912);
nor I_72363 (I1232714,I772906,I772906);
not I_72364 (I1232731,I1232714);
nand I_72365 (I1232456,I1232598,I1232731);
DFFARX1 I_72366 (I1232714,I2507,I1232482,I1232471,);
nor I_72367 (I1232776,I772915,I772909);
nor I_72368 (I1232793,I1232776,I772927);
and I_72369 (I1232810,I1232793,I1232697);
DFFARX1 I_72370 (I1232810,I2507,I1232482,I1232468,);
nor I_72371 (I1232465,I1232776,I1232632);
or I_72372 (I1232462,I1232714,I1232776);
nor I_72373 (I1232869,I772915,I772930);
DFFARX1 I_72374 (I1232869,I2507,I1232482,I1232895,);
not I_72375 (I1232903,I1232895);
nand I_72376 (I1232920,I1232903,I1232581);
nor I_72377 (I1232937,I1232920,I772927);
DFFARX1 I_72378 (I1232937,I2507,I1232482,I1232450,);
nor I_72379 (I1232968,I1232903,I1232632);
nor I_72380 (I1232459,I1232776,I1232968);
not I_72381 (I1233026,I2514);
DFFARX1 I_72382 (I869183,I2507,I1233026,I1233052,);
nand I_72383 (I1233060,I1233052,I869177);
DFFARX1 I_72384 (I869180,I2507,I1233026,I1233086,);
DFFARX1 I_72385 (I1233086,I2507,I1233026,I1233103,);
not I_72386 (I1233018,I1233103);
not I_72387 (I1233125,I869186);
nor I_72388 (I1233142,I869186,I869180);
not I_72389 (I1233159,I869189);
nand I_72390 (I1233176,I1233125,I1233159);
nor I_72391 (I1233193,I869189,I869186);
and I_72392 (I1232997,I1233193,I1233060);
not I_72393 (I1233224,I869198);
nand I_72394 (I1233241,I1233224,I869192);
nor I_72395 (I1233258,I869198,I869195);
not I_72396 (I1233275,I1233258);
nand I_72397 (I1233000,I1233142,I1233275);
DFFARX1 I_72398 (I1233258,I2507,I1233026,I1233015,);
nor I_72399 (I1233320,I869177,I869189);
nor I_72400 (I1233337,I1233320,I869180);
and I_72401 (I1233354,I1233337,I1233241);
DFFARX1 I_72402 (I1233354,I2507,I1233026,I1233012,);
nor I_72403 (I1233009,I1233320,I1233176);
or I_72404 (I1233006,I1233258,I1233320);
nor I_72405 (I1233413,I869177,I869183);
DFFARX1 I_72406 (I1233413,I2507,I1233026,I1233439,);
not I_72407 (I1233447,I1233439);
nand I_72408 (I1233464,I1233447,I1233125);
nor I_72409 (I1233481,I1233464,I869180);
DFFARX1 I_72410 (I1233481,I2507,I1233026,I1232994,);
nor I_72411 (I1233512,I1233447,I1233176);
nor I_72412 (I1233003,I1233320,I1233512);
not I_72413 (I1233570,I2514);
DFFARX1 I_72414 (I209144,I2507,I1233570,I1233596,);
nand I_72415 (I1233604,I1233596,I209159);
DFFARX1 I_72416 (I209156,I2507,I1233570,I1233630,);
DFFARX1 I_72417 (I1233630,I2507,I1233570,I1233647,);
not I_72418 (I1233562,I1233647);
not I_72419 (I1233669,I209135);
nor I_72420 (I1233686,I209135,I209141);
not I_72421 (I1233703,I209147);
nand I_72422 (I1233720,I1233669,I1233703);
nor I_72423 (I1233737,I209147,I209135);
and I_72424 (I1233541,I1233737,I1233604);
not I_72425 (I1233768,I209153);
nand I_72426 (I1233785,I1233768,I209135);
nor I_72427 (I1233802,I209153,I209138);
not I_72428 (I1233819,I1233802);
nand I_72429 (I1233544,I1233686,I1233819);
DFFARX1 I_72430 (I1233802,I2507,I1233570,I1233559,);
nor I_72431 (I1233864,I209138,I209147);
nor I_72432 (I1233881,I1233864,I209141);
and I_72433 (I1233898,I1233881,I1233785);
DFFARX1 I_72434 (I1233898,I2507,I1233570,I1233556,);
nor I_72435 (I1233553,I1233864,I1233720);
or I_72436 (I1233550,I1233802,I1233864);
nor I_72437 (I1233957,I209138,I209150);
DFFARX1 I_72438 (I1233957,I2507,I1233570,I1233983,);
not I_72439 (I1233991,I1233983);
nand I_72440 (I1234008,I1233991,I1233669);
nor I_72441 (I1234025,I1234008,I209141);
DFFARX1 I_72442 (I1234025,I2507,I1233570,I1233538,);
nor I_72443 (I1234056,I1233991,I1233720);
nor I_72444 (I1233547,I1233864,I1234056);
not I_72445 (I1234114,I2514);
DFFARX1 I_72446 (I598371,I2507,I1234114,I1234140,);
nand I_72447 (I1234148,I1234140,I598359);
DFFARX1 I_72448 (I598365,I2507,I1234114,I1234174,);
DFFARX1 I_72449 (I1234174,I2507,I1234114,I1234191,);
not I_72450 (I1234106,I1234191);
not I_72451 (I1234213,I598350);
nor I_72452 (I1234230,I598350,I598362);
not I_72453 (I1234247,I598353);
nand I_72454 (I1234264,I1234213,I1234247);
nor I_72455 (I1234281,I598353,I598350);
and I_72456 (I1234085,I1234281,I1234148);
not I_72457 (I1234312,I598368);
nand I_72458 (I1234329,I1234312,I598350);
nor I_72459 (I1234346,I598368,I598374);
not I_72460 (I1234363,I1234346);
nand I_72461 (I1234088,I1234230,I1234363);
DFFARX1 I_72462 (I1234346,I2507,I1234114,I1234103,);
nor I_72463 (I1234408,I598356,I598353);
nor I_72464 (I1234425,I1234408,I598362);
and I_72465 (I1234442,I1234425,I1234329);
DFFARX1 I_72466 (I1234442,I2507,I1234114,I1234100,);
nor I_72467 (I1234097,I1234408,I1234264);
or I_72468 (I1234094,I1234346,I1234408);
nor I_72469 (I1234501,I598356,I598353);
DFFARX1 I_72470 (I1234501,I2507,I1234114,I1234527,);
not I_72471 (I1234535,I1234527);
nand I_72472 (I1234552,I1234535,I1234213);
nor I_72473 (I1234569,I1234552,I598362);
DFFARX1 I_72474 (I1234569,I2507,I1234114,I1234082,);
nor I_72475 (I1234600,I1234535,I1234264);
nor I_72476 (I1234091,I1234408,I1234600);
not I_72477 (I1234658,I2514);
DFFARX1 I_72478 (I708173,I2507,I1234658,I1234684,);
nand I_72479 (I1234692,I1234684,I708188);
DFFARX1 I_72480 (I708182,I2507,I1234658,I1234718,);
DFFARX1 I_72481 (I1234718,I2507,I1234658,I1234735,);
not I_72482 (I1234650,I1234735);
not I_72483 (I1234757,I708185);
nor I_72484 (I1234774,I708185,I708191);
not I_72485 (I1234791,I708173);
nand I_72486 (I1234808,I1234757,I1234791);
nor I_72487 (I1234825,I708173,I708185);
and I_72488 (I1234629,I1234825,I1234692);
not I_72489 (I1234856,I708170);
nand I_72490 (I1234873,I1234856,I708176);
nor I_72491 (I1234890,I708170,I708170);
not I_72492 (I1234907,I1234890);
nand I_72493 (I1234632,I1234774,I1234907);
DFFARX1 I_72494 (I1234890,I2507,I1234658,I1234647,);
nor I_72495 (I1234952,I708179,I708173);
nor I_72496 (I1234969,I1234952,I708191);
and I_72497 (I1234986,I1234969,I1234873);
DFFARX1 I_72498 (I1234986,I2507,I1234658,I1234644,);
nor I_72499 (I1234641,I1234952,I1234808);
or I_72500 (I1234638,I1234890,I1234952);
nor I_72501 (I1235045,I708179,I708194);
DFFARX1 I_72502 (I1235045,I2507,I1234658,I1235071,);
not I_72503 (I1235079,I1235071);
nand I_72504 (I1235096,I1235079,I1234757);
nor I_72505 (I1235113,I1235096,I708191);
DFFARX1 I_72506 (I1235113,I2507,I1234658,I1234626,);
nor I_72507 (I1235144,I1235079,I1234808);
nor I_72508 (I1234635,I1234952,I1235144);
not I_72509 (I1235202,I2514);
DFFARX1 I_72510 (I1100588,I2507,I1235202,I1235228,);
nand I_72511 (I1235236,I1235228,I1100567);
DFFARX1 I_72512 (I1100564,I2507,I1235202,I1235262,);
DFFARX1 I_72513 (I1235262,I2507,I1235202,I1235279,);
not I_72514 (I1235194,I1235279);
not I_72515 (I1235301,I1100576);
nor I_72516 (I1235318,I1100576,I1100585);
not I_72517 (I1235335,I1100573);
nand I_72518 (I1235352,I1235301,I1235335);
nor I_72519 (I1235369,I1100573,I1100576);
and I_72520 (I1235173,I1235369,I1235236);
not I_72521 (I1235400,I1100582);
nand I_72522 (I1235417,I1235400,I1100579);
nor I_72523 (I1235434,I1100582,I1100564);
not I_72524 (I1235451,I1235434);
nand I_72525 (I1235176,I1235318,I1235451);
DFFARX1 I_72526 (I1235434,I2507,I1235202,I1235191,);
nor I_72527 (I1235496,I1100567,I1100573);
nor I_72528 (I1235513,I1235496,I1100585);
and I_72529 (I1235530,I1235513,I1235417);
DFFARX1 I_72530 (I1235530,I2507,I1235202,I1235188,);
nor I_72531 (I1235185,I1235496,I1235352);
or I_72532 (I1235182,I1235434,I1235496);
nor I_72533 (I1235589,I1100567,I1100570);
DFFARX1 I_72534 (I1235589,I2507,I1235202,I1235615,);
not I_72535 (I1235623,I1235615);
nand I_72536 (I1235640,I1235623,I1235301);
nor I_72537 (I1235657,I1235640,I1100585);
DFFARX1 I_72538 (I1235657,I2507,I1235202,I1235170,);
nor I_72539 (I1235688,I1235623,I1235352);
nor I_72540 (I1235179,I1235496,I1235688);
not I_72541 (I1235746,I2514);
DFFARX1 I_72542 (I468647,I2507,I1235746,I1235772,);
nand I_72543 (I1235780,I1235772,I468644);
DFFARX1 I_72544 (I468623,I2507,I1235746,I1235806,);
DFFARX1 I_72545 (I1235806,I2507,I1235746,I1235823,);
not I_72546 (I1235738,I1235823);
not I_72547 (I1235845,I468638);
nor I_72548 (I1235862,I468638,I468641);
not I_72549 (I1235879,I468632);
nand I_72550 (I1235896,I1235845,I1235879);
nor I_72551 (I1235913,I468632,I468638);
and I_72552 (I1235717,I1235913,I1235780);
not I_72553 (I1235944,I468629);
nand I_72554 (I1235961,I1235944,I468650);
nor I_72555 (I1235978,I468629,I468626);
not I_72556 (I1235995,I1235978);
nand I_72557 (I1235720,I1235862,I1235995);
DFFARX1 I_72558 (I1235978,I2507,I1235746,I1235735,);
nor I_72559 (I1236040,I468635,I468632);
nor I_72560 (I1236057,I1236040,I468641);
and I_72561 (I1236074,I1236057,I1235961);
DFFARX1 I_72562 (I1236074,I2507,I1235746,I1235732,);
nor I_72563 (I1235729,I1236040,I1235896);
or I_72564 (I1235726,I1235978,I1236040);
nor I_72565 (I1236133,I468635,I468623);
DFFARX1 I_72566 (I1236133,I2507,I1235746,I1236159,);
not I_72567 (I1236167,I1236159);
nand I_72568 (I1236184,I1236167,I1235845);
nor I_72569 (I1236201,I1236184,I468641);
DFFARX1 I_72570 (I1236201,I2507,I1235746,I1235714,);
nor I_72571 (I1236232,I1236167,I1235896);
nor I_72572 (I1235723,I1236040,I1236232);
not I_72573 (I1236290,I2514);
DFFARX1 I_72574 (I784336,I2507,I1236290,I1236316,);
nand I_72575 (I1236324,I1236316,I784330);
DFFARX1 I_72576 (I784333,I2507,I1236290,I1236350,);
DFFARX1 I_72577 (I1236350,I2507,I1236290,I1236367,);
not I_72578 (I1236282,I1236367);
not I_72579 (I1236389,I784339);
nor I_72580 (I1236406,I784339,I784333);
not I_72581 (I1236423,I784342);
nand I_72582 (I1236440,I1236389,I1236423);
nor I_72583 (I1236457,I784342,I784339);
and I_72584 (I1236261,I1236457,I1236324);
not I_72585 (I1236488,I784351);
nand I_72586 (I1236505,I1236488,I784345);
nor I_72587 (I1236522,I784351,I784348);
not I_72588 (I1236539,I1236522);
nand I_72589 (I1236264,I1236406,I1236539);
DFFARX1 I_72590 (I1236522,I2507,I1236290,I1236279,);
nor I_72591 (I1236584,I784330,I784342);
nor I_72592 (I1236601,I1236584,I784333);
and I_72593 (I1236618,I1236601,I1236505);
DFFARX1 I_72594 (I1236618,I2507,I1236290,I1236276,);
nor I_72595 (I1236273,I1236584,I1236440);
or I_72596 (I1236270,I1236522,I1236584);
nor I_72597 (I1236677,I784330,I784336);
DFFARX1 I_72598 (I1236677,I2507,I1236290,I1236703,);
not I_72599 (I1236711,I1236703);
nand I_72600 (I1236728,I1236711,I1236389);
nor I_72601 (I1236745,I1236728,I784333);
DFFARX1 I_72602 (I1236745,I2507,I1236290,I1236258,);
nor I_72603 (I1236776,I1236711,I1236440);
nor I_72604 (I1236267,I1236584,I1236776);
not I_72605 (I1236834,I2514);
DFFARX1 I_72606 (I66475,I2507,I1236834,I1236860,);
nand I_72607 (I1236868,I1236860,I66457);
DFFARX1 I_72608 (I66454,I2507,I1236834,I1236894,);
DFFARX1 I_72609 (I1236894,I2507,I1236834,I1236911,);
not I_72610 (I1236826,I1236911);
not I_72611 (I1236933,I66472);
nor I_72612 (I1236950,I66472,I66466);
not I_72613 (I1236967,I66454);
nand I_72614 (I1236984,I1236933,I1236967);
nor I_72615 (I1237001,I66454,I66472);
and I_72616 (I1236805,I1237001,I1236868);
not I_72617 (I1237032,I66463);
nand I_72618 (I1237049,I1237032,I66469);
nor I_72619 (I1237066,I66463,I66457);
not I_72620 (I1237083,I1237066);
nand I_72621 (I1236808,I1236950,I1237083);
DFFARX1 I_72622 (I1237066,I2507,I1236834,I1236823,);
nor I_72623 (I1237128,I66460,I66454);
nor I_72624 (I1237145,I1237128,I66466);
and I_72625 (I1237162,I1237145,I1237049);
DFFARX1 I_72626 (I1237162,I2507,I1236834,I1236820,);
nor I_72627 (I1236817,I1237128,I1236984);
or I_72628 (I1236814,I1237066,I1237128);
nor I_72629 (I1237221,I66460,I66478);
DFFARX1 I_72630 (I1237221,I2507,I1236834,I1237247,);
not I_72631 (I1237255,I1237247);
nand I_72632 (I1237272,I1237255,I1236933);
nor I_72633 (I1237289,I1237272,I66466);
DFFARX1 I_72634 (I1237289,I2507,I1236834,I1236802,);
nor I_72635 (I1237320,I1237255,I1236984);
nor I_72636 (I1236811,I1237128,I1237320);
not I_72637 (I1237378,I2514);
DFFARX1 I_72638 (I1124864,I2507,I1237378,I1237404,);
nand I_72639 (I1237412,I1237404,I1124843);
DFFARX1 I_72640 (I1124840,I2507,I1237378,I1237438,);
DFFARX1 I_72641 (I1237438,I2507,I1237378,I1237455,);
not I_72642 (I1237370,I1237455);
not I_72643 (I1237477,I1124852);
nor I_72644 (I1237494,I1124852,I1124861);
not I_72645 (I1237511,I1124849);
nand I_72646 (I1237528,I1237477,I1237511);
nor I_72647 (I1237545,I1124849,I1124852);
and I_72648 (I1237349,I1237545,I1237412);
not I_72649 (I1237576,I1124858);
nand I_72650 (I1237593,I1237576,I1124855);
nor I_72651 (I1237610,I1124858,I1124840);
not I_72652 (I1237627,I1237610);
nand I_72653 (I1237352,I1237494,I1237627);
DFFARX1 I_72654 (I1237610,I2507,I1237378,I1237367,);
nor I_72655 (I1237672,I1124843,I1124849);
nor I_72656 (I1237689,I1237672,I1124861);
and I_72657 (I1237706,I1237689,I1237593);
DFFARX1 I_72658 (I1237706,I2507,I1237378,I1237364,);
nor I_72659 (I1237361,I1237672,I1237528);
or I_72660 (I1237358,I1237610,I1237672);
nor I_72661 (I1237765,I1124843,I1124846);
DFFARX1 I_72662 (I1237765,I2507,I1237378,I1237791,);
not I_72663 (I1237799,I1237791);
nand I_72664 (I1237816,I1237799,I1237477);
nor I_72665 (I1237833,I1237816,I1124861);
DFFARX1 I_72666 (I1237833,I2507,I1237378,I1237346,);
nor I_72667 (I1237864,I1237799,I1237528);
nor I_72668 (I1237355,I1237672,I1237864);
not I_72669 (I1237922,I2514);
DFFARX1 I_72670 (I560223,I2507,I1237922,I1237948,);
nand I_72671 (I1237956,I1237948,I560211);
DFFARX1 I_72672 (I560217,I2507,I1237922,I1237982,);
DFFARX1 I_72673 (I1237982,I2507,I1237922,I1237999,);
not I_72674 (I1237914,I1237999);
not I_72675 (I1238021,I560202);
nor I_72676 (I1238038,I560202,I560214);
not I_72677 (I1238055,I560205);
nand I_72678 (I1238072,I1238021,I1238055);
nor I_72679 (I1238089,I560205,I560202);
and I_72680 (I1237893,I1238089,I1237956);
not I_72681 (I1238120,I560220);
nand I_72682 (I1238137,I1238120,I560202);
nor I_72683 (I1238154,I560220,I560226);
not I_72684 (I1238171,I1238154);
nand I_72685 (I1237896,I1238038,I1238171);
DFFARX1 I_72686 (I1238154,I2507,I1237922,I1237911,);
nor I_72687 (I1238216,I560208,I560205);
nor I_72688 (I1238233,I1238216,I560214);
and I_72689 (I1238250,I1238233,I1238137);
DFFARX1 I_72690 (I1238250,I2507,I1237922,I1237908,);
nor I_72691 (I1237905,I1238216,I1238072);
or I_72692 (I1237902,I1238154,I1238216);
nor I_72693 (I1238309,I560208,I560205);
DFFARX1 I_72694 (I1238309,I2507,I1237922,I1238335,);
not I_72695 (I1238343,I1238335);
nand I_72696 (I1238360,I1238343,I1238021);
nor I_72697 (I1238377,I1238360,I560214);
DFFARX1 I_72698 (I1238377,I2507,I1237922,I1237890,);
nor I_72699 (I1238408,I1238343,I1238072);
nor I_72700 (I1237899,I1238216,I1238408);
not I_72701 (I1238466,I2514);
DFFARX1 I_72702 (I595481,I2507,I1238466,I1238492,);
nand I_72703 (I1238500,I1238492,I595469);
DFFARX1 I_72704 (I595475,I2507,I1238466,I1238526,);
DFFARX1 I_72705 (I1238526,I2507,I1238466,I1238543,);
not I_72706 (I1238458,I1238543);
not I_72707 (I1238565,I595460);
nor I_72708 (I1238582,I595460,I595472);
not I_72709 (I1238599,I595463);
nand I_72710 (I1238616,I1238565,I1238599);
nor I_72711 (I1238633,I595463,I595460);
and I_72712 (I1238437,I1238633,I1238500);
not I_72713 (I1238664,I595478);
nand I_72714 (I1238681,I1238664,I595460);
nor I_72715 (I1238698,I595478,I595484);
not I_72716 (I1238715,I1238698);
nand I_72717 (I1238440,I1238582,I1238715);
DFFARX1 I_72718 (I1238698,I2507,I1238466,I1238455,);
nor I_72719 (I1238760,I595466,I595463);
nor I_72720 (I1238777,I1238760,I595472);
and I_72721 (I1238794,I1238777,I1238681);
DFFARX1 I_72722 (I1238794,I2507,I1238466,I1238452,);
nor I_72723 (I1238449,I1238760,I1238616);
or I_72724 (I1238446,I1238698,I1238760);
nor I_72725 (I1238853,I595466,I595463);
DFFARX1 I_72726 (I1238853,I2507,I1238466,I1238879,);
not I_72727 (I1238887,I1238879);
nand I_72728 (I1238904,I1238887,I1238565);
nor I_72729 (I1238921,I1238904,I595472);
DFFARX1 I_72730 (I1238921,I2507,I1238466,I1238434,);
nor I_72731 (I1238952,I1238887,I1238616);
nor I_72732 (I1238443,I1238760,I1238952);
not I_72733 (I1239010,I2514);
DFFARX1 I_72734 (I849684,I2507,I1239010,I1239036,);
nand I_72735 (I1239044,I1239036,I849678);
DFFARX1 I_72736 (I849681,I2507,I1239010,I1239070,);
DFFARX1 I_72737 (I1239070,I2507,I1239010,I1239087,);
not I_72738 (I1239002,I1239087);
not I_72739 (I1239109,I849687);
nor I_72740 (I1239126,I849687,I849681);
not I_72741 (I1239143,I849690);
nand I_72742 (I1239160,I1239109,I1239143);
nor I_72743 (I1239177,I849690,I849687);
and I_72744 (I1238981,I1239177,I1239044);
not I_72745 (I1239208,I849699);
nand I_72746 (I1239225,I1239208,I849693);
nor I_72747 (I1239242,I849699,I849696);
not I_72748 (I1239259,I1239242);
nand I_72749 (I1238984,I1239126,I1239259);
DFFARX1 I_72750 (I1239242,I2507,I1239010,I1238999,);
nor I_72751 (I1239304,I849678,I849690);
nor I_72752 (I1239321,I1239304,I849681);
and I_72753 (I1239338,I1239321,I1239225);
DFFARX1 I_72754 (I1239338,I2507,I1239010,I1238996,);
nor I_72755 (I1238993,I1239304,I1239160);
or I_72756 (I1238990,I1239242,I1239304);
nor I_72757 (I1239397,I849678,I849684);
DFFARX1 I_72758 (I1239397,I2507,I1239010,I1239423,);
not I_72759 (I1239431,I1239423);
nand I_72760 (I1239448,I1239431,I1239109);
nor I_72761 (I1239465,I1239448,I849681);
DFFARX1 I_72762 (I1239465,I2507,I1239010,I1238978,);
nor I_72763 (I1239496,I1239431,I1239160);
nor I_72764 (I1238987,I1239304,I1239496);
not I_72765 (I1239554,I2514);
DFFARX1 I_72766 (I67002,I2507,I1239554,I1239580,);
nand I_72767 (I1239588,I1239580,I66984);
DFFARX1 I_72768 (I66981,I2507,I1239554,I1239614,);
DFFARX1 I_72769 (I1239614,I2507,I1239554,I1239631,);
not I_72770 (I1239546,I1239631);
not I_72771 (I1239653,I66999);
nor I_72772 (I1239670,I66999,I66993);
not I_72773 (I1239687,I66981);
nand I_72774 (I1239704,I1239653,I1239687);
nor I_72775 (I1239721,I66981,I66999);
and I_72776 (I1239525,I1239721,I1239588);
not I_72777 (I1239752,I66990);
nand I_72778 (I1239769,I1239752,I66996);
nor I_72779 (I1239786,I66990,I66984);
not I_72780 (I1239803,I1239786);
nand I_72781 (I1239528,I1239670,I1239803);
DFFARX1 I_72782 (I1239786,I2507,I1239554,I1239543,);
nor I_72783 (I1239848,I66987,I66981);
nor I_72784 (I1239865,I1239848,I66993);
and I_72785 (I1239882,I1239865,I1239769);
DFFARX1 I_72786 (I1239882,I2507,I1239554,I1239540,);
nor I_72787 (I1239537,I1239848,I1239704);
or I_72788 (I1239534,I1239786,I1239848);
nor I_72789 (I1239941,I66987,I67005);
DFFARX1 I_72790 (I1239941,I2507,I1239554,I1239967,);
not I_72791 (I1239975,I1239967);
nand I_72792 (I1239992,I1239975,I1239653);
nor I_72793 (I1240009,I1239992,I66993);
DFFARX1 I_72794 (I1240009,I2507,I1239554,I1239522,);
nor I_72795 (I1240040,I1239975,I1239704);
nor I_72796 (I1239531,I1239848,I1240040);
not I_72797 (I1240098,I2514);
DFFARX1 I_72798 (I1089028,I2507,I1240098,I1240124,);
nand I_72799 (I1240132,I1240124,I1089007);
DFFARX1 I_72800 (I1089004,I2507,I1240098,I1240158,);
DFFARX1 I_72801 (I1240158,I2507,I1240098,I1240175,);
not I_72802 (I1240090,I1240175);
not I_72803 (I1240197,I1089016);
nor I_72804 (I1240214,I1089016,I1089025);
not I_72805 (I1240231,I1089013);
nand I_72806 (I1240248,I1240197,I1240231);
nor I_72807 (I1240265,I1089013,I1089016);
and I_72808 (I1240069,I1240265,I1240132);
not I_72809 (I1240296,I1089022);
nand I_72810 (I1240313,I1240296,I1089019);
nor I_72811 (I1240330,I1089022,I1089004);
not I_72812 (I1240347,I1240330);
nand I_72813 (I1240072,I1240214,I1240347);
DFFARX1 I_72814 (I1240330,I2507,I1240098,I1240087,);
nor I_72815 (I1240392,I1089007,I1089013);
nor I_72816 (I1240409,I1240392,I1089025);
and I_72817 (I1240426,I1240409,I1240313);
DFFARX1 I_72818 (I1240426,I2507,I1240098,I1240084,);
nor I_72819 (I1240081,I1240392,I1240248);
or I_72820 (I1240078,I1240330,I1240392);
nor I_72821 (I1240485,I1089007,I1089010);
DFFARX1 I_72822 (I1240485,I2507,I1240098,I1240511,);
not I_72823 (I1240519,I1240511);
nand I_72824 (I1240536,I1240519,I1240197);
nor I_72825 (I1240553,I1240536,I1089025);
DFFARX1 I_72826 (I1240553,I2507,I1240098,I1240066,);
nor I_72827 (I1240584,I1240519,I1240248);
nor I_72828 (I1240075,I1240392,I1240584);
not I_72829 (I1240642,I2514);
DFFARX1 I_72830 (I802781,I2507,I1240642,I1240668,);
nand I_72831 (I1240676,I1240668,I802775);
DFFARX1 I_72832 (I802778,I2507,I1240642,I1240702,);
DFFARX1 I_72833 (I1240702,I2507,I1240642,I1240719,);
not I_72834 (I1240634,I1240719);
not I_72835 (I1240741,I802784);
nor I_72836 (I1240758,I802784,I802778);
not I_72837 (I1240775,I802787);
nand I_72838 (I1240792,I1240741,I1240775);
nor I_72839 (I1240809,I802787,I802784);
and I_72840 (I1240613,I1240809,I1240676);
not I_72841 (I1240840,I802796);
nand I_72842 (I1240857,I1240840,I802790);
nor I_72843 (I1240874,I802796,I802793);
not I_72844 (I1240891,I1240874);
nand I_72845 (I1240616,I1240758,I1240891);
DFFARX1 I_72846 (I1240874,I2507,I1240642,I1240631,);
nor I_72847 (I1240936,I802775,I802787);
nor I_72848 (I1240953,I1240936,I802778);
and I_72849 (I1240970,I1240953,I1240857);
DFFARX1 I_72850 (I1240970,I2507,I1240642,I1240628,);
nor I_72851 (I1240625,I1240936,I1240792);
or I_72852 (I1240622,I1240874,I1240936);
nor I_72853 (I1241029,I802775,I802781);
DFFARX1 I_72854 (I1241029,I2507,I1240642,I1241055,);
not I_72855 (I1241063,I1241055);
nand I_72856 (I1241080,I1241063,I1240741);
nor I_72857 (I1241097,I1241080,I802778);
DFFARX1 I_72858 (I1241097,I2507,I1240642,I1240610,);
nor I_72859 (I1241128,I1241063,I1240792);
nor I_72860 (I1240619,I1240936,I1241128);
not I_72861 (I1241186,I2514);
DFFARX1 I_72862 (I312388,I2507,I1241186,I1241212,);
nand I_72863 (I1241220,I1241212,I312391);
DFFARX1 I_72864 (I312385,I2507,I1241186,I1241246,);
DFFARX1 I_72865 (I1241246,I2507,I1241186,I1241263,);
not I_72866 (I1241178,I1241263);
not I_72867 (I1241285,I312394);
nor I_72868 (I1241302,I312394,I312379);
not I_72869 (I1241319,I312403);
nand I_72870 (I1241336,I1241285,I1241319);
nor I_72871 (I1241353,I312403,I312394);
and I_72872 (I1241157,I1241353,I1241220);
not I_72873 (I1241384,I312382);
nand I_72874 (I1241401,I1241384,I312400);
nor I_72875 (I1241418,I312382,I312376);
not I_72876 (I1241435,I1241418);
nand I_72877 (I1241160,I1241302,I1241435);
DFFARX1 I_72878 (I1241418,I2507,I1241186,I1241175,);
nor I_72879 (I1241480,I312397,I312403);
nor I_72880 (I1241497,I1241480,I312379);
and I_72881 (I1241514,I1241497,I1241401);
DFFARX1 I_72882 (I1241514,I2507,I1241186,I1241172,);
nor I_72883 (I1241169,I1241480,I1241336);
or I_72884 (I1241166,I1241418,I1241480);
nor I_72885 (I1241573,I312397,I312376);
DFFARX1 I_72886 (I1241573,I2507,I1241186,I1241599,);
not I_72887 (I1241607,I1241599);
nand I_72888 (I1241624,I1241607,I1241285);
nor I_72889 (I1241641,I1241624,I312379);
DFFARX1 I_72890 (I1241641,I2507,I1241186,I1241154,);
nor I_72891 (I1241672,I1241607,I1241336);
nor I_72892 (I1241163,I1241480,I1241672);
not I_72893 (I1241730,I2514);
DFFARX1 I_72894 (I581031,I2507,I1241730,I1241756,);
nand I_72895 (I1241764,I1241756,I581019);
DFFARX1 I_72896 (I581025,I2507,I1241730,I1241790,);
DFFARX1 I_72897 (I1241790,I2507,I1241730,I1241807,);
not I_72898 (I1241722,I1241807);
not I_72899 (I1241829,I581010);
nor I_72900 (I1241846,I581010,I581022);
not I_72901 (I1241863,I581013);
nand I_72902 (I1241880,I1241829,I1241863);
nor I_72903 (I1241897,I581013,I581010);
and I_72904 (I1241701,I1241897,I1241764);
not I_72905 (I1241928,I581028);
nand I_72906 (I1241945,I1241928,I581010);
nor I_72907 (I1241962,I581028,I581034);
not I_72908 (I1241979,I1241962);
nand I_72909 (I1241704,I1241846,I1241979);
DFFARX1 I_72910 (I1241962,I2507,I1241730,I1241719,);
nor I_72911 (I1242024,I581016,I581013);
nor I_72912 (I1242041,I1242024,I581022);
and I_72913 (I1242058,I1242041,I1241945);
DFFARX1 I_72914 (I1242058,I2507,I1241730,I1241716,);
nor I_72915 (I1241713,I1242024,I1241880);
or I_72916 (I1241710,I1241962,I1242024);
nor I_72917 (I1242117,I581016,I581013);
DFFARX1 I_72918 (I1242117,I2507,I1241730,I1242143,);
not I_72919 (I1242151,I1242143);
nand I_72920 (I1242168,I1242151,I1241829);
nor I_72921 (I1242185,I1242168,I581022);
DFFARX1 I_72922 (I1242185,I2507,I1241730,I1241698,);
nor I_72923 (I1242216,I1242151,I1241880);
nor I_72924 (I1241707,I1242024,I1242216);
not I_72925 (I1242274,I2514);
DFFARX1 I_72926 (I343481,I2507,I1242274,I1242300,);
nand I_72927 (I1242308,I1242300,I343484);
DFFARX1 I_72928 (I343478,I2507,I1242274,I1242334,);
DFFARX1 I_72929 (I1242334,I2507,I1242274,I1242351,);
not I_72930 (I1242266,I1242351);
not I_72931 (I1242373,I343487);
nor I_72932 (I1242390,I343487,I343472);
not I_72933 (I1242407,I343496);
nand I_72934 (I1242424,I1242373,I1242407);
nor I_72935 (I1242441,I343496,I343487);
and I_72936 (I1242245,I1242441,I1242308);
not I_72937 (I1242472,I343475);
nand I_72938 (I1242489,I1242472,I343493);
nor I_72939 (I1242506,I343475,I343469);
not I_72940 (I1242523,I1242506);
nand I_72941 (I1242248,I1242390,I1242523);
DFFARX1 I_72942 (I1242506,I2507,I1242274,I1242263,);
nor I_72943 (I1242568,I343490,I343496);
nor I_72944 (I1242585,I1242568,I343472);
and I_72945 (I1242602,I1242585,I1242489);
DFFARX1 I_72946 (I1242602,I2507,I1242274,I1242260,);
nor I_72947 (I1242257,I1242568,I1242424);
or I_72948 (I1242254,I1242506,I1242568);
nor I_72949 (I1242661,I343490,I343469);
DFFARX1 I_72950 (I1242661,I2507,I1242274,I1242687,);
not I_72951 (I1242695,I1242687);
nand I_72952 (I1242712,I1242695,I1242373);
nor I_72953 (I1242729,I1242712,I343472);
DFFARX1 I_72954 (I1242729,I2507,I1242274,I1242242,);
nor I_72955 (I1242760,I1242695,I1242424);
nor I_72956 (I1242251,I1242568,I1242760);
not I_72957 (I1242818,I2514);
DFFARX1 I_72958 (I517294,I2507,I1242818,I1242844,);
nand I_72959 (I1242852,I1242844,I517318);
DFFARX1 I_72960 (I517297,I2507,I1242818,I1242878,);
DFFARX1 I_72961 (I1242878,I2507,I1242818,I1242895,);
not I_72962 (I1242810,I1242895);
not I_72963 (I1242917,I517300);
nor I_72964 (I1242934,I517300,I517315);
not I_72965 (I1242951,I517306);
nand I_72966 (I1242968,I1242917,I1242951);
nor I_72967 (I1242985,I517306,I517300);
and I_72968 (I1242789,I1242985,I1242852);
not I_72969 (I1243016,I517303);
nand I_72970 (I1243033,I1243016,I517297);
nor I_72971 (I1243050,I517303,I517312);
not I_72972 (I1243067,I1243050);
nand I_72973 (I1242792,I1242934,I1243067);
DFFARX1 I_72974 (I1243050,I2507,I1242818,I1242807,);
nor I_72975 (I1243112,I517309,I517306);
nor I_72976 (I1243129,I1243112,I517315);
and I_72977 (I1243146,I1243129,I1243033);
DFFARX1 I_72978 (I1243146,I2507,I1242818,I1242804,);
nor I_72979 (I1242801,I1243112,I1242968);
or I_72980 (I1242798,I1243050,I1243112);
nor I_72981 (I1243205,I517309,I517294);
DFFARX1 I_72982 (I1243205,I2507,I1242818,I1243231,);
not I_72983 (I1243239,I1243231);
nand I_72984 (I1243256,I1243239,I1242917);
nor I_72985 (I1243273,I1243256,I517315);
DFFARX1 I_72986 (I1243273,I2507,I1242818,I1242786,);
nor I_72987 (I1243304,I1243239,I1242968);
nor I_72988 (I1242795,I1243112,I1243304);
not I_72989 (I1243362,I2514);
DFFARX1 I_72990 (I50138,I2507,I1243362,I1243388,);
nand I_72991 (I1243396,I1243388,I50120);
DFFARX1 I_72992 (I50117,I2507,I1243362,I1243422,);
DFFARX1 I_72993 (I1243422,I2507,I1243362,I1243439,);
not I_72994 (I1243354,I1243439);
not I_72995 (I1243461,I50135);
nor I_72996 (I1243478,I50135,I50129);
not I_72997 (I1243495,I50117);
nand I_72998 (I1243512,I1243461,I1243495);
nor I_72999 (I1243529,I50117,I50135);
and I_73000 (I1243333,I1243529,I1243396);
not I_73001 (I1243560,I50126);
nand I_73002 (I1243577,I1243560,I50132);
nor I_73003 (I1243594,I50126,I50120);
not I_73004 (I1243611,I1243594);
nand I_73005 (I1243336,I1243478,I1243611);
DFFARX1 I_73006 (I1243594,I2507,I1243362,I1243351,);
nor I_73007 (I1243656,I50123,I50117);
nor I_73008 (I1243673,I1243656,I50129);
and I_73009 (I1243690,I1243673,I1243577);
DFFARX1 I_73010 (I1243690,I2507,I1243362,I1243348,);
nor I_73011 (I1243345,I1243656,I1243512);
or I_73012 (I1243342,I1243594,I1243656);
nor I_73013 (I1243749,I50123,I50141);
DFFARX1 I_73014 (I1243749,I2507,I1243362,I1243775,);
not I_73015 (I1243783,I1243775);
nand I_73016 (I1243800,I1243783,I1243461);
nor I_73017 (I1243817,I1243800,I50129);
DFFARX1 I_73018 (I1243817,I2507,I1243362,I1243330,);
nor I_73019 (I1243848,I1243783,I1243512);
nor I_73020 (I1243339,I1243656,I1243848);
not I_73021 (I1243906,I2514);
DFFARX1 I_73022 (I1202316,I2507,I1243906,I1243932,);
nand I_73023 (I1243940,I1243932,I1202295);
DFFARX1 I_73024 (I1202292,I2507,I1243906,I1243966,);
DFFARX1 I_73025 (I1243966,I2507,I1243906,I1243983,);
not I_73026 (I1243898,I1243983);
not I_73027 (I1244005,I1202304);
nor I_73028 (I1244022,I1202304,I1202313);
not I_73029 (I1244039,I1202301);
nand I_73030 (I1244056,I1244005,I1244039);
nor I_73031 (I1244073,I1202301,I1202304);
and I_73032 (I1243877,I1244073,I1243940);
not I_73033 (I1244104,I1202310);
nand I_73034 (I1244121,I1244104,I1202307);
nor I_73035 (I1244138,I1202310,I1202292);
not I_73036 (I1244155,I1244138);
nand I_73037 (I1243880,I1244022,I1244155);
DFFARX1 I_73038 (I1244138,I2507,I1243906,I1243895,);
nor I_73039 (I1244200,I1202295,I1202301);
nor I_73040 (I1244217,I1244200,I1202313);
and I_73041 (I1244234,I1244217,I1244121);
DFFARX1 I_73042 (I1244234,I2507,I1243906,I1243892,);
nor I_73043 (I1243889,I1244200,I1244056);
or I_73044 (I1243886,I1244138,I1244200);
nor I_73045 (I1244293,I1202295,I1202298);
DFFARX1 I_73046 (I1244293,I2507,I1243906,I1244319,);
not I_73047 (I1244327,I1244319);
nand I_73048 (I1244344,I1244327,I1244005);
nor I_73049 (I1244361,I1244344,I1202313);
DFFARX1 I_73050 (I1244361,I2507,I1243906,I1243874,);
nor I_73051 (I1244392,I1244327,I1244056);
nor I_73052 (I1243883,I1244200,I1244392);
not I_73053 (I1244450,I2514);
DFFARX1 I_73054 (I942481,I2507,I1244450,I1244476,);
nand I_73055 (I1244484,I1244476,I942481);
DFFARX1 I_73056 (I942493,I2507,I1244450,I1244510,);
DFFARX1 I_73057 (I1244510,I2507,I1244450,I1244527,);
not I_73058 (I1244442,I1244527);
not I_73059 (I1244549,I942487);
nor I_73060 (I1244566,I942487,I942508);
not I_73061 (I1244583,I942496);
nand I_73062 (I1244600,I1244549,I1244583);
nor I_73063 (I1244617,I942496,I942487);
and I_73064 (I1244421,I1244617,I1244484);
not I_73065 (I1244648,I942490);
nand I_73066 (I1244665,I1244648,I942505);
nor I_73067 (I1244682,I942490,I942499);
not I_73068 (I1244699,I1244682);
nand I_73069 (I1244424,I1244566,I1244699);
DFFARX1 I_73070 (I1244682,I2507,I1244450,I1244439,);
nor I_73071 (I1244744,I942502,I942496);
nor I_73072 (I1244761,I1244744,I942508);
and I_73073 (I1244778,I1244761,I1244665);
DFFARX1 I_73074 (I1244778,I2507,I1244450,I1244436,);
nor I_73075 (I1244433,I1244744,I1244600);
or I_73076 (I1244430,I1244682,I1244744);
nor I_73077 (I1244837,I942502,I942484);
DFFARX1 I_73078 (I1244837,I2507,I1244450,I1244863,);
not I_73079 (I1244871,I1244863);
nand I_73080 (I1244888,I1244871,I1244549);
nor I_73081 (I1244905,I1244888,I942508);
DFFARX1 I_73082 (I1244905,I2507,I1244450,I1244418,);
nor I_73083 (I1244936,I1244871,I1244600);
nor I_73084 (I1244427,I1244744,I1244936);
not I_73085 (I1244994,I2514);
DFFARX1 I_73086 (I357183,I2507,I1244994,I1245020,);
nand I_73087 (I1245028,I1245020,I357186);
DFFARX1 I_73088 (I357180,I2507,I1244994,I1245054,);
DFFARX1 I_73089 (I1245054,I2507,I1244994,I1245071,);
not I_73090 (I1244986,I1245071);
not I_73091 (I1245093,I357189);
nor I_73092 (I1245110,I357189,I357174);
not I_73093 (I1245127,I357198);
nand I_73094 (I1245144,I1245093,I1245127);
nor I_73095 (I1245161,I357198,I357189);
and I_73096 (I1244965,I1245161,I1245028);
not I_73097 (I1245192,I357177);
nand I_73098 (I1245209,I1245192,I357195);
nor I_73099 (I1245226,I357177,I357171);
not I_73100 (I1245243,I1245226);
nand I_73101 (I1244968,I1245110,I1245243);
DFFARX1 I_73102 (I1245226,I2507,I1244994,I1244983,);
nor I_73103 (I1245288,I357192,I357198);
nor I_73104 (I1245305,I1245288,I357174);
and I_73105 (I1245322,I1245305,I1245209);
DFFARX1 I_73106 (I1245322,I2507,I1244994,I1244980,);
nor I_73107 (I1244977,I1245288,I1245144);
or I_73108 (I1244974,I1245226,I1245288);
nor I_73109 (I1245381,I357192,I357171);
DFFARX1 I_73110 (I1245381,I2507,I1244994,I1245407,);
not I_73111 (I1245415,I1245407);
nand I_73112 (I1245432,I1245415,I1245093);
nor I_73113 (I1245449,I1245432,I357174);
DFFARX1 I_73114 (I1245449,I2507,I1244994,I1244962,);
nor I_73115 (I1245480,I1245415,I1245144);
nor I_73116 (I1244971,I1245288,I1245480);
not I_73117 (I1245538,I2514);
DFFARX1 I_73118 (I187129,I2507,I1245538,I1245564,);
nand I_73119 (I1245572,I1245564,I187144);
DFFARX1 I_73120 (I187141,I2507,I1245538,I1245598,);
DFFARX1 I_73121 (I1245598,I2507,I1245538,I1245615,);
not I_73122 (I1245530,I1245615);
not I_73123 (I1245637,I187120);
nor I_73124 (I1245654,I187120,I187126);
not I_73125 (I1245671,I187132);
nand I_73126 (I1245688,I1245637,I1245671);
nor I_73127 (I1245705,I187132,I187120);
and I_73128 (I1245509,I1245705,I1245572);
not I_73129 (I1245736,I187138);
nand I_73130 (I1245753,I1245736,I187120);
nor I_73131 (I1245770,I187138,I187123);
not I_73132 (I1245787,I1245770);
nand I_73133 (I1245512,I1245654,I1245787);
DFFARX1 I_73134 (I1245770,I2507,I1245538,I1245527,);
nor I_73135 (I1245832,I187123,I187132);
nor I_73136 (I1245849,I1245832,I187126);
and I_73137 (I1245866,I1245849,I1245753);
DFFARX1 I_73138 (I1245866,I2507,I1245538,I1245524,);
nor I_73139 (I1245521,I1245832,I1245688);
or I_73140 (I1245518,I1245770,I1245832);
nor I_73141 (I1245925,I187123,I187135);
DFFARX1 I_73142 (I1245925,I2507,I1245538,I1245951,);
not I_73143 (I1245959,I1245951);
nand I_73144 (I1245976,I1245959,I1245637);
nor I_73145 (I1245993,I1245976,I187126);
DFFARX1 I_73146 (I1245993,I2507,I1245538,I1245506,);
nor I_73147 (I1246024,I1245959,I1245688);
nor I_73148 (I1245515,I1245832,I1246024);
not I_73149 (I1246082,I2514);
DFFARX1 I_73150 (I1194224,I2507,I1246082,I1246108,);
nand I_73151 (I1246116,I1246108,I1194203);
DFFARX1 I_73152 (I1194200,I2507,I1246082,I1246142,);
DFFARX1 I_73153 (I1246142,I2507,I1246082,I1246159,);
not I_73154 (I1246074,I1246159);
not I_73155 (I1246181,I1194212);
nor I_73156 (I1246198,I1194212,I1194221);
not I_73157 (I1246215,I1194209);
nand I_73158 (I1246232,I1246181,I1246215);
nor I_73159 (I1246249,I1194209,I1194212);
and I_73160 (I1246053,I1246249,I1246116);
not I_73161 (I1246280,I1194218);
nand I_73162 (I1246297,I1246280,I1194215);
nor I_73163 (I1246314,I1194218,I1194200);
not I_73164 (I1246331,I1246314);
nand I_73165 (I1246056,I1246198,I1246331);
DFFARX1 I_73166 (I1246314,I2507,I1246082,I1246071,);
nor I_73167 (I1246376,I1194203,I1194209);
nor I_73168 (I1246393,I1246376,I1194221);
and I_73169 (I1246410,I1246393,I1246297);
DFFARX1 I_73170 (I1246410,I2507,I1246082,I1246068,);
nor I_73171 (I1246065,I1246376,I1246232);
or I_73172 (I1246062,I1246314,I1246376);
nor I_73173 (I1246469,I1194203,I1194206);
DFFARX1 I_73174 (I1246469,I2507,I1246082,I1246495,);
not I_73175 (I1246503,I1246495);
nand I_73176 (I1246520,I1246503,I1246181);
nor I_73177 (I1246537,I1246520,I1194221);
DFFARX1 I_73178 (I1246537,I2507,I1246082,I1246050,);
nor I_73179 (I1246568,I1246503,I1246232);
nor I_73180 (I1246059,I1246376,I1246568);
not I_73181 (I1246626,I2514);
DFFARX1 I_73182 (I1054478,I2507,I1246626,I1246652,);
nand I_73183 (I1246660,I1246652,I1054466);
DFFARX1 I_73184 (I1054460,I2507,I1246626,I1246686,);
DFFARX1 I_73185 (I1246686,I2507,I1246626,I1246703,);
not I_73186 (I1246618,I1246703);
not I_73187 (I1246725,I1054460);
nor I_73188 (I1246742,I1054460,I1054472);
not I_73189 (I1246759,I1054469);
nand I_73190 (I1246776,I1246725,I1246759);
nor I_73191 (I1246793,I1054469,I1054460);
and I_73192 (I1246597,I1246793,I1246660);
not I_73193 (I1246824,I1054463);
nand I_73194 (I1246841,I1246824,I1054475);
nor I_73195 (I1246858,I1054463,I1054481);
not I_73196 (I1246875,I1246858);
nand I_73197 (I1246600,I1246742,I1246875);
DFFARX1 I_73198 (I1246858,I2507,I1246626,I1246615,);
nor I_73199 (I1246920,I1054466,I1054469);
nor I_73200 (I1246937,I1246920,I1054472);
and I_73201 (I1246954,I1246937,I1246841);
DFFARX1 I_73202 (I1246954,I2507,I1246626,I1246612,);
nor I_73203 (I1246609,I1246920,I1246776);
or I_73204 (I1246606,I1246858,I1246920);
nor I_73205 (I1247013,I1054466,I1054463);
DFFARX1 I_73206 (I1247013,I2507,I1246626,I1247039,);
not I_73207 (I1247047,I1247039);
nand I_73208 (I1247064,I1247047,I1246725);
nor I_73209 (I1247081,I1247064,I1054472);
DFFARX1 I_73210 (I1247081,I2507,I1246626,I1246594,);
nor I_73211 (I1247112,I1247047,I1246776);
nor I_73212 (I1246603,I1246920,I1247112);
not I_73213 (I1247170,I2514);
DFFARX1 I_73214 (I443079,I2507,I1247170,I1247196,);
nand I_73215 (I1247204,I1247196,I443076);
DFFARX1 I_73216 (I443055,I2507,I1247170,I1247230,);
DFFARX1 I_73217 (I1247230,I2507,I1247170,I1247247,);
not I_73218 (I1247162,I1247247);
not I_73219 (I1247269,I443070);
nor I_73220 (I1247286,I443070,I443073);
not I_73221 (I1247303,I443064);
nand I_73222 (I1247320,I1247269,I1247303);
nor I_73223 (I1247337,I443064,I443070);
and I_73224 (I1247141,I1247337,I1247204);
not I_73225 (I1247368,I443061);
nand I_73226 (I1247385,I1247368,I443082);
nor I_73227 (I1247402,I443061,I443058);
not I_73228 (I1247419,I1247402);
nand I_73229 (I1247144,I1247286,I1247419);
DFFARX1 I_73230 (I1247402,I2507,I1247170,I1247159,);
nor I_73231 (I1247464,I443067,I443064);
nor I_73232 (I1247481,I1247464,I443073);
and I_73233 (I1247498,I1247481,I1247385);
DFFARX1 I_73234 (I1247498,I2507,I1247170,I1247156,);
nor I_73235 (I1247153,I1247464,I1247320);
or I_73236 (I1247150,I1247402,I1247464);
nor I_73237 (I1247557,I443067,I443055);
DFFARX1 I_73238 (I1247557,I2507,I1247170,I1247583,);
not I_73239 (I1247591,I1247583);
nand I_73240 (I1247608,I1247591,I1247269);
nor I_73241 (I1247625,I1247608,I443073);
DFFARX1 I_73242 (I1247625,I2507,I1247170,I1247138,);
nor I_73243 (I1247656,I1247591,I1247320);
nor I_73244 (I1247147,I1247464,I1247656);
not I_73245 (I1247714,I2514);
DFFARX1 I_73246 (I606463,I2507,I1247714,I1247740,);
nand I_73247 (I1247748,I1247740,I606451);
DFFARX1 I_73248 (I606457,I2507,I1247714,I1247774,);
DFFARX1 I_73249 (I1247774,I2507,I1247714,I1247791,);
not I_73250 (I1247706,I1247791);
not I_73251 (I1247813,I606442);
nor I_73252 (I1247830,I606442,I606454);
not I_73253 (I1247847,I606445);
nand I_73254 (I1247864,I1247813,I1247847);
nor I_73255 (I1247881,I606445,I606442);
and I_73256 (I1247685,I1247881,I1247748);
not I_73257 (I1247912,I606460);
nand I_73258 (I1247929,I1247912,I606442);
nor I_73259 (I1247946,I606460,I606466);
not I_73260 (I1247963,I1247946);
nand I_73261 (I1247688,I1247830,I1247963);
DFFARX1 I_73262 (I1247946,I2507,I1247714,I1247703,);
nor I_73263 (I1248008,I606448,I606445);
nor I_73264 (I1248025,I1248008,I606454);
and I_73265 (I1248042,I1248025,I1247929);
DFFARX1 I_73266 (I1248042,I2507,I1247714,I1247700,);
nor I_73267 (I1247697,I1248008,I1247864);
or I_73268 (I1247694,I1247946,I1248008);
nor I_73269 (I1248101,I606448,I606445);
DFFARX1 I_73270 (I1248101,I2507,I1247714,I1248127,);
not I_73271 (I1248135,I1248127);
nand I_73272 (I1248152,I1248135,I1247813);
nor I_73273 (I1248169,I1248152,I606454);
DFFARX1 I_73274 (I1248169,I2507,I1247714,I1247682,);
nor I_73275 (I1248200,I1248135,I1247864);
nor I_73276 (I1247691,I1248008,I1248200);
not I_73277 (I1248258,I2514);
DFFARX1 I_73278 (I880777,I2507,I1248258,I1248284,);
nand I_73279 (I1248292,I1248284,I880771);
DFFARX1 I_73280 (I880774,I2507,I1248258,I1248318,);
DFFARX1 I_73281 (I1248318,I2507,I1248258,I1248335,);
not I_73282 (I1248250,I1248335);
not I_73283 (I1248357,I880780);
nor I_73284 (I1248374,I880780,I880774);
not I_73285 (I1248391,I880783);
nand I_73286 (I1248408,I1248357,I1248391);
nor I_73287 (I1248425,I880783,I880780);
and I_73288 (I1248229,I1248425,I1248292);
not I_73289 (I1248456,I880792);
nand I_73290 (I1248473,I1248456,I880786);
nor I_73291 (I1248490,I880792,I880789);
not I_73292 (I1248507,I1248490);
nand I_73293 (I1248232,I1248374,I1248507);
DFFARX1 I_73294 (I1248490,I2507,I1248258,I1248247,);
nor I_73295 (I1248552,I880771,I880783);
nor I_73296 (I1248569,I1248552,I880774);
and I_73297 (I1248586,I1248569,I1248473);
DFFARX1 I_73298 (I1248586,I2507,I1248258,I1248244,);
nor I_73299 (I1248241,I1248552,I1248408);
or I_73300 (I1248238,I1248490,I1248552);
nor I_73301 (I1248645,I880771,I880777);
DFFARX1 I_73302 (I1248645,I2507,I1248258,I1248671,);
not I_73303 (I1248679,I1248671);
nand I_73304 (I1248696,I1248679,I1248357);
nor I_73305 (I1248713,I1248696,I880774);
DFFARX1 I_73306 (I1248713,I2507,I1248258,I1248226,);
nor I_73307 (I1248744,I1248679,I1248408);
nor I_73308 (I1248235,I1248552,I1248744);
not I_73309 (I1248802,I2514);
DFFARX1 I_73310 (I428391,I2507,I1248802,I1248828,);
nand I_73311 (I1248836,I1248828,I428388);
DFFARX1 I_73312 (I428367,I2507,I1248802,I1248862,);
DFFARX1 I_73313 (I1248862,I2507,I1248802,I1248879,);
not I_73314 (I1248794,I1248879);
not I_73315 (I1248901,I428382);
nor I_73316 (I1248918,I428382,I428385);
not I_73317 (I1248935,I428376);
nand I_73318 (I1248952,I1248901,I1248935);
nor I_73319 (I1248969,I428376,I428382);
and I_73320 (I1248773,I1248969,I1248836);
not I_73321 (I1249000,I428373);
nand I_73322 (I1249017,I1249000,I428394);
nor I_73323 (I1249034,I428373,I428370);
not I_73324 (I1249051,I1249034);
nand I_73325 (I1248776,I1248918,I1249051);
DFFARX1 I_73326 (I1249034,I2507,I1248802,I1248791,);
nor I_73327 (I1249096,I428379,I428376);
nor I_73328 (I1249113,I1249096,I428385);
and I_73329 (I1249130,I1249113,I1249017);
DFFARX1 I_73330 (I1249130,I2507,I1248802,I1248788,);
nor I_73331 (I1248785,I1249096,I1248952);
or I_73332 (I1248782,I1249034,I1249096);
nor I_73333 (I1249189,I428379,I428367);
DFFARX1 I_73334 (I1249189,I2507,I1248802,I1249215,);
not I_73335 (I1249223,I1249215);
nand I_73336 (I1249240,I1249223,I1248901);
nor I_73337 (I1249257,I1249240,I428385);
DFFARX1 I_73338 (I1249257,I2507,I1248802,I1248770,);
nor I_73339 (I1249288,I1249223,I1248952);
nor I_73340 (I1248779,I1249096,I1249288);
not I_73341 (I1249346,I2514);
DFFARX1 I_73342 (I124972,I2507,I1249346,I1249372,);
nand I_73343 (I1249380,I1249372,I124954);
DFFARX1 I_73344 (I124951,I2507,I1249346,I1249406,);
DFFARX1 I_73345 (I1249406,I2507,I1249346,I1249423,);
not I_73346 (I1249338,I1249423);
not I_73347 (I1249445,I124969);
nor I_73348 (I1249462,I124969,I124963);
not I_73349 (I1249479,I124951);
nand I_73350 (I1249496,I1249445,I1249479);
nor I_73351 (I1249513,I124951,I124969);
and I_73352 (I1249317,I1249513,I1249380);
not I_73353 (I1249544,I124960);
nand I_73354 (I1249561,I1249544,I124966);
nor I_73355 (I1249578,I124960,I124954);
not I_73356 (I1249595,I1249578);
nand I_73357 (I1249320,I1249462,I1249595);
DFFARX1 I_73358 (I1249578,I2507,I1249346,I1249335,);
nor I_73359 (I1249640,I124957,I124951);
nor I_73360 (I1249657,I1249640,I124963);
and I_73361 (I1249674,I1249657,I1249561);
DFFARX1 I_73362 (I1249674,I2507,I1249346,I1249332,);
nor I_73363 (I1249329,I1249640,I1249496);
or I_73364 (I1249326,I1249578,I1249640);
nor I_73365 (I1249733,I124957,I124975);
DFFARX1 I_73366 (I1249733,I2507,I1249346,I1249759,);
not I_73367 (I1249767,I1249759);
nand I_73368 (I1249784,I1249767,I1249445);
nor I_73369 (I1249801,I1249784,I124963);
DFFARX1 I_73370 (I1249801,I2507,I1249346,I1249314,);
nor I_73371 (I1249832,I1249767,I1249496);
nor I_73372 (I1249323,I1249640,I1249832);
not I_73373 (I1249890,I2514);
DFFARX1 I_73374 (I383239,I2507,I1249890,I1249916,);
nand I_73375 (I1249924,I1249916,I383236);
DFFARX1 I_73376 (I383215,I2507,I1249890,I1249950,);
DFFARX1 I_73377 (I1249950,I2507,I1249890,I1249967,);
not I_73378 (I1249882,I1249967);
not I_73379 (I1249989,I383230);
nor I_73380 (I1250006,I383230,I383233);
not I_73381 (I1250023,I383224);
nand I_73382 (I1250040,I1249989,I1250023);
nor I_73383 (I1250057,I383224,I383230);
and I_73384 (I1249861,I1250057,I1249924);
not I_73385 (I1250088,I383221);
nand I_73386 (I1250105,I1250088,I383242);
nor I_73387 (I1250122,I383221,I383218);
not I_73388 (I1250139,I1250122);
nand I_73389 (I1249864,I1250006,I1250139);
DFFARX1 I_73390 (I1250122,I2507,I1249890,I1249879,);
nor I_73391 (I1250184,I383227,I383224);
nor I_73392 (I1250201,I1250184,I383233);
and I_73393 (I1250218,I1250201,I1250105);
DFFARX1 I_73394 (I1250218,I2507,I1249890,I1249876,);
nor I_73395 (I1249873,I1250184,I1250040);
or I_73396 (I1249870,I1250122,I1250184);
nor I_73397 (I1250277,I383227,I383215);
DFFARX1 I_73398 (I1250277,I2507,I1249890,I1250303,);
not I_73399 (I1250311,I1250303);
nand I_73400 (I1250328,I1250311,I1249989);
nor I_73401 (I1250345,I1250328,I383233);
DFFARX1 I_73402 (I1250345,I2507,I1249890,I1249858,);
nor I_73403 (I1250376,I1250311,I1250040);
nor I_73404 (I1249867,I1250184,I1250376);
not I_73405 (I1250434,I2514);
DFFARX1 I_73406 (I1015769,I2507,I1250434,I1250460,);
nand I_73407 (I1250468,I1250460,I1015757);
DFFARX1 I_73408 (I1015751,I2507,I1250434,I1250494,);
DFFARX1 I_73409 (I1250494,I2507,I1250434,I1250511,);
not I_73410 (I1250426,I1250511);
not I_73411 (I1250533,I1015751);
nor I_73412 (I1250550,I1015751,I1015763);
not I_73413 (I1250567,I1015760);
nand I_73414 (I1250584,I1250533,I1250567);
nor I_73415 (I1250601,I1015760,I1015751);
and I_73416 (I1250405,I1250601,I1250468);
not I_73417 (I1250632,I1015754);
nand I_73418 (I1250649,I1250632,I1015766);
nor I_73419 (I1250666,I1015754,I1015772);
not I_73420 (I1250683,I1250666);
nand I_73421 (I1250408,I1250550,I1250683);
DFFARX1 I_73422 (I1250666,I2507,I1250434,I1250423,);
nor I_73423 (I1250728,I1015757,I1015760);
nor I_73424 (I1250745,I1250728,I1015763);
and I_73425 (I1250762,I1250745,I1250649);
DFFARX1 I_73426 (I1250762,I2507,I1250434,I1250420,);
nor I_73427 (I1250417,I1250728,I1250584);
or I_73428 (I1250414,I1250666,I1250728);
nor I_73429 (I1250821,I1015757,I1015754);
DFFARX1 I_73430 (I1250821,I2507,I1250434,I1250847,);
not I_73431 (I1250855,I1250847);
nand I_73432 (I1250872,I1250855,I1250533);
nor I_73433 (I1250889,I1250872,I1015763);
DFFARX1 I_73434 (I1250889,I2507,I1250434,I1250402,);
nor I_73435 (I1250920,I1250855,I1250584);
nor I_73436 (I1250411,I1250728,I1250920);
not I_73437 (I1250978,I2514);
DFFARX1 I_73438 (I862332,I2507,I1250978,I1251004,);
nand I_73439 (I1251012,I1251004,I862326);
DFFARX1 I_73440 (I862329,I2507,I1250978,I1251038,);
DFFARX1 I_73441 (I1251038,I2507,I1250978,I1251055,);
not I_73442 (I1250970,I1251055);
not I_73443 (I1251077,I862335);
nor I_73444 (I1251094,I862335,I862329);
not I_73445 (I1251111,I862338);
nand I_73446 (I1251128,I1251077,I1251111);
nor I_73447 (I1251145,I862338,I862335);
and I_73448 (I1250949,I1251145,I1251012);
not I_73449 (I1251176,I862347);
nand I_73450 (I1251193,I1251176,I862341);
nor I_73451 (I1251210,I862347,I862344);
not I_73452 (I1251227,I1251210);
nand I_73453 (I1250952,I1251094,I1251227);
DFFARX1 I_73454 (I1251210,I2507,I1250978,I1250967,);
nor I_73455 (I1251272,I862326,I862338);
nor I_73456 (I1251289,I1251272,I862329);
and I_73457 (I1251306,I1251289,I1251193);
DFFARX1 I_73458 (I1251306,I2507,I1250978,I1250964,);
nor I_73459 (I1250961,I1251272,I1251128);
or I_73460 (I1250958,I1251210,I1251272);
nor I_73461 (I1251365,I862326,I862332);
DFFARX1 I_73462 (I1251365,I2507,I1250978,I1251391,);
not I_73463 (I1251399,I1251391);
nand I_73464 (I1251416,I1251399,I1251077);
nor I_73465 (I1251433,I1251416,I862329);
DFFARX1 I_73466 (I1251433,I2507,I1250978,I1250946,);
nor I_73467 (I1251464,I1251399,I1251128);
nor I_73468 (I1250955,I1251272,I1251464);
not I_73469 (I1251522,I2514);
DFFARX1 I_73470 (I300267,I2507,I1251522,I1251548,);
nand I_73471 (I1251556,I1251548,I300270);
DFFARX1 I_73472 (I300264,I2507,I1251522,I1251582,);
DFFARX1 I_73473 (I1251582,I2507,I1251522,I1251599,);
not I_73474 (I1251514,I1251599);
not I_73475 (I1251621,I300273);
nor I_73476 (I1251638,I300273,I300258);
not I_73477 (I1251655,I300282);
nand I_73478 (I1251672,I1251621,I1251655);
nor I_73479 (I1251689,I300282,I300273);
and I_73480 (I1251493,I1251689,I1251556);
not I_73481 (I1251720,I300261);
nand I_73482 (I1251737,I1251720,I300279);
nor I_73483 (I1251754,I300261,I300255);
not I_73484 (I1251771,I1251754);
nand I_73485 (I1251496,I1251638,I1251771);
DFFARX1 I_73486 (I1251754,I2507,I1251522,I1251511,);
nor I_73487 (I1251816,I300276,I300282);
nor I_73488 (I1251833,I1251816,I300258);
and I_73489 (I1251850,I1251833,I1251737);
DFFARX1 I_73490 (I1251850,I2507,I1251522,I1251508,);
nor I_73491 (I1251505,I1251816,I1251672);
or I_73492 (I1251502,I1251754,I1251816);
nor I_73493 (I1251909,I300276,I300255);
DFFARX1 I_73494 (I1251909,I2507,I1251522,I1251935,);
not I_73495 (I1251943,I1251935);
nand I_73496 (I1251960,I1251943,I1251621);
nor I_73497 (I1251977,I1251960,I300258);
DFFARX1 I_73498 (I1251977,I2507,I1251522,I1251490,);
nor I_73499 (I1252008,I1251943,I1251672);
nor I_73500 (I1251499,I1251816,I1252008);
not I_73501 (I1252066,I2514);
DFFARX1 I_73502 (I954109,I2507,I1252066,I1252092,);
nand I_73503 (I1252100,I1252092,I954109);
DFFARX1 I_73504 (I954121,I2507,I1252066,I1252126,);
DFFARX1 I_73505 (I1252126,I2507,I1252066,I1252143,);
not I_73506 (I1252058,I1252143);
not I_73507 (I1252165,I954115);
nor I_73508 (I1252182,I954115,I954136);
not I_73509 (I1252199,I954124);
nand I_73510 (I1252216,I1252165,I1252199);
nor I_73511 (I1252233,I954124,I954115);
and I_73512 (I1252037,I1252233,I1252100);
not I_73513 (I1252264,I954118);
nand I_73514 (I1252281,I1252264,I954133);
nor I_73515 (I1252298,I954118,I954127);
not I_73516 (I1252315,I1252298);
nand I_73517 (I1252040,I1252182,I1252315);
DFFARX1 I_73518 (I1252298,I2507,I1252066,I1252055,);
nor I_73519 (I1252360,I954130,I954124);
nor I_73520 (I1252377,I1252360,I954136);
and I_73521 (I1252394,I1252377,I1252281);
DFFARX1 I_73522 (I1252394,I2507,I1252066,I1252052,);
nor I_73523 (I1252049,I1252360,I1252216);
or I_73524 (I1252046,I1252298,I1252360);
nor I_73525 (I1252453,I954130,I954112);
DFFARX1 I_73526 (I1252453,I2507,I1252066,I1252479,);
not I_73527 (I1252487,I1252479);
nand I_73528 (I1252504,I1252487,I1252165);
nor I_73529 (I1252521,I1252504,I954136);
DFFARX1 I_73530 (I1252521,I2507,I1252066,I1252034,);
nor I_73531 (I1252552,I1252487,I1252216);
nor I_73532 (I1252043,I1252360,I1252552);
not I_73533 (I1252610,I2514);
DFFARX1 I_73534 (I924393,I2507,I1252610,I1252636,);
nand I_73535 (I1252644,I1252636,I924393);
DFFARX1 I_73536 (I924405,I2507,I1252610,I1252670,);
DFFARX1 I_73537 (I1252670,I2507,I1252610,I1252687,);
not I_73538 (I1252602,I1252687);
not I_73539 (I1252709,I924399);
nor I_73540 (I1252726,I924399,I924420);
not I_73541 (I1252743,I924408);
nand I_73542 (I1252760,I1252709,I1252743);
nor I_73543 (I1252777,I924408,I924399);
and I_73544 (I1252581,I1252777,I1252644);
not I_73545 (I1252808,I924402);
nand I_73546 (I1252825,I1252808,I924417);
nor I_73547 (I1252842,I924402,I924411);
not I_73548 (I1252859,I1252842);
nand I_73549 (I1252584,I1252726,I1252859);
DFFARX1 I_73550 (I1252842,I2507,I1252610,I1252599,);
nor I_73551 (I1252904,I924414,I924408);
nor I_73552 (I1252921,I1252904,I924420);
and I_73553 (I1252938,I1252921,I1252825);
DFFARX1 I_73554 (I1252938,I2507,I1252610,I1252596,);
nor I_73555 (I1252593,I1252904,I1252760);
or I_73556 (I1252590,I1252842,I1252904);
nor I_73557 (I1252997,I924414,I924396);
DFFARX1 I_73558 (I1252997,I2507,I1252610,I1253023,);
not I_73559 (I1253031,I1253023);
nand I_73560 (I1253048,I1253031,I1252709);
nor I_73561 (I1253065,I1253048,I924420);
DFFARX1 I_73562 (I1253065,I2507,I1252610,I1252578,);
nor I_73563 (I1253096,I1253031,I1252760);
nor I_73564 (I1252587,I1252904,I1253096);
not I_73565 (I1253154,I2514);
DFFARX1 I_73566 (I60151,I2507,I1253154,I1253180,);
nand I_73567 (I1253188,I1253180,I60133);
DFFARX1 I_73568 (I60130,I2507,I1253154,I1253214,);
DFFARX1 I_73569 (I1253214,I2507,I1253154,I1253231,);
not I_73570 (I1253146,I1253231);
not I_73571 (I1253253,I60148);
nor I_73572 (I1253270,I60148,I60142);
not I_73573 (I1253287,I60130);
nand I_73574 (I1253304,I1253253,I1253287);
nor I_73575 (I1253321,I60130,I60148);
and I_73576 (I1253125,I1253321,I1253188);
not I_73577 (I1253352,I60139);
nand I_73578 (I1253369,I1253352,I60145);
nor I_73579 (I1253386,I60139,I60133);
not I_73580 (I1253403,I1253386);
nand I_73581 (I1253128,I1253270,I1253403);
DFFARX1 I_73582 (I1253386,I2507,I1253154,I1253143,);
nor I_73583 (I1253448,I60136,I60130);
nor I_73584 (I1253465,I1253448,I60142);
and I_73585 (I1253482,I1253465,I1253369);
DFFARX1 I_73586 (I1253482,I2507,I1253154,I1253140,);
nor I_73587 (I1253137,I1253448,I1253304);
or I_73588 (I1253134,I1253386,I1253448);
nor I_73589 (I1253541,I60136,I60154);
DFFARX1 I_73590 (I1253541,I2507,I1253154,I1253567,);
not I_73591 (I1253575,I1253567);
nand I_73592 (I1253592,I1253575,I1253253);
nor I_73593 (I1253609,I1253592,I60142);
DFFARX1 I_73594 (I1253609,I2507,I1253154,I1253122,);
nor I_73595 (I1253640,I1253575,I1253304);
nor I_73596 (I1253131,I1253448,I1253640);
not I_73597 (I1253698,I2514);
DFFARX1 I_73598 (I1087872,I2507,I1253698,I1253724,);
nand I_73599 (I1253732,I1253724,I1087851);
DFFARX1 I_73600 (I1087848,I2507,I1253698,I1253758,);
DFFARX1 I_73601 (I1253758,I2507,I1253698,I1253775,);
not I_73602 (I1253690,I1253775);
not I_73603 (I1253797,I1087860);
nor I_73604 (I1253814,I1087860,I1087869);
not I_73605 (I1253831,I1087857);
nand I_73606 (I1253848,I1253797,I1253831);
nor I_73607 (I1253865,I1087857,I1087860);
and I_73608 (I1253669,I1253865,I1253732);
not I_73609 (I1253896,I1087866);
nand I_73610 (I1253913,I1253896,I1087863);
nor I_73611 (I1253930,I1087866,I1087848);
not I_73612 (I1253947,I1253930);
nand I_73613 (I1253672,I1253814,I1253947);
DFFARX1 I_73614 (I1253930,I2507,I1253698,I1253687,);
nor I_73615 (I1253992,I1087851,I1087857);
nor I_73616 (I1254009,I1253992,I1087869);
and I_73617 (I1254026,I1254009,I1253913);
DFFARX1 I_73618 (I1254026,I2507,I1253698,I1253684,);
nor I_73619 (I1253681,I1253992,I1253848);
or I_73620 (I1253678,I1253930,I1253992);
nor I_73621 (I1254085,I1087851,I1087854);
DFFARX1 I_73622 (I1254085,I2507,I1253698,I1254111,);
not I_73623 (I1254119,I1254111);
nand I_73624 (I1254136,I1254119,I1253797);
nor I_73625 (I1254153,I1254136,I1087869);
DFFARX1 I_73626 (I1254153,I2507,I1253698,I1253666,);
nor I_73627 (I1254184,I1254119,I1253848);
nor I_73628 (I1253675,I1253992,I1254184);
not I_73629 (I1254242,I2514);
DFFARX1 I_73630 (I17979,I2507,I1254242,I1254268,);
nand I_73631 (I1254276,I1254268,I17973);
DFFARX1 I_73632 (I17994,I2507,I1254242,I1254302,);
DFFARX1 I_73633 (I1254302,I2507,I1254242,I1254319,);
not I_73634 (I1254234,I1254319);
not I_73635 (I1254341,I17982);
nor I_73636 (I1254358,I17982,I17991);
not I_73637 (I1254375,I17970);
nand I_73638 (I1254392,I1254341,I1254375);
nor I_73639 (I1254409,I17970,I17982);
and I_73640 (I1254213,I1254409,I1254276);
not I_73641 (I1254440,I17988);
nand I_73642 (I1254457,I1254440,I17976);
nor I_73643 (I1254474,I17988,I17970);
not I_73644 (I1254491,I1254474);
nand I_73645 (I1254216,I1254358,I1254491);
DFFARX1 I_73646 (I1254474,I2507,I1254242,I1254231,);
nor I_73647 (I1254536,I17973,I17970);
nor I_73648 (I1254553,I1254536,I17991);
and I_73649 (I1254570,I1254553,I1254457);
DFFARX1 I_73650 (I1254570,I2507,I1254242,I1254228,);
nor I_73651 (I1254225,I1254536,I1254392);
or I_73652 (I1254222,I1254474,I1254536);
nor I_73653 (I1254629,I17973,I17985);
DFFARX1 I_73654 (I1254629,I2507,I1254242,I1254655,);
not I_73655 (I1254663,I1254655);
nand I_73656 (I1254680,I1254663,I1254341);
nor I_73657 (I1254697,I1254680,I17991);
DFFARX1 I_73658 (I1254697,I2507,I1254242,I1254210,);
nor I_73659 (I1254728,I1254663,I1254392);
nor I_73660 (I1254219,I1254536,I1254728);
not I_73661 (I1254786,I2514);
DFFARX1 I_73662 (I276546,I2507,I1254786,I1254812,);
nand I_73663 (I1254820,I1254812,I276567);
not I_73664 (I1254837,I1254820);
DFFARX1 I_73665 (I276561,I2507,I1254786,I1254863,);
not I_73666 (I1254871,I1254863);
not I_73667 (I1254888,I276549);
or I_73668 (I1254905,I276564,I276549);
nor I_73669 (I1254922,I276564,I276549);
or I_73670 (I1254939,I276555,I276564);
DFFARX1 I_73671 (I1254939,I2507,I1254786,I1254778,);
not I_73672 (I1254970,I276543);
nand I_73673 (I1254987,I1254970,I276540);
nand I_73674 (I1255004,I1254888,I1254987);
and I_73675 (I1254757,I1254871,I1255004);
nor I_73676 (I1255035,I276543,I276552);
and I_73677 (I1255052,I1254871,I1255035);
nor I_73678 (I1254763,I1254837,I1255052);
DFFARX1 I_73679 (I1255035,I2507,I1254786,I1255092,);
not I_73680 (I1255100,I1255092);
nor I_73681 (I1254772,I1254871,I1255100);
or I_73682 (I1255131,I1254939,I276558);
nor I_73683 (I1255148,I276558,I276555);
nand I_73684 (I1255165,I1255004,I1255148);
nand I_73685 (I1255182,I1255131,I1255165);
DFFARX1 I_73686 (I1255182,I2507,I1254786,I1254775,);
nor I_73687 (I1255213,I1255148,I1254905);
DFFARX1 I_73688 (I1255213,I2507,I1254786,I1254754,);
nor I_73689 (I1255244,I276558,I276540);
DFFARX1 I_73690 (I1255244,I2507,I1254786,I1255270,);
DFFARX1 I_73691 (I1255270,I2507,I1254786,I1254769,);
not I_73692 (I1255292,I1255270);
nand I_73693 (I1254766,I1255292,I1254820);
nand I_73694 (I1254760,I1255292,I1254922);
not I_73695 (I1255364,I2514);
DFFARX1 I_73696 (I1187860,I2507,I1255364,I1255390,);
nand I_73697 (I1255398,I1255390,I1187845);
not I_73698 (I1255415,I1255398);
DFFARX1 I_73699 (I1187848,I2507,I1255364,I1255441,);
not I_73700 (I1255449,I1255441);
not I_73701 (I1255466,I1187863);
or I_73702 (I1255483,I1187866,I1187863);
nor I_73703 (I1255500,I1187866,I1187863);
or I_73704 (I1255517,I1187842,I1187866);
DFFARX1 I_73705 (I1255517,I2507,I1255364,I1255356,);
not I_73706 (I1255548,I1187854);
nand I_73707 (I1255565,I1255548,I1187857);
nand I_73708 (I1255582,I1255466,I1255565);
and I_73709 (I1255335,I1255449,I1255582);
nor I_73710 (I1255613,I1187854,I1187851);
and I_73711 (I1255630,I1255449,I1255613);
nor I_73712 (I1255341,I1255415,I1255630);
DFFARX1 I_73713 (I1255613,I2507,I1255364,I1255670,);
not I_73714 (I1255678,I1255670);
nor I_73715 (I1255350,I1255449,I1255678);
or I_73716 (I1255709,I1255517,I1187842);
nor I_73717 (I1255726,I1187842,I1187842);
nand I_73718 (I1255743,I1255582,I1255726);
nand I_73719 (I1255760,I1255709,I1255743);
DFFARX1 I_73720 (I1255760,I2507,I1255364,I1255353,);
nor I_73721 (I1255791,I1255726,I1255483);
DFFARX1 I_73722 (I1255791,I2507,I1255364,I1255332,);
nor I_73723 (I1255822,I1187842,I1187845);
DFFARX1 I_73724 (I1255822,I2507,I1255364,I1255848,);
DFFARX1 I_73725 (I1255848,I2507,I1255364,I1255347,);
not I_73726 (I1255870,I1255848);
nand I_73727 (I1255344,I1255870,I1255398);
nand I_73728 (I1255338,I1255870,I1255500);
not I_73729 (I1255942,I2514);
DFFARX1 I_73730 (I146675,I2507,I1255942,I1255968,);
nand I_73731 (I1255976,I1255968,I146684);
not I_73732 (I1255993,I1255976);
DFFARX1 I_73733 (I146666,I2507,I1255942,I1256019,);
not I_73734 (I1256027,I1256019);
not I_73735 (I1256044,I146672);
or I_73736 (I1256061,I146681,I146672);
nor I_73737 (I1256078,I146681,I146672);
or I_73738 (I1256095,I146669,I146681);
DFFARX1 I_73739 (I1256095,I2507,I1255942,I1255934,);
not I_73740 (I1256126,I146687);
nand I_73741 (I1256143,I1256126,I146660);
nand I_73742 (I1256160,I1256044,I1256143);
and I_73743 (I1255913,I1256027,I1256160);
nor I_73744 (I1256191,I146687,I146663);
and I_73745 (I1256208,I1256027,I1256191);
nor I_73746 (I1255919,I1255993,I1256208);
DFFARX1 I_73747 (I1256191,I2507,I1255942,I1256248,);
not I_73748 (I1256256,I1256248);
nor I_73749 (I1255928,I1256027,I1256256);
or I_73750 (I1256287,I1256095,I146678);
nor I_73751 (I1256304,I146678,I146669);
nand I_73752 (I1256321,I1256160,I1256304);
nand I_73753 (I1256338,I1256287,I1256321);
DFFARX1 I_73754 (I1256338,I2507,I1255942,I1255931,);
nor I_73755 (I1256369,I1256304,I1256061);
DFFARX1 I_73756 (I1256369,I2507,I1255942,I1255910,);
nor I_73757 (I1256400,I146678,I146660);
DFFARX1 I_73758 (I1256400,I2507,I1255942,I1256426,);
DFFARX1 I_73759 (I1256426,I2507,I1255942,I1255925,);
not I_73760 (I1256448,I1256426);
nand I_73761 (I1255922,I1256448,I1255976);
nand I_73762 (I1255916,I1256448,I1256078);
not I_73763 (I1256520,I2514);
DFFARX1 I_73764 (I803832,I2507,I1256520,I1256546,);
nand I_73765 (I1256554,I1256546,I803832);
not I_73766 (I1256571,I1256554);
DFFARX1 I_73767 (I803838,I2507,I1256520,I1256597,);
not I_73768 (I1256605,I1256597);
not I_73769 (I1256622,I803850);
or I_73770 (I1256639,I803835,I803850);
nor I_73771 (I1256656,I803835,I803850);
or I_73772 (I1256673,I803829,I803835);
DFFARX1 I_73773 (I1256673,I2507,I1256520,I1256512,);
not I_73774 (I1256704,I803847);
nand I_73775 (I1256721,I1256704,I803841);
nand I_73776 (I1256738,I1256622,I1256721);
and I_73777 (I1256491,I1256605,I1256738);
nor I_73778 (I1256769,I803847,I803829);
and I_73779 (I1256786,I1256605,I1256769);
nor I_73780 (I1256497,I1256571,I1256786);
DFFARX1 I_73781 (I1256769,I2507,I1256520,I1256826,);
not I_73782 (I1256834,I1256826);
nor I_73783 (I1256506,I1256605,I1256834);
or I_73784 (I1256865,I1256673,I803844);
nor I_73785 (I1256882,I803844,I803829);
nand I_73786 (I1256899,I1256738,I1256882);
nand I_73787 (I1256916,I1256865,I1256899);
DFFARX1 I_73788 (I1256916,I2507,I1256520,I1256509,);
nor I_73789 (I1256947,I1256882,I1256639);
DFFARX1 I_73790 (I1256947,I2507,I1256520,I1256488,);
nor I_73791 (I1256978,I803844,I803835);
DFFARX1 I_73792 (I1256978,I2507,I1256520,I1257004,);
DFFARX1 I_73793 (I1257004,I2507,I1256520,I1256503,);
not I_73794 (I1257026,I1257004);
nand I_73795 (I1256500,I1257026,I1256554);
nand I_73796 (I1256494,I1257026,I1256656);
not I_73797 (I1257098,I2514);
DFFARX1 I_73798 (I212110,I2507,I1257098,I1257124,);
nand I_73799 (I1257132,I1257124,I212113);
not I_73800 (I1257149,I1257132);
DFFARX1 I_73801 (I212122,I2507,I1257098,I1257175,);
not I_73802 (I1257183,I1257175);
not I_73803 (I1257200,I212125);
or I_73804 (I1257217,I212116,I212125);
nor I_73805 (I1257234,I212116,I212125);
or I_73806 (I1257251,I212128,I212116);
DFFARX1 I_73807 (I1257251,I2507,I1257098,I1257090,);
not I_73808 (I1257282,I212113);
nand I_73809 (I1257299,I1257282,I212119);
nand I_73810 (I1257316,I1257200,I1257299);
and I_73811 (I1257069,I1257183,I1257316);
nor I_73812 (I1257347,I212113,I212131);
and I_73813 (I1257364,I1257183,I1257347);
nor I_73814 (I1257075,I1257149,I1257364);
DFFARX1 I_73815 (I1257347,I2507,I1257098,I1257404,);
not I_73816 (I1257412,I1257404);
nor I_73817 (I1257084,I1257183,I1257412);
or I_73818 (I1257443,I1257251,I212110);
nor I_73819 (I1257460,I212110,I212128);
nand I_73820 (I1257477,I1257316,I1257460);
nand I_73821 (I1257494,I1257443,I1257477);
DFFARX1 I_73822 (I1257494,I2507,I1257098,I1257087,);
nor I_73823 (I1257525,I1257460,I1257217);
DFFARX1 I_73824 (I1257525,I2507,I1257098,I1257066,);
nor I_73825 (I1257556,I212110,I212134);
DFFARX1 I_73826 (I1257556,I2507,I1257098,I1257582,);
DFFARX1 I_73827 (I1257582,I2507,I1257098,I1257081,);
not I_73828 (I1257604,I1257582);
nand I_73829 (I1257078,I1257604,I1257132);
nand I_73830 (I1257072,I1257604,I1257234);
not I_73831 (I1257676,I2514);
DFFARX1 I_73832 (I854951,I2507,I1257676,I1257702,);
nand I_73833 (I1257710,I1257702,I854951);
not I_73834 (I1257727,I1257710);
DFFARX1 I_73835 (I854957,I2507,I1257676,I1257753,);
not I_73836 (I1257761,I1257753);
not I_73837 (I1257778,I854969);
or I_73838 (I1257795,I854954,I854969);
nor I_73839 (I1257812,I854954,I854969);
or I_73840 (I1257829,I854948,I854954);
DFFARX1 I_73841 (I1257829,I2507,I1257676,I1257668,);
not I_73842 (I1257860,I854966);
nand I_73843 (I1257877,I1257860,I854960);
nand I_73844 (I1257894,I1257778,I1257877);
and I_73845 (I1257647,I1257761,I1257894);
nor I_73846 (I1257925,I854966,I854948);
and I_73847 (I1257942,I1257761,I1257925);
nor I_73848 (I1257653,I1257727,I1257942);
DFFARX1 I_73849 (I1257925,I2507,I1257676,I1257982,);
not I_73850 (I1257990,I1257982);
nor I_73851 (I1257662,I1257761,I1257990);
or I_73852 (I1258021,I1257829,I854963);
nor I_73853 (I1258038,I854963,I854948);
nand I_73854 (I1258055,I1257894,I1258038);
nand I_73855 (I1258072,I1258021,I1258055);
DFFARX1 I_73856 (I1258072,I2507,I1257676,I1257665,);
nor I_73857 (I1258103,I1258038,I1257795);
DFFARX1 I_73858 (I1258103,I2507,I1257676,I1257644,);
nor I_73859 (I1258134,I854963,I854954);
DFFARX1 I_73860 (I1258134,I2507,I1257676,I1258160,);
DFFARX1 I_73861 (I1258160,I2507,I1257676,I1257659,);
not I_73862 (I1258182,I1258160);
nand I_73863 (I1257656,I1258182,I1257710);
nand I_73864 (I1257650,I1258182,I1257812);
not I_73865 (I1258254,I2514);
DFFARX1 I_73866 (I634186,I2507,I1258254,I1258280,);
nand I_73867 (I1258288,I1258280,I634189);
not I_73868 (I1258305,I1258288);
DFFARX1 I_73869 (I634201,I2507,I1258254,I1258331,);
not I_73870 (I1258339,I1258331);
not I_73871 (I1258356,I634186);
or I_73872 (I1258373,I634195,I634186);
nor I_73873 (I1258390,I634195,I634186);
or I_73874 (I1258407,I634204,I634195);
DFFARX1 I_73875 (I1258407,I2507,I1258254,I1258246,);
not I_73876 (I1258438,I634207);
nand I_73877 (I1258455,I1258438,I634189);
nand I_73878 (I1258472,I1258356,I1258455);
and I_73879 (I1258225,I1258339,I1258472);
nor I_73880 (I1258503,I634207,I634192);
and I_73881 (I1258520,I1258339,I1258503);
nor I_73882 (I1258231,I1258305,I1258520);
DFFARX1 I_73883 (I1258503,I2507,I1258254,I1258560,);
not I_73884 (I1258568,I1258560);
nor I_73885 (I1258240,I1258339,I1258568);
or I_73886 (I1258599,I1258407,I634198);
nor I_73887 (I1258616,I634198,I634204);
nand I_73888 (I1258633,I1258472,I1258616);
nand I_73889 (I1258650,I1258599,I1258633);
DFFARX1 I_73890 (I1258650,I2507,I1258254,I1258243,);
nor I_73891 (I1258681,I1258616,I1258373);
DFFARX1 I_73892 (I1258681,I2507,I1258254,I1258222,);
nor I_73893 (I1258712,I634198,I634210);
DFFARX1 I_73894 (I1258712,I2507,I1258254,I1258738,);
DFFARX1 I_73895 (I1258738,I2507,I1258254,I1258237,);
not I_73896 (I1258760,I1258738);
nand I_73897 (I1258234,I1258760,I1258288);
nand I_73898 (I1258228,I1258760,I1258390);
not I_73899 (I1258832,I2514);
DFFARX1 I_73900 (I667710,I2507,I1258832,I1258858,);
nand I_73901 (I1258866,I1258858,I667713);
not I_73902 (I1258883,I1258866);
DFFARX1 I_73903 (I667725,I2507,I1258832,I1258909,);
not I_73904 (I1258917,I1258909);
not I_73905 (I1258934,I667710);
or I_73906 (I1258951,I667719,I667710);
nor I_73907 (I1258968,I667719,I667710);
or I_73908 (I1258985,I667728,I667719);
DFFARX1 I_73909 (I1258985,I2507,I1258832,I1258824,);
not I_73910 (I1259016,I667731);
nand I_73911 (I1259033,I1259016,I667713);
nand I_73912 (I1259050,I1258934,I1259033);
and I_73913 (I1258803,I1258917,I1259050);
nor I_73914 (I1259081,I667731,I667716);
and I_73915 (I1259098,I1258917,I1259081);
nor I_73916 (I1258809,I1258883,I1259098);
DFFARX1 I_73917 (I1259081,I2507,I1258832,I1259138,);
not I_73918 (I1259146,I1259138);
nor I_73919 (I1258818,I1258917,I1259146);
or I_73920 (I1259177,I1258985,I667722);
nor I_73921 (I1259194,I667722,I667728);
nand I_73922 (I1259211,I1259050,I1259194);
nand I_73923 (I1259228,I1259177,I1259211);
DFFARX1 I_73924 (I1259228,I2507,I1258832,I1258821,);
nor I_73925 (I1259259,I1259194,I1258951);
DFFARX1 I_73926 (I1259259,I2507,I1258832,I1258800,);
nor I_73927 (I1259290,I667722,I667734);
DFFARX1 I_73928 (I1259290,I2507,I1258832,I1259316,);
DFFARX1 I_73929 (I1259316,I2507,I1258832,I1258815,);
not I_73930 (I1259338,I1259316);
nand I_73931 (I1258812,I1259338,I1258866);
nand I_73932 (I1258806,I1259338,I1258968);
not I_73933 (I1259410,I2514);
DFFARX1 I_73934 (I968973,I2507,I1259410,I1259436,);
nand I_73935 (I1259444,I1259436,I968994);
not I_73936 (I1259461,I1259444);
DFFARX1 I_73937 (I968967,I2507,I1259410,I1259487,);
not I_73938 (I1259495,I1259487);
not I_73939 (I1259512,I968988);
or I_73940 (I1259529,I968979,I968988);
nor I_73941 (I1259546,I968979,I968988);
or I_73942 (I1259563,I968982,I968979);
DFFARX1 I_73943 (I1259563,I2507,I1259410,I1259402,);
not I_73944 (I1259594,I968970);
nand I_73945 (I1259611,I1259594,I968985);
nand I_73946 (I1259628,I1259512,I1259611);
and I_73947 (I1259381,I1259495,I1259628);
nor I_73948 (I1259659,I968970,I968967);
and I_73949 (I1259676,I1259495,I1259659);
nor I_73950 (I1259387,I1259461,I1259676);
DFFARX1 I_73951 (I1259659,I2507,I1259410,I1259716,);
not I_73952 (I1259724,I1259716);
nor I_73953 (I1259396,I1259495,I1259724);
or I_73954 (I1259755,I1259563,I968991);
nor I_73955 (I1259772,I968991,I968982);
nand I_73956 (I1259789,I1259628,I1259772);
nand I_73957 (I1259806,I1259755,I1259789);
DFFARX1 I_73958 (I1259806,I2507,I1259410,I1259399,);
nor I_73959 (I1259837,I1259772,I1259529);
DFFARX1 I_73960 (I1259837,I2507,I1259410,I1259378,);
nor I_73961 (I1259868,I968991,I968976);
DFFARX1 I_73962 (I1259868,I2507,I1259410,I1259894,);
DFFARX1 I_73963 (I1259894,I2507,I1259410,I1259393,);
not I_73964 (I1259916,I1259894);
nand I_73965 (I1259390,I1259916,I1259444);
nand I_73966 (I1259384,I1259916,I1259546);
not I_73967 (I1259988,I2514);
DFFARX1 I_73968 (I401714,I2507,I1259988,I1260014,);
nand I_73969 (I1260022,I1260014,I401723);
not I_73970 (I1260039,I1260022);
DFFARX1 I_73971 (I401711,I2507,I1259988,I1260065,);
not I_73972 (I1260073,I1260065);
not I_73973 (I1260090,I401717);
or I_73974 (I1260107,I401711,I401717);
nor I_73975 (I1260124,I401711,I401717);
or I_73976 (I1260141,I401726,I401711);
DFFARX1 I_73977 (I1260141,I2507,I1259988,I1259980,);
not I_73978 (I1260172,I401720);
nand I_73979 (I1260189,I1260172,I401735);
nand I_73980 (I1260206,I1260090,I1260189);
and I_73981 (I1259959,I1260073,I1260206);
nor I_73982 (I1260237,I401720,I401738);
and I_73983 (I1260254,I1260073,I1260237);
nor I_73984 (I1259965,I1260039,I1260254);
DFFARX1 I_73985 (I1260237,I2507,I1259988,I1260294,);
not I_73986 (I1260302,I1260294);
nor I_73987 (I1259974,I1260073,I1260302);
or I_73988 (I1260333,I1260141,I401729);
nor I_73989 (I1260350,I401729,I401726);
nand I_73990 (I1260367,I1260206,I1260350);
nand I_73991 (I1260384,I1260333,I1260367);
DFFARX1 I_73992 (I1260384,I2507,I1259988,I1259977,);
nor I_73993 (I1260415,I1260350,I1260107);
DFFARX1 I_73994 (I1260415,I2507,I1259988,I1259956,);
nor I_73995 (I1260446,I401729,I401732);
DFFARX1 I_73996 (I1260446,I2507,I1259988,I1260472,);
DFFARX1 I_73997 (I1260472,I2507,I1259988,I1259971,);
not I_73998 (I1260494,I1260472);
nand I_73999 (I1259968,I1260494,I1260022);
nand I_74000 (I1259962,I1260494,I1260124);
not I_74001 (I1260566,I2514);
DFFARX1 I_74002 (I1297510,I2507,I1260566,I1260592,);
nand I_74003 (I1260600,I1260592,I1297504);
not I_74004 (I1260617,I1260600);
DFFARX1 I_74005 (I1297519,I2507,I1260566,I1260643,);
not I_74006 (I1260651,I1260643);
not I_74007 (I1260668,I1297495);
or I_74008 (I1260685,I1297492,I1297495);
nor I_74009 (I1260702,I1297492,I1297495);
or I_74010 (I1260719,I1297498,I1297492);
DFFARX1 I_74011 (I1260719,I2507,I1260566,I1260558,);
not I_74012 (I1260750,I1297492);
nand I_74013 (I1260767,I1260750,I1297507);
nand I_74014 (I1260784,I1260668,I1260767);
and I_74015 (I1260537,I1260651,I1260784);
nor I_74016 (I1260815,I1297492,I1297501);
and I_74017 (I1260832,I1260651,I1260815);
nor I_74018 (I1260543,I1260617,I1260832);
DFFARX1 I_74019 (I1260815,I2507,I1260566,I1260872,);
not I_74020 (I1260880,I1260872);
nor I_74021 (I1260552,I1260651,I1260880);
or I_74022 (I1260911,I1260719,I1297516);
nor I_74023 (I1260928,I1297516,I1297498);
nand I_74024 (I1260945,I1260784,I1260928);
nand I_74025 (I1260962,I1260911,I1260945);
DFFARX1 I_74026 (I1260962,I2507,I1260566,I1260555,);
nor I_74027 (I1260993,I1260928,I1260685);
DFFARX1 I_74028 (I1260993,I2507,I1260566,I1260534,);
nor I_74029 (I1261024,I1297516,I1297513);
DFFARX1 I_74030 (I1261024,I2507,I1260566,I1261050,);
DFFARX1 I_74031 (I1261050,I2507,I1260566,I1260549,);
not I_74032 (I1261072,I1261050);
nand I_74033 (I1260546,I1261072,I1260600);
nand I_74034 (I1260540,I1261072,I1260702);
not I_74035 (I1261144,I2514);
DFFARX1 I_74036 (I1187282,I2507,I1261144,I1261170,);
nand I_74037 (I1261178,I1261170,I1187267);
not I_74038 (I1261195,I1261178);
DFFARX1 I_74039 (I1187270,I2507,I1261144,I1261221,);
not I_74040 (I1261229,I1261221);
not I_74041 (I1261246,I1187285);
or I_74042 (I1261263,I1187288,I1187285);
nor I_74043 (I1261280,I1187288,I1187285);
or I_74044 (I1261297,I1187264,I1187288);
DFFARX1 I_74045 (I1261297,I2507,I1261144,I1261136,);
not I_74046 (I1261328,I1187276);
nand I_74047 (I1261345,I1261328,I1187279);
nand I_74048 (I1261362,I1261246,I1261345);
and I_74049 (I1261115,I1261229,I1261362);
nor I_74050 (I1261393,I1187276,I1187273);
and I_74051 (I1261410,I1261229,I1261393);
nor I_74052 (I1261121,I1261195,I1261410);
DFFARX1 I_74053 (I1261393,I2507,I1261144,I1261450,);
not I_74054 (I1261458,I1261450);
nor I_74055 (I1261130,I1261229,I1261458);
or I_74056 (I1261489,I1261297,I1187264);
nor I_74057 (I1261506,I1187264,I1187264);
nand I_74058 (I1261523,I1261362,I1261506);
nand I_74059 (I1261540,I1261489,I1261523);
DFFARX1 I_74060 (I1261540,I2507,I1261144,I1261133,);
nor I_74061 (I1261571,I1261506,I1261263);
DFFARX1 I_74062 (I1261571,I2507,I1261144,I1261112,);
nor I_74063 (I1261602,I1187264,I1187267);
DFFARX1 I_74064 (I1261602,I2507,I1261144,I1261628,);
DFFARX1 I_74065 (I1261628,I2507,I1261144,I1261127,);
not I_74066 (I1261650,I1261628);
nand I_74067 (I1261124,I1261650,I1261178);
nand I_74068 (I1261118,I1261650,I1261280);
not I_74069 (I1261722,I2514);
DFFARX1 I_74070 (I15868,I2507,I1261722,I1261748,);
nand I_74071 (I1261756,I1261748,I15862);
not I_74072 (I1261773,I1261756);
DFFARX1 I_74073 (I15880,I2507,I1261722,I1261799,);
not I_74074 (I1261807,I1261799);
not I_74075 (I1261824,I15883);
or I_74076 (I1261841,I15886,I15883);
nor I_74077 (I1261858,I15886,I15883);
or I_74078 (I1261875,I15871,I15886);
DFFARX1 I_74079 (I1261875,I2507,I1261722,I1261714,);
not I_74080 (I1261906,I15874);
nand I_74081 (I1261923,I1261906,I15877);
nand I_74082 (I1261940,I1261824,I1261923);
and I_74083 (I1261693,I1261807,I1261940);
nor I_74084 (I1261971,I15874,I15865);
and I_74085 (I1261988,I1261807,I1261971);
nor I_74086 (I1261699,I1261773,I1261988);
DFFARX1 I_74087 (I1261971,I2507,I1261722,I1262028,);
not I_74088 (I1262036,I1262028);
nor I_74089 (I1261708,I1261807,I1262036);
or I_74090 (I1262067,I1261875,I15865);
nor I_74091 (I1262084,I15865,I15871);
nand I_74092 (I1262101,I1261940,I1262084);
nand I_74093 (I1262118,I1262067,I1262101);
DFFARX1 I_74094 (I1262118,I2507,I1261722,I1261711,);
nor I_74095 (I1262149,I1262084,I1261841);
DFFARX1 I_74096 (I1262149,I2507,I1261722,I1261690,);
nor I_74097 (I1262180,I15865,I15862);
DFFARX1 I_74098 (I1262180,I2507,I1261722,I1262206,);
DFFARX1 I_74099 (I1262206,I2507,I1261722,I1261705,);
not I_74100 (I1262228,I1262206);
nand I_74101 (I1261702,I1262228,I1261756);
nand I_74102 (I1261696,I1262228,I1261858);
not I_74103 (I1262300,I2514);
DFFARX1 I_74104 (I121274,I2507,I1262300,I1262326,);
nand I_74105 (I1262334,I1262326,I121265);
not I_74106 (I1262351,I1262334);
DFFARX1 I_74107 (I121262,I2507,I1262300,I1262377,);
not I_74108 (I1262385,I1262377);
not I_74109 (I1262402,I121271);
or I_74110 (I1262419,I121262,I121271);
nor I_74111 (I1262436,I121262,I121271);
or I_74112 (I1262453,I121268,I121262);
DFFARX1 I_74113 (I1262453,I2507,I1262300,I1262292,);
not I_74114 (I1262484,I121277);
nand I_74115 (I1262501,I1262484,I121286);
nand I_74116 (I1262518,I1262402,I1262501);
and I_74117 (I1262271,I1262385,I1262518);
nor I_74118 (I1262549,I121277,I121280);
and I_74119 (I1262566,I1262385,I1262549);
nor I_74120 (I1262277,I1262351,I1262566);
DFFARX1 I_74121 (I1262549,I2507,I1262300,I1262606,);
not I_74122 (I1262614,I1262606);
nor I_74123 (I1262286,I1262385,I1262614);
or I_74124 (I1262645,I1262453,I121265);
nor I_74125 (I1262662,I121265,I121268);
nand I_74126 (I1262679,I1262518,I1262662);
nand I_74127 (I1262696,I1262645,I1262679);
DFFARX1 I_74128 (I1262696,I2507,I1262300,I1262289,);
nor I_74129 (I1262727,I1262662,I1262419);
DFFARX1 I_74130 (I1262727,I2507,I1262300,I1262268,);
nor I_74131 (I1262758,I121265,I121283);
DFFARX1 I_74132 (I1262758,I2507,I1262300,I1262784,);
DFFARX1 I_74133 (I1262784,I2507,I1262300,I1262283,);
not I_74134 (I1262806,I1262784);
nand I_74135 (I1262280,I1262806,I1262334);
nand I_74136 (I1262274,I1262806,I1262436);
not I_74137 (I1262878,I2514);
DFFARX1 I_74138 (I790130,I2507,I1262878,I1262904,);
nand I_74139 (I1262912,I1262904,I790130);
not I_74140 (I1262929,I1262912);
DFFARX1 I_74141 (I790136,I2507,I1262878,I1262955,);
not I_74142 (I1262963,I1262955);
not I_74143 (I1262980,I790148);
or I_74144 (I1262997,I790133,I790148);
nor I_74145 (I1263014,I790133,I790148);
or I_74146 (I1263031,I790127,I790133);
DFFARX1 I_74147 (I1263031,I2507,I1262878,I1262870,);
not I_74148 (I1263062,I790145);
nand I_74149 (I1263079,I1263062,I790139);
nand I_74150 (I1263096,I1262980,I1263079);
and I_74151 (I1262849,I1262963,I1263096);
nor I_74152 (I1263127,I790145,I790127);
and I_74153 (I1263144,I1262963,I1263127);
nor I_74154 (I1262855,I1262929,I1263144);
DFFARX1 I_74155 (I1263127,I2507,I1262878,I1263184,);
not I_74156 (I1263192,I1263184);
nor I_74157 (I1262864,I1262963,I1263192);
or I_74158 (I1263223,I1263031,I790142);
nor I_74159 (I1263240,I790142,I790127);
nand I_74160 (I1263257,I1263096,I1263240);
nand I_74161 (I1263274,I1263223,I1263257);
DFFARX1 I_74162 (I1263274,I2507,I1262878,I1262867,);
nor I_74163 (I1263305,I1263240,I1262997);
DFFARX1 I_74164 (I1263305,I2507,I1262878,I1262846,);
nor I_74165 (I1263336,I790142,I790133);
DFFARX1 I_74166 (I1263336,I2507,I1262878,I1263362,);
DFFARX1 I_74167 (I1263362,I2507,I1262878,I1262861,);
not I_74168 (I1263384,I1263362);
nand I_74169 (I1262858,I1263384,I1262912);
nand I_74170 (I1262852,I1263384,I1263014);
not I_74171 (I1263456,I2514);
DFFARX1 I_74172 (I776955,I2507,I1263456,I1263482,);
nand I_74173 (I1263490,I1263482,I776955);
not I_74174 (I1263507,I1263490);
DFFARX1 I_74175 (I776961,I2507,I1263456,I1263533,);
not I_74176 (I1263541,I1263533);
not I_74177 (I1263558,I776973);
or I_74178 (I1263575,I776958,I776973);
nor I_74179 (I1263592,I776958,I776973);
or I_74180 (I1263609,I776952,I776958);
DFFARX1 I_74181 (I1263609,I2507,I1263456,I1263448,);
not I_74182 (I1263640,I776970);
nand I_74183 (I1263657,I1263640,I776964);
nand I_74184 (I1263674,I1263558,I1263657);
and I_74185 (I1263427,I1263541,I1263674);
nor I_74186 (I1263705,I776970,I776952);
and I_74187 (I1263722,I1263541,I1263705);
nor I_74188 (I1263433,I1263507,I1263722);
DFFARX1 I_74189 (I1263705,I2507,I1263456,I1263762,);
not I_74190 (I1263770,I1263762);
nor I_74191 (I1263442,I1263541,I1263770);
or I_74192 (I1263801,I1263609,I776967);
nor I_74193 (I1263818,I776967,I776952);
nand I_74194 (I1263835,I1263674,I1263818);
nand I_74195 (I1263852,I1263801,I1263835);
DFFARX1 I_74196 (I1263852,I2507,I1263456,I1263445,);
nor I_74197 (I1263883,I1263818,I1263575);
DFFARX1 I_74198 (I1263883,I2507,I1263456,I1263424,);
nor I_74199 (I1263914,I776967,I776958);
DFFARX1 I_74200 (I1263914,I2507,I1263456,I1263940,);
DFFARX1 I_74201 (I1263940,I2507,I1263456,I1263439,);
not I_74202 (I1263962,I1263940);
nand I_74203 (I1263436,I1263962,I1263490);
nand I_74204 (I1263430,I1263962,I1263592);
not I_74205 (I1264034,I2514);
DFFARX1 I_74206 (I40637,I2507,I1264034,I1264060,);
nand I_74207 (I1264068,I1264060,I40631);
not I_74208 (I1264085,I1264068);
DFFARX1 I_74209 (I40649,I2507,I1264034,I1264111,);
not I_74210 (I1264119,I1264111);
not I_74211 (I1264136,I40652);
or I_74212 (I1264153,I40655,I40652);
nor I_74213 (I1264170,I40655,I40652);
or I_74214 (I1264187,I40640,I40655);
DFFARX1 I_74215 (I1264187,I2507,I1264034,I1264026,);
not I_74216 (I1264218,I40643);
nand I_74217 (I1264235,I1264218,I40646);
nand I_74218 (I1264252,I1264136,I1264235);
and I_74219 (I1264005,I1264119,I1264252);
nor I_74220 (I1264283,I40643,I40634);
and I_74221 (I1264300,I1264119,I1264283);
nor I_74222 (I1264011,I1264085,I1264300);
DFFARX1 I_74223 (I1264283,I2507,I1264034,I1264340,);
not I_74224 (I1264348,I1264340);
nor I_74225 (I1264020,I1264119,I1264348);
or I_74226 (I1264379,I1264187,I40634);
nor I_74227 (I1264396,I40634,I40640);
nand I_74228 (I1264413,I1264252,I1264396);
nand I_74229 (I1264430,I1264379,I1264413);
DFFARX1 I_74230 (I1264430,I2507,I1264034,I1264023,);
nor I_74231 (I1264461,I1264396,I1264153);
DFFARX1 I_74232 (I1264461,I2507,I1264034,I1264002,);
nor I_74233 (I1264492,I40634,I40631);
DFFARX1 I_74234 (I1264492,I2507,I1264034,I1264518,);
DFFARX1 I_74235 (I1264518,I2507,I1264034,I1264017,);
not I_74236 (I1264540,I1264518);
nand I_74237 (I1264014,I1264540,I1264068);
nand I_74238 (I1264008,I1264540,I1264170);
not I_74239 (I1264612,I2514);
DFFARX1 I_74240 (I153800,I2507,I1264612,I1264638,);
nand I_74241 (I1264646,I1264638,I153803);
not I_74242 (I1264663,I1264646);
DFFARX1 I_74243 (I153812,I2507,I1264612,I1264689,);
not I_74244 (I1264697,I1264689);
not I_74245 (I1264714,I153815);
or I_74246 (I1264731,I153806,I153815);
nor I_74247 (I1264748,I153806,I153815);
or I_74248 (I1264765,I153818,I153806);
DFFARX1 I_74249 (I1264765,I2507,I1264612,I1264604,);
not I_74250 (I1264796,I153803);
nand I_74251 (I1264813,I1264796,I153809);
nand I_74252 (I1264830,I1264714,I1264813);
and I_74253 (I1264583,I1264697,I1264830);
nor I_74254 (I1264861,I153803,I153821);
and I_74255 (I1264878,I1264697,I1264861);
nor I_74256 (I1264589,I1264663,I1264878);
DFFARX1 I_74257 (I1264861,I2507,I1264612,I1264918,);
not I_74258 (I1264926,I1264918);
nor I_74259 (I1264598,I1264697,I1264926);
or I_74260 (I1264957,I1264765,I153800);
nor I_74261 (I1264974,I153800,I153818);
nand I_74262 (I1264991,I1264830,I1264974);
nand I_74263 (I1265008,I1264957,I1264991);
DFFARX1 I_74264 (I1265008,I2507,I1264612,I1264601,);
nor I_74265 (I1265039,I1264974,I1264731);
DFFARX1 I_74266 (I1265039,I2507,I1264612,I1264580,);
nor I_74267 (I1265070,I153800,I153824);
DFFARX1 I_74268 (I1265070,I2507,I1264612,I1265096,);
DFFARX1 I_74269 (I1265096,I2507,I1264612,I1264595,);
not I_74270 (I1265118,I1265096);
nand I_74271 (I1264592,I1265118,I1264646);
nand I_74272 (I1264586,I1265118,I1264748);
not I_74273 (I1265190,I2514);
DFFARX1 I_74274 (I379410,I2507,I1265190,I1265216,);
nand I_74275 (I1265224,I1265216,I379419);
not I_74276 (I1265241,I1265224);
DFFARX1 I_74277 (I379407,I2507,I1265190,I1265267,);
not I_74278 (I1265275,I1265267);
not I_74279 (I1265292,I379413);
or I_74280 (I1265309,I379407,I379413);
nor I_74281 (I1265326,I379407,I379413);
or I_74282 (I1265343,I379422,I379407);
DFFARX1 I_74283 (I1265343,I2507,I1265190,I1265182,);
not I_74284 (I1265374,I379416);
nand I_74285 (I1265391,I1265374,I379431);
nand I_74286 (I1265408,I1265292,I1265391);
and I_74287 (I1265161,I1265275,I1265408);
nor I_74288 (I1265439,I379416,I379434);
and I_74289 (I1265456,I1265275,I1265439);
nor I_74290 (I1265167,I1265241,I1265456);
DFFARX1 I_74291 (I1265439,I2507,I1265190,I1265496,);
not I_74292 (I1265504,I1265496);
nor I_74293 (I1265176,I1265275,I1265504);
or I_74294 (I1265535,I1265343,I379425);
nor I_74295 (I1265552,I379425,I379422);
nand I_74296 (I1265569,I1265408,I1265552);
nand I_74297 (I1265586,I1265535,I1265569);
DFFARX1 I_74298 (I1265586,I2507,I1265190,I1265179,);
nor I_74299 (I1265617,I1265552,I1265309);
DFFARX1 I_74300 (I1265617,I2507,I1265190,I1265158,);
nor I_74301 (I1265648,I379425,I379428);
DFFARX1 I_74302 (I1265648,I2507,I1265190,I1265674,);
DFFARX1 I_74303 (I1265674,I2507,I1265190,I1265173,);
not I_74304 (I1265696,I1265674);
nand I_74305 (I1265170,I1265696,I1265224);
nand I_74306 (I1265164,I1265696,I1265326);
not I_74307 (I1265768,I2514);
DFFARX1 I_74308 (I505394,I2507,I1265768,I1265794,);
nand I_74309 (I1265802,I1265794,I505403);
not I_74310 (I1265819,I1265802);
DFFARX1 I_74311 (I505415,I2507,I1265768,I1265845,);
not I_74312 (I1265853,I1265845);
not I_74313 (I1265870,I505406);
or I_74314 (I1265887,I505400,I505406);
nor I_74315 (I1265904,I505400,I505406);
or I_74316 (I1265921,I505394,I505400);
DFFARX1 I_74317 (I1265921,I2507,I1265768,I1265760,);
not I_74318 (I1265952,I505397);
nand I_74319 (I1265969,I1265952,I505409);
nand I_74320 (I1265986,I1265870,I1265969);
and I_74321 (I1265739,I1265853,I1265986);
nor I_74322 (I1266017,I505397,I505418);
and I_74323 (I1266034,I1265853,I1266017);
nor I_74324 (I1265745,I1265819,I1266034);
DFFARX1 I_74325 (I1266017,I2507,I1265768,I1266074,);
not I_74326 (I1266082,I1266074);
nor I_74327 (I1265754,I1265853,I1266082);
or I_74328 (I1266113,I1265921,I505412);
nor I_74329 (I1266130,I505412,I505394);
nand I_74330 (I1266147,I1265986,I1266130);
nand I_74331 (I1266164,I1266113,I1266147);
DFFARX1 I_74332 (I1266164,I2507,I1265768,I1265757,);
nor I_74333 (I1266195,I1266130,I1265887);
DFFARX1 I_74334 (I1266195,I2507,I1265768,I1265736,);
nor I_74335 (I1266226,I505412,I505397);
DFFARX1 I_74336 (I1266226,I2507,I1265768,I1266252,);
DFFARX1 I_74337 (I1266252,I2507,I1265768,I1265751,);
not I_74338 (I1266274,I1266252);
nand I_74339 (I1265748,I1266274,I1265802);
nand I_74340 (I1265742,I1266274,I1265904);
not I_74341 (I1266346,I2514);
DFFARX1 I_74342 (I530979,I2507,I1266346,I1266372,);
nand I_74343 (I1266380,I1266372,I530988);
not I_74344 (I1266397,I1266380);
DFFARX1 I_74345 (I531000,I2507,I1266346,I1266423,);
not I_74346 (I1266431,I1266423);
not I_74347 (I1266448,I530991);
or I_74348 (I1266465,I530985,I530991);
nor I_74349 (I1266482,I530985,I530991);
or I_74350 (I1266499,I530979,I530985);
DFFARX1 I_74351 (I1266499,I2507,I1266346,I1266338,);
not I_74352 (I1266530,I530982);
nand I_74353 (I1266547,I1266530,I530994);
nand I_74354 (I1266564,I1266448,I1266547);
and I_74355 (I1266317,I1266431,I1266564);
nor I_74356 (I1266595,I530982,I531003);
and I_74357 (I1266612,I1266431,I1266595);
nor I_74358 (I1266323,I1266397,I1266612);
DFFARX1 I_74359 (I1266595,I2507,I1266346,I1266652,);
not I_74360 (I1266660,I1266652);
nor I_74361 (I1266332,I1266431,I1266660);
or I_74362 (I1266691,I1266499,I530997);
nor I_74363 (I1266708,I530997,I530979);
nand I_74364 (I1266725,I1266564,I1266708);
nand I_74365 (I1266742,I1266691,I1266725);
DFFARX1 I_74366 (I1266742,I2507,I1266346,I1266335,);
nor I_74367 (I1266773,I1266708,I1266465);
DFFARX1 I_74368 (I1266773,I2507,I1266346,I1266314,);
nor I_74369 (I1266804,I530997,I530982);
DFFARX1 I_74370 (I1266804,I2507,I1266346,I1266830,);
DFFARX1 I_74371 (I1266830,I2507,I1266346,I1266329,);
not I_74372 (I1266852,I1266830);
nand I_74373 (I1266326,I1266852,I1266380);
nand I_74374 (I1266320,I1266852,I1266482);
not I_74375 (I1266924,I2514);
DFFARX1 I_74376 (I341894,I2507,I1266924,I1266950,);
nand I_74377 (I1266958,I1266950,I341915);
not I_74378 (I1266975,I1266958);
DFFARX1 I_74379 (I341909,I2507,I1266924,I1267001,);
not I_74380 (I1267009,I1267001);
not I_74381 (I1267026,I341897);
or I_74382 (I1267043,I341912,I341897);
nor I_74383 (I1267060,I341912,I341897);
or I_74384 (I1267077,I341903,I341912);
DFFARX1 I_74385 (I1267077,I2507,I1266924,I1266916,);
not I_74386 (I1267108,I341891);
nand I_74387 (I1267125,I1267108,I341888);
nand I_74388 (I1267142,I1267026,I1267125);
and I_74389 (I1266895,I1267009,I1267142);
nor I_74390 (I1267173,I341891,I341900);
and I_74391 (I1267190,I1267009,I1267173);
nor I_74392 (I1266901,I1266975,I1267190);
DFFARX1 I_74393 (I1267173,I2507,I1266924,I1267230,);
not I_74394 (I1267238,I1267230);
nor I_74395 (I1266910,I1267009,I1267238);
or I_74396 (I1267269,I1267077,I341906);
nor I_74397 (I1267286,I341906,I341903);
nand I_74398 (I1267303,I1267142,I1267286);
nand I_74399 (I1267320,I1267269,I1267303);
DFFARX1 I_74400 (I1267320,I2507,I1266924,I1266913,);
nor I_74401 (I1267351,I1267286,I1267043);
DFFARX1 I_74402 (I1267351,I2507,I1266924,I1266892,);
nor I_74403 (I1267382,I341906,I341888);
DFFARX1 I_74404 (I1267382,I2507,I1266924,I1267408,);
DFFARX1 I_74405 (I1267408,I2507,I1266924,I1266907,);
not I_74406 (I1267430,I1267408);
nand I_74407 (I1266904,I1267430,I1266958);
nand I_74408 (I1266898,I1267430,I1267060);
not I_74409 (I1267502,I2514);
DFFARX1 I_74410 (I1159538,I2507,I1267502,I1267528,);
nand I_74411 (I1267536,I1267528,I1159523);
not I_74412 (I1267553,I1267536);
DFFARX1 I_74413 (I1159526,I2507,I1267502,I1267579,);
not I_74414 (I1267587,I1267579);
not I_74415 (I1267604,I1159541);
or I_74416 (I1267621,I1159544,I1159541);
nor I_74417 (I1267638,I1159544,I1159541);
or I_74418 (I1267655,I1159520,I1159544);
DFFARX1 I_74419 (I1267655,I2507,I1267502,I1267494,);
not I_74420 (I1267686,I1159532);
nand I_74421 (I1267703,I1267686,I1159535);
nand I_74422 (I1267720,I1267604,I1267703);
and I_74423 (I1267473,I1267587,I1267720);
nor I_74424 (I1267751,I1159532,I1159529);
and I_74425 (I1267768,I1267587,I1267751);
nor I_74426 (I1267479,I1267553,I1267768);
DFFARX1 I_74427 (I1267751,I2507,I1267502,I1267808,);
not I_74428 (I1267816,I1267808);
nor I_74429 (I1267488,I1267587,I1267816);
or I_74430 (I1267847,I1267655,I1159520);
nor I_74431 (I1267864,I1159520,I1159520);
nand I_74432 (I1267881,I1267720,I1267864);
nand I_74433 (I1267898,I1267847,I1267881);
DFFARX1 I_74434 (I1267898,I2507,I1267502,I1267491,);
nor I_74435 (I1267929,I1267864,I1267621);
DFFARX1 I_74436 (I1267929,I2507,I1267502,I1267470,);
nor I_74437 (I1267960,I1159520,I1159523);
DFFARX1 I_74438 (I1267960,I2507,I1267502,I1267986,);
DFFARX1 I_74439 (I1267986,I2507,I1267502,I1267485,);
not I_74440 (I1268008,I1267986);
nand I_74441 (I1267482,I1268008,I1267536);
nand I_74442 (I1267476,I1268008,I1267638);
not I_74443 (I1268080,I2514);
DFFARX1 I_74444 (I1094802,I2507,I1268080,I1268106,);
nand I_74445 (I1268114,I1268106,I1094787);
not I_74446 (I1268131,I1268114);
DFFARX1 I_74447 (I1094790,I2507,I1268080,I1268157,);
not I_74448 (I1268165,I1268157);
not I_74449 (I1268182,I1094805);
or I_74450 (I1268199,I1094808,I1094805);
nor I_74451 (I1268216,I1094808,I1094805);
or I_74452 (I1268233,I1094784,I1094808);
DFFARX1 I_74453 (I1268233,I2507,I1268080,I1268072,);
not I_74454 (I1268264,I1094796);
nand I_74455 (I1268281,I1268264,I1094799);
nand I_74456 (I1268298,I1268182,I1268281);
and I_74457 (I1268051,I1268165,I1268298);
nor I_74458 (I1268329,I1094796,I1094793);
and I_74459 (I1268346,I1268165,I1268329);
nor I_74460 (I1268057,I1268131,I1268346);
DFFARX1 I_74461 (I1268329,I2507,I1268080,I1268386,);
not I_74462 (I1268394,I1268386);
nor I_74463 (I1268066,I1268165,I1268394);
or I_74464 (I1268425,I1268233,I1094784);
nor I_74465 (I1268442,I1094784,I1094784);
nand I_74466 (I1268459,I1268298,I1268442);
nand I_74467 (I1268476,I1268425,I1268459);
DFFARX1 I_74468 (I1268476,I2507,I1268080,I1268069,);
nor I_74469 (I1268507,I1268442,I1268199);
DFFARX1 I_74470 (I1268507,I2507,I1268080,I1268048,);
nor I_74471 (I1268538,I1094784,I1094787);
DFFARX1 I_74472 (I1268538,I2507,I1268080,I1268564,);
DFFARX1 I_74473 (I1268564,I2507,I1268080,I1268063,);
not I_74474 (I1268586,I1268564);
nand I_74475 (I1268060,I1268586,I1268114);
nand I_74476 (I1268054,I1268586,I1268216);
not I_74477 (I1268658,I2514);
DFFARX1 I_74478 (I1084976,I2507,I1268658,I1268684,);
nand I_74479 (I1268692,I1268684,I1084961);
not I_74480 (I1268709,I1268692);
DFFARX1 I_74481 (I1084964,I2507,I1268658,I1268735,);
not I_74482 (I1268743,I1268735);
not I_74483 (I1268760,I1084979);
or I_74484 (I1268777,I1084982,I1084979);
nor I_74485 (I1268794,I1084982,I1084979);
or I_74486 (I1268811,I1084958,I1084982);
DFFARX1 I_74487 (I1268811,I2507,I1268658,I1268650,);
not I_74488 (I1268842,I1084970);
nand I_74489 (I1268859,I1268842,I1084973);
nand I_74490 (I1268876,I1268760,I1268859);
and I_74491 (I1268629,I1268743,I1268876);
nor I_74492 (I1268907,I1084970,I1084967);
and I_74493 (I1268924,I1268743,I1268907);
nor I_74494 (I1268635,I1268709,I1268924);
DFFARX1 I_74495 (I1268907,I2507,I1268658,I1268964,);
not I_74496 (I1268972,I1268964);
nor I_74497 (I1268644,I1268743,I1268972);
or I_74498 (I1269003,I1268811,I1084958);
nor I_74499 (I1269020,I1084958,I1084958);
nand I_74500 (I1269037,I1268876,I1269020);
nand I_74501 (I1269054,I1269003,I1269037);
DFFARX1 I_74502 (I1269054,I2507,I1268658,I1268647,);
nor I_74503 (I1269085,I1269020,I1268777);
DFFARX1 I_74504 (I1269085,I2507,I1268658,I1268626,);
nor I_74505 (I1269116,I1084958,I1084961);
DFFARX1 I_74506 (I1269116,I2507,I1268658,I1269142,);
DFFARX1 I_74507 (I1269142,I2507,I1268658,I1268641,);
not I_74508 (I1269164,I1269142);
nand I_74509 (I1268638,I1269164,I1268692);
nand I_74510 (I1268632,I1269164,I1268794);
not I_74511 (I1269236,I2514);
DFFARX1 I_74512 (I865491,I2507,I1269236,I1269262,);
nand I_74513 (I1269270,I1269262,I865491);
not I_74514 (I1269287,I1269270);
DFFARX1 I_74515 (I865497,I2507,I1269236,I1269313,);
not I_74516 (I1269321,I1269313);
not I_74517 (I1269338,I865509);
or I_74518 (I1269355,I865494,I865509);
nor I_74519 (I1269372,I865494,I865509);
or I_74520 (I1269389,I865488,I865494);
DFFARX1 I_74521 (I1269389,I2507,I1269236,I1269228,);
not I_74522 (I1269420,I865506);
nand I_74523 (I1269437,I1269420,I865500);
nand I_74524 (I1269454,I1269338,I1269437);
and I_74525 (I1269207,I1269321,I1269454);
nor I_74526 (I1269485,I865506,I865488);
and I_74527 (I1269502,I1269321,I1269485);
nor I_74528 (I1269213,I1269287,I1269502);
DFFARX1 I_74529 (I1269485,I2507,I1269236,I1269542,);
not I_74530 (I1269550,I1269542);
nor I_74531 (I1269222,I1269321,I1269550);
or I_74532 (I1269581,I1269389,I865503);
nor I_74533 (I1269598,I865503,I865488);
nand I_74534 (I1269615,I1269454,I1269598);
nand I_74535 (I1269632,I1269581,I1269615);
DFFARX1 I_74536 (I1269632,I2507,I1269236,I1269225,);
nor I_74537 (I1269663,I1269598,I1269355);
DFFARX1 I_74538 (I1269663,I2507,I1269236,I1269204,);
nor I_74539 (I1269694,I865503,I865494);
DFFARX1 I_74540 (I1269694,I2507,I1269236,I1269720,);
DFFARX1 I_74541 (I1269720,I2507,I1269236,I1269219,);
not I_74542 (I1269742,I1269720);
nand I_74543 (I1269216,I1269742,I1269270);
nand I_74544 (I1269210,I1269742,I1269372);
not I_74545 (I1269814,I2514);
DFFARX1 I_74546 (I1972,I2507,I1269814,I1269840,);
nand I_74547 (I1269848,I1269840,I1788);
not I_74548 (I1269865,I1269848);
DFFARX1 I_74549 (I2012,I2507,I1269814,I1269891,);
not I_74550 (I1269899,I1269891);
not I_74551 (I1269916,I2292);
or I_74552 (I1269933,I1836,I2292);
nor I_74553 (I1269950,I1836,I2292);
or I_74554 (I1269967,I1804,I1836);
DFFARX1 I_74555 (I1269967,I2507,I1269814,I1269806,);
not I_74556 (I1269998,I1420);
nand I_74557 (I1270015,I1269998,I2084);
nand I_74558 (I1270032,I1269916,I1270015);
and I_74559 (I1269785,I1269899,I1270032);
nor I_74560 (I1270063,I1420,I2164);
and I_74561 (I1270080,I1269899,I1270063);
nor I_74562 (I1269791,I1269865,I1270080);
DFFARX1 I_74563 (I1270063,I2507,I1269814,I1270120,);
not I_74564 (I1270128,I1270120);
nor I_74565 (I1269800,I1269899,I1270128);
or I_74566 (I1270159,I1269967,I2356);
nor I_74567 (I1270176,I2356,I1804);
nand I_74568 (I1270193,I1270032,I1270176);
nand I_74569 (I1270210,I1270159,I1270193);
DFFARX1 I_74570 (I1270210,I2507,I1269814,I1269803,);
nor I_74571 (I1270241,I1270176,I1269933);
DFFARX1 I_74572 (I1270241,I2507,I1269814,I1269782,);
nor I_74573 (I1270272,I2356,I1964);
DFFARX1 I_74574 (I1270272,I2507,I1269814,I1270298,);
DFFARX1 I_74575 (I1270298,I2507,I1269814,I1269797,);
not I_74576 (I1270320,I1270298);
nand I_74577 (I1269794,I1270320,I1269848);
nand I_74578 (I1269788,I1270320,I1269950);
not I_74579 (I1270392,I2514);
DFFARX1 I_74580 (I969619,I2507,I1270392,I1270418,);
nand I_74581 (I1270426,I1270418,I969640);
not I_74582 (I1270443,I1270426);
DFFARX1 I_74583 (I969613,I2507,I1270392,I1270469,);
not I_74584 (I1270477,I1270469);
not I_74585 (I1270494,I969634);
or I_74586 (I1270511,I969625,I969634);
nor I_74587 (I1270528,I969625,I969634);
or I_74588 (I1270545,I969628,I969625);
DFFARX1 I_74589 (I1270545,I2507,I1270392,I1270384,);
not I_74590 (I1270576,I969616);
nand I_74591 (I1270593,I1270576,I969631);
nand I_74592 (I1270610,I1270494,I1270593);
and I_74593 (I1270363,I1270477,I1270610);
nor I_74594 (I1270641,I969616,I969613);
and I_74595 (I1270658,I1270477,I1270641);
nor I_74596 (I1270369,I1270443,I1270658);
DFFARX1 I_74597 (I1270641,I2507,I1270392,I1270698,);
not I_74598 (I1270706,I1270698);
nor I_74599 (I1270378,I1270477,I1270706);
or I_74600 (I1270737,I1270545,I969637);
nor I_74601 (I1270754,I969637,I969628);
nand I_74602 (I1270771,I1270610,I1270754);
nand I_74603 (I1270788,I1270737,I1270771);
DFFARX1 I_74604 (I1270788,I2507,I1270392,I1270381,);
nor I_74605 (I1270819,I1270754,I1270511);
DFFARX1 I_74606 (I1270819,I2507,I1270392,I1270360,);
nor I_74607 (I1270850,I969637,I969622);
DFFARX1 I_74608 (I1270850,I2507,I1270392,I1270876,);
DFFARX1 I_74609 (I1270876,I2507,I1270392,I1270375,);
not I_74610 (I1270898,I1270876);
nand I_74611 (I1270372,I1270898,I1270426);
nand I_74612 (I1270366,I1270898,I1270528);
not I_74613 (I1270970,I2514);
DFFARX1 I_74614 (I1239537,I2507,I1270970,I1270996,);
nand I_74615 (I1271004,I1270996,I1239546);
not I_74616 (I1271021,I1271004);
DFFARX1 I_74617 (I1239522,I2507,I1270970,I1271047,);
not I_74618 (I1271055,I1271047);
not I_74619 (I1271072,I1239525);
or I_74620 (I1271089,I1239522,I1239525);
nor I_74621 (I1271106,I1239522,I1239525);
or I_74622 (I1271123,I1239540,I1239522);
DFFARX1 I_74623 (I1271123,I2507,I1270970,I1270962,);
not I_74624 (I1271154,I1239528);
nand I_74625 (I1271171,I1271154,I1239543);
nand I_74626 (I1271188,I1271072,I1271171);
and I_74627 (I1270941,I1271055,I1271188);
nor I_74628 (I1271219,I1239528,I1239531);
and I_74629 (I1271236,I1271055,I1271219);
nor I_74630 (I1270947,I1271021,I1271236);
DFFARX1 I_74631 (I1271219,I2507,I1270970,I1271276,);
not I_74632 (I1271284,I1271276);
nor I_74633 (I1270956,I1271055,I1271284);
or I_74634 (I1271315,I1271123,I1239534);
nor I_74635 (I1271332,I1239534,I1239540);
nand I_74636 (I1271349,I1271188,I1271332);
nand I_74637 (I1271366,I1271315,I1271349);
DFFARX1 I_74638 (I1271366,I2507,I1270970,I1270959,);
nor I_74639 (I1271397,I1271332,I1271089);
DFFARX1 I_74640 (I1271397,I2507,I1270970,I1270938,);
nor I_74641 (I1271428,I1239534,I1239525);
DFFARX1 I_74642 (I1271428,I2507,I1270970,I1271454,);
DFFARX1 I_74643 (I1271454,I2507,I1270970,I1270953,);
not I_74644 (I1271476,I1271454);
nand I_74645 (I1270950,I1271476,I1271004);
nand I_74646 (I1270944,I1271476,I1271106);
not I_74647 (I1271548,I2514);
DFFARX1 I_74648 (I650370,I2507,I1271548,I1271574,);
nand I_74649 (I1271582,I1271574,I650373);
not I_74650 (I1271599,I1271582);
DFFARX1 I_74651 (I650385,I2507,I1271548,I1271625,);
not I_74652 (I1271633,I1271625);
not I_74653 (I1271650,I650370);
or I_74654 (I1271667,I650379,I650370);
nor I_74655 (I1271684,I650379,I650370);
or I_74656 (I1271701,I650388,I650379);
DFFARX1 I_74657 (I1271701,I2507,I1271548,I1271540,);
not I_74658 (I1271732,I650391);
nand I_74659 (I1271749,I1271732,I650373);
nand I_74660 (I1271766,I1271650,I1271749);
and I_74661 (I1271519,I1271633,I1271766);
nor I_74662 (I1271797,I650391,I650376);
and I_74663 (I1271814,I1271633,I1271797);
nor I_74664 (I1271525,I1271599,I1271814);
DFFARX1 I_74665 (I1271797,I2507,I1271548,I1271854,);
not I_74666 (I1271862,I1271854);
nor I_74667 (I1271534,I1271633,I1271862);
or I_74668 (I1271893,I1271701,I650382);
nor I_74669 (I1271910,I650382,I650388);
nand I_74670 (I1271927,I1271766,I1271910);
nand I_74671 (I1271944,I1271893,I1271927);
DFFARX1 I_74672 (I1271944,I2507,I1271548,I1271537,);
nor I_74673 (I1271975,I1271910,I1271667);
DFFARX1 I_74674 (I1271975,I2507,I1271548,I1271516,);
nor I_74675 (I1272006,I650382,I650394);
DFFARX1 I_74676 (I1272006,I2507,I1271548,I1272032,);
DFFARX1 I_74677 (I1272032,I2507,I1271548,I1271531,);
not I_74678 (I1272054,I1272032);
nand I_74679 (I1271528,I1272054,I1271582);
nand I_74680 (I1271522,I1272054,I1271684);
not I_74681 (I1272126,I2514);
DFFARX1 I_74682 (I1317831,I2507,I1272126,I1272152,);
nand I_74683 (I1272160,I1272152,I1317822);
not I_74684 (I1272177,I1272160);
DFFARX1 I_74685 (I1317807,I2507,I1272126,I1272203,);
not I_74686 (I1272211,I1272203);
not I_74687 (I1272228,I1317810);
or I_74688 (I1272245,I1317819,I1317810);
nor I_74689 (I1272262,I1317819,I1317810);
or I_74690 (I1272279,I1317816,I1317819);
DFFARX1 I_74691 (I1272279,I2507,I1272126,I1272118,);
not I_74692 (I1272310,I1317828);
nand I_74693 (I1272327,I1272310,I1317807);
nand I_74694 (I1272344,I1272228,I1272327);
and I_74695 (I1272097,I1272211,I1272344);
nor I_74696 (I1272375,I1317828,I1317813);
and I_74697 (I1272392,I1272211,I1272375);
nor I_74698 (I1272103,I1272177,I1272392);
DFFARX1 I_74699 (I1272375,I2507,I1272126,I1272432,);
not I_74700 (I1272440,I1272432);
nor I_74701 (I1272112,I1272211,I1272440);
or I_74702 (I1272471,I1272279,I1317834);
nor I_74703 (I1272488,I1317834,I1317816);
nand I_74704 (I1272505,I1272344,I1272488);
nand I_74705 (I1272522,I1272471,I1272505);
DFFARX1 I_74706 (I1272522,I2507,I1272126,I1272115,);
nor I_74707 (I1272553,I1272488,I1272245);
DFFARX1 I_74708 (I1272553,I2507,I1272126,I1272094,);
nor I_74709 (I1272584,I1317834,I1317825);
DFFARX1 I_74710 (I1272584,I2507,I1272126,I1272610,);
DFFARX1 I_74711 (I1272610,I2507,I1272126,I1272109,);
not I_74712 (I1272632,I1272610);
nand I_74713 (I1272106,I1272632,I1272160);
nand I_74714 (I1272100,I1272632,I1272262);
not I_74715 (I1272704,I2514);
DFFARX1 I_74716 (I748630,I2507,I1272704,I1272730,);
nand I_74717 (I1272738,I1272730,I748633);
not I_74718 (I1272755,I1272738);
DFFARX1 I_74719 (I748645,I2507,I1272704,I1272781,);
not I_74720 (I1272789,I1272781);
not I_74721 (I1272806,I748630);
or I_74722 (I1272823,I748639,I748630);
nor I_74723 (I1272840,I748639,I748630);
or I_74724 (I1272857,I748648,I748639);
DFFARX1 I_74725 (I1272857,I2507,I1272704,I1272696,);
not I_74726 (I1272888,I748651);
nand I_74727 (I1272905,I1272888,I748633);
nand I_74728 (I1272922,I1272806,I1272905);
and I_74729 (I1272675,I1272789,I1272922);
nor I_74730 (I1272953,I748651,I748636);
and I_74731 (I1272970,I1272789,I1272953);
nor I_74732 (I1272681,I1272755,I1272970);
DFFARX1 I_74733 (I1272953,I2507,I1272704,I1273010,);
not I_74734 (I1273018,I1273010);
nor I_74735 (I1272690,I1272789,I1273018);
or I_74736 (I1273049,I1272857,I748642);
nor I_74737 (I1273066,I748642,I748648);
nand I_74738 (I1273083,I1272922,I1273066);
nand I_74739 (I1273100,I1273049,I1273083);
DFFARX1 I_74740 (I1273100,I2507,I1272704,I1272693,);
nor I_74741 (I1273131,I1273066,I1272823);
DFFARX1 I_74742 (I1273131,I2507,I1272704,I1272672,);
nor I_74743 (I1273162,I748642,I748654);
DFFARX1 I_74744 (I1273162,I2507,I1272704,I1273188,);
DFFARX1 I_74745 (I1273188,I2507,I1272704,I1272687,);
not I_74746 (I1273210,I1273188);
nand I_74747 (I1272684,I1273210,I1272738);
nand I_74748 (I1272678,I1273210,I1272840);
not I_74749 (I1273282,I2514);
DFFARX1 I_74750 (I62250,I2507,I1273282,I1273308,);
nand I_74751 (I1273316,I1273308,I62241);
not I_74752 (I1273333,I1273316);
DFFARX1 I_74753 (I62238,I2507,I1273282,I1273359,);
not I_74754 (I1273367,I1273359);
not I_74755 (I1273384,I62247);
or I_74756 (I1273401,I62238,I62247);
nor I_74757 (I1273418,I62238,I62247);
or I_74758 (I1273435,I62244,I62238);
DFFARX1 I_74759 (I1273435,I2507,I1273282,I1273274,);
not I_74760 (I1273466,I62253);
nand I_74761 (I1273483,I1273466,I62262);
nand I_74762 (I1273500,I1273384,I1273483);
and I_74763 (I1273253,I1273367,I1273500);
nor I_74764 (I1273531,I62253,I62256);
and I_74765 (I1273548,I1273367,I1273531);
nor I_74766 (I1273259,I1273333,I1273548);
DFFARX1 I_74767 (I1273531,I2507,I1273282,I1273588,);
not I_74768 (I1273596,I1273588);
nor I_74769 (I1273268,I1273367,I1273596);
or I_74770 (I1273627,I1273435,I62241);
nor I_74771 (I1273644,I62241,I62244);
nand I_74772 (I1273661,I1273500,I1273644);
nand I_74773 (I1273678,I1273627,I1273661);
DFFARX1 I_74774 (I1273678,I2507,I1273282,I1273271,);
nor I_74775 (I1273709,I1273644,I1273401);
DFFARX1 I_74776 (I1273709,I2507,I1273282,I1273250,);
nor I_74777 (I1273740,I62241,I62259);
DFFARX1 I_74778 (I1273740,I2507,I1273282,I1273766,);
DFFARX1 I_74779 (I1273766,I2507,I1273282,I1273265,);
not I_74780 (I1273788,I1273766);
nand I_74781 (I1273262,I1273788,I1273316);
nand I_74782 (I1273256,I1273788,I1273418);
not I_74783 (I1273860,I2514);
DFFARX1 I_74784 (I546911,I2507,I1273860,I1273886,);
nand I_74785 (I1273894,I1273886,I546926);
not I_74786 (I1273911,I1273894);
DFFARX1 I_74787 (I546908,I2507,I1273860,I1273937,);
not I_74788 (I1273945,I1273937);
not I_74789 (I1273962,I546917);
or I_74790 (I1273979,I546911,I546917);
nor I_74791 (I1273996,I546911,I546917);
or I_74792 (I1274013,I546908,I546911);
DFFARX1 I_74793 (I1274013,I2507,I1273860,I1273852,);
not I_74794 (I1274044,I546929);
nand I_74795 (I1274061,I1274044,I546932);
nand I_74796 (I1274078,I1273962,I1274061);
and I_74797 (I1273831,I1273945,I1274078);
nor I_74798 (I1274109,I546929,I546914);
and I_74799 (I1274126,I1273945,I1274109);
nor I_74800 (I1273837,I1273911,I1274126);
DFFARX1 I_74801 (I1274109,I2507,I1273860,I1274166,);
not I_74802 (I1274174,I1274166);
nor I_74803 (I1273846,I1273945,I1274174);
or I_74804 (I1274205,I1274013,I546920);
nor I_74805 (I1274222,I546920,I546908);
nand I_74806 (I1274239,I1274078,I1274222);
nand I_74807 (I1274256,I1274205,I1274239);
DFFARX1 I_74808 (I1274256,I2507,I1273860,I1273849,);
nor I_74809 (I1274287,I1274222,I1273979);
DFFARX1 I_74810 (I1274287,I2507,I1273860,I1273828,);
nor I_74811 (I1274318,I546920,I546923);
DFFARX1 I_74812 (I1274318,I2507,I1273860,I1274344,);
DFFARX1 I_74813 (I1274344,I2507,I1273860,I1273843,);
not I_74814 (I1274366,I1274344);
nand I_74815 (I1273840,I1274366,I1273894);
nand I_74816 (I1273834,I1274366,I1273996);
not I_74817 (I1274438,I2514);
DFFARX1 I_74818 (I1134106,I2507,I1274438,I1274464,);
nand I_74819 (I1274472,I1274464,I1134091);
not I_74820 (I1274489,I1274472);
DFFARX1 I_74821 (I1134094,I2507,I1274438,I1274515,);
not I_74822 (I1274523,I1274515);
not I_74823 (I1274540,I1134109);
or I_74824 (I1274557,I1134112,I1134109);
nor I_74825 (I1274574,I1134112,I1134109);
or I_74826 (I1274591,I1134088,I1134112);
DFFARX1 I_74827 (I1274591,I2507,I1274438,I1274430,);
not I_74828 (I1274622,I1134100);
nand I_74829 (I1274639,I1274622,I1134103);
nand I_74830 (I1274656,I1274540,I1274639);
and I_74831 (I1274409,I1274523,I1274656);
nor I_74832 (I1274687,I1134100,I1134097);
and I_74833 (I1274704,I1274523,I1274687);
nor I_74834 (I1274415,I1274489,I1274704);
DFFARX1 I_74835 (I1274687,I2507,I1274438,I1274744,);
not I_74836 (I1274752,I1274744);
nor I_74837 (I1274424,I1274523,I1274752);
or I_74838 (I1274783,I1274591,I1134088);
nor I_74839 (I1274800,I1134088,I1134088);
nand I_74840 (I1274817,I1274656,I1274800);
nand I_74841 (I1274834,I1274783,I1274817);
DFFARX1 I_74842 (I1274834,I2507,I1274438,I1274427,);
nor I_74843 (I1274865,I1274800,I1274557);
DFFARX1 I_74844 (I1274865,I2507,I1274438,I1274406,);
nor I_74845 (I1274896,I1134088,I1134091);
DFFARX1 I_74846 (I1274896,I2507,I1274438,I1274922,);
DFFARX1 I_74847 (I1274922,I2507,I1274438,I1274421,);
not I_74848 (I1274944,I1274922);
nand I_74849 (I1274418,I1274944,I1274472);
nand I_74850 (I1274412,I1274944,I1274574);
not I_74851 (I1275016,I2514);
DFFARX1 I_74852 (I808575,I2507,I1275016,I1275042,);
nand I_74853 (I1275050,I1275042,I808575);
not I_74854 (I1275067,I1275050);
DFFARX1 I_74855 (I808581,I2507,I1275016,I1275093,);
not I_74856 (I1275101,I1275093);
not I_74857 (I1275118,I808593);
or I_74858 (I1275135,I808578,I808593);
nor I_74859 (I1275152,I808578,I808593);
or I_74860 (I1275169,I808572,I808578);
DFFARX1 I_74861 (I1275169,I2507,I1275016,I1275008,);
not I_74862 (I1275200,I808590);
nand I_74863 (I1275217,I1275200,I808584);
nand I_74864 (I1275234,I1275118,I1275217);
and I_74865 (I1274987,I1275101,I1275234);
nor I_74866 (I1275265,I808590,I808572);
and I_74867 (I1275282,I1275101,I1275265);
nor I_74868 (I1274993,I1275067,I1275282);
DFFARX1 I_74869 (I1275265,I2507,I1275016,I1275322,);
not I_74870 (I1275330,I1275322);
nor I_74871 (I1275002,I1275101,I1275330);
or I_74872 (I1275361,I1275169,I808587);
nor I_74873 (I1275378,I808587,I808572);
nand I_74874 (I1275395,I1275234,I1275378);
nand I_74875 (I1275412,I1275361,I1275395);
DFFARX1 I_74876 (I1275412,I2507,I1275016,I1275005,);
nor I_74877 (I1275443,I1275378,I1275135);
DFFARX1 I_74878 (I1275443,I2507,I1275016,I1274984,);
nor I_74879 (I1275474,I808587,I808578);
DFFARX1 I_74880 (I1275474,I2507,I1275016,I1275500,);
DFFARX1 I_74881 (I1275500,I2507,I1275016,I1274999,);
not I_74882 (I1275522,I1275500);
nand I_74883 (I1274996,I1275522,I1275050);
nand I_74884 (I1274990,I1275522,I1275152);
not I_74885 (I1275594,I2514);
DFFARX1 I_74886 (I424018,I2507,I1275594,I1275620,);
nand I_74887 (I1275628,I1275620,I424027);
not I_74888 (I1275645,I1275628);
DFFARX1 I_74889 (I424015,I2507,I1275594,I1275671,);
not I_74890 (I1275679,I1275671);
not I_74891 (I1275696,I424021);
or I_74892 (I1275713,I424015,I424021);
nor I_74893 (I1275730,I424015,I424021);
or I_74894 (I1275747,I424030,I424015);
DFFARX1 I_74895 (I1275747,I2507,I1275594,I1275586,);
not I_74896 (I1275778,I424024);
nand I_74897 (I1275795,I1275778,I424039);
nand I_74898 (I1275812,I1275696,I1275795);
and I_74899 (I1275565,I1275679,I1275812);
nor I_74900 (I1275843,I424024,I424042);
and I_74901 (I1275860,I1275679,I1275843);
nor I_74902 (I1275571,I1275645,I1275860);
DFFARX1 I_74903 (I1275843,I2507,I1275594,I1275900,);
not I_74904 (I1275908,I1275900);
nor I_74905 (I1275580,I1275679,I1275908);
or I_74906 (I1275939,I1275747,I424033);
nor I_74907 (I1275956,I424033,I424030);
nand I_74908 (I1275973,I1275812,I1275956);
nand I_74909 (I1275990,I1275939,I1275973);
DFFARX1 I_74910 (I1275990,I2507,I1275594,I1275583,);
nor I_74911 (I1276021,I1275956,I1275713);
DFFARX1 I_74912 (I1276021,I2507,I1275594,I1275562,);
nor I_74913 (I1276052,I424033,I424036);
DFFARX1 I_74914 (I1276052,I2507,I1275594,I1276078,);
DFFARX1 I_74915 (I1276078,I2507,I1275594,I1275577,);
not I_74916 (I1276100,I1276078);
nand I_74917 (I1275574,I1276100,I1275628);
nand I_74918 (I1275568,I1276100,I1275730);
not I_74919 (I1276172,I2514);
DFFARX1 I_74920 (I1009028,I2507,I1276172,I1276198,);
nand I_74921 (I1276206,I1276198,I1009025);
not I_74922 (I1276223,I1276206);
DFFARX1 I_74923 (I1009025,I2507,I1276172,I1276249,);
not I_74924 (I1276257,I1276249);
not I_74925 (I1276274,I1009022);
or I_74926 (I1276291,I1009031,I1009022);
nor I_74927 (I1276308,I1009031,I1009022);
or I_74928 (I1276325,I1009034,I1009031);
DFFARX1 I_74929 (I1276325,I2507,I1276172,I1276164,);
not I_74930 (I1276356,I1009022);
nand I_74931 (I1276373,I1276356,I1009019);
nand I_74932 (I1276390,I1276274,I1276373);
and I_74933 (I1276143,I1276257,I1276390);
nor I_74934 (I1276421,I1009022,I1009037);
and I_74935 (I1276438,I1276257,I1276421);
nor I_74936 (I1276149,I1276223,I1276438);
DFFARX1 I_74937 (I1276421,I2507,I1276172,I1276478,);
not I_74938 (I1276486,I1276478);
nor I_74939 (I1276158,I1276257,I1276486);
or I_74940 (I1276517,I1276325,I1009040);
nor I_74941 (I1276534,I1009040,I1009034);
nand I_74942 (I1276551,I1276390,I1276534);
nand I_74943 (I1276568,I1276517,I1276551);
DFFARX1 I_74944 (I1276568,I2507,I1276172,I1276161,);
nor I_74945 (I1276599,I1276534,I1276291);
DFFARX1 I_74946 (I1276599,I2507,I1276172,I1276140,);
nor I_74947 (I1276630,I1009040,I1009019);
DFFARX1 I_74948 (I1276630,I2507,I1276172,I1276656,);
DFFARX1 I_74949 (I1276656,I2507,I1276172,I1276155,);
not I_74950 (I1276678,I1276656);
nand I_74951 (I1276152,I1276678,I1276206);
nand I_74952 (I1276146,I1276678,I1276308);
not I_74953 (I1276750,I2514);
DFFARX1 I_74954 (I282870,I2507,I1276750,I1276776,);
nand I_74955 (I1276784,I1276776,I282891);
not I_74956 (I1276801,I1276784);
DFFARX1 I_74957 (I282885,I2507,I1276750,I1276827,);
not I_74958 (I1276835,I1276827);
not I_74959 (I1276852,I282873);
or I_74960 (I1276869,I282888,I282873);
nor I_74961 (I1276886,I282888,I282873);
or I_74962 (I1276903,I282879,I282888);
DFFARX1 I_74963 (I1276903,I2507,I1276750,I1276742,);
not I_74964 (I1276934,I282867);
nand I_74965 (I1276951,I1276934,I282864);
nand I_74966 (I1276968,I1276852,I1276951);
and I_74967 (I1276721,I1276835,I1276968);
nor I_74968 (I1276999,I282867,I282876);
and I_74969 (I1277016,I1276835,I1276999);
nor I_74970 (I1276727,I1276801,I1277016);
DFFARX1 I_74971 (I1276999,I2507,I1276750,I1277056,);
not I_74972 (I1277064,I1277056);
nor I_74973 (I1276736,I1276835,I1277064);
or I_74974 (I1277095,I1276903,I282882);
nor I_74975 (I1277112,I282882,I282879);
nand I_74976 (I1277129,I1276968,I1277112);
nand I_74977 (I1277146,I1277095,I1277129);
DFFARX1 I_74978 (I1277146,I2507,I1276750,I1276739,);
nor I_74979 (I1277177,I1277112,I1276869);
DFFARX1 I_74980 (I1277177,I2507,I1276750,I1276718,);
nor I_74981 (I1277208,I282882,I282864);
DFFARX1 I_74982 (I1277208,I2507,I1276750,I1277234,);
DFFARX1 I_74983 (I1277234,I2507,I1276750,I1276733,);
not I_74984 (I1277256,I1277234);
nand I_74985 (I1276730,I1277256,I1276784);
nand I_74986 (I1276724,I1277256,I1276886);
not I_74987 (I1277328,I2514);
DFFARX1 I_74988 (I390834,I2507,I1277328,I1277354,);
nand I_74989 (I1277362,I1277354,I390843);
not I_74990 (I1277379,I1277362);
DFFARX1 I_74991 (I390831,I2507,I1277328,I1277405,);
not I_74992 (I1277413,I1277405);
not I_74993 (I1277430,I390837);
or I_74994 (I1277447,I390831,I390837);
nor I_74995 (I1277464,I390831,I390837);
or I_74996 (I1277481,I390846,I390831);
DFFARX1 I_74997 (I1277481,I2507,I1277328,I1277320,);
not I_74998 (I1277512,I390840);
nand I_74999 (I1277529,I1277512,I390855);
nand I_75000 (I1277546,I1277430,I1277529);
and I_75001 (I1277299,I1277413,I1277546);
nor I_75002 (I1277577,I390840,I390858);
and I_75003 (I1277594,I1277413,I1277577);
nor I_75004 (I1277305,I1277379,I1277594);
DFFARX1 I_75005 (I1277577,I2507,I1277328,I1277634,);
not I_75006 (I1277642,I1277634);
nor I_75007 (I1277314,I1277413,I1277642);
or I_75008 (I1277673,I1277481,I390849);
nor I_75009 (I1277690,I390849,I390846);
nand I_75010 (I1277707,I1277546,I1277690);
nand I_75011 (I1277724,I1277673,I1277707);
DFFARX1 I_75012 (I1277724,I2507,I1277328,I1277317,);
nor I_75013 (I1277755,I1277690,I1277447);
DFFARX1 I_75014 (I1277755,I2507,I1277328,I1277296,);
nor I_75015 (I1277786,I390849,I390852);
DFFARX1 I_75016 (I1277786,I2507,I1277328,I1277812,);
DFFARX1 I_75017 (I1277812,I2507,I1277328,I1277311,);
not I_75018 (I1277834,I1277812);
nand I_75019 (I1277308,I1277834,I1277362);
nand I_75020 (I1277302,I1277834,I1277464);
not I_75021 (I1277906,I2514);
DFFARX1 I_75022 (I532764,I2507,I1277906,I1277932,);
nand I_75023 (I1277940,I1277932,I532773);
not I_75024 (I1277957,I1277940);
DFFARX1 I_75025 (I532785,I2507,I1277906,I1277983,);
not I_75026 (I1277991,I1277983);
not I_75027 (I1278008,I532776);
or I_75028 (I1278025,I532770,I532776);
nor I_75029 (I1278042,I532770,I532776);
or I_75030 (I1278059,I532764,I532770);
DFFARX1 I_75031 (I1278059,I2507,I1277906,I1277898,);
not I_75032 (I1278090,I532767);
nand I_75033 (I1278107,I1278090,I532779);
nand I_75034 (I1278124,I1278008,I1278107);
and I_75035 (I1277877,I1277991,I1278124);
nor I_75036 (I1278155,I532767,I532788);
and I_75037 (I1278172,I1277991,I1278155);
nor I_75038 (I1277883,I1277957,I1278172);
DFFARX1 I_75039 (I1278155,I2507,I1277906,I1278212,);
not I_75040 (I1278220,I1278212);
nor I_75041 (I1277892,I1277991,I1278220);
or I_75042 (I1278251,I1278059,I532782);
nor I_75043 (I1278268,I532782,I532764);
nand I_75044 (I1278285,I1278124,I1278268);
nand I_75045 (I1278302,I1278251,I1278285);
DFFARX1 I_75046 (I1278302,I2507,I1277906,I1277895,);
nor I_75047 (I1278333,I1278268,I1278025);
DFFARX1 I_75048 (I1278333,I2507,I1277906,I1277874,);
nor I_75049 (I1278364,I532782,I532767);
DFFARX1 I_75050 (I1278364,I2507,I1277906,I1278390,);
DFFARX1 I_75051 (I1278390,I2507,I1277906,I1277889,);
not I_75052 (I1278412,I1278390);
nand I_75053 (I1277886,I1278412,I1277940);
nand I_75054 (I1277880,I1278412,I1278042);
not I_75055 (I1278484,I2514);
DFFARX1 I_75056 (I754410,I2507,I1278484,I1278510,);
nand I_75057 (I1278518,I1278510,I754413);
not I_75058 (I1278535,I1278518);
DFFARX1 I_75059 (I754425,I2507,I1278484,I1278561,);
not I_75060 (I1278569,I1278561);
not I_75061 (I1278586,I754410);
or I_75062 (I1278603,I754419,I754410);
nor I_75063 (I1278620,I754419,I754410);
or I_75064 (I1278637,I754428,I754419);
DFFARX1 I_75065 (I1278637,I2507,I1278484,I1278476,);
not I_75066 (I1278668,I754431);
nand I_75067 (I1278685,I1278668,I754413);
nand I_75068 (I1278702,I1278586,I1278685);
and I_75069 (I1278455,I1278569,I1278702);
nor I_75070 (I1278733,I754431,I754416);
and I_75071 (I1278750,I1278569,I1278733);
nor I_75072 (I1278461,I1278535,I1278750);
DFFARX1 I_75073 (I1278733,I2507,I1278484,I1278790,);
not I_75074 (I1278798,I1278790);
nor I_75075 (I1278470,I1278569,I1278798);
or I_75076 (I1278829,I1278637,I754422);
nor I_75077 (I1278846,I754422,I754428);
nand I_75078 (I1278863,I1278702,I1278846);
nand I_75079 (I1278880,I1278829,I1278863);
DFFARX1 I_75080 (I1278880,I2507,I1278484,I1278473,);
nor I_75081 (I1278911,I1278846,I1278603);
DFFARX1 I_75082 (I1278911,I2507,I1278484,I1278452,);
nor I_75083 (I1278942,I754422,I754434);
DFFARX1 I_75084 (I1278942,I2507,I1278484,I1278968,);
DFFARX1 I_75085 (I1278968,I2507,I1278484,I1278467,);
not I_75086 (I1278990,I1278968);
nand I_75087 (I1278464,I1278990,I1278518);
nand I_75088 (I1278458,I1278990,I1278620);
not I_75089 (I1279062,I2514);
DFFARX1 I_75090 (I147865,I2507,I1279062,I1279088,);
nand I_75091 (I1279096,I1279088,I147874);
not I_75092 (I1279113,I1279096);
DFFARX1 I_75093 (I147856,I2507,I1279062,I1279139,);
not I_75094 (I1279147,I1279139);
not I_75095 (I1279164,I147862);
or I_75096 (I1279181,I147871,I147862);
nor I_75097 (I1279198,I147871,I147862);
or I_75098 (I1279215,I147859,I147871);
DFFARX1 I_75099 (I1279215,I2507,I1279062,I1279054,);
not I_75100 (I1279246,I147877);
nand I_75101 (I1279263,I1279246,I147850);
nand I_75102 (I1279280,I1279164,I1279263);
and I_75103 (I1279033,I1279147,I1279280);
nor I_75104 (I1279311,I147877,I147853);
and I_75105 (I1279328,I1279147,I1279311);
nor I_75106 (I1279039,I1279113,I1279328);
DFFARX1 I_75107 (I1279311,I2507,I1279062,I1279368,);
not I_75108 (I1279376,I1279368);
nor I_75109 (I1279048,I1279147,I1279376);
or I_75110 (I1279407,I1279215,I147868);
nor I_75111 (I1279424,I147868,I147859);
nand I_75112 (I1279441,I1279280,I1279424);
nand I_75113 (I1279458,I1279407,I1279441);
DFFARX1 I_75114 (I1279458,I2507,I1279062,I1279051,);
nor I_75115 (I1279489,I1279424,I1279181);
DFFARX1 I_75116 (I1279489,I2507,I1279062,I1279030,);
nor I_75117 (I1279520,I147868,I147850);
DFFARX1 I_75118 (I1279520,I2507,I1279062,I1279546,);
DFFARX1 I_75119 (I1279546,I2507,I1279062,I1279045,);
not I_75120 (I1279568,I1279546);
nand I_75121 (I1279042,I1279568,I1279096);
nand I_75122 (I1279036,I1279568,I1279198);
not I_75123 (I1279640,I2514);
DFFARX1 I_75124 (I505989,I2507,I1279640,I1279666,);
nand I_75125 (I1279674,I1279666,I505998);
not I_75126 (I1279691,I1279674);
DFFARX1 I_75127 (I506010,I2507,I1279640,I1279717,);
not I_75128 (I1279725,I1279717);
not I_75129 (I1279742,I506001);
or I_75130 (I1279759,I505995,I506001);
nor I_75131 (I1279776,I505995,I506001);
or I_75132 (I1279793,I505989,I505995);
DFFARX1 I_75133 (I1279793,I2507,I1279640,I1279632,);
not I_75134 (I1279824,I505992);
nand I_75135 (I1279841,I1279824,I506004);
nand I_75136 (I1279858,I1279742,I1279841);
and I_75137 (I1279611,I1279725,I1279858);
nor I_75138 (I1279889,I505992,I506013);
and I_75139 (I1279906,I1279725,I1279889);
nor I_75140 (I1279617,I1279691,I1279906);
DFFARX1 I_75141 (I1279889,I2507,I1279640,I1279946,);
not I_75142 (I1279954,I1279946);
nor I_75143 (I1279626,I1279725,I1279954);
or I_75144 (I1279985,I1279793,I506007);
nor I_75145 (I1280002,I506007,I505989);
nand I_75146 (I1280019,I1279858,I1280002);
nand I_75147 (I1280036,I1279985,I1280019);
DFFARX1 I_75148 (I1280036,I2507,I1279640,I1279629,);
nor I_75149 (I1280067,I1280002,I1279759);
DFFARX1 I_75150 (I1280067,I2507,I1279640,I1279608,);
nor I_75151 (I1280098,I506007,I505992);
DFFARX1 I_75152 (I1280098,I2507,I1279640,I1280124,);
DFFARX1 I_75153 (I1280124,I2507,I1279640,I1279623,);
not I_75154 (I1280146,I1280124);
nand I_75155 (I1279620,I1280146,I1279674);
nand I_75156 (I1279614,I1280146,I1279776);
not I_75157 (I1280218,I2514);
DFFARX1 I_75158 (I1328541,I2507,I1280218,I1280244,);
nand I_75159 (I1280252,I1280244,I1328532);
not I_75160 (I1280269,I1280252);
DFFARX1 I_75161 (I1328517,I2507,I1280218,I1280295,);
not I_75162 (I1280303,I1280295);
not I_75163 (I1280320,I1328520);
or I_75164 (I1280337,I1328529,I1328520);
nor I_75165 (I1280354,I1328529,I1328520);
or I_75166 (I1280371,I1328526,I1328529);
DFFARX1 I_75167 (I1280371,I2507,I1280218,I1280210,);
not I_75168 (I1280402,I1328538);
nand I_75169 (I1280419,I1280402,I1328517);
nand I_75170 (I1280436,I1280320,I1280419);
and I_75171 (I1280189,I1280303,I1280436);
nor I_75172 (I1280467,I1328538,I1328523);
and I_75173 (I1280484,I1280303,I1280467);
nor I_75174 (I1280195,I1280269,I1280484);
DFFARX1 I_75175 (I1280467,I2507,I1280218,I1280524,);
not I_75176 (I1280532,I1280524);
nor I_75177 (I1280204,I1280303,I1280532);
or I_75178 (I1280563,I1280371,I1328544);
nor I_75179 (I1280580,I1328544,I1328526);
nand I_75180 (I1280597,I1280436,I1280580);
nand I_75181 (I1280614,I1280563,I1280597);
DFFARX1 I_75182 (I1280614,I2507,I1280218,I1280207,);
nor I_75183 (I1280645,I1280580,I1280337);
DFFARX1 I_75184 (I1280645,I2507,I1280218,I1280186,);
nor I_75185 (I1280676,I1328544,I1328535);
DFFARX1 I_75186 (I1280676,I2507,I1280218,I1280702,);
DFFARX1 I_75187 (I1280702,I2507,I1280218,I1280201,);
not I_75188 (I1280724,I1280702);
nand I_75189 (I1280198,I1280724,I1280252);
nand I_75190 (I1280192,I1280724,I1280354);
not I_75191 (I1280796,I2514);
DFFARX1 I_75192 (I282343,I2507,I1280796,I1280822,);
nand I_75193 (I1280830,I1280822,I282364);
not I_75194 (I1280847,I1280830);
DFFARX1 I_75195 (I282358,I2507,I1280796,I1280873,);
not I_75196 (I1280881,I1280873);
not I_75197 (I1280898,I282346);
or I_75198 (I1280915,I282361,I282346);
nor I_75199 (I1280932,I282361,I282346);
or I_75200 (I1280949,I282352,I282361);
DFFARX1 I_75201 (I1280949,I2507,I1280796,I1280788,);
not I_75202 (I1280980,I282340);
nand I_75203 (I1280997,I1280980,I282337);
nand I_75204 (I1281014,I1280898,I1280997);
and I_75205 (I1280767,I1280881,I1281014);
nor I_75206 (I1281045,I282340,I282349);
and I_75207 (I1281062,I1280881,I1281045);
nor I_75208 (I1280773,I1280847,I1281062);
DFFARX1 I_75209 (I1281045,I2507,I1280796,I1281102,);
not I_75210 (I1281110,I1281102);
nor I_75211 (I1280782,I1280881,I1281110);
or I_75212 (I1281141,I1280949,I282355);
nor I_75213 (I1281158,I282355,I282352);
nand I_75214 (I1281175,I1281014,I1281158);
nand I_75215 (I1281192,I1281141,I1281175);
DFFARX1 I_75216 (I1281192,I2507,I1280796,I1280785,);
nor I_75217 (I1281223,I1281158,I1280915);
DFFARX1 I_75218 (I1281223,I2507,I1280796,I1280764,);
nor I_75219 (I1281254,I282355,I282337);
DFFARX1 I_75220 (I1281254,I2507,I1280796,I1281280,);
DFFARX1 I_75221 (I1281280,I2507,I1280796,I1280779,);
not I_75222 (I1281302,I1281280);
nand I_75223 (I1280776,I1281302,I1280830);
nand I_75224 (I1280770,I1281302,I1280932);
not I_75225 (I1281374,I2514);
DFFARX1 I_75226 (I1161272,I2507,I1281374,I1281400,);
nand I_75227 (I1281408,I1281400,I1161257);
not I_75228 (I1281425,I1281408);
DFFARX1 I_75229 (I1161260,I2507,I1281374,I1281451,);
not I_75230 (I1281459,I1281451);
not I_75231 (I1281476,I1161275);
or I_75232 (I1281493,I1161278,I1161275);
nor I_75233 (I1281510,I1161278,I1161275);
or I_75234 (I1281527,I1161254,I1161278);
DFFARX1 I_75235 (I1281527,I2507,I1281374,I1281366,);
not I_75236 (I1281558,I1161266);
nand I_75237 (I1281575,I1281558,I1161269);
nand I_75238 (I1281592,I1281476,I1281575);
and I_75239 (I1281345,I1281459,I1281592);
nor I_75240 (I1281623,I1161266,I1161263);
and I_75241 (I1281640,I1281459,I1281623);
nor I_75242 (I1281351,I1281425,I1281640);
DFFARX1 I_75243 (I1281623,I2507,I1281374,I1281680,);
not I_75244 (I1281688,I1281680);
nor I_75245 (I1281360,I1281459,I1281688);
or I_75246 (I1281719,I1281527,I1161254);
nor I_75247 (I1281736,I1161254,I1161254);
nand I_75248 (I1281753,I1281592,I1281736);
nand I_75249 (I1281770,I1281719,I1281753);
DFFARX1 I_75250 (I1281770,I2507,I1281374,I1281363,);
nor I_75251 (I1281801,I1281736,I1281493);
DFFARX1 I_75252 (I1281801,I2507,I1281374,I1281342,);
nor I_75253 (I1281832,I1161254,I1161257);
DFFARX1 I_75254 (I1281832,I2507,I1281374,I1281858,);
DFFARX1 I_75255 (I1281858,I2507,I1281374,I1281357,);
not I_75256 (I1281880,I1281858);
nand I_75257 (I1281354,I1281880,I1281408);
nand I_75258 (I1281348,I1281880,I1281510);
not I_75259 (I1281952,I2514);
DFFARX1 I_75260 (I221630,I2507,I1281952,I1281978,);
nand I_75261 (I1281986,I1281978,I221633);
not I_75262 (I1282003,I1281986);
DFFARX1 I_75263 (I221642,I2507,I1281952,I1282029,);
not I_75264 (I1282037,I1282029);
not I_75265 (I1282054,I221645);
or I_75266 (I1282071,I221636,I221645);
nor I_75267 (I1282088,I221636,I221645);
or I_75268 (I1282105,I221648,I221636);
DFFARX1 I_75269 (I1282105,I2507,I1281952,I1281944,);
not I_75270 (I1282136,I221633);
nand I_75271 (I1282153,I1282136,I221639);
nand I_75272 (I1282170,I1282054,I1282153);
and I_75273 (I1281923,I1282037,I1282170);
nor I_75274 (I1282201,I221633,I221651);
and I_75275 (I1282218,I1282037,I1282201);
nor I_75276 (I1281929,I1282003,I1282218);
DFFARX1 I_75277 (I1282201,I2507,I1281952,I1282258,);
not I_75278 (I1282266,I1282258);
nor I_75279 (I1281938,I1282037,I1282266);
or I_75280 (I1282297,I1282105,I221630);
nor I_75281 (I1282314,I221630,I221648);
nand I_75282 (I1282331,I1282170,I1282314);
nand I_75283 (I1282348,I1282297,I1282331);
DFFARX1 I_75284 (I1282348,I2507,I1281952,I1281941,);
nor I_75285 (I1282379,I1282314,I1282071);
DFFARX1 I_75286 (I1282379,I2507,I1281952,I1281920,);
nor I_75287 (I1282410,I221630,I221654);
DFFARX1 I_75288 (I1282410,I2507,I1281952,I1282436,);
DFFARX1 I_75289 (I1282436,I2507,I1281952,I1281935,);
not I_75290 (I1282458,I1282436);
nand I_75291 (I1281932,I1282458,I1281986);
nand I_75292 (I1281926,I1282458,I1282088);
not I_75293 (I1282530,I2514);
DFFARX1 I_75294 (I1103472,I2507,I1282530,I1282556,);
nand I_75295 (I1282564,I1282556,I1103457);
not I_75296 (I1282581,I1282564);
DFFARX1 I_75297 (I1103460,I2507,I1282530,I1282607,);
not I_75298 (I1282615,I1282607);
not I_75299 (I1282632,I1103475);
or I_75300 (I1282649,I1103478,I1103475);
nor I_75301 (I1282666,I1103478,I1103475);
or I_75302 (I1282683,I1103454,I1103478);
DFFARX1 I_75303 (I1282683,I2507,I1282530,I1282522,);
not I_75304 (I1282714,I1103466);
nand I_75305 (I1282731,I1282714,I1103469);
nand I_75306 (I1282748,I1282632,I1282731);
and I_75307 (I1282501,I1282615,I1282748);
nor I_75308 (I1282779,I1103466,I1103463);
and I_75309 (I1282796,I1282615,I1282779);
nor I_75310 (I1282507,I1282581,I1282796);
DFFARX1 I_75311 (I1282779,I2507,I1282530,I1282836,);
not I_75312 (I1282844,I1282836);
nor I_75313 (I1282516,I1282615,I1282844);
or I_75314 (I1282875,I1282683,I1103454);
nor I_75315 (I1282892,I1103454,I1103454);
nand I_75316 (I1282909,I1282748,I1282892);
nand I_75317 (I1282926,I1282875,I1282909);
DFFARX1 I_75318 (I1282926,I2507,I1282530,I1282519,);
nor I_75319 (I1282957,I1282892,I1282649);
DFFARX1 I_75320 (I1282957,I2507,I1282530,I1282498,);
nor I_75321 (I1282988,I1103454,I1103457);
DFFARX1 I_75322 (I1282988,I2507,I1282530,I1283014,);
DFFARX1 I_75323 (I1283014,I2507,I1282530,I1282513,);
not I_75324 (I1283036,I1283014);
nand I_75325 (I1282510,I1283036,I1282564);
nand I_75326 (I1282504,I1283036,I1282666);
not I_75327 (I1283108,I2514);
DFFARX1 I_75328 (I539309,I2507,I1283108,I1283134,);
nand I_75329 (I1283142,I1283134,I539318);
not I_75330 (I1283159,I1283142);
DFFARX1 I_75331 (I539330,I2507,I1283108,I1283185,);
not I_75332 (I1283193,I1283185);
not I_75333 (I1283210,I539321);
or I_75334 (I1283227,I539315,I539321);
nor I_75335 (I1283244,I539315,I539321);
or I_75336 (I1283261,I539309,I539315);
DFFARX1 I_75337 (I1283261,I2507,I1283108,I1283100,);
not I_75338 (I1283292,I539312);
nand I_75339 (I1283309,I1283292,I539324);
nand I_75340 (I1283326,I1283210,I1283309);
and I_75341 (I1283079,I1283193,I1283326);
nor I_75342 (I1283357,I539312,I539333);
and I_75343 (I1283374,I1283193,I1283357);
nor I_75344 (I1283085,I1283159,I1283374);
DFFARX1 I_75345 (I1283357,I2507,I1283108,I1283414,);
not I_75346 (I1283422,I1283414);
nor I_75347 (I1283094,I1283193,I1283422);
or I_75348 (I1283453,I1283261,I539327);
nor I_75349 (I1283470,I539327,I539309);
nand I_75350 (I1283487,I1283326,I1283470);
nand I_75351 (I1283504,I1283453,I1283487);
DFFARX1 I_75352 (I1283504,I2507,I1283108,I1283097,);
nor I_75353 (I1283535,I1283470,I1283227);
DFFARX1 I_75354 (I1283535,I2507,I1283108,I1283076,);
nor I_75355 (I1283566,I539327,I539312);
DFFARX1 I_75356 (I1283566,I2507,I1283108,I1283592,);
DFFARX1 I_75357 (I1283592,I2507,I1283108,I1283091,);
not I_75358 (I1283614,I1283592);
nand I_75359 (I1283088,I1283614,I1283142);
nand I_75360 (I1283082,I1283614,I1283244);
not I_75361 (I1283686,I2514);
DFFARX1 I_75362 (I1176300,I2507,I1283686,I1283712,);
nand I_75363 (I1283720,I1283712,I1176285);
not I_75364 (I1283737,I1283720);
DFFARX1 I_75365 (I1176288,I2507,I1283686,I1283763,);
not I_75366 (I1283771,I1283763);
not I_75367 (I1283788,I1176303);
or I_75368 (I1283805,I1176306,I1176303);
nor I_75369 (I1283822,I1176306,I1176303);
or I_75370 (I1283839,I1176282,I1176306);
DFFARX1 I_75371 (I1283839,I2507,I1283686,I1283678,);
not I_75372 (I1283870,I1176294);
nand I_75373 (I1283887,I1283870,I1176297);
nand I_75374 (I1283904,I1283788,I1283887);
and I_75375 (I1283657,I1283771,I1283904);
nor I_75376 (I1283935,I1176294,I1176291);
and I_75377 (I1283952,I1283771,I1283935);
nor I_75378 (I1283663,I1283737,I1283952);
DFFARX1 I_75379 (I1283935,I2507,I1283686,I1283992,);
not I_75380 (I1284000,I1283992);
nor I_75381 (I1283672,I1283771,I1284000);
or I_75382 (I1284031,I1283839,I1176282);
nor I_75383 (I1284048,I1176282,I1176282);
nand I_75384 (I1284065,I1283904,I1284048);
nand I_75385 (I1284082,I1284031,I1284065);
DFFARX1 I_75386 (I1284082,I2507,I1283686,I1283675,);
nor I_75387 (I1284113,I1284048,I1283805);
DFFARX1 I_75388 (I1284113,I2507,I1283686,I1283654,);
nor I_75389 (I1284144,I1176282,I1176285);
DFFARX1 I_75390 (I1284144,I2507,I1283686,I1284170,);
DFFARX1 I_75391 (I1284170,I2507,I1283686,I1283669,);
not I_75392 (I1284192,I1284170);
nand I_75393 (I1283666,I1284192,I1283720);
nand I_75394 (I1283660,I1284192,I1283822);
not I_75395 (I1284264,I2514);
DFFARX1 I_75396 (I1374356,I2507,I1284264,I1284290,);
nand I_75397 (I1284298,I1284290,I1374347);
not I_75398 (I1284315,I1284298);
DFFARX1 I_75399 (I1374332,I2507,I1284264,I1284341,);
not I_75400 (I1284349,I1284341);
not I_75401 (I1284366,I1374335);
or I_75402 (I1284383,I1374344,I1374335);
nor I_75403 (I1284400,I1374344,I1374335);
or I_75404 (I1284417,I1374341,I1374344);
DFFARX1 I_75405 (I1284417,I2507,I1284264,I1284256,);
not I_75406 (I1284448,I1374353);
nand I_75407 (I1284465,I1284448,I1374332);
nand I_75408 (I1284482,I1284366,I1284465);
and I_75409 (I1284235,I1284349,I1284482);
nor I_75410 (I1284513,I1374353,I1374338);
and I_75411 (I1284530,I1284349,I1284513);
nor I_75412 (I1284241,I1284315,I1284530);
DFFARX1 I_75413 (I1284513,I2507,I1284264,I1284570,);
not I_75414 (I1284578,I1284570);
nor I_75415 (I1284250,I1284349,I1284578);
or I_75416 (I1284609,I1284417,I1374359);
nor I_75417 (I1284626,I1374359,I1374341);
nand I_75418 (I1284643,I1284482,I1284626);
nand I_75419 (I1284660,I1284609,I1284643);
DFFARX1 I_75420 (I1284660,I2507,I1284264,I1284253,);
nor I_75421 (I1284691,I1284626,I1284383);
DFFARX1 I_75422 (I1284691,I2507,I1284264,I1284232,);
nor I_75423 (I1284722,I1374359,I1374350);
DFFARX1 I_75424 (I1284722,I2507,I1284264,I1284748,);
DFFARX1 I_75425 (I1284748,I2507,I1284264,I1284247,);
not I_75426 (I1284770,I1284748);
nand I_75427 (I1284244,I1284770,I1284298);
nand I_75428 (I1284238,I1284770,I1284400);
not I_75429 (I1284842,I2514);
DFFARX1 I_75430 (I532169,I2507,I1284842,I1284868,);
nand I_75431 (I1284876,I1284868,I532178);
not I_75432 (I1284893,I1284876);
DFFARX1 I_75433 (I532190,I2507,I1284842,I1284919,);
not I_75434 (I1284927,I1284919);
not I_75435 (I1284944,I532181);
or I_75436 (I1284961,I532175,I532181);
nor I_75437 (I1284978,I532175,I532181);
or I_75438 (I1284995,I532169,I532175);
DFFARX1 I_75439 (I1284995,I2507,I1284842,I1284834,);
not I_75440 (I1285026,I532172);
nand I_75441 (I1285043,I1285026,I532184);
nand I_75442 (I1285060,I1284944,I1285043);
and I_75443 (I1284813,I1284927,I1285060);
nor I_75444 (I1285091,I532172,I532193);
and I_75445 (I1285108,I1284927,I1285091);
nor I_75446 (I1284819,I1284893,I1285108);
DFFARX1 I_75447 (I1285091,I2507,I1284842,I1285148,);
not I_75448 (I1285156,I1285148);
nor I_75449 (I1284828,I1284927,I1285156);
or I_75450 (I1285187,I1284995,I532187);
nor I_75451 (I1285204,I532187,I532169);
nand I_75452 (I1285221,I1285060,I1285204);
nand I_75453 (I1285238,I1285187,I1285221);
DFFARX1 I_75454 (I1285238,I2507,I1284842,I1284831,);
nor I_75455 (I1285269,I1285204,I1284961);
DFFARX1 I_75456 (I1285269,I2507,I1284842,I1284810,);
nor I_75457 (I1285300,I532187,I532172);
DFFARX1 I_75458 (I1285300,I2507,I1284842,I1285326,);
DFFARX1 I_75459 (I1285326,I2507,I1284842,I1284825,);
not I_75460 (I1285348,I1285326);
nand I_75461 (I1284822,I1285348,I1284876);
nand I_75462 (I1284816,I1285348,I1284978);
not I_75463 (I1285420,I2514);
DFFARX1 I_75464 (I990291,I2507,I1285420,I1285446,);
nand I_75465 (I1285454,I1285446,I990312);
not I_75466 (I1285471,I1285454);
DFFARX1 I_75467 (I990285,I2507,I1285420,I1285497,);
not I_75468 (I1285505,I1285497);
not I_75469 (I1285522,I990306);
or I_75470 (I1285539,I990297,I990306);
nor I_75471 (I1285556,I990297,I990306);
or I_75472 (I1285573,I990300,I990297);
DFFARX1 I_75473 (I1285573,I2507,I1285420,I1285412,);
not I_75474 (I1285604,I990288);
nand I_75475 (I1285621,I1285604,I990303);
nand I_75476 (I1285638,I1285522,I1285621);
and I_75477 (I1285391,I1285505,I1285638);
nor I_75478 (I1285669,I990288,I990285);
and I_75479 (I1285686,I1285505,I1285669);
nor I_75480 (I1285397,I1285471,I1285686);
DFFARX1 I_75481 (I1285669,I2507,I1285420,I1285726,);
not I_75482 (I1285734,I1285726);
nor I_75483 (I1285406,I1285505,I1285734);
or I_75484 (I1285765,I1285573,I990309);
nor I_75485 (I1285782,I990309,I990300);
nand I_75486 (I1285799,I1285638,I1285782);
nand I_75487 (I1285816,I1285765,I1285799);
DFFARX1 I_75488 (I1285816,I2507,I1285420,I1285409,);
nor I_75489 (I1285847,I1285782,I1285539);
DFFARX1 I_75490 (I1285847,I2507,I1285420,I1285388,);
nor I_75491 (I1285878,I990309,I990294);
DFFARX1 I_75492 (I1285878,I2507,I1285420,I1285904,);
DFFARX1 I_75493 (I1285904,I2507,I1285420,I1285403,);
not I_75494 (I1285926,I1285904);
nand I_75495 (I1285400,I1285926,I1285454);
nand I_75496 (I1285394,I1285926,I1285556);
not I_75497 (I1285998,I2514);
DFFARX1 I_75498 (I1006441,I2507,I1285998,I1286024,);
nand I_75499 (I1286032,I1286024,I1006462);
not I_75500 (I1286049,I1286032);
DFFARX1 I_75501 (I1006435,I2507,I1285998,I1286075,);
not I_75502 (I1286083,I1286075);
not I_75503 (I1286100,I1006456);
or I_75504 (I1286117,I1006447,I1006456);
nor I_75505 (I1286134,I1006447,I1006456);
or I_75506 (I1286151,I1006450,I1006447);
DFFARX1 I_75507 (I1286151,I2507,I1285998,I1285990,);
not I_75508 (I1286182,I1006438);
nand I_75509 (I1286199,I1286182,I1006453);
nand I_75510 (I1286216,I1286100,I1286199);
and I_75511 (I1285969,I1286083,I1286216);
nor I_75512 (I1286247,I1006438,I1006435);
and I_75513 (I1286264,I1286083,I1286247);
nor I_75514 (I1285975,I1286049,I1286264);
DFFARX1 I_75515 (I1286247,I2507,I1285998,I1286304,);
not I_75516 (I1286312,I1286304);
nor I_75517 (I1285984,I1286083,I1286312);
or I_75518 (I1286343,I1286151,I1006459);
nor I_75519 (I1286360,I1006459,I1006450);
nand I_75520 (I1286377,I1286216,I1286360);
nand I_75521 (I1286394,I1286343,I1286377);
DFFARX1 I_75522 (I1286394,I2507,I1285998,I1285987,);
nor I_75523 (I1286425,I1286360,I1286117);
DFFARX1 I_75524 (I1286425,I2507,I1285998,I1285966,);
nor I_75525 (I1286456,I1006459,I1006444);
DFFARX1 I_75526 (I1286456,I2507,I1285998,I1286482,);
DFFARX1 I_75527 (I1286482,I2507,I1285998,I1285981,);
not I_75528 (I1286504,I1286482);
nand I_75529 (I1285978,I1286504,I1286032);
nand I_75530 (I1285972,I1286504,I1286134);
not I_75531 (I1286576,I2514);
DFFARX1 I_75532 (I1038200,I2507,I1286576,I1286602,);
nand I_75533 (I1286610,I1286602,I1038197);
not I_75534 (I1286627,I1286610);
DFFARX1 I_75535 (I1038197,I2507,I1286576,I1286653,);
not I_75536 (I1286661,I1286653);
not I_75537 (I1286678,I1038194);
or I_75538 (I1286695,I1038203,I1038194);
nor I_75539 (I1286712,I1038203,I1038194);
or I_75540 (I1286729,I1038206,I1038203);
DFFARX1 I_75541 (I1286729,I2507,I1286576,I1286568,);
not I_75542 (I1286760,I1038194);
nand I_75543 (I1286777,I1286760,I1038191);
nand I_75544 (I1286794,I1286678,I1286777);
and I_75545 (I1286547,I1286661,I1286794);
nor I_75546 (I1286825,I1038194,I1038209);
and I_75547 (I1286842,I1286661,I1286825);
nor I_75548 (I1286553,I1286627,I1286842);
DFFARX1 I_75549 (I1286825,I2507,I1286576,I1286882,);
not I_75550 (I1286890,I1286882);
nor I_75551 (I1286562,I1286661,I1286890);
or I_75552 (I1286921,I1286729,I1038212);
nor I_75553 (I1286938,I1038212,I1038206);
nand I_75554 (I1286955,I1286794,I1286938);
nand I_75555 (I1286972,I1286921,I1286955);
DFFARX1 I_75556 (I1286972,I2507,I1286576,I1286565,);
nor I_75557 (I1287003,I1286938,I1286695);
DFFARX1 I_75558 (I1287003,I2507,I1286576,I1286544,);
nor I_75559 (I1287034,I1038212,I1038191);
DFFARX1 I_75560 (I1287034,I2507,I1286576,I1287060,);
DFFARX1 I_75561 (I1287060,I2507,I1286576,I1286559,);
not I_75562 (I1287082,I1287060);
nand I_75563 (I1286556,I1287082,I1286610);
nand I_75564 (I1286550,I1287082,I1286712);
not I_75565 (I1287154,I2514);
DFFARX1 I_75566 (I529194,I2507,I1287154,I1287180,);
nand I_75567 (I1287188,I1287180,I529203);
not I_75568 (I1287205,I1287188);
DFFARX1 I_75569 (I529215,I2507,I1287154,I1287231,);
not I_75570 (I1287239,I1287231);
not I_75571 (I1287256,I529206);
or I_75572 (I1287273,I529200,I529206);
nor I_75573 (I1287290,I529200,I529206);
or I_75574 (I1287307,I529194,I529200);
DFFARX1 I_75575 (I1287307,I2507,I1287154,I1287146,);
not I_75576 (I1287338,I529197);
nand I_75577 (I1287355,I1287338,I529209);
nand I_75578 (I1287372,I1287256,I1287355);
and I_75579 (I1287125,I1287239,I1287372);
nor I_75580 (I1287403,I529197,I529218);
and I_75581 (I1287420,I1287239,I1287403);
nor I_75582 (I1287131,I1287205,I1287420);
DFFARX1 I_75583 (I1287403,I2507,I1287154,I1287460,);
not I_75584 (I1287468,I1287460);
nor I_75585 (I1287140,I1287239,I1287468);
or I_75586 (I1287499,I1287307,I529212);
nor I_75587 (I1287516,I529212,I529194);
nand I_75588 (I1287533,I1287372,I1287516);
nand I_75589 (I1287550,I1287499,I1287533);
DFFARX1 I_75590 (I1287550,I2507,I1287154,I1287143,);
nor I_75591 (I1287581,I1287516,I1287273);
DFFARX1 I_75592 (I1287581,I2507,I1287154,I1287122,);
nor I_75593 (I1287612,I529212,I529197);
DFFARX1 I_75594 (I1287612,I2507,I1287154,I1287638,);
DFFARX1 I_75595 (I1287638,I2507,I1287154,I1287137,);
not I_75596 (I1287660,I1287638);
nand I_75597 (I1287134,I1287660,I1287188);
nand I_75598 (I1287128,I1287660,I1287290);
not I_75599 (I1287732,I2514);
DFFARX1 I_75600 (I635920,I2507,I1287732,I1287758,);
nand I_75601 (I1287766,I1287758,I635923);
not I_75602 (I1287783,I1287766);
DFFARX1 I_75603 (I635935,I2507,I1287732,I1287809,);
not I_75604 (I1287817,I1287809);
not I_75605 (I1287834,I635920);
or I_75606 (I1287851,I635929,I635920);
nor I_75607 (I1287868,I635929,I635920);
or I_75608 (I1287885,I635938,I635929);
DFFARX1 I_75609 (I1287885,I2507,I1287732,I1287724,);
not I_75610 (I1287916,I635941);
nand I_75611 (I1287933,I1287916,I635923);
nand I_75612 (I1287950,I1287834,I1287933);
and I_75613 (I1287703,I1287817,I1287950);
nor I_75614 (I1287981,I635941,I635926);
and I_75615 (I1287998,I1287817,I1287981);
nor I_75616 (I1287709,I1287783,I1287998);
DFFARX1 I_75617 (I1287981,I2507,I1287732,I1288038,);
not I_75618 (I1288046,I1288038);
nor I_75619 (I1287718,I1287817,I1288046);
or I_75620 (I1288077,I1287885,I635932);
nor I_75621 (I1288094,I635932,I635938);
nand I_75622 (I1288111,I1287950,I1288094);
nand I_75623 (I1288128,I1288077,I1288111);
DFFARX1 I_75624 (I1288128,I2507,I1287732,I1287721,);
nor I_75625 (I1288159,I1288094,I1287851);
DFFARX1 I_75626 (I1288159,I2507,I1287732,I1287700,);
nor I_75627 (I1288190,I635932,I635944);
DFFARX1 I_75628 (I1288190,I2507,I1287732,I1288216,);
DFFARX1 I_75629 (I1288216,I2507,I1287732,I1287715,);
not I_75630 (I1288238,I1288216);
nand I_75631 (I1287712,I1288238,I1287766);
nand I_75632 (I1287706,I1288238,I1287868);
not I_75633 (I1288310,I2514);
DFFARX1 I_75634 (I951531,I2507,I1288310,I1288336,);
nand I_75635 (I1288344,I1288336,I951552);
not I_75636 (I1288361,I1288344);
DFFARX1 I_75637 (I951525,I2507,I1288310,I1288387,);
not I_75638 (I1288395,I1288387);
not I_75639 (I1288412,I951546);
or I_75640 (I1288429,I951537,I951546);
nor I_75641 (I1288446,I951537,I951546);
or I_75642 (I1288463,I951540,I951537);
DFFARX1 I_75643 (I1288463,I2507,I1288310,I1288302,);
not I_75644 (I1288494,I951528);
nand I_75645 (I1288511,I1288494,I951543);
nand I_75646 (I1288528,I1288412,I1288511);
and I_75647 (I1288281,I1288395,I1288528);
nor I_75648 (I1288559,I951528,I951525);
and I_75649 (I1288576,I1288395,I1288559);
nor I_75650 (I1288287,I1288361,I1288576);
DFFARX1 I_75651 (I1288559,I2507,I1288310,I1288616,);
not I_75652 (I1288624,I1288616);
nor I_75653 (I1288296,I1288395,I1288624);
or I_75654 (I1288655,I1288463,I951549);
nor I_75655 (I1288672,I951549,I951540);
nand I_75656 (I1288689,I1288528,I1288672);
nand I_75657 (I1288706,I1288655,I1288689);
DFFARX1 I_75658 (I1288706,I2507,I1288310,I1288299,);
nor I_75659 (I1288737,I1288672,I1288429);
DFFARX1 I_75660 (I1288737,I2507,I1288310,I1288278,);
nor I_75661 (I1288768,I951549,I951534);
DFFARX1 I_75662 (I1288768,I2507,I1288310,I1288794,);
DFFARX1 I_75663 (I1288794,I2507,I1288310,I1288293,);
not I_75664 (I1288816,I1288794);
nand I_75665 (I1288290,I1288816,I1288344);
nand I_75666 (I1288284,I1288816,I1288446);
not I_75667 (I1288888,I2514);
DFFARX1 I_75668 (I784860,I2507,I1288888,I1288914,);
nand I_75669 (I1288922,I1288914,I784860);
not I_75670 (I1288939,I1288922);
DFFARX1 I_75671 (I784866,I2507,I1288888,I1288965,);
not I_75672 (I1288973,I1288965);
not I_75673 (I1288990,I784878);
or I_75674 (I1289007,I784863,I784878);
nor I_75675 (I1289024,I784863,I784878);
or I_75676 (I1289041,I784857,I784863);
DFFARX1 I_75677 (I1289041,I2507,I1288888,I1288880,);
not I_75678 (I1289072,I784875);
nand I_75679 (I1289089,I1289072,I784869);
nand I_75680 (I1289106,I1288990,I1289089);
and I_75681 (I1288859,I1288973,I1289106);
nor I_75682 (I1289137,I784875,I784857);
and I_75683 (I1289154,I1288973,I1289137);
nor I_75684 (I1288865,I1288939,I1289154);
DFFARX1 I_75685 (I1289137,I2507,I1288888,I1289194,);
not I_75686 (I1289202,I1289194);
nor I_75687 (I1288874,I1288973,I1289202);
or I_75688 (I1289233,I1289041,I784872);
nor I_75689 (I1289250,I784872,I784857);
nand I_75690 (I1289267,I1289106,I1289250);
nand I_75691 (I1289284,I1289233,I1289267);
DFFARX1 I_75692 (I1289284,I2507,I1288888,I1288877,);
nor I_75693 (I1289315,I1289250,I1289007);
DFFARX1 I_75694 (I1289315,I2507,I1288888,I1288856,);
nor I_75695 (I1289346,I784872,I784863);
DFFARX1 I_75696 (I1289346,I2507,I1288888,I1289372,);
DFFARX1 I_75697 (I1289372,I2507,I1288888,I1288871,);
not I_75698 (I1289394,I1289372);
nand I_75699 (I1288868,I1289394,I1288922);
nand I_75700 (I1288862,I1289394,I1289024);
not I_75701 (I1289466,I2514);
DFFARX1 I_75702 (I893391,I2507,I1289466,I1289492,);
nand I_75703 (I1289500,I1289492,I893412);
not I_75704 (I1289517,I1289500);
DFFARX1 I_75705 (I893385,I2507,I1289466,I1289543,);
not I_75706 (I1289551,I1289543);
not I_75707 (I1289568,I893406);
or I_75708 (I1289585,I893397,I893406);
nor I_75709 (I1289602,I893397,I893406);
or I_75710 (I1289619,I893400,I893397);
DFFARX1 I_75711 (I1289619,I2507,I1289466,I1289458,);
not I_75712 (I1289650,I893388);
nand I_75713 (I1289667,I1289650,I893403);
nand I_75714 (I1289684,I1289568,I1289667);
and I_75715 (I1289437,I1289551,I1289684);
nor I_75716 (I1289715,I893388,I893385);
and I_75717 (I1289732,I1289551,I1289715);
nor I_75718 (I1289443,I1289517,I1289732);
DFFARX1 I_75719 (I1289715,I2507,I1289466,I1289772,);
not I_75720 (I1289780,I1289772);
nor I_75721 (I1289452,I1289551,I1289780);
or I_75722 (I1289811,I1289619,I893409);
nor I_75723 (I1289828,I893409,I893400);
nand I_75724 (I1289845,I1289684,I1289828);
nand I_75725 (I1289862,I1289811,I1289845);
DFFARX1 I_75726 (I1289862,I2507,I1289466,I1289455,);
nor I_75727 (I1289893,I1289828,I1289585);
DFFARX1 I_75728 (I1289893,I2507,I1289466,I1289434,);
nor I_75729 (I1289924,I893409,I893394);
DFFARX1 I_75730 (I1289924,I2507,I1289466,I1289950,);
DFFARX1 I_75731 (I1289950,I2507,I1289466,I1289449,);
not I_75732 (I1289972,I1289950);
nand I_75733 (I1289446,I1289972,I1289500);
nand I_75734 (I1289440,I1289972,I1289602);
not I_75735 (I1290044,I2514);
DFFARX1 I_75736 (I1111564,I2507,I1290044,I1290070,);
nand I_75737 (I1290078,I1290070,I1111549);
not I_75738 (I1290095,I1290078);
DFFARX1 I_75739 (I1111552,I2507,I1290044,I1290121,);
not I_75740 (I1290129,I1290121);
not I_75741 (I1290146,I1111567);
or I_75742 (I1290163,I1111570,I1111567);
nor I_75743 (I1290180,I1111570,I1111567);
or I_75744 (I1290197,I1111546,I1111570);
DFFARX1 I_75745 (I1290197,I2507,I1290044,I1290036,);
not I_75746 (I1290228,I1111558);
nand I_75747 (I1290245,I1290228,I1111561);
nand I_75748 (I1290262,I1290146,I1290245);
and I_75749 (I1290015,I1290129,I1290262);
nor I_75750 (I1290293,I1111558,I1111555);
and I_75751 (I1290310,I1290129,I1290293);
nor I_75752 (I1290021,I1290095,I1290310);
DFFARX1 I_75753 (I1290293,I2507,I1290044,I1290350,);
not I_75754 (I1290358,I1290350);
nor I_75755 (I1290030,I1290129,I1290358);
or I_75756 (I1290389,I1290197,I1111546);
nor I_75757 (I1290406,I1111546,I1111546);
nand I_75758 (I1290423,I1290262,I1290406);
nand I_75759 (I1290440,I1290389,I1290423);
DFFARX1 I_75760 (I1290440,I2507,I1290044,I1290033,);
nor I_75761 (I1290471,I1290406,I1290163);
DFFARX1 I_75762 (I1290471,I2507,I1290044,I1290012,);
nor I_75763 (I1290502,I1111546,I1111549);
DFFARX1 I_75764 (I1290502,I2507,I1290044,I1290528,);
DFFARX1 I_75765 (I1290528,I2507,I1290044,I1290027,);
not I_75766 (I1290550,I1290528);
nand I_75767 (I1290024,I1290550,I1290078);
nand I_75768 (I1290018,I1290550,I1290180);
not I_75769 (I1290622,I2514);
DFFARX1 I_75770 (I1298071,I2507,I1290622,I1290648,);
nand I_75771 (I1290656,I1290648,I1298065);
not I_75772 (I1290673,I1290656);
DFFARX1 I_75773 (I1298080,I2507,I1290622,I1290699,);
not I_75774 (I1290707,I1290699);
not I_75775 (I1290724,I1298056);
or I_75776 (I1290741,I1298053,I1298056);
nor I_75777 (I1290758,I1298053,I1298056);
or I_75778 (I1290775,I1298059,I1298053);
DFFARX1 I_75779 (I1290775,I2507,I1290622,I1290614,);
not I_75780 (I1290806,I1298053);
nand I_75781 (I1290823,I1290806,I1298068);
nand I_75782 (I1290840,I1290724,I1290823);
and I_75783 (I1290593,I1290707,I1290840);
nor I_75784 (I1290871,I1298053,I1298062);
and I_75785 (I1290888,I1290707,I1290871);
nor I_75786 (I1290599,I1290673,I1290888);
DFFARX1 I_75787 (I1290871,I2507,I1290622,I1290928,);
not I_75788 (I1290936,I1290928);
nor I_75789 (I1290608,I1290707,I1290936);
or I_75790 (I1290967,I1290775,I1298077);
nor I_75791 (I1290984,I1298077,I1298059);
nand I_75792 (I1291001,I1290840,I1290984);
nand I_75793 (I1291018,I1290967,I1291001);
DFFARX1 I_75794 (I1291018,I2507,I1290622,I1290611,);
nor I_75795 (I1291049,I1290984,I1290741);
DFFARX1 I_75796 (I1291049,I2507,I1290622,I1290590,);
nor I_75797 (I1291080,I1298077,I1298074);
DFFARX1 I_75798 (I1291080,I2507,I1290622,I1291106,);
DFFARX1 I_75799 (I1291106,I2507,I1290622,I1290605,);
not I_75800 (I1291128,I1291106);
nand I_75801 (I1290602,I1291128,I1290656);
nand I_75802 (I1290596,I1291128,I1290758);
not I_75803 (I1291200,I2514);
DFFARX1 I_75804 (I926983,I2507,I1291200,I1291226,);
nand I_75805 (I1291234,I1291226,I927004);
not I_75806 (I1291251,I1291234);
DFFARX1 I_75807 (I926977,I2507,I1291200,I1291277,);
not I_75808 (I1291285,I1291277);
not I_75809 (I1291302,I926998);
or I_75810 (I1291319,I926989,I926998);
nor I_75811 (I1291336,I926989,I926998);
or I_75812 (I1291353,I926992,I926989);
DFFARX1 I_75813 (I1291353,I2507,I1291200,I1291192,);
not I_75814 (I1291384,I926980);
nand I_75815 (I1291401,I1291384,I926995);
nand I_75816 (I1291418,I1291302,I1291401);
and I_75817 (I1291171,I1291285,I1291418);
nor I_75818 (I1291449,I926980,I926977);
and I_75819 (I1291466,I1291285,I1291449);
nor I_75820 (I1291177,I1291251,I1291466);
DFFARX1 I_75821 (I1291449,I2507,I1291200,I1291506,);
not I_75822 (I1291514,I1291506);
nor I_75823 (I1291186,I1291285,I1291514);
or I_75824 (I1291545,I1291353,I927001);
nor I_75825 (I1291562,I927001,I926992);
nand I_75826 (I1291579,I1291418,I1291562);
nand I_75827 (I1291596,I1291545,I1291579);
DFFARX1 I_75828 (I1291596,I2507,I1291200,I1291189,);
nor I_75829 (I1291627,I1291562,I1291319);
DFFARX1 I_75830 (I1291627,I2507,I1291200,I1291168,);
nor I_75831 (I1291658,I927001,I926986);
DFFARX1 I_75832 (I1291658,I2507,I1291200,I1291684,);
DFFARX1 I_75833 (I1291684,I2507,I1291200,I1291183,);
not I_75834 (I1291706,I1291684);
nand I_75835 (I1291180,I1291706,I1291234);
nand I_75836 (I1291174,I1291706,I1291336);
not I_75837 (I1291778,I2514);
DFFARX1 I_75838 (I801724,I2507,I1291778,I1291804,);
nand I_75839 (I1291812,I1291804,I801724);
not I_75840 (I1291829,I1291812);
DFFARX1 I_75841 (I801730,I2507,I1291778,I1291855,);
not I_75842 (I1291863,I1291855);
not I_75843 (I1291880,I801742);
or I_75844 (I1291897,I801727,I801742);
nor I_75845 (I1291914,I801727,I801742);
or I_75846 (I1291931,I801721,I801727);
DFFARX1 I_75847 (I1291931,I2507,I1291778,I1291770,);
not I_75848 (I1291962,I801739);
nand I_75849 (I1291979,I1291962,I801733);
nand I_75850 (I1291996,I1291880,I1291979);
and I_75851 (I1291749,I1291863,I1291996);
nor I_75852 (I1292027,I801739,I801721);
and I_75853 (I1292044,I1291863,I1292027);
nor I_75854 (I1291755,I1291829,I1292044);
DFFARX1 I_75855 (I1292027,I2507,I1291778,I1292084,);
not I_75856 (I1292092,I1292084);
nor I_75857 (I1291764,I1291863,I1292092);
or I_75858 (I1292123,I1291931,I801736);
nor I_75859 (I1292140,I801736,I801721);
nand I_75860 (I1292157,I1291996,I1292140);
nand I_75861 (I1292174,I1292123,I1292157);
DFFARX1 I_75862 (I1292174,I2507,I1291778,I1291767,);
nor I_75863 (I1292205,I1292140,I1291897);
DFFARX1 I_75864 (I1292205,I2507,I1291778,I1291746,);
nor I_75865 (I1292236,I801736,I801727);
DFFARX1 I_75866 (I1292236,I2507,I1291778,I1292262,);
DFFARX1 I_75867 (I1292262,I2507,I1291778,I1291761,);
not I_75868 (I1292284,I1292262);
nand I_75869 (I1291758,I1292284,I1291812);
nand I_75870 (I1291752,I1292284,I1291914);
not I_75871 (I1292356,I2514);
DFFARX1 I_75872 (I281816,I2507,I1292356,I1292382,);
nand I_75873 (I1292390,I1292382,I281837);
not I_75874 (I1292407,I1292390);
DFFARX1 I_75875 (I281831,I2507,I1292356,I1292433,);
not I_75876 (I1292441,I1292433);
not I_75877 (I1292458,I281819);
or I_75878 (I1292475,I281834,I281819);
nor I_75879 (I1292492,I281834,I281819);
or I_75880 (I1292509,I281825,I281834);
DFFARX1 I_75881 (I1292509,I2507,I1292356,I1292348,);
not I_75882 (I1292540,I281813);
nand I_75883 (I1292557,I1292540,I281810);
nand I_75884 (I1292574,I1292458,I1292557);
and I_75885 (I1292327,I1292441,I1292574);
nor I_75886 (I1292605,I281813,I281822);
and I_75887 (I1292622,I1292441,I1292605);
nor I_75888 (I1292333,I1292407,I1292622);
DFFARX1 I_75889 (I1292605,I2507,I1292356,I1292662,);
not I_75890 (I1292670,I1292662);
nor I_75891 (I1292342,I1292441,I1292670);
or I_75892 (I1292701,I1292509,I281828);
nor I_75893 (I1292718,I281828,I281825);
nand I_75894 (I1292735,I1292574,I1292718);
nand I_75895 (I1292752,I1292701,I1292735);
DFFARX1 I_75896 (I1292752,I2507,I1292356,I1292345,);
nor I_75897 (I1292783,I1292718,I1292475);
DFFARX1 I_75898 (I1292783,I2507,I1292356,I1292324,);
nor I_75899 (I1292814,I281828,I281810);
DFFARX1 I_75900 (I1292814,I2507,I1292356,I1292840,);
DFFARX1 I_75901 (I1292840,I2507,I1292356,I1292339,);
not I_75902 (I1292862,I1292840);
nand I_75903 (I1292336,I1292862,I1292390);
nand I_75904 (I1292330,I1292862,I1292492);
not I_75905 (I1292934,I2514);
DFFARX1 I_75906 (I1333896,I2507,I1292934,I1292960,);
nand I_75907 (I1292968,I1292960,I1333887);
not I_75908 (I1292985,I1292968);
DFFARX1 I_75909 (I1333872,I2507,I1292934,I1293011,);
not I_75910 (I1293019,I1293011);
not I_75911 (I1293036,I1333875);
or I_75912 (I1293053,I1333884,I1333875);
nor I_75913 (I1293070,I1333884,I1333875);
or I_75914 (I1293087,I1333881,I1333884);
DFFARX1 I_75915 (I1293087,I2507,I1292934,I1292926,);
not I_75916 (I1293118,I1333893);
nand I_75917 (I1293135,I1293118,I1333872);
nand I_75918 (I1293152,I1293036,I1293135);
and I_75919 (I1292905,I1293019,I1293152);
nor I_75920 (I1293183,I1333893,I1333878);
and I_75921 (I1293200,I1293019,I1293183);
nor I_75922 (I1292911,I1292985,I1293200);
DFFARX1 I_75923 (I1293183,I2507,I1292934,I1293240,);
not I_75924 (I1293248,I1293240);
nor I_75925 (I1292920,I1293019,I1293248);
or I_75926 (I1293279,I1293087,I1333899);
nor I_75927 (I1293296,I1333899,I1333881);
nand I_75928 (I1293313,I1293152,I1293296);
nand I_75929 (I1293330,I1293279,I1293313);
DFFARX1 I_75930 (I1293330,I2507,I1292934,I1292923,);
nor I_75931 (I1293361,I1293296,I1293053);
DFFARX1 I_75932 (I1293361,I2507,I1292934,I1292902,);
nor I_75933 (I1293392,I1333899,I1333890);
DFFARX1 I_75934 (I1293392,I2507,I1292934,I1293418,);
DFFARX1 I_75935 (I1293418,I2507,I1292934,I1292917,);
not I_75936 (I1293440,I1293418);
nand I_75937 (I1292914,I1293440,I1292968);
nand I_75938 (I1292908,I1293440,I1293070);
not I_75939 (I1293512,I2514);
DFFARX1 I_75940 (I465362,I2507,I1293512,I1293538,);
nand I_75941 (I1293546,I1293538,I465371);
not I_75942 (I1293563,I1293546);
DFFARX1 I_75943 (I465359,I2507,I1293512,I1293589,);
not I_75944 (I1293597,I1293589);
not I_75945 (I1293614,I465365);
or I_75946 (I1293631,I465359,I465365);
nor I_75947 (I1293648,I465359,I465365);
or I_75948 (I1293665,I465374,I465359);
DFFARX1 I_75949 (I1293665,I2507,I1293512,I1293504,);
not I_75950 (I1293696,I465368);
nand I_75951 (I1293713,I1293696,I465383);
nand I_75952 (I1293730,I1293614,I1293713);
and I_75953 (I1293483,I1293597,I1293730);
nor I_75954 (I1293761,I465368,I465386);
and I_75955 (I1293778,I1293597,I1293761);
nor I_75956 (I1293489,I1293563,I1293778);
DFFARX1 I_75957 (I1293761,I2507,I1293512,I1293818,);
not I_75958 (I1293826,I1293818);
nor I_75959 (I1293498,I1293597,I1293826);
or I_75960 (I1293857,I1293665,I465377);
nor I_75961 (I1293874,I465377,I465374);
nand I_75962 (I1293891,I1293730,I1293874);
nand I_75963 (I1293908,I1293857,I1293891);
DFFARX1 I_75964 (I1293908,I2507,I1293512,I1293501,);
nor I_75965 (I1293939,I1293874,I1293631);
DFFARX1 I_75966 (I1293939,I2507,I1293512,I1293480,);
nor I_75967 (I1293970,I465377,I465380);
DFFARX1 I_75968 (I1293970,I2507,I1293512,I1293996,);
DFFARX1 I_75969 (I1293996,I2507,I1293512,I1293495,);
not I_75970 (I1294018,I1293996);
nand I_75971 (I1293492,I1294018,I1293546);
nand I_75972 (I1293486,I1294018,I1293648);
not I_75973 (I1294090,I2514);
DFFARX1 I_75974 (I1018565,I2507,I1294090,I1294116,);
nand I_75975 (I1294124,I1294116,I1018562);
not I_75976 (I1294141,I1294124);
DFFARX1 I_75977 (I1018562,I2507,I1294090,I1294167,);
not I_75978 (I1294175,I1294167);
not I_75979 (I1294192,I1018559);
or I_75980 (I1294209,I1018568,I1018559);
nor I_75981 (I1294226,I1018568,I1018559);
or I_75982 (I1294243,I1018571,I1018568);
DFFARX1 I_75983 (I1294243,I2507,I1294090,I1294082,);
not I_75984 (I1294274,I1018559);
nand I_75985 (I1294291,I1294274,I1018556);
nand I_75986 (I1294308,I1294192,I1294291);
and I_75987 (I1294061,I1294175,I1294308);
nor I_75988 (I1294339,I1018559,I1018574);
and I_75989 (I1294356,I1294175,I1294339);
nor I_75990 (I1294067,I1294141,I1294356);
DFFARX1 I_75991 (I1294339,I2507,I1294090,I1294396,);
not I_75992 (I1294404,I1294396);
nor I_75993 (I1294076,I1294175,I1294404);
or I_75994 (I1294435,I1294243,I1018577);
nor I_75995 (I1294452,I1018577,I1018571);
nand I_75996 (I1294469,I1294308,I1294452);
nand I_75997 (I1294486,I1294435,I1294469);
DFFARX1 I_75998 (I1294486,I2507,I1294090,I1294079,);
nor I_75999 (I1294517,I1294452,I1294209);
DFFARX1 I_76000 (I1294517,I2507,I1294090,I1294058,);
nor I_76001 (I1294548,I1018577,I1018556);
DFFARX1 I_76002 (I1294548,I2507,I1294090,I1294574,);
DFFARX1 I_76003 (I1294574,I2507,I1294090,I1294073,);
not I_76004 (I1294596,I1294574);
nand I_76005 (I1294070,I1294596,I1294124);
nand I_76006 (I1294064,I1294596,I1294226);
not I_76007 (I1294668,I2514);
DFFARX1 I_76008 (I27462,I2507,I1294668,I1294694,);
nand I_76009 (I1294702,I1294694,I27456);
not I_76010 (I1294719,I1294702);
DFFARX1 I_76011 (I27474,I2507,I1294668,I1294745,);
not I_76012 (I1294753,I1294745);
not I_76013 (I1294770,I27477);
or I_76014 (I1294787,I27480,I27477);
nor I_76015 (I1294804,I27480,I27477);
or I_76016 (I1294821,I27465,I27480);
DFFARX1 I_76017 (I1294821,I2507,I1294668,I1294660,);
not I_76018 (I1294852,I27468);
nand I_76019 (I1294869,I1294852,I27471);
nand I_76020 (I1294886,I1294770,I1294869);
and I_76021 (I1294639,I1294753,I1294886);
nor I_76022 (I1294917,I27468,I27459);
and I_76023 (I1294934,I1294753,I1294917);
nor I_76024 (I1294645,I1294719,I1294934);
DFFARX1 I_76025 (I1294917,I2507,I1294668,I1294974,);
not I_76026 (I1294982,I1294974);
nor I_76027 (I1294654,I1294753,I1294982);
or I_76028 (I1295013,I1294821,I27459);
nor I_76029 (I1295030,I27459,I27465);
nand I_76030 (I1295047,I1294886,I1295030);
nand I_76031 (I1295064,I1295013,I1295047);
DFFARX1 I_76032 (I1295064,I2507,I1294668,I1294657,);
nor I_76033 (I1295095,I1295030,I1294787);
DFFARX1 I_76034 (I1295095,I2507,I1294668,I1294636,);
nor I_76035 (I1295126,I27459,I27456);
DFFARX1 I_76036 (I1295126,I2507,I1294668,I1295152,);
DFFARX1 I_76037 (I1295152,I2507,I1294668,I1294651,);
not I_76038 (I1295174,I1295152);
nand I_76039 (I1294648,I1295174,I1294702);
nand I_76040 (I1294642,I1295174,I1294804);
not I_76041 (I1295246,I2514);
DFFARX1 I_76042 (I1326756,I2507,I1295246,I1295272,);
nand I_76043 (I1295280,I1295272,I1326747);
not I_76044 (I1295297,I1295280);
DFFARX1 I_76045 (I1326732,I2507,I1295246,I1295323,);
not I_76046 (I1295331,I1295323);
not I_76047 (I1295348,I1326735);
or I_76048 (I1295365,I1326744,I1326735);
nor I_76049 (I1295382,I1326744,I1326735);
or I_76050 (I1295399,I1326741,I1326744);
DFFARX1 I_76051 (I1295399,I2507,I1295246,I1295238,);
not I_76052 (I1295430,I1326753);
nand I_76053 (I1295447,I1295430,I1326732);
nand I_76054 (I1295464,I1295348,I1295447);
and I_76055 (I1295217,I1295331,I1295464);
nor I_76056 (I1295495,I1326753,I1326738);
and I_76057 (I1295512,I1295331,I1295495);
nor I_76058 (I1295223,I1295297,I1295512);
DFFARX1 I_76059 (I1295495,I2507,I1295246,I1295552,);
not I_76060 (I1295560,I1295552);
nor I_76061 (I1295232,I1295331,I1295560);
or I_76062 (I1295591,I1295399,I1326759);
nor I_76063 (I1295608,I1326759,I1326741);
nand I_76064 (I1295625,I1295464,I1295608);
nand I_76065 (I1295642,I1295591,I1295625);
DFFARX1 I_76066 (I1295642,I2507,I1295246,I1295235,);
nor I_76067 (I1295673,I1295608,I1295365);
DFFARX1 I_76068 (I1295673,I2507,I1295246,I1295214,);
nor I_76069 (I1295704,I1326759,I1326750);
DFFARX1 I_76070 (I1295704,I2507,I1295246,I1295730,);
DFFARX1 I_76071 (I1295730,I2507,I1295246,I1295229,);
not I_76072 (I1295752,I1295730);
nand I_76073 (I1295226,I1295752,I1295280);
nand I_76074 (I1295220,I1295752,I1295382);
not I_76075 (I1295824,I2514);
DFFARX1 I_76076 (I582169,I2507,I1295824,I1295850,);
nand I_76077 (I1295858,I1295850,I582184);
not I_76078 (I1295875,I1295858);
DFFARX1 I_76079 (I582166,I2507,I1295824,I1295901,);
not I_76080 (I1295909,I1295901);
not I_76081 (I1295926,I582175);
or I_76082 (I1295943,I582169,I582175);
nor I_76083 (I1295960,I582169,I582175);
or I_76084 (I1295977,I582166,I582169);
DFFARX1 I_76085 (I1295977,I2507,I1295824,I1295816,);
not I_76086 (I1296008,I582187);
nand I_76087 (I1296025,I1296008,I582190);
nand I_76088 (I1296042,I1295926,I1296025);
and I_76089 (I1295795,I1295909,I1296042);
nor I_76090 (I1296073,I582187,I582172);
and I_76091 (I1296090,I1295909,I1296073);
nor I_76092 (I1295801,I1295875,I1296090);
DFFARX1 I_76093 (I1296073,I2507,I1295824,I1296130,);
not I_76094 (I1296138,I1296130);
nor I_76095 (I1295810,I1295909,I1296138);
or I_76096 (I1296169,I1295977,I582178);
nor I_76097 (I1296186,I582178,I582166);
nand I_76098 (I1296203,I1296042,I1296186);
nand I_76099 (I1296220,I1296169,I1296203);
DFFARX1 I_76100 (I1296220,I2507,I1295824,I1295813,);
nor I_76101 (I1296251,I1296186,I1295943);
DFFARX1 I_76102 (I1296251,I2507,I1295824,I1295792,);
nor I_76103 (I1296282,I582178,I582181);
DFFARX1 I_76104 (I1296282,I2507,I1295824,I1296308,);
DFFARX1 I_76105 (I1296308,I2507,I1295824,I1295807,);
not I_76106 (I1296330,I1296308);
nand I_76107 (I1295804,I1296330,I1295858);
nand I_76108 (I1295798,I1296330,I1295960);
not I_76109 (I1296405,I2514);
DFFARX1 I_76110 (I1017446,I2507,I1296405,I1296431,);
nand I_76111 (I1296439,I1296431,I1017449);
not I_76112 (I1296456,I1296439);
DFFARX1 I_76113 (I1017437,I2507,I1296405,I1296482,);
not I_76114 (I1296490,I1296482);
nor I_76115 (I1296507,I1017455,I1017452);
not I_76116 (I1296524,I1296507);
DFFARX1 I_76117 (I1296524,I2507,I1296405,I1296391,);
or I_76118 (I1296555,I1017434,I1017455);
DFFARX1 I_76119 (I1296555,I2507,I1296405,I1296394,);
not I_76120 (I1296586,I1017434);
nor I_76121 (I1296603,I1296586,I1017437);
nor I_76122 (I1296620,I1296603,I1017452);
nor I_76123 (I1296637,I1017437,I1017440);
nor I_76124 (I1296654,I1296490,I1296637);
nor I_76125 (I1296379,I1296456,I1296654);
not I_76126 (I1296685,I1296637);
nand I_76127 (I1296382,I1296685,I1296439);
nand I_76128 (I1296376,I1296685,I1296507);
nor I_76129 (I1296373,I1296637,I1296620);
nor I_76130 (I1296744,I1017443,I1017434);
not I_76131 (I1296761,I1296744);
DFFARX1 I_76132 (I1296744,I2507,I1296405,I1296787,);
not I_76133 (I1296397,I1296787);
nor I_76134 (I1296809,I1017443,I1017440);
DFFARX1 I_76135 (I1296809,I2507,I1296405,I1296835,);
and I_76136 (I1296843,I1296835,I1017455);
nor I_76137 (I1296860,I1296843,I1296761);
DFFARX1 I_76138 (I1296860,I2507,I1296405,I1296388,);
nor I_76139 (I1296891,I1296835,I1296620);
DFFARX1 I_76140 (I1296891,I2507,I1296405,I1296370,);
nor I_76141 (I1296385,I1296835,I1296524);
not I_76142 (I1296966,I2514);
DFFARX1 I_76143 (I960593,I2507,I1296966,I1296992,);
nand I_76144 (I1297000,I1296992,I960575);
not I_76145 (I1297017,I1297000);
DFFARX1 I_76146 (I960587,I2507,I1296966,I1297043,);
not I_76147 (I1297051,I1297043);
nor I_76148 (I1297068,I960569,I960569);
not I_76149 (I1297085,I1297068);
DFFARX1 I_76150 (I1297085,I2507,I1296966,I1296952,);
or I_76151 (I1297116,I960581,I960569);
DFFARX1 I_76152 (I1297116,I2507,I1296966,I1296955,);
not I_76153 (I1297147,I960596);
nor I_76154 (I1297164,I1297147,I960584);
nor I_76155 (I1297181,I1297164,I960569);
nor I_76156 (I1297198,I960584,I960572);
nor I_76157 (I1297215,I1297051,I1297198);
nor I_76158 (I1296940,I1297017,I1297215);
not I_76159 (I1297246,I1297198);
nand I_76160 (I1296943,I1297246,I1297000);
nand I_76161 (I1296937,I1297246,I1297068);
nor I_76162 (I1296934,I1297198,I1297181);
nor I_76163 (I1297305,I960578,I960581);
not I_76164 (I1297322,I1297305);
DFFARX1 I_76165 (I1297305,I2507,I1296966,I1297348,);
not I_76166 (I1296958,I1297348);
nor I_76167 (I1297370,I960578,I960590);
DFFARX1 I_76168 (I1297370,I2507,I1296966,I1297396,);
and I_76169 (I1297404,I1297396,I960569);
nor I_76170 (I1297421,I1297404,I1297322);
DFFARX1 I_76171 (I1297421,I2507,I1296966,I1296949,);
nor I_76172 (I1297452,I1297396,I1297181);
DFFARX1 I_76173 (I1297452,I2507,I1296966,I1296931,);
nor I_76174 (I1296946,I1297396,I1297085);
not I_76175 (I1297527,I2514);
DFFARX1 I_76176 (I58573,I2507,I1297527,I1297553,);
nand I_76177 (I1297561,I1297553,I58564);
not I_76178 (I1297578,I1297561);
DFFARX1 I_76179 (I58552,I2507,I1297527,I1297604,);
not I_76180 (I1297612,I1297604);
nor I_76181 (I1297629,I58555,I58552);
not I_76182 (I1297646,I1297629);
DFFARX1 I_76183 (I1297646,I2507,I1297527,I1297513,);
or I_76184 (I1297677,I58549,I58555);
DFFARX1 I_76185 (I1297677,I2507,I1297527,I1297516,);
not I_76186 (I1297708,I58558);
nor I_76187 (I1297725,I1297708,I58549);
nor I_76188 (I1297742,I1297725,I58552);
nor I_76189 (I1297759,I58549,I58561);
nor I_76190 (I1297776,I1297612,I1297759);
nor I_76191 (I1297501,I1297578,I1297776);
not I_76192 (I1297807,I1297759);
nand I_76193 (I1297504,I1297807,I1297561);
nand I_76194 (I1297498,I1297807,I1297629);
nor I_76195 (I1297495,I1297759,I1297742);
nor I_76196 (I1297866,I58567,I58549);
not I_76197 (I1297883,I1297866);
DFFARX1 I_76198 (I1297866,I2507,I1297527,I1297909,);
not I_76199 (I1297519,I1297909);
nor I_76200 (I1297931,I58567,I58570);
DFFARX1 I_76201 (I1297931,I2507,I1297527,I1297957,);
and I_76202 (I1297965,I1297957,I58555);
nor I_76203 (I1297982,I1297965,I1297883);
DFFARX1 I_76204 (I1297982,I2507,I1297527,I1297510,);
nor I_76205 (I1298013,I1297957,I1297742);
DFFARX1 I_76206 (I1298013,I2507,I1297527,I1297492,);
nor I_76207 (I1297507,I1297957,I1297646);
not I_76208 (I1298088,I2514);
DFFARX1 I_76209 (I835452,I2507,I1298088,I1298114,);
nand I_76210 (I1298122,I1298114,I835470);
not I_76211 (I1298139,I1298122);
DFFARX1 I_76212 (I835449,I2507,I1298088,I1298165,);
not I_76213 (I1298173,I1298165);
nor I_76214 (I1298190,I835464,I835458);
not I_76215 (I1298207,I1298190);
DFFARX1 I_76216 (I1298207,I2507,I1298088,I1298074,);
or I_76217 (I1298238,I835455,I835464);
DFFARX1 I_76218 (I1298238,I2507,I1298088,I1298077,);
not I_76219 (I1298269,I835455);
nor I_76220 (I1298286,I1298269,I835461);
nor I_76221 (I1298303,I1298286,I835458);
nor I_76222 (I1298320,I835461,I835449);
nor I_76223 (I1298337,I1298173,I1298320);
nor I_76224 (I1298062,I1298139,I1298337);
not I_76225 (I1298368,I1298320);
nand I_76226 (I1298065,I1298368,I1298122);
nand I_76227 (I1298059,I1298368,I1298190);
nor I_76228 (I1298056,I1298320,I1298303);
nor I_76229 (I1298427,I835452,I835455);
not I_76230 (I1298444,I1298427);
DFFARX1 I_76231 (I1298427,I2507,I1298088,I1298470,);
not I_76232 (I1298080,I1298470);
nor I_76233 (I1298492,I835452,I835467);
DFFARX1 I_76234 (I1298492,I2507,I1298088,I1298518,);
and I_76235 (I1298526,I1298518,I835464);
nor I_76236 (I1298543,I1298526,I1298444);
DFFARX1 I_76237 (I1298543,I2507,I1298088,I1298071,);
nor I_76238 (I1298574,I1298518,I1298303);
DFFARX1 I_76239 (I1298574,I2507,I1298088,I1298053,);
nor I_76240 (I1298068,I1298518,I1298207);
not I_76241 (I1298649,I2514);
DFFARX1 I_76242 (I558492,I2507,I1298649,I1298675,);
nand I_76243 (I1298683,I1298675,I558471);
not I_76244 (I1298700,I1298683);
DFFARX1 I_76245 (I558483,I2507,I1298649,I1298726,);
not I_76246 (I1298734,I1298726);
nor I_76247 (I1298751,I558471,I558480);
not I_76248 (I1298768,I1298751);
DFFARX1 I_76249 (I1298768,I2507,I1298649,I1298635,);
or I_76250 (I1298799,I558474,I558471);
DFFARX1 I_76251 (I1298799,I2507,I1298649,I1298638,);
not I_76252 (I1298830,I558477);
nor I_76253 (I1298847,I1298830,I558468);
nor I_76254 (I1298864,I1298847,I558480);
nor I_76255 (I1298881,I558468,I558486);
nor I_76256 (I1298898,I1298734,I1298881);
nor I_76257 (I1298623,I1298700,I1298898);
not I_76258 (I1298929,I1298881);
nand I_76259 (I1298626,I1298929,I1298683);
nand I_76260 (I1298620,I1298929,I1298751);
nor I_76261 (I1298617,I1298881,I1298864);
nor I_76262 (I1298988,I558489,I558474);
not I_76263 (I1299005,I1298988);
DFFARX1 I_76264 (I1298988,I2507,I1298649,I1299031,);
not I_76265 (I1298641,I1299031);
nor I_76266 (I1299053,I558489,I558468);
DFFARX1 I_76267 (I1299053,I2507,I1298649,I1299079,);
and I_76268 (I1299087,I1299079,I558471);
nor I_76269 (I1299104,I1299087,I1299005);
DFFARX1 I_76270 (I1299104,I2507,I1298649,I1298632,);
nor I_76271 (I1299135,I1299079,I1298864);
DFFARX1 I_76272 (I1299135,I2507,I1298649,I1298614,);
nor I_76273 (I1298629,I1299079,I1298768);
not I_76274 (I1299210,I2514);
DFFARX1 I_76275 (I1325557,I2507,I1299210,I1299236,);
nand I_76276 (I1299244,I1299236,I1325551);
not I_76277 (I1299261,I1299244);
DFFARX1 I_76278 (I1325569,I2507,I1299210,I1299287,);
not I_76279 (I1299295,I1299287);
nor I_76280 (I1299312,I1325554,I1325545);
not I_76281 (I1299329,I1299312);
DFFARX1 I_76282 (I1299329,I2507,I1299210,I1299196,);
or I_76283 (I1299360,I1325560,I1325554);
DFFARX1 I_76284 (I1299360,I2507,I1299210,I1299199,);
not I_76285 (I1299391,I1325563);
nor I_76286 (I1299408,I1299391,I1325566);
nor I_76287 (I1299425,I1299408,I1325545);
nor I_76288 (I1299442,I1325566,I1325548);
nor I_76289 (I1299459,I1299295,I1299442);
nor I_76290 (I1299184,I1299261,I1299459);
not I_76291 (I1299490,I1299442);
nand I_76292 (I1299187,I1299490,I1299244);
nand I_76293 (I1299181,I1299490,I1299312);
nor I_76294 (I1299178,I1299442,I1299425);
nor I_76295 (I1299549,I1325542,I1325560);
not I_76296 (I1299566,I1299549);
DFFARX1 I_76297 (I1299549,I2507,I1299210,I1299592,);
not I_76298 (I1299202,I1299592);
nor I_76299 (I1299614,I1325542,I1325542);
DFFARX1 I_76300 (I1299614,I2507,I1299210,I1299640,);
and I_76301 (I1299648,I1299640,I1325554);
nor I_76302 (I1299665,I1299648,I1299566);
DFFARX1 I_76303 (I1299665,I2507,I1299210,I1299193,);
nor I_76304 (I1299696,I1299640,I1299425);
DFFARX1 I_76305 (I1299696,I2507,I1299210,I1299175,);
nor I_76306 (I1299190,I1299640,I1299329);
not I_76307 (I1299771,I2514);
DFFARX1 I_76308 (I817007,I2507,I1299771,I1299797,);
nand I_76309 (I1299805,I1299797,I817025);
not I_76310 (I1299822,I1299805);
DFFARX1 I_76311 (I817004,I2507,I1299771,I1299848,);
not I_76312 (I1299856,I1299848);
nor I_76313 (I1299873,I817019,I817013);
not I_76314 (I1299890,I1299873);
DFFARX1 I_76315 (I1299890,I2507,I1299771,I1299757,);
or I_76316 (I1299921,I817010,I817019);
DFFARX1 I_76317 (I1299921,I2507,I1299771,I1299760,);
not I_76318 (I1299952,I817010);
nor I_76319 (I1299969,I1299952,I817016);
nor I_76320 (I1299986,I1299969,I817013);
nor I_76321 (I1300003,I817016,I817004);
nor I_76322 (I1300020,I1299856,I1300003);
nor I_76323 (I1299745,I1299822,I1300020);
not I_76324 (I1300051,I1300003);
nand I_76325 (I1299748,I1300051,I1299805);
nand I_76326 (I1299742,I1300051,I1299873);
nor I_76327 (I1299739,I1300003,I1299986);
nor I_76328 (I1300110,I817007,I817010);
not I_76329 (I1300127,I1300110);
DFFARX1 I_76330 (I1300110,I2507,I1299771,I1300153,);
not I_76331 (I1299763,I1300153);
nor I_76332 (I1300175,I817007,I817022);
DFFARX1 I_76333 (I1300175,I2507,I1299771,I1300201,);
and I_76334 (I1300209,I1300201,I817019);
nor I_76335 (I1300226,I1300209,I1300127);
DFFARX1 I_76336 (I1300226,I2507,I1299771,I1299754,);
nor I_76337 (I1300257,I1300201,I1299986);
DFFARX1 I_76338 (I1300257,I2507,I1299771,I1299736,);
nor I_76339 (I1299751,I1300201,I1299890);
not I_76340 (I1300332,I2514);
DFFARX1 I_76341 (I332423,I2507,I1300332,I1300358,);
nand I_76342 (I1300366,I1300358,I332402);
not I_76343 (I1300383,I1300366);
DFFARX1 I_76344 (I332411,I2507,I1300332,I1300409,);
not I_76345 (I1300417,I1300409);
nor I_76346 (I1300434,I332405,I332417);
not I_76347 (I1300451,I1300434);
DFFARX1 I_76348 (I1300451,I2507,I1300332,I1300318,);
or I_76349 (I1300482,I332408,I332405);
DFFARX1 I_76350 (I1300482,I2507,I1300332,I1300321,);
not I_76351 (I1300513,I332429);
nor I_76352 (I1300530,I1300513,I332414);
nor I_76353 (I1300547,I1300530,I332417);
nor I_76354 (I1300564,I332414,I332402);
nor I_76355 (I1300581,I1300417,I1300564);
nor I_76356 (I1300306,I1300383,I1300581);
not I_76357 (I1300612,I1300564);
nand I_76358 (I1300309,I1300612,I1300366);
nand I_76359 (I1300303,I1300612,I1300434);
nor I_76360 (I1300300,I1300564,I1300547);
nor I_76361 (I1300671,I332420,I332408);
not I_76362 (I1300688,I1300671);
DFFARX1 I_76363 (I1300671,I2507,I1300332,I1300714,);
not I_76364 (I1300324,I1300714);
nor I_76365 (I1300736,I332420,I332426);
DFFARX1 I_76366 (I1300736,I2507,I1300332,I1300762,);
and I_76367 (I1300770,I1300762,I332405);
nor I_76368 (I1300787,I1300770,I1300688);
DFFARX1 I_76369 (I1300787,I2507,I1300332,I1300315,);
nor I_76370 (I1300818,I1300762,I1300547);
DFFARX1 I_76371 (I1300818,I2507,I1300332,I1300297,);
nor I_76372 (I1300312,I1300762,I1300451);
not I_76373 (I1300893,I2514);
DFFARX1 I_76374 (I1341622,I2507,I1300893,I1300919,);
nand I_76375 (I1300927,I1300919,I1341616);
not I_76376 (I1300944,I1300927);
DFFARX1 I_76377 (I1341634,I2507,I1300893,I1300970,);
not I_76378 (I1300978,I1300970);
nor I_76379 (I1300995,I1341619,I1341610);
not I_76380 (I1301012,I1300995);
DFFARX1 I_76381 (I1301012,I2507,I1300893,I1300879,);
or I_76382 (I1301043,I1341625,I1341619);
DFFARX1 I_76383 (I1301043,I2507,I1300893,I1300882,);
not I_76384 (I1301074,I1341628);
nor I_76385 (I1301091,I1301074,I1341631);
nor I_76386 (I1301108,I1301091,I1341610);
nor I_76387 (I1301125,I1341631,I1341613);
nor I_76388 (I1301142,I1300978,I1301125);
nor I_76389 (I1300867,I1300944,I1301142);
not I_76390 (I1301173,I1301125);
nand I_76391 (I1300870,I1301173,I1300927);
nand I_76392 (I1300864,I1301173,I1300995);
nor I_76393 (I1300861,I1301125,I1301108);
nor I_76394 (I1301232,I1341607,I1341625);
not I_76395 (I1301249,I1301232);
DFFARX1 I_76396 (I1301232,I2507,I1300893,I1301275,);
not I_76397 (I1300885,I1301275);
nor I_76398 (I1301297,I1341607,I1341607);
DFFARX1 I_76399 (I1301297,I2507,I1300893,I1301323,);
and I_76400 (I1301331,I1301323,I1341619);
nor I_76401 (I1301348,I1301331,I1301249);
DFFARX1 I_76402 (I1301348,I2507,I1300893,I1300876,);
nor I_76403 (I1301379,I1301323,I1301108);
DFFARX1 I_76404 (I1301379,I2507,I1300893,I1300858,);
nor I_76405 (I1300873,I1301323,I1301012);
not I_76406 (I1301454,I2514);
DFFARX1 I_76407 (I1152587,I2507,I1301454,I1301480,);
nand I_76408 (I1301488,I1301480,I1152584);
not I_76409 (I1301505,I1301488);
DFFARX1 I_76410 (I1152587,I2507,I1301454,I1301531,);
not I_76411 (I1301539,I1301531);
nor I_76412 (I1301556,I1152605,I1152599);
not I_76413 (I1301573,I1301556);
DFFARX1 I_76414 (I1301573,I2507,I1301454,I1301440,);
or I_76415 (I1301604,I1152608,I1152605);
DFFARX1 I_76416 (I1301604,I2507,I1301454,I1301443,);
not I_76417 (I1301635,I1152596);
nor I_76418 (I1301652,I1301635,I1152593);
nor I_76419 (I1301669,I1301652,I1152599);
nor I_76420 (I1301686,I1152593,I1152584);
nor I_76421 (I1301703,I1301539,I1301686);
nor I_76422 (I1301428,I1301505,I1301703);
not I_76423 (I1301734,I1301686);
nand I_76424 (I1301431,I1301734,I1301488);
nand I_76425 (I1301425,I1301734,I1301556);
nor I_76426 (I1301422,I1301686,I1301669);
nor I_76427 (I1301793,I1152590,I1152608);
not I_76428 (I1301810,I1301793);
DFFARX1 I_76429 (I1301793,I2507,I1301454,I1301836,);
not I_76430 (I1301446,I1301836);
nor I_76431 (I1301858,I1152590,I1152602);
DFFARX1 I_76432 (I1301858,I2507,I1301454,I1301884,);
and I_76433 (I1301892,I1301884,I1152605);
nor I_76434 (I1301909,I1301892,I1301810);
DFFARX1 I_76435 (I1301909,I2507,I1301454,I1301437,);
nor I_76436 (I1301940,I1301884,I1301669);
DFFARX1 I_76437 (I1301940,I2507,I1301454,I1301419,);
nor I_76438 (I1301434,I1301884,I1301573);
not I_76439 (I1302015,I2514);
DFFARX1 I_76440 (I1205185,I2507,I1302015,I1302041,);
nand I_76441 (I1302049,I1302041,I1205182);
not I_76442 (I1302066,I1302049);
DFFARX1 I_76443 (I1205185,I2507,I1302015,I1302092,);
not I_76444 (I1302100,I1302092);
nor I_76445 (I1302117,I1205203,I1205197);
not I_76446 (I1302134,I1302117);
DFFARX1 I_76447 (I1302134,I2507,I1302015,I1302001,);
or I_76448 (I1302165,I1205206,I1205203);
DFFARX1 I_76449 (I1302165,I2507,I1302015,I1302004,);
not I_76450 (I1302196,I1205194);
nor I_76451 (I1302213,I1302196,I1205191);
nor I_76452 (I1302230,I1302213,I1205197);
nor I_76453 (I1302247,I1205191,I1205182);
nor I_76454 (I1302264,I1302100,I1302247);
nor I_76455 (I1301989,I1302066,I1302264);
not I_76456 (I1302295,I1302247);
nand I_76457 (I1301992,I1302295,I1302049);
nand I_76458 (I1301986,I1302295,I1302117);
nor I_76459 (I1301983,I1302247,I1302230);
nor I_76460 (I1302354,I1205188,I1205206);
not I_76461 (I1302371,I1302354);
DFFARX1 I_76462 (I1302354,I2507,I1302015,I1302397,);
not I_76463 (I1302007,I1302397);
nor I_76464 (I1302419,I1205188,I1205200);
DFFARX1 I_76465 (I1302419,I2507,I1302015,I1302445,);
and I_76466 (I1302453,I1302445,I1205203);
nor I_76467 (I1302470,I1302453,I1302371);
DFFARX1 I_76468 (I1302470,I2507,I1302015,I1301998,);
nor I_76469 (I1302501,I1302445,I1302230);
DFFARX1 I_76470 (I1302501,I2507,I1302015,I1301980,);
nor I_76471 (I1301995,I1302445,I1302134);
not I_76472 (I1302576,I2514);
DFFARX1 I_76473 (I724372,I2507,I1302576,I1302602,);
nand I_76474 (I1302610,I1302602,I724357);
not I_76475 (I1302627,I1302610);
DFFARX1 I_76476 (I724375,I2507,I1302576,I1302653,);
not I_76477 (I1302661,I1302653);
nor I_76478 (I1302678,I724354,I724369);
not I_76479 (I1302695,I1302678);
DFFARX1 I_76480 (I1302695,I2507,I1302576,I1302562,);
or I_76481 (I1302726,I724366,I724354);
DFFARX1 I_76482 (I1302726,I2507,I1302576,I1302565,);
not I_76483 (I1302757,I724354);
nor I_76484 (I1302774,I1302757,I724363);
nor I_76485 (I1302791,I1302774,I724369);
nor I_76486 (I1302808,I724363,I724357);
nor I_76487 (I1302825,I1302661,I1302808);
nor I_76488 (I1302550,I1302627,I1302825);
not I_76489 (I1302856,I1302808);
nand I_76490 (I1302553,I1302856,I1302610);
nand I_76491 (I1302547,I1302856,I1302678);
nor I_76492 (I1302544,I1302808,I1302791);
nor I_76493 (I1302915,I724360,I724366);
not I_76494 (I1302932,I1302915);
DFFARX1 I_76495 (I1302915,I2507,I1302576,I1302958,);
not I_76496 (I1302568,I1302958);
nor I_76497 (I1302980,I724360,I724378);
DFFARX1 I_76498 (I1302980,I2507,I1302576,I1303006,);
and I_76499 (I1303014,I1303006,I724354);
nor I_76500 (I1303031,I1303014,I1302932);
DFFARX1 I_76501 (I1303031,I2507,I1302576,I1302559,);
nor I_76502 (I1303062,I1303006,I1302791);
DFFARX1 I_76503 (I1303062,I2507,I1302576,I1302541,);
nor I_76504 (I1302556,I1303006,I1302695);
not I_76505 (I1303137,I2514);
DFFARX1 I_76506 (I676398,I2507,I1303137,I1303163,);
nand I_76507 (I1303171,I1303163,I676383);
not I_76508 (I1303188,I1303171);
DFFARX1 I_76509 (I676401,I2507,I1303137,I1303214,);
not I_76510 (I1303222,I1303214);
nor I_76511 (I1303239,I676380,I676395);
not I_76512 (I1303256,I1303239);
DFFARX1 I_76513 (I1303256,I2507,I1303137,I1303123,);
or I_76514 (I1303287,I676392,I676380);
DFFARX1 I_76515 (I1303287,I2507,I1303137,I1303126,);
not I_76516 (I1303318,I676380);
nor I_76517 (I1303335,I1303318,I676389);
nor I_76518 (I1303352,I1303335,I676395);
nor I_76519 (I1303369,I676389,I676383);
nor I_76520 (I1303386,I1303222,I1303369);
nor I_76521 (I1303111,I1303188,I1303386);
not I_76522 (I1303417,I1303369);
nand I_76523 (I1303114,I1303417,I1303171);
nand I_76524 (I1303108,I1303417,I1303239);
nor I_76525 (I1303105,I1303369,I1303352);
nor I_76526 (I1303476,I676386,I676392);
not I_76527 (I1303493,I1303476);
DFFARX1 I_76528 (I1303476,I2507,I1303137,I1303519,);
not I_76529 (I1303129,I1303519);
nor I_76530 (I1303541,I676386,I676404);
DFFARX1 I_76531 (I1303541,I2507,I1303137,I1303567,);
and I_76532 (I1303575,I1303567,I676380);
nor I_76533 (I1303592,I1303575,I1303493);
DFFARX1 I_76534 (I1303592,I2507,I1303137,I1303120,);
nor I_76535 (I1303623,I1303567,I1303352);
DFFARX1 I_76536 (I1303623,I2507,I1303137,I1303102,);
nor I_76537 (I1303117,I1303567,I1303256);
not I_76538 (I1303698,I2514);
DFFARX1 I_76539 (I1339837,I2507,I1303698,I1303724,);
nand I_76540 (I1303732,I1303724,I1339831);
not I_76541 (I1303749,I1303732);
DFFARX1 I_76542 (I1339849,I2507,I1303698,I1303775,);
not I_76543 (I1303783,I1303775);
nor I_76544 (I1303800,I1339834,I1339825);
not I_76545 (I1303817,I1303800);
DFFARX1 I_76546 (I1303817,I2507,I1303698,I1303684,);
or I_76547 (I1303848,I1339840,I1339834);
DFFARX1 I_76548 (I1303848,I2507,I1303698,I1303687,);
not I_76549 (I1303879,I1339843);
nor I_76550 (I1303896,I1303879,I1339846);
nor I_76551 (I1303913,I1303896,I1339825);
nor I_76552 (I1303930,I1339846,I1339828);
nor I_76553 (I1303947,I1303783,I1303930);
nor I_76554 (I1303672,I1303749,I1303947);
not I_76555 (I1303978,I1303930);
nand I_76556 (I1303675,I1303978,I1303732);
nand I_76557 (I1303669,I1303978,I1303800);
nor I_76558 (I1303666,I1303930,I1303913);
nor I_76559 (I1304037,I1339822,I1339840);
not I_76560 (I1304054,I1304037);
DFFARX1 I_76561 (I1304037,I2507,I1303698,I1304080,);
not I_76562 (I1303690,I1304080);
nor I_76563 (I1304102,I1339822,I1339822);
DFFARX1 I_76564 (I1304102,I2507,I1303698,I1304128,);
and I_76565 (I1304136,I1304128,I1339834);
nor I_76566 (I1304153,I1304136,I1304054);
DFFARX1 I_76567 (I1304153,I2507,I1303698,I1303681,);
nor I_76568 (I1304184,I1304128,I1303913);
DFFARX1 I_76569 (I1304184,I2507,I1303698,I1303663,);
nor I_76570 (I1303678,I1304128,I1303817);
not I_76571 (I1304259,I2514);
DFFARX1 I_76572 (I415332,I2507,I1304259,I1304285,);
nand I_76573 (I1304293,I1304285,I415314);
not I_76574 (I1304310,I1304293);
DFFARX1 I_76575 (I415311,I2507,I1304259,I1304336,);
not I_76576 (I1304344,I1304336);
nor I_76577 (I1304361,I415317,I415311);
not I_76578 (I1304378,I1304361);
DFFARX1 I_76579 (I1304378,I2507,I1304259,I1304245,);
or I_76580 (I1304409,I415320,I415317);
DFFARX1 I_76581 (I1304409,I2507,I1304259,I1304248,);
not I_76582 (I1304440,I415326);
nor I_76583 (I1304457,I1304440,I415338);
nor I_76584 (I1304474,I1304457,I415311);
nor I_76585 (I1304491,I415338,I415323);
nor I_76586 (I1304508,I1304344,I1304491);
nor I_76587 (I1304233,I1304310,I1304508);
not I_76588 (I1304539,I1304491);
nand I_76589 (I1304236,I1304539,I1304293);
nand I_76590 (I1304230,I1304539,I1304361);
nor I_76591 (I1304227,I1304491,I1304474);
nor I_76592 (I1304598,I415329,I415320);
not I_76593 (I1304615,I1304598);
DFFARX1 I_76594 (I1304598,I2507,I1304259,I1304641,);
not I_76595 (I1304251,I1304641);
nor I_76596 (I1304663,I415329,I415335);
DFFARX1 I_76597 (I1304663,I2507,I1304259,I1304689,);
and I_76598 (I1304697,I1304689,I415317);
nor I_76599 (I1304714,I1304697,I1304615);
DFFARX1 I_76600 (I1304714,I2507,I1304259,I1304242,);
nor I_76601 (I1304745,I1304689,I1304474);
DFFARX1 I_76602 (I1304745,I2507,I1304259,I1304224,);
nor I_76603 (I1304239,I1304689,I1304378);
not I_76604 (I1304820,I2514);
DFFARX1 I_76605 (I1147963,I2507,I1304820,I1304846,);
nand I_76606 (I1304854,I1304846,I1147960);
not I_76607 (I1304871,I1304854);
DFFARX1 I_76608 (I1147963,I2507,I1304820,I1304897,);
not I_76609 (I1304905,I1304897);
nor I_76610 (I1304922,I1147981,I1147975);
not I_76611 (I1304939,I1304922);
DFFARX1 I_76612 (I1304939,I2507,I1304820,I1304806,);
or I_76613 (I1304970,I1147984,I1147981);
DFFARX1 I_76614 (I1304970,I2507,I1304820,I1304809,);
not I_76615 (I1305001,I1147972);
nor I_76616 (I1305018,I1305001,I1147969);
nor I_76617 (I1305035,I1305018,I1147975);
nor I_76618 (I1305052,I1147969,I1147960);
nor I_76619 (I1305069,I1304905,I1305052);
nor I_76620 (I1304794,I1304871,I1305069);
not I_76621 (I1305100,I1305052);
nand I_76622 (I1304797,I1305100,I1304854);
nand I_76623 (I1304791,I1305100,I1304922);
nor I_76624 (I1304788,I1305052,I1305035);
nor I_76625 (I1305159,I1147966,I1147984);
not I_76626 (I1305176,I1305159);
DFFARX1 I_76627 (I1305159,I2507,I1304820,I1305202,);
not I_76628 (I1304812,I1305202);
nor I_76629 (I1305224,I1147966,I1147978);
DFFARX1 I_76630 (I1305224,I2507,I1304820,I1305250,);
and I_76631 (I1305258,I1305250,I1147981);
nor I_76632 (I1305275,I1305258,I1305176);
DFFARX1 I_76633 (I1305275,I2507,I1304820,I1304803,);
nor I_76634 (I1305306,I1305250,I1305035);
DFFARX1 I_76635 (I1305306,I2507,I1304820,I1304785,);
nor I_76636 (I1304800,I1305250,I1304939);
not I_76637 (I1305381,I2514);
DFFARX1 I_76638 (I848627,I2507,I1305381,I1305407,);
nand I_76639 (I1305415,I1305407,I848645);
not I_76640 (I1305432,I1305415);
DFFARX1 I_76641 (I848624,I2507,I1305381,I1305458,);
not I_76642 (I1305466,I1305458);
nor I_76643 (I1305483,I848639,I848633);
not I_76644 (I1305500,I1305483);
DFFARX1 I_76645 (I1305500,I2507,I1305381,I1305367,);
or I_76646 (I1305531,I848630,I848639);
DFFARX1 I_76647 (I1305531,I2507,I1305381,I1305370,);
not I_76648 (I1305562,I848630);
nor I_76649 (I1305579,I1305562,I848636);
nor I_76650 (I1305596,I1305579,I848633);
nor I_76651 (I1305613,I848636,I848624);
nor I_76652 (I1305630,I1305466,I1305613);
nor I_76653 (I1305355,I1305432,I1305630);
not I_76654 (I1305661,I1305613);
nand I_76655 (I1305358,I1305661,I1305415);
nand I_76656 (I1305352,I1305661,I1305483);
nor I_76657 (I1305349,I1305613,I1305596);
nor I_76658 (I1305720,I848627,I848630);
not I_76659 (I1305737,I1305720);
DFFARX1 I_76660 (I1305720,I2507,I1305381,I1305763,);
not I_76661 (I1305373,I1305763);
nor I_76662 (I1305785,I848627,I848642);
DFFARX1 I_76663 (I1305785,I2507,I1305381,I1305811,);
and I_76664 (I1305819,I1305811,I848639);
nor I_76665 (I1305836,I1305819,I1305737);
DFFARX1 I_76666 (I1305836,I2507,I1305381,I1305364,);
nor I_76667 (I1305867,I1305811,I1305596);
DFFARX1 I_76668 (I1305867,I2507,I1305381,I1305346,);
nor I_76669 (I1305361,I1305811,I1305500);
not I_76670 (I1305942,I2514);
DFFARX1 I_76671 (I274453,I2507,I1305942,I1305968,);
DFFARX1 I_76672 (I274447,I2507,I1305942,I1305985,);
not I_76673 (I1305993,I1305985);
nor I_76674 (I1305910,I1305968,I1305993);
DFFARX1 I_76675 (I1305993,I2507,I1305942,I1305925,);
nor I_76676 (I1306038,I274435,I274456);
and I_76677 (I1306055,I1306038,I274450);
nor I_76678 (I1306072,I1306055,I274435);
not I_76679 (I1306089,I274435);
and I_76680 (I1306106,I1306089,I274432);
nand I_76681 (I1306123,I1306106,I274444);
nor I_76682 (I1306140,I1306089,I1306123);
DFFARX1 I_76683 (I1306140,I2507,I1305942,I1305907,);
not I_76684 (I1306171,I1306123);
nand I_76685 (I1306188,I1305993,I1306171);
nand I_76686 (I1305919,I1306055,I1306171);
DFFARX1 I_76687 (I1306089,I2507,I1305942,I1305934,);
not I_76688 (I1306233,I274459);
nor I_76689 (I1306250,I1306233,I274432);
nor I_76690 (I1306267,I1306250,I1306072);
DFFARX1 I_76691 (I1306267,I2507,I1305942,I1305931,);
not I_76692 (I1306298,I1306250);
DFFARX1 I_76693 (I1306298,I2507,I1305942,I1306324,);
not I_76694 (I1306332,I1306324);
nor I_76695 (I1305928,I1306332,I1306250);
nor I_76696 (I1306363,I1306233,I274441);
and I_76697 (I1306380,I1306363,I274438);
or I_76698 (I1306397,I1306380,I274432);
DFFARX1 I_76699 (I1306397,I2507,I1305942,I1306423,);
not I_76700 (I1306431,I1306423);
nand I_76701 (I1306448,I1306431,I1306171);
not I_76702 (I1305922,I1306448);
nand I_76703 (I1305916,I1306448,I1306188);
nand I_76704 (I1305913,I1306431,I1306055);
not I_76705 (I1306537,I2514);
DFFARX1 I_76706 (I970911,I2507,I1306537,I1306563,);
DFFARX1 I_76707 (I970929,I2507,I1306537,I1306580,);
not I_76708 (I1306588,I1306580);
nor I_76709 (I1306505,I1306563,I1306588);
DFFARX1 I_76710 (I1306588,I2507,I1306537,I1306520,);
nor I_76711 (I1306633,I970908,I970920);
and I_76712 (I1306650,I1306633,I970905);
nor I_76713 (I1306667,I1306650,I970908);
not I_76714 (I1306684,I970908);
and I_76715 (I1306701,I1306684,I970914);
nand I_76716 (I1306718,I1306701,I970926);
nor I_76717 (I1306735,I1306684,I1306718);
DFFARX1 I_76718 (I1306735,I2507,I1306537,I1306502,);
not I_76719 (I1306766,I1306718);
nand I_76720 (I1306783,I1306588,I1306766);
nand I_76721 (I1306514,I1306650,I1306766);
DFFARX1 I_76722 (I1306684,I2507,I1306537,I1306529,);
not I_76723 (I1306828,I970917);
nor I_76724 (I1306845,I1306828,I970914);
nor I_76725 (I1306862,I1306845,I1306667);
DFFARX1 I_76726 (I1306862,I2507,I1306537,I1306526,);
not I_76727 (I1306893,I1306845);
DFFARX1 I_76728 (I1306893,I2507,I1306537,I1306919,);
not I_76729 (I1306927,I1306919);
nor I_76730 (I1306523,I1306927,I1306845);
nor I_76731 (I1306958,I1306828,I970905);
and I_76732 (I1306975,I1306958,I970932);
or I_76733 (I1306992,I1306975,I970923);
DFFARX1 I_76734 (I1306992,I2507,I1306537,I1307018,);
not I_76735 (I1307026,I1307018);
nand I_76736 (I1307043,I1307026,I1306766);
not I_76737 (I1306517,I1307043);
nand I_76738 (I1306511,I1307043,I1306783);
nand I_76739 (I1306508,I1307026,I1306650);
not I_76740 (I1307132,I2514);
DFFARX1 I_76741 (I422383,I2507,I1307132,I1307158,);
DFFARX1 I_76742 (I422389,I2507,I1307132,I1307175,);
not I_76743 (I1307183,I1307175);
nor I_76744 (I1307100,I1307158,I1307183);
DFFARX1 I_76745 (I1307183,I2507,I1307132,I1307115,);
nor I_76746 (I1307228,I422398,I422383);
and I_76747 (I1307245,I1307228,I422410);
nor I_76748 (I1307262,I1307245,I422398);
not I_76749 (I1307279,I422398);
and I_76750 (I1307296,I1307279,I422386);
nand I_76751 (I1307313,I1307296,I422407);
nor I_76752 (I1307330,I1307279,I1307313);
DFFARX1 I_76753 (I1307330,I2507,I1307132,I1307097,);
not I_76754 (I1307361,I1307313);
nand I_76755 (I1307378,I1307183,I1307361);
nand I_76756 (I1307109,I1307245,I1307361);
DFFARX1 I_76757 (I1307279,I2507,I1307132,I1307124,);
not I_76758 (I1307423,I422395);
nor I_76759 (I1307440,I1307423,I422386);
nor I_76760 (I1307457,I1307440,I1307262);
DFFARX1 I_76761 (I1307457,I2507,I1307132,I1307121,);
not I_76762 (I1307488,I1307440);
DFFARX1 I_76763 (I1307488,I2507,I1307132,I1307514,);
not I_76764 (I1307522,I1307514);
nor I_76765 (I1307118,I1307522,I1307440);
nor I_76766 (I1307553,I1307423,I422392);
and I_76767 (I1307570,I1307553,I422404);
or I_76768 (I1307587,I1307570,I422401);
DFFARX1 I_76769 (I1307587,I2507,I1307132,I1307613,);
not I_76770 (I1307621,I1307613);
nand I_76771 (I1307638,I1307621,I1307361);
not I_76772 (I1307112,I1307638);
nand I_76773 (I1307106,I1307638,I1307378);
nand I_76774 (I1307103,I1307621,I1307245);
not I_76775 (I1307727,I2514);
DFFARX1 I_76776 (I1211234,I2507,I1307727,I1307753,);
DFFARX1 I_76777 (I1211237,I2507,I1307727,I1307770,);
not I_76778 (I1307778,I1307770);
nor I_76779 (I1307695,I1307753,I1307778);
DFFARX1 I_76780 (I1307778,I2507,I1307727,I1307710,);
nor I_76781 (I1307823,I1211237,I1211252);
and I_76782 (I1307840,I1307823,I1211246);
nor I_76783 (I1307857,I1307840,I1211237);
not I_76784 (I1307874,I1211237);
and I_76785 (I1307891,I1307874,I1211255);
nand I_76786 (I1307908,I1307891,I1211243);
nor I_76787 (I1307925,I1307874,I1307908);
DFFARX1 I_76788 (I1307925,I2507,I1307727,I1307692,);
not I_76789 (I1307956,I1307908);
nand I_76790 (I1307973,I1307778,I1307956);
nand I_76791 (I1307704,I1307840,I1307956);
DFFARX1 I_76792 (I1307874,I2507,I1307727,I1307719,);
not I_76793 (I1308018,I1211249);
nor I_76794 (I1308035,I1308018,I1211255);
nor I_76795 (I1308052,I1308035,I1307857);
DFFARX1 I_76796 (I1308052,I2507,I1307727,I1307716,);
not I_76797 (I1308083,I1308035);
DFFARX1 I_76798 (I1308083,I2507,I1307727,I1308109,);
not I_76799 (I1308117,I1308109);
nor I_76800 (I1307713,I1308117,I1308035);
nor I_76801 (I1308148,I1308018,I1211234);
and I_76802 (I1308165,I1308148,I1211258);
or I_76803 (I1308182,I1308165,I1211240);
DFFARX1 I_76804 (I1308182,I2507,I1307727,I1308208,);
not I_76805 (I1308216,I1308208);
nand I_76806 (I1308233,I1308216,I1307956);
not I_76807 (I1307707,I1308233);
nand I_76808 (I1307701,I1308233,I1307973);
nand I_76809 (I1307698,I1308216,I1307840);
not I_76810 (I1308322,I2514);
DFFARX1 I_76811 (I124445,I2507,I1308322,I1308348,);
DFFARX1 I_76812 (I124433,I2507,I1308322,I1308365,);
not I_76813 (I1308373,I1308365);
nor I_76814 (I1308290,I1308348,I1308373);
DFFARX1 I_76815 (I1308373,I2507,I1308322,I1308305,);
nor I_76816 (I1308418,I124424,I124448);
and I_76817 (I1308435,I1308418,I124427);
nor I_76818 (I1308452,I1308435,I124424);
not I_76819 (I1308469,I124424);
and I_76820 (I1308486,I1308469,I124430);
nand I_76821 (I1308503,I1308486,I124442);
nor I_76822 (I1308520,I1308469,I1308503);
DFFARX1 I_76823 (I1308520,I2507,I1308322,I1308287,);
not I_76824 (I1308551,I1308503);
nand I_76825 (I1308568,I1308373,I1308551);
nand I_76826 (I1308299,I1308435,I1308551);
DFFARX1 I_76827 (I1308469,I2507,I1308322,I1308314,);
not I_76828 (I1308613,I124424);
nor I_76829 (I1308630,I1308613,I124430);
nor I_76830 (I1308647,I1308630,I1308452);
DFFARX1 I_76831 (I1308647,I2507,I1308322,I1308311,);
not I_76832 (I1308678,I1308630);
DFFARX1 I_76833 (I1308678,I2507,I1308322,I1308704,);
not I_76834 (I1308712,I1308704);
nor I_76835 (I1308308,I1308712,I1308630);
nor I_76836 (I1308743,I1308613,I124427);
and I_76837 (I1308760,I1308743,I124436);
or I_76838 (I1308777,I1308760,I124439);
DFFARX1 I_76839 (I1308777,I2507,I1308322,I1308803,);
not I_76840 (I1308811,I1308803);
nand I_76841 (I1308828,I1308811,I1308551);
not I_76842 (I1308302,I1308828);
nand I_76843 (I1308296,I1308828,I1308568);
nand I_76844 (I1308293,I1308811,I1308435);
not I_76845 (I1308917,I2514);
DFFARX1 I_76846 (I803311,I2507,I1308917,I1308943,);
DFFARX1 I_76847 (I803308,I2507,I1308917,I1308960,);
not I_76848 (I1308968,I1308960);
nor I_76849 (I1308885,I1308943,I1308968);
DFFARX1 I_76850 (I1308968,I2507,I1308917,I1308900,);
nor I_76851 (I1309013,I803323,I803305);
and I_76852 (I1309030,I1309013,I803302);
nor I_76853 (I1309047,I1309030,I803323);
not I_76854 (I1309064,I803323);
and I_76855 (I1309081,I1309064,I803308);
nand I_76856 (I1309098,I1309081,I803320);
nor I_76857 (I1309115,I1309064,I1309098);
DFFARX1 I_76858 (I1309115,I2507,I1308917,I1308882,);
not I_76859 (I1309146,I1309098);
nand I_76860 (I1309163,I1308968,I1309146);
nand I_76861 (I1308894,I1309030,I1309146);
DFFARX1 I_76862 (I1309064,I2507,I1308917,I1308909,);
not I_76863 (I1309208,I803314);
nor I_76864 (I1309225,I1309208,I803308);
nor I_76865 (I1309242,I1309225,I1309047);
DFFARX1 I_76866 (I1309242,I2507,I1308917,I1308906,);
not I_76867 (I1309273,I1309225);
DFFARX1 I_76868 (I1309273,I2507,I1308917,I1309299,);
not I_76869 (I1309307,I1309299);
nor I_76870 (I1308903,I1309307,I1309225);
nor I_76871 (I1309338,I1309208,I803302);
and I_76872 (I1309355,I1309338,I803317);
or I_76873 (I1309372,I1309355,I803305);
DFFARX1 I_76874 (I1309372,I2507,I1308917,I1309398,);
not I_76875 (I1309406,I1309398);
nand I_76876 (I1309423,I1309406,I1309146);
not I_76877 (I1308897,I1309423);
nand I_76878 (I1308891,I1309423,I1309163);
nand I_76879 (I1308888,I1309406,I1309030);
not I_76880 (I1309512,I2514);
DFFARX1 I_76881 (I43811,I2507,I1309512,I1309538,);
DFFARX1 I_76882 (I43793,I2507,I1309512,I1309555,);
not I_76883 (I1309563,I1309555);
nor I_76884 (I1309480,I1309538,I1309563);
DFFARX1 I_76885 (I1309563,I2507,I1309512,I1309495,);
nor I_76886 (I1309608,I43793,I43808);
and I_76887 (I1309625,I1309608,I43802);
nor I_76888 (I1309642,I1309625,I43793);
not I_76889 (I1309659,I43793);
and I_76890 (I1309676,I1309659,I43796);
nand I_76891 (I1309693,I1309676,I43799);
nor I_76892 (I1309710,I1309659,I1309693);
DFFARX1 I_76893 (I1309710,I2507,I1309512,I1309477,);
not I_76894 (I1309741,I1309693);
nand I_76895 (I1309758,I1309563,I1309741);
nand I_76896 (I1309489,I1309625,I1309741);
DFFARX1 I_76897 (I1309659,I2507,I1309512,I1309504,);
not I_76898 (I1309803,I43805);
nor I_76899 (I1309820,I1309803,I43796);
nor I_76900 (I1309837,I1309820,I1309642);
DFFARX1 I_76901 (I1309837,I2507,I1309512,I1309501,);
not I_76902 (I1309868,I1309820);
DFFARX1 I_76903 (I1309868,I2507,I1309512,I1309894,);
not I_76904 (I1309902,I1309894);
nor I_76905 (I1309498,I1309902,I1309820);
nor I_76906 (I1309933,I1309803,I43817);
and I_76907 (I1309950,I1309933,I43814);
or I_76908 (I1309967,I1309950,I43796);
DFFARX1 I_76909 (I1309967,I2507,I1309512,I1309993,);
not I_76910 (I1310001,I1309993);
nand I_76911 (I1310018,I1310001,I1309741);
not I_76912 (I1309492,I1310018);
nand I_76913 (I1309486,I1310018,I1309758);
nand I_76914 (I1309483,I1310001,I1309625);
not I_76915 (I1310107,I2514);
DFFARX1 I_76916 (I1270956,I2507,I1310107,I1310133,);
DFFARX1 I_76917 (I1270947,I2507,I1310107,I1310150,);
not I_76918 (I1310158,I1310150);
nor I_76919 (I1310075,I1310133,I1310158);
DFFARX1 I_76920 (I1310158,I2507,I1310107,I1310090,);
nor I_76921 (I1310203,I1270938,I1270953);
and I_76922 (I1310220,I1310203,I1270941);
nor I_76923 (I1310237,I1310220,I1270938);
not I_76924 (I1310254,I1270938);
and I_76925 (I1310271,I1310254,I1270944);
nand I_76926 (I1310288,I1310271,I1270962);
nor I_76927 (I1310305,I1310254,I1310288);
DFFARX1 I_76928 (I1310305,I2507,I1310107,I1310072,);
not I_76929 (I1310336,I1310288);
nand I_76930 (I1310353,I1310158,I1310336);
nand I_76931 (I1310084,I1310220,I1310336);
DFFARX1 I_76932 (I1310254,I2507,I1310107,I1310099,);
not I_76933 (I1310398,I1270938);
nor I_76934 (I1310415,I1310398,I1270944);
nor I_76935 (I1310432,I1310415,I1310237);
DFFARX1 I_76936 (I1310432,I2507,I1310107,I1310096,);
not I_76937 (I1310463,I1310415);
DFFARX1 I_76938 (I1310463,I2507,I1310107,I1310489,);
not I_76939 (I1310497,I1310489);
nor I_76940 (I1310093,I1310497,I1310415);
nor I_76941 (I1310528,I1310398,I1270941);
and I_76942 (I1310545,I1310528,I1270950);
or I_76943 (I1310562,I1310545,I1270959);
DFFARX1 I_76944 (I1310562,I2507,I1310107,I1310588,);
not I_76945 (I1310596,I1310588);
nand I_76946 (I1310613,I1310596,I1310336);
not I_76947 (I1310087,I1310613);
nand I_76948 (I1310081,I1310613,I1310353);
nand I_76949 (I1310078,I1310596,I1310220);
not I_76950 (I1310702,I2514);
DFFARX1 I_76951 (I867605,I2507,I1310702,I1310728,);
DFFARX1 I_76952 (I867602,I2507,I1310702,I1310745,);
not I_76953 (I1310753,I1310745);
nor I_76954 (I1310670,I1310728,I1310753);
DFFARX1 I_76955 (I1310753,I2507,I1310702,I1310685,);
nor I_76956 (I1310798,I867617,I867599);
and I_76957 (I1310815,I1310798,I867596);
nor I_76958 (I1310832,I1310815,I867617);
not I_76959 (I1310849,I867617);
and I_76960 (I1310866,I1310849,I867602);
nand I_76961 (I1310883,I1310866,I867614);
nor I_76962 (I1310900,I1310849,I1310883);
DFFARX1 I_76963 (I1310900,I2507,I1310702,I1310667,);
not I_76964 (I1310931,I1310883);
nand I_76965 (I1310948,I1310753,I1310931);
nand I_76966 (I1310679,I1310815,I1310931);
DFFARX1 I_76967 (I1310849,I2507,I1310702,I1310694,);
not I_76968 (I1310993,I867608);
nor I_76969 (I1311010,I1310993,I867602);
nor I_76970 (I1311027,I1311010,I1310832);
DFFARX1 I_76971 (I1311027,I2507,I1310702,I1310691,);
not I_76972 (I1311058,I1311010);
DFFARX1 I_76973 (I1311058,I2507,I1310702,I1311084,);
not I_76974 (I1311092,I1311084);
nor I_76975 (I1310688,I1311092,I1311010);
nor I_76976 (I1311123,I1310993,I867596);
and I_76977 (I1311140,I1311123,I867611);
or I_76978 (I1311157,I1311140,I867599);
DFFARX1 I_76979 (I1311157,I2507,I1310702,I1311183,);
not I_76980 (I1311191,I1311183);
nand I_76981 (I1311208,I1311191,I1310931);
not I_76982 (I1310682,I1311208);
nand I_76983 (I1310676,I1311208,I1310948);
nand I_76984 (I1310673,I1311191,I1310815);
not I_76985 (I1311297,I2514);
DFFARX1 I_76986 (I354030,I2507,I1311297,I1311323,);
DFFARX1 I_76987 (I354024,I2507,I1311297,I1311340,);
not I_76988 (I1311348,I1311340);
nor I_76989 (I1311265,I1311323,I1311348);
DFFARX1 I_76990 (I1311348,I2507,I1311297,I1311280,);
nor I_76991 (I1311393,I354012,I354033);
and I_76992 (I1311410,I1311393,I354027);
nor I_76993 (I1311427,I1311410,I354012);
not I_76994 (I1311444,I354012);
and I_76995 (I1311461,I1311444,I354009);
nand I_76996 (I1311478,I1311461,I354021);
nor I_76997 (I1311495,I1311444,I1311478);
DFFARX1 I_76998 (I1311495,I2507,I1311297,I1311262,);
not I_76999 (I1311526,I1311478);
nand I_77000 (I1311543,I1311348,I1311526);
nand I_77001 (I1311274,I1311410,I1311526);
DFFARX1 I_77002 (I1311444,I2507,I1311297,I1311289,);
not I_77003 (I1311588,I354036);
nor I_77004 (I1311605,I1311588,I354009);
nor I_77005 (I1311622,I1311605,I1311427);
DFFARX1 I_77006 (I1311622,I2507,I1311297,I1311286,);
not I_77007 (I1311653,I1311605);
DFFARX1 I_77008 (I1311653,I2507,I1311297,I1311679,);
not I_77009 (I1311687,I1311679);
nor I_77010 (I1311283,I1311687,I1311605);
nor I_77011 (I1311718,I1311588,I354018);
and I_77012 (I1311735,I1311718,I354015);
or I_77013 (I1311752,I1311735,I354009);
DFFARX1 I_77014 (I1311752,I2507,I1311297,I1311778,);
not I_77015 (I1311786,I1311778);
nand I_77016 (I1311803,I1311786,I1311526);
not I_77017 (I1311277,I1311803);
nand I_77018 (I1311271,I1311803,I1311543);
nand I_77019 (I1311268,I1311786,I1311410);
not I_77020 (I1311892,I2514);
DFFARX1 I_77021 (I1158945,I2507,I1311892,I1311918,);
DFFARX1 I_77022 (I1158957,I2507,I1311892,I1311935,);
not I_77023 (I1311943,I1311935);
nor I_77024 (I1311860,I1311918,I1311943);
DFFARX1 I_77025 (I1311943,I2507,I1311892,I1311875,);
nor I_77026 (I1311988,I1158954,I1158948);
and I_77027 (I1312005,I1311988,I1158942);
nor I_77028 (I1312022,I1312005,I1158954);
not I_77029 (I1312039,I1158954);
and I_77030 (I1312056,I1312039,I1158951);
nand I_77031 (I1312073,I1312056,I1158942);
nor I_77032 (I1312090,I1312039,I1312073);
DFFARX1 I_77033 (I1312090,I2507,I1311892,I1311857,);
not I_77034 (I1312121,I1312073);
nand I_77035 (I1312138,I1311943,I1312121);
nand I_77036 (I1311869,I1312005,I1312121);
DFFARX1 I_77037 (I1312039,I2507,I1311892,I1311884,);
not I_77038 (I1312183,I1158966);
nor I_77039 (I1312200,I1312183,I1158951);
nor I_77040 (I1312217,I1312200,I1312022);
DFFARX1 I_77041 (I1312217,I2507,I1311892,I1311881,);
not I_77042 (I1312248,I1312200);
DFFARX1 I_77043 (I1312248,I2507,I1311892,I1312274,);
not I_77044 (I1312282,I1312274);
nor I_77045 (I1311878,I1312282,I1312200);
nor I_77046 (I1312313,I1312183,I1158960);
and I_77047 (I1312330,I1312313,I1158963);
or I_77048 (I1312347,I1312330,I1158945);
DFFARX1 I_77049 (I1312347,I2507,I1311892,I1312373,);
not I_77050 (I1312381,I1312373);
nand I_77051 (I1312398,I1312381,I1312121);
not I_77052 (I1311872,I1312398);
nand I_77053 (I1311866,I1312398,I1312138);
nand I_77054 (I1311863,I1312381,I1312005);
not I_77055 (I1312487,I2514);
DFFARX1 I_77056 (I1009592,I2507,I1312487,I1312513,);
DFFARX1 I_77057 (I1009583,I2507,I1312487,I1312530,);
not I_77058 (I1312538,I1312530);
nor I_77059 (I1312455,I1312513,I1312538);
DFFARX1 I_77060 (I1312538,I2507,I1312487,I1312470,);
nor I_77061 (I1312583,I1009589,I1009598);
and I_77062 (I1312600,I1312583,I1009601);
nor I_77063 (I1312617,I1312600,I1009589);
not I_77064 (I1312634,I1009589);
and I_77065 (I1312651,I1312634,I1009580);
nand I_77066 (I1312668,I1312651,I1009586);
nor I_77067 (I1312685,I1312634,I1312668);
DFFARX1 I_77068 (I1312685,I2507,I1312487,I1312452,);
not I_77069 (I1312716,I1312668);
nand I_77070 (I1312733,I1312538,I1312716);
nand I_77071 (I1312464,I1312600,I1312716);
DFFARX1 I_77072 (I1312634,I2507,I1312487,I1312479,);
not I_77073 (I1312778,I1009595);
nor I_77074 (I1312795,I1312778,I1009580);
nor I_77075 (I1312812,I1312795,I1312617);
DFFARX1 I_77076 (I1312812,I2507,I1312487,I1312476,);
not I_77077 (I1312843,I1312795);
DFFARX1 I_77078 (I1312843,I2507,I1312487,I1312869,);
not I_77079 (I1312877,I1312869);
nor I_77080 (I1312473,I1312877,I1312795);
nor I_77081 (I1312908,I1312778,I1009580);
and I_77082 (I1312925,I1312908,I1009583);
or I_77083 (I1312942,I1312925,I1009586);
DFFARX1 I_77084 (I1312942,I2507,I1312487,I1312968,);
not I_77085 (I1312976,I1312968);
nand I_77086 (I1312993,I1312976,I1312716);
not I_77087 (I1312467,I1312993);
nand I_77088 (I1312461,I1312993,I1312733);
nand I_77089 (I1312458,I1312976,I1312600);
not I_77090 (I1313082,I2514);
DFFARX1 I_77091 (I666575,I2507,I1313082,I1313108,);
DFFARX1 I_77092 (I666557,I2507,I1313082,I1313125,);
not I_77093 (I1313133,I1313125);
nor I_77094 (I1313050,I1313108,I1313133);
DFFARX1 I_77095 (I1313133,I2507,I1313082,I1313065,);
nor I_77096 (I1313178,I666563,I666566);
and I_77097 (I1313195,I1313178,I666554);
nor I_77098 (I1313212,I1313195,I666563);
not I_77099 (I1313229,I666563);
and I_77100 (I1313246,I1313229,I666572);
nand I_77101 (I1313263,I1313246,I666560);
nor I_77102 (I1313280,I1313229,I1313263);
DFFARX1 I_77103 (I1313280,I2507,I1313082,I1313047,);
not I_77104 (I1313311,I1313263);
nand I_77105 (I1313328,I1313133,I1313311);
nand I_77106 (I1313059,I1313195,I1313311);
DFFARX1 I_77107 (I1313229,I2507,I1313082,I1313074,);
not I_77108 (I1313373,I666557);
nor I_77109 (I1313390,I1313373,I666572);
nor I_77110 (I1313407,I1313390,I1313212);
DFFARX1 I_77111 (I1313407,I2507,I1313082,I1313071,);
not I_77112 (I1313438,I1313390);
DFFARX1 I_77113 (I1313438,I2507,I1313082,I1313464,);
not I_77114 (I1313472,I1313464);
nor I_77115 (I1313068,I1313472,I1313390);
nor I_77116 (I1313503,I1313373,I666569);
and I_77117 (I1313520,I1313503,I666578);
or I_77118 (I1313537,I1313520,I666554);
DFFARX1 I_77119 (I1313537,I2507,I1313082,I1313563,);
not I_77120 (I1313571,I1313563);
nand I_77121 (I1313588,I1313571,I1313311);
not I_77122 (I1313062,I1313588);
nand I_77123 (I1313056,I1313588,I1313328);
nand I_77124 (I1313053,I1313571,I1313195);
not I_77125 (I1313677,I2514);
DFFARX1 I_77126 (I721485,I2507,I1313677,I1313703,);
DFFARX1 I_77127 (I721467,I2507,I1313677,I1313720,);
not I_77128 (I1313728,I1313720);
nor I_77129 (I1313645,I1313703,I1313728);
DFFARX1 I_77130 (I1313728,I2507,I1313677,I1313660,);
nor I_77131 (I1313773,I721473,I721476);
and I_77132 (I1313790,I1313773,I721464);
nor I_77133 (I1313807,I1313790,I721473);
not I_77134 (I1313824,I721473);
and I_77135 (I1313841,I1313824,I721482);
nand I_77136 (I1313858,I1313841,I721470);
nor I_77137 (I1313875,I1313824,I1313858);
DFFARX1 I_77138 (I1313875,I2507,I1313677,I1313642,);
not I_77139 (I1313906,I1313858);
nand I_77140 (I1313923,I1313728,I1313906);
nand I_77141 (I1313654,I1313790,I1313906);
DFFARX1 I_77142 (I1313824,I2507,I1313677,I1313669,);
not I_77143 (I1313968,I721467);
nor I_77144 (I1313985,I1313968,I721482);
nor I_77145 (I1314002,I1313985,I1313807);
DFFARX1 I_77146 (I1314002,I2507,I1313677,I1313666,);
not I_77147 (I1314033,I1313985);
DFFARX1 I_77148 (I1314033,I2507,I1313677,I1314059,);
not I_77149 (I1314067,I1314059);
nor I_77150 (I1313663,I1314067,I1313985);
nor I_77151 (I1314098,I1313968,I721479);
and I_77152 (I1314115,I1314098,I721488);
or I_77153 (I1314132,I1314115,I721464);
DFFARX1 I_77154 (I1314132,I2507,I1313677,I1314158,);
not I_77155 (I1314166,I1314158);
nand I_77156 (I1314183,I1314166,I1313906);
not I_77157 (I1313657,I1314183);
nand I_77158 (I1313651,I1314183,I1313923);
nand I_77159 (I1313648,I1314166,I1313790);
not I_77160 (I1314272,I2514);
DFFARX1 I_77161 (I109162,I2507,I1314272,I1314298,);
DFFARX1 I_77162 (I109150,I2507,I1314272,I1314315,);
not I_77163 (I1314323,I1314315);
nor I_77164 (I1314240,I1314298,I1314323);
DFFARX1 I_77165 (I1314323,I2507,I1314272,I1314255,);
nor I_77166 (I1314368,I109141,I109165);
and I_77167 (I1314385,I1314368,I109144);
nor I_77168 (I1314402,I1314385,I109141);
not I_77169 (I1314419,I109141);
and I_77170 (I1314436,I1314419,I109147);
nand I_77171 (I1314453,I1314436,I109159);
nor I_77172 (I1314470,I1314419,I1314453);
DFFARX1 I_77173 (I1314470,I2507,I1314272,I1314237,);
not I_77174 (I1314501,I1314453);
nand I_77175 (I1314518,I1314323,I1314501);
nand I_77176 (I1314249,I1314385,I1314501);
DFFARX1 I_77177 (I1314419,I2507,I1314272,I1314264,);
not I_77178 (I1314563,I109141);
nor I_77179 (I1314580,I1314563,I109147);
nor I_77180 (I1314597,I1314580,I1314402);
DFFARX1 I_77181 (I1314597,I2507,I1314272,I1314261,);
not I_77182 (I1314628,I1314580);
DFFARX1 I_77183 (I1314628,I2507,I1314272,I1314654,);
not I_77184 (I1314662,I1314654);
nor I_77185 (I1314258,I1314662,I1314580);
nor I_77186 (I1314693,I1314563,I109144);
and I_77187 (I1314710,I1314693,I109153);
or I_77188 (I1314727,I1314710,I109156);
DFFARX1 I_77189 (I1314727,I2507,I1314272,I1314753,);
not I_77190 (I1314761,I1314753);
nand I_77191 (I1314778,I1314761,I1314501);
not I_77192 (I1314252,I1314778);
nand I_77193 (I1314246,I1314778,I1314518);
nand I_77194 (I1314243,I1314761,I1314385);
not I_77195 (I1314867,I2514);
DFFARX1 I_77196 (I987707,I2507,I1314867,I1314893,);
DFFARX1 I_77197 (I987725,I2507,I1314867,I1314910,);
not I_77198 (I1314918,I1314910);
nor I_77199 (I1314835,I1314893,I1314918);
DFFARX1 I_77200 (I1314918,I2507,I1314867,I1314850,);
nor I_77201 (I1314963,I987704,I987716);
and I_77202 (I1314980,I1314963,I987701);
nor I_77203 (I1314997,I1314980,I987704);
not I_77204 (I1315014,I987704);
and I_77205 (I1315031,I1315014,I987710);
nand I_77206 (I1315048,I1315031,I987722);
nor I_77207 (I1315065,I1315014,I1315048);
DFFARX1 I_77208 (I1315065,I2507,I1314867,I1314832,);
not I_77209 (I1315096,I1315048);
nand I_77210 (I1315113,I1314918,I1315096);
nand I_77211 (I1314844,I1314980,I1315096);
DFFARX1 I_77212 (I1315014,I2507,I1314867,I1314859,);
not I_77213 (I1315158,I987713);
nor I_77214 (I1315175,I1315158,I987710);
nor I_77215 (I1315192,I1315175,I1314997);
DFFARX1 I_77216 (I1315192,I2507,I1314867,I1314856,);
not I_77217 (I1315223,I1315175);
DFFARX1 I_77218 (I1315223,I2507,I1314867,I1315249,);
not I_77219 (I1315257,I1315249);
nor I_77220 (I1314853,I1315257,I1315175);
nor I_77221 (I1315288,I1315158,I987701);
and I_77222 (I1315305,I1315288,I987728);
or I_77223 (I1315322,I1315305,I987719);
DFFARX1 I_77224 (I1315322,I2507,I1314867,I1315348,);
not I_77225 (I1315356,I1315348);
nand I_77226 (I1315373,I1315356,I1315096);
not I_77227 (I1314847,I1315373);
nand I_77228 (I1314841,I1315373,I1315113);
nand I_77229 (I1314838,I1315356,I1314980);
not I_77230 (I1315462,I2514);
DFFARX1 I_77231 (I193665,I2507,I1315462,I1315488,);
DFFARX1 I_77232 (I193668,I2507,I1315462,I1315505,);
not I_77233 (I1315513,I1315505);
nor I_77234 (I1315430,I1315488,I1315513);
DFFARX1 I_77235 (I1315513,I2507,I1315462,I1315445,);
nor I_77236 (I1315558,I193674,I193668);
and I_77237 (I1315575,I1315558,I193671);
nor I_77238 (I1315592,I1315575,I193674);
not I_77239 (I1315609,I193674);
and I_77240 (I1315626,I1315609,I193665);
nand I_77241 (I1315643,I1315626,I193683);
nor I_77242 (I1315660,I1315609,I1315643);
DFFARX1 I_77243 (I1315660,I2507,I1315462,I1315427,);
not I_77244 (I1315691,I1315643);
nand I_77245 (I1315708,I1315513,I1315691);
nand I_77246 (I1315439,I1315575,I1315691);
DFFARX1 I_77247 (I1315609,I2507,I1315462,I1315454,);
not I_77248 (I1315753,I193677);
nor I_77249 (I1315770,I1315753,I193665);
nor I_77250 (I1315787,I1315770,I1315592);
DFFARX1 I_77251 (I1315787,I2507,I1315462,I1315451,);
not I_77252 (I1315818,I1315770);
DFFARX1 I_77253 (I1315818,I2507,I1315462,I1315844,);
not I_77254 (I1315852,I1315844);
nor I_77255 (I1315448,I1315852,I1315770);
nor I_77256 (I1315883,I1315753,I193680);
and I_77257 (I1315900,I1315883,I193686);
or I_77258 (I1315917,I1315900,I193689);
DFFARX1 I_77259 (I1315917,I2507,I1315462,I1315943,);
not I_77260 (I1315951,I1315943);
nand I_77261 (I1315968,I1315951,I1315691);
not I_77262 (I1315442,I1315968);
nand I_77263 (I1315436,I1315968,I1315708);
nand I_77264 (I1315433,I1315951,I1315575);
not I_77265 (I1316057,I2514);
DFFARX1 I_77266 (I440879,I2507,I1316057,I1316083,);
DFFARX1 I_77267 (I440885,I2507,I1316057,I1316100,);
not I_77268 (I1316108,I1316100);
nor I_77269 (I1316025,I1316083,I1316108);
DFFARX1 I_77270 (I1316108,I2507,I1316057,I1316040,);
nor I_77271 (I1316153,I440894,I440879);
and I_77272 (I1316170,I1316153,I440906);
nor I_77273 (I1316187,I1316170,I440894);
not I_77274 (I1316204,I440894);
and I_77275 (I1316221,I1316204,I440882);
nand I_77276 (I1316238,I1316221,I440903);
nor I_77277 (I1316255,I1316204,I1316238);
DFFARX1 I_77278 (I1316255,I2507,I1316057,I1316022,);
not I_77279 (I1316286,I1316238);
nand I_77280 (I1316303,I1316108,I1316286);
nand I_77281 (I1316034,I1316170,I1316286);
DFFARX1 I_77282 (I1316204,I2507,I1316057,I1316049,);
not I_77283 (I1316348,I440891);
nor I_77284 (I1316365,I1316348,I440882);
nor I_77285 (I1316382,I1316365,I1316187);
DFFARX1 I_77286 (I1316382,I2507,I1316057,I1316046,);
not I_77287 (I1316413,I1316365);
DFFARX1 I_77288 (I1316413,I2507,I1316057,I1316439,);
not I_77289 (I1316447,I1316439);
nor I_77290 (I1316043,I1316447,I1316365);
nor I_77291 (I1316478,I1316348,I440888);
and I_77292 (I1316495,I1316478,I440900);
or I_77293 (I1316512,I1316495,I440897);
DFFARX1 I_77294 (I1316512,I2507,I1316057,I1316538,);
not I_77295 (I1316546,I1316538);
nand I_77296 (I1316563,I1316546,I1316286);
not I_77297 (I1316037,I1316563);
nand I_77298 (I1316031,I1316563,I1316303);
nand I_77299 (I1316028,I1316546,I1316170);
not I_77300 (I1316652,I2514);
DFFARX1 I_77301 (I152015,I2507,I1316652,I1316678,);
DFFARX1 I_77302 (I152018,I2507,I1316652,I1316695,);
not I_77303 (I1316703,I1316695);
nor I_77304 (I1316620,I1316678,I1316703);
DFFARX1 I_77305 (I1316703,I2507,I1316652,I1316635,);
nor I_77306 (I1316748,I152024,I152018);
and I_77307 (I1316765,I1316748,I152021);
nor I_77308 (I1316782,I1316765,I152024);
not I_77309 (I1316799,I152024);
and I_77310 (I1316816,I1316799,I152015);
nand I_77311 (I1316833,I1316816,I152033);
nor I_77312 (I1316850,I1316799,I1316833);
DFFARX1 I_77313 (I1316850,I2507,I1316652,I1316617,);
not I_77314 (I1316881,I1316833);
nand I_77315 (I1316898,I1316703,I1316881);
nand I_77316 (I1316629,I1316765,I1316881);
DFFARX1 I_77317 (I1316799,I2507,I1316652,I1316644,);
not I_77318 (I1316943,I152027);
nor I_77319 (I1316960,I1316943,I152015);
nor I_77320 (I1316977,I1316960,I1316782);
DFFARX1 I_77321 (I1316977,I2507,I1316652,I1316641,);
not I_77322 (I1317008,I1316960);
DFFARX1 I_77323 (I1317008,I2507,I1316652,I1317034,);
not I_77324 (I1317042,I1317034);
nor I_77325 (I1316638,I1317042,I1316960);
nor I_77326 (I1317073,I1316943,I152030);
and I_77327 (I1317090,I1317073,I152036);
or I_77328 (I1317107,I1317090,I152039);
DFFARX1 I_77329 (I1317107,I2507,I1316652,I1317133,);
not I_77330 (I1317141,I1317133);
nand I_77331 (I1317158,I1317141,I1316881);
not I_77332 (I1316632,I1317158);
nand I_77333 (I1316626,I1317158,I1316898);
nand I_77334 (I1316623,I1317141,I1316765);
not I_77335 (I1317247,I2514);
DFFARX1 I_77336 (I1172239,I2507,I1317247,I1317273,);
DFFARX1 I_77337 (I1172251,I2507,I1317247,I1317290,);
not I_77338 (I1317298,I1317290);
nor I_77339 (I1317215,I1317273,I1317298);
DFFARX1 I_77340 (I1317298,I2507,I1317247,I1317230,);
nor I_77341 (I1317343,I1172248,I1172242);
and I_77342 (I1317360,I1317343,I1172236);
nor I_77343 (I1317377,I1317360,I1172248);
not I_77344 (I1317394,I1172248);
and I_77345 (I1317411,I1317394,I1172245);
nand I_77346 (I1317428,I1317411,I1172236);
nor I_77347 (I1317445,I1317394,I1317428);
DFFARX1 I_77348 (I1317445,I2507,I1317247,I1317212,);
not I_77349 (I1317476,I1317428);
nand I_77350 (I1317493,I1317298,I1317476);
nand I_77351 (I1317224,I1317360,I1317476);
DFFARX1 I_77352 (I1317394,I2507,I1317247,I1317239,);
not I_77353 (I1317538,I1172260);
nor I_77354 (I1317555,I1317538,I1172245);
nor I_77355 (I1317572,I1317555,I1317377);
DFFARX1 I_77356 (I1317572,I2507,I1317247,I1317236,);
not I_77357 (I1317603,I1317555);
DFFARX1 I_77358 (I1317603,I2507,I1317247,I1317629,);
not I_77359 (I1317637,I1317629);
nor I_77360 (I1317233,I1317637,I1317555);
nor I_77361 (I1317668,I1317538,I1172254);
and I_77362 (I1317685,I1317668,I1172257);
or I_77363 (I1317702,I1317685,I1172239);
DFFARX1 I_77364 (I1317702,I2507,I1317247,I1317728,);
not I_77365 (I1317736,I1317728);
nand I_77366 (I1317753,I1317736,I1317476);
not I_77367 (I1317227,I1317753);
nand I_77368 (I1317221,I1317753,I1317493);
nand I_77369 (I1317218,I1317736,I1317360);
not I_77370 (I1317842,I2514);
DFFARX1 I_77371 (I615133,I2507,I1317842,I1317868,);
DFFARX1 I_77372 (I615127,I2507,I1317842,I1317885,);
not I_77373 (I1317893,I1317885);
nor I_77374 (I1317810,I1317868,I1317893);
DFFARX1 I_77375 (I1317893,I2507,I1317842,I1317825,);
nor I_77376 (I1317938,I615124,I615115);
and I_77377 (I1317955,I1317938,I615112);
nor I_77378 (I1317972,I1317955,I615124);
not I_77379 (I1317989,I615124);
and I_77380 (I1318006,I1317989,I615118);
nand I_77381 (I1318023,I1318006,I615130);
nor I_77382 (I1318040,I1317989,I1318023);
DFFARX1 I_77383 (I1318040,I2507,I1317842,I1317807,);
not I_77384 (I1318071,I1318023);
nand I_77385 (I1318088,I1317893,I1318071);
nand I_77386 (I1317819,I1317955,I1318071);
DFFARX1 I_77387 (I1317989,I2507,I1317842,I1317834,);
not I_77388 (I1318133,I615136);
nor I_77389 (I1318150,I1318133,I615118);
nor I_77390 (I1318167,I1318150,I1317972);
DFFARX1 I_77391 (I1318167,I2507,I1317842,I1317831,);
not I_77392 (I1318198,I1318150);
DFFARX1 I_77393 (I1318198,I2507,I1317842,I1318224,);
not I_77394 (I1318232,I1318224);
nor I_77395 (I1317828,I1318232,I1318150);
nor I_77396 (I1318263,I1318133,I615115);
and I_77397 (I1318280,I1318263,I615121);
or I_77398 (I1318297,I1318280,I615112);
DFFARX1 I_77399 (I1318297,I2507,I1317842,I1318323,);
not I_77400 (I1318331,I1318323);
nand I_77401 (I1318348,I1318331,I1318071);
not I_77402 (I1317822,I1318348);
nand I_77403 (I1317816,I1318348,I1318088);
nand I_77404 (I1317813,I1318331,I1317955);
not I_77405 (I1318437,I2514);
DFFARX1 I_77406 (I629583,I2507,I1318437,I1318463,);
DFFARX1 I_77407 (I629565,I2507,I1318437,I1318480,);
not I_77408 (I1318488,I1318480);
nor I_77409 (I1318405,I1318463,I1318488);
DFFARX1 I_77410 (I1318488,I2507,I1318437,I1318420,);
nor I_77411 (I1318533,I629571,I629574);
and I_77412 (I1318550,I1318533,I629562);
nor I_77413 (I1318567,I1318550,I629571);
not I_77414 (I1318584,I629571);
and I_77415 (I1318601,I1318584,I629580);
nand I_77416 (I1318618,I1318601,I629568);
nor I_77417 (I1318635,I1318584,I1318618);
DFFARX1 I_77418 (I1318635,I2507,I1318437,I1318402,);
not I_77419 (I1318666,I1318618);
nand I_77420 (I1318683,I1318488,I1318666);
nand I_77421 (I1318414,I1318550,I1318666);
DFFARX1 I_77422 (I1318584,I2507,I1318437,I1318429,);
not I_77423 (I1318728,I629565);
nor I_77424 (I1318745,I1318728,I629580);
nor I_77425 (I1318762,I1318745,I1318567);
DFFARX1 I_77426 (I1318762,I2507,I1318437,I1318426,);
not I_77427 (I1318793,I1318745);
DFFARX1 I_77428 (I1318793,I2507,I1318437,I1318819,);
not I_77429 (I1318827,I1318819);
nor I_77430 (I1318423,I1318827,I1318745);
nor I_77431 (I1318858,I1318728,I629577);
and I_77432 (I1318875,I1318858,I629586);
or I_77433 (I1318892,I1318875,I629562);
DFFARX1 I_77434 (I1318892,I2507,I1318437,I1318918,);
not I_77435 (I1318926,I1318918);
nand I_77436 (I1318943,I1318926,I1318666);
not I_77437 (I1318417,I1318943);
nand I_77438 (I1318411,I1318943,I1318683);
nand I_77439 (I1318408,I1318926,I1318550);
not I_77440 (I1319032,I2514);
DFFARX1 I_77441 (I374583,I2507,I1319032,I1319058,);
DFFARX1 I_77442 (I374577,I2507,I1319032,I1319075,);
not I_77443 (I1319083,I1319075);
nor I_77444 (I1319000,I1319058,I1319083);
DFFARX1 I_77445 (I1319083,I2507,I1319032,I1319015,);
nor I_77446 (I1319128,I374565,I374586);
and I_77447 (I1319145,I1319128,I374580);
nor I_77448 (I1319162,I1319145,I374565);
not I_77449 (I1319179,I374565);
and I_77450 (I1319196,I1319179,I374562);
nand I_77451 (I1319213,I1319196,I374574);
nor I_77452 (I1319230,I1319179,I1319213);
DFFARX1 I_77453 (I1319230,I2507,I1319032,I1318997,);
not I_77454 (I1319261,I1319213);
nand I_77455 (I1319278,I1319083,I1319261);
nand I_77456 (I1319009,I1319145,I1319261);
DFFARX1 I_77457 (I1319179,I2507,I1319032,I1319024,);
not I_77458 (I1319323,I374589);
nor I_77459 (I1319340,I1319323,I374562);
nor I_77460 (I1319357,I1319340,I1319162);
DFFARX1 I_77461 (I1319357,I2507,I1319032,I1319021,);
not I_77462 (I1319388,I1319340);
DFFARX1 I_77463 (I1319388,I2507,I1319032,I1319414,);
not I_77464 (I1319422,I1319414);
nor I_77465 (I1319018,I1319422,I1319340);
nor I_77466 (I1319453,I1319323,I374571);
and I_77467 (I1319470,I1319453,I374568);
or I_77468 (I1319487,I1319470,I374562);
DFFARX1 I_77469 (I1319487,I2507,I1319032,I1319513,);
not I_77470 (I1319521,I1319513);
nand I_77471 (I1319538,I1319521,I1319261);
not I_77472 (I1319012,I1319538);
nand I_77473 (I1319006,I1319538,I1319278);
nand I_77474 (I1319003,I1319521,I1319145);
not I_77475 (I1319627,I2514);
DFFARX1 I_77476 (I844417,I2507,I1319627,I1319653,);
DFFARX1 I_77477 (I844414,I2507,I1319627,I1319670,);
not I_77478 (I1319678,I1319670);
nor I_77479 (I1319595,I1319653,I1319678);
DFFARX1 I_77480 (I1319678,I2507,I1319627,I1319610,);
nor I_77481 (I1319723,I844429,I844411);
and I_77482 (I1319740,I1319723,I844408);
nor I_77483 (I1319757,I1319740,I844429);
not I_77484 (I1319774,I844429);
and I_77485 (I1319791,I1319774,I844414);
nand I_77486 (I1319808,I1319791,I844426);
nor I_77487 (I1319825,I1319774,I1319808);
DFFARX1 I_77488 (I1319825,I2507,I1319627,I1319592,);
not I_77489 (I1319856,I1319808);
nand I_77490 (I1319873,I1319678,I1319856);
nand I_77491 (I1319604,I1319740,I1319856);
DFFARX1 I_77492 (I1319774,I2507,I1319627,I1319619,);
not I_77493 (I1319918,I844420);
nor I_77494 (I1319935,I1319918,I844414);
nor I_77495 (I1319952,I1319935,I1319757);
DFFARX1 I_77496 (I1319952,I2507,I1319627,I1319616,);
not I_77497 (I1319983,I1319935);
DFFARX1 I_77498 (I1319983,I2507,I1319627,I1320009,);
not I_77499 (I1320017,I1320009);
nor I_77500 (I1319613,I1320017,I1319935);
nor I_77501 (I1320048,I1319918,I844408);
and I_77502 (I1320065,I1320048,I844423);
or I_77503 (I1320082,I1320065,I844411);
DFFARX1 I_77504 (I1320082,I2507,I1319627,I1320108,);
not I_77505 (I1320116,I1320108);
nand I_77506 (I1320133,I1320116,I1319856);
not I_77507 (I1319607,I1320133);
nand I_77508 (I1319601,I1320133,I1319873);
nand I_77509 (I1319598,I1320116,I1319740);
not I_77510 (I1320222,I2514);
DFFARX1 I_77511 (I93352,I2507,I1320222,I1320248,);
DFFARX1 I_77512 (I93340,I2507,I1320222,I1320265,);
not I_77513 (I1320273,I1320265);
nor I_77514 (I1320190,I1320248,I1320273);
DFFARX1 I_77515 (I1320273,I2507,I1320222,I1320205,);
nor I_77516 (I1320318,I93331,I93355);
and I_77517 (I1320335,I1320318,I93334);
nor I_77518 (I1320352,I1320335,I93331);
not I_77519 (I1320369,I93331);
and I_77520 (I1320386,I1320369,I93337);
nand I_77521 (I1320403,I1320386,I93349);
nor I_77522 (I1320420,I1320369,I1320403);
DFFARX1 I_77523 (I1320420,I2507,I1320222,I1320187,);
not I_77524 (I1320451,I1320403);
nand I_77525 (I1320468,I1320273,I1320451);
nand I_77526 (I1320199,I1320335,I1320451);
DFFARX1 I_77527 (I1320369,I2507,I1320222,I1320214,);
not I_77528 (I1320513,I93331);
nor I_77529 (I1320530,I1320513,I93337);
nor I_77530 (I1320547,I1320530,I1320352);
DFFARX1 I_77531 (I1320547,I2507,I1320222,I1320211,);
not I_77532 (I1320578,I1320530);
DFFARX1 I_77533 (I1320578,I2507,I1320222,I1320604,);
not I_77534 (I1320612,I1320604);
nor I_77535 (I1320208,I1320612,I1320530);
nor I_77536 (I1320643,I1320513,I93334);
and I_77537 (I1320660,I1320643,I93343);
or I_77538 (I1320677,I1320660,I93346);
DFFARX1 I_77539 (I1320677,I2507,I1320222,I1320703,);
not I_77540 (I1320711,I1320703);
nand I_77541 (I1320728,I1320711,I1320451);
not I_77542 (I1320202,I1320728);
nand I_77543 (I1320196,I1320728,I1320468);
nand I_77544 (I1320193,I1320711,I1320335);
not I_77545 (I1320817,I2514);
DFFARX1 I_77546 (I1032032,I2507,I1320817,I1320843,);
DFFARX1 I_77547 (I1032023,I2507,I1320817,I1320860,);
not I_77548 (I1320868,I1320860);
nor I_77549 (I1320785,I1320843,I1320868);
DFFARX1 I_77550 (I1320868,I2507,I1320817,I1320800,);
nor I_77551 (I1320913,I1032029,I1032038);
and I_77552 (I1320930,I1320913,I1032041);
nor I_77553 (I1320947,I1320930,I1032029);
not I_77554 (I1320964,I1032029);
and I_77555 (I1320981,I1320964,I1032020);
nand I_77556 (I1320998,I1320981,I1032026);
nor I_77557 (I1321015,I1320964,I1320998);
DFFARX1 I_77558 (I1321015,I2507,I1320817,I1320782,);
not I_77559 (I1321046,I1320998);
nand I_77560 (I1321063,I1320868,I1321046);
nand I_77561 (I1320794,I1320930,I1321046);
DFFARX1 I_77562 (I1320964,I2507,I1320817,I1320809,);
not I_77563 (I1321108,I1032035);
nor I_77564 (I1321125,I1321108,I1032020);
nor I_77565 (I1321142,I1321125,I1320947);
DFFARX1 I_77566 (I1321142,I2507,I1320817,I1320806,);
not I_77567 (I1321173,I1321125);
DFFARX1 I_77568 (I1321173,I2507,I1320817,I1321199,);
not I_77569 (I1321207,I1321199);
nor I_77570 (I1320803,I1321207,I1321125);
nor I_77571 (I1321238,I1321108,I1032020);
and I_77572 (I1321255,I1321238,I1032023);
or I_77573 (I1321272,I1321255,I1032026);
DFFARX1 I_77574 (I1321272,I2507,I1320817,I1321298,);
not I_77575 (I1321306,I1321298);
nand I_77576 (I1321323,I1321306,I1321046);
not I_77577 (I1320797,I1321323);
nand I_77578 (I1320791,I1321323,I1321063);
nand I_77579 (I1320788,I1321306,I1320930);
not I_77580 (I1321412,I2514);
DFFARX1 I_77581 (I30636,I2507,I1321412,I1321438,);
DFFARX1 I_77582 (I30618,I2507,I1321412,I1321455,);
not I_77583 (I1321463,I1321455);
nor I_77584 (I1321380,I1321438,I1321463);
DFFARX1 I_77585 (I1321463,I2507,I1321412,I1321395,);
nor I_77586 (I1321508,I30618,I30633);
and I_77587 (I1321525,I1321508,I30627);
nor I_77588 (I1321542,I1321525,I30618);
not I_77589 (I1321559,I30618);
and I_77590 (I1321576,I1321559,I30621);
nand I_77591 (I1321593,I1321576,I30624);
nor I_77592 (I1321610,I1321559,I1321593);
DFFARX1 I_77593 (I1321610,I2507,I1321412,I1321377,);
not I_77594 (I1321641,I1321593);
nand I_77595 (I1321658,I1321463,I1321641);
nand I_77596 (I1321389,I1321525,I1321641);
DFFARX1 I_77597 (I1321559,I2507,I1321412,I1321404,);
not I_77598 (I1321703,I30630);
nor I_77599 (I1321720,I1321703,I30621);
nor I_77600 (I1321737,I1321720,I1321542);
DFFARX1 I_77601 (I1321737,I2507,I1321412,I1321401,);
not I_77602 (I1321768,I1321720);
DFFARX1 I_77603 (I1321768,I2507,I1321412,I1321794,);
not I_77604 (I1321802,I1321794);
nor I_77605 (I1321398,I1321802,I1321720);
nor I_77606 (I1321833,I1321703,I30642);
and I_77607 (I1321850,I1321833,I30639);
or I_77608 (I1321867,I1321850,I30621);
DFFARX1 I_77609 (I1321867,I2507,I1321412,I1321893,);
not I_77610 (I1321901,I1321893);
nand I_77611 (I1321918,I1321901,I1321641);
not I_77612 (I1321392,I1321918);
nand I_77613 (I1321386,I1321918,I1321658);
nand I_77614 (I1321383,I1321901,I1321525);
not I_77615 (I1322007,I2514);
DFFARX1 I_77616 (I709925,I2507,I1322007,I1322033,);
DFFARX1 I_77617 (I709907,I2507,I1322007,I1322050,);
not I_77618 (I1322058,I1322050);
nor I_77619 (I1321975,I1322033,I1322058);
DFFARX1 I_77620 (I1322058,I2507,I1322007,I1321990,);
nor I_77621 (I1322103,I709913,I709916);
and I_77622 (I1322120,I1322103,I709904);
nor I_77623 (I1322137,I1322120,I709913);
not I_77624 (I1322154,I709913);
and I_77625 (I1322171,I1322154,I709922);
nand I_77626 (I1322188,I1322171,I709910);
nor I_77627 (I1322205,I1322154,I1322188);
DFFARX1 I_77628 (I1322205,I2507,I1322007,I1321972,);
not I_77629 (I1322236,I1322188);
nand I_77630 (I1322253,I1322058,I1322236);
nand I_77631 (I1321984,I1322120,I1322236);
DFFARX1 I_77632 (I1322154,I2507,I1322007,I1321999,);
not I_77633 (I1322298,I709907);
nor I_77634 (I1322315,I1322298,I709922);
nor I_77635 (I1322332,I1322315,I1322137);
DFFARX1 I_77636 (I1322332,I2507,I1322007,I1321996,);
not I_77637 (I1322363,I1322315);
DFFARX1 I_77638 (I1322363,I2507,I1322007,I1322389,);
not I_77639 (I1322397,I1322389);
nor I_77640 (I1321993,I1322397,I1322315);
nor I_77641 (I1322428,I1322298,I709919);
and I_77642 (I1322445,I1322428,I709928);
or I_77643 (I1322462,I1322445,I709904);
DFFARX1 I_77644 (I1322462,I2507,I1322007,I1322488,);
not I_77645 (I1322496,I1322488);
nand I_77646 (I1322513,I1322496,I1322236);
not I_77647 (I1321987,I1322513);
nand I_77648 (I1321981,I1322513,I1322253);
nand I_77649 (I1321978,I1322496,I1322120);
not I_77650 (I1322602,I2514);
DFFARX1 I_77651 (I504799,I2507,I1322602,I1322628,);
DFFARX1 I_77652 (I504802,I2507,I1322602,I1322645,);
not I_77653 (I1322653,I1322645);
nor I_77654 (I1322570,I1322628,I1322653);
DFFARX1 I_77655 (I1322653,I2507,I1322602,I1322585,);
nor I_77656 (I1322698,I504805,I504823);
and I_77657 (I1322715,I1322698,I504808);
nor I_77658 (I1322732,I1322715,I504805);
not I_77659 (I1322749,I504805);
and I_77660 (I1322766,I1322749,I504817);
nand I_77661 (I1322783,I1322766,I504820);
nor I_77662 (I1322800,I1322749,I1322783);
DFFARX1 I_77663 (I1322800,I2507,I1322602,I1322567,);
not I_77664 (I1322831,I1322783);
nand I_77665 (I1322848,I1322653,I1322831);
nand I_77666 (I1322579,I1322715,I1322831);
DFFARX1 I_77667 (I1322749,I2507,I1322602,I1322594,);
not I_77668 (I1322893,I504811);
nor I_77669 (I1322910,I1322893,I504817);
nor I_77670 (I1322927,I1322910,I1322732);
DFFARX1 I_77671 (I1322927,I2507,I1322602,I1322591,);
not I_77672 (I1322958,I1322910);
DFFARX1 I_77673 (I1322958,I2507,I1322602,I1322984,);
not I_77674 (I1322992,I1322984);
nor I_77675 (I1322588,I1322992,I1322910);
nor I_77676 (I1323023,I1322893,I504799);
and I_77677 (I1323040,I1323023,I504814);
or I_77678 (I1323057,I1323040,I504802);
DFFARX1 I_77679 (I1323057,I2507,I1322602,I1323083,);
not I_77680 (I1323091,I1323083);
nand I_77681 (I1323108,I1323091,I1322831);
not I_77682 (I1322582,I1323108);
nand I_77683 (I1322576,I1323108,I1322848);
nand I_77684 (I1322573,I1323091,I1322715);
not I_77685 (I1323197,I2514);
DFFARX1 I_77686 (I930859,I2507,I1323197,I1323223,);
DFFARX1 I_77687 (I930877,I2507,I1323197,I1323240,);
not I_77688 (I1323248,I1323240);
nor I_77689 (I1323165,I1323223,I1323248);
DFFARX1 I_77690 (I1323248,I2507,I1323197,I1323180,);
nor I_77691 (I1323293,I930856,I930868);
and I_77692 (I1323310,I1323293,I930853);
nor I_77693 (I1323327,I1323310,I930856);
not I_77694 (I1323344,I930856);
and I_77695 (I1323361,I1323344,I930862);
nand I_77696 (I1323378,I1323361,I930874);
nor I_77697 (I1323395,I1323344,I1323378);
DFFARX1 I_77698 (I1323395,I2507,I1323197,I1323162,);
not I_77699 (I1323426,I1323378);
nand I_77700 (I1323443,I1323248,I1323426);
nand I_77701 (I1323174,I1323310,I1323426);
DFFARX1 I_77702 (I1323344,I2507,I1323197,I1323189,);
not I_77703 (I1323488,I930865);
nor I_77704 (I1323505,I1323488,I930862);
nor I_77705 (I1323522,I1323505,I1323327);
DFFARX1 I_77706 (I1323522,I2507,I1323197,I1323186,);
not I_77707 (I1323553,I1323505);
DFFARX1 I_77708 (I1323553,I2507,I1323197,I1323579,);
not I_77709 (I1323587,I1323579);
nor I_77710 (I1323183,I1323587,I1323505);
nor I_77711 (I1323618,I1323488,I930853);
and I_77712 (I1323635,I1323618,I930880);
or I_77713 (I1323652,I1323635,I930871);
DFFARX1 I_77714 (I1323652,I2507,I1323197,I1323678,);
not I_77715 (I1323686,I1323678);
nand I_77716 (I1323703,I1323686,I1323426);
not I_77717 (I1323177,I1323703);
nand I_77718 (I1323171,I1323703,I1323443);
nand I_77719 (I1323168,I1323686,I1323310);
not I_77720 (I1323792,I2514);
DFFARX1 I_77721 (I402799,I2507,I1323792,I1323818,);
DFFARX1 I_77722 (I402805,I2507,I1323792,I1323835,);
not I_77723 (I1323843,I1323835);
nor I_77724 (I1323760,I1323818,I1323843);
DFFARX1 I_77725 (I1323843,I2507,I1323792,I1323775,);
nor I_77726 (I1323888,I402814,I402799);
and I_77727 (I1323905,I1323888,I402826);
nor I_77728 (I1323922,I1323905,I402814);
not I_77729 (I1323939,I402814);
and I_77730 (I1323956,I1323939,I402802);
nand I_77731 (I1323973,I1323956,I402823);
nor I_77732 (I1323990,I1323939,I1323973);
DFFARX1 I_77733 (I1323990,I2507,I1323792,I1323757,);
not I_77734 (I1324021,I1323973);
nand I_77735 (I1324038,I1323843,I1324021);
nand I_77736 (I1323769,I1323905,I1324021);
DFFARX1 I_77737 (I1323939,I2507,I1323792,I1323784,);
not I_77738 (I1324083,I402811);
nor I_77739 (I1324100,I1324083,I402802);
nor I_77740 (I1324117,I1324100,I1323922);
DFFARX1 I_77741 (I1324117,I2507,I1323792,I1323781,);
not I_77742 (I1324148,I1324100);
DFFARX1 I_77743 (I1324148,I2507,I1323792,I1324174,);
not I_77744 (I1324182,I1324174);
nor I_77745 (I1323778,I1324182,I1324100);
nor I_77746 (I1324213,I1324083,I402808);
and I_77747 (I1324230,I1324213,I402820);
or I_77748 (I1324247,I1324230,I402817);
DFFARX1 I_77749 (I1324247,I2507,I1323792,I1324273,);
not I_77750 (I1324281,I1324273);
nand I_77751 (I1324298,I1324281,I1324021);
not I_77752 (I1323772,I1324298);
nand I_77753 (I1323766,I1324298,I1324038);
nand I_77754 (I1323763,I1324281,I1323905);
not I_77755 (I1324387,I2514);
DFFARX1 I_77756 (I179980,I2507,I1324387,I1324413,);
DFFARX1 I_77757 (I179983,I2507,I1324387,I1324430,);
not I_77758 (I1324438,I1324430);
nor I_77759 (I1324355,I1324413,I1324438);
DFFARX1 I_77760 (I1324438,I2507,I1324387,I1324370,);
nor I_77761 (I1324483,I179989,I179983);
and I_77762 (I1324500,I1324483,I179986);
nor I_77763 (I1324517,I1324500,I179989);
not I_77764 (I1324534,I179989);
and I_77765 (I1324551,I1324534,I179980);
nand I_77766 (I1324568,I1324551,I179998);
nor I_77767 (I1324585,I1324534,I1324568);
DFFARX1 I_77768 (I1324585,I2507,I1324387,I1324352,);
not I_77769 (I1324616,I1324568);
nand I_77770 (I1324633,I1324438,I1324616);
nand I_77771 (I1324364,I1324500,I1324616);
DFFARX1 I_77772 (I1324534,I2507,I1324387,I1324379,);
not I_77773 (I1324678,I179992);
nor I_77774 (I1324695,I1324678,I179980);
nor I_77775 (I1324712,I1324695,I1324517);
DFFARX1 I_77776 (I1324712,I2507,I1324387,I1324376,);
not I_77777 (I1324743,I1324695);
DFFARX1 I_77778 (I1324743,I2507,I1324387,I1324769,);
not I_77779 (I1324777,I1324769);
nor I_77780 (I1324373,I1324777,I1324695);
nor I_77781 (I1324808,I1324678,I179995);
and I_77782 (I1324825,I1324808,I180001);
or I_77783 (I1324842,I1324825,I180004);
DFFARX1 I_77784 (I1324842,I2507,I1324387,I1324868,);
not I_77785 (I1324876,I1324868);
nand I_77786 (I1324893,I1324876,I1324616);
not I_77787 (I1324367,I1324893);
nand I_77788 (I1324361,I1324893,I1324633);
nand I_77789 (I1324358,I1324876,I1324500);
not I_77790 (I1324982,I2514);
DFFARX1 I_77791 (I1038764,I2507,I1324982,I1325008,);
DFFARX1 I_77792 (I1038755,I2507,I1324982,I1325025,);
not I_77793 (I1325033,I1325025);
nor I_77794 (I1324950,I1325008,I1325033);
DFFARX1 I_77795 (I1325033,I2507,I1324982,I1324965,);
nor I_77796 (I1325078,I1038761,I1038770);
and I_77797 (I1325095,I1325078,I1038773);
nor I_77798 (I1325112,I1325095,I1038761);
not I_77799 (I1325129,I1038761);
and I_77800 (I1325146,I1325129,I1038752);
nand I_77801 (I1325163,I1325146,I1038758);
nor I_77802 (I1325180,I1325129,I1325163);
DFFARX1 I_77803 (I1325180,I2507,I1324982,I1324947,);
not I_77804 (I1325211,I1325163);
nand I_77805 (I1325228,I1325033,I1325211);
nand I_77806 (I1324959,I1325095,I1325211);
DFFARX1 I_77807 (I1325129,I2507,I1324982,I1324974,);
not I_77808 (I1325273,I1038767);
nor I_77809 (I1325290,I1325273,I1038752);
nor I_77810 (I1325307,I1325290,I1325112);
DFFARX1 I_77811 (I1325307,I2507,I1324982,I1324971,);
not I_77812 (I1325338,I1325290);
DFFARX1 I_77813 (I1325338,I2507,I1324982,I1325364,);
not I_77814 (I1325372,I1325364);
nor I_77815 (I1324968,I1325372,I1325290);
nor I_77816 (I1325403,I1325273,I1038752);
and I_77817 (I1325420,I1325403,I1038755);
or I_77818 (I1325437,I1325420,I1038758);
DFFARX1 I_77819 (I1325437,I2507,I1324982,I1325463,);
not I_77820 (I1325471,I1325463);
nand I_77821 (I1325488,I1325471,I1325211);
not I_77822 (I1324962,I1325488);
nand I_77823 (I1324956,I1325488,I1325228);
nand I_77824 (I1324953,I1325471,I1325095);
not I_77825 (I1325577,I2514);
DFFARX1 I_77826 (I349287,I2507,I1325577,I1325603,);
DFFARX1 I_77827 (I349281,I2507,I1325577,I1325620,);
not I_77828 (I1325628,I1325620);
nor I_77829 (I1325545,I1325603,I1325628);
DFFARX1 I_77830 (I1325628,I2507,I1325577,I1325560,);
nor I_77831 (I1325673,I349269,I349290);
and I_77832 (I1325690,I1325673,I349284);
nor I_77833 (I1325707,I1325690,I349269);
not I_77834 (I1325724,I349269);
and I_77835 (I1325741,I1325724,I349266);
nand I_77836 (I1325758,I1325741,I349278);
nor I_77837 (I1325775,I1325724,I1325758);
DFFARX1 I_77838 (I1325775,I2507,I1325577,I1325542,);
not I_77839 (I1325806,I1325758);
nand I_77840 (I1325823,I1325628,I1325806);
nand I_77841 (I1325554,I1325690,I1325806);
DFFARX1 I_77842 (I1325724,I2507,I1325577,I1325569,);
not I_77843 (I1325868,I349293);
nor I_77844 (I1325885,I1325868,I349266);
nor I_77845 (I1325902,I1325885,I1325707);
DFFARX1 I_77846 (I1325902,I2507,I1325577,I1325566,);
not I_77847 (I1325933,I1325885);
DFFARX1 I_77848 (I1325933,I2507,I1325577,I1325959,);
not I_77849 (I1325967,I1325959);
nor I_77850 (I1325563,I1325967,I1325885);
nor I_77851 (I1325998,I1325868,I349275);
and I_77852 (I1326015,I1325998,I349272);
or I_77853 (I1326032,I1326015,I349266);
DFFARX1 I_77854 (I1326032,I2507,I1325577,I1326058,);
not I_77855 (I1326066,I1326058);
nand I_77856 (I1326083,I1326066,I1325806);
not I_77857 (I1325557,I1326083);
nand I_77858 (I1325551,I1326083,I1325823);
nand I_77859 (I1325548,I1326066,I1325690);
not I_77860 (I1326172,I2514);
DFFARX1 I_77861 (I693163,I2507,I1326172,I1326198,);
DFFARX1 I_77862 (I693145,I2507,I1326172,I1326215,);
not I_77863 (I1326223,I1326215);
nor I_77864 (I1326140,I1326198,I1326223);
DFFARX1 I_77865 (I1326223,I2507,I1326172,I1326155,);
nor I_77866 (I1326268,I693151,I693154);
and I_77867 (I1326285,I1326268,I693142);
nor I_77868 (I1326302,I1326285,I693151);
not I_77869 (I1326319,I693151);
and I_77870 (I1326336,I1326319,I693160);
nand I_77871 (I1326353,I1326336,I693148);
nor I_77872 (I1326370,I1326319,I1326353);
DFFARX1 I_77873 (I1326370,I2507,I1326172,I1326137,);
not I_77874 (I1326401,I1326353);
nand I_77875 (I1326418,I1326223,I1326401);
nand I_77876 (I1326149,I1326285,I1326401);
DFFARX1 I_77877 (I1326319,I2507,I1326172,I1326164,);
not I_77878 (I1326463,I693145);
nor I_77879 (I1326480,I1326463,I693160);
nor I_77880 (I1326497,I1326480,I1326302);
DFFARX1 I_77881 (I1326497,I2507,I1326172,I1326161,);
not I_77882 (I1326528,I1326480);
DFFARX1 I_77883 (I1326528,I2507,I1326172,I1326554,);
not I_77884 (I1326562,I1326554);
nor I_77885 (I1326158,I1326562,I1326480);
nor I_77886 (I1326593,I1326463,I693157);
and I_77887 (I1326610,I1326593,I693166);
or I_77888 (I1326627,I1326610,I693142);
DFFARX1 I_77889 (I1326627,I2507,I1326172,I1326653,);
not I_77890 (I1326661,I1326653);
nand I_77891 (I1326678,I1326661,I1326401);
not I_77892 (I1326152,I1326678);
nand I_77893 (I1326146,I1326678,I1326418);
nand I_77894 (I1326143,I1326661,I1326285);
not I_77895 (I1326767,I2514);
DFFARX1 I_77896 (I538119,I2507,I1326767,I1326793,);
DFFARX1 I_77897 (I538122,I2507,I1326767,I1326810,);
not I_77898 (I1326818,I1326810);
nor I_77899 (I1326735,I1326793,I1326818);
DFFARX1 I_77900 (I1326818,I2507,I1326767,I1326750,);
nor I_77901 (I1326863,I538125,I538143);
and I_77902 (I1326880,I1326863,I538128);
nor I_77903 (I1326897,I1326880,I538125);
not I_77904 (I1326914,I538125);
and I_77905 (I1326931,I1326914,I538137);
nand I_77906 (I1326948,I1326931,I538140);
nor I_77907 (I1326965,I1326914,I1326948);
DFFARX1 I_77908 (I1326965,I2507,I1326767,I1326732,);
not I_77909 (I1326996,I1326948);
nand I_77910 (I1327013,I1326818,I1326996);
nand I_77911 (I1326744,I1326880,I1326996);
DFFARX1 I_77912 (I1326914,I2507,I1326767,I1326759,);
not I_77913 (I1327058,I538131);
nor I_77914 (I1327075,I1327058,I538137);
nor I_77915 (I1327092,I1327075,I1326897);
DFFARX1 I_77916 (I1327092,I2507,I1326767,I1326756,);
not I_77917 (I1327123,I1327075);
DFFARX1 I_77918 (I1327123,I2507,I1326767,I1327149,);
not I_77919 (I1327157,I1327149);
nor I_77920 (I1326753,I1327157,I1327075);
nor I_77921 (I1327188,I1327058,I538119);
and I_77922 (I1327205,I1327188,I538134);
or I_77923 (I1327222,I1327205,I538122);
DFFARX1 I_77924 (I1327222,I2507,I1326767,I1327248,);
not I_77925 (I1327256,I1327248);
nand I_77926 (I1327273,I1327256,I1326996);
not I_77927 (I1326747,I1327273);
nand I_77928 (I1326741,I1327273,I1327013);
nand I_77929 (I1326738,I1327256,I1326880);
not I_77930 (I1327362,I2514);
DFFARX1 I_77931 (I316613,I2507,I1327362,I1327388,);
DFFARX1 I_77932 (I316607,I2507,I1327362,I1327405,);
not I_77933 (I1327413,I1327405);
nor I_77934 (I1327330,I1327388,I1327413);
DFFARX1 I_77935 (I1327413,I2507,I1327362,I1327345,);
nor I_77936 (I1327458,I316595,I316616);
and I_77937 (I1327475,I1327458,I316610);
nor I_77938 (I1327492,I1327475,I316595);
not I_77939 (I1327509,I316595);
and I_77940 (I1327526,I1327509,I316592);
nand I_77941 (I1327543,I1327526,I316604);
nor I_77942 (I1327560,I1327509,I1327543);
DFFARX1 I_77943 (I1327560,I2507,I1327362,I1327327,);
not I_77944 (I1327591,I1327543);
nand I_77945 (I1327608,I1327413,I1327591);
nand I_77946 (I1327339,I1327475,I1327591);
DFFARX1 I_77947 (I1327509,I2507,I1327362,I1327354,);
not I_77948 (I1327653,I316619);
nor I_77949 (I1327670,I1327653,I316592);
nor I_77950 (I1327687,I1327670,I1327492);
DFFARX1 I_77951 (I1327687,I2507,I1327362,I1327351,);
not I_77952 (I1327718,I1327670);
DFFARX1 I_77953 (I1327718,I2507,I1327362,I1327744,);
not I_77954 (I1327752,I1327744);
nor I_77955 (I1327348,I1327752,I1327670);
nor I_77956 (I1327783,I1327653,I316601);
and I_77957 (I1327800,I1327783,I316598);
or I_77958 (I1327817,I1327800,I316592);
DFFARX1 I_77959 (I1327817,I2507,I1327362,I1327843,);
not I_77960 (I1327851,I1327843);
nand I_77961 (I1327868,I1327851,I1327591);
not I_77962 (I1327342,I1327868);
nand I_77963 (I1327336,I1327868,I1327608);
nand I_77964 (I1327333,I1327851,I1327475);
not I_77965 (I1327957,I2514);
DFFARX1 I_77966 (I206160,I2507,I1327957,I1327983,);
DFFARX1 I_77967 (I206163,I2507,I1327957,I1328000,);
not I_77968 (I1328008,I1328000);
nor I_77969 (I1327925,I1327983,I1328008);
DFFARX1 I_77970 (I1328008,I2507,I1327957,I1327940,);
nor I_77971 (I1328053,I206169,I206163);
and I_77972 (I1328070,I1328053,I206166);
nor I_77973 (I1328087,I1328070,I206169);
not I_77974 (I1328104,I206169);
and I_77975 (I1328121,I1328104,I206160);
nand I_77976 (I1328138,I1328121,I206178);
nor I_77977 (I1328155,I1328104,I1328138);
DFFARX1 I_77978 (I1328155,I2507,I1327957,I1327922,);
not I_77979 (I1328186,I1328138);
nand I_77980 (I1328203,I1328008,I1328186);
nand I_77981 (I1327934,I1328070,I1328186);
DFFARX1 I_77982 (I1328104,I2507,I1327957,I1327949,);
not I_77983 (I1328248,I206172);
nor I_77984 (I1328265,I1328248,I206160);
nor I_77985 (I1328282,I1328265,I1328087);
DFFARX1 I_77986 (I1328282,I2507,I1327957,I1327946,);
not I_77987 (I1328313,I1328265);
DFFARX1 I_77988 (I1328313,I2507,I1327957,I1328339,);
not I_77989 (I1328347,I1328339);
nor I_77990 (I1327943,I1328347,I1328265);
nor I_77991 (I1328378,I1328248,I206175);
and I_77992 (I1328395,I1328378,I206181);
or I_77993 (I1328412,I1328395,I206184);
DFFARX1 I_77994 (I1328412,I2507,I1327957,I1328438,);
not I_77995 (I1328446,I1328438);
nand I_77996 (I1328463,I1328446,I1328186);
not I_77997 (I1327937,I1328463);
nand I_77998 (I1327931,I1328463,I1328203);
nand I_77999 (I1327928,I1328446,I1328070);
not I_78000 (I1328552,I2514);
DFFARX1 I_78001 (I1105191,I2507,I1328552,I1328578,);
DFFARX1 I_78002 (I1105203,I2507,I1328552,I1328595,);
not I_78003 (I1328603,I1328595);
nor I_78004 (I1328520,I1328578,I1328603);
DFFARX1 I_78005 (I1328603,I2507,I1328552,I1328535,);
nor I_78006 (I1328648,I1105200,I1105194);
and I_78007 (I1328665,I1328648,I1105188);
nor I_78008 (I1328682,I1328665,I1105200);
not I_78009 (I1328699,I1105200);
and I_78010 (I1328716,I1328699,I1105197);
nand I_78011 (I1328733,I1328716,I1105188);
nor I_78012 (I1328750,I1328699,I1328733);
DFFARX1 I_78013 (I1328750,I2507,I1328552,I1328517,);
not I_78014 (I1328781,I1328733);
nand I_78015 (I1328798,I1328603,I1328781);
nand I_78016 (I1328529,I1328665,I1328781);
DFFARX1 I_78017 (I1328699,I2507,I1328552,I1328544,);
not I_78018 (I1328843,I1105212);
nor I_78019 (I1328860,I1328843,I1105197);
nor I_78020 (I1328877,I1328860,I1328682);
DFFARX1 I_78021 (I1328877,I2507,I1328552,I1328541,);
not I_78022 (I1328908,I1328860);
DFFARX1 I_78023 (I1328908,I2507,I1328552,I1328934,);
not I_78024 (I1328942,I1328934);
nor I_78025 (I1328538,I1328942,I1328860);
nor I_78026 (I1328973,I1328843,I1105206);
and I_78027 (I1328990,I1328973,I1105209);
or I_78028 (I1329007,I1328990,I1105191);
DFFARX1 I_78029 (I1329007,I2507,I1328552,I1329033,);
not I_78030 (I1329041,I1329033);
nand I_78031 (I1329058,I1329041,I1328781);
not I_78032 (I1328532,I1329058);
nand I_78033 (I1328526,I1329058,I1328798);
nand I_78034 (I1328523,I1329041,I1328665);
not I_78035 (I1329147,I2514);
DFFARX1 I_78036 (I234720,I2507,I1329147,I1329173,);
DFFARX1 I_78037 (I234723,I2507,I1329147,I1329190,);
not I_78038 (I1329198,I1329190);
nor I_78039 (I1329115,I1329173,I1329198);
DFFARX1 I_78040 (I1329198,I2507,I1329147,I1329130,);
nor I_78041 (I1329243,I234729,I234723);
and I_78042 (I1329260,I1329243,I234726);
nor I_78043 (I1329277,I1329260,I234729);
not I_78044 (I1329294,I234729);
and I_78045 (I1329311,I1329294,I234720);
nand I_78046 (I1329328,I1329311,I234738);
nor I_78047 (I1329345,I1329294,I1329328);
DFFARX1 I_78048 (I1329345,I2507,I1329147,I1329112,);
not I_78049 (I1329376,I1329328);
nand I_78050 (I1329393,I1329198,I1329376);
nand I_78051 (I1329124,I1329260,I1329376);
DFFARX1 I_78052 (I1329294,I2507,I1329147,I1329139,);
not I_78053 (I1329438,I234732);
nor I_78054 (I1329455,I1329438,I234720);
nor I_78055 (I1329472,I1329455,I1329277);
DFFARX1 I_78056 (I1329472,I2507,I1329147,I1329136,);
not I_78057 (I1329503,I1329455);
DFFARX1 I_78058 (I1329503,I2507,I1329147,I1329529,);
not I_78059 (I1329537,I1329529);
nor I_78060 (I1329133,I1329537,I1329455);
nor I_78061 (I1329568,I1329438,I234735);
and I_78062 (I1329585,I1329568,I234741);
or I_78063 (I1329602,I1329585,I234744);
DFFARX1 I_78064 (I1329602,I2507,I1329147,I1329628,);
not I_78065 (I1329636,I1329628);
nand I_78066 (I1329653,I1329636,I1329376);
not I_78067 (I1329127,I1329653);
nand I_78068 (I1329121,I1329653,I1329393);
nand I_78069 (I1329118,I1329636,I1329260);
not I_78070 (I1329742,I2514);
DFFARX1 I_78071 (I413135,I2507,I1329742,I1329768,);
DFFARX1 I_78072 (I413141,I2507,I1329742,I1329785,);
not I_78073 (I1329793,I1329785);
nor I_78074 (I1329710,I1329768,I1329793);
DFFARX1 I_78075 (I1329793,I2507,I1329742,I1329725,);
nor I_78076 (I1329838,I413150,I413135);
and I_78077 (I1329855,I1329838,I413162);
nor I_78078 (I1329872,I1329855,I413150);
not I_78079 (I1329889,I413150);
and I_78080 (I1329906,I1329889,I413138);
nand I_78081 (I1329923,I1329906,I413159);
nor I_78082 (I1329940,I1329889,I1329923);
DFFARX1 I_78083 (I1329940,I2507,I1329742,I1329707,);
not I_78084 (I1329971,I1329923);
nand I_78085 (I1329988,I1329793,I1329971);
nand I_78086 (I1329719,I1329855,I1329971);
DFFARX1 I_78087 (I1329889,I2507,I1329742,I1329734,);
not I_78088 (I1330033,I413147);
nor I_78089 (I1330050,I1330033,I413138);
nor I_78090 (I1330067,I1330050,I1329872);
DFFARX1 I_78091 (I1330067,I2507,I1329742,I1329731,);
not I_78092 (I1330098,I1330050);
DFFARX1 I_78093 (I1330098,I2507,I1329742,I1330124,);
not I_78094 (I1330132,I1330124);
nor I_78095 (I1329728,I1330132,I1330050);
nor I_78096 (I1330163,I1330033,I413144);
and I_78097 (I1330180,I1330163,I413156);
or I_78098 (I1330197,I1330180,I413153);
DFFARX1 I_78099 (I1330197,I2507,I1329742,I1330223,);
not I_78100 (I1330231,I1330223);
nand I_78101 (I1330248,I1330231,I1329971);
not I_78102 (I1329722,I1330248);
nand I_78103 (I1329716,I1330248,I1329988);
nand I_78104 (I1329713,I1330231,I1329855);
not I_78105 (I1330337,I2514);
DFFARX1 I_78106 (I824391,I2507,I1330337,I1330363,);
DFFARX1 I_78107 (I824388,I2507,I1330337,I1330380,);
not I_78108 (I1330388,I1330380);
nor I_78109 (I1330305,I1330363,I1330388);
DFFARX1 I_78110 (I1330388,I2507,I1330337,I1330320,);
nor I_78111 (I1330433,I824403,I824385);
and I_78112 (I1330450,I1330433,I824382);
nor I_78113 (I1330467,I1330450,I824403);
not I_78114 (I1330484,I824403);
and I_78115 (I1330501,I1330484,I824388);
nand I_78116 (I1330518,I1330501,I824400);
nor I_78117 (I1330535,I1330484,I1330518);
DFFARX1 I_78118 (I1330535,I2507,I1330337,I1330302,);
not I_78119 (I1330566,I1330518);
nand I_78120 (I1330583,I1330388,I1330566);
nand I_78121 (I1330314,I1330450,I1330566);
DFFARX1 I_78122 (I1330484,I2507,I1330337,I1330329,);
not I_78123 (I1330628,I824394);
nor I_78124 (I1330645,I1330628,I824388);
nor I_78125 (I1330662,I1330645,I1330467);
DFFARX1 I_78126 (I1330662,I2507,I1330337,I1330326,);
not I_78127 (I1330693,I1330645);
DFFARX1 I_78128 (I1330693,I2507,I1330337,I1330719,);
not I_78129 (I1330727,I1330719);
nor I_78130 (I1330323,I1330727,I1330645);
nor I_78131 (I1330758,I1330628,I824382);
and I_78132 (I1330775,I1330758,I824397);
or I_78133 (I1330792,I1330775,I824385);
DFFARX1 I_78134 (I1330792,I2507,I1330337,I1330818,);
not I_78135 (I1330826,I1330818);
nand I_78136 (I1330843,I1330826,I1330566);
not I_78137 (I1330317,I1330843);
nand I_78138 (I1330311,I1330843,I1330583);
nand I_78139 (I1330308,I1330826,I1330450);
not I_78140 (I1330932,I2514);
DFFARX1 I_78141 (I296587,I2507,I1330932,I1330958,);
DFFARX1 I_78142 (I296581,I2507,I1330932,I1330975,);
not I_78143 (I1330983,I1330975);
nor I_78144 (I1330900,I1330958,I1330983);
DFFARX1 I_78145 (I1330983,I2507,I1330932,I1330915,);
nor I_78146 (I1331028,I296569,I296590);
and I_78147 (I1331045,I1331028,I296584);
nor I_78148 (I1331062,I1331045,I296569);
not I_78149 (I1331079,I296569);
and I_78150 (I1331096,I1331079,I296566);
nand I_78151 (I1331113,I1331096,I296578);
nor I_78152 (I1331130,I1331079,I1331113);
DFFARX1 I_78153 (I1331130,I2507,I1330932,I1330897,);
not I_78154 (I1331161,I1331113);
nand I_78155 (I1331178,I1330983,I1331161);
nand I_78156 (I1330909,I1331045,I1331161);
DFFARX1 I_78157 (I1331079,I2507,I1330932,I1330924,);
not I_78158 (I1331223,I296593);
nor I_78159 (I1331240,I1331223,I296566);
nor I_78160 (I1331257,I1331240,I1331062);
DFFARX1 I_78161 (I1331257,I2507,I1330932,I1330921,);
not I_78162 (I1331288,I1331240);
DFFARX1 I_78163 (I1331288,I2507,I1330932,I1331314,);
not I_78164 (I1331322,I1331314);
nor I_78165 (I1330918,I1331322,I1331240);
nor I_78166 (I1331353,I1331223,I296575);
and I_78167 (I1331370,I1331353,I296572);
or I_78168 (I1331387,I1331370,I296566);
DFFARX1 I_78169 (I1331387,I2507,I1330932,I1331413,);
not I_78170 (I1331421,I1331413);
nand I_78171 (I1331438,I1331421,I1331161);
not I_78172 (I1330912,I1331438);
nand I_78173 (I1330906,I1331438,I1331178);
nand I_78174 (I1330903,I1331421,I1331045);
not I_78175 (I1331527,I2514);
DFFARX1 I_78176 (I1174551,I2507,I1331527,I1331553,);
DFFARX1 I_78177 (I1174563,I2507,I1331527,I1331570,);
not I_78178 (I1331578,I1331570);
nor I_78179 (I1331495,I1331553,I1331578);
DFFARX1 I_78180 (I1331578,I2507,I1331527,I1331510,);
nor I_78181 (I1331623,I1174560,I1174554);
and I_78182 (I1331640,I1331623,I1174548);
nor I_78183 (I1331657,I1331640,I1174560);
not I_78184 (I1331674,I1174560);
and I_78185 (I1331691,I1331674,I1174557);
nand I_78186 (I1331708,I1331691,I1174548);
nor I_78187 (I1331725,I1331674,I1331708);
DFFARX1 I_78188 (I1331725,I2507,I1331527,I1331492,);
not I_78189 (I1331756,I1331708);
nand I_78190 (I1331773,I1331578,I1331756);
nand I_78191 (I1331504,I1331640,I1331756);
DFFARX1 I_78192 (I1331674,I2507,I1331527,I1331519,);
not I_78193 (I1331818,I1174572);
nor I_78194 (I1331835,I1331818,I1174557);
nor I_78195 (I1331852,I1331835,I1331657);
DFFARX1 I_78196 (I1331852,I2507,I1331527,I1331516,);
not I_78197 (I1331883,I1331835);
DFFARX1 I_78198 (I1331883,I2507,I1331527,I1331909,);
not I_78199 (I1331917,I1331909);
nor I_78200 (I1331513,I1331917,I1331835);
nor I_78201 (I1331948,I1331818,I1174566);
and I_78202 (I1331965,I1331948,I1174569);
or I_78203 (I1331982,I1331965,I1174551);
DFFARX1 I_78204 (I1331982,I2507,I1331527,I1332008,);
not I_78205 (I1332016,I1332008);
nand I_78206 (I1332033,I1332016,I1331756);
not I_78207 (I1331507,I1332033);
nand I_78208 (I1331501,I1332033,I1331773);
nand I_78209 (I1331498,I1332016,I1331640);
not I_78210 (I1332122,I2514);
DFFARX1 I_78211 (I1216674,I2507,I1332122,I1332148,);
DFFARX1 I_78212 (I1216677,I2507,I1332122,I1332165,);
not I_78213 (I1332173,I1332165);
nor I_78214 (I1332090,I1332148,I1332173);
DFFARX1 I_78215 (I1332173,I2507,I1332122,I1332105,);
nor I_78216 (I1332218,I1216677,I1216692);
and I_78217 (I1332235,I1332218,I1216686);
nor I_78218 (I1332252,I1332235,I1216677);
not I_78219 (I1332269,I1216677);
and I_78220 (I1332286,I1332269,I1216695);
nand I_78221 (I1332303,I1332286,I1216683);
nor I_78222 (I1332320,I1332269,I1332303);
DFFARX1 I_78223 (I1332320,I2507,I1332122,I1332087,);
not I_78224 (I1332351,I1332303);
nand I_78225 (I1332368,I1332173,I1332351);
nand I_78226 (I1332099,I1332235,I1332351);
DFFARX1 I_78227 (I1332269,I2507,I1332122,I1332114,);
not I_78228 (I1332413,I1216689);
nor I_78229 (I1332430,I1332413,I1216695);
nor I_78230 (I1332447,I1332430,I1332252);
DFFARX1 I_78231 (I1332447,I2507,I1332122,I1332111,);
not I_78232 (I1332478,I1332430);
DFFARX1 I_78233 (I1332478,I2507,I1332122,I1332504,);
not I_78234 (I1332512,I1332504);
nor I_78235 (I1332108,I1332512,I1332430);
nor I_78236 (I1332543,I1332413,I1216674);
and I_78237 (I1332560,I1332543,I1216698);
or I_78238 (I1332577,I1332560,I1216680);
DFFARX1 I_78239 (I1332577,I2507,I1332122,I1332603,);
not I_78240 (I1332611,I1332603);
nand I_78241 (I1332628,I1332611,I1332351);
not I_78242 (I1332102,I1332628);
nand I_78243 (I1332096,I1332628,I1332368);
nand I_78244 (I1332093,I1332611,I1332235);
not I_78245 (I1332717,I2514);
DFFARX1 I_78246 (I871294,I2507,I1332717,I1332743,);
DFFARX1 I_78247 (I871291,I2507,I1332717,I1332760,);
not I_78248 (I1332768,I1332760);
nor I_78249 (I1332685,I1332743,I1332768);
DFFARX1 I_78250 (I1332768,I2507,I1332717,I1332700,);
nor I_78251 (I1332813,I871306,I871288);
and I_78252 (I1332830,I1332813,I871285);
nor I_78253 (I1332847,I1332830,I871306);
not I_78254 (I1332864,I871306);
and I_78255 (I1332881,I1332864,I871291);
nand I_78256 (I1332898,I1332881,I871303);
nor I_78257 (I1332915,I1332864,I1332898);
DFFARX1 I_78258 (I1332915,I2507,I1332717,I1332682,);
not I_78259 (I1332946,I1332898);
nand I_78260 (I1332963,I1332768,I1332946);
nand I_78261 (I1332694,I1332830,I1332946);
DFFARX1 I_78262 (I1332864,I2507,I1332717,I1332709,);
not I_78263 (I1333008,I871297);
nor I_78264 (I1333025,I1333008,I871291);
nor I_78265 (I1333042,I1333025,I1332847);
DFFARX1 I_78266 (I1333042,I2507,I1332717,I1332706,);
not I_78267 (I1333073,I1333025);
DFFARX1 I_78268 (I1333073,I2507,I1332717,I1333099,);
not I_78269 (I1333107,I1333099);
nor I_78270 (I1332703,I1333107,I1333025);
nor I_78271 (I1333138,I1333008,I871285);
and I_78272 (I1333155,I1333138,I871300);
or I_78273 (I1333172,I1333155,I871288);
DFFARX1 I_78274 (I1333172,I2507,I1332717,I1333198,);
not I_78275 (I1333206,I1333198);
nand I_78276 (I1333223,I1333206,I1332946);
not I_78277 (I1332697,I1333223);
nand I_78278 (I1332691,I1333223,I1332963);
nand I_78279 (I1332688,I1333206,I1332830);
not I_78280 (I1333312,I2514);
DFFARX1 I_78281 (I994167,I2507,I1333312,I1333338,);
DFFARX1 I_78282 (I994185,I2507,I1333312,I1333355,);
not I_78283 (I1333363,I1333355);
nor I_78284 (I1333280,I1333338,I1333363);
DFFARX1 I_78285 (I1333363,I2507,I1333312,I1333295,);
nor I_78286 (I1333408,I994164,I994176);
and I_78287 (I1333425,I1333408,I994161);
nor I_78288 (I1333442,I1333425,I994164);
not I_78289 (I1333459,I994164);
and I_78290 (I1333476,I1333459,I994170);
nand I_78291 (I1333493,I1333476,I994182);
nor I_78292 (I1333510,I1333459,I1333493);
DFFARX1 I_78293 (I1333510,I2507,I1333312,I1333277,);
not I_78294 (I1333541,I1333493);
nand I_78295 (I1333558,I1333363,I1333541);
nand I_78296 (I1333289,I1333425,I1333541);
DFFARX1 I_78297 (I1333459,I2507,I1333312,I1333304,);
not I_78298 (I1333603,I994173);
nor I_78299 (I1333620,I1333603,I994170);
nor I_78300 (I1333637,I1333620,I1333442);
DFFARX1 I_78301 (I1333637,I2507,I1333312,I1333301,);
not I_78302 (I1333668,I1333620);
DFFARX1 I_78303 (I1333668,I2507,I1333312,I1333694,);
not I_78304 (I1333702,I1333694);
nor I_78305 (I1333298,I1333702,I1333620);
nor I_78306 (I1333733,I1333603,I994161);
and I_78307 (I1333750,I1333733,I994188);
or I_78308 (I1333767,I1333750,I994179);
DFFARX1 I_78309 (I1333767,I2507,I1333312,I1333793,);
not I_78310 (I1333801,I1333793);
nand I_78311 (I1333818,I1333801,I1333541);
not I_78312 (I1333292,I1333818);
nand I_78313 (I1333286,I1333818,I1333558);
nand I_78314 (I1333283,I1333801,I1333425);
not I_78315 (I1333907,I2514);
DFFARX1 I_78316 (I900497,I2507,I1333907,I1333933,);
DFFARX1 I_78317 (I900515,I2507,I1333907,I1333950,);
not I_78318 (I1333958,I1333950);
nor I_78319 (I1333875,I1333933,I1333958);
DFFARX1 I_78320 (I1333958,I2507,I1333907,I1333890,);
nor I_78321 (I1334003,I900494,I900506);
and I_78322 (I1334020,I1334003,I900491);
nor I_78323 (I1334037,I1334020,I900494);
not I_78324 (I1334054,I900494);
and I_78325 (I1334071,I1334054,I900500);
nand I_78326 (I1334088,I1334071,I900512);
nor I_78327 (I1334105,I1334054,I1334088);
DFFARX1 I_78328 (I1334105,I2507,I1333907,I1333872,);
not I_78329 (I1334136,I1334088);
nand I_78330 (I1334153,I1333958,I1334136);
nand I_78331 (I1333884,I1334020,I1334136);
DFFARX1 I_78332 (I1334054,I2507,I1333907,I1333899,);
not I_78333 (I1334198,I900503);
nor I_78334 (I1334215,I1334198,I900500);
nor I_78335 (I1334232,I1334215,I1334037);
DFFARX1 I_78336 (I1334232,I2507,I1333907,I1333896,);
not I_78337 (I1334263,I1334215);
DFFARX1 I_78338 (I1334263,I2507,I1333907,I1334289,);
not I_78339 (I1334297,I1334289);
nor I_78340 (I1333893,I1334297,I1334215);
nor I_78341 (I1334328,I1334198,I900491);
and I_78342 (I1334345,I1334328,I900518);
or I_78343 (I1334362,I1334345,I900509);
DFFARX1 I_78344 (I1334362,I2507,I1333907,I1334388,);
not I_78345 (I1334396,I1334388);
nand I_78346 (I1334413,I1334396,I1334136);
not I_78347 (I1333887,I1334413);
nand I_78348 (I1333881,I1334413,I1334153);
nand I_78349 (I1333878,I1334396,I1334020);
not I_78350 (I1334502,I2514);
DFFARX1 I_78351 (I232935,I2507,I1334502,I1334528,);
DFFARX1 I_78352 (I232938,I2507,I1334502,I1334545,);
not I_78353 (I1334553,I1334545);
nor I_78354 (I1334470,I1334528,I1334553);
DFFARX1 I_78355 (I1334553,I2507,I1334502,I1334485,);
nor I_78356 (I1334598,I232944,I232938);
and I_78357 (I1334615,I1334598,I232941);
nor I_78358 (I1334632,I1334615,I232944);
not I_78359 (I1334649,I232944);
and I_78360 (I1334666,I1334649,I232935);
nand I_78361 (I1334683,I1334666,I232953);
nor I_78362 (I1334700,I1334649,I1334683);
DFFARX1 I_78363 (I1334700,I2507,I1334502,I1334467,);
not I_78364 (I1334731,I1334683);
nand I_78365 (I1334748,I1334553,I1334731);
nand I_78366 (I1334479,I1334615,I1334731);
DFFARX1 I_78367 (I1334649,I2507,I1334502,I1334494,);
not I_78368 (I1334793,I232947);
nor I_78369 (I1334810,I1334793,I232935);
nor I_78370 (I1334827,I1334810,I1334632);
DFFARX1 I_78371 (I1334827,I2507,I1334502,I1334491,);
not I_78372 (I1334858,I1334810);
DFFARX1 I_78373 (I1334858,I2507,I1334502,I1334884,);
not I_78374 (I1334892,I1334884);
nor I_78375 (I1334488,I1334892,I1334810);
nor I_78376 (I1334923,I1334793,I232950);
and I_78377 (I1334940,I1334923,I232956);
or I_78378 (I1334957,I1334940,I232959);
DFFARX1 I_78379 (I1334957,I2507,I1334502,I1334983,);
not I_78380 (I1334991,I1334983);
nand I_78381 (I1335008,I1334991,I1334731);
not I_78382 (I1334482,I1335008);
nand I_78383 (I1334476,I1335008,I1334748);
nand I_78384 (I1334473,I1334991,I1334615);
not I_78385 (I1335097,I2514);
DFFARX1 I_78386 (I707613,I2507,I1335097,I1335123,);
DFFARX1 I_78387 (I707595,I2507,I1335097,I1335140,);
not I_78388 (I1335148,I1335140);
nor I_78389 (I1335065,I1335123,I1335148);
DFFARX1 I_78390 (I1335148,I2507,I1335097,I1335080,);
nor I_78391 (I1335193,I707601,I707604);
and I_78392 (I1335210,I1335193,I707592);
nor I_78393 (I1335227,I1335210,I707601);
not I_78394 (I1335244,I707601);
and I_78395 (I1335261,I1335244,I707610);
nand I_78396 (I1335278,I1335261,I707598);
nor I_78397 (I1335295,I1335244,I1335278);
DFFARX1 I_78398 (I1335295,I2507,I1335097,I1335062,);
not I_78399 (I1335326,I1335278);
nand I_78400 (I1335343,I1335148,I1335326);
nand I_78401 (I1335074,I1335210,I1335326);
DFFARX1 I_78402 (I1335244,I2507,I1335097,I1335089,);
not I_78403 (I1335388,I707595);
nor I_78404 (I1335405,I1335388,I707610);
nor I_78405 (I1335422,I1335405,I1335227);
DFFARX1 I_78406 (I1335422,I2507,I1335097,I1335086,);
not I_78407 (I1335453,I1335405);
DFFARX1 I_78408 (I1335453,I2507,I1335097,I1335479,);
not I_78409 (I1335487,I1335479);
nor I_78410 (I1335083,I1335487,I1335405);
nor I_78411 (I1335518,I1335388,I707607);
and I_78412 (I1335535,I1335518,I707616);
or I_78413 (I1335552,I1335535,I707592);
DFFARX1 I_78414 (I1335552,I2507,I1335097,I1335578,);
not I_78415 (I1335586,I1335578);
nand I_78416 (I1335603,I1335586,I1335326);
not I_78417 (I1335077,I1335603);
nand I_78418 (I1335071,I1335603,I1335343);
nand I_78419 (I1335068,I1335586,I1335210);
not I_78420 (I1335692,I2514);
DFFARX1 I_78421 (I277615,I2507,I1335692,I1335718,);
DFFARX1 I_78422 (I277609,I2507,I1335692,I1335735,);
not I_78423 (I1335743,I1335735);
nor I_78424 (I1335660,I1335718,I1335743);
DFFARX1 I_78425 (I1335743,I2507,I1335692,I1335675,);
nor I_78426 (I1335788,I277597,I277618);
and I_78427 (I1335805,I1335788,I277612);
nor I_78428 (I1335822,I1335805,I277597);
not I_78429 (I1335839,I277597);
and I_78430 (I1335856,I1335839,I277594);
nand I_78431 (I1335873,I1335856,I277606);
nor I_78432 (I1335890,I1335839,I1335873);
DFFARX1 I_78433 (I1335890,I2507,I1335692,I1335657,);
not I_78434 (I1335921,I1335873);
nand I_78435 (I1335938,I1335743,I1335921);
nand I_78436 (I1335669,I1335805,I1335921);
DFFARX1 I_78437 (I1335839,I2507,I1335692,I1335684,);
not I_78438 (I1335983,I277621);
nor I_78439 (I1336000,I1335983,I277594);
nor I_78440 (I1336017,I1336000,I1335822);
DFFARX1 I_78441 (I1336017,I2507,I1335692,I1335681,);
not I_78442 (I1336048,I1336000);
DFFARX1 I_78443 (I1336048,I2507,I1335692,I1336074,);
not I_78444 (I1336082,I1336074);
nor I_78445 (I1335678,I1336082,I1336000);
nor I_78446 (I1336113,I1335983,I277603);
and I_78447 (I1336130,I1336113,I277600);
or I_78448 (I1336147,I1336130,I277594);
DFFARX1 I_78449 (I1336147,I2507,I1335692,I1336173,);
not I_78450 (I1336181,I1336173);
nand I_78451 (I1336198,I1336181,I1335921);
not I_78452 (I1335672,I1336198);
nand I_78453 (I1335666,I1336198,I1335938);
nand I_78454 (I1335663,I1336181,I1335805);
not I_78455 (I1336287,I2514);
DFFARX1 I_78456 (I421839,I2507,I1336287,I1336313,);
DFFARX1 I_78457 (I421845,I2507,I1336287,I1336330,);
not I_78458 (I1336338,I1336330);
nor I_78459 (I1336255,I1336313,I1336338);
DFFARX1 I_78460 (I1336338,I2507,I1336287,I1336270,);
nor I_78461 (I1336383,I421854,I421839);
and I_78462 (I1336400,I1336383,I421866);
nor I_78463 (I1336417,I1336400,I421854);
not I_78464 (I1336434,I421854);
and I_78465 (I1336451,I1336434,I421842);
nand I_78466 (I1336468,I1336451,I421863);
nor I_78467 (I1336485,I1336434,I1336468);
DFFARX1 I_78468 (I1336485,I2507,I1336287,I1336252,);
not I_78469 (I1336516,I1336468);
nand I_78470 (I1336533,I1336338,I1336516);
nand I_78471 (I1336264,I1336400,I1336516);
DFFARX1 I_78472 (I1336434,I2507,I1336287,I1336279,);
not I_78473 (I1336578,I421851);
nor I_78474 (I1336595,I1336578,I421842);
nor I_78475 (I1336612,I1336595,I1336417);
DFFARX1 I_78476 (I1336612,I2507,I1336287,I1336276,);
not I_78477 (I1336643,I1336595);
DFFARX1 I_78478 (I1336643,I2507,I1336287,I1336669,);
not I_78479 (I1336677,I1336669);
nor I_78480 (I1336273,I1336677,I1336595);
nor I_78481 (I1336708,I1336578,I421848);
and I_78482 (I1336725,I1336708,I421860);
or I_78483 (I1336742,I1336725,I421857);
DFFARX1 I_78484 (I1336742,I2507,I1336287,I1336768,);
not I_78485 (I1336776,I1336768);
nand I_78486 (I1336793,I1336776,I1336516);
not I_78487 (I1336267,I1336793);
nand I_78488 (I1336261,I1336793,I1336533);
nand I_78489 (I1336258,I1336776,I1336400);
not I_78490 (I1336882,I2514);
DFFARX1 I_78491 (I320302,I2507,I1336882,I1336908,);
DFFARX1 I_78492 (I320296,I2507,I1336882,I1336925,);
not I_78493 (I1336933,I1336925);
nor I_78494 (I1336850,I1336908,I1336933);
DFFARX1 I_78495 (I1336933,I2507,I1336882,I1336865,);
nor I_78496 (I1336978,I320284,I320305);
and I_78497 (I1336995,I1336978,I320299);
nor I_78498 (I1337012,I1336995,I320284);
not I_78499 (I1337029,I320284);
and I_78500 (I1337046,I1337029,I320281);
nand I_78501 (I1337063,I1337046,I320293);
nor I_78502 (I1337080,I1337029,I1337063);
DFFARX1 I_78503 (I1337080,I2507,I1336882,I1336847,);
not I_78504 (I1337111,I1337063);
nand I_78505 (I1337128,I1336933,I1337111);
nand I_78506 (I1336859,I1336995,I1337111);
DFFARX1 I_78507 (I1337029,I2507,I1336882,I1336874,);
not I_78508 (I1337173,I320308);
nor I_78509 (I1337190,I1337173,I320281);
nor I_78510 (I1337207,I1337190,I1337012);
DFFARX1 I_78511 (I1337207,I2507,I1336882,I1336871,);
not I_78512 (I1337238,I1337190);
DFFARX1 I_78513 (I1337238,I2507,I1336882,I1337264,);
not I_78514 (I1337272,I1337264);
nor I_78515 (I1336868,I1337272,I1337190);
nor I_78516 (I1337303,I1337173,I320290);
and I_78517 (I1337320,I1337303,I320287);
or I_78518 (I1337337,I1337320,I320281);
DFFARX1 I_78519 (I1337337,I2507,I1336882,I1337363,);
not I_78520 (I1337371,I1337363);
nand I_78521 (I1337388,I1337371,I1337111);
not I_78522 (I1336862,I1337388);
nand I_78523 (I1336856,I1337388,I1337128);
nand I_78524 (I1336853,I1337371,I1336995);
not I_78525 (I1337477,I2514);
DFFARX1 I_78526 (I868659,I2507,I1337477,I1337503,);
DFFARX1 I_78527 (I868656,I2507,I1337477,I1337520,);
not I_78528 (I1337528,I1337520);
nor I_78529 (I1337445,I1337503,I1337528);
DFFARX1 I_78530 (I1337528,I2507,I1337477,I1337460,);
nor I_78531 (I1337573,I868671,I868653);
and I_78532 (I1337590,I1337573,I868650);
nor I_78533 (I1337607,I1337590,I868671);
not I_78534 (I1337624,I868671);
and I_78535 (I1337641,I1337624,I868656);
nand I_78536 (I1337658,I1337641,I868668);
nor I_78537 (I1337675,I1337624,I1337658);
DFFARX1 I_78538 (I1337675,I2507,I1337477,I1337442,);
not I_78539 (I1337706,I1337658);
nand I_78540 (I1337723,I1337528,I1337706);
nand I_78541 (I1337454,I1337590,I1337706);
DFFARX1 I_78542 (I1337624,I2507,I1337477,I1337469,);
not I_78543 (I1337768,I868662);
nor I_78544 (I1337785,I1337768,I868656);
nor I_78545 (I1337802,I1337785,I1337607);
DFFARX1 I_78546 (I1337802,I2507,I1337477,I1337466,);
not I_78547 (I1337833,I1337785);
DFFARX1 I_78548 (I1337833,I2507,I1337477,I1337859,);
not I_78549 (I1337867,I1337859);
nor I_78550 (I1337463,I1337867,I1337785);
nor I_78551 (I1337898,I1337768,I868650);
and I_78552 (I1337915,I1337898,I868665);
or I_78553 (I1337932,I1337915,I868653);
DFFARX1 I_78554 (I1337932,I2507,I1337477,I1337958,);
not I_78555 (I1337966,I1337958);
nand I_78556 (I1337983,I1337966,I1337706);
not I_78557 (I1337457,I1337983);
nand I_78558 (I1337451,I1337983,I1337723);
nand I_78559 (I1337448,I1337966,I1337590);
not I_78560 (I1338072,I2514);
DFFARX1 I_78561 (I195450,I2507,I1338072,I1338098,);
DFFARX1 I_78562 (I195453,I2507,I1338072,I1338115,);
not I_78563 (I1338123,I1338115);
nor I_78564 (I1338040,I1338098,I1338123);
DFFARX1 I_78565 (I1338123,I2507,I1338072,I1338055,);
nor I_78566 (I1338168,I195459,I195453);
and I_78567 (I1338185,I1338168,I195456);
nor I_78568 (I1338202,I1338185,I195459);
not I_78569 (I1338219,I195459);
and I_78570 (I1338236,I1338219,I195450);
nand I_78571 (I1338253,I1338236,I195468);
nor I_78572 (I1338270,I1338219,I1338253);
DFFARX1 I_78573 (I1338270,I2507,I1338072,I1338037,);
not I_78574 (I1338301,I1338253);
nand I_78575 (I1338318,I1338123,I1338301);
nand I_78576 (I1338049,I1338185,I1338301);
DFFARX1 I_78577 (I1338219,I2507,I1338072,I1338064,);
not I_78578 (I1338363,I195462);
nor I_78579 (I1338380,I1338363,I195450);
nor I_78580 (I1338397,I1338380,I1338202);
DFFARX1 I_78581 (I1338397,I2507,I1338072,I1338061,);
not I_78582 (I1338428,I1338380);
DFFARX1 I_78583 (I1338428,I2507,I1338072,I1338454,);
not I_78584 (I1338462,I1338454);
nor I_78585 (I1338058,I1338462,I1338380);
nor I_78586 (I1338493,I1338363,I195465);
and I_78587 (I1338510,I1338493,I195471);
or I_78588 (I1338527,I1338510,I195474);
DFFARX1 I_78589 (I1338527,I2507,I1338072,I1338553,);
not I_78590 (I1338561,I1338553);
nand I_78591 (I1338578,I1338561,I1338301);
not I_78592 (I1338052,I1338578);
nand I_78593 (I1338046,I1338578,I1338318);
nand I_78594 (I1338043,I1338561,I1338185);
not I_78595 (I1338667,I2514);
DFFARX1 I_78596 (I993521,I2507,I1338667,I1338693,);
DFFARX1 I_78597 (I993539,I2507,I1338667,I1338710,);
not I_78598 (I1338718,I1338710);
nor I_78599 (I1338635,I1338693,I1338718);
DFFARX1 I_78600 (I1338718,I2507,I1338667,I1338650,);
nor I_78601 (I1338763,I993518,I993530);
and I_78602 (I1338780,I1338763,I993515);
nor I_78603 (I1338797,I1338780,I993518);
not I_78604 (I1338814,I993518);
and I_78605 (I1338831,I1338814,I993524);
nand I_78606 (I1338848,I1338831,I993536);
nor I_78607 (I1338865,I1338814,I1338848);
DFFARX1 I_78608 (I1338865,I2507,I1338667,I1338632,);
not I_78609 (I1338896,I1338848);
nand I_78610 (I1338913,I1338718,I1338896);
nand I_78611 (I1338644,I1338780,I1338896);
DFFARX1 I_78612 (I1338814,I2507,I1338667,I1338659,);
not I_78613 (I1338958,I993527);
nor I_78614 (I1338975,I1338958,I993524);
nor I_78615 (I1338992,I1338975,I1338797);
DFFARX1 I_78616 (I1338992,I2507,I1338667,I1338656,);
not I_78617 (I1339023,I1338975);
DFFARX1 I_78618 (I1339023,I2507,I1338667,I1339049,);
not I_78619 (I1339057,I1339049);
nor I_78620 (I1338653,I1339057,I1338975);
nor I_78621 (I1339088,I1338958,I993515);
and I_78622 (I1339105,I1339088,I993542);
or I_78623 (I1339122,I1339105,I993533);
DFFARX1 I_78624 (I1339122,I2507,I1338667,I1339148,);
not I_78625 (I1339156,I1339148);
nand I_78626 (I1339173,I1339156,I1338896);
not I_78627 (I1338647,I1339173);
nand I_78628 (I1338641,I1339173,I1338913);
nand I_78629 (I1338638,I1339156,I1338780);
not I_78630 (I1339262,I2514);
DFFARX1 I_78631 (I642877,I2507,I1339262,I1339288,);
DFFARX1 I_78632 (I642859,I2507,I1339262,I1339305,);
not I_78633 (I1339313,I1339305);
nor I_78634 (I1339230,I1339288,I1339313);
DFFARX1 I_78635 (I1339313,I2507,I1339262,I1339245,);
nor I_78636 (I1339358,I642865,I642868);
and I_78637 (I1339375,I1339358,I642856);
nor I_78638 (I1339392,I1339375,I642865);
not I_78639 (I1339409,I642865);
and I_78640 (I1339426,I1339409,I642874);
nand I_78641 (I1339443,I1339426,I642862);
nor I_78642 (I1339460,I1339409,I1339443);
DFFARX1 I_78643 (I1339460,I2507,I1339262,I1339227,);
not I_78644 (I1339491,I1339443);
nand I_78645 (I1339508,I1339313,I1339491);
nand I_78646 (I1339239,I1339375,I1339491);
DFFARX1 I_78647 (I1339409,I2507,I1339262,I1339254,);
not I_78648 (I1339553,I642859);
nor I_78649 (I1339570,I1339553,I642874);
nor I_78650 (I1339587,I1339570,I1339392);
DFFARX1 I_78651 (I1339587,I2507,I1339262,I1339251,);
not I_78652 (I1339618,I1339570);
DFFARX1 I_78653 (I1339618,I2507,I1339262,I1339644,);
not I_78654 (I1339652,I1339644);
nor I_78655 (I1339248,I1339652,I1339570);
nor I_78656 (I1339683,I1339553,I642871);
and I_78657 (I1339700,I1339683,I642880);
or I_78658 (I1339717,I1339700,I642856);
DFFARX1 I_78659 (I1339717,I2507,I1339262,I1339743,);
not I_78660 (I1339751,I1339743);
nand I_78661 (I1339768,I1339751,I1339491);
not I_78662 (I1339242,I1339768);
nand I_78663 (I1339236,I1339768,I1339508);
nand I_78664 (I1339233,I1339751,I1339375);
not I_78665 (I1339857,I2514);
DFFARX1 I_78666 (I808054,I2507,I1339857,I1339883,);
DFFARX1 I_78667 (I808051,I2507,I1339857,I1339900,);
not I_78668 (I1339908,I1339900);
nor I_78669 (I1339825,I1339883,I1339908);
DFFARX1 I_78670 (I1339908,I2507,I1339857,I1339840,);
nor I_78671 (I1339953,I808066,I808048);
and I_78672 (I1339970,I1339953,I808045);
nor I_78673 (I1339987,I1339970,I808066);
not I_78674 (I1340004,I808066);
and I_78675 (I1340021,I1340004,I808051);
nand I_78676 (I1340038,I1340021,I808063);
nor I_78677 (I1340055,I1340004,I1340038);
DFFARX1 I_78678 (I1340055,I2507,I1339857,I1339822,);
not I_78679 (I1340086,I1340038);
nand I_78680 (I1340103,I1339908,I1340086);
nand I_78681 (I1339834,I1339970,I1340086);
DFFARX1 I_78682 (I1340004,I2507,I1339857,I1339849,);
not I_78683 (I1340148,I808057);
nor I_78684 (I1340165,I1340148,I808051);
nor I_78685 (I1340182,I1340165,I1339987);
DFFARX1 I_78686 (I1340182,I2507,I1339857,I1339846,);
not I_78687 (I1340213,I1340165);
DFFARX1 I_78688 (I1340213,I2507,I1339857,I1340239,);
not I_78689 (I1340247,I1340239);
nor I_78690 (I1339843,I1340247,I1340165);
nor I_78691 (I1340278,I1340148,I808045);
and I_78692 (I1340295,I1340278,I808060);
or I_78693 (I1340312,I1340295,I808048);
DFFARX1 I_78694 (I1340312,I2507,I1339857,I1340338,);
not I_78695 (I1340346,I1340338);
nand I_78696 (I1340363,I1340346,I1340086);
not I_78697 (I1339837,I1340363);
nand I_78698 (I1339831,I1340363,I1340103);
nand I_78699 (I1339828,I1340346,I1339970);
not I_78700 (I1340452,I2514);
DFFARX1 I_78701 (I1051106,I2507,I1340452,I1340478,);
DFFARX1 I_78702 (I1051097,I2507,I1340452,I1340495,);
not I_78703 (I1340503,I1340495);
nor I_78704 (I1340420,I1340478,I1340503);
DFFARX1 I_78705 (I1340503,I2507,I1340452,I1340435,);
nor I_78706 (I1340548,I1051103,I1051112);
and I_78707 (I1340565,I1340548,I1051115);
nor I_78708 (I1340582,I1340565,I1051103);
not I_78709 (I1340599,I1051103);
and I_78710 (I1340616,I1340599,I1051094);
nand I_78711 (I1340633,I1340616,I1051100);
nor I_78712 (I1340650,I1340599,I1340633);
DFFARX1 I_78713 (I1340650,I2507,I1340452,I1340417,);
not I_78714 (I1340681,I1340633);
nand I_78715 (I1340698,I1340503,I1340681);
nand I_78716 (I1340429,I1340565,I1340681);
DFFARX1 I_78717 (I1340599,I2507,I1340452,I1340444,);
not I_78718 (I1340743,I1051109);
nor I_78719 (I1340760,I1340743,I1051094);
nor I_78720 (I1340777,I1340760,I1340582);
DFFARX1 I_78721 (I1340777,I2507,I1340452,I1340441,);
not I_78722 (I1340808,I1340760);
DFFARX1 I_78723 (I1340808,I2507,I1340452,I1340834,);
not I_78724 (I1340842,I1340834);
nor I_78725 (I1340438,I1340842,I1340760);
nor I_78726 (I1340873,I1340743,I1051094);
and I_78727 (I1340890,I1340873,I1051097);
or I_78728 (I1340907,I1340890,I1051100);
DFFARX1 I_78729 (I1340907,I2507,I1340452,I1340933,);
not I_78730 (I1340941,I1340933);
nand I_78731 (I1340958,I1340941,I1340681);
not I_78732 (I1340432,I1340958);
nand I_78733 (I1340426,I1340958,I1340698);
nand I_78734 (I1340423,I1340941,I1340565);
not I_78735 (I1341047,I2514);
DFFARX1 I_78736 (I81758,I2507,I1341047,I1341073,);
DFFARX1 I_78737 (I81746,I2507,I1341047,I1341090,);
not I_78738 (I1341098,I1341090);
nor I_78739 (I1341015,I1341073,I1341098);
DFFARX1 I_78740 (I1341098,I2507,I1341047,I1341030,);
nor I_78741 (I1341143,I81737,I81761);
and I_78742 (I1341160,I1341143,I81740);
nor I_78743 (I1341177,I1341160,I81737);
not I_78744 (I1341194,I81737);
and I_78745 (I1341211,I1341194,I81743);
nand I_78746 (I1341228,I1341211,I81755);
nor I_78747 (I1341245,I1341194,I1341228);
DFFARX1 I_78748 (I1341245,I2507,I1341047,I1341012,);
not I_78749 (I1341276,I1341228);
nand I_78750 (I1341293,I1341098,I1341276);
nand I_78751 (I1341024,I1341160,I1341276);
DFFARX1 I_78752 (I1341194,I2507,I1341047,I1341039,);
not I_78753 (I1341338,I81737);
nor I_78754 (I1341355,I1341338,I81743);
nor I_78755 (I1341372,I1341355,I1341177);
DFFARX1 I_78756 (I1341372,I2507,I1341047,I1341036,);
not I_78757 (I1341403,I1341355);
DFFARX1 I_78758 (I1341403,I2507,I1341047,I1341429,);
not I_78759 (I1341437,I1341429);
nor I_78760 (I1341033,I1341437,I1341355);
nor I_78761 (I1341468,I1341338,I81740);
and I_78762 (I1341485,I1341468,I81749);
or I_78763 (I1341502,I1341485,I81752);
DFFARX1 I_78764 (I1341502,I2507,I1341047,I1341528,);
not I_78765 (I1341536,I1341528);
nand I_78766 (I1341553,I1341536,I1341276);
not I_78767 (I1341027,I1341553);
nand I_78768 (I1341021,I1341553,I1341293);
nand I_78769 (I1341018,I1341536,I1341160);
not I_78770 (I1341642,I2514);
DFFARX1 I_78771 (I1001273,I2507,I1341642,I1341668,);
DFFARX1 I_78772 (I1001291,I2507,I1341642,I1341685,);
not I_78773 (I1341693,I1341685);
nor I_78774 (I1341610,I1341668,I1341693);
DFFARX1 I_78775 (I1341693,I2507,I1341642,I1341625,);
nor I_78776 (I1341738,I1001270,I1001282);
and I_78777 (I1341755,I1341738,I1001267);
nor I_78778 (I1341772,I1341755,I1001270);
not I_78779 (I1341789,I1001270);
and I_78780 (I1341806,I1341789,I1001276);
nand I_78781 (I1341823,I1341806,I1001288);
nor I_78782 (I1341840,I1341789,I1341823);
DFFARX1 I_78783 (I1341840,I2507,I1341642,I1341607,);
not I_78784 (I1341871,I1341823);
nand I_78785 (I1341888,I1341693,I1341871);
nand I_78786 (I1341619,I1341755,I1341871);
DFFARX1 I_78787 (I1341789,I2507,I1341642,I1341634,);
not I_78788 (I1341933,I1001279);
nor I_78789 (I1341950,I1341933,I1001276);
nor I_78790 (I1341967,I1341950,I1341772);
DFFARX1 I_78791 (I1341967,I2507,I1341642,I1341631,);
not I_78792 (I1341998,I1341950);
DFFARX1 I_78793 (I1341998,I2507,I1341642,I1342024,);
not I_78794 (I1342032,I1342024);
nor I_78795 (I1341628,I1342032,I1341950);
nor I_78796 (I1342063,I1341933,I1001267);
and I_78797 (I1342080,I1342063,I1001294);
or I_78798 (I1342097,I1342080,I1001285);
DFFARX1 I_78799 (I1342097,I2507,I1341642,I1342123,);
not I_78800 (I1342131,I1342123);
nand I_78801 (I1342148,I1342131,I1341871);
not I_78802 (I1341622,I1342148);
nand I_78803 (I1341616,I1342148,I1341888);
nand I_78804 (I1341613,I1342131,I1341755);
not I_78805 (I1342237,I2514);
DFFARX1 I_78806 (I672933,I2507,I1342237,I1342263,);
DFFARX1 I_78807 (I672915,I2507,I1342237,I1342280,);
not I_78808 (I1342288,I1342280);
nor I_78809 (I1342205,I1342263,I1342288);
DFFARX1 I_78810 (I1342288,I2507,I1342237,I1342220,);
nor I_78811 (I1342333,I672921,I672924);
and I_78812 (I1342350,I1342333,I672912);
nor I_78813 (I1342367,I1342350,I672921);
not I_78814 (I1342384,I672921);
and I_78815 (I1342401,I1342384,I672930);
nand I_78816 (I1342418,I1342401,I672918);
nor I_78817 (I1342435,I1342384,I1342418);
DFFARX1 I_78818 (I1342435,I2507,I1342237,I1342202,);
not I_78819 (I1342466,I1342418);
nand I_78820 (I1342483,I1342288,I1342466);
nand I_78821 (I1342214,I1342350,I1342466);
DFFARX1 I_78822 (I1342384,I2507,I1342237,I1342229,);
not I_78823 (I1342528,I672915);
nor I_78824 (I1342545,I1342528,I672930);
nor I_78825 (I1342562,I1342545,I1342367);
DFFARX1 I_78826 (I1342562,I2507,I1342237,I1342226,);
not I_78827 (I1342593,I1342545);
DFFARX1 I_78828 (I1342593,I2507,I1342237,I1342619,);
not I_78829 (I1342627,I1342619);
nor I_78830 (I1342223,I1342627,I1342545);
nor I_78831 (I1342658,I1342528,I672927);
and I_78832 (I1342675,I1342658,I672936);
or I_78833 (I1342692,I1342675,I672912);
DFFARX1 I_78834 (I1342692,I2507,I1342237,I1342718,);
not I_78835 (I1342726,I1342718);
nand I_78836 (I1342743,I1342726,I1342466);
not I_78837 (I1342217,I1342743);
nand I_78838 (I1342211,I1342743,I1342483);
nand I_78839 (I1342208,I1342726,I1342350);
not I_78840 (I1342832,I2514);
DFFARX1 I_78841 (I141329,I2507,I1342832,I1342858,);
DFFARX1 I_78842 (I141305,I2507,I1342832,I1342875,);
not I_78843 (I1342883,I1342875);
nor I_78844 (I1342800,I1342858,I1342883);
DFFARX1 I_78845 (I1342883,I2507,I1342832,I1342815,);
nor I_78846 (I1342928,I141332,I141314);
and I_78847 (I1342945,I1342928,I141326);
nor I_78848 (I1342962,I1342945,I141332);
not I_78849 (I1342979,I141332);
and I_78850 (I1342996,I1342979,I141308);
nand I_78851 (I1343013,I1342996,I141323);
nor I_78852 (I1343030,I1342979,I1343013);
DFFARX1 I_78853 (I1343030,I2507,I1342832,I1342797,);
not I_78854 (I1343061,I1343013);
nand I_78855 (I1343078,I1342883,I1343061);
nand I_78856 (I1342809,I1342945,I1343061);
DFFARX1 I_78857 (I1342979,I2507,I1342832,I1342824,);
not I_78858 (I1343123,I141317);
nor I_78859 (I1343140,I1343123,I141308);
nor I_78860 (I1343157,I1343140,I1342962);
DFFARX1 I_78861 (I1343157,I2507,I1342832,I1342821,);
not I_78862 (I1343188,I1343140);
DFFARX1 I_78863 (I1343188,I2507,I1342832,I1343214,);
not I_78864 (I1343222,I1343214);
nor I_78865 (I1342818,I1343222,I1343140);
nor I_78866 (I1343253,I1343123,I141320);
and I_78867 (I1343270,I1343253,I141311);
or I_78868 (I1343287,I1343270,I141305);
DFFARX1 I_78869 (I1343287,I2507,I1342832,I1343313,);
not I_78870 (I1343321,I1343313);
nand I_78871 (I1343338,I1343321,I1343061);
not I_78872 (I1342812,I1343338);
nand I_78873 (I1342806,I1343338,I1343078);
nand I_78874 (I1342803,I1343321,I1342945);
not I_78875 (I1343427,I2514);
DFFARX1 I_78876 (I1113861,I2507,I1343427,I1343453,);
DFFARX1 I_78877 (I1113873,I2507,I1343427,I1343470,);
not I_78878 (I1343478,I1343470);
nor I_78879 (I1343395,I1343453,I1343478);
DFFARX1 I_78880 (I1343478,I2507,I1343427,I1343410,);
nor I_78881 (I1343523,I1113870,I1113864);
and I_78882 (I1343540,I1343523,I1113858);
nor I_78883 (I1343557,I1343540,I1113870);
not I_78884 (I1343574,I1113870);
and I_78885 (I1343591,I1343574,I1113867);
nand I_78886 (I1343608,I1343591,I1113858);
nor I_78887 (I1343625,I1343574,I1343608);
DFFARX1 I_78888 (I1343625,I2507,I1343427,I1343392,);
not I_78889 (I1343656,I1343608);
nand I_78890 (I1343673,I1343478,I1343656);
nand I_78891 (I1343404,I1343540,I1343656);
DFFARX1 I_78892 (I1343574,I2507,I1343427,I1343419,);
not I_78893 (I1343718,I1113882);
nor I_78894 (I1343735,I1343718,I1113867);
nor I_78895 (I1343752,I1343735,I1343557);
DFFARX1 I_78896 (I1343752,I2507,I1343427,I1343416,);
not I_78897 (I1343783,I1343735);
DFFARX1 I_78898 (I1343783,I2507,I1343427,I1343809,);
not I_78899 (I1343817,I1343809);
nor I_78900 (I1343413,I1343817,I1343735);
nor I_78901 (I1343848,I1343718,I1113876);
and I_78902 (I1343865,I1343848,I1113879);
or I_78903 (I1343882,I1343865,I1113861);
DFFARX1 I_78904 (I1343882,I2507,I1343427,I1343908,);
not I_78905 (I1343916,I1343908);
nand I_78906 (I1343933,I1343916,I1343656);
not I_78907 (I1343407,I1343933);
nand I_78908 (I1343401,I1343933,I1343673);
nand I_78909 (I1343398,I1343916,I1343540);
not I_78910 (I1344022,I2514);
DFFARX1 I_78911 (I1224834,I2507,I1344022,I1344048,);
DFFARX1 I_78912 (I1224837,I2507,I1344022,I1344065,);
not I_78913 (I1344073,I1344065);
nor I_78914 (I1343990,I1344048,I1344073);
DFFARX1 I_78915 (I1344073,I2507,I1344022,I1344005,);
nor I_78916 (I1344118,I1224837,I1224852);
and I_78917 (I1344135,I1344118,I1224846);
nor I_78918 (I1344152,I1344135,I1224837);
not I_78919 (I1344169,I1224837);
and I_78920 (I1344186,I1344169,I1224855);
nand I_78921 (I1344203,I1344186,I1224843);
nor I_78922 (I1344220,I1344169,I1344203);
DFFARX1 I_78923 (I1344220,I2507,I1344022,I1343987,);
not I_78924 (I1344251,I1344203);
nand I_78925 (I1344268,I1344073,I1344251);
nand I_78926 (I1343999,I1344135,I1344251);
DFFARX1 I_78927 (I1344169,I2507,I1344022,I1344014,);
not I_78928 (I1344313,I1224849);
nor I_78929 (I1344330,I1344313,I1224855);
nor I_78930 (I1344347,I1344330,I1344152);
DFFARX1 I_78931 (I1344347,I2507,I1344022,I1344011,);
not I_78932 (I1344378,I1344330);
DFFARX1 I_78933 (I1344378,I2507,I1344022,I1344404,);
not I_78934 (I1344412,I1344404);
nor I_78935 (I1344008,I1344412,I1344330);
nor I_78936 (I1344443,I1344313,I1224834);
and I_78937 (I1344460,I1344443,I1224858);
or I_78938 (I1344477,I1344460,I1224840);
DFFARX1 I_78939 (I1344477,I2507,I1344022,I1344503,);
not I_78940 (I1344511,I1344503);
nand I_78941 (I1344528,I1344511,I1344251);
not I_78942 (I1344002,I1344528);
nand I_78943 (I1343996,I1344528,I1344268);
nand I_78944 (I1343993,I1344511,I1344135);
not I_78945 (I1344617,I2514);
DFFARX1 I_78946 (I502419,I2507,I1344617,I1344643,);
DFFARX1 I_78947 (I502422,I2507,I1344617,I1344660,);
not I_78948 (I1344668,I1344660);
nor I_78949 (I1344585,I1344643,I1344668);
DFFARX1 I_78950 (I1344668,I2507,I1344617,I1344600,);
nor I_78951 (I1344713,I502425,I502443);
and I_78952 (I1344730,I1344713,I502428);
nor I_78953 (I1344747,I1344730,I502425);
not I_78954 (I1344764,I502425);
and I_78955 (I1344781,I1344764,I502437);
nand I_78956 (I1344798,I1344781,I502440);
nor I_78957 (I1344815,I1344764,I1344798);
DFFARX1 I_78958 (I1344815,I2507,I1344617,I1344582,);
not I_78959 (I1344846,I1344798);
nand I_78960 (I1344863,I1344668,I1344846);
nand I_78961 (I1344594,I1344730,I1344846);
DFFARX1 I_78962 (I1344764,I2507,I1344617,I1344609,);
not I_78963 (I1344908,I502431);
nor I_78964 (I1344925,I1344908,I502437);
nor I_78965 (I1344942,I1344925,I1344747);
DFFARX1 I_78966 (I1344942,I2507,I1344617,I1344606,);
not I_78967 (I1344973,I1344925);
DFFARX1 I_78968 (I1344973,I2507,I1344617,I1344999,);
not I_78969 (I1345007,I1344999);
nor I_78970 (I1344603,I1345007,I1344925);
nor I_78971 (I1345038,I1344908,I502419);
and I_78972 (I1345055,I1345038,I502434);
or I_78973 (I1345072,I1345055,I502422);
DFFARX1 I_78974 (I1345072,I2507,I1344617,I1345098,);
not I_78975 (I1345106,I1345098);
nand I_78976 (I1345123,I1345106,I1344846);
not I_78977 (I1344597,I1345123);
nand I_78978 (I1344591,I1345123,I1344863);
nand I_78979 (I1344588,I1345106,I1344730);
not I_78980 (I1345212,I2514);
DFFARX1 I_78981 (I1135825,I2507,I1345212,I1345238,);
DFFARX1 I_78982 (I1135837,I2507,I1345212,I1345255,);
not I_78983 (I1345263,I1345255);
nor I_78984 (I1345180,I1345238,I1345263);
DFFARX1 I_78985 (I1345263,I2507,I1345212,I1345195,);
nor I_78986 (I1345308,I1135834,I1135828);
and I_78987 (I1345325,I1345308,I1135822);
nor I_78988 (I1345342,I1345325,I1135834);
not I_78989 (I1345359,I1135834);
and I_78990 (I1345376,I1345359,I1135831);
nand I_78991 (I1345393,I1345376,I1135822);
nor I_78992 (I1345410,I1345359,I1345393);
DFFARX1 I_78993 (I1345410,I2507,I1345212,I1345177,);
not I_78994 (I1345441,I1345393);
nand I_78995 (I1345458,I1345263,I1345441);
nand I_78996 (I1345189,I1345325,I1345441);
DFFARX1 I_78997 (I1345359,I2507,I1345212,I1345204,);
not I_78998 (I1345503,I1135846);
nor I_78999 (I1345520,I1345503,I1135831);
nor I_79000 (I1345537,I1345520,I1345342);
DFFARX1 I_79001 (I1345537,I2507,I1345212,I1345201,);
not I_79002 (I1345568,I1345520);
DFFARX1 I_79003 (I1345568,I2507,I1345212,I1345594,);
not I_79004 (I1345602,I1345594);
nor I_79005 (I1345198,I1345602,I1345520);
nor I_79006 (I1345633,I1345503,I1135840);
and I_79007 (I1345650,I1345633,I1135843);
or I_79008 (I1345667,I1345650,I1135825);
DFFARX1 I_79009 (I1345667,I2507,I1345212,I1345693,);
not I_79010 (I1345701,I1345693);
nand I_79011 (I1345718,I1345701,I1345441);
not I_79012 (I1345192,I1345718);
nand I_79013 (I1345186,I1345718,I1345458);
nand I_79014 (I1345183,I1345701,I1345325);
not I_79015 (I1345807,I2514);
DFFARX1 I_79016 (I324518,I2507,I1345807,I1345833,);
DFFARX1 I_79017 (I324512,I2507,I1345807,I1345850,);
not I_79018 (I1345858,I1345850);
nor I_79019 (I1345775,I1345833,I1345858);
DFFARX1 I_79020 (I1345858,I2507,I1345807,I1345790,);
nor I_79021 (I1345903,I324500,I324521);
and I_79022 (I1345920,I1345903,I324515);
nor I_79023 (I1345937,I1345920,I324500);
not I_79024 (I1345954,I324500);
and I_79025 (I1345971,I1345954,I324497);
nand I_79026 (I1345988,I1345971,I324509);
nor I_79027 (I1346005,I1345954,I1345988);
DFFARX1 I_79028 (I1346005,I2507,I1345807,I1345772,);
not I_79029 (I1346036,I1345988);
nand I_79030 (I1346053,I1345858,I1346036);
nand I_79031 (I1345784,I1345920,I1346036);
DFFARX1 I_79032 (I1345954,I2507,I1345807,I1345799,);
not I_79033 (I1346098,I324524);
nor I_79034 (I1346115,I1346098,I324497);
nor I_79035 (I1346132,I1346115,I1345937);
DFFARX1 I_79036 (I1346132,I2507,I1345807,I1345796,);
not I_79037 (I1346163,I1346115);
DFFARX1 I_79038 (I1346163,I2507,I1345807,I1346189,);
not I_79039 (I1346197,I1346189);
nor I_79040 (I1345793,I1346197,I1346115);
nor I_79041 (I1346228,I1346098,I324506);
and I_79042 (I1346245,I1346228,I324503);
or I_79043 (I1346262,I1346245,I324497);
DFFARX1 I_79044 (I1346262,I2507,I1345807,I1346288,);
not I_79045 (I1346296,I1346288);
nand I_79046 (I1346313,I1346296,I1346036);
not I_79047 (I1345787,I1346313);
nand I_79048 (I1345781,I1346313,I1346053);
nand I_79049 (I1345778,I1346296,I1345920);
not I_79050 (I1346402,I2514);
DFFARX1 I_79051 (I895329,I2507,I1346402,I1346428,);
DFFARX1 I_79052 (I895347,I2507,I1346402,I1346445,);
not I_79053 (I1346453,I1346445);
nor I_79054 (I1346370,I1346428,I1346453);
DFFARX1 I_79055 (I1346453,I2507,I1346402,I1346385,);
nor I_79056 (I1346498,I895326,I895338);
and I_79057 (I1346515,I1346498,I895323);
nor I_79058 (I1346532,I1346515,I895326);
not I_79059 (I1346549,I895326);
and I_79060 (I1346566,I1346549,I895332);
nand I_79061 (I1346583,I1346566,I895344);
nor I_79062 (I1346600,I1346549,I1346583);
DFFARX1 I_79063 (I1346600,I2507,I1346402,I1346367,);
not I_79064 (I1346631,I1346583);
nand I_79065 (I1346648,I1346453,I1346631);
nand I_79066 (I1346379,I1346515,I1346631);
DFFARX1 I_79067 (I1346549,I2507,I1346402,I1346394,);
not I_79068 (I1346693,I895335);
nor I_79069 (I1346710,I1346693,I895332);
nor I_79070 (I1346727,I1346710,I1346532);
DFFARX1 I_79071 (I1346727,I2507,I1346402,I1346391,);
not I_79072 (I1346758,I1346710);
DFFARX1 I_79073 (I1346758,I2507,I1346402,I1346784,);
not I_79074 (I1346792,I1346784);
nor I_79075 (I1346388,I1346792,I1346710);
nor I_79076 (I1346823,I1346693,I895323);
and I_79077 (I1346840,I1346823,I895350);
or I_79078 (I1346857,I1346840,I895341);
DFFARX1 I_79079 (I1346857,I2507,I1346402,I1346883,);
not I_79080 (I1346891,I1346883);
nand I_79081 (I1346908,I1346891,I1346631);
not I_79082 (I1346382,I1346908);
nand I_79083 (I1346376,I1346908,I1346648);
nand I_79084 (I1346373,I1346891,I1346515);
not I_79085 (I1346997,I2514);
DFFARX1 I_79086 (I1053350,I2507,I1346997,I1347023,);
DFFARX1 I_79087 (I1053341,I2507,I1346997,I1347040,);
not I_79088 (I1347048,I1347040);
nor I_79089 (I1346965,I1347023,I1347048);
DFFARX1 I_79090 (I1347048,I2507,I1346997,I1346980,);
nor I_79091 (I1347093,I1053347,I1053356);
and I_79092 (I1347110,I1347093,I1053359);
nor I_79093 (I1347127,I1347110,I1053347);
not I_79094 (I1347144,I1053347);
and I_79095 (I1347161,I1347144,I1053338);
nand I_79096 (I1347178,I1347161,I1053344);
nor I_79097 (I1347195,I1347144,I1347178);
DFFARX1 I_79098 (I1347195,I2507,I1346997,I1346962,);
not I_79099 (I1347226,I1347178);
nand I_79100 (I1347243,I1347048,I1347226);
nand I_79101 (I1346974,I1347110,I1347226);
DFFARX1 I_79102 (I1347144,I2507,I1346997,I1346989,);
not I_79103 (I1347288,I1053353);
nor I_79104 (I1347305,I1347288,I1053338);
nor I_79105 (I1347322,I1347305,I1347127);
DFFARX1 I_79106 (I1347322,I2507,I1346997,I1346986,);
not I_79107 (I1347353,I1347305);
DFFARX1 I_79108 (I1347353,I2507,I1346997,I1347379,);
not I_79109 (I1347387,I1347379);
nor I_79110 (I1346983,I1347387,I1347305);
nor I_79111 (I1347418,I1347288,I1053338);
and I_79112 (I1347435,I1347418,I1053341);
or I_79113 (I1347452,I1347435,I1053344);
DFFARX1 I_79114 (I1347452,I2507,I1346997,I1347478,);
not I_79115 (I1347486,I1347478);
nand I_79116 (I1347503,I1347486,I1347226);
not I_79117 (I1346977,I1347503);
nand I_79118 (I1346971,I1347503,I1347243);
nand I_79119 (I1346968,I1347486,I1347110);
not I_79120 (I1347592,I2514);
DFFARX1 I_79121 (I1016885,I2507,I1347592,I1347618,);
DFFARX1 I_79122 (I1016876,I2507,I1347592,I1347635,);
not I_79123 (I1347643,I1347635);
nor I_79124 (I1347560,I1347618,I1347643);
DFFARX1 I_79125 (I1347643,I2507,I1347592,I1347575,);
nor I_79126 (I1347688,I1016882,I1016891);
and I_79127 (I1347705,I1347688,I1016894);
nor I_79128 (I1347722,I1347705,I1016882);
not I_79129 (I1347739,I1016882);
and I_79130 (I1347756,I1347739,I1016873);
nand I_79131 (I1347773,I1347756,I1016879);
nor I_79132 (I1347790,I1347739,I1347773);
DFFARX1 I_79133 (I1347790,I2507,I1347592,I1347557,);
not I_79134 (I1347821,I1347773);
nand I_79135 (I1347838,I1347643,I1347821);
nand I_79136 (I1347569,I1347705,I1347821);
DFFARX1 I_79137 (I1347739,I2507,I1347592,I1347584,);
not I_79138 (I1347883,I1016888);
nor I_79139 (I1347900,I1347883,I1016873);
nor I_79140 (I1347917,I1347900,I1347722);
DFFARX1 I_79141 (I1347917,I2507,I1347592,I1347581,);
not I_79142 (I1347948,I1347900);
DFFARX1 I_79143 (I1347948,I2507,I1347592,I1347974,);
not I_79144 (I1347982,I1347974);
nor I_79145 (I1347578,I1347982,I1347900);
nor I_79146 (I1348013,I1347883,I1016873);
and I_79147 (I1348030,I1348013,I1016876);
or I_79148 (I1348047,I1348030,I1016879);
DFFARX1 I_79149 (I1348047,I2507,I1347592,I1348073,);
not I_79150 (I1348081,I1348073);
nand I_79151 (I1348098,I1348081,I1347821);
not I_79152 (I1347572,I1348098);
nand I_79153 (I1347566,I1348098,I1347838);
nand I_79154 (I1347563,I1348081,I1347705);
not I_79155 (I1348187,I2514);
DFFARX1 I_79156 (I154395,I2507,I1348187,I1348213,);
DFFARX1 I_79157 (I154398,I2507,I1348187,I1348230,);
not I_79158 (I1348238,I1348230);
nor I_79159 (I1348155,I1348213,I1348238);
DFFARX1 I_79160 (I1348238,I2507,I1348187,I1348170,);
nor I_79161 (I1348283,I154404,I154398);
and I_79162 (I1348300,I1348283,I154401);
nor I_79163 (I1348317,I1348300,I154404);
not I_79164 (I1348334,I154404);
and I_79165 (I1348351,I1348334,I154395);
nand I_79166 (I1348368,I1348351,I154413);
nor I_79167 (I1348385,I1348334,I1348368);
DFFARX1 I_79168 (I1348385,I2507,I1348187,I1348152,);
not I_79169 (I1348416,I1348368);
nand I_79170 (I1348433,I1348238,I1348416);
nand I_79171 (I1348164,I1348300,I1348416);
DFFARX1 I_79172 (I1348334,I2507,I1348187,I1348179,);
not I_79173 (I1348478,I154407);
nor I_79174 (I1348495,I1348478,I154395);
nor I_79175 (I1348512,I1348495,I1348317);
DFFARX1 I_79176 (I1348512,I2507,I1348187,I1348176,);
not I_79177 (I1348543,I1348495);
DFFARX1 I_79178 (I1348543,I2507,I1348187,I1348569,);
not I_79179 (I1348577,I1348569);
nor I_79180 (I1348173,I1348577,I1348495);
nor I_79181 (I1348608,I1348478,I154410);
and I_79182 (I1348625,I1348608,I154416);
or I_79183 (I1348642,I1348625,I154419);
DFFARX1 I_79184 (I1348642,I2507,I1348187,I1348668,);
not I_79185 (I1348676,I1348668);
nand I_79186 (I1348693,I1348676,I1348416);
not I_79187 (I1348167,I1348693);
nand I_79188 (I1348161,I1348693,I1348433);
nand I_79189 (I1348158,I1348676,I1348300);
not I_79190 (I1348782,I2514);
DFFARX1 I_79191 (I56989,I2507,I1348782,I1348808,);
DFFARX1 I_79192 (I56977,I2507,I1348782,I1348825,);
not I_79193 (I1348833,I1348825);
nor I_79194 (I1348750,I1348808,I1348833);
DFFARX1 I_79195 (I1348833,I2507,I1348782,I1348765,);
nor I_79196 (I1348878,I56968,I56992);
and I_79197 (I1348895,I1348878,I56971);
nor I_79198 (I1348912,I1348895,I56968);
not I_79199 (I1348929,I56968);
and I_79200 (I1348946,I1348929,I56974);
nand I_79201 (I1348963,I1348946,I56986);
nor I_79202 (I1348980,I1348929,I1348963);
DFFARX1 I_79203 (I1348980,I2507,I1348782,I1348747,);
not I_79204 (I1349011,I1348963);
nand I_79205 (I1349028,I1348833,I1349011);
nand I_79206 (I1348759,I1348895,I1349011);
DFFARX1 I_79207 (I1348929,I2507,I1348782,I1348774,);
not I_79208 (I1349073,I56968);
nor I_79209 (I1349090,I1349073,I56974);
nor I_79210 (I1349107,I1349090,I1348912);
DFFARX1 I_79211 (I1349107,I2507,I1348782,I1348771,);
not I_79212 (I1349138,I1349090);
DFFARX1 I_79213 (I1349138,I2507,I1348782,I1349164,);
not I_79214 (I1349172,I1349164);
nor I_79215 (I1348768,I1349172,I1349090);
nor I_79216 (I1349203,I1349073,I56971);
and I_79217 (I1349220,I1349203,I56980);
or I_79218 (I1349237,I1349220,I56983);
DFFARX1 I_79219 (I1349237,I2507,I1348782,I1349263,);
not I_79220 (I1349271,I1349263);
nand I_79221 (I1349288,I1349271,I1349011);
not I_79222 (I1348762,I1349288);
nand I_79223 (I1348756,I1349288,I1349028);
nand I_79224 (I1348753,I1349271,I1348895);
not I_79225 (I1349377,I2514);
DFFARX1 I_79226 (I830715,I2507,I1349377,I1349403,);
DFFARX1 I_79227 (I830712,I2507,I1349377,I1349420,);
not I_79228 (I1349428,I1349420);
nor I_79229 (I1349345,I1349403,I1349428);
DFFARX1 I_79230 (I1349428,I2507,I1349377,I1349360,);
nor I_79231 (I1349473,I830727,I830709);
and I_79232 (I1349490,I1349473,I830706);
nor I_79233 (I1349507,I1349490,I830727);
not I_79234 (I1349524,I830727);
and I_79235 (I1349541,I1349524,I830712);
nand I_79236 (I1349558,I1349541,I830724);
nor I_79237 (I1349575,I1349524,I1349558);
DFFARX1 I_79238 (I1349575,I2507,I1349377,I1349342,);
not I_79239 (I1349606,I1349558);
nand I_79240 (I1349623,I1349428,I1349606);
nand I_79241 (I1349354,I1349490,I1349606);
DFFARX1 I_79242 (I1349524,I2507,I1349377,I1349369,);
not I_79243 (I1349668,I830718);
nor I_79244 (I1349685,I1349668,I830712);
nor I_79245 (I1349702,I1349685,I1349507);
DFFARX1 I_79246 (I1349702,I2507,I1349377,I1349366,);
not I_79247 (I1349733,I1349685);
DFFARX1 I_79248 (I1349733,I2507,I1349377,I1349759,);
not I_79249 (I1349767,I1349759);
nor I_79250 (I1349363,I1349767,I1349685);
nor I_79251 (I1349798,I1349668,I830706);
and I_79252 (I1349815,I1349798,I830721);
or I_79253 (I1349832,I1349815,I830709);
DFFARX1 I_79254 (I1349832,I2507,I1349377,I1349858,);
not I_79255 (I1349866,I1349858);
nand I_79256 (I1349883,I1349866,I1349606);
not I_79257 (I1349357,I1349883);
nand I_79258 (I1349351,I1349883,I1349623);
nand I_79259 (I1349348,I1349866,I1349490);
not I_79260 (I1349972,I2514);
DFFARX1 I_79261 (I1144495,I2507,I1349972,I1349998,);
DFFARX1 I_79262 (I1144507,I2507,I1349972,I1350015,);
not I_79263 (I1350023,I1350015);
nor I_79264 (I1349940,I1349998,I1350023);
DFFARX1 I_79265 (I1350023,I2507,I1349972,I1349955,);
nor I_79266 (I1350068,I1144504,I1144498);
and I_79267 (I1350085,I1350068,I1144492);
nor I_79268 (I1350102,I1350085,I1144504);
not I_79269 (I1350119,I1144504);
and I_79270 (I1350136,I1350119,I1144501);
nand I_79271 (I1350153,I1350136,I1144492);
nor I_79272 (I1350170,I1350119,I1350153);
DFFARX1 I_79273 (I1350170,I2507,I1349972,I1349937,);
not I_79274 (I1350201,I1350153);
nand I_79275 (I1350218,I1350023,I1350201);
nand I_79276 (I1349949,I1350085,I1350201);
DFFARX1 I_79277 (I1350119,I2507,I1349972,I1349964,);
not I_79278 (I1350263,I1144516);
nor I_79279 (I1350280,I1350263,I1144501);
nor I_79280 (I1350297,I1350280,I1350102);
DFFARX1 I_79281 (I1350297,I2507,I1349972,I1349961,);
not I_79282 (I1350328,I1350280);
DFFARX1 I_79283 (I1350328,I2507,I1349972,I1350354,);
not I_79284 (I1350362,I1350354);
nor I_79285 (I1349958,I1350362,I1350280);
nor I_79286 (I1350393,I1350263,I1144510);
and I_79287 (I1350410,I1350393,I1144513);
or I_79288 (I1350427,I1350410,I1144495);
DFFARX1 I_79289 (I1350427,I2507,I1349972,I1350453,);
not I_79290 (I1350461,I1350453);
nand I_79291 (I1350478,I1350461,I1350201);
not I_79292 (I1349952,I1350478);
nand I_79293 (I1349946,I1350478,I1350218);
nand I_79294 (I1349943,I1350461,I1350085);
not I_79295 (I1350567,I2514);
DFFARX1 I_79296 (I369313,I2507,I1350567,I1350593,);
DFFARX1 I_79297 (I369307,I2507,I1350567,I1350610,);
not I_79298 (I1350618,I1350610);
nor I_79299 (I1350535,I1350593,I1350618);
DFFARX1 I_79300 (I1350618,I2507,I1350567,I1350550,);
nor I_79301 (I1350663,I369295,I369316);
and I_79302 (I1350680,I1350663,I369310);
nor I_79303 (I1350697,I1350680,I369295);
not I_79304 (I1350714,I369295);
and I_79305 (I1350731,I1350714,I369292);
nand I_79306 (I1350748,I1350731,I369304);
nor I_79307 (I1350765,I1350714,I1350748);
DFFARX1 I_79308 (I1350765,I2507,I1350567,I1350532,);
not I_79309 (I1350796,I1350748);
nand I_79310 (I1350813,I1350618,I1350796);
nand I_79311 (I1350544,I1350680,I1350796);
DFFARX1 I_79312 (I1350714,I2507,I1350567,I1350559,);
not I_79313 (I1350858,I369319);
nor I_79314 (I1350875,I1350858,I369292);
nor I_79315 (I1350892,I1350875,I1350697);
DFFARX1 I_79316 (I1350892,I2507,I1350567,I1350556,);
not I_79317 (I1350923,I1350875);
DFFARX1 I_79318 (I1350923,I2507,I1350567,I1350949,);
not I_79319 (I1350957,I1350949);
nor I_79320 (I1350553,I1350957,I1350875);
nor I_79321 (I1350988,I1350858,I369301);
and I_79322 (I1351005,I1350988,I369298);
or I_79323 (I1351022,I1351005,I369292);
DFFARX1 I_79324 (I1351022,I2507,I1350567,I1351048,);
not I_79325 (I1351056,I1351048);
nand I_79326 (I1351073,I1351056,I1350796);
not I_79327 (I1350547,I1351073);
nand I_79328 (I1350541,I1351073,I1350813);
nand I_79329 (I1350538,I1351056,I1350680);
not I_79330 (I1351162,I2514);
DFFARX1 I_79331 (I1044374,I2507,I1351162,I1351188,);
DFFARX1 I_79332 (I1044365,I2507,I1351162,I1351205,);
not I_79333 (I1351213,I1351205);
nor I_79334 (I1351130,I1351188,I1351213);
DFFARX1 I_79335 (I1351213,I2507,I1351162,I1351145,);
nor I_79336 (I1351258,I1044371,I1044380);
and I_79337 (I1351275,I1351258,I1044383);
nor I_79338 (I1351292,I1351275,I1044371);
not I_79339 (I1351309,I1044371);
and I_79340 (I1351326,I1351309,I1044362);
nand I_79341 (I1351343,I1351326,I1044368);
nor I_79342 (I1351360,I1351309,I1351343);
DFFARX1 I_79343 (I1351360,I2507,I1351162,I1351127,);
not I_79344 (I1351391,I1351343);
nand I_79345 (I1351408,I1351213,I1351391);
nand I_79346 (I1351139,I1351275,I1351391);
DFFARX1 I_79347 (I1351309,I2507,I1351162,I1351154,);
not I_79348 (I1351453,I1044377);
nor I_79349 (I1351470,I1351453,I1044362);
nor I_79350 (I1351487,I1351470,I1351292);
DFFARX1 I_79351 (I1351487,I2507,I1351162,I1351151,);
not I_79352 (I1351518,I1351470);
DFFARX1 I_79353 (I1351518,I2507,I1351162,I1351544,);
not I_79354 (I1351552,I1351544);
nor I_79355 (I1351148,I1351552,I1351470);
nor I_79356 (I1351583,I1351453,I1044362);
and I_79357 (I1351600,I1351583,I1044365);
or I_79358 (I1351617,I1351600,I1044368);
DFFARX1 I_79359 (I1351617,I2507,I1351162,I1351643,);
not I_79360 (I1351651,I1351643);
nand I_79361 (I1351668,I1351651,I1351391);
not I_79362 (I1351142,I1351668);
nand I_79363 (I1351136,I1351668,I1351408);
nand I_79364 (I1351133,I1351651,I1351275);
not I_79365 (I1351757,I2514);
DFFARX1 I_79366 (I92825,I2507,I1351757,I1351783,);
DFFARX1 I_79367 (I92813,I2507,I1351757,I1351800,);
not I_79368 (I1351808,I1351800);
nor I_79369 (I1351725,I1351783,I1351808);
DFFARX1 I_79370 (I1351808,I2507,I1351757,I1351740,);
nor I_79371 (I1351853,I92804,I92828);
and I_79372 (I1351870,I1351853,I92807);
nor I_79373 (I1351887,I1351870,I92804);
not I_79374 (I1351904,I92804);
and I_79375 (I1351921,I1351904,I92810);
nand I_79376 (I1351938,I1351921,I92822);
nor I_79377 (I1351955,I1351904,I1351938);
DFFARX1 I_79378 (I1351955,I2507,I1351757,I1351722,);
not I_79379 (I1351986,I1351938);
nand I_79380 (I1352003,I1351808,I1351986);
nand I_79381 (I1351734,I1351870,I1351986);
DFFARX1 I_79382 (I1351904,I2507,I1351757,I1351749,);
not I_79383 (I1352048,I92804);
nor I_79384 (I1352065,I1352048,I92810);
nor I_79385 (I1352082,I1352065,I1351887);
DFFARX1 I_79386 (I1352082,I2507,I1351757,I1351746,);
not I_79387 (I1352113,I1352065);
DFFARX1 I_79388 (I1352113,I2507,I1351757,I1352139,);
not I_79389 (I1352147,I1352139);
nor I_79390 (I1351743,I1352147,I1352065);
nor I_79391 (I1352178,I1352048,I92807);
and I_79392 (I1352195,I1352178,I92816);
or I_79393 (I1352212,I1352195,I92819);
DFFARX1 I_79394 (I1352212,I2507,I1351757,I1352238,);
not I_79395 (I1352246,I1352238);
nand I_79396 (I1352263,I1352246,I1351986);
not I_79397 (I1351737,I1352263);
nand I_79398 (I1351731,I1352263,I1352003);
nand I_79399 (I1351728,I1352246,I1351870);
not I_79400 (I1352352,I2514);
DFFARX1 I_79401 (I988999,I2507,I1352352,I1352378,);
DFFARX1 I_79402 (I989017,I2507,I1352352,I1352395,);
not I_79403 (I1352403,I1352395);
nor I_79404 (I1352320,I1352378,I1352403);
DFFARX1 I_79405 (I1352403,I2507,I1352352,I1352335,);
nor I_79406 (I1352448,I988996,I989008);
and I_79407 (I1352465,I1352448,I988993);
nor I_79408 (I1352482,I1352465,I988996);
not I_79409 (I1352499,I988996);
and I_79410 (I1352516,I1352499,I989002);
nand I_79411 (I1352533,I1352516,I989014);
nor I_79412 (I1352550,I1352499,I1352533);
DFFARX1 I_79413 (I1352550,I2507,I1352352,I1352317,);
not I_79414 (I1352581,I1352533);
nand I_79415 (I1352598,I1352403,I1352581);
nand I_79416 (I1352329,I1352465,I1352581);
DFFARX1 I_79417 (I1352499,I2507,I1352352,I1352344,);
not I_79418 (I1352643,I989005);
nor I_79419 (I1352660,I1352643,I989002);
nor I_79420 (I1352677,I1352660,I1352482);
DFFARX1 I_79421 (I1352677,I2507,I1352352,I1352341,);
not I_79422 (I1352708,I1352660);
DFFARX1 I_79423 (I1352708,I2507,I1352352,I1352734,);
not I_79424 (I1352742,I1352734);
nor I_79425 (I1352338,I1352742,I1352660);
nor I_79426 (I1352773,I1352643,I988993);
and I_79427 (I1352790,I1352773,I989020);
or I_79428 (I1352807,I1352790,I989011);
DFFARX1 I_79429 (I1352807,I2507,I1352352,I1352833,);
not I_79430 (I1352841,I1352833);
nand I_79431 (I1352858,I1352841,I1352581);
not I_79432 (I1352332,I1352858);
nand I_79433 (I1352326,I1352858,I1352598);
nand I_79434 (I1352323,I1352841,I1352465);
not I_79435 (I1352947,I2514);
DFFARX1 I_79436 (I216870,I2507,I1352947,I1352973,);
DFFARX1 I_79437 (I216873,I2507,I1352947,I1352990,);
not I_79438 (I1352998,I1352990);
nor I_79439 (I1352915,I1352973,I1352998);
DFFARX1 I_79440 (I1352998,I2507,I1352947,I1352930,);
nor I_79441 (I1353043,I216879,I216873);
and I_79442 (I1353060,I1353043,I216876);
nor I_79443 (I1353077,I1353060,I216879);
not I_79444 (I1353094,I216879);
and I_79445 (I1353111,I1353094,I216870);
nand I_79446 (I1353128,I1353111,I216888);
nor I_79447 (I1353145,I1353094,I1353128);
DFFARX1 I_79448 (I1353145,I2507,I1352947,I1352912,);
not I_79449 (I1353176,I1353128);
nand I_79450 (I1353193,I1352998,I1353176);
nand I_79451 (I1352924,I1353060,I1353176);
DFFARX1 I_79452 (I1353094,I2507,I1352947,I1352939,);
not I_79453 (I1353238,I216882);
nor I_79454 (I1353255,I1353238,I216870);
nor I_79455 (I1353272,I1353255,I1353077);
DFFARX1 I_79456 (I1353272,I2507,I1352947,I1352936,);
not I_79457 (I1353303,I1353255);
DFFARX1 I_79458 (I1353303,I2507,I1352947,I1353329,);
not I_79459 (I1353337,I1353329);
nor I_79460 (I1352933,I1353337,I1353255);
nor I_79461 (I1353368,I1353238,I216885);
and I_79462 (I1353385,I1353368,I216891);
or I_79463 (I1353402,I1353385,I216894);
DFFARX1 I_79464 (I1353402,I2507,I1352947,I1353428,);
not I_79465 (I1353436,I1353428);
nand I_79466 (I1353453,I1353436,I1353176);
not I_79467 (I1352927,I1353453);
nand I_79468 (I1352921,I1353453,I1353193);
nand I_79469 (I1352918,I1353436,I1353060);
not I_79470 (I1353542,I2514);
DFFARX1 I_79471 (I788555,I2507,I1353542,I1353568,);
DFFARX1 I_79472 (I788552,I2507,I1353542,I1353585,);
not I_79473 (I1353593,I1353585);
nor I_79474 (I1353510,I1353568,I1353593);
DFFARX1 I_79475 (I1353593,I2507,I1353542,I1353525,);
nor I_79476 (I1353638,I788567,I788549);
and I_79477 (I1353655,I1353638,I788546);
nor I_79478 (I1353672,I1353655,I788567);
not I_79479 (I1353689,I788567);
and I_79480 (I1353706,I1353689,I788552);
nand I_79481 (I1353723,I1353706,I788564);
nor I_79482 (I1353740,I1353689,I1353723);
DFFARX1 I_79483 (I1353740,I2507,I1353542,I1353507,);
not I_79484 (I1353771,I1353723);
nand I_79485 (I1353788,I1353593,I1353771);
nand I_79486 (I1353519,I1353655,I1353771);
DFFARX1 I_79487 (I1353689,I2507,I1353542,I1353534,);
not I_79488 (I1353833,I788558);
nor I_79489 (I1353850,I1353833,I788552);
nor I_79490 (I1353867,I1353850,I1353672);
DFFARX1 I_79491 (I1353867,I2507,I1353542,I1353531,);
not I_79492 (I1353898,I1353850);
DFFARX1 I_79493 (I1353898,I2507,I1353542,I1353924,);
not I_79494 (I1353932,I1353924);
nor I_79495 (I1353528,I1353932,I1353850);
nor I_79496 (I1353963,I1353833,I788546);
and I_79497 (I1353980,I1353963,I788561);
or I_79498 (I1353997,I1353980,I788549);
DFFARX1 I_79499 (I1353997,I2507,I1353542,I1354023,);
not I_79500 (I1354031,I1354023);
nand I_79501 (I1354048,I1354031,I1353771);
not I_79502 (I1353522,I1354048);
nand I_79503 (I1353516,I1354048,I1353788);
nand I_79504 (I1353513,I1354031,I1353655);
not I_79505 (I1354137,I2514);
DFFARX1 I_79506 (I639987,I2507,I1354137,I1354163,);
DFFARX1 I_79507 (I639969,I2507,I1354137,I1354180,);
not I_79508 (I1354188,I1354180);
nor I_79509 (I1354105,I1354163,I1354188);
DFFARX1 I_79510 (I1354188,I2507,I1354137,I1354120,);
nor I_79511 (I1354233,I639975,I639978);
and I_79512 (I1354250,I1354233,I639966);
nor I_79513 (I1354267,I1354250,I639975);
not I_79514 (I1354284,I639975);
and I_79515 (I1354301,I1354284,I639984);
nand I_79516 (I1354318,I1354301,I639972);
nor I_79517 (I1354335,I1354284,I1354318);
DFFARX1 I_79518 (I1354335,I2507,I1354137,I1354102,);
not I_79519 (I1354366,I1354318);
nand I_79520 (I1354383,I1354188,I1354366);
nand I_79521 (I1354114,I1354250,I1354366);
DFFARX1 I_79522 (I1354284,I2507,I1354137,I1354129,);
not I_79523 (I1354428,I639969);
nor I_79524 (I1354445,I1354428,I639984);
nor I_79525 (I1354462,I1354445,I1354267);
DFFARX1 I_79526 (I1354462,I2507,I1354137,I1354126,);
not I_79527 (I1354493,I1354445);
DFFARX1 I_79528 (I1354493,I2507,I1354137,I1354519,);
not I_79529 (I1354527,I1354519);
nor I_79530 (I1354123,I1354527,I1354445);
nor I_79531 (I1354558,I1354428,I639981);
and I_79532 (I1354575,I1354558,I639990);
or I_79533 (I1354592,I1354575,I639966);
DFFARX1 I_79534 (I1354592,I2507,I1354137,I1354618,);
not I_79535 (I1354626,I1354618);
nand I_79536 (I1354643,I1354626,I1354366);
not I_79537 (I1354117,I1354643);
nand I_79538 (I1354111,I1354643,I1354383);
nand I_79539 (I1354108,I1354626,I1354250);
not I_79540 (I1354732,I2514);
DFFARX1 I_79541 (I692585,I2507,I1354732,I1354758,);
DFFARX1 I_79542 (I692567,I2507,I1354732,I1354775,);
not I_79543 (I1354783,I1354775);
nor I_79544 (I1354700,I1354758,I1354783);
DFFARX1 I_79545 (I1354783,I2507,I1354732,I1354715,);
nor I_79546 (I1354828,I692573,I692576);
and I_79547 (I1354845,I1354828,I692564);
nor I_79548 (I1354862,I1354845,I692573);
not I_79549 (I1354879,I692573);
and I_79550 (I1354896,I1354879,I692582);
nand I_79551 (I1354913,I1354896,I692570);
nor I_79552 (I1354930,I1354879,I1354913);
DFFARX1 I_79553 (I1354930,I2507,I1354732,I1354697,);
not I_79554 (I1354961,I1354913);
nand I_79555 (I1354978,I1354783,I1354961);
nand I_79556 (I1354709,I1354845,I1354961);
DFFARX1 I_79557 (I1354879,I2507,I1354732,I1354724,);
not I_79558 (I1355023,I692567);
nor I_79559 (I1355040,I1355023,I692582);
nor I_79560 (I1355057,I1355040,I1354862);
DFFARX1 I_79561 (I1355057,I2507,I1354732,I1354721,);
not I_79562 (I1355088,I1355040);
DFFARX1 I_79563 (I1355088,I2507,I1354732,I1355114,);
not I_79564 (I1355122,I1355114);
nor I_79565 (I1354718,I1355122,I1355040);
nor I_79566 (I1355153,I1355023,I692579);
and I_79567 (I1355170,I1355153,I692588);
or I_79568 (I1355187,I1355170,I692564);
DFFARX1 I_79569 (I1355187,I2507,I1354732,I1355213,);
not I_79570 (I1355221,I1355213);
nand I_79571 (I1355238,I1355221,I1354961);
not I_79572 (I1354712,I1355238);
nand I_79573 (I1354706,I1355238,I1354978);
nand I_79574 (I1354703,I1355221,I1354845);
not I_79575 (I1355327,I2514);
DFFARX1 I_79576 (I577563,I2507,I1355327,I1355353,);
DFFARX1 I_79577 (I577557,I2507,I1355327,I1355370,);
not I_79578 (I1355378,I1355370);
nor I_79579 (I1355295,I1355353,I1355378);
DFFARX1 I_79580 (I1355378,I2507,I1355327,I1355310,);
nor I_79581 (I1355423,I577554,I577545);
and I_79582 (I1355440,I1355423,I577542);
nor I_79583 (I1355457,I1355440,I577554);
not I_79584 (I1355474,I577554);
and I_79585 (I1355491,I1355474,I577548);
nand I_79586 (I1355508,I1355491,I577560);
nor I_79587 (I1355525,I1355474,I1355508);
DFFARX1 I_79588 (I1355525,I2507,I1355327,I1355292,);
not I_79589 (I1355556,I1355508);
nand I_79590 (I1355573,I1355378,I1355556);
nand I_79591 (I1355304,I1355440,I1355556);
DFFARX1 I_79592 (I1355474,I2507,I1355327,I1355319,);
not I_79593 (I1355618,I577566);
nor I_79594 (I1355635,I1355618,I577548);
nor I_79595 (I1355652,I1355635,I1355457);
DFFARX1 I_79596 (I1355652,I2507,I1355327,I1355316,);
not I_79597 (I1355683,I1355635);
DFFARX1 I_79598 (I1355683,I2507,I1355327,I1355709,);
not I_79599 (I1355717,I1355709);
nor I_79600 (I1355313,I1355717,I1355635);
nor I_79601 (I1355748,I1355618,I577545);
and I_79602 (I1355765,I1355748,I577551);
or I_79603 (I1355782,I1355765,I577542);
DFFARX1 I_79604 (I1355782,I2507,I1355327,I1355808,);
not I_79605 (I1355816,I1355808);
nand I_79606 (I1355833,I1355816,I1355556);
not I_79607 (I1355307,I1355833);
nand I_79608 (I1355301,I1355833,I1355573);
nand I_79609 (I1355298,I1355816,I1355440);
not I_79610 (I1355922,I2514);
DFFARX1 I_79611 (I454479,I2507,I1355922,I1355948,);
DFFARX1 I_79612 (I454485,I2507,I1355922,I1355965,);
not I_79613 (I1355973,I1355965);
nor I_79614 (I1355890,I1355948,I1355973);
DFFARX1 I_79615 (I1355973,I2507,I1355922,I1355905,);
nor I_79616 (I1356018,I454494,I454479);
and I_79617 (I1356035,I1356018,I454506);
nor I_79618 (I1356052,I1356035,I454494);
not I_79619 (I1356069,I454494);
and I_79620 (I1356086,I1356069,I454482);
nand I_79621 (I1356103,I1356086,I454503);
nor I_79622 (I1356120,I1356069,I1356103);
DFFARX1 I_79623 (I1356120,I2507,I1355922,I1355887,);
not I_79624 (I1356151,I1356103);
nand I_79625 (I1356168,I1355973,I1356151);
nand I_79626 (I1355899,I1356035,I1356151);
DFFARX1 I_79627 (I1356069,I2507,I1355922,I1355914,);
not I_79628 (I1356213,I454491);
nor I_79629 (I1356230,I1356213,I454482);
nor I_79630 (I1356247,I1356230,I1356052);
DFFARX1 I_79631 (I1356247,I2507,I1355922,I1355911,);
not I_79632 (I1356278,I1356230);
DFFARX1 I_79633 (I1356278,I2507,I1355922,I1356304,);
not I_79634 (I1356312,I1356304);
nor I_79635 (I1355908,I1356312,I1356230);
nor I_79636 (I1356343,I1356213,I454488);
and I_79637 (I1356360,I1356343,I454500);
or I_79638 (I1356377,I1356360,I454497);
DFFARX1 I_79639 (I1356377,I2507,I1355922,I1356403,);
not I_79640 (I1356411,I1356403);
nand I_79641 (I1356428,I1356411,I1356151);
not I_79642 (I1355902,I1356428);
nand I_79643 (I1355896,I1356428,I1356168);
nand I_79644 (I1355893,I1356411,I1356035);
not I_79645 (I1356517,I2514);
DFFARX1 I_79646 (I928275,I2507,I1356517,I1356543,);
DFFARX1 I_79647 (I928293,I2507,I1356517,I1356560,);
not I_79648 (I1356568,I1356560);
nor I_79649 (I1356485,I1356543,I1356568);
DFFARX1 I_79650 (I1356568,I2507,I1356517,I1356500,);
nor I_79651 (I1356613,I928272,I928284);
and I_79652 (I1356630,I1356613,I928269);
nor I_79653 (I1356647,I1356630,I928272);
not I_79654 (I1356664,I928272);
and I_79655 (I1356681,I1356664,I928278);
nand I_79656 (I1356698,I1356681,I928290);
nor I_79657 (I1356715,I1356664,I1356698);
DFFARX1 I_79658 (I1356715,I2507,I1356517,I1356482,);
not I_79659 (I1356746,I1356698);
nand I_79660 (I1356763,I1356568,I1356746);
nand I_79661 (I1356494,I1356630,I1356746);
DFFARX1 I_79662 (I1356664,I2507,I1356517,I1356509,);
not I_79663 (I1356808,I928281);
nor I_79664 (I1356825,I1356808,I928278);
nor I_79665 (I1356842,I1356825,I1356647);
DFFARX1 I_79666 (I1356842,I2507,I1356517,I1356506,);
not I_79667 (I1356873,I1356825);
DFFARX1 I_79668 (I1356873,I2507,I1356517,I1356899,);
not I_79669 (I1356907,I1356899);
nor I_79670 (I1356503,I1356907,I1356825);
nor I_79671 (I1356938,I1356808,I928269);
and I_79672 (I1356955,I1356938,I928296);
or I_79673 (I1356972,I1356955,I928287);
DFFARX1 I_79674 (I1356972,I2507,I1356517,I1356998,);
not I_79675 (I1357006,I1356998);
nand I_79676 (I1357023,I1357006,I1356746);
not I_79677 (I1356497,I1357023);
nand I_79678 (I1356491,I1357023,I1356763);
nand I_79679 (I1356488,I1357006,I1356630);
not I_79680 (I1357112,I2514);
DFFARX1 I_79681 (I433263,I2507,I1357112,I1357138,);
DFFARX1 I_79682 (I433269,I2507,I1357112,I1357155,);
not I_79683 (I1357163,I1357155);
nor I_79684 (I1357080,I1357138,I1357163);
DFFARX1 I_79685 (I1357163,I2507,I1357112,I1357095,);
nor I_79686 (I1357208,I433278,I433263);
and I_79687 (I1357225,I1357208,I433290);
nor I_79688 (I1357242,I1357225,I433278);
not I_79689 (I1357259,I433278);
and I_79690 (I1357276,I1357259,I433266);
nand I_79691 (I1357293,I1357276,I433287);
nor I_79692 (I1357310,I1357259,I1357293);
DFFARX1 I_79693 (I1357310,I2507,I1357112,I1357077,);
not I_79694 (I1357341,I1357293);
nand I_79695 (I1357358,I1357163,I1357341);
nand I_79696 (I1357089,I1357225,I1357341);
DFFARX1 I_79697 (I1357259,I2507,I1357112,I1357104,);
not I_79698 (I1357403,I433275);
nor I_79699 (I1357420,I1357403,I433266);
nor I_79700 (I1357437,I1357420,I1357242);
DFFARX1 I_79701 (I1357437,I2507,I1357112,I1357101,);
not I_79702 (I1357468,I1357420);
DFFARX1 I_79703 (I1357468,I2507,I1357112,I1357494,);
not I_79704 (I1357502,I1357494);
nor I_79705 (I1357098,I1357502,I1357420);
nor I_79706 (I1357533,I1357403,I433272);
and I_79707 (I1357550,I1357533,I433284);
or I_79708 (I1357567,I1357550,I433281);
DFFARX1 I_79709 (I1357567,I2507,I1357112,I1357593,);
not I_79710 (I1357601,I1357593);
nand I_79711 (I1357618,I1357601,I1357341);
not I_79712 (I1357092,I1357618);
nand I_79713 (I1357086,I1357618,I1357358);
nand I_79714 (I1357083,I1357601,I1357225);
not I_79715 (I1357707,I2514);
DFFARX1 I_79716 (I930213,I2507,I1357707,I1357733,);
DFFARX1 I_79717 (I930231,I2507,I1357707,I1357750,);
not I_79718 (I1357758,I1357750);
nor I_79719 (I1357675,I1357733,I1357758);
DFFARX1 I_79720 (I1357758,I2507,I1357707,I1357690,);
nor I_79721 (I1357803,I930210,I930222);
and I_79722 (I1357820,I1357803,I930207);
nor I_79723 (I1357837,I1357820,I930210);
not I_79724 (I1357854,I930210);
and I_79725 (I1357871,I1357854,I930216);
nand I_79726 (I1357888,I1357871,I930228);
nor I_79727 (I1357905,I1357854,I1357888);
DFFARX1 I_79728 (I1357905,I2507,I1357707,I1357672,);
not I_79729 (I1357936,I1357888);
nand I_79730 (I1357953,I1357758,I1357936);
nand I_79731 (I1357684,I1357820,I1357936);
DFFARX1 I_79732 (I1357854,I2507,I1357707,I1357699,);
not I_79733 (I1357998,I930219);
nor I_79734 (I1358015,I1357998,I930216);
nor I_79735 (I1358032,I1358015,I1357837);
DFFARX1 I_79736 (I1358032,I2507,I1357707,I1357696,);
not I_79737 (I1358063,I1358015);
DFFARX1 I_79738 (I1358063,I2507,I1357707,I1358089,);
not I_79739 (I1358097,I1358089);
nor I_79740 (I1357693,I1358097,I1358015);
nor I_79741 (I1358128,I1357998,I930207);
and I_79742 (I1358145,I1358128,I930234);
or I_79743 (I1358162,I1358145,I930225);
DFFARX1 I_79744 (I1358162,I2507,I1357707,I1358188,);
not I_79745 (I1358196,I1358188);
nand I_79746 (I1358213,I1358196,I1357936);
not I_79747 (I1357687,I1358213);
nand I_79748 (I1357681,I1358213,I1357953);
nand I_79749 (I1357678,I1358196,I1357820);
not I_79750 (I1358302,I2514);
DFFARX1 I_79751 (I364043,I2507,I1358302,I1358328,);
DFFARX1 I_79752 (I364037,I2507,I1358302,I1358345,);
not I_79753 (I1358353,I1358345);
nor I_79754 (I1358270,I1358328,I1358353);
DFFARX1 I_79755 (I1358353,I2507,I1358302,I1358285,);
nor I_79756 (I1358398,I364025,I364046);
and I_79757 (I1358415,I1358398,I364040);
nor I_79758 (I1358432,I1358415,I364025);
not I_79759 (I1358449,I364025);
and I_79760 (I1358466,I1358449,I364022);
nand I_79761 (I1358483,I1358466,I364034);
nor I_79762 (I1358500,I1358449,I1358483);
DFFARX1 I_79763 (I1358500,I2507,I1358302,I1358267,);
not I_79764 (I1358531,I1358483);
nand I_79765 (I1358548,I1358353,I1358531);
nand I_79766 (I1358279,I1358415,I1358531);
DFFARX1 I_79767 (I1358449,I2507,I1358302,I1358294,);
not I_79768 (I1358593,I364049);
nor I_79769 (I1358610,I1358593,I364022);
nor I_79770 (I1358627,I1358610,I1358432);
DFFARX1 I_79771 (I1358627,I2507,I1358302,I1358291,);
not I_79772 (I1358658,I1358610);
DFFARX1 I_79773 (I1358658,I2507,I1358302,I1358684,);
not I_79774 (I1358692,I1358684);
nor I_79775 (I1358288,I1358692,I1358610);
nor I_79776 (I1358723,I1358593,I364031);
and I_79777 (I1358740,I1358723,I364028);
or I_79778 (I1358757,I1358740,I364022);
DFFARX1 I_79779 (I1358757,I2507,I1358302,I1358783,);
not I_79780 (I1358791,I1358783);
nand I_79781 (I1358808,I1358791,I1358531);
not I_79782 (I1358282,I1358808);
nand I_79783 (I1358276,I1358808,I1358548);
nand I_79784 (I1358273,I1358791,I1358415);
not I_79785 (I1358897,I2514);
DFFARX1 I_79786 (I1141605,I2507,I1358897,I1358923,);
DFFARX1 I_79787 (I1141617,I2507,I1358897,I1358940,);
not I_79788 (I1358948,I1358940);
nor I_79789 (I1358865,I1358923,I1358948);
DFFARX1 I_79790 (I1358948,I2507,I1358897,I1358880,);
nor I_79791 (I1358993,I1141614,I1141608);
and I_79792 (I1359010,I1358993,I1141602);
nor I_79793 (I1359027,I1359010,I1141614);
not I_79794 (I1359044,I1141614);
and I_79795 (I1359061,I1359044,I1141611);
nand I_79796 (I1359078,I1359061,I1141602);
nor I_79797 (I1359095,I1359044,I1359078);
DFFARX1 I_79798 (I1359095,I2507,I1358897,I1358862,);
not I_79799 (I1359126,I1359078);
nand I_79800 (I1359143,I1358948,I1359126);
nand I_79801 (I1358874,I1359010,I1359126);
DFFARX1 I_79802 (I1359044,I2507,I1358897,I1358889,);
not I_79803 (I1359188,I1141626);
nor I_79804 (I1359205,I1359188,I1141611);
nor I_79805 (I1359222,I1359205,I1359027);
DFFARX1 I_79806 (I1359222,I2507,I1358897,I1358886,);
not I_79807 (I1359253,I1359205);
DFFARX1 I_79808 (I1359253,I2507,I1358897,I1359279,);
not I_79809 (I1359287,I1359279);
nor I_79810 (I1358883,I1359287,I1359205);
nor I_79811 (I1359318,I1359188,I1141620);
and I_79812 (I1359335,I1359318,I1141623);
or I_79813 (I1359352,I1359335,I1141605);
DFFARX1 I_79814 (I1359352,I2507,I1358897,I1359378,);
not I_79815 (I1359386,I1359378);
nand I_79816 (I1359403,I1359386,I1359126);
not I_79817 (I1358877,I1359403);
nand I_79818 (I1358871,I1359403,I1359143);
nand I_79819 (I1358868,I1359386,I1359010);
not I_79820 (I1359492,I2514);
DFFARX1 I_79821 (I527409,I2507,I1359492,I1359518,);
DFFARX1 I_79822 (I527412,I2507,I1359492,I1359535,);
not I_79823 (I1359543,I1359535);
nor I_79824 (I1359460,I1359518,I1359543);
DFFARX1 I_79825 (I1359543,I2507,I1359492,I1359475,);
nor I_79826 (I1359588,I527415,I527433);
and I_79827 (I1359605,I1359588,I527418);
nor I_79828 (I1359622,I1359605,I527415);
not I_79829 (I1359639,I527415);
and I_79830 (I1359656,I1359639,I527427);
nand I_79831 (I1359673,I1359656,I527430);
nor I_79832 (I1359690,I1359639,I1359673);
DFFARX1 I_79833 (I1359690,I2507,I1359492,I1359457,);
not I_79834 (I1359721,I1359673);
nand I_79835 (I1359738,I1359543,I1359721);
nand I_79836 (I1359469,I1359605,I1359721);
DFFARX1 I_79837 (I1359639,I2507,I1359492,I1359484,);
not I_79838 (I1359783,I527421);
nor I_79839 (I1359800,I1359783,I527427);
nor I_79840 (I1359817,I1359800,I1359622);
DFFARX1 I_79841 (I1359817,I2507,I1359492,I1359481,);
not I_79842 (I1359848,I1359800);
DFFARX1 I_79843 (I1359848,I2507,I1359492,I1359874,);
not I_79844 (I1359882,I1359874);
nor I_79845 (I1359478,I1359882,I1359800);
nor I_79846 (I1359913,I1359783,I527409);
and I_79847 (I1359930,I1359913,I527424);
or I_79848 (I1359947,I1359930,I527412);
DFFARX1 I_79849 (I1359947,I2507,I1359492,I1359973,);
not I_79850 (I1359981,I1359973);
nand I_79851 (I1359998,I1359981,I1359721);
not I_79852 (I1359472,I1359998);
nand I_79853 (I1359466,I1359998,I1359738);
nand I_79854 (I1359463,I1359981,I1359605);
not I_79855 (I1360087,I2514);
DFFARX1 I_79856 (I356665,I2507,I1360087,I1360113,);
DFFARX1 I_79857 (I356659,I2507,I1360087,I1360130,);
not I_79858 (I1360138,I1360130);
nor I_79859 (I1360055,I1360113,I1360138);
DFFARX1 I_79860 (I1360138,I2507,I1360087,I1360070,);
nor I_79861 (I1360183,I356647,I356668);
and I_79862 (I1360200,I1360183,I356662);
nor I_79863 (I1360217,I1360200,I356647);
not I_79864 (I1360234,I356647);
and I_79865 (I1360251,I1360234,I356644);
nand I_79866 (I1360268,I1360251,I356656);
nor I_79867 (I1360285,I1360234,I1360268);
DFFARX1 I_79868 (I1360285,I2507,I1360087,I1360052,);
not I_79869 (I1360316,I1360268);
nand I_79870 (I1360333,I1360138,I1360316);
nand I_79871 (I1360064,I1360200,I1360316);
DFFARX1 I_79872 (I1360234,I2507,I1360087,I1360079,);
not I_79873 (I1360378,I356671);
nor I_79874 (I1360395,I1360378,I356644);
nor I_79875 (I1360412,I1360395,I1360217);
DFFARX1 I_79876 (I1360412,I2507,I1360087,I1360076,);
not I_79877 (I1360443,I1360395);
DFFARX1 I_79878 (I1360443,I2507,I1360087,I1360469,);
not I_79879 (I1360477,I1360469);
nor I_79880 (I1360073,I1360477,I1360395);
nor I_79881 (I1360508,I1360378,I356653);
and I_79882 (I1360525,I1360508,I356650);
or I_79883 (I1360542,I1360525,I356644);
DFFARX1 I_79884 (I1360542,I2507,I1360087,I1360568,);
not I_79885 (I1360576,I1360568);
nand I_79886 (I1360593,I1360576,I1360316);
not I_79887 (I1360067,I1360593);
nand I_79888 (I1360061,I1360593,I1360333);
nand I_79889 (I1360058,I1360576,I1360200);
not I_79890 (I1360682,I2514);
DFFARX1 I_79891 (I97041,I2507,I1360682,I1360708,);
DFFARX1 I_79892 (I97029,I2507,I1360682,I1360725,);
not I_79893 (I1360733,I1360725);
nor I_79894 (I1360650,I1360708,I1360733);
DFFARX1 I_79895 (I1360733,I2507,I1360682,I1360665,);
nor I_79896 (I1360778,I97020,I97044);
and I_79897 (I1360795,I1360778,I97023);
nor I_79898 (I1360812,I1360795,I97020);
not I_79899 (I1360829,I97020);
and I_79900 (I1360846,I1360829,I97026);
nand I_79901 (I1360863,I1360846,I97038);
nor I_79902 (I1360880,I1360829,I1360863);
DFFARX1 I_79903 (I1360880,I2507,I1360682,I1360647,);
not I_79904 (I1360911,I1360863);
nand I_79905 (I1360928,I1360733,I1360911);
nand I_79906 (I1360659,I1360795,I1360911);
DFFARX1 I_79907 (I1360829,I2507,I1360682,I1360674,);
not I_79908 (I1360973,I97020);
nor I_79909 (I1360990,I1360973,I97026);
nor I_79910 (I1361007,I1360990,I1360812);
DFFARX1 I_79911 (I1361007,I2507,I1360682,I1360671,);
not I_79912 (I1361038,I1360990);
DFFARX1 I_79913 (I1361038,I2507,I1360682,I1361064,);
not I_79914 (I1361072,I1361064);
nor I_79915 (I1360668,I1361072,I1360990);
nor I_79916 (I1361103,I1360973,I97023);
and I_79917 (I1361120,I1361103,I97032);
or I_79918 (I1361137,I1361120,I97035);
DFFARX1 I_79919 (I1361137,I2507,I1360682,I1361163,);
not I_79920 (I1361171,I1361163);
nand I_79921 (I1361188,I1361171,I1360911);
not I_79922 (I1360662,I1361188);
nand I_79923 (I1360656,I1361188,I1360928);
nand I_79924 (I1360653,I1361171,I1360795);
not I_79925 (I1361277,I2514);
DFFARX1 I_79926 (I1010714,I2507,I1361277,I1361303,);
DFFARX1 I_79927 (I1010705,I2507,I1361277,I1361320,);
not I_79928 (I1361328,I1361320);
nor I_79929 (I1361245,I1361303,I1361328);
DFFARX1 I_79930 (I1361328,I2507,I1361277,I1361260,);
nor I_79931 (I1361373,I1010711,I1010720);
and I_79932 (I1361390,I1361373,I1010723);
nor I_79933 (I1361407,I1361390,I1010711);
not I_79934 (I1361424,I1010711);
and I_79935 (I1361441,I1361424,I1010702);
nand I_79936 (I1361458,I1361441,I1010708);
nor I_79937 (I1361475,I1361424,I1361458);
DFFARX1 I_79938 (I1361475,I2507,I1361277,I1361242,);
not I_79939 (I1361506,I1361458);
nand I_79940 (I1361523,I1361328,I1361506);
nand I_79941 (I1361254,I1361390,I1361506);
DFFARX1 I_79942 (I1361424,I2507,I1361277,I1361269,);
not I_79943 (I1361568,I1010717);
nor I_79944 (I1361585,I1361568,I1010702);
nor I_79945 (I1361602,I1361585,I1361407);
DFFARX1 I_79946 (I1361602,I2507,I1361277,I1361266,);
not I_79947 (I1361633,I1361585);
DFFARX1 I_79948 (I1361633,I2507,I1361277,I1361659,);
not I_79949 (I1361667,I1361659);
nor I_79950 (I1361263,I1361667,I1361585);
nor I_79951 (I1361698,I1361568,I1010702);
and I_79952 (I1361715,I1361698,I1010705);
or I_79953 (I1361732,I1361715,I1010708);
DFFARX1 I_79954 (I1361732,I2507,I1361277,I1361758,);
not I_79955 (I1361766,I1361758);
nand I_79956 (I1361783,I1361766,I1361506);
not I_79957 (I1361257,I1361783);
nand I_79958 (I1361251,I1361783,I1361523);
nand I_79959 (I1361248,I1361766,I1361390);
not I_79960 (I1361872,I2514);
DFFARX1 I_79961 (I858119,I2507,I1361872,I1361898,);
DFFARX1 I_79962 (I858116,I2507,I1361872,I1361915,);
not I_79963 (I1361923,I1361915);
nor I_79964 (I1361840,I1361898,I1361923);
DFFARX1 I_79965 (I1361923,I2507,I1361872,I1361855,);
nor I_79966 (I1361968,I858131,I858113);
and I_79967 (I1361985,I1361968,I858110);
nor I_79968 (I1362002,I1361985,I858131);
not I_79969 (I1362019,I858131);
and I_79970 (I1362036,I1362019,I858116);
nand I_79971 (I1362053,I1362036,I858128);
nor I_79972 (I1362070,I1362019,I1362053);
DFFARX1 I_79973 (I1362070,I2507,I1361872,I1361837,);
not I_79974 (I1362101,I1362053);
nand I_79975 (I1362118,I1361923,I1362101);
nand I_79976 (I1361849,I1361985,I1362101);
DFFARX1 I_79977 (I1362019,I2507,I1361872,I1361864,);
not I_79978 (I1362163,I858122);
nor I_79979 (I1362180,I1362163,I858116);
nor I_79980 (I1362197,I1362180,I1362002);
DFFARX1 I_79981 (I1362197,I2507,I1361872,I1361861,);
not I_79982 (I1362228,I1362180);
DFFARX1 I_79983 (I1362228,I2507,I1361872,I1362254,);
not I_79984 (I1362262,I1362254);
nor I_79985 (I1361858,I1362262,I1362180);
nor I_79986 (I1362293,I1362163,I858110);
and I_79987 (I1362310,I1362293,I858125);
or I_79988 (I1362327,I1362310,I858113);
DFFARX1 I_79989 (I1362327,I2507,I1361872,I1362353,);
not I_79990 (I1362361,I1362353);
nand I_79991 (I1362378,I1362361,I1362101);
not I_79992 (I1361852,I1362378);
nand I_79993 (I1361846,I1362378,I1362118);
nand I_79994 (I1361843,I1362361,I1361985);
not I_79995 (I1362467,I2514);
DFFARX1 I_79996 (I818067,I2507,I1362467,I1362493,);
DFFARX1 I_79997 (I818064,I2507,I1362467,I1362510,);
not I_79998 (I1362518,I1362510);
nor I_79999 (I1362435,I1362493,I1362518);
DFFARX1 I_80000 (I1362518,I2507,I1362467,I1362450,);
nor I_80001 (I1362563,I818079,I818061);
and I_80002 (I1362580,I1362563,I818058);
nor I_80003 (I1362597,I1362580,I818079);
not I_80004 (I1362614,I818079);
and I_80005 (I1362631,I1362614,I818064);
nand I_80006 (I1362648,I1362631,I818076);
nor I_80007 (I1362665,I1362614,I1362648);
DFFARX1 I_80008 (I1362665,I2507,I1362467,I1362432,);
not I_80009 (I1362696,I1362648);
nand I_80010 (I1362713,I1362518,I1362696);
nand I_80011 (I1362444,I1362580,I1362696);
DFFARX1 I_80012 (I1362614,I2507,I1362467,I1362459,);
not I_80013 (I1362758,I818070);
nor I_80014 (I1362775,I1362758,I818064);
nor I_80015 (I1362792,I1362775,I1362597);
DFFARX1 I_80016 (I1362792,I2507,I1362467,I1362456,);
not I_80017 (I1362823,I1362775);
DFFARX1 I_80018 (I1362823,I2507,I1362467,I1362849,);
not I_80019 (I1362857,I1362849);
nor I_80020 (I1362453,I1362857,I1362775);
nor I_80021 (I1362888,I1362758,I818058);
and I_80022 (I1362905,I1362888,I818073);
or I_80023 (I1362922,I1362905,I818061);
DFFARX1 I_80024 (I1362922,I2507,I1362467,I1362948,);
not I_80025 (I1362956,I1362948);
nand I_80026 (I1362973,I1362956,I1362696);
not I_80027 (I1362447,I1362973);
nand I_80028 (I1362441,I1362973,I1362713);
nand I_80029 (I1362438,I1362956,I1362580);
not I_80030 (I1363062,I2514);
DFFARX1 I_80031 (I1273268,I2507,I1363062,I1363088,);
DFFARX1 I_80032 (I1273259,I2507,I1363062,I1363105,);
not I_80033 (I1363113,I1363105);
nor I_80034 (I1363030,I1363088,I1363113);
DFFARX1 I_80035 (I1363113,I2507,I1363062,I1363045,);
nor I_80036 (I1363158,I1273250,I1273265);
and I_80037 (I1363175,I1363158,I1273253);
nor I_80038 (I1363192,I1363175,I1273250);
not I_80039 (I1363209,I1273250);
and I_80040 (I1363226,I1363209,I1273256);
nand I_80041 (I1363243,I1363226,I1273274);
nor I_80042 (I1363260,I1363209,I1363243);
DFFARX1 I_80043 (I1363260,I2507,I1363062,I1363027,);
not I_80044 (I1363291,I1363243);
nand I_80045 (I1363308,I1363113,I1363291);
nand I_80046 (I1363039,I1363175,I1363291);
DFFARX1 I_80047 (I1363209,I2507,I1363062,I1363054,);
not I_80048 (I1363353,I1273250);
nor I_80049 (I1363370,I1363353,I1273256);
nor I_80050 (I1363387,I1363370,I1363192);
DFFARX1 I_80051 (I1363387,I2507,I1363062,I1363051,);
not I_80052 (I1363418,I1363370);
DFFARX1 I_80053 (I1363418,I2507,I1363062,I1363444,);
not I_80054 (I1363452,I1363444);
nor I_80055 (I1363048,I1363452,I1363370);
nor I_80056 (I1363483,I1363353,I1273253);
and I_80057 (I1363500,I1363483,I1273262);
or I_80058 (I1363517,I1363500,I1273271);
DFFARX1 I_80059 (I1363517,I2507,I1363062,I1363543,);
not I_80060 (I1363551,I1363543);
nand I_80061 (I1363568,I1363551,I1363291);
not I_80062 (I1363042,I1363568);
nand I_80063 (I1363036,I1363568,I1363308);
nand I_80064 (I1363033,I1363551,I1363175);
not I_80065 (I1363657,I2514);
DFFARX1 I_80066 (I1087273,I2507,I1363657,I1363683,);
DFFARX1 I_80067 (I1087285,I2507,I1363657,I1363700,);
not I_80068 (I1363708,I1363700);
nor I_80069 (I1363625,I1363683,I1363708);
DFFARX1 I_80070 (I1363708,I2507,I1363657,I1363640,);
nor I_80071 (I1363753,I1087282,I1087276);
and I_80072 (I1363770,I1363753,I1087270);
nor I_80073 (I1363787,I1363770,I1087282);
not I_80074 (I1363804,I1087282);
and I_80075 (I1363821,I1363804,I1087279);
nand I_80076 (I1363838,I1363821,I1087270);
nor I_80077 (I1363855,I1363804,I1363838);
DFFARX1 I_80078 (I1363855,I2507,I1363657,I1363622,);
not I_80079 (I1363886,I1363838);
nand I_80080 (I1363903,I1363708,I1363886);
nand I_80081 (I1363634,I1363770,I1363886);
DFFARX1 I_80082 (I1363804,I2507,I1363657,I1363649,);
not I_80083 (I1363948,I1087294);
nor I_80084 (I1363965,I1363948,I1087279);
nor I_80085 (I1363982,I1363965,I1363787);
DFFARX1 I_80086 (I1363982,I2507,I1363657,I1363646,);
not I_80087 (I1364013,I1363965);
DFFARX1 I_80088 (I1364013,I2507,I1363657,I1364039,);
not I_80089 (I1364047,I1364039);
nor I_80090 (I1363643,I1364047,I1363965);
nor I_80091 (I1364078,I1363948,I1087288);
and I_80092 (I1364095,I1364078,I1087291);
or I_80093 (I1364112,I1364095,I1087273);
DFFARX1 I_80094 (I1364112,I2507,I1363657,I1364138,);
not I_80095 (I1364146,I1364138);
nand I_80096 (I1364163,I1364146,I1363886);
not I_80097 (I1363637,I1364163);
nand I_80098 (I1363631,I1364163,I1363903);
nand I_80099 (I1363628,I1364146,I1363770);
not I_80100 (I1364252,I2514);
DFFARX1 I_80101 (I996751,I2507,I1364252,I1364278,);
DFFARX1 I_80102 (I996769,I2507,I1364252,I1364295,);
not I_80103 (I1364303,I1364295);
nor I_80104 (I1364220,I1364278,I1364303);
DFFARX1 I_80105 (I1364303,I2507,I1364252,I1364235,);
nor I_80106 (I1364348,I996748,I996760);
and I_80107 (I1364365,I1364348,I996745);
nor I_80108 (I1364382,I1364365,I996748);
not I_80109 (I1364399,I996748);
and I_80110 (I1364416,I1364399,I996754);
nand I_80111 (I1364433,I1364416,I996766);
nor I_80112 (I1364450,I1364399,I1364433);
DFFARX1 I_80113 (I1364450,I2507,I1364252,I1364217,);
not I_80114 (I1364481,I1364433);
nand I_80115 (I1364498,I1364303,I1364481);
nand I_80116 (I1364229,I1364365,I1364481);
DFFARX1 I_80117 (I1364399,I2507,I1364252,I1364244,);
not I_80118 (I1364543,I996757);
nor I_80119 (I1364560,I1364543,I996754);
nor I_80120 (I1364577,I1364560,I1364382);
DFFARX1 I_80121 (I1364577,I2507,I1364252,I1364241,);
not I_80122 (I1364608,I1364560);
DFFARX1 I_80123 (I1364608,I2507,I1364252,I1364634,);
not I_80124 (I1364642,I1364634);
nor I_80125 (I1364238,I1364642,I1364560);
nor I_80126 (I1364673,I1364543,I996745);
and I_80127 (I1364690,I1364673,I996772);
or I_80128 (I1364707,I1364690,I996763);
DFFARX1 I_80129 (I1364707,I2507,I1364252,I1364733,);
not I_80130 (I1364741,I1364733);
nand I_80131 (I1364758,I1364741,I1364481);
not I_80132 (I1364232,I1364758);
nand I_80133 (I1364226,I1364758,I1364498);
nand I_80134 (I1364223,I1364741,I1364365);
not I_80135 (I1364847,I2514);
DFFARX1 I_80136 (I275507,I2507,I1364847,I1364873,);
DFFARX1 I_80137 (I275501,I2507,I1364847,I1364890,);
not I_80138 (I1364898,I1364890);
nor I_80139 (I1364815,I1364873,I1364898);
DFFARX1 I_80140 (I1364898,I2507,I1364847,I1364830,);
nor I_80141 (I1364943,I275489,I275510);
and I_80142 (I1364960,I1364943,I275504);
nor I_80143 (I1364977,I1364960,I275489);
not I_80144 (I1364994,I275489);
and I_80145 (I1365011,I1364994,I275486);
nand I_80146 (I1365028,I1365011,I275498);
nor I_80147 (I1365045,I1364994,I1365028);
DFFARX1 I_80148 (I1365045,I2507,I1364847,I1364812,);
not I_80149 (I1365076,I1365028);
nand I_80150 (I1365093,I1364898,I1365076);
nand I_80151 (I1364824,I1364960,I1365076);
DFFARX1 I_80152 (I1364994,I2507,I1364847,I1364839,);
not I_80153 (I1365138,I275513);
nor I_80154 (I1365155,I1365138,I275486);
nor I_80155 (I1365172,I1365155,I1364977);
DFFARX1 I_80156 (I1365172,I2507,I1364847,I1364836,);
not I_80157 (I1365203,I1365155);
DFFARX1 I_80158 (I1365203,I2507,I1364847,I1365229,);
not I_80159 (I1365237,I1365229);
nor I_80160 (I1364833,I1365237,I1365155);
nor I_80161 (I1365268,I1365138,I275495);
and I_80162 (I1365285,I1365268,I275492);
or I_80163 (I1365302,I1365285,I275486);
DFFARX1 I_80164 (I1365302,I2507,I1364847,I1365328,);
not I_80165 (I1365336,I1365328);
nand I_80166 (I1365353,I1365336,I1365076);
not I_80167 (I1364827,I1365353);
nand I_80168 (I1364821,I1365353,I1365093);
nand I_80169 (I1364818,I1365336,I1364960);
not I_80170 (I1365442,I2514);
DFFARX1 I_80171 (I442511,I2507,I1365442,I1365468,);
DFFARX1 I_80172 (I442517,I2507,I1365442,I1365485,);
not I_80173 (I1365493,I1365485);
nor I_80174 (I1365410,I1365468,I1365493);
DFFARX1 I_80175 (I1365493,I2507,I1365442,I1365425,);
nor I_80176 (I1365538,I442526,I442511);
and I_80177 (I1365555,I1365538,I442538);
nor I_80178 (I1365572,I1365555,I442526);
not I_80179 (I1365589,I442526);
and I_80180 (I1365606,I1365589,I442514);
nand I_80181 (I1365623,I1365606,I442535);
nor I_80182 (I1365640,I1365589,I1365623);
DFFARX1 I_80183 (I1365640,I2507,I1365442,I1365407,);
not I_80184 (I1365671,I1365623);
nand I_80185 (I1365688,I1365493,I1365671);
nand I_80186 (I1365419,I1365555,I1365671);
DFFARX1 I_80187 (I1365589,I2507,I1365442,I1365434,);
not I_80188 (I1365733,I442523);
nor I_80189 (I1365750,I1365733,I442514);
nor I_80190 (I1365767,I1365750,I1365572);
DFFARX1 I_80191 (I1365767,I2507,I1365442,I1365431,);
not I_80192 (I1365798,I1365750);
DFFARX1 I_80193 (I1365798,I2507,I1365442,I1365824,);
not I_80194 (I1365832,I1365824);
nor I_80195 (I1365428,I1365832,I1365750);
nor I_80196 (I1365863,I1365733,I442520);
and I_80197 (I1365880,I1365863,I442532);
or I_80198 (I1365897,I1365880,I442529);
DFFARX1 I_80199 (I1365897,I2507,I1365442,I1365923,);
not I_80200 (I1365931,I1365923);
nand I_80201 (I1365948,I1365931,I1365671);
not I_80202 (I1365422,I1365948);
nand I_80203 (I1365416,I1365948,I1365688);
nand I_80204 (I1365413,I1365931,I1365555);
not I_80205 (I1366037,I2514);
DFFARX1 I_80206 (I742871,I2507,I1366037,I1366063,);
DFFARX1 I_80207 (I742853,I2507,I1366037,I1366080,);
not I_80208 (I1366088,I1366080);
nor I_80209 (I1366005,I1366063,I1366088);
DFFARX1 I_80210 (I1366088,I2507,I1366037,I1366020,);
nor I_80211 (I1366133,I742859,I742862);
and I_80212 (I1366150,I1366133,I742850);
nor I_80213 (I1366167,I1366150,I742859);
not I_80214 (I1366184,I742859);
and I_80215 (I1366201,I1366184,I742868);
nand I_80216 (I1366218,I1366201,I742856);
nor I_80217 (I1366235,I1366184,I1366218);
DFFARX1 I_80218 (I1366235,I2507,I1366037,I1366002,);
not I_80219 (I1366266,I1366218);
nand I_80220 (I1366283,I1366088,I1366266);
nand I_80221 (I1366014,I1366150,I1366266);
DFFARX1 I_80222 (I1366184,I2507,I1366037,I1366029,);
not I_80223 (I1366328,I742853);
nor I_80224 (I1366345,I1366328,I742868);
nor I_80225 (I1366362,I1366345,I1366167);
DFFARX1 I_80226 (I1366362,I2507,I1366037,I1366026,);
not I_80227 (I1366393,I1366345);
DFFARX1 I_80228 (I1366393,I2507,I1366037,I1366419,);
not I_80229 (I1366427,I1366419);
nor I_80230 (I1366023,I1366427,I1366345);
nor I_80231 (I1366458,I1366328,I742865);
and I_80232 (I1366475,I1366458,I742874);
or I_80233 (I1366492,I1366475,I742850);
DFFARX1 I_80234 (I1366492,I2507,I1366037,I1366518,);
not I_80235 (I1366526,I1366518);
nand I_80236 (I1366543,I1366526,I1366266);
not I_80237 (I1366017,I1366543);
nand I_80238 (I1366011,I1366543,I1366283);
nand I_80239 (I1366008,I1366526,I1366150);
not I_80240 (I1366632,I2514);
DFFARX1 I_80241 (I366678,I2507,I1366632,I1366658,);
DFFARX1 I_80242 (I366672,I2507,I1366632,I1366675,);
not I_80243 (I1366683,I1366675);
nor I_80244 (I1366600,I1366658,I1366683);
DFFARX1 I_80245 (I1366683,I2507,I1366632,I1366615,);
nor I_80246 (I1366728,I366660,I366681);
and I_80247 (I1366745,I1366728,I366675);
nor I_80248 (I1366762,I1366745,I366660);
not I_80249 (I1366779,I366660);
and I_80250 (I1366796,I1366779,I366657);
nand I_80251 (I1366813,I1366796,I366669);
nor I_80252 (I1366830,I1366779,I1366813);
DFFARX1 I_80253 (I1366830,I2507,I1366632,I1366597,);
not I_80254 (I1366861,I1366813);
nand I_80255 (I1366878,I1366683,I1366861);
nand I_80256 (I1366609,I1366745,I1366861);
DFFARX1 I_80257 (I1366779,I2507,I1366632,I1366624,);
not I_80258 (I1366923,I366684);
nor I_80259 (I1366940,I1366923,I366657);
nor I_80260 (I1366957,I1366940,I1366762);
DFFARX1 I_80261 (I1366957,I2507,I1366632,I1366621,);
not I_80262 (I1366988,I1366940);
DFFARX1 I_80263 (I1366988,I2507,I1366632,I1367014,);
not I_80264 (I1367022,I1367014);
nor I_80265 (I1366618,I1367022,I1366940);
nor I_80266 (I1367053,I1366923,I366666);
and I_80267 (I1367070,I1367053,I366663);
or I_80268 (I1367087,I1367070,I366657);
DFFARX1 I_80269 (I1367087,I2507,I1366632,I1367113,);
not I_80270 (I1367121,I1367113);
nand I_80271 (I1367138,I1367121,I1366861);
not I_80272 (I1366612,I1367138);
nand I_80273 (I1366606,I1367138,I1366878);
nand I_80274 (I1366603,I1367121,I1366745);
not I_80275 (I1367227,I2514);
DFFARX1 I_80276 (I150230,I2507,I1367227,I1367253,);
DFFARX1 I_80277 (I150233,I2507,I1367227,I1367270,);
not I_80278 (I1367278,I1367270);
nor I_80279 (I1367195,I1367253,I1367278);
DFFARX1 I_80280 (I1367278,I2507,I1367227,I1367210,);
nor I_80281 (I1367323,I150239,I150233);
and I_80282 (I1367340,I1367323,I150236);
nor I_80283 (I1367357,I1367340,I150239);
not I_80284 (I1367374,I150239);
and I_80285 (I1367391,I1367374,I150230);
nand I_80286 (I1367408,I1367391,I150248);
nor I_80287 (I1367425,I1367374,I1367408);
DFFARX1 I_80288 (I1367425,I2507,I1367227,I1367192,);
not I_80289 (I1367456,I1367408);
nand I_80290 (I1367473,I1367278,I1367456);
nand I_80291 (I1367204,I1367340,I1367456);
DFFARX1 I_80292 (I1367374,I2507,I1367227,I1367219,);
not I_80293 (I1367518,I150242);
nor I_80294 (I1367535,I1367518,I150230);
nor I_80295 (I1367552,I1367535,I1367357);
DFFARX1 I_80296 (I1367552,I2507,I1367227,I1367216,);
not I_80297 (I1367583,I1367535);
DFFARX1 I_80298 (I1367583,I2507,I1367227,I1367609,);
not I_80299 (I1367617,I1367609);
nor I_80300 (I1367213,I1367617,I1367535);
nor I_80301 (I1367648,I1367518,I150245);
and I_80302 (I1367665,I1367648,I150251);
or I_80303 (I1367682,I1367665,I150254);
DFFARX1 I_80304 (I1367682,I2507,I1367227,I1367708,);
not I_80305 (I1367716,I1367708);
nand I_80306 (I1367733,I1367716,I1367456);
not I_80307 (I1367207,I1367733);
nand I_80308 (I1367201,I1367733,I1367473);
nand I_80309 (I1367198,I1367716,I1367340);
not I_80310 (I1367822,I2514);
DFFARX1 I_80311 (I288155,I2507,I1367822,I1367848,);
DFFARX1 I_80312 (I288149,I2507,I1367822,I1367865,);
not I_80313 (I1367873,I1367865);
nor I_80314 (I1367790,I1367848,I1367873);
DFFARX1 I_80315 (I1367873,I2507,I1367822,I1367805,);
nor I_80316 (I1367918,I288137,I288158);
and I_80317 (I1367935,I1367918,I288152);
nor I_80318 (I1367952,I1367935,I288137);
not I_80319 (I1367969,I288137);
and I_80320 (I1367986,I1367969,I288134);
nand I_80321 (I1368003,I1367986,I288146);
nor I_80322 (I1368020,I1367969,I1368003);
DFFARX1 I_80323 (I1368020,I2507,I1367822,I1367787,);
not I_80324 (I1368051,I1368003);
nand I_80325 (I1368068,I1367873,I1368051);
nand I_80326 (I1367799,I1367935,I1368051);
DFFARX1 I_80327 (I1367969,I2507,I1367822,I1367814,);
not I_80328 (I1368113,I288161);
nor I_80329 (I1368130,I1368113,I288134);
nor I_80330 (I1368147,I1368130,I1367952);
DFFARX1 I_80331 (I1368147,I2507,I1367822,I1367811,);
not I_80332 (I1368178,I1368130);
DFFARX1 I_80333 (I1368178,I2507,I1367822,I1368204,);
not I_80334 (I1368212,I1368204);
nor I_80335 (I1367808,I1368212,I1368130);
nor I_80336 (I1368243,I1368113,I288143);
and I_80337 (I1368260,I1368243,I288140);
or I_80338 (I1368277,I1368260,I288134);
DFFARX1 I_80339 (I1368277,I2507,I1367822,I1368303,);
not I_80340 (I1368311,I1368303);
nand I_80341 (I1368328,I1368311,I1368051);
not I_80342 (I1367802,I1368328);
nand I_80343 (I1367796,I1368328,I1368068);
nand I_80344 (I1367793,I1368311,I1367935);
not I_80345 (I1368417,I2514);
DFFARX1 I_80346 (I679291,I2507,I1368417,I1368443,);
DFFARX1 I_80347 (I679273,I2507,I1368417,I1368460,);
not I_80348 (I1368468,I1368460);
nor I_80349 (I1368385,I1368443,I1368468);
DFFARX1 I_80350 (I1368468,I2507,I1368417,I1368400,);
nor I_80351 (I1368513,I679279,I679282);
and I_80352 (I1368530,I1368513,I679270);
nor I_80353 (I1368547,I1368530,I679279);
not I_80354 (I1368564,I679279);
and I_80355 (I1368581,I1368564,I679288);
nand I_80356 (I1368598,I1368581,I679276);
nor I_80357 (I1368615,I1368564,I1368598);
DFFARX1 I_80358 (I1368615,I2507,I1368417,I1368382,);
not I_80359 (I1368646,I1368598);
nand I_80360 (I1368663,I1368468,I1368646);
nand I_80361 (I1368394,I1368530,I1368646);
DFFARX1 I_80362 (I1368564,I2507,I1368417,I1368409,);
not I_80363 (I1368708,I679273);
nor I_80364 (I1368725,I1368708,I679288);
nor I_80365 (I1368742,I1368725,I1368547);
DFFARX1 I_80366 (I1368742,I2507,I1368417,I1368406,);
not I_80367 (I1368773,I1368725);
DFFARX1 I_80368 (I1368773,I2507,I1368417,I1368799,);
not I_80369 (I1368807,I1368799);
nor I_80370 (I1368403,I1368807,I1368725);
nor I_80371 (I1368838,I1368708,I679285);
and I_80372 (I1368855,I1368838,I679294);
or I_80373 (I1368872,I1368855,I679270);
DFFARX1 I_80374 (I1368872,I2507,I1368417,I1368898,);
not I_80375 (I1368906,I1368898);
nand I_80376 (I1368923,I1368906,I1368646);
not I_80377 (I1368397,I1368923);
nand I_80378 (I1368391,I1368923,I1368663);
nand I_80379 (I1368388,I1368906,I1368530);
not I_80380 (I1369012,I2514);
DFFARX1 I_80381 (I87555,I2507,I1369012,I1369038,);
DFFARX1 I_80382 (I87543,I2507,I1369012,I1369055,);
not I_80383 (I1369063,I1369055);
nor I_80384 (I1368980,I1369038,I1369063);
DFFARX1 I_80385 (I1369063,I2507,I1369012,I1368995,);
nor I_80386 (I1369108,I87534,I87558);
and I_80387 (I1369125,I1369108,I87537);
nor I_80388 (I1369142,I1369125,I87534);
not I_80389 (I1369159,I87534);
and I_80390 (I1369176,I1369159,I87540);
nand I_80391 (I1369193,I1369176,I87552);
nor I_80392 (I1369210,I1369159,I1369193);
DFFARX1 I_80393 (I1369210,I2507,I1369012,I1368977,);
not I_80394 (I1369241,I1369193);
nand I_80395 (I1369258,I1369063,I1369241);
nand I_80396 (I1368989,I1369125,I1369241);
DFFARX1 I_80397 (I1369159,I2507,I1369012,I1369004,);
not I_80398 (I1369303,I87534);
nor I_80399 (I1369320,I1369303,I87540);
nor I_80400 (I1369337,I1369320,I1369142);
DFFARX1 I_80401 (I1369337,I2507,I1369012,I1369001,);
not I_80402 (I1369368,I1369320);
DFFARX1 I_80403 (I1369368,I2507,I1369012,I1369394,);
not I_80404 (I1369402,I1369394);
nor I_80405 (I1368998,I1369402,I1369320);
nor I_80406 (I1369433,I1369303,I87537);
and I_80407 (I1369450,I1369433,I87546);
or I_80408 (I1369467,I1369450,I87549);
DFFARX1 I_80409 (I1369467,I2507,I1369012,I1369493,);
not I_80410 (I1369501,I1369493);
nand I_80411 (I1369518,I1369501,I1369241);
not I_80412 (I1368992,I1369518);
nand I_80413 (I1368986,I1369518,I1369258);
nand I_80414 (I1368983,I1369501,I1369125);
not I_80415 (I1369607,I2514);
DFFARX1 I_80416 (I1127733,I2507,I1369607,I1369633,);
DFFARX1 I_80417 (I1127745,I2507,I1369607,I1369650,);
not I_80418 (I1369658,I1369650);
nor I_80419 (I1369575,I1369633,I1369658);
DFFARX1 I_80420 (I1369658,I2507,I1369607,I1369590,);
nor I_80421 (I1369703,I1127742,I1127736);
and I_80422 (I1369720,I1369703,I1127730);
nor I_80423 (I1369737,I1369720,I1127742);
not I_80424 (I1369754,I1127742);
and I_80425 (I1369771,I1369754,I1127739);
nand I_80426 (I1369788,I1369771,I1127730);
nor I_80427 (I1369805,I1369754,I1369788);
DFFARX1 I_80428 (I1369805,I2507,I1369607,I1369572,);
not I_80429 (I1369836,I1369788);
nand I_80430 (I1369853,I1369658,I1369836);
nand I_80431 (I1369584,I1369720,I1369836);
DFFARX1 I_80432 (I1369754,I2507,I1369607,I1369599,);
not I_80433 (I1369898,I1127754);
nor I_80434 (I1369915,I1369898,I1127739);
nor I_80435 (I1369932,I1369915,I1369737);
DFFARX1 I_80436 (I1369932,I2507,I1369607,I1369596,);
not I_80437 (I1369963,I1369915);
DFFARX1 I_80438 (I1369963,I2507,I1369607,I1369989,);
not I_80439 (I1369997,I1369989);
nor I_80440 (I1369593,I1369997,I1369915);
nor I_80441 (I1370028,I1369898,I1127748);
and I_80442 (I1370045,I1370028,I1127751);
or I_80443 (I1370062,I1370045,I1127733);
DFFARX1 I_80444 (I1370062,I2507,I1369607,I1370088,);
not I_80445 (I1370096,I1370088);
nand I_80446 (I1370113,I1370096,I1369836);
not I_80447 (I1369587,I1370113);
nand I_80448 (I1369581,I1370113,I1369853);
nand I_80449 (I1369578,I1370096,I1369720);
not I_80450 (I1370202,I2514);
DFFARX1 I_80451 (I471887,I2507,I1370202,I1370228,);
DFFARX1 I_80452 (I471893,I2507,I1370202,I1370245,);
not I_80453 (I1370253,I1370245);
nor I_80454 (I1370170,I1370228,I1370253);
DFFARX1 I_80455 (I1370253,I2507,I1370202,I1370185,);
nor I_80456 (I1370298,I471902,I471887);
and I_80457 (I1370315,I1370298,I471914);
nor I_80458 (I1370332,I1370315,I471902);
not I_80459 (I1370349,I471902);
and I_80460 (I1370366,I1370349,I471890);
nand I_80461 (I1370383,I1370366,I471911);
nor I_80462 (I1370400,I1370349,I1370383);
DFFARX1 I_80463 (I1370400,I2507,I1370202,I1370167,);
not I_80464 (I1370431,I1370383);
nand I_80465 (I1370448,I1370253,I1370431);
nand I_80466 (I1370179,I1370315,I1370431);
DFFARX1 I_80467 (I1370349,I2507,I1370202,I1370194,);
not I_80468 (I1370493,I471899);
nor I_80469 (I1370510,I1370493,I471890);
nor I_80470 (I1370527,I1370510,I1370332);
DFFARX1 I_80471 (I1370527,I2507,I1370202,I1370191,);
not I_80472 (I1370558,I1370510);
DFFARX1 I_80473 (I1370558,I2507,I1370202,I1370584,);
not I_80474 (I1370592,I1370584);
nor I_80475 (I1370188,I1370592,I1370510);
nor I_80476 (I1370623,I1370493,I471896);
and I_80477 (I1370640,I1370623,I471908);
or I_80478 (I1370657,I1370640,I471905);
DFFARX1 I_80479 (I1370657,I2507,I1370202,I1370683,);
not I_80480 (I1370691,I1370683);
nand I_80481 (I1370708,I1370691,I1370431);
not I_80482 (I1370182,I1370708);
nand I_80483 (I1370176,I1370708,I1370448);
nand I_80484 (I1370173,I1370691,I1370315);
not I_80485 (I1370797,I2514);
DFFARX1 I_80486 (I71218,I2507,I1370797,I1370823,);
DFFARX1 I_80487 (I71206,I2507,I1370797,I1370840,);
not I_80488 (I1370848,I1370840);
nor I_80489 (I1370765,I1370823,I1370848);
DFFARX1 I_80490 (I1370848,I2507,I1370797,I1370780,);
nor I_80491 (I1370893,I71197,I71221);
and I_80492 (I1370910,I1370893,I71200);
nor I_80493 (I1370927,I1370910,I71197);
not I_80494 (I1370944,I71197);
and I_80495 (I1370961,I1370944,I71203);
nand I_80496 (I1370978,I1370961,I71215);
nor I_80497 (I1370995,I1370944,I1370978);
DFFARX1 I_80498 (I1370995,I2507,I1370797,I1370762,);
not I_80499 (I1371026,I1370978);
nand I_80500 (I1371043,I1370848,I1371026);
nand I_80501 (I1370774,I1370910,I1371026);
DFFARX1 I_80502 (I1370944,I2507,I1370797,I1370789,);
not I_80503 (I1371088,I71197);
nor I_80504 (I1371105,I1371088,I71203);
nor I_80505 (I1371122,I1371105,I1370927);
DFFARX1 I_80506 (I1371122,I2507,I1370797,I1370786,);
not I_80507 (I1371153,I1371105);
DFFARX1 I_80508 (I1371153,I2507,I1370797,I1371179,);
not I_80509 (I1371187,I1371179);
nor I_80510 (I1370783,I1371187,I1371105);
nor I_80511 (I1371218,I1371088,I71200);
and I_80512 (I1371235,I1371218,I71209);
or I_80513 (I1371252,I1371235,I71212);
DFFARX1 I_80514 (I1371252,I2507,I1370797,I1371278,);
not I_80515 (I1371286,I1371278);
nand I_80516 (I1371303,I1371286,I1371026);
not I_80517 (I1370777,I1371303);
nand I_80518 (I1370771,I1371303,I1371043);
nand I_80519 (I1370768,I1371286,I1370910);
not I_80520 (I1371392,I2514);
DFFARX1 I_80521 (I425103,I2507,I1371392,I1371418,);
DFFARX1 I_80522 (I425109,I2507,I1371392,I1371435,);
not I_80523 (I1371443,I1371435);
nor I_80524 (I1371360,I1371418,I1371443);
DFFARX1 I_80525 (I1371443,I2507,I1371392,I1371375,);
nor I_80526 (I1371488,I425118,I425103);
and I_80527 (I1371505,I1371488,I425130);
nor I_80528 (I1371522,I1371505,I425118);
not I_80529 (I1371539,I425118);
and I_80530 (I1371556,I1371539,I425106);
nand I_80531 (I1371573,I1371556,I425127);
nor I_80532 (I1371590,I1371539,I1371573);
DFFARX1 I_80533 (I1371590,I2507,I1371392,I1371357,);
not I_80534 (I1371621,I1371573);
nand I_80535 (I1371638,I1371443,I1371621);
nand I_80536 (I1371369,I1371505,I1371621);
DFFARX1 I_80537 (I1371539,I2507,I1371392,I1371384,);
not I_80538 (I1371683,I425115);
nor I_80539 (I1371700,I1371683,I425106);
nor I_80540 (I1371717,I1371700,I1371522);
DFFARX1 I_80541 (I1371717,I2507,I1371392,I1371381,);
not I_80542 (I1371748,I1371700);
DFFARX1 I_80543 (I1371748,I2507,I1371392,I1371774,);
not I_80544 (I1371782,I1371774);
nor I_80545 (I1371378,I1371782,I1371700);
nor I_80546 (I1371813,I1371683,I425112);
and I_80547 (I1371830,I1371813,I425124);
or I_80548 (I1371847,I1371830,I425121);
DFFARX1 I_80549 (I1371847,I2507,I1371392,I1371873,);
not I_80550 (I1371881,I1371873);
nand I_80551 (I1371898,I1371881,I1371621);
not I_80552 (I1371372,I1371898);
nand I_80553 (I1371366,I1371898,I1371638);
nand I_80554 (I1371363,I1371881,I1371505);
not I_80555 (I1371987,I2514);
DFFARX1 I_80556 (I618601,I2507,I1371987,I1372013,);
DFFARX1 I_80557 (I618595,I2507,I1371987,I1372030,);
not I_80558 (I1372038,I1372030);
nor I_80559 (I1371955,I1372013,I1372038);
DFFARX1 I_80560 (I1372038,I2507,I1371987,I1371970,);
nor I_80561 (I1372083,I618592,I618583);
and I_80562 (I1372100,I1372083,I618580);
nor I_80563 (I1372117,I1372100,I618592);
not I_80564 (I1372134,I618592);
and I_80565 (I1372151,I1372134,I618586);
nand I_80566 (I1372168,I1372151,I618598);
nor I_80567 (I1372185,I1372134,I1372168);
DFFARX1 I_80568 (I1372185,I2507,I1371987,I1371952,);
not I_80569 (I1372216,I1372168);
nand I_80570 (I1372233,I1372038,I1372216);
nand I_80571 (I1371964,I1372100,I1372216);
DFFARX1 I_80572 (I1372134,I2507,I1371987,I1371979,);
not I_80573 (I1372278,I618604);
nor I_80574 (I1372295,I1372278,I618586);
nor I_80575 (I1372312,I1372295,I1372117);
DFFARX1 I_80576 (I1372312,I2507,I1371987,I1371976,);
not I_80577 (I1372343,I1372295);
DFFARX1 I_80578 (I1372343,I2507,I1371987,I1372369,);
not I_80579 (I1372377,I1372369);
nor I_80580 (I1371973,I1372377,I1372295);
nor I_80581 (I1372408,I1372278,I618583);
and I_80582 (I1372425,I1372408,I618589);
or I_80583 (I1372442,I1372425,I618580);
DFFARX1 I_80584 (I1372442,I2507,I1371987,I1372468,);
not I_80585 (I1372476,I1372468);
nand I_80586 (I1372493,I1372476,I1372216);
not I_80587 (I1371967,I1372493);
nand I_80588 (I1371961,I1372493,I1372233);
nand I_80589 (I1371958,I1372476,I1372100);
not I_80590 (I1372582,I2514);
DFFARX1 I_80591 (I37487,I2507,I1372582,I1372608,);
DFFARX1 I_80592 (I37469,I2507,I1372582,I1372625,);
not I_80593 (I1372633,I1372625);
nor I_80594 (I1372550,I1372608,I1372633);
DFFARX1 I_80595 (I1372633,I2507,I1372582,I1372565,);
nor I_80596 (I1372678,I37469,I37484);
and I_80597 (I1372695,I1372678,I37478);
nor I_80598 (I1372712,I1372695,I37469);
not I_80599 (I1372729,I37469);
and I_80600 (I1372746,I1372729,I37472);
nand I_80601 (I1372763,I1372746,I37475);
nor I_80602 (I1372780,I1372729,I1372763);
DFFARX1 I_80603 (I1372780,I2507,I1372582,I1372547,);
not I_80604 (I1372811,I1372763);
nand I_80605 (I1372828,I1372633,I1372811);
nand I_80606 (I1372559,I1372695,I1372811);
DFFARX1 I_80607 (I1372729,I2507,I1372582,I1372574,);
not I_80608 (I1372873,I37481);
nor I_80609 (I1372890,I1372873,I37472);
nor I_80610 (I1372907,I1372890,I1372712);
DFFARX1 I_80611 (I1372907,I2507,I1372582,I1372571,);
not I_80612 (I1372938,I1372890);
DFFARX1 I_80613 (I1372938,I2507,I1372582,I1372964,);
not I_80614 (I1372972,I1372964);
nor I_80615 (I1372568,I1372972,I1372890);
nor I_80616 (I1373003,I1372873,I37493);
and I_80617 (I1373020,I1373003,I37490);
or I_80618 (I1373037,I1373020,I37472);
DFFARX1 I_80619 (I1373037,I2507,I1372582,I1373063,);
not I_80620 (I1373071,I1373063);
nand I_80621 (I1373088,I1373071,I1372811);
not I_80622 (I1372562,I1373088);
nand I_80623 (I1372556,I1373088,I1372828);
nand I_80624 (I1372553,I1373071,I1372695);
not I_80625 (I1373177,I2514);
DFFARX1 I_80626 (I305019,I2507,I1373177,I1373203,);
DFFARX1 I_80627 (I305013,I2507,I1373177,I1373220,);
not I_80628 (I1373228,I1373220);
nor I_80629 (I1373145,I1373203,I1373228);
DFFARX1 I_80630 (I1373228,I2507,I1373177,I1373160,);
nor I_80631 (I1373273,I305001,I305022);
and I_80632 (I1373290,I1373273,I305016);
nor I_80633 (I1373307,I1373290,I305001);
not I_80634 (I1373324,I305001);
and I_80635 (I1373341,I1373324,I304998);
nand I_80636 (I1373358,I1373341,I305010);
nor I_80637 (I1373375,I1373324,I1373358);
DFFARX1 I_80638 (I1373375,I2507,I1373177,I1373142,);
not I_80639 (I1373406,I1373358);
nand I_80640 (I1373423,I1373228,I1373406);
nand I_80641 (I1373154,I1373290,I1373406);
DFFARX1 I_80642 (I1373324,I2507,I1373177,I1373169,);
not I_80643 (I1373468,I305025);
nor I_80644 (I1373485,I1373468,I304998);
nor I_80645 (I1373502,I1373485,I1373307);
DFFARX1 I_80646 (I1373502,I2507,I1373177,I1373166,);
not I_80647 (I1373533,I1373485);
DFFARX1 I_80648 (I1373533,I2507,I1373177,I1373559,);
not I_80649 (I1373567,I1373559);
nor I_80650 (I1373163,I1373567,I1373485);
nor I_80651 (I1373598,I1373468,I305007);
and I_80652 (I1373615,I1373598,I305004);
or I_80653 (I1373632,I1373615,I304998);
DFFARX1 I_80654 (I1373632,I2507,I1373177,I1373658,);
not I_80655 (I1373666,I1373658);
nand I_80656 (I1373683,I1373666,I1373406);
not I_80657 (I1373157,I1373683);
nand I_80658 (I1373151,I1373683,I1373423);
nand I_80659 (I1373148,I1373666,I1373290);
not I_80660 (I1373772,I2514);
DFFARX1 I_80661 (I918585,I2507,I1373772,I1373798,);
DFFARX1 I_80662 (I918603,I2507,I1373772,I1373815,);
not I_80663 (I1373823,I1373815);
nor I_80664 (I1373740,I1373798,I1373823);
DFFARX1 I_80665 (I1373823,I2507,I1373772,I1373755,);
nor I_80666 (I1373868,I918582,I918594);
and I_80667 (I1373885,I1373868,I918579);
nor I_80668 (I1373902,I1373885,I918582);
not I_80669 (I1373919,I918582);
and I_80670 (I1373936,I1373919,I918588);
nand I_80671 (I1373953,I1373936,I918600);
nor I_80672 (I1373970,I1373919,I1373953);
DFFARX1 I_80673 (I1373970,I2507,I1373772,I1373737,);
not I_80674 (I1374001,I1373953);
nand I_80675 (I1374018,I1373823,I1374001);
nand I_80676 (I1373749,I1373885,I1374001);
DFFARX1 I_80677 (I1373919,I2507,I1373772,I1373764,);
not I_80678 (I1374063,I918591);
nor I_80679 (I1374080,I1374063,I918588);
nor I_80680 (I1374097,I1374080,I1373902);
DFFARX1 I_80681 (I1374097,I2507,I1373772,I1373761,);
not I_80682 (I1374128,I1374080);
DFFARX1 I_80683 (I1374128,I2507,I1373772,I1374154,);
not I_80684 (I1374162,I1374154);
nor I_80685 (I1373758,I1374162,I1374080);
nor I_80686 (I1374193,I1374063,I918579);
and I_80687 (I1374210,I1374193,I918606);
or I_80688 (I1374227,I1374210,I918597);
DFFARX1 I_80689 (I1374227,I2507,I1373772,I1374253,);
not I_80690 (I1374261,I1374253);
nand I_80691 (I1374278,I1374261,I1374001);
not I_80692 (I1373752,I1374278);
nand I_80693 (I1373746,I1374278,I1374018);
nand I_80694 (I1373743,I1374261,I1373885);
not I_80695 (I1374367,I2514);
DFFARX1 I_80696 (I719173,I2507,I1374367,I1374393,);
DFFARX1 I_80697 (I719155,I2507,I1374367,I1374410,);
not I_80698 (I1374418,I1374410);
nor I_80699 (I1374335,I1374393,I1374418);
DFFARX1 I_80700 (I1374418,I2507,I1374367,I1374350,);
nor I_80701 (I1374463,I719161,I719164);
and I_80702 (I1374480,I1374463,I719152);
nor I_80703 (I1374497,I1374480,I719161);
not I_80704 (I1374514,I719161);
and I_80705 (I1374531,I1374514,I719170);
nand I_80706 (I1374548,I1374531,I719158);
nor I_80707 (I1374565,I1374514,I1374548);
DFFARX1 I_80708 (I1374565,I2507,I1374367,I1374332,);
not I_80709 (I1374596,I1374548);
nand I_80710 (I1374613,I1374418,I1374596);
nand I_80711 (I1374344,I1374480,I1374596);
DFFARX1 I_80712 (I1374514,I2507,I1374367,I1374359,);
not I_80713 (I1374658,I719155);
nor I_80714 (I1374675,I1374658,I719170);
nor I_80715 (I1374692,I1374675,I1374497);
DFFARX1 I_80716 (I1374692,I2507,I1374367,I1374356,);
not I_80717 (I1374723,I1374675);
DFFARX1 I_80718 (I1374723,I2507,I1374367,I1374749,);
not I_80719 (I1374757,I1374749);
nor I_80720 (I1374353,I1374757,I1374675);
nor I_80721 (I1374788,I1374658,I719167);
and I_80722 (I1374805,I1374788,I719176);
or I_80723 (I1374822,I1374805,I719152);
DFFARX1 I_80724 (I1374822,I2507,I1374367,I1374848,);
not I_80725 (I1374856,I1374848);
nand I_80726 (I1374873,I1374856,I1374596);
not I_80727 (I1374347,I1374873);
nand I_80728 (I1374341,I1374873,I1374613);
nand I_80729 (I1374338,I1374856,I1374480);
not I_80730 (I1374962,I2514);
DFFARX1 I_80731 (I125499,I2507,I1374962,I1374988,);
DFFARX1 I_80732 (I125487,I2507,I1374962,I1375005,);
not I_80733 (I1375013,I1375005);
nor I_80734 (I1374930,I1374988,I1375013);
DFFARX1 I_80735 (I1375013,I2507,I1374962,I1374945,);
nor I_80736 (I1375058,I125478,I125502);
and I_80737 (I1375075,I1375058,I125481);
nor I_80738 (I1375092,I1375075,I125478);
not I_80739 (I1375109,I125478);
and I_80740 (I1375126,I1375109,I125484);
nand I_80741 (I1375143,I1375126,I125496);
nor I_80742 (I1375160,I1375109,I1375143);
DFFARX1 I_80743 (I1375160,I2507,I1374962,I1374927,);
not I_80744 (I1375191,I1375143);
nand I_80745 (I1375208,I1375013,I1375191);
nand I_80746 (I1374939,I1375075,I1375191);
DFFARX1 I_80747 (I1375109,I2507,I1374962,I1374954,);
not I_80748 (I1375253,I125478);
nor I_80749 (I1375270,I1375253,I125484);
nor I_80750 (I1375287,I1375270,I1375092);
DFFARX1 I_80751 (I1375287,I2507,I1374962,I1374951,);
not I_80752 (I1375318,I1375270);
DFFARX1 I_80753 (I1375318,I2507,I1374962,I1375344,);
not I_80754 (I1375352,I1375344);
nor I_80755 (I1374948,I1375352,I1375270);
nor I_80756 (I1375383,I1375253,I125481);
and I_80757 (I1375400,I1375383,I125490);
or I_80758 (I1375417,I1375400,I125493);
DFFARX1 I_80759 (I1375417,I2507,I1374962,I1375443,);
not I_80760 (I1375451,I1375443);
nand I_80761 (I1375468,I1375451,I1375191);
not I_80762 (I1374942,I1375468);
nand I_80763 (I1374936,I1375468,I1375208);
nand I_80764 (I1374933,I1375451,I1375075);
not I_80765 (I1375557,I2514);
DFFARX1 I_80766 (I906311,I2507,I1375557,I1375583,);
DFFARX1 I_80767 (I906329,I2507,I1375557,I1375600,);
not I_80768 (I1375608,I1375600);
nor I_80769 (I1375525,I1375583,I1375608);
DFFARX1 I_80770 (I1375608,I2507,I1375557,I1375540,);
nor I_80771 (I1375653,I906308,I906320);
and I_80772 (I1375670,I1375653,I906305);
nor I_80773 (I1375687,I1375670,I906308);
not I_80774 (I1375704,I906308);
and I_80775 (I1375721,I1375704,I906314);
nand I_80776 (I1375738,I1375721,I906326);
nor I_80777 (I1375755,I1375704,I1375738);
DFFARX1 I_80778 (I1375755,I2507,I1375557,I1375522,);
not I_80779 (I1375786,I1375738);
nand I_80780 (I1375803,I1375608,I1375786);
nand I_80781 (I1375534,I1375670,I1375786);
DFFARX1 I_80782 (I1375704,I2507,I1375557,I1375549,);
not I_80783 (I1375848,I906317);
nor I_80784 (I1375865,I1375848,I906314);
nor I_80785 (I1375882,I1375865,I1375687);
DFFARX1 I_80786 (I1375882,I2507,I1375557,I1375546,);
not I_80787 (I1375913,I1375865);
DFFARX1 I_80788 (I1375913,I2507,I1375557,I1375939,);
not I_80789 (I1375947,I1375939);
nor I_80790 (I1375543,I1375947,I1375865);
nor I_80791 (I1375978,I1375848,I906305);
and I_80792 (I1375995,I1375978,I906332);
or I_80793 (I1376012,I1375995,I906323);
DFFARX1 I_80794 (I1376012,I2507,I1375557,I1376038,);
not I_80795 (I1376046,I1376038);
nand I_80796 (I1376063,I1376046,I1375786);
not I_80797 (I1375537,I1376063);
nand I_80798 (I1375531,I1376063,I1375803);
nand I_80799 (I1375528,I1376046,I1375670);
not I_80800 (I1376152,I2514);
DFFARX1 I_80801 (I932797,I2507,I1376152,I1376178,);
DFFARX1 I_80802 (I932815,I2507,I1376152,I1376195,);
not I_80803 (I1376203,I1376195);
nor I_80804 (I1376120,I1376178,I1376203);
DFFARX1 I_80805 (I1376203,I2507,I1376152,I1376135,);
nor I_80806 (I1376248,I932794,I932806);
and I_80807 (I1376265,I1376248,I932791);
nor I_80808 (I1376282,I1376265,I932794);
not I_80809 (I1376299,I932794);
and I_80810 (I1376316,I1376299,I932800);
nand I_80811 (I1376333,I1376316,I932812);
nor I_80812 (I1376350,I1376299,I1376333);
DFFARX1 I_80813 (I1376350,I2507,I1376152,I1376117,);
not I_80814 (I1376381,I1376333);
nand I_80815 (I1376398,I1376203,I1376381);
nand I_80816 (I1376129,I1376265,I1376381);
DFFARX1 I_80817 (I1376299,I2507,I1376152,I1376144,);
not I_80818 (I1376443,I932803);
nor I_80819 (I1376460,I1376443,I932800);
nor I_80820 (I1376477,I1376460,I1376282);
DFFARX1 I_80821 (I1376477,I2507,I1376152,I1376141,);
not I_80822 (I1376508,I1376460);
DFFARX1 I_80823 (I1376508,I2507,I1376152,I1376534,);
not I_80824 (I1376542,I1376534);
nor I_80825 (I1376138,I1376542,I1376460);
nor I_80826 (I1376573,I1376443,I932791);
and I_80827 (I1376590,I1376573,I932818);
or I_80828 (I1376607,I1376590,I932809);
DFFARX1 I_80829 (I1376607,I2507,I1376152,I1376633,);
not I_80830 (I1376641,I1376633);
nand I_80831 (I1376658,I1376641,I1376381);
not I_80832 (I1376132,I1376658);
nand I_80833 (I1376126,I1376658,I1376398);
nand I_80834 (I1376123,I1376641,I1376265);
not I_80835 (I1376747,I2514);
DFFARX1 I_80836 (I711659,I2507,I1376747,I1376773,);
DFFARX1 I_80837 (I711641,I2507,I1376747,I1376790,);
not I_80838 (I1376798,I1376790);
nor I_80839 (I1376715,I1376773,I1376798);
DFFARX1 I_80840 (I1376798,I2507,I1376747,I1376730,);
nor I_80841 (I1376843,I711647,I711650);
and I_80842 (I1376860,I1376843,I711638);
nor I_80843 (I1376877,I1376860,I711647);
not I_80844 (I1376894,I711647);
and I_80845 (I1376911,I1376894,I711656);
nand I_80846 (I1376928,I1376911,I711644);
nor I_80847 (I1376945,I1376894,I1376928);
DFFARX1 I_80848 (I1376945,I2507,I1376747,I1376712,);
not I_80849 (I1376976,I1376928);
nand I_80850 (I1376993,I1376798,I1376976);
nand I_80851 (I1376724,I1376860,I1376976);
DFFARX1 I_80852 (I1376894,I2507,I1376747,I1376739,);
not I_80853 (I1377038,I711641);
nor I_80854 (I1377055,I1377038,I711656);
nor I_80855 (I1377072,I1377055,I1376877);
DFFARX1 I_80856 (I1377072,I2507,I1376747,I1376736,);
not I_80857 (I1377103,I1377055);
DFFARX1 I_80858 (I1377103,I2507,I1376747,I1377129,);
not I_80859 (I1377137,I1377129);
nor I_80860 (I1376733,I1377137,I1377055);
nor I_80861 (I1377168,I1377038,I711653);
and I_80862 (I1377185,I1377168,I711662);
or I_80863 (I1377202,I1377185,I711638);
DFFARX1 I_80864 (I1377202,I2507,I1376747,I1377228,);
not I_80865 (I1377236,I1377228);
nand I_80866 (I1377253,I1377236,I1376976);
not I_80867 (I1376727,I1377253);
nand I_80868 (I1376721,I1377253,I1376993);
nand I_80869 (I1376718,I1377236,I1376860);
not I_80870 (I1377342,I2514);
DFFARX1 I_80871 (I1104035,I2507,I1377342,I1377368,);
DFFARX1 I_80872 (I1104047,I2507,I1377342,I1377385,);
not I_80873 (I1377393,I1377385);
nor I_80874 (I1377310,I1377368,I1377393);
DFFARX1 I_80875 (I1377393,I2507,I1377342,I1377325,);
nor I_80876 (I1377438,I1104044,I1104038);
and I_80877 (I1377455,I1377438,I1104032);
nor I_80878 (I1377472,I1377455,I1104044);
not I_80879 (I1377489,I1104044);
and I_80880 (I1377506,I1377489,I1104041);
nand I_80881 (I1377523,I1377506,I1104032);
nor I_80882 (I1377540,I1377489,I1377523);
DFFARX1 I_80883 (I1377540,I2507,I1377342,I1377307,);
not I_80884 (I1377571,I1377523);
nand I_80885 (I1377588,I1377393,I1377571);
nand I_80886 (I1377319,I1377455,I1377571);
DFFARX1 I_80887 (I1377489,I2507,I1377342,I1377334,);
not I_80888 (I1377633,I1104056);
nor I_80889 (I1377650,I1377633,I1104041);
nor I_80890 (I1377667,I1377650,I1377472);
DFFARX1 I_80891 (I1377667,I2507,I1377342,I1377331,);
not I_80892 (I1377698,I1377650);
DFFARX1 I_80893 (I1377698,I2507,I1377342,I1377724,);
not I_80894 (I1377732,I1377724);
nor I_80895 (I1377328,I1377732,I1377650);
nor I_80896 (I1377763,I1377633,I1104050);
and I_80897 (I1377780,I1377763,I1104053);
or I_80898 (I1377797,I1377780,I1104035);
DFFARX1 I_80899 (I1377797,I2507,I1377342,I1377823,);
not I_80900 (I1377831,I1377823);
nand I_80901 (I1377848,I1377831,I1377571);
not I_80902 (I1377322,I1377848);
nand I_80903 (I1377316,I1377848,I1377588);
nand I_80904 (I1377313,I1377831,I1377455);
not I_80905 (I1377937,I2514);
DFFARX1 I_80906 (I132350,I2507,I1377937,I1377963,);
DFFARX1 I_80907 (I132338,I2507,I1377937,I1377980,);
not I_80908 (I1377988,I1377980);
nor I_80909 (I1377905,I1377963,I1377988);
DFFARX1 I_80910 (I1377988,I2507,I1377937,I1377920,);
nor I_80911 (I1378033,I132329,I132353);
and I_80912 (I1378050,I1378033,I132332);
nor I_80913 (I1378067,I1378050,I132329);
not I_80914 (I1378084,I132329);
and I_80915 (I1378101,I1378084,I132335);
nand I_80916 (I1378118,I1378101,I132347);
nor I_80917 (I1378135,I1378084,I1378118);
DFFARX1 I_80918 (I1378135,I2507,I1377937,I1377902,);
not I_80919 (I1378166,I1378118);
nand I_80920 (I1378183,I1377988,I1378166);
nand I_80921 (I1377914,I1378050,I1378166);
DFFARX1 I_80922 (I1378084,I2507,I1377937,I1377929,);
not I_80923 (I1378228,I132329);
nor I_80924 (I1378245,I1378228,I132335);
nor I_80925 (I1378262,I1378245,I1378067);
DFFARX1 I_80926 (I1378262,I2507,I1377937,I1377926,);
not I_80927 (I1378293,I1378245);
DFFARX1 I_80928 (I1378293,I2507,I1377937,I1378319,);
not I_80929 (I1378327,I1378319);
nor I_80930 (I1377923,I1378327,I1378245);
nor I_80931 (I1378358,I1378228,I132332);
and I_80932 (I1378375,I1378358,I132341);
or I_80933 (I1378392,I1378375,I132344);
DFFARX1 I_80934 (I1378392,I2507,I1377937,I1378418,);
not I_80935 (I1378426,I1378418);
nand I_80936 (I1378443,I1378426,I1378166);
not I_80937 (I1377917,I1378443);
nand I_80938 (I1377911,I1378443,I1378183);
nand I_80939 (I1377908,I1378426,I1378050);
not I_80940 (I1378532,I2514);
DFFARX1 I_80941 (I123918,I2507,I1378532,I1378558,);
DFFARX1 I_80942 (I123906,I2507,I1378532,I1378575,);
not I_80943 (I1378583,I1378575);
nor I_80944 (I1378500,I1378558,I1378583);
DFFARX1 I_80945 (I1378583,I2507,I1378532,I1378515,);
nor I_80946 (I1378628,I123897,I123921);
and I_80947 (I1378645,I1378628,I123900);
nor I_80948 (I1378662,I1378645,I123897);
not I_80949 (I1378679,I123897);
and I_80950 (I1378696,I1378679,I123903);
nand I_80951 (I1378713,I1378696,I123915);
nor I_80952 (I1378730,I1378679,I1378713);
DFFARX1 I_80953 (I1378730,I2507,I1378532,I1378497,);
not I_80954 (I1378761,I1378713);
nand I_80955 (I1378778,I1378583,I1378761);
nand I_80956 (I1378509,I1378645,I1378761);
DFFARX1 I_80957 (I1378679,I2507,I1378532,I1378524,);
not I_80958 (I1378823,I123897);
nor I_80959 (I1378840,I1378823,I123903);
nor I_80960 (I1378857,I1378840,I1378662);
DFFARX1 I_80961 (I1378857,I2507,I1378532,I1378521,);
not I_80962 (I1378888,I1378840);
DFFARX1 I_80963 (I1378888,I2507,I1378532,I1378914,);
not I_80964 (I1378922,I1378914);
nor I_80965 (I1378518,I1378922,I1378840);
nor I_80966 (I1378953,I1378823,I123900);
and I_80967 (I1378970,I1378953,I123909);
or I_80968 (I1378987,I1378970,I123912);
DFFARX1 I_80969 (I1378987,I2507,I1378532,I1379013,);
not I_80970 (I1379021,I1379013);
nand I_80971 (I1379038,I1379021,I1378761);
not I_80972 (I1378512,I1379038);
nand I_80973 (I1378506,I1379038,I1378778);
nand I_80974 (I1378503,I1379021,I1378645);
not I_80975 (I1379127,I2514);
DFFARX1 I_80976 (I59624,I2507,I1379127,I1379153,);
DFFARX1 I_80977 (I59612,I2507,I1379127,I1379170,);
not I_80978 (I1379178,I1379170);
nor I_80979 (I1379095,I1379153,I1379178);
DFFARX1 I_80980 (I1379178,I2507,I1379127,I1379110,);
nor I_80981 (I1379223,I59603,I59627);
and I_80982 (I1379240,I1379223,I59606);
nor I_80983 (I1379257,I1379240,I59603);
not I_80984 (I1379274,I59603);
and I_80985 (I1379291,I1379274,I59609);
nand I_80986 (I1379308,I1379291,I59621);
nor I_80987 (I1379325,I1379274,I1379308);
DFFARX1 I_80988 (I1379325,I2507,I1379127,I1379092,);
not I_80989 (I1379356,I1379308);
nand I_80990 (I1379373,I1379178,I1379356);
nand I_80991 (I1379104,I1379240,I1379356);
DFFARX1 I_80992 (I1379274,I2507,I1379127,I1379119,);
not I_80993 (I1379418,I59603);
nor I_80994 (I1379435,I1379418,I59609);
nor I_80995 (I1379452,I1379435,I1379257);
DFFARX1 I_80996 (I1379452,I2507,I1379127,I1379116,);
not I_80997 (I1379483,I1379435);
DFFARX1 I_80998 (I1379483,I2507,I1379127,I1379509,);
not I_80999 (I1379517,I1379509);
nor I_81000 (I1379113,I1379517,I1379435);
nor I_81001 (I1379548,I1379418,I59606);
and I_81002 (I1379565,I1379548,I59615);
or I_81003 (I1379582,I1379565,I59618);
DFFARX1 I_81004 (I1379582,I2507,I1379127,I1379608,);
not I_81005 (I1379616,I1379608);
nand I_81006 (I1379633,I1379616,I1379356);
not I_81007 (I1379107,I1379633);
nand I_81008 (I1379101,I1379633,I1379373);
nand I_81009 (I1379098,I1379616,I1379240);
not I_81010 (I1379722,I2514);
DFFARX1 I_81011 (I166890,I2507,I1379722,I1379748,);
DFFARX1 I_81012 (I166893,I2507,I1379722,I1379765,);
not I_81013 (I1379773,I1379765);
nor I_81014 (I1379690,I1379748,I1379773);
DFFARX1 I_81015 (I1379773,I2507,I1379722,I1379705,);
nor I_81016 (I1379818,I166899,I166893);
and I_81017 (I1379835,I1379818,I166896);
nor I_81018 (I1379852,I1379835,I166899);
not I_81019 (I1379869,I166899);
and I_81020 (I1379886,I1379869,I166890);
nand I_81021 (I1379903,I1379886,I166908);
nor I_81022 (I1379920,I1379869,I1379903);
DFFARX1 I_81023 (I1379920,I2507,I1379722,I1379687,);
not I_81024 (I1379951,I1379903);
nand I_81025 (I1379968,I1379773,I1379951);
nand I_81026 (I1379699,I1379835,I1379951);
DFFARX1 I_81027 (I1379869,I2507,I1379722,I1379714,);
not I_81028 (I1380013,I166902);
nor I_81029 (I1380030,I1380013,I166890);
nor I_81030 (I1380047,I1380030,I1379852);
DFFARX1 I_81031 (I1380047,I2507,I1379722,I1379711,);
not I_81032 (I1380078,I1380030);
DFFARX1 I_81033 (I1380078,I2507,I1379722,I1380104,);
not I_81034 (I1380112,I1380104);
nor I_81035 (I1379708,I1380112,I1380030);
nor I_81036 (I1380143,I1380013,I166905);
and I_81037 (I1380160,I1380143,I166911);
or I_81038 (I1380177,I1380160,I166914);
DFFARX1 I_81039 (I1380177,I2507,I1379722,I1380203,);
not I_81040 (I1380211,I1380203);
nand I_81041 (I1380228,I1380211,I1379951);
not I_81042 (I1379702,I1380228);
nand I_81043 (I1379696,I1380228,I1379968);
nand I_81044 (I1379693,I1380211,I1379835);
not I_81045 (I1380317,I2514);
DFFARX1 I_81046 (I761945,I2507,I1380317,I1380343,);
DFFARX1 I_81047 (I761927,I2507,I1380317,I1380360,);
not I_81048 (I1380368,I1380360);
nor I_81049 (I1380285,I1380343,I1380368);
DFFARX1 I_81050 (I1380368,I2507,I1380317,I1380300,);
nor I_81051 (I1380413,I761933,I761936);
and I_81052 (I1380430,I1380413,I761924);
nor I_81053 (I1380447,I1380430,I761933);
not I_81054 (I1380464,I761933);
and I_81055 (I1380481,I1380464,I761942);
nand I_81056 (I1380498,I1380481,I761930);
nor I_81057 (I1380515,I1380464,I1380498);
DFFARX1 I_81058 (I1380515,I2507,I1380317,I1380282,);
not I_81059 (I1380546,I1380498);
nand I_81060 (I1380563,I1380368,I1380546);
nand I_81061 (I1380294,I1380430,I1380546);
DFFARX1 I_81062 (I1380464,I2507,I1380317,I1380309,);
not I_81063 (I1380608,I761927);
nor I_81064 (I1380625,I1380608,I761942);
nor I_81065 (I1380642,I1380625,I1380447);
DFFARX1 I_81066 (I1380642,I2507,I1380317,I1380306,);
not I_81067 (I1380673,I1380625);
DFFARX1 I_81068 (I1380673,I2507,I1380317,I1380699,);
not I_81069 (I1380707,I1380699);
nor I_81070 (I1380303,I1380707,I1380625);
nor I_81071 (I1380738,I1380608,I761939);
and I_81072 (I1380755,I1380738,I761948);
or I_81073 (I1380772,I1380755,I761924);
DFFARX1 I_81074 (I1380772,I2507,I1380317,I1380798,);
not I_81075 (I1380806,I1380798);
nand I_81076 (I1380823,I1380806,I1380546);
not I_81077 (I1380297,I1380823);
nand I_81078 (I1380291,I1380823,I1380563);
nand I_81079 (I1380288,I1380806,I1380430);
not I_81080 (I1380912,I2514);
DFFARX1 I_81081 (I825445,I2507,I1380912,I1380938,);
DFFARX1 I_81082 (I825442,I2507,I1380912,I1380955,);
not I_81083 (I1380963,I1380955);
nor I_81084 (I1380880,I1380938,I1380963);
DFFARX1 I_81085 (I1380963,I2507,I1380912,I1380895,);
nor I_81086 (I1381008,I825457,I825439);
and I_81087 (I1381025,I1381008,I825436);
nor I_81088 (I1381042,I1381025,I825457);
not I_81089 (I1381059,I825457);
and I_81090 (I1381076,I1381059,I825442);
nand I_81091 (I1381093,I1381076,I825454);
nor I_81092 (I1381110,I1381059,I1381093);
DFFARX1 I_81093 (I1381110,I2507,I1380912,I1380877,);
not I_81094 (I1381141,I1381093);
nand I_81095 (I1381158,I1380963,I1381141);
nand I_81096 (I1380889,I1381025,I1381141);
DFFARX1 I_81097 (I1381059,I2507,I1380912,I1380904,);
not I_81098 (I1381203,I825448);
nor I_81099 (I1381220,I1381203,I825442);
nor I_81100 (I1381237,I1381220,I1381042);
DFFARX1 I_81101 (I1381237,I2507,I1380912,I1380901,);
not I_81102 (I1381268,I1381220);
DFFARX1 I_81103 (I1381268,I2507,I1380912,I1381294,);
not I_81104 (I1381302,I1381294);
nor I_81105 (I1380898,I1381302,I1381220);
nor I_81106 (I1381333,I1381203,I825436);
and I_81107 (I1381350,I1381333,I825451);
or I_81108 (I1381367,I1381350,I825439);
DFFARX1 I_81109 (I1381367,I2507,I1380912,I1381393,);
not I_81110 (I1381401,I1381393);
nand I_81111 (I1381418,I1381401,I1381141);
not I_81112 (I1380892,I1381418);
nand I_81113 (I1380886,I1381418,I1381158);
nand I_81114 (I1380883,I1381401,I1381025);
not I_81115 (I1381507,I2514);
DFFARX1 I_81116 (I1005149,I2507,I1381507,I1381533,);
DFFARX1 I_81117 (I1005167,I2507,I1381507,I1381550,);
not I_81118 (I1381558,I1381550);
nor I_81119 (I1381475,I1381533,I1381558);
DFFARX1 I_81120 (I1381558,I2507,I1381507,I1381490,);
nor I_81121 (I1381603,I1005146,I1005158);
and I_81122 (I1381620,I1381603,I1005143);
nor I_81123 (I1381637,I1381620,I1005146);
not I_81124 (I1381654,I1005146);
and I_81125 (I1381671,I1381654,I1005152);
nand I_81126 (I1381688,I1381671,I1005164);
nor I_81127 (I1381705,I1381654,I1381688);
DFFARX1 I_81128 (I1381705,I2507,I1381507,I1381472,);
not I_81129 (I1381736,I1381688);
nand I_81130 (I1381753,I1381558,I1381736);
nand I_81131 (I1381484,I1381620,I1381736);
DFFARX1 I_81132 (I1381654,I2507,I1381507,I1381499,);
not I_81133 (I1381798,I1005155);
nor I_81134 (I1381815,I1381798,I1005152);
nor I_81135 (I1381832,I1381815,I1381637);
DFFARX1 I_81136 (I1381832,I2507,I1381507,I1381496,);
not I_81137 (I1381863,I1381815);
DFFARX1 I_81138 (I1381863,I2507,I1381507,I1381889,);
not I_81139 (I1381897,I1381889);
nor I_81140 (I1381493,I1381897,I1381815);
nor I_81141 (I1381928,I1381798,I1005143);
and I_81142 (I1381945,I1381928,I1005170);
or I_81143 (I1381962,I1381945,I1005161);
DFFARX1 I_81144 (I1381962,I2507,I1381507,I1381988,);
not I_81145 (I1381996,I1381988);
nand I_81146 (I1382013,I1381996,I1381736);
not I_81147 (I1381487,I1382013);
nand I_81148 (I1381481,I1382013,I1381753);
nand I_81149 (I1381478,I1381996,I1381620);
not I_81150 (I1382102,I2514);
DFFARX1 I_81151 (I1022495,I2507,I1382102,I1382128,);
DFFARX1 I_81152 (I1022486,I2507,I1382102,I1382145,);
not I_81153 (I1382153,I1382145);
nor I_81154 (I1382070,I1382128,I1382153);
DFFARX1 I_81155 (I1382153,I2507,I1382102,I1382085,);
nor I_81156 (I1382198,I1022492,I1022501);
and I_81157 (I1382215,I1382198,I1022504);
nor I_81158 (I1382232,I1382215,I1022492);
not I_81159 (I1382249,I1022492);
and I_81160 (I1382266,I1382249,I1022483);
nand I_81161 (I1382283,I1382266,I1022489);
nor I_81162 (I1382300,I1382249,I1382283);
DFFARX1 I_81163 (I1382300,I2507,I1382102,I1382067,);
not I_81164 (I1382331,I1382283);
nand I_81165 (I1382348,I1382153,I1382331);
nand I_81166 (I1382079,I1382215,I1382331);
DFFARX1 I_81167 (I1382249,I2507,I1382102,I1382094,);
not I_81168 (I1382393,I1022498);
nor I_81169 (I1382410,I1382393,I1022483);
nor I_81170 (I1382427,I1382410,I1382232);
DFFARX1 I_81171 (I1382427,I2507,I1382102,I1382091,);
not I_81172 (I1382458,I1382410);
DFFARX1 I_81173 (I1382458,I2507,I1382102,I1382484,);
not I_81174 (I1382492,I1382484);
nor I_81175 (I1382088,I1382492,I1382410);
nor I_81176 (I1382523,I1382393,I1022483);
and I_81177 (I1382540,I1382523,I1022486);
or I_81178 (I1382557,I1382540,I1022489);
DFFARX1 I_81179 (I1382557,I2507,I1382102,I1382583,);
not I_81180 (I1382591,I1382583);
nand I_81181 (I1382608,I1382591,I1382331);
not I_81182 (I1382082,I1382608);
nand I_81183 (I1382076,I1382608,I1382348);
nand I_81184 (I1382073,I1382591,I1382215);
not I_81185 (I1382697,I2514);
DFFARX1 I_81186 (I49084,I2507,I1382697,I1382723,);
DFFARX1 I_81187 (I49072,I2507,I1382697,I1382740,);
not I_81188 (I1382748,I1382740);
nor I_81189 (I1382665,I1382723,I1382748);
DFFARX1 I_81190 (I1382748,I2507,I1382697,I1382680,);
nor I_81191 (I1382793,I49063,I49087);
and I_81192 (I1382810,I1382793,I49066);
nor I_81193 (I1382827,I1382810,I49063);
not I_81194 (I1382844,I49063);
and I_81195 (I1382861,I1382844,I49069);
nand I_81196 (I1382878,I1382861,I49081);
nor I_81197 (I1382895,I1382844,I1382878);
DFFARX1 I_81198 (I1382895,I2507,I1382697,I1382662,);
not I_81199 (I1382926,I1382878);
nand I_81200 (I1382943,I1382748,I1382926);
nand I_81201 (I1382674,I1382810,I1382926);
DFFARX1 I_81202 (I1382844,I2507,I1382697,I1382689,);
not I_81203 (I1382988,I49063);
nor I_81204 (I1383005,I1382988,I49069);
nor I_81205 (I1383022,I1383005,I1382827);
DFFARX1 I_81206 (I1383022,I2507,I1382697,I1382686,);
not I_81207 (I1383053,I1383005);
DFFARX1 I_81208 (I1383053,I2507,I1382697,I1383079,);
not I_81209 (I1383087,I1383079);
nor I_81210 (I1382683,I1383087,I1383005);
nor I_81211 (I1383118,I1382988,I49066);
and I_81212 (I1383135,I1383118,I49075);
or I_81213 (I1383152,I1383135,I49078);
DFFARX1 I_81214 (I1383152,I2507,I1382697,I1383178,);
not I_81215 (I1383186,I1383178);
nand I_81216 (I1383203,I1383186,I1382926);
not I_81217 (I1382677,I1383203);
nand I_81218 (I1382671,I1383203,I1382943);
nand I_81219 (I1382668,I1383186,I1382810);
not I_81220 (I1383292,I2514);
DFFARX1 I_81221 (I539904,I2507,I1383292,I1383318,);
DFFARX1 I_81222 (I539907,I2507,I1383292,I1383335,);
not I_81223 (I1383343,I1383335);
nor I_81224 (I1383260,I1383318,I1383343);
DFFARX1 I_81225 (I1383343,I2507,I1383292,I1383275,);
nor I_81226 (I1383388,I539910,I539928);
and I_81227 (I1383405,I1383388,I539913);
nor I_81228 (I1383422,I1383405,I539910);
not I_81229 (I1383439,I539910);
and I_81230 (I1383456,I1383439,I539922);
nand I_81231 (I1383473,I1383456,I539925);
nor I_81232 (I1383490,I1383439,I1383473);
DFFARX1 I_81233 (I1383490,I2507,I1383292,I1383257,);
not I_81234 (I1383521,I1383473);
nand I_81235 (I1383538,I1383343,I1383521);
nand I_81236 (I1383269,I1383405,I1383521);
DFFARX1 I_81237 (I1383439,I2507,I1383292,I1383284,);
not I_81238 (I1383583,I539916);
nor I_81239 (I1383600,I1383583,I539922);
nor I_81240 (I1383617,I1383600,I1383422);
DFFARX1 I_81241 (I1383617,I2507,I1383292,I1383281,);
not I_81242 (I1383648,I1383600);
DFFARX1 I_81243 (I1383648,I2507,I1383292,I1383674,);
not I_81244 (I1383682,I1383674);
nor I_81245 (I1383278,I1383682,I1383600);
nor I_81246 (I1383713,I1383583,I539904);
and I_81247 (I1383730,I1383713,I539919);
or I_81248 (I1383747,I1383730,I539907);
DFFARX1 I_81249 (I1383747,I2507,I1383292,I1383773,);
not I_81250 (I1383781,I1383773);
nand I_81251 (I1383798,I1383781,I1383521);
not I_81252 (I1383272,I1383798);
nand I_81253 (I1383266,I1383798,I1383538);
nand I_81254 (I1383263,I1383781,I1383405);
not I_81255 (I1383887,I2514);
DFFARX1 I_81256 (I48027,I2507,I1383887,I1383913,);
DFFARX1 I_81257 (I48009,I2507,I1383887,I1383930,);
not I_81258 (I1383938,I1383930);
nor I_81259 (I1383855,I1383913,I1383938);
DFFARX1 I_81260 (I1383938,I2507,I1383887,I1383870,);
nor I_81261 (I1383983,I48009,I48024);
and I_81262 (I1384000,I1383983,I48018);
nor I_81263 (I1384017,I1384000,I48009);
not I_81264 (I1384034,I48009);
and I_81265 (I1384051,I1384034,I48012);
nand I_81266 (I1384068,I1384051,I48015);
nor I_81267 (I1384085,I1384034,I1384068);
DFFARX1 I_81268 (I1384085,I2507,I1383887,I1383852,);
not I_81269 (I1384116,I1384068);
nand I_81270 (I1384133,I1383938,I1384116);
nand I_81271 (I1383864,I1384000,I1384116);
DFFARX1 I_81272 (I1384034,I2507,I1383887,I1383879,);
not I_81273 (I1384178,I48021);
nor I_81274 (I1384195,I1384178,I48012);
nor I_81275 (I1384212,I1384195,I1384017);
DFFARX1 I_81276 (I1384212,I2507,I1383887,I1383876,);
not I_81277 (I1384243,I1384195);
DFFARX1 I_81278 (I1384243,I2507,I1383887,I1384269,);
not I_81279 (I1384277,I1384269);
nor I_81280 (I1383873,I1384277,I1384195);
nor I_81281 (I1384308,I1384178,I48033);
and I_81282 (I1384325,I1384308,I48030);
or I_81283 (I1384342,I1384325,I48012);
DFFARX1 I_81284 (I1384342,I2507,I1383887,I1384368,);
not I_81285 (I1384376,I1384368);
nand I_81286 (I1384393,I1384376,I1384116);
not I_81287 (I1383867,I1384393);
nand I_81288 (I1383861,I1384393,I1384133);
nand I_81289 (I1383858,I1384376,I1384000);
not I_81290 (I1384482,I2514);
DFFARX1 I_81291 (I391919,I2507,I1384482,I1384508,);
DFFARX1 I_81292 (I391925,I2507,I1384482,I1384525,);
not I_81293 (I1384533,I1384525);
nor I_81294 (I1384450,I1384508,I1384533);
DFFARX1 I_81295 (I1384533,I2507,I1384482,I1384465,);
nor I_81296 (I1384578,I391934,I391919);
and I_81297 (I1384595,I1384578,I391946);
nor I_81298 (I1384612,I1384595,I391934);
not I_81299 (I1384629,I391934);
and I_81300 (I1384646,I1384629,I391922);
nand I_81301 (I1384663,I1384646,I391943);
nor I_81302 (I1384680,I1384629,I1384663);
DFFARX1 I_81303 (I1384680,I2507,I1384482,I1384447,);
not I_81304 (I1384711,I1384663);
nand I_81305 (I1384728,I1384533,I1384711);
nand I_81306 (I1384459,I1384595,I1384711);
DFFARX1 I_81307 (I1384629,I2507,I1384482,I1384474,);
not I_81308 (I1384773,I391931);
nor I_81309 (I1384790,I1384773,I391922);
nor I_81310 (I1384807,I1384790,I1384612);
DFFARX1 I_81311 (I1384807,I2507,I1384482,I1384471,);
not I_81312 (I1384838,I1384790);
DFFARX1 I_81313 (I1384838,I2507,I1384482,I1384864,);
not I_81314 (I1384872,I1384864);
nor I_81315 (I1384468,I1384872,I1384790);
nor I_81316 (I1384903,I1384773,I391928);
and I_81317 (I1384920,I1384903,I391940);
or I_81318 (I1384937,I1384920,I391937);
DFFARX1 I_81319 (I1384937,I2507,I1384482,I1384963,);
not I_81320 (I1384971,I1384963);
nand I_81321 (I1384988,I1384971,I1384711);
not I_81322 (I1384462,I1384988);
nand I_81323 (I1384456,I1384988,I1384728);
nand I_81324 (I1384453,I1384971,I1384595);
not I_81325 (I1385077,I2514);
DFFARX1 I_81326 (I165105,I2507,I1385077,I1385103,);
DFFARX1 I_81327 (I165108,I2507,I1385077,I1385120,);
not I_81328 (I1385128,I1385120);
nor I_81329 (I1385045,I1385103,I1385128);
DFFARX1 I_81330 (I1385128,I2507,I1385077,I1385060,);
nor I_81331 (I1385173,I165114,I165108);
and I_81332 (I1385190,I1385173,I165111);
nor I_81333 (I1385207,I1385190,I165114);
not I_81334 (I1385224,I165114);
and I_81335 (I1385241,I1385224,I165105);
nand I_81336 (I1385258,I1385241,I165123);
nor I_81337 (I1385275,I1385224,I1385258);
DFFARX1 I_81338 (I1385275,I2507,I1385077,I1385042,);
not I_81339 (I1385306,I1385258);
nand I_81340 (I1385323,I1385128,I1385306);
nand I_81341 (I1385054,I1385190,I1385306);
DFFARX1 I_81342 (I1385224,I2507,I1385077,I1385069,);
not I_81343 (I1385368,I165117);
nor I_81344 (I1385385,I1385368,I165105);
nor I_81345 (I1385402,I1385385,I1385207);
DFFARX1 I_81346 (I1385402,I2507,I1385077,I1385066,);
not I_81347 (I1385433,I1385385);
DFFARX1 I_81348 (I1385433,I2507,I1385077,I1385459,);
not I_81349 (I1385467,I1385459);
nor I_81350 (I1385063,I1385467,I1385385);
nor I_81351 (I1385498,I1385368,I165120);
and I_81352 (I1385515,I1385498,I165126);
or I_81353 (I1385532,I1385515,I165129);
DFFARX1 I_81354 (I1385532,I2507,I1385077,I1385558,);
not I_81355 (I1385566,I1385558);
nand I_81356 (I1385583,I1385566,I1385306);
not I_81357 (I1385057,I1385583);
nand I_81358 (I1385051,I1385583,I1385323);
nand I_81359 (I1385048,I1385566,I1385190);
not I_81360 (I1385672,I2514);
DFFARX1 I_81361 (I662529,I2507,I1385672,I1385698,);
DFFARX1 I_81362 (I662511,I2507,I1385672,I1385715,);
not I_81363 (I1385723,I1385715);
nor I_81364 (I1385640,I1385698,I1385723);
DFFARX1 I_81365 (I1385723,I2507,I1385672,I1385655,);
nor I_81366 (I1385768,I662517,I662520);
and I_81367 (I1385785,I1385768,I662508);
nor I_81368 (I1385802,I1385785,I662517);
not I_81369 (I1385819,I662517);
and I_81370 (I1385836,I1385819,I662526);
nand I_81371 (I1385853,I1385836,I662514);
nor I_81372 (I1385870,I1385819,I1385853);
DFFARX1 I_81373 (I1385870,I2507,I1385672,I1385637,);
not I_81374 (I1385901,I1385853);
nand I_81375 (I1385918,I1385723,I1385901);
nand I_81376 (I1385649,I1385785,I1385901);
DFFARX1 I_81377 (I1385819,I2507,I1385672,I1385664,);
not I_81378 (I1385963,I662511);
nor I_81379 (I1385980,I1385963,I662526);
nor I_81380 (I1385997,I1385980,I1385802);
DFFARX1 I_81381 (I1385997,I2507,I1385672,I1385661,);
not I_81382 (I1386028,I1385980);
DFFARX1 I_81383 (I1386028,I2507,I1385672,I1386054,);
not I_81384 (I1386062,I1386054);
nor I_81385 (I1385658,I1386062,I1385980);
nor I_81386 (I1386093,I1385963,I662523);
and I_81387 (I1386110,I1386093,I662532);
or I_81388 (I1386127,I1386110,I662508);
DFFARX1 I_81389 (I1386127,I2507,I1385672,I1386153,);
not I_81390 (I1386161,I1386153);
nand I_81391 (I1386178,I1386161,I1385901);
not I_81392 (I1385652,I1386178);
nand I_81393 (I1385646,I1386178,I1385918);
nand I_81394 (I1385643,I1386161,I1385785);
not I_81395 (I1386267,I2514);
DFFARX1 I_81396 (I861281,I2507,I1386267,I1386293,);
DFFARX1 I_81397 (I861278,I2507,I1386267,I1386310,);
not I_81398 (I1386318,I1386310);
nor I_81399 (I1386235,I1386293,I1386318);
DFFARX1 I_81400 (I1386318,I2507,I1386267,I1386250,);
nor I_81401 (I1386363,I861293,I861275);
and I_81402 (I1386380,I1386363,I861272);
nor I_81403 (I1386397,I1386380,I861293);
not I_81404 (I1386414,I861293);
and I_81405 (I1386431,I1386414,I861278);
nand I_81406 (I1386448,I1386431,I861290);
nor I_81407 (I1386465,I1386414,I1386448);
DFFARX1 I_81408 (I1386465,I2507,I1386267,I1386232,);
not I_81409 (I1386496,I1386448);
nand I_81410 (I1386513,I1386318,I1386496);
nand I_81411 (I1386244,I1386380,I1386496);
DFFARX1 I_81412 (I1386414,I2507,I1386267,I1386259,);
not I_81413 (I1386558,I861284);
nor I_81414 (I1386575,I1386558,I861278);
nor I_81415 (I1386592,I1386575,I1386397);
DFFARX1 I_81416 (I1386592,I2507,I1386267,I1386256,);
not I_81417 (I1386623,I1386575);
DFFARX1 I_81418 (I1386623,I2507,I1386267,I1386649,);
not I_81419 (I1386657,I1386649);
nor I_81420 (I1386253,I1386657,I1386575);
nor I_81421 (I1386688,I1386558,I861272);
and I_81422 (I1386705,I1386688,I861287);
or I_81423 (I1386722,I1386705,I861275);
DFFARX1 I_81424 (I1386722,I2507,I1386267,I1386748,);
not I_81425 (I1386756,I1386748);
nand I_81426 (I1386773,I1386756,I1386496);
not I_81427 (I1386247,I1386773);
nand I_81428 (I1386241,I1386773,I1386513);
nand I_81429 (I1386238,I1386756,I1386380);
not I_81430 (I1386862,I2514);
DFFARX1 I_81431 (I1191313,I2507,I1386862,I1386888,);
DFFARX1 I_81432 (I1191325,I2507,I1386862,I1386905,);
not I_81433 (I1386913,I1386905);
nor I_81434 (I1386830,I1386888,I1386913);
DFFARX1 I_81435 (I1386913,I2507,I1386862,I1386845,);
nor I_81436 (I1386958,I1191322,I1191316);
and I_81437 (I1386975,I1386958,I1191310);
nor I_81438 (I1386992,I1386975,I1191322);
not I_81439 (I1387009,I1191322);
and I_81440 (I1387026,I1387009,I1191319);
nand I_81441 (I1387043,I1387026,I1191310);
nor I_81442 (I1387060,I1387009,I1387043);
DFFARX1 I_81443 (I1387060,I2507,I1386862,I1386827,);
not I_81444 (I1387091,I1387043);
nand I_81445 (I1387108,I1386913,I1387091);
nand I_81446 (I1386839,I1386975,I1387091);
DFFARX1 I_81447 (I1387009,I2507,I1386862,I1386854,);
not I_81448 (I1387153,I1191334);
nor I_81449 (I1387170,I1387153,I1191319);
nor I_81450 (I1387187,I1387170,I1386992);
DFFARX1 I_81451 (I1387187,I2507,I1386862,I1386851,);
not I_81452 (I1387218,I1387170);
DFFARX1 I_81453 (I1387218,I2507,I1386862,I1387244,);
not I_81454 (I1387252,I1387244);
nor I_81455 (I1386848,I1387252,I1387170);
nor I_81456 (I1387283,I1387153,I1191328);
and I_81457 (I1387300,I1387283,I1191331);
or I_81458 (I1387317,I1387300,I1191313);
DFFARX1 I_81459 (I1387317,I2507,I1386862,I1387343,);
not I_81460 (I1387351,I1387343);
nand I_81461 (I1387368,I1387351,I1387091);
not I_81462 (I1386842,I1387368);
nand I_81463 (I1386836,I1387368,I1387108);
nand I_81464 (I1386833,I1387351,I1386975);
not I_81465 (I1387457,I2514);
DFFARX1 I_81466 (I971557,I2507,I1387457,I1387483,);
DFFARX1 I_81467 (I971575,I2507,I1387457,I1387500,);
not I_81468 (I1387508,I1387500);
nor I_81469 (I1387425,I1387483,I1387508);
DFFARX1 I_81470 (I1387508,I2507,I1387457,I1387440,);
nor I_81471 (I1387553,I971554,I971566);
and I_81472 (I1387570,I1387553,I971551);
nor I_81473 (I1387587,I1387570,I971554);
not I_81474 (I1387604,I971554);
and I_81475 (I1387621,I1387604,I971560);
nand I_81476 (I1387638,I1387621,I971572);
nor I_81477 (I1387655,I1387604,I1387638);
DFFARX1 I_81478 (I1387655,I2507,I1387457,I1387422,);
not I_81479 (I1387686,I1387638);
nand I_81480 (I1387703,I1387508,I1387686);
nand I_81481 (I1387434,I1387570,I1387686);
DFFARX1 I_81482 (I1387604,I2507,I1387457,I1387449,);
not I_81483 (I1387748,I971563);
nor I_81484 (I1387765,I1387748,I971560);
nor I_81485 (I1387782,I1387765,I1387587);
DFFARX1 I_81486 (I1387782,I2507,I1387457,I1387446,);
not I_81487 (I1387813,I1387765);
DFFARX1 I_81488 (I1387813,I2507,I1387457,I1387839,);
not I_81489 (I1387847,I1387839);
nor I_81490 (I1387443,I1387847,I1387765);
nor I_81491 (I1387878,I1387748,I971551);
and I_81492 (I1387895,I1387878,I971578);
or I_81493 (I1387912,I1387895,I971569);
DFFARX1 I_81494 (I1387912,I2507,I1387457,I1387938,);
not I_81495 (I1387946,I1387938);
nand I_81496 (I1387963,I1387946,I1387686);
not I_81497 (I1387437,I1387963);
nand I_81498 (I1387431,I1387963,I1387703);
nand I_81499 (I1387428,I1387946,I1387570);
not I_81500 (I1388052,I2514);
DFFARX1 I_81501 (I1293498,I2507,I1388052,I1388078,);
DFFARX1 I_81502 (I1293489,I2507,I1388052,I1388095,);
not I_81503 (I1388103,I1388095);
nor I_81504 (I1388020,I1388078,I1388103);
DFFARX1 I_81505 (I1388103,I2507,I1388052,I1388035,);
nor I_81506 (I1388148,I1293480,I1293495);
and I_81507 (I1388165,I1388148,I1293483);
nor I_81508 (I1388182,I1388165,I1293480);
not I_81509 (I1388199,I1293480);
and I_81510 (I1388216,I1388199,I1293486);
nand I_81511 (I1388233,I1388216,I1293504);
nor I_81512 (I1388250,I1388199,I1388233);
DFFARX1 I_81513 (I1388250,I2507,I1388052,I1388017,);
not I_81514 (I1388281,I1388233);
nand I_81515 (I1388298,I1388103,I1388281);
nand I_81516 (I1388029,I1388165,I1388281);
DFFARX1 I_81517 (I1388199,I2507,I1388052,I1388044,);
not I_81518 (I1388343,I1293480);
nor I_81519 (I1388360,I1388343,I1293486);
nor I_81520 (I1388377,I1388360,I1388182);
DFFARX1 I_81521 (I1388377,I2507,I1388052,I1388041,);
not I_81522 (I1388408,I1388360);
DFFARX1 I_81523 (I1388408,I2507,I1388052,I1388434,);
not I_81524 (I1388442,I1388434);
nor I_81525 (I1388038,I1388442,I1388360);
nor I_81526 (I1388473,I1388343,I1293483);
and I_81527 (I1388490,I1388473,I1293492);
or I_81528 (I1388507,I1388490,I1293501);
DFFARX1 I_81529 (I1388507,I2507,I1388052,I1388533,);
not I_81530 (I1388541,I1388533);
nand I_81531 (I1388558,I1388541,I1388281);
not I_81532 (I1388032,I1388558);
nand I_81533 (I1388026,I1388558,I1388298);
nand I_81534 (I1388023,I1388541,I1388165);
not I_81535 (I1388647,I2514);
DFFARX1 I_81536 (I210920,I2507,I1388647,I1388673,);
DFFARX1 I_81537 (I210923,I2507,I1388647,I1388690,);
not I_81538 (I1388698,I1388690);
nor I_81539 (I1388615,I1388673,I1388698);
DFFARX1 I_81540 (I1388698,I2507,I1388647,I1388630,);
nor I_81541 (I1388743,I210929,I210923);
and I_81542 (I1388760,I1388743,I210926);
nor I_81543 (I1388777,I1388760,I210929);
not I_81544 (I1388794,I210929);
and I_81545 (I1388811,I1388794,I210920);
nand I_81546 (I1388828,I1388811,I210938);
nor I_81547 (I1388845,I1388794,I1388828);
DFFARX1 I_81548 (I1388845,I2507,I1388647,I1388612,);
not I_81549 (I1388876,I1388828);
nand I_81550 (I1388893,I1388698,I1388876);
nand I_81551 (I1388624,I1388760,I1388876);
DFFARX1 I_81552 (I1388794,I2507,I1388647,I1388639,);
not I_81553 (I1388938,I210932);
nor I_81554 (I1388955,I1388938,I210920);
nor I_81555 (I1388972,I1388955,I1388777);
DFFARX1 I_81556 (I1388972,I2507,I1388647,I1388636,);
not I_81557 (I1389003,I1388955);
DFFARX1 I_81558 (I1389003,I2507,I1388647,I1389029,);
not I_81559 (I1389037,I1389029);
nor I_81560 (I1388633,I1389037,I1388955);
nor I_81561 (I1389068,I1388938,I210935);
and I_81562 (I1389085,I1389068,I210941);
or I_81563 (I1389102,I1389085,I210944);
DFFARX1 I_81564 (I1389102,I2507,I1388647,I1389128,);
not I_81565 (I1389136,I1389128);
nand I_81566 (I1389153,I1389136,I1388876);
not I_81567 (I1388627,I1389153);
nand I_81568 (I1388621,I1389153,I1388893);
nand I_81569 (I1388618,I1389136,I1388760);
not I_81570 (I1389242,I2514);
DFFARX1 I_81571 (I701255,I2507,I1389242,I1389268,);
DFFARX1 I_81572 (I701237,I2507,I1389242,I1389285,);
not I_81573 (I1389293,I1389285);
nor I_81574 (I1389210,I1389268,I1389293);
DFFARX1 I_81575 (I1389293,I2507,I1389242,I1389225,);
nor I_81576 (I1389338,I701243,I701246);
and I_81577 (I1389355,I1389338,I701234);
nor I_81578 (I1389372,I1389355,I701243);
not I_81579 (I1389389,I701243);
and I_81580 (I1389406,I1389389,I701252);
nand I_81581 (I1389423,I1389406,I701240);
nor I_81582 (I1389440,I1389389,I1389423);
DFFARX1 I_81583 (I1389440,I2507,I1389242,I1389207,);
not I_81584 (I1389471,I1389423);
nand I_81585 (I1389488,I1389293,I1389471);
nand I_81586 (I1389219,I1389355,I1389471);
DFFARX1 I_81587 (I1389389,I2507,I1389242,I1389234,);
not I_81588 (I1389533,I701237);
nor I_81589 (I1389550,I1389533,I701252);
nor I_81590 (I1389567,I1389550,I1389372);
DFFARX1 I_81591 (I1389567,I2507,I1389242,I1389231,);
not I_81592 (I1389598,I1389550);
DFFARX1 I_81593 (I1389598,I2507,I1389242,I1389624,);
not I_81594 (I1389632,I1389624);
nor I_81595 (I1389228,I1389632,I1389550);
nor I_81596 (I1389663,I1389533,I701249);
and I_81597 (I1389680,I1389663,I701258);
or I_81598 (I1389697,I1389680,I701234);
DFFARX1 I_81599 (I1389697,I2507,I1389242,I1389723,);
not I_81600 (I1389731,I1389723);
nand I_81601 (I1389748,I1389731,I1389471);
not I_81602 (I1389222,I1389748);
nand I_81603 (I1389216,I1389748,I1389488);
nand I_81604 (I1389213,I1389731,I1389355);
not I_81605 (I1389837,I2514);
DFFARX1 I_81606 (I511344,I2507,I1389837,I1389863,);
DFFARX1 I_81607 (I511347,I2507,I1389837,I1389880,);
not I_81608 (I1389888,I1389880);
nor I_81609 (I1389805,I1389863,I1389888);
DFFARX1 I_81610 (I1389888,I2507,I1389837,I1389820,);
nor I_81611 (I1389933,I511350,I511368);
and I_81612 (I1389950,I1389933,I511353);
nor I_81613 (I1389967,I1389950,I511350);
not I_81614 (I1389984,I511350);
and I_81615 (I1390001,I1389984,I511362);
nand I_81616 (I1390018,I1390001,I511365);
nor I_81617 (I1390035,I1389984,I1390018);
DFFARX1 I_81618 (I1390035,I2507,I1389837,I1389802,);
not I_81619 (I1390066,I1390018);
nand I_81620 (I1390083,I1389888,I1390066);
nand I_81621 (I1389814,I1389950,I1390066);
DFFARX1 I_81622 (I1389984,I2507,I1389837,I1389829,);
not I_81623 (I1390128,I511356);
nor I_81624 (I1390145,I1390128,I511362);
nor I_81625 (I1390162,I1390145,I1389967);
DFFARX1 I_81626 (I1390162,I2507,I1389837,I1389826,);
not I_81627 (I1390193,I1390145);
DFFARX1 I_81628 (I1390193,I2507,I1389837,I1390219,);
not I_81629 (I1390227,I1390219);
nor I_81630 (I1389823,I1390227,I1390145);
nor I_81631 (I1390258,I1390128,I511344);
and I_81632 (I1390275,I1390258,I511359);
or I_81633 (I1390292,I1390275,I511347);
DFFARX1 I_81634 (I1390292,I2507,I1389837,I1390318,);
not I_81635 (I1390326,I1390318);
nand I_81636 (I1390343,I1390326,I1390066);
not I_81637 (I1389817,I1390343);
nand I_81638 (I1389811,I1390343,I1390083);
nand I_81639 (I1389808,I1390326,I1389950);
not I_81640 (I1390432,I2514);
DFFARX1 I_81641 (I1117329,I2507,I1390432,I1390458,);
DFFARX1 I_81642 (I1117341,I2507,I1390432,I1390475,);
not I_81643 (I1390483,I1390475);
nor I_81644 (I1390400,I1390458,I1390483);
DFFARX1 I_81645 (I1390483,I2507,I1390432,I1390415,);
nor I_81646 (I1390528,I1117338,I1117332);
and I_81647 (I1390545,I1390528,I1117326);
nor I_81648 (I1390562,I1390545,I1117338);
not I_81649 (I1390579,I1117338);
and I_81650 (I1390596,I1390579,I1117335);
nand I_81651 (I1390613,I1390596,I1117326);
nor I_81652 (I1390630,I1390579,I1390613);
DFFARX1 I_81653 (I1390630,I2507,I1390432,I1390397,);
not I_81654 (I1390661,I1390613);
nand I_81655 (I1390678,I1390483,I1390661);
nand I_81656 (I1390409,I1390545,I1390661);
DFFARX1 I_81657 (I1390579,I2507,I1390432,I1390424,);
not I_81658 (I1390723,I1117350);
nor I_81659 (I1390740,I1390723,I1117335);
nor I_81660 (I1390757,I1390740,I1390562);
DFFARX1 I_81661 (I1390757,I2507,I1390432,I1390421,);
not I_81662 (I1390788,I1390740);
DFFARX1 I_81663 (I1390788,I2507,I1390432,I1390814,);
not I_81664 (I1390822,I1390814);
nor I_81665 (I1390418,I1390822,I1390740);
nor I_81666 (I1390853,I1390723,I1117344);
and I_81667 (I1390870,I1390853,I1117347);
or I_81668 (I1390887,I1390870,I1117329);
DFFARX1 I_81669 (I1390887,I2507,I1390432,I1390913,);
not I_81670 (I1390921,I1390913);
nand I_81671 (I1390938,I1390921,I1390661);
not I_81672 (I1390412,I1390938);
nand I_81673 (I1390406,I1390938,I1390678);
nand I_81674 (I1390403,I1390921,I1390545);
not I_81675 (I1391027,I2514);
DFFARX1 I_81676 (I619757,I2507,I1391027,I1391053,);
DFFARX1 I_81677 (I619751,I2507,I1391027,I1391070,);
not I_81678 (I1391078,I1391070);
nor I_81679 (I1390995,I1391053,I1391078);
DFFARX1 I_81680 (I1391078,I2507,I1391027,I1391010,);
nor I_81681 (I1391123,I619748,I619739);
and I_81682 (I1391140,I1391123,I619736);
nor I_81683 (I1391157,I1391140,I619748);
not I_81684 (I1391174,I619748);
and I_81685 (I1391191,I1391174,I619742);
nand I_81686 (I1391208,I1391191,I619754);
nor I_81687 (I1391225,I1391174,I1391208);
DFFARX1 I_81688 (I1391225,I2507,I1391027,I1390992,);
not I_81689 (I1391256,I1391208);
nand I_81690 (I1391273,I1391078,I1391256);
nand I_81691 (I1391004,I1391140,I1391256);
DFFARX1 I_81692 (I1391174,I2507,I1391027,I1391019,);
not I_81693 (I1391318,I619760);
nor I_81694 (I1391335,I1391318,I619742);
nor I_81695 (I1391352,I1391335,I1391157);
DFFARX1 I_81696 (I1391352,I2507,I1391027,I1391016,);
not I_81697 (I1391383,I1391335);
DFFARX1 I_81698 (I1391383,I2507,I1391027,I1391409,);
not I_81699 (I1391417,I1391409);
nor I_81700 (I1391013,I1391417,I1391335);
nor I_81701 (I1391448,I1391318,I619739);
and I_81702 (I1391465,I1391448,I619745);
or I_81703 (I1391482,I1391465,I619736);
DFFARX1 I_81704 (I1391482,I2507,I1391027,I1391508,);
not I_81705 (I1391516,I1391508);
nand I_81706 (I1391533,I1391516,I1391256);
not I_81707 (I1391007,I1391533);
nand I_81708 (I1391001,I1391533,I1391273);
nand I_81709 (I1390998,I1391516,I1391140);
not I_81710 (I1391622,I2514);
DFFARX1 I_81711 (I352449,I2507,I1391622,I1391648,);
DFFARX1 I_81712 (I352443,I2507,I1391622,I1391665,);
not I_81713 (I1391673,I1391665);
nor I_81714 (I1391590,I1391648,I1391673);
DFFARX1 I_81715 (I1391673,I2507,I1391622,I1391605,);
nor I_81716 (I1391718,I352431,I352452);
and I_81717 (I1391735,I1391718,I352446);
nor I_81718 (I1391752,I1391735,I352431);
not I_81719 (I1391769,I352431);
and I_81720 (I1391786,I1391769,I352428);
nand I_81721 (I1391803,I1391786,I352440);
nor I_81722 (I1391820,I1391769,I1391803);
DFFARX1 I_81723 (I1391820,I2507,I1391622,I1391587,);
not I_81724 (I1391851,I1391803);
nand I_81725 (I1391868,I1391673,I1391851);
nand I_81726 (I1391599,I1391735,I1391851);
DFFARX1 I_81727 (I1391769,I2507,I1391622,I1391614,);
not I_81728 (I1391913,I352455);
nor I_81729 (I1391930,I1391913,I352428);
nor I_81730 (I1391947,I1391930,I1391752);
DFFARX1 I_81731 (I1391947,I2507,I1391622,I1391611,);
not I_81732 (I1391978,I1391930);
DFFARX1 I_81733 (I1391978,I2507,I1391622,I1392004,);
not I_81734 (I1392012,I1392004);
nor I_81735 (I1391608,I1392012,I1391930);
nor I_81736 (I1392043,I1391913,I352437);
and I_81737 (I1392060,I1392043,I352434);
or I_81738 (I1392077,I1392060,I352428);
DFFARX1 I_81739 (I1392077,I2507,I1391622,I1392103,);
not I_81740 (I1392111,I1392103);
nand I_81741 (I1392128,I1392111,I1391851);
not I_81742 (I1391602,I1392128);
nand I_81743 (I1391596,I1392128,I1391868);
nand I_81744 (I1391593,I1392111,I1391735);
not I_81745 (I1392217,I2514);
DFFARX1 I_81746 (I179385,I2507,I1392217,I1392243,);
DFFARX1 I_81747 (I179388,I2507,I1392217,I1392260,);
not I_81748 (I1392268,I1392260);
nor I_81749 (I1392185,I1392243,I1392268);
DFFARX1 I_81750 (I1392268,I2507,I1392217,I1392200,);
nor I_81751 (I1392313,I179394,I179388);
and I_81752 (I1392330,I1392313,I179391);
nor I_81753 (I1392347,I1392330,I179394);
not I_81754 (I1392364,I179394);
and I_81755 (I1392381,I1392364,I179385);
nand I_81756 (I1392398,I1392381,I179403);
nor I_81757 (I1392415,I1392364,I1392398);
DFFARX1 I_81758 (I1392415,I2507,I1392217,I1392182,);
not I_81759 (I1392446,I1392398);
nand I_81760 (I1392463,I1392268,I1392446);
nand I_81761 (I1392194,I1392330,I1392446);
DFFARX1 I_81762 (I1392364,I2507,I1392217,I1392209,);
not I_81763 (I1392508,I179397);
nor I_81764 (I1392525,I1392508,I179385);
nor I_81765 (I1392542,I1392525,I1392347);
DFFARX1 I_81766 (I1392542,I2507,I1392217,I1392206,);
not I_81767 (I1392573,I1392525);
DFFARX1 I_81768 (I1392573,I2507,I1392217,I1392599,);
not I_81769 (I1392607,I1392599);
nor I_81770 (I1392203,I1392607,I1392525);
nor I_81771 (I1392638,I1392508,I179400);
and I_81772 (I1392655,I1392638,I179406);
or I_81773 (I1392672,I1392655,I179409);
DFFARX1 I_81774 (I1392672,I2507,I1392217,I1392698,);
not I_81775 (I1392706,I1392698);
nand I_81776 (I1392723,I1392706,I1392446);
not I_81777 (I1392197,I1392723);
nand I_81778 (I1392191,I1392723,I1392463);
nand I_81779 (I1392188,I1392706,I1392330);
not I_81780 (I1392812,I2514);
DFFARX1 I_81781 (I862862,I2507,I1392812,I1392838,);
DFFARX1 I_81782 (I862859,I2507,I1392812,I1392855,);
not I_81783 (I1392863,I1392855);
nor I_81784 (I1392780,I1392838,I1392863);
DFFARX1 I_81785 (I1392863,I2507,I1392812,I1392795,);
nor I_81786 (I1392908,I862874,I862856);
and I_81787 (I1392925,I1392908,I862853);
nor I_81788 (I1392942,I1392925,I862874);
not I_81789 (I1392959,I862874);
and I_81790 (I1392976,I1392959,I862859);
nand I_81791 (I1392993,I1392976,I862871);
nor I_81792 (I1393010,I1392959,I1392993);
DFFARX1 I_81793 (I1393010,I2507,I1392812,I1392777,);
not I_81794 (I1393041,I1392993);
nand I_81795 (I1393058,I1392863,I1393041);
nand I_81796 (I1392789,I1392925,I1393041);
DFFARX1 I_81797 (I1392959,I2507,I1392812,I1392804,);
not I_81798 (I1393103,I862865);
nor I_81799 (I1393120,I1393103,I862859);
nor I_81800 (I1393137,I1393120,I1392942);
DFFARX1 I_81801 (I1393137,I2507,I1392812,I1392801,);
not I_81802 (I1393168,I1393120);
DFFARX1 I_81803 (I1393168,I2507,I1392812,I1393194,);
not I_81804 (I1393202,I1393194);
nor I_81805 (I1392798,I1393202,I1393120);
nor I_81806 (I1393233,I1393103,I862853);
and I_81807 (I1393250,I1393233,I862868);
or I_81808 (I1393267,I1393250,I862856);
DFFARX1 I_81809 (I1393267,I2507,I1392812,I1393293,);
not I_81810 (I1393301,I1393293);
nand I_81811 (I1393318,I1393301,I1393041);
not I_81812 (I1392792,I1393318);
nand I_81813 (I1392786,I1393318,I1393058);
nand I_81814 (I1392783,I1393301,I1392925);
not I_81815 (I1393407,I2514);
DFFARX1 I_81816 (I982539,I2507,I1393407,I1393433,);
DFFARX1 I_81817 (I982557,I2507,I1393407,I1393450,);
not I_81818 (I1393458,I1393450);
nor I_81819 (I1393375,I1393433,I1393458);
DFFARX1 I_81820 (I1393458,I2507,I1393407,I1393390,);
nor I_81821 (I1393503,I982536,I982548);
and I_81822 (I1393520,I1393503,I982533);
nor I_81823 (I1393537,I1393520,I982536);
not I_81824 (I1393554,I982536);
and I_81825 (I1393571,I1393554,I982542);
nand I_81826 (I1393588,I1393571,I982554);
nor I_81827 (I1393605,I1393554,I1393588);
DFFARX1 I_81828 (I1393605,I2507,I1393407,I1393372,);
not I_81829 (I1393636,I1393588);
nand I_81830 (I1393653,I1393458,I1393636);
nand I_81831 (I1393384,I1393520,I1393636);
DFFARX1 I_81832 (I1393554,I2507,I1393407,I1393399,);
not I_81833 (I1393698,I982545);
nor I_81834 (I1393715,I1393698,I982542);
nor I_81835 (I1393732,I1393715,I1393537);
DFFARX1 I_81836 (I1393732,I2507,I1393407,I1393396,);
not I_81837 (I1393763,I1393715);
DFFARX1 I_81838 (I1393763,I2507,I1393407,I1393789,);
not I_81839 (I1393797,I1393789);
nor I_81840 (I1393393,I1393797,I1393715);
nor I_81841 (I1393828,I1393698,I982533);
and I_81842 (I1393845,I1393828,I982560);
or I_81843 (I1393862,I1393845,I982551);
DFFARX1 I_81844 (I1393862,I2507,I1393407,I1393888,);
not I_81845 (I1393896,I1393888);
nand I_81846 (I1393913,I1393896,I1393636);
not I_81847 (I1393387,I1393913);
nand I_81848 (I1393381,I1393913,I1393653);
nand I_81849 (I1393378,I1393896,I1393520);
not I_81850 (I1394002,I2514);
DFFARX1 I_81851 (I214490,I2507,I1394002,I1394028,);
DFFARX1 I_81852 (I214493,I2507,I1394002,I1394045,);
not I_81853 (I1394053,I1394045);
nor I_81854 (I1393970,I1394028,I1394053);
DFFARX1 I_81855 (I1394053,I2507,I1394002,I1393985,);
nor I_81856 (I1394098,I214499,I214493);
and I_81857 (I1394115,I1394098,I214496);
nor I_81858 (I1394132,I1394115,I214499);
not I_81859 (I1394149,I214499);
and I_81860 (I1394166,I1394149,I214490);
nand I_81861 (I1394183,I1394166,I214508);
nor I_81862 (I1394200,I1394149,I1394183);
DFFARX1 I_81863 (I1394200,I2507,I1394002,I1393967,);
not I_81864 (I1394231,I1394183);
nand I_81865 (I1394248,I1394053,I1394231);
nand I_81866 (I1393979,I1394115,I1394231);
DFFARX1 I_81867 (I1394149,I2507,I1394002,I1393994,);
not I_81868 (I1394293,I214502);
nor I_81869 (I1394310,I1394293,I214490);
nor I_81870 (I1394327,I1394310,I1394132);
DFFARX1 I_81871 (I1394327,I2507,I1394002,I1393991,);
not I_81872 (I1394358,I1394310);
DFFARX1 I_81873 (I1394358,I2507,I1394002,I1394384,);
not I_81874 (I1394392,I1394384);
nor I_81875 (I1393988,I1394392,I1394310);
nor I_81876 (I1394423,I1394293,I214505);
and I_81877 (I1394440,I1394423,I214511);
or I_81878 (I1394457,I1394440,I214514);
DFFARX1 I_81879 (I1394457,I2507,I1394002,I1394483,);
not I_81880 (I1394491,I1394483);
nand I_81881 (I1394508,I1394491,I1394231);
not I_81882 (I1393982,I1394508);
nand I_81883 (I1393976,I1394508,I1394248);
nand I_81884 (I1393973,I1394491,I1394115);
not I_81885 (I1394597,I2514);
DFFARX1 I_81886 (I675245,I2507,I1394597,I1394623,);
DFFARX1 I_81887 (I675227,I2507,I1394597,I1394640,);
not I_81888 (I1394648,I1394640);
nor I_81889 (I1394565,I1394623,I1394648);
DFFARX1 I_81890 (I1394648,I2507,I1394597,I1394580,);
nor I_81891 (I1394693,I675233,I675236);
and I_81892 (I1394710,I1394693,I675224);
nor I_81893 (I1394727,I1394710,I675233);
not I_81894 (I1394744,I675233);
and I_81895 (I1394761,I1394744,I675242);
nand I_81896 (I1394778,I1394761,I675230);
nor I_81897 (I1394795,I1394744,I1394778);
DFFARX1 I_81898 (I1394795,I2507,I1394597,I1394562,);
not I_81899 (I1394826,I1394778);
nand I_81900 (I1394843,I1394648,I1394826);
nand I_81901 (I1394574,I1394710,I1394826);
DFFARX1 I_81902 (I1394744,I2507,I1394597,I1394589,);
not I_81903 (I1394888,I675227);
nor I_81904 (I1394905,I1394888,I675242);
nor I_81905 (I1394922,I1394905,I1394727);
DFFARX1 I_81906 (I1394922,I2507,I1394597,I1394586,);
not I_81907 (I1394953,I1394905);
DFFARX1 I_81908 (I1394953,I2507,I1394597,I1394979,);
not I_81909 (I1394987,I1394979);
nor I_81910 (I1394583,I1394987,I1394905);
nor I_81911 (I1395018,I1394888,I675239);
and I_81912 (I1395035,I1395018,I675248);
or I_81913 (I1395052,I1395035,I675224);
DFFARX1 I_81914 (I1395052,I2507,I1394597,I1395078,);
not I_81915 (I1395086,I1395078);
nand I_81916 (I1395103,I1395086,I1394826);
not I_81917 (I1394577,I1395103);
nand I_81918 (I1394571,I1395103,I1394843);
nand I_81919 (I1394568,I1395086,I1394710);
not I_81920 (I1395192,I2514);
DFFARX1 I_81921 (I453935,I2507,I1395192,I1395218,);
DFFARX1 I_81922 (I453941,I2507,I1395192,I1395235,);
not I_81923 (I1395243,I1395235);
nor I_81924 (I1395160,I1395218,I1395243);
DFFARX1 I_81925 (I1395243,I2507,I1395192,I1395175,);
nor I_81926 (I1395288,I453950,I453935);
and I_81927 (I1395305,I1395288,I453962);
nor I_81928 (I1395322,I1395305,I453950);
not I_81929 (I1395339,I453950);
and I_81930 (I1395356,I1395339,I453938);
nand I_81931 (I1395373,I1395356,I453959);
nor I_81932 (I1395390,I1395339,I1395373);
DFFARX1 I_81933 (I1395390,I2507,I1395192,I1395157,);
not I_81934 (I1395421,I1395373);
nand I_81935 (I1395438,I1395243,I1395421);
nand I_81936 (I1395169,I1395305,I1395421);
DFFARX1 I_81937 (I1395339,I2507,I1395192,I1395184,);
not I_81938 (I1395483,I453947);
nor I_81939 (I1395500,I1395483,I453938);
nor I_81940 (I1395517,I1395500,I1395322);
DFFARX1 I_81941 (I1395517,I2507,I1395192,I1395181,);
not I_81942 (I1395548,I1395500);
DFFARX1 I_81943 (I1395548,I2507,I1395192,I1395574,);
not I_81944 (I1395582,I1395574);
nor I_81945 (I1395178,I1395582,I1395500);
nor I_81946 (I1395613,I1395483,I453944);
and I_81947 (I1395630,I1395613,I453956);
or I_81948 (I1395647,I1395630,I453953);
DFFARX1 I_81949 (I1395647,I2507,I1395192,I1395673,);
not I_81950 (I1395681,I1395673);
nand I_81951 (I1395698,I1395681,I1395421);
not I_81952 (I1395172,I1395698);
nand I_81953 (I1395166,I1395698,I1395438);
nand I_81954 (I1395163,I1395681,I1395305);
not I_81955 (I1395787,I2514);
DFFARX1 I_81956 (I263913,I2507,I1395787,I1395813,);
DFFARX1 I_81957 (I263907,I2507,I1395787,I1395830,);
not I_81958 (I1395838,I1395830);
nor I_81959 (I1395755,I1395813,I1395838);
DFFARX1 I_81960 (I1395838,I2507,I1395787,I1395770,);
nor I_81961 (I1395883,I263895,I263916);
and I_81962 (I1395900,I1395883,I263910);
nor I_81963 (I1395917,I1395900,I263895);
not I_81964 (I1395934,I263895);
and I_81965 (I1395951,I1395934,I263892);
nand I_81966 (I1395968,I1395951,I263904);
nor I_81967 (I1395985,I1395934,I1395968);
DFFARX1 I_81968 (I1395985,I2507,I1395787,I1395752,);
not I_81969 (I1396016,I1395968);
nand I_81970 (I1396033,I1395838,I1396016);
nand I_81971 (I1395764,I1395900,I1396016);
DFFARX1 I_81972 (I1395934,I2507,I1395787,I1395779,);
not I_81973 (I1396078,I263919);
nor I_81974 (I1396095,I1396078,I263892);
nor I_81975 (I1396112,I1396095,I1395917);
DFFARX1 I_81976 (I1396112,I2507,I1395787,I1395776,);
not I_81977 (I1396143,I1396095);
DFFARX1 I_81978 (I1396143,I2507,I1395787,I1396169,);
not I_81979 (I1396177,I1396169);
nor I_81980 (I1395773,I1396177,I1396095);
nor I_81981 (I1396208,I1396078,I263901);
and I_81982 (I1396225,I1396208,I263898);
or I_81983 (I1396242,I1396225,I263892);
DFFARX1 I_81984 (I1396242,I2507,I1395787,I1396268,);
not I_81985 (I1396276,I1396268);
nand I_81986 (I1396293,I1396276,I1396016);
not I_81987 (I1395767,I1396293);
nand I_81988 (I1395761,I1396293,I1396033);
nand I_81989 (I1395758,I1396276,I1395900);
endmodule


