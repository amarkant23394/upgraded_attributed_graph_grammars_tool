module test_I14004(I1477,I12493,I1470,I12191,I14004);
input I1477,I12493,I1470,I12191;
output I14004;
wire I11935,I11950,I12208,I13775,I13987,I11973,I13970,I11941;
DFFARX1 I_0(I12208,I1470,I11973,,,I11935,);
DFFARX1 I_1(I12493,I1470,I11973,,,I11950,);
DFFARX1 I_2(I13987,I1470,I13775,,,I14004,);
DFFARX1 I_3(I12191,I1470,I11973,,,I12208,);
not I_4(I13775,I1477);
and I_5(I13987,I13970,I11941);
not I_6(I11973,I1477);
nand I_7(I13970,I11935,I11950);
DFFARX1 I_8(I12208,I1470,I11973,,,I11941,);
endmodule


