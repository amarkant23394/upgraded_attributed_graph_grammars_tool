module test_I1393(I1287,I1215,I1223,I1393);
input I1287,I1215,I1223;
output I1393;
wire I1376;
nor I_0(I1376,I1215,I1223);
nand I_1(I1393,I1376,I1287);
endmodule


