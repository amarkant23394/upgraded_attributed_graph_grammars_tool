module test_I16934(I12584,I12930,I1477,I1470,I16934);
input I12584,I12930,I1477,I1470;
output I16934;
wire I12602,I15109,I14945,I16818,I15126,I14965,I15372;
not I_0(I12602,I12930);
DFFARX1 I_1(I14945,I1470,I16818,,,I16934,);
not I_2(I15109,I12584);
nand I_3(I14945,I15372,I15126);
not I_4(I16818,I1477);
not I_5(I15126,I15109);
not I_6(I14965,I1477);
DFFARX1 I_7(I12602,I1470,I14965,,,I15372,);
endmodule


