module test_I9638(I8527,I1477,I5737,I1470,I5740,I9638);
input I8527,I1477,I5737,I1470,I5740;
output I9638;
wire I8202,I8496,I8216,I8298,I5719,I8377,I8250,I8315,I9491,I8181,I8360,I8592,I8205,I8462,I9576,I8267,I9621;
nand I_0(I8202,I8267,I8496);
nor I_1(I8496,I8462,I8377);
not I_2(I8216,I1477);
nor I_3(I9638,I9621,I9576);
nor I_4(I8298,I5719);
DFFARX1 I_5(I1470,,,I5719,);
not I_6(I8377,I8360);
nor I_7(I8250,I5719);
nand I_8(I8315,I8298,I5740);
not I_9(I9491,I1477);
and I_10(I8181,I8360,I8592);
not I_11(I8360,I5719);
DFFARX1 I_12(I8527,I1470,I8216,,,I8592,);
not I_13(I8205,I8315);
DFFARX1 I_14(I1470,I8216,,,I8462,);
nor I_15(I9576,I8181,I8202);
nand I_16(I8267,I8250,I5737);
DFFARX1 I_17(I8205,I1470,I9491,,,I9621,);
endmodule


