module test_I12174(I7621,I1477,I7850,I1470,I12174);
input I7621,I1477,I7850,I1470;
output I12174;
wire I7556,I12140,I10219,I10583,I10014,I10052,I12157,I10490,I10017,I10035;
nand I_0(I7556,I7621,I7850);
not I_1(I12140,I10014);
DFFARX1 I_2(I1470,I10052,,,I10219,);
DFFARX1 I_3(I10490,I1470,I10052,,,I10583,);
DFFARX1 I_4(I10219,I1470,I10052,,,I10014,);
not I_5(I10052,I1477);
nor I_6(I12157,I12140,I10035);
DFFARX1 I_7(I7556,I1470,I10052,,,I10490,);
and I_8(I10017,I10490,I10583);
and I_9(I12174,I12157,I10017);
not I_10(I10035,I10490);
endmodule


