module test_I1507(I1215,I1423,I1455,I1507);
input I1215,I1423,I1455;
output I1507;
wire I1637,I1586,I1603,I1535;
not I_0(I1637,I1215);
nor I_1(I1507,I1603,I1637);
nor I_2(I1586,I1535,I1215);
nand I_3(I1603,I1586,I1423);
not I_4(I1535,I1455);
endmodule


