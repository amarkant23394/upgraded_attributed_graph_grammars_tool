module test_I3521(I1477,I1470,I1832,I3521);
input I1477,I1470,I1832;
output I3521;
wire I1518,I1486,I1801,I1784,I2038,I3504,I2021,I1849,I1495,I1489,I2103,I3487,I1767;
not I_0(I1518,I1477);
DFFARX1 I_1(I1832,I1470,I1518,,,I1486,);
DFFARX1 I_2(I1767,I1470,I1518,,,I1801,);
nor I_3(I1784,I1767);
not I_4(I2038,I2021);
nor I_5(I3521,I3504,I1495);
and I_6(I3504,I3487,I1489);
DFFARX1 I_7(I1470,I1518,,,I2021,);
and I_8(I1849,I1832,I1784);
DFFARX1 I_9(I2103,I1470,I1518,,,I1495,);
not I_10(I1489,I1801);
or I_11(I2103,I2038,I1849);
not I_12(I3487,I1486);
DFFARX1 I_13(I1470,I1518,,,I1767,);
endmodule


