module test_final(G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_569_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0,n4_1_l_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_0,blif_clk_net_1_r_4,n6_4,G42_1_r_0,);
nor I_1(n_572_1_r_0,IN_5_1_l_0,n23_0);
nand I_2(n_573_1_r_0,n21_0,n22_0);
nand I_3(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_4(n_569_1_r_0,n21_0,n26_0);
nor I_5(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_6(N3_2_r_0,blif_clk_net_1_r_4,n6_4,G199_2_r_0,);
DFFARX1 I_7(N1_4_r_0,blif_clk_net_1_r_4,n6_4,G199_4_r_0,);
DFFARX1 I_8(n2_0,blif_clk_net_1_r_4,n6_4,G214_4_r_0,);
nor I_9(n4_1_l_0,G18_1_l_0,IN_1_1_l_0);
DFFARX1 I_10(n4_1_l_0,blif_clk_net_1_r_4,n6_4,n37_0,);
DFFARX1 I_11(IN_1_3_l_0,blif_clk_net_1_r_4,n6_4,n38_0,);
not I_12(n20_0,n38_0);
DFFARX1 I_13(IN_2_3_l_0,blif_clk_net_1_r_4,n6_4,ACVQN1_3_l_0,);
nor I_14(n4_1_r_0,IN_10_1_l_0,n23_0);
nor I_15(N3_2_r_0,n31_0,n32_0);
nor I_16(N1_4_r_0,n29_0,n32_0);
not I_17(n2_0,n31_0);
nor I_18(n21_0,IN_9_1_l_0,n37_0);
not I_19(n22_0,IN_5_1_l_0);
nand I_20(n23_0,n20_0,n30_0);
nand I_21(n24_0,n38_0,n25_0);
nor I_22(n25_0,IN_9_1_l_0,IN_10_1_l_0);
not I_23(n26_0,IN_10_1_l_0);
not I_24(n27_0,n29_0);
nor I_25(n28_0,G15_1_l_0,IN_7_1_l_0);
nand I_26(n29_0,n26_0,n33_0);
not I_27(n30_0,IN_9_1_l_0);
nand I_28(n31_0,IN_4_3_l_0,ACVQN1_3_l_0);
and I_29(n32_0,n35_0,n36_0);
nand I_30(n33_0,IN_4_1_l_0,n34_0);
not I_31(n34_0,G15_1_l_0);
nor I_32(n35_0,G18_1_l_0,G15_1_l_0);
nor I_33(n36_0,IN_5_1_l_0,IN_7_1_l_0);
DFFARX1 I_34(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_35(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_36(n_573_1_r_4,n16_4,G199_2_r_0);
nor I_37(n_549_1_r_4,n22_4,n23_4);
nand I_38(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_39(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_40(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_41(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_42(P6_5_r_4,P6_5_r_internal_4);
or I_43(n_431_0_l_4,n26_4,n_573_1_r_0);
not I_44(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_45(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_46(n_573_1_r_0,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_47(n16_4,ACVQN1_5_l_4);
DFFARX1 I_48(n_572_1_r_0,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_49(n17_4,n17_internal_4);
nor I_50(n4_1_r_4,n30_4,n31_4);
nand I_51(n19_4,n33_4,G42_1_r_0);
DFFARX1 I_52(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_53(n15_4,n15_internal_4);
DFFARX1 I_54(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_55(n20_4,n16_4,G214_4_r_0);
nor I_56(n21_4,n_549_1_r_0,G199_2_r_0);
nand I_57(n22_4,G78_0_l_4,n25_4);
nand I_58(n23_4,n24_4,G214_4_r_0);
not I_59(n24_4,G199_2_r_0);
not I_60(n25_4,n_549_1_r_0);
and I_61(n26_4,n27_4,G42_1_r_0);
nor I_62(n27_4,n28_4,n_572_1_r_0);
not I_63(n28_4,G42_1_r_0);
not I_64(n29_4,n30_4);
nand I_65(n30_4,n32_4,G199_4_r_0);
nand I_66(n31_4,n25_4,G214_4_r_0);
nor I_67(n32_4,n33_4,G199_2_r_0);
not I_68(n33_4,n_42_2_r_0);
endmodule


