module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_7_r_2,n10_2,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_7_r_2,n10_2,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_7_r_2,n10_2,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_7_r_2,n10_2,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
nor I_43(N1371_0_r_2,n32_2,n35_2);
nor I_44(N1508_0_r_2,n32_2,n55_2);
not I_45(N1372_1_r_2,n54_2);
nor I_46(N1508_1_r_2,n59_2,n54_2);
nor I_47(N6147_2_r_2,n42_2,n43_2);
nor I_48(N1507_6_r_2,n40_2,n53_2);
nor I_49(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_50(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_51(n_572_7_r_2,n36_2,n37_2);
or I_52(n_573_7_r_2,n34_2,n35_2);
nor I_53(n_549_7_r_2,n40_2,n41_2);
nand I_54(n_569_7_r_2,n38_2,n39_2);
nor I_55(n_452_7_r_2,n59_2,n35_2);
nor I_56(n4_7_l_2,n_42_8_r_9,N1372_4_r_9);
not I_57(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_58(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_59(n33_2,n59_2);
and I_60(N3_8_l_2,n49_2,G199_8_r_9);
DFFARX1 I_61(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_62(n32_2,n32_internal_2);
nor I_63(n4_7_r_2,n59_2,n36_2);
not I_64(n34_2,n39_2);
nor I_65(n35_2,n_547_5_r_9,N6134_9_r_9);
nor I_66(n36_2,N6147_2_r_9,N1372_4_r_9);
or I_67(n37_2,N1508_4_r_9,G78_5_r_9);
not I_68(n38_2,n40_2);
nand I_69(n39_2,n45_2,n57_2);
nor I_70(n40_2,n47_2,G78_5_r_9);
nor I_71(n41_2,n32_2,n36_2);
not I_72(n42_2,n53_2);
nand I_73(n43_2,n44_2,n45_2);
nand I_74(n44_2,n38_2,n46_2);
not I_75(n45_2,G78_5_r_9);
nand I_76(n46_2,n47_2,n48_2);
nand I_77(n47_2,G199_8_r_9,N6147_9_r_9);
or I_78(n48_2,n_576_5_r_9,n_547_5_r_9);
nand I_79(n49_2,n_547_5_r_9,n_42_8_r_9);
nand I_80(n50_2,n51_2,n52_2);
not I_81(n51_2,n47_2);
nand I_82(n52_2,n38_2,n53_2);
nor I_83(n53_2,N6147_2_r_9,N1508_4_r_9);
nand I_84(n54_2,n42_2,n56_2);
nor I_85(n55_2,n34_2,n56_2);
nor I_86(n56_2,n_576_5_r_9,n_547_5_r_9);
nand I_87(n57_2,n58_2,N1372_4_r_9);
not I_88(n58_2,n_576_5_r_9);
endmodule


