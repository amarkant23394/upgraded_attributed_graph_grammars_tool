module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_7_r_1,n9_1,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_7_r_1,n9_1,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
and I_35(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_36(N1508_0_r_1,n40_1,n44_1);
nor I_37(N1507_6_r_1,n43_1,n49_1);
nor I_38(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_39(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_40(n_572_7_r_1,n29_1,n30_1);
not I_41(n_573_7_r_1,n_452_7_r_1);
nor I_42(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_43(n_569_7_r_1,n30_1,n31_1);
nor I_44(n_452_7_r_1,n30_1,n32_1);
nor I_45(N6147_9_r_1,n35_1,n36_1);
nand I_46(N6134_9_r_1,n38_1,n39_1);
not I_47(I_BUFF_1_9_r_1,n40_1);
nor I_48(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_49(n9_1,blif_reset_net_7_r_1);
nor I_50(n29_1,n34_1,n_569_7_r_0);
nor I_51(n30_1,n33_1,n34_1);
nor I_52(n31_1,n54_1,n_573_7_r_0);
not I_53(n32_1,n48_1);
nor I_54(n33_1,N1371_0_r_0,G78_5_r_0);
not I_55(n34_1,G42_7_r_0);
nor I_56(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_57(n36_1,n29_1);
not I_58(n37_1,n41_1);
nand I_59(n38_1,I_BUFF_1_9_r_1,N1508_0_r_0);
nand I_60(n39_1,n37_1,n40_1);
nand I_61(n40_1,n_429_or_0_5_r_0,n_549_7_r_0);
nand I_62(n41_1,n52_1,n_547_5_r_0);
or I_63(n42_1,n36_1,n43_1);
nor I_64(n43_1,n32_1,n49_1);
nand I_65(n44_1,n45_1,n46_1);
nand I_66(n45_1,n47_1,n48_1);
not I_67(n46_1,N1508_0_r_0);
not I_68(n47_1,n31_1);
nand I_69(n48_1,n50_1,n_576_5_r_0);
nor I_70(n49_1,n41_1,n47_1);
and I_71(n50_1,n51_1,G78_5_r_0);
nand I_72(n51_1,n52_1,n53_1);
nand I_73(n52_1,N1371_0_r_0,n_429_or_0_5_r_0);
not I_74(n53_1,n_547_5_r_0);
or I_75(n54_1,N1508_0_r_0,n_572_7_r_0);
nor I_76(n55_1,n29_1,N1508_0_r_0);
endmodule


