module test_I17611(I15897,I13908,I1477,I1470,I17611);
input I15897,I13908,I1477,I1470;
output I17611;
wire I13752,I15928,I13743,I15576,I15832,I14162,I16052,I15628,I13749,I15611,I16007,I17594,I15591,I16069;
DFFARX1 I_0(I1470,,,I13752,);
DFFARX1 I_1(I1470,I15611,,,I15928,);
nor I_2(I17611,I17594,I15591);
DFFARX1 I_3(I1470,,,I13743,);
DFFARX1 I_4(I16007,I1470,I15611,,,I15576,);
nand I_5(I15832,I15628,I13749);
DFFARX1 I_6(I1470,,,I14162,);
DFFARX1 I_7(I13752,I1470,I15611,,,I16052,);
not I_8(I15628,I13743);
nand I_9(I13749,I14162,I13908);
not I_10(I15611,I1477);
or I_11(I16007,I15928,I15897);
not I_12(I17594,I15576);
nor I_13(I15591,I16069,I15832);
not I_14(I16069,I16052);
endmodule


