module test_I5317(I1492,I3470,I1477,I1470,I3589,I1498,I5317);
input I1492,I3470,I1477,I1470,I3589,I1498;
output I5317;
wire I3374,I3388,I3702,I3747,I3620,I1483,I3668,I3365,I3877,I3685,I3356,I5283,I5300;
nand I_0(I3374,I3620,I3877);
not I_1(I3388,I1477);
DFFARX1 I_2(I3685,I1470,I3388,,,I3702,);
DFFARX1 I_3(I1470,I3388,,,I3747,);
nor I_4(I3620,I1492,I1483);
DFFARX1 I_5(I1470,,,I1483,);
DFFARX1 I_6(I1470,I3388,,,I3668,);
not I_7(I3365,I3702);
nor I_8(I3877,I3747,I3470);
and I_9(I5317,I5300,I3365);
and I_10(I3685,I3668,I1498);
DFFARX1 I_11(I3589,I1470,I3388,,,I3356,);
not I_12(I5283,I3356);
nor I_13(I5300,I5283,I3374);
endmodule


