module test_c6288_5_106(IN_1,IN_2,IN_3,N1371,N1372,N1508);
input IN_1,IN_2,IN_3;
output N1371,N1372,N1508;
wire N591,N1311;
and I_0(N591,IN_1,IN_2);
not I_1(N1311,N591);
nor I_2(N1371,N591,N1311);
not I_3(N1372,N1311);
nor I_4(N1508,N1311,IN_3);
endmodule


