module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2,n4_7_l_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
nor I_0(N1371_0_r_2,n32_2,n35_2);
nor I_1(N1508_0_r_2,n32_2,n55_2);
not I_2(N1372_1_r_2,n54_2);
nor I_3(N1508_1_r_2,n59_2,n54_2);
nor I_4(N6147_2_r_2,n42_2,n43_2);
nor I_5(N1507_6_r_2,n40_2,n53_2);
nor I_6(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_7(n4_7_r_2,blif_clk_net_7_r_4,n6_4,G42_7_r_2,);
nor I_8(n_572_7_r_2,n36_2,n37_2);
or I_9(n_573_7_r_2,n34_2,n35_2);
nor I_10(n_549_7_r_2,n40_2,n41_2);
nand I_11(n_569_7_r_2,n38_2,n39_2);
nor I_12(n_452_7_r_2,n59_2,n35_2);
nor I_13(n4_7_l_2,G18_7_l_2,IN_1_7_l_2);
DFFARX1 I_14(n4_7_l_2,blif_clk_net_7_r_4,n6_4,n59_2,);
not I_15(n33_2,n59_2);
and I_16(N3_8_l_2,IN_6_8_l_2,n49_2);
DFFARX1 I_17(N3_8_l_2,blif_clk_net_7_r_4,n6_4,n32_internal_2,);
not I_18(n32_2,n32_internal_2);
nor I_19(n4_7_r_2,n59_2,n36_2);
not I_20(n34_2,n39_2);
nor I_21(n35_2,IN_1_8_l_2,IN_3_8_l_2);
nor I_22(n36_2,G18_7_l_2,IN_5_7_l_2);
or I_23(n37_2,IN_9_7_l_2,IN_10_7_l_2);
not I_24(n38_2,n40_2);
nand I_25(n39_2,n45_2,n57_2);
nor I_26(n40_2,IN_3_1_l_2,n47_2);
nor I_27(n41_2,n32_2,n36_2);
not I_28(n42_2,n53_2);
nand I_29(n43_2,n44_2,n45_2);
nand I_30(n44_2,n38_2,n46_2);
not I_31(n45_2,IN_10_7_l_2);
nand I_32(n46_2,n47_2,n48_2);
nand I_33(n47_2,IN_1_1_l_2,IN_2_1_l_2);
or I_34(n48_2,G15_7_l_2,IN_7_7_l_2);
nand I_35(n49_2,IN_2_8_l_2,IN_3_8_l_2);
nand I_36(n50_2,n51_2,n52_2);
not I_37(n51_2,n47_2);
nand I_38(n52_2,n38_2,n53_2);
nor I_39(n53_2,IN_5_7_l_2,IN_9_7_l_2);
nand I_40(n54_2,n42_2,n56_2);
nor I_41(n55_2,n34_2,n56_2);
nor I_42(n56_2,G15_7_l_2,IN_7_7_l_2);
nand I_43(n57_2,IN_4_7_l_2,n58_2);
not I_44(n58_2,G15_7_l_2);
nor I_45(N1371_0_r_4,n25_4,N6147_2_r_2);
not I_46(N1508_0_r_4,n25_4);
nor I_47(N1507_6_r_4,n32_4,n33_4);
nor I_48(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_49(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_50(n_572_7_r_4,n_573_7_r_4);
nand I_51(n_573_7_r_4,n21_4,n22_4);
nor I_52(n_549_7_r_4,n24_4,N6147_2_r_2);
nand I_53(n_569_7_r_4,n22_4,n23_4);
nor I_54(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_55(N6147_9_r_4,n28_4);
nor I_56(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_57(I_BUFF_1_9_r_4,n21_4);
nor I_58(n4_7_r_4,N6147_9_r_4,N6147_2_r_2);
not I_59(n6_4,blif_reset_net_7_r_4);
nand I_60(n21_4,n39_4,n40_4);
or I_61(n22_4,n31_4,N1508_6_r_2);
not I_62(n23_4,N6147_2_r_2);
nor I_63(n24_4,n25_4,n26_4);
nand I_64(n25_4,N1371_0_r_2,N1508_0_r_2);
nand I_65(n26_4,n21_4,n27_4);
nand I_66(n27_4,n36_4,n37_4);
nand I_67(n28_4,n38_4,n_572_7_r_2);
nand I_68(n29_4,N1508_0_r_4,n30_4);
nand I_69(n30_4,n34_4,n35_4);
nor I_70(n31_4,N1372_1_r_2,n_569_7_r_2);
not I_71(n32_4,n30_4);
nor I_72(n33_4,n21_4,n28_4);
nand I_73(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_74(n35_4,N1508_0_r_4,n27_4);
not I_75(n36_4,n_549_7_r_2);
nand I_76(n37_4,n_573_7_r_2,N1371_0_r_2);
or I_77(n38_4,N1372_1_r_2,n_569_7_r_2);
nor I_78(n39_4,N1507_6_r_2,G42_7_r_2);
or I_79(n40_4,n41_4,N1508_1_r_2);
nor I_80(n41_4,N1508_0_r_2,n_452_7_r_2);
endmodule


