module test_I1639(I1255,I1294,I1207,I1301,I1639);
input I1255,I1294,I1207,I1301;
output I1639;
wire I1622,I1342;
DFFARX1 I_0(I1255,I1294,I1342,,,I1622,);
not I_1(I1342,I1301);
and I_2(I1639,I1622,I1207);
endmodule


