module test_I2393(I1477,I1470,I1375,I2393);
input I1477,I1470,I1375;
output I2393;
wire I2181,I2345;
not I_0(I2181,I1477);
DFFARX1 I_1(I1375,I1470,I2181,,,I2345,);
DFFARX1 I_2(I2345,I1470,I2181,,,I2393,);
endmodule


