module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7,n_452_7_r_7,n4_7_l_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N1371_0_r_7,n53_7,n52_7);
nor I_1(N1508_0_r_7,n51_7,n52_7);
nand I_2(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_3(n_431_5_r_7,blif_clk_net_7_r_12,n8_12,G78_5_r_7,);
nand I_4(n_576_5_r_7,n31_7,n32_7);
nor I_5(n_102_5_r_7,IN_5_7_l_7,IN_9_7_l_7);
nand I_6(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_7(n4_7_r_7,blif_clk_net_7_r_12,n8_12,G42_7_r_7,);
nor I_8(n_572_7_r_7,n54_7,n33_7);
nand I_9(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_10(n_549_7_r_7,n53_7,n36_7);
nand I_11(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_12(n_452_7_r_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_13(n4_7_l_7,G18_7_l_7,IN_1_7_l_7);
DFFARX1 I_14(n4_7_l_7,blif_clk_net_7_r_12,n8_12,n53_7,);
not I_15(n30_7,n53_7);
and I_16(N3_8_l_7,IN_6_8_l_7,n50_7);
DFFARX1 I_17(N3_8_l_7,blif_clk_net_7_r_12,n8_12,n54_7,);
nand I_18(n_431_5_r_7,n40_7,n41_7);
nor I_19(n4_7_r_7,n54_7,n49_7);
and I_20(n31_7,n_102_5_r_7,n39_7);
not I_21(n32_7,G18_7_l_7);
nor I_22(n33_7,IN_10_7_l_7,n34_7);
and I_23(n34_7,IN_4_7_l_7,n35_7);
not I_24(n35_7,G15_7_l_7);
nor I_25(n36_7,G18_7_l_7,n37_7);
or I_26(n37_7,IN_5_7_l_7,n54_7);
or I_27(n38_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_28(n39_7,IN_3_1_l_7,n_452_7_r_7);
nand I_29(n40_7,n46_7,n47_7);
nand I_30(n41_7,n42_7,n43_7);
nor I_31(n42_7,n44_7,n45_7);
nor I_32(n43_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_33(n44_7,G15_7_l_7,IN_7_7_l_7);
nor I_34(n45_7,IN_9_7_l_7,IN_10_7_l_7);
nand I_35(n46_7,IN_4_7_l_7,n35_7);
not I_36(n47_7,IN_10_7_l_7);
or I_37(n48_7,IN_3_1_l_7,n_452_7_r_7);
not I_38(n49_7,n_452_7_r_7);
nand I_39(n50_7,IN_2_8_l_7,IN_3_8_l_7);
and I_40(n51_7,n_452_7_r_7,n45_7);
not I_41(n52_7,n44_7);
nor I_42(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_43(N1508_0_r_12,n30_12,n37_12);
nor I_44(N1507_6_r_12,n25_12,n39_12);
nor I_45(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_46(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_47(n_572_7_r_12,n23_12,n24_12);
nand I_48(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_49(n_549_7_r_12,n27_12,n28_12);
nand I_50(n_569_7_r_12,n25_12,n26_12);
nand I_51(n_452_7_r_12,n_573_7_r_7,n_549_7_r_7);
nand I_52(N6147_9_r_12,n30_12,n31_12);
nor I_53(N6134_9_r_12,n35_12,n36_12);
not I_54(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_55(n1_12,n_573_7_r_12);
not I_56(n8_12,blif_reset_net_7_r_12);
not I_57(n23_12,n36_12);
nor I_58(n24_12,n_452_7_r_12,N1508_0_r_7);
nand I_59(n25_12,n23_12,n40_12);
not I_60(n26_12,n35_12);
not I_61(n27_12,N6134_9_r_12);
nand I_62(n28_12,n26_12,n29_12);
not I_63(n29_12,n24_12);
nand I_64(n30_12,n33_12,n41_12);
nand I_65(n31_12,n32_12,n33_12);
nor I_66(n32_12,n26_12,n34_12);
nor I_67(n33_12,n_429_or_0_5_r_7,N1371_0_r_7);
nor I_68(n34_12,n42_12,n_429_or_0_5_r_7);
nor I_69(n35_12,n38_12,G78_5_r_7);
nand I_70(n36_12,n_547_5_r_7,n_572_7_r_7);
nand I_71(n37_12,n23_12,n35_12);
or I_72(n38_12,n_576_5_r_7,G78_5_r_7);
not I_73(n39_12,n30_12);
or I_74(n40_12,N1371_0_r_7,N1508_0_r_7);
nor I_75(n41_12,n34_12,n36_12);
nor I_76(n42_12,G42_7_r_7,n_569_7_r_7);
endmodule


