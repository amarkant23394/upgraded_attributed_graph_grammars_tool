module test_I14404(I1477,I11395,I13231,I11429,I1470,I13409,I14404);
input I1477,I11395,I13231,I11429,I1470,I13409;
output I14404;
wire I13183,I13525,I13171,I13601,I13186,I13460,I14387,I13197,I11299,I13248,I13426,I11272,I13508,I13491;
nand I_0(I13183,I13601,I13525);
nor I_1(I13525,I13508,I13426);
nand I_2(I13171,I13248,I13460);
DFFARX1 I_3(I11299,I1470,I13197,,,I13601,);
nor I_4(I13186,I13601,I13508);
not I_5(I13460,I13426);
nand I_6(I14387,I13171,I13186);
not I_7(I13197,I1477);
nor I_8(I11299,I11395,I11429);
DFFARX1 I_9(I13231,I1470,I13197,,,I13248,);
DFFARX1 I_10(I13409,I1470,I13197,,,I13426,);
DFFARX1 I_11(I1470,,,I11272,);
and I_12(I14404,I14387,I13183);
and I_13(I13508,I13491,I11272);
DFFARX1 I_14(I1470,I13197,,,I13491,);
endmodule


