module test_I12670(I10797,I1477,I1470,I11201,I12670);
input I10797,I1477,I1470,I11201;
output I12670;
wire I12619,I10612,I11009,I10647,I11167,I11057,I10627,I10639,I11150,I12636,I12653;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
DFFARX1 I_2(I11009,I1470,I10647,,,I10612,);
DFFARX1 I_3(I1470,I10647,,,I11009,);
not I_4(I10647,I1477);
not I_5(I11167,I11150);
nor I_6(I11057,I11009,I10797);
nand I_7(I10627,I11167,I11057);
DFFARX1 I_8(I11201,I1470,I10647,,,I10639,);
DFFARX1 I_9(I1470,I10647,,,I11150,);
nand I_10(I12636,I10612,I10639);
and I_11(I12653,I12636,I10627);
endmodule


