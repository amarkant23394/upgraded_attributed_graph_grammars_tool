module test_I9465(I8267,I1477,I8360,I8496,I1470,I8315,I9465);
input I8267,I1477,I8360,I8496,I1470,I8315;
output I9465;
wire I9576,I8202,I8181,I9638,I8216,I8623,I9816,I8705,I8592,I8205,I9621,I8193,I9491;
nor I_0(I9576,I8181,I8202);
nand I_1(I8202,I8267,I8496);
and I_2(I8181,I8360,I8592);
nand I_3(I9465,I9816,I9638);
nor I_4(I9638,I9621,I9576);
not I_5(I8216,I1477);
DFFARX1 I_6(I1470,I8216,,,I8623,);
DFFARX1 I_7(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_8(I8623,I1470,I8216,,,I8705,);
DFFARX1 I_9(I1470,I8216,,,I8592,);
not I_10(I8205,I8315);
DFFARX1 I_11(I8205,I1470,I9491,,,I9621,);
not I_12(I8193,I8705);
not I_13(I9491,I1477);
endmodule


