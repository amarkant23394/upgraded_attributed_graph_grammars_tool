module test_I5768(I4544,I2328,I2181,I2170,I2557,I2509,I1470,I5768);
input I4544,I2328,I2181,I2170,I2557,I2509,I1470;
output I5768;
wire I2167,I4629,I4595,I4869,I2149,I2633,I2143,I4886,I4530,I4807,I2173,I4515,I4824,I4612;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
DFFARX1 I_2(I1470,I4544,,,I4595,);
DFFARX1 I_3(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_4(I1470,I2181,,,I2149,);
DFFARX1 I_5(I1470,I2181,,,I2633,);
DFFARX1 I_6(I2557,I1470,I2181,,,I2143,);
and I_7(I4886,I4869,I4612);
nand I_8(I5768,I4530,I4515);
nor I_9(I4530,I4824,I4886);
DFFARX1 I_10(I2170,I1470,I4544,,,I4807,);
nand I_11(I2173,I2557,I2509);
not I_12(I4515,I4629);
and I_13(I4824,I4807,I2143);
not I_14(I4612,I4595);
endmodule


