module test_final(IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_6,blif_reset_net_5_r_6,N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,G78_5_r_6,n_576_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_6,blif_reset_net_5_r_6;
output N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,G78_5_r_6,n_576_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_102_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4,n_431_5_r_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n_429_or_0_5_r_6,n_102_5_r_6,n_431_5_r_6,n6_6,n24_6,n25_6,n26_6,n27_6,n28_6,n29_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6;
nor I_0(N1371_0_r_4,n25_4,n29_4);
nor I_1(N1508_0_r_4,n25_4,n32_4);
nor I_2(N6147_2_r_4,n24_4,n31_4);
or I_3(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_4(n_431_5_r_4,blif_clk_net_5_r_6,n6_6,G78_5_r_4,);
nand I_5(n_576_5_r_4,n22_4,n23_4);
nand I_6(n_102_5_r_4,n34_4,n35_4);
nand I_7(n_547_5_r_4,n26_4,n27_4);
nor I_8(N1507_6_r_4,n27_4,n30_4);
nor I_9(N1508_6_r_4,n30_4,n33_4);
nand I_10(n_431_5_r_4,n_102_5_r_4,n28_4);
nor I_11(n22_4,n24_4,n25_4);
nor I_12(n23_4,IN_1_3_l_4,n37_4);
not I_13(n24_4,n_102_5_r_4);
nand I_14(n25_4,IN_1_1_l_4,IN_2_1_l_4);
nor I_15(n26_4,n23_4,n24_4);
not I_16(n27_4,n25_4);
nand I_17(n28_4,n23_4,n29_4);
nor I_18(n29_4,IN_3_1_l_4,n25_4);
not I_19(n30_4,n29_4);
nor I_20(n31_4,N1371_0_r_4,n32_4);
nor I_21(n32_4,n23_4,n29_4);
nand I_22(n33_4,n23_4,n24_4);
nor I_23(n34_4,IN_1_2_l_4,IN_2_2_l_4);
or I_24(n35_4,IN_5_2_l_4,n36_4);
nor I_25(n36_4,IN_3_2_l_4,IN_4_2_l_4);
or I_26(n37_4,IN_2_3_l_4,IN_3_3_l_4);
nor I_27(N1371_0_r_6,n26_6,n38_6);
not I_28(N1508_0_r_6,n38_6);
nor I_29(N6147_3_r_6,n30_6,n35_6);
nand I_30(n_429_or_0_5_r_6,n30_6,n32_6);
DFFARX1 I_31(n_431_5_r_6,blif_clk_net_5_r_6,n6_6,G78_5_r_6,);
nand I_32(n_576_5_r_6,n24_6,n25_6);
not I_33(n_102_5_r_6,n26_6);
or I_34(n_547_5_r_6,n_429_or_0_5_r_6,n26_6);
not I_35(N1372_10_r_6,n37_6);
nor I_36(N1508_10_r_6,n36_6,n37_6);
nand I_37(n_431_5_r_6,n_102_5_r_6,n28_6);
not I_38(n6_6,blif_reset_net_5_r_6);
nor I_39(n24_6,n33_6,n34_6);
nor I_40(n25_6,n26_6,n27_6);
nor I_41(n26_6,n40_6,N6147_2_r_4);
nand I_42(n27_6,n_576_5_r_4,N1508_0_r_4);
nand I_43(n28_6,n29_6,n30_6);
nor I_44(n29_6,n31_6,N1508_0_r_4);
not I_45(n30_6,n27_6);
nor I_46(n31_6,n39_6,n40_6);
nor I_47(n32_6,n24_6,N1508_0_r_4);
not I_48(n33_6,N1508_6_r_4);
not I_49(n34_6,n_429_or_0_5_r_4);
or I_50(n35_6,n26_6,n31_6);
and I_51(n36_6,n38_6,N1508_0_r_4);
nand I_52(n37_6,n30_6,n31_6);
nand I_53(n38_6,n41_6,n_429_or_0_5_r_4);
nor I_54(n39_6,n_547_5_r_4,N1507_6_r_4);
not I_55(n40_6,G78_5_r_4);
nor I_56(n41_6,n33_6,n42_6);
nor I_57(n42_6,N6147_2_r_4,n_429_or_0_5_r_4);
endmodule


