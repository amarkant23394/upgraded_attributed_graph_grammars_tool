module test_I16486(I14350,I16257,I1477,I1470,I14825,I14359,I16486);
input I14350,I16257,I1477,I1470,I14825,I14359;
output I16486;
wire I16308,I14362,I16452,I16291,I16469,I16240,I16274,I16435,I14370,I14332;
not I_0(I16308,I16291);
DFFARX1 I_1(I14825,I1470,I14370,,,I14362,);
and I_2(I16452,I16435,I14362);
DFFARX1 I_3(I16274,I1470,I16240,,,I16291,);
nor I_4(I16486,I16469,I16308);
DFFARX1 I_5(I16452,I1470,I16240,,,I16469,);
not I_6(I16240,I1477);
and I_7(I16274,I16257,I14332);
nand I_8(I16435,I14359,I14350);
not I_9(I14370,I1477);
DFFARX1 I_10(I1470,I14370,,,I14332,);
endmodule


