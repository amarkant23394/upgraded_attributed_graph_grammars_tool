module test_I8205(I6265,I5751,I5785,I1470,I8205);
input I6265,I5751,I5785,I1470;
output I8205;
wire I8233,I5802,I8298,I5719,I5740,I8315,I5722;
not I_0(I8205,I8315);
not I_1(I8233,I5722);
DFFARX1 I_2(I5785,I1470,I5751,,,I5802,);
nor I_3(I8298,I8233,I5719);
DFFARX1 I_4(I6265,I1470,I5751,,,I5719,);
not I_5(I5740,I5802);
nand I_6(I8315,I8298,I5740);
DFFARX1 I_7(I1470,I5751,,,I5722,);
endmodule


