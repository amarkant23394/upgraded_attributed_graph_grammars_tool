module test_I7286(I1477,I5204,I1470,I5249,I7286);
input I1477,I5204,I1470,I5249;
output I7286;
wire I5105,I5351,I5073,I6992,I6975,I5625,I5368,I5070,I5067,I6907,I5481,I7269,I5097,I5642,I6924;
not I_0(I5105,I1477);
DFFARX1 I_1(I1470,I5105,,,I5351,);
DFFARX1 I_2(I1470,I5105,,,I5073,);
nand I_3(I6992,I6975,I5097);
nor I_4(I6975,I6924,I5070);
DFFARX1 I_5(I1470,I5105,,,I5625,);
nor I_6(I5368,I5351,I5204);
and I_7(I5070,I5249,I5481);
DFFARX1 I_8(I5642,I1470,I5105,,,I5067,);
not I_9(I6907,I1477);
DFFARX1 I_10(I1470,I5105,,,I5481,);
DFFARX1 I_11(I5067,I1470,I6907,,,I7269,);
nand I_12(I5097,I5642,I5368);
nor I_13(I7286,I7269,I6992);
not I_14(I5642,I5625);
not I_15(I6924,I5073);
endmodule


