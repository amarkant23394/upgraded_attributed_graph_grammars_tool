module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_7_r_5,n7_5,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_5,n28_5,n46_5);
nand I_40(N1508_0_r_5,n26_5,n43_5);
not I_41(N1372_1_r_5,n43_5);
nor I_42(N1508_1_r_5,n30_5,n43_5);
nor I_43(N6147_2_r_5,n29_5,n32_5);
nor I_44(N1507_6_r_5,n26_5,n44_5);
nor I_45(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_46(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_47(n_572_7_r_5,n27_5,n28_5);
nand I_48(n_573_7_r_5,n26_5,n27_5);
nand I_49(n_549_7_r_5,N1508_6_r_15,n_429_or_0_5_r_15);
nand I_50(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_51(n_452_7_r_5,n29_5);
nor I_52(n4_7_r_5,n30_5,n31_5);
not I_53(n7_5,blif_reset_net_7_r_5);
not I_54(n26_5,n35_5);
nand I_55(n27_5,n40_5,n41_5);
nand I_56(n28_5,n_429_or_0_5_r_15,n_547_5_r_15);
nand I_57(n29_5,n27_5,n33_5);
nor I_58(n30_5,n45_5,N1508_1_r_15);
not I_59(n31_5,n_549_7_r_5);
nor I_60(n32_5,n34_5,n35_5);
not I_61(n33_5,n30_5);
nor I_62(n34_5,n31_5,n36_5);
nor I_63(n35_5,n28_5,G78_5_r_15);
not I_64(n36_5,n28_5);
nand I_65(n37_5,n36_5,n38_5);
nand I_66(n38_5,n26_5,n39_5);
nand I_67(n39_5,n30_5,n31_5);
nor I_68(n40_5,N1372_4_r_15,G78_5_r_15);
or I_69(n41_5,n42_5,N1508_1_r_15);
nor I_70(n42_5,N1372_4_r_15,n_576_5_r_15);
nand I_71(n43_5,n36_5,n46_5);
nor I_72(n44_5,n_549_7_r_5,n33_5);
or I_73(n45_5,N1507_6_r_15,N1508_4_r_15);
and I_74(n46_5,n31_5,n47_5);
or I_75(n47_5,N1508_4_r_15,n_576_5_r_15);
endmodule


