module test_final(G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8,n_431_0_l_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_8,blif_clk_net_1_r_15,n4_15,G42_1_r_8,);
nor I_1(n_572_1_r_8,n39_8,n23_8);
and I_2(n_549_1_r_8,n38_8,n23_8);
nand I_3(n_569_1_r_8,n38_8,n24_8);
nor I_4(n_452_1_r_8,n25_8,n26_8);
nor I_5(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_6(N3_2_r_8,blif_clk_net_1_r_15,n4_15,G199_2_r_8,);
DFFARX1 I_7(N1_4_r_8,blif_clk_net_1_r_15,n4_15,G199_4_r_8,);
DFFARX1 I_8(G78_0_l_8,blif_clk_net_1_r_15,n4_15,G214_4_r_8,);
or I_9(n_431_0_l_8,IN_8_0_l_8,n29_8);
DFFARX1 I_10(n_431_0_l_8,blif_clk_net_1_r_15,n4_15,G78_0_l_8,);
not I_11(n19_8,G78_0_l_8);
DFFARX1 I_12(IN_2_5_l_8,blif_clk_net_1_r_15,n4_15,n39_8,);
not I_13(n22_8,n39_8);
DFFARX1 I_14(IN_1_5_l_8,blif_clk_net_1_r_15,n4_15,n38_8,);
nor I_15(n4_1_r_8,G78_0_l_8,n33_8);
nor I_16(N3_2_r_8,n22_8,n35_8);
nor I_17(N1_4_r_8,n27_8,n37_8);
nand I_18(n23_8,IN_7_0_l_8,n32_8);
not I_19(n24_8,n23_8);
nand I_20(n25_8,IN_11_0_l_8,n36_8);
nand I_21(n26_8,n27_8,n28_8);
nor I_22(n27_8,IN_5_0_l_8,n31_8);
not I_23(n28_8,G2_0_l_8);
and I_24(n29_8,IN_2_0_l_8,n30_8);
nor I_25(n30_8,IN_4_0_l_8,n31_8);
not I_26(n31_8,G1_0_l_8);
and I_27(n32_8,IN_5_0_l_8,n28_8);
nand I_28(n33_8,n28_8,n34_8);
not I_29(n34_8,n25_8);
nor I_30(n35_8,G2_0_l_8,n34_8);
not I_31(n36_8,IN_10_0_l_8);
nor I_32(n37_8,n19_8,n38_8);
DFFARX1 I_33(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_34(n_572_1_r_15,n17_15,n19_15);
nand I_35(n_573_1_r_15,n15_15,n18_15);
nor I_36(n_549_1_r_15,n21_15,n22_15);
nand I_37(n_569_1_r_15,n15_15,n20_15);
nor I_38(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_39(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_40(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_41(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_42(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_43(n4_1_l_15,n_452_1_r_8,n_42_2_r_8);
not I_44(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_45(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_46(n15_15,G42_1_l_15);
DFFARX1 I_47(G42_1_r_8,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_48(n17_15,n17_internal_15);
DFFARX1 I_49(n_572_1_r_8,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_50(n_572_1_l_15,n_549_1_r_8,G199_4_r_8);
DFFARX1 I_51(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_52(n14_15,n14_internal_15);
nand I_53(N1_4_r_15,n25_15,n26_15);
or I_54(n_573_1_l_15,n_572_1_r_8,G42_1_r_8);
nor I_55(n18_15,n_572_1_r_8,n_569_1_r_8);
nand I_56(n19_15,n27_15,n28_15);
nand I_57(n20_15,n30_15,G199_2_r_8);
not I_58(n21_15,n20_15);
and I_59(n22_15,n17_15,n_572_1_l_15);
nor I_60(n23_15,n_452_1_r_8,G42_1_r_8);
or I_61(n24_15,n_572_1_r_8,n_569_1_r_8);
or I_62(n25_15,n_573_1_l_15,n_452_1_r_8);
nand I_63(n26_15,n19_15,n23_15);
not I_64(n27_15,n_569_1_r_8);
nand I_65(n28_15,n29_15,G214_4_r_8);
not I_66(n29_15,G199_4_r_8);
endmodule


