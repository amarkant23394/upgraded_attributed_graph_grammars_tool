module test_I8770(I1477,I6127,I6079,I1470,I5881,I8298,I5740,I8770);
input I1477,I6127,I6079,I1470,I5881,I8298,I5740;
output I8770;
wire I8674,I8640,I8216,I8753,I8623,I5743,I8657,I5915,I5731,I8315,I8736;
or I_0(I8770,I8753,I8674);
and I_1(I8674,I8623,I8657);
not I_2(I8640,I8623);
not I_3(I8216,I1477);
not I_4(I8753,I8736);
DFFARX1 I_5(I5743,I1470,I8216,,,I8623,);
nand I_6(I5743,I6127,I6079);
nor I_7(I8657,I8315,I8640);
DFFARX1 I_8(I1470,,,I5915,);
nand I_9(I5731,I5915,I5881);
nand I_10(I8315,I8298,I5740);
DFFARX1 I_11(I5731,I1470,I8216,,,I8736,);
endmodule


