module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_14,blif_reset_net_7_r_14,N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_7_r_14,blif_reset_net_7_r_14;
output N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,I_BUFF_1_9_r_14,N3_8_l_14,n8_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_7_r_14,n8_14,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_14,n47_14,n30_14);
nor I_40(N1508_0_r_14,n30_14,n41_14);
nor I_41(N1507_6_r_14,n37_14,n44_14);
nor I_42(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_43(n4_7_r_14,blif_clk_net_7_r_14,n8_14,G42_7_r_14,);
nor I_44(n_572_7_r_14,n28_14,n29_14);
nand I_45(n_573_7_r_14,n26_14,n27_14);
nor I_46(n_549_7_r_14,n31_14,n32_14);
nand I_47(n_569_7_r_14,n26_14,n30_14);
nor I_48(n_452_7_r_14,n47_14,n28_14);
nor I_49(N6147_9_r_14,n36_14,n37_14);
nor I_50(N6134_9_r_14,n28_14,n36_14);
not I_51(I_BUFF_1_9_r_14,n26_14);
and I_52(N3_8_l_14,n38_14,N1372_4_r_15);
not I_53(n8_14,blif_reset_net_7_r_14);
DFFARX1 I_54(N3_8_l_14,blif_clk_net_7_r_14,n8_14,n47_14,);
nor I_55(n4_7_r_14,n47_14,n35_14);
nand I_56(n26_14,n_576_5_r_15,n_547_5_r_15);
not I_57(n27_14,n28_14);
nor I_58(n28_14,n43_14,G78_5_r_15);
not I_59(n29_14,n33_14);
not I_60(n30_14,n31_14);
nor I_61(n31_14,n46_14,N1372_4_r_15);
and I_62(n32_14,n33_14,n34_14);
nand I_63(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_64(n34_14,n42_14,n43_14);
nor I_65(n35_14,N1508_1_r_15,G78_5_r_15);
nor I_66(n36_14,n47_14,n34_14);
not I_67(n37_14,n35_14);
nand I_68(n38_14,N1508_4_r_15,G78_5_r_15);
nand I_69(n39_14,n29_14,n40_14);
nand I_70(n40_14,n27_14,n37_14);
nor I_71(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_72(n42_14,N1507_6_r_15,n_576_5_r_15);
not I_73(n43_14,N1508_6_r_15);
nor I_74(n44_14,n27_14,n33_14);
or I_75(n45_14,N1508_4_r_15,n_429_or_0_5_r_15);
or I_76(n46_14,N1508_1_r_15,n_429_or_0_5_r_15);
endmodule


