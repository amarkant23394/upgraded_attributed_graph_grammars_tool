module test_I10732(I8202,I1477,I8181,I8205,I1470,I10732);
input I8202,I1477,I8181,I8205,I1470;
output I10732;
wire I10664,I9559,I9471,I10715,I9542,I9638,I9816,I9771,I8178,I8193,I9491,I9477,I9754,I8705,I9833,I9576,I9465,I9621,I9689;
not I_0(I10664,I9471);
not I_1(I9559,I9542);
nor I_2(I9471,I9689,I9542);
nor I_3(I10715,I10664,I9477);
DFFARX1 I_4(I1470,I9491,,,I9542,);
nor I_5(I9638,I9621,I9576);
DFFARX1 I_6(I8193,I1470,I9491,,,I9816,);
and I_7(I9771,I9754,I8178);
DFFARX1 I_8(I1470,,,I8178,);
nand I_9(I10732,I10715,I9465);
not I_10(I8193,I8705);
not I_11(I9491,I1477);
nor I_12(I9477,I9771,I9833);
DFFARX1 I_13(I1470,I9491,,,I9754,);
DFFARX1 I_14(I1470,,,I8705,);
and I_15(I9833,I9816,I9559);
nor I_16(I9576,I8181,I8202);
nand I_17(I9465,I9816,I9638);
DFFARX1 I_18(I8205,I1470,I9491,,,I9621,);
DFFARX1 I_19(I1470,I9491,,,I9689,);
endmodule


