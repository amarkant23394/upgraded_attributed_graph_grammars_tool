module test_I15485(I12831,I1477,I10766,I1470,I10732,I15485);
input I12831,I1477,I10766,I1470,I10732;
output I15485;
wire I12619,I12913,I13023,I12930,I12605,I12947,I10636,I14965,I12848,I10609;
not I_0(I12619,I1477);
DFFARX1 I_1(I1470,I12619,,,I12913,);
DFFARX1 I_2(I10636,I1470,I12619,,,I13023,);
and I_3(I12930,I12913,I10609);
nand I_4(I12605,I13023,I12947);
nor I_5(I12947,I12930,I12848);
nor I_6(I10636,I10732,I10766);
not I_7(I14965,I1477);
DFFARX1 I_8(I12831,I1470,I12619,,,I12848,);
DFFARX1 I_9(I12605,I1470,I14965,,,I15485,);
DFFARX1 I_10(I1470,,,I10609,);
endmodule


