module test_I5079(I3798,I1477,I3521,I3405,I1470,I5079);
input I3798,I1477,I3521,I3405,I1470;
output I5079;
wire I5156,I3388,I3359,I3371,I5139,I3380,I3846,I3815,I3747,I5105;
nand I_0(I5156,I5139,I3371);
not I_1(I3388,I1477);
DFFARX1 I_2(I3747,I1470,I3388,,,I3359,);
DFFARX1 I_3(I3815,I1470,I3388,,,I3371,);
nor I_4(I5139,I3380,I3359);
nand I_5(I3380,I3521,I3846);
nor I_6(I3846,I3747);
or I_7(I3815,I3405,I3798);
DFFARX1 I_8(I5156,I1470,I5105,,,I5079,);
DFFARX1 I_9(I1470,I3388,,,I3747,);
not I_10(I5105,I1477);
endmodule


