module test_I9480(I8527,I1477,I8315,I5737,I1470,I9480);
input I8527,I1477,I8315,I5737,I1470;
output I9480;
wire I8202,I8753,I8496,I8216,I9771,I8178,I5719,I8377,I8250,I9491,I8181,I8360,I9754,I8592,I8736,I8462,I8187,I9576,I8267;
nand I_0(I8202,I8267,I8496);
not I_1(I8753,I8736);
nor I_2(I8496,I8462,I8377);
not I_3(I8216,I1477);
or I_4(I9480,I9771,I9576);
and I_5(I9771,I9754,I8178);
DFFARX1 I_6(I8753,I1470,I8216,,,I8178,);
DFFARX1 I_7(I1470,,,I5719,);
not I_8(I8377,I8360);
nor I_9(I8250,I5719);
not I_10(I9491,I1477);
and I_11(I8181,I8360,I8592);
not I_12(I8360,I5719);
DFFARX1 I_13(I8187,I1470,I9491,,,I9754,);
DFFARX1 I_14(I8527,I1470,I8216,,,I8592,);
DFFARX1 I_15(I1470,I8216,,,I8736,);
DFFARX1 I_16(I1470,I8216,,,I8462,);
DFFARX1 I_17(I8315,I1470,I8216,,,I8187,);
nor I_18(I9576,I8181,I8202);
nand I_19(I8267,I8250,I5737);
endmodule


