module test_I13755(I1477,I12058,I12380,I11944,I12304,I1470,I13755);
input I1477,I12058,I12380,I11944,I12304,I1470;
output I13755;
wire I11935,I13908,I14004,I13891,I11941,I12208,I13987,I13775,I13843,I11965,I11950,I11973,I13970,I11959,I13925;
DFFARX1 I_0(I12208,I1470,I11973,,,I11935,);
not I_1(I13908,I13891);
DFFARX1 I_2(I13987,I1470,I13775,,,I14004,);
DFFARX1 I_3(I11944,I1470,I13775,,,I13891,);
DFFARX1 I_4(I12208,I1470,I11973,,,I11941,);
DFFARX1 I_5(I1470,I11973,,,I12208,);
and I_6(I13987,I13970,I11941);
not I_7(I13775,I1477);
nor I_8(I13843,I11959,I11965);
DFFARX1 I_9(I12304,I1470,I11973,,,I11965,);
nand I_10(I13755,I14004,I13925);
DFFARX1 I_11(I1470,I11973,,,I11950,);
not I_12(I11973,I1477);
nand I_13(I13970,I11935,I11950);
nand I_14(I11959,I12058,I12380);
nor I_15(I13925,I13843,I13908);
endmodule


