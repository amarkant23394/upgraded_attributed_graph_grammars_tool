module test_I3379(I2234,I1294,I1301,I3379);
input I2234,I1294,I1301;
output I3379;
wire I2548,I2583,I1902,I2203,I2945;
not I_0(I3379,I2548);
DFFARX1 I_1(I2945,I1294,I2583,,,I2548,);
not I_2(I2583,I1301);
and I_3(I1902,I2234,I2203);
DFFARX1 I_4(I1294,,,I2203,);
DFFARX1 I_5(I1902,I1294,I2583,,,I2945,);
endmodule


