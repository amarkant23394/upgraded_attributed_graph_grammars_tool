module test_I6781(I2810,I2742,I3124,I1477,I1470,I2751,I6781);
input I2810,I2742,I3124,I1477,I1470,I2751;
output I6781;
wire I2727,I6329,I4113,I4308,I4068,I4130,I3957,I2724,I3983;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
nand I_1(I2727,I2810,I3124);
not I_2(I6329,I1477);
DFFARX1 I_3(I2751,I1470,I3983,,,I4113,);
DFFARX1 I_4(I2727,I1470,I3983,,,I4308,);
nor I_5(I4068,I2742,I2724);
nor I_6(I4130,I4113,I4068);
nand I_7(I3957,I4308,I4130);
DFFARX1 I_8(I1470,,,I2724,);
not I_9(I3983,I1477);
endmodule


