module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_2,blif_reset_net_1_r_2,G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_2,blif_reset_net_1_r_2;
output G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_573_1_r_2,N3_2_l_2,n5_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_2,n5_2,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_2,n5_2,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_2,n5_2,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_2,n5_2,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_2,blif_clk_net_1_r_2,n5_2,G42_1_r_2,);
nor I_32(n_572_1_r_2,n26_2,n18_2);
nand I_33(n_573_1_r_2,n17_2,n19_2);
nor I_34(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_35(n_569_1_r_2,n13_2,n19_2);
not I_36(n_452_1_r_2,n_573_1_r_2);
nor I_37(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_38(N3_2_r_2,blif_clk_net_1_r_2,n5_2,G199_2_r_2,);
DFFARX1 I_39(ACVQN2_3_l_2,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_2,);
not I_40(P6_5_r_2,P6_5_r_internal_2);
and I_41(N3_2_l_2,n24_2,n_569_1_r_14);
not I_42(n5_2,blif_reset_net_1_r_2);
DFFARX1 I_43(N3_2_l_2,blif_clk_net_1_r_2,n5_2,G199_2_l_2,);
not I_44(n13_2,G199_2_l_2);
DFFARX1 I_45(G42_1_r_14,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_2,);
DFFARX1 I_46(P6_5_r_14,blif_clk_net_1_r_2,n5_2,n16_2,);
and I_47(N1_4_l_2,n25_2,G199_2_r_14);
DFFARX1 I_48(N1_4_l_2,blif_clk_net_1_r_2,n5_2,n26_2,);
DFFARX1 I_49(G42_1_r_14,blif_clk_net_1_r_2,n5_2,n17_internal_2,);
not I_50(n17_2,n17_internal_2);
nor I_51(n4_1_r_2,n26_2,n22_2);
nor I_52(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_53(G199_2_l_2,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_2,);
nor I_54(n18_2,n_573_1_r_14,ACVQN1_5_r_14);
nand I_55(n19_2,n16_2,n_572_1_r_14);
nor I_56(n20_2,n26_2,n21_2);
not I_57(n21_2,n18_2);
and I_58(n22_2,n16_2,n_572_1_r_14);
nor I_59(n23_2,n13_2,n21_2);
nand I_60(n24_2,n_42_2_r_14,ACVQN1_5_r_14);
nand I_61(n25_2,n_572_1_r_14,n_549_1_r_14);
endmodule


