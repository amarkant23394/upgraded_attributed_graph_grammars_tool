module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_7_r_12,n8_12,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
nor I_39(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_40(N1508_0_r_12,n30_12,n37_12);
nor I_41(N1507_6_r_12,n25_12,n39_12);
nor I_42(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_43(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_44(n_572_7_r_12,n23_12,n24_12);
nand I_45(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_46(n_549_7_r_12,n27_12,n28_12);
nand I_47(n_569_7_r_12,n25_12,n26_12);
nand I_48(n_452_7_r_12,N1508_10_r_6,N1508_0_r_6);
nand I_49(N6147_9_r_12,n30_12,n31_12);
nor I_50(N6134_9_r_12,n35_12,n36_12);
not I_51(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_52(n1_12,n_573_7_r_12);
not I_53(n8_12,blif_reset_net_7_r_12);
not I_54(n23_12,n36_12);
nor I_55(n24_12,n_452_7_r_12,N1372_1_r_6);
nand I_56(n25_12,n23_12,n40_12);
not I_57(n26_12,n35_12);
not I_58(n27_12,N6134_9_r_12);
nand I_59(n28_12,n26_12,n29_12);
not I_60(n29_12,n24_12);
nand I_61(n30_12,n33_12,n41_12);
nand I_62(n31_12,n32_12,n33_12);
nor I_63(n32_12,n26_12,n34_12);
nor I_64(n33_12,N1508_1_r_6,N6134_9_r_6);
nor I_65(n34_12,n42_12,N1508_0_r_6);
nor I_66(n35_12,n38_12,N1507_6_r_6);
nand I_67(n36_12,N6147_9_r_6,N1372_1_r_6);
nand I_68(n37_12,n23_12,n35_12);
or I_69(n38_12,N1371_0_r_6,N1508_6_r_6);
not I_70(n39_12,n30_12);
or I_71(n40_12,G199_8_r_6,N1371_0_r_6);
nor I_72(n41_12,n34_12,n36_12);
nor I_73(n42_12,n_42_8_r_6,N1372_10_r_6);
endmodule


