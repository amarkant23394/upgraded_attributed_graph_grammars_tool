module test_I11508(I9148,I6992,I1477,I7057,I1470,I6887,I11508);
input I9148,I6992,I1477,I7057,I1470,I6887;
output I11508;
wire I9320,I11491,I6875,I8827,I8842,I9303,I8862,I6881,I8879,I9258,I9179,I9083;
not I_0(I9320,I9303);
not I_1(I11491,I8827);
DFFARX1 I_2(I1470,,,I6875,);
nor I_3(I11508,I11491,I8842);
DFFARX1 I_4(I9258,I1470,I8862,,,I8827,);
nor I_5(I8842,I9320,I9083);
DFFARX1 I_6(I6875,I1470,I8862,,,I9303,);
not I_7(I8862,I1477);
nand I_8(I6881,I6992,I7057);
not I_9(I8879,I6887);
or I_10(I9258,I9179,I9148);
DFFARX1 I_11(I1470,I8862,,,I9179,);
nand I_12(I9083,I8879,I6881);
endmodule


