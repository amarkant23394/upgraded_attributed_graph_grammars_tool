module test_I12913(I9462,I9465,I9864,I10715,I10862,I1470_clk,I1477_rst,I12913);
input I9462,I9465,I9864,I10715,I10862,I1470_clk,I1477_rst;
output I12913;
wire I10879,I12619_rst,I10732,I11009,I10647,I11026,I10633,I9468,I10896,I9491_rst;
or I_0(I10879,I10862,I9462);
not I_1(I12619_rst,I1477_rst);
nand I_2(I10732,I10715,I9465);
DFFARX1 I_3 (I9468,I10647,I1470_clk,);
not I_4(I10647,I1477_rst);
nor I_5(I11026,I11009,I10732);
nand I_6(I10633,I10896,I11026);
DFFARX1 I_7 (I9864,I1470_clk,I9491_rst,I9468);
DFFARX1 I_8 (I10879,I10647,I1470_clk,);
not I_9(I9491_rst,I1477_rst);
DFFARX1 I_10 (I10633,I1470_clk,I12619_rst,I12913);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule