module test_final(IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_5,blif_reset_net_1_r_5,G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5);
input IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_5,blif_reset_net_1_r_5;
output G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5;
wire G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1,N3_2_l_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1,N3_2_l_5,n5_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5;
DFFARX1 I_0(n4_1_r_1,blif_clk_net_1_r_5,n5_5,G42_1_r_1,);
nor I_1(n_572_1_r_1,n26_1,n19_1);
nand I_2(n_573_1_r_1,n16_1,n18_1);
nor I_3(n_549_1_r_1,n20_1,n21_1);
nor I_4(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_5(G199_4_l_1,blif_clk_net_1_r_5,n5_5,ACVQN2_3_r_1,);
nor I_6(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_7(N1_4_r_1,blif_clk_net_1_r_5,n5_5,G199_4_r_1,);
DFFARX1 I_8(G199_4_l_1,blif_clk_net_1_r_5,n5_5,G214_4_r_1,);
and I_9(N3_2_l_1,IN_6_2_l_1,n23_1);
DFFARX1 I_10(N3_2_l_1,blif_clk_net_1_r_5,n5_5,n26_1,);
not I_11(n17_1,n26_1);
DFFARX1 I_12(IN_1_3_l_1,blif_clk_net_1_r_5,n5_5,n16_internal_1,);
not I_13(n16_1,n16_internal_1);
DFFARX1 I_14(IN_2_3_l_1,blif_clk_net_1_r_5,n5_5,ACVQN1_3_l_1,);
and I_15(N1_4_l_1,IN_6_4_l_1,n25_1);
DFFARX1 I_16(N1_4_l_1,blif_clk_net_1_r_5,n5_5,G199_4_l_1,);
DFFARX1 I_17(IN_3_4_l_1,blif_clk_net_1_r_5,n5_5,G214_4_l_1,);
nor I_18(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_19(G214_4_l_1,blif_clk_net_1_r_5,n5_5,n14_internal_1,);
not I_20(n14_1,n14_internal_1);
nor I_21(N1_4_r_1,n17_1,n24_1);
nand I_22(n18_1,IN_4_3_l_1,ACVQN1_3_l_1);
nor I_23(n19_1,IN_1_2_l_1,IN_3_2_l_1);
not I_24(n20_1,n18_1);
nor I_25(n21_1,n26_1,n22_1);
not I_26(n22_1,n19_1);
nand I_27(n23_1,IN_2_2_l_1,IN_3_2_l_1);
nor I_28(n24_1,n18_1,n22_1);
nand I_29(n25_1,IN_1_4_l_1,IN_2_4_l_1);
DFFARX1 I_30(n4_1_r_5,blif_clk_net_1_r_5,n5_5,G42_1_r_5,);
nor I_31(n_572_1_r_5,n21_5,n22_5);
nand I_32(n_573_1_r_5,n13_5,n16_5);
nor I_33(n_549_1_r_5,n21_5,n17_5);
nand I_34(n_569_1_r_5,n13_5,n15_5);
nor I_35(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_36(G199_2_l_5,blif_clk_net_1_r_5,n5_5,ACVQN2_3_r_5,);
nor I_37(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_38(n_42_2_l_5,blif_clk_net_1_r_5,n5_5,ACVQN1_5_r_5,);
not I_39(P6_5_r_5,P6_5_r_internal_5);
and I_40(N3_2_l_5,n19_5,n_452_1_r_1);
not I_41(n5_5,blif_reset_net_1_r_5);
DFFARX1 I_42(N3_2_l_5,blif_clk_net_1_r_5,n5_5,G199_2_l_5,);
DFFARX1 I_43(n_549_1_r_1,blif_clk_net_1_r_5,n5_5,ACVQN2_3_l_5,);
not I_44(n13_5,ACVQN2_3_l_5);
DFFARX1 I_45(n_573_1_r_1,blif_clk_net_1_r_5,n5_5,ACVQN1_3_l_5,);
and I_46(N1_4_l_5,n20_5,G42_1_r_1);
DFFARX1 I_47(N1_4_l_5,blif_clk_net_1_r_5,n5_5,n21_5,);
not I_48(n15_5,n21_5);
DFFARX1 I_49(G42_1_r_1,blif_clk_net_1_r_5,n5_5,n22_5,);
nor I_50(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_51(ACVQN2_3_l_5,blif_clk_net_1_r_5,n5_5,n11_internal_5,);
not I_52(n11_5,n11_internal_5);
nor I_53(n_42_2_l_5,n_572_1_r_1,n_266_and_0_3_r_1);
not I_54(n1_5,n18_5);
DFFARX1 I_55(n1_5,blif_clk_net_1_r_5,n5_5,P6_5_r_internal_5,);
not I_56(n16_5,n_42_2_l_5);
nor I_57(n17_5,n22_5,n18_5);
nand I_58(n18_5,ACVQN1_3_l_5,ACVQN2_3_r_1);
nand I_59(n19_5,n_572_1_r_1,G199_4_r_1);
nand I_60(n20_5,G214_4_r_1,n_572_1_r_1);
endmodule


