module test_I7156(I3368,I1477,I5204,I1470,I7088,I5249,I7156);
input I3368,I1477,I5204,I1470,I7088,I5249;
output I7156;
wire I5076,I7122,I5266,I5079,I5105,I7105,I5085,I6907,I5512,I7139;
DFFARX1 I_0(I5204,I1470,I5105,,,I5076,);
and I_1(I7122,I7105,I5076);
not I_2(I5266,I5249);
DFFARX1 I_3(I1470,I5105,,,I5079,);
not I_4(I5105,I1477);
DFFARX1 I_5(I7139,I1470,I6907,,,I7156,);
nor I_6(I7105,I7088,I5079);
nand I_7(I5085,I5512,I5266);
not I_8(I6907,I1477);
DFFARX1 I_9(I3368,I1470,I5105,,,I5512,);
or I_10(I7139,I7122,I5085);
endmodule


