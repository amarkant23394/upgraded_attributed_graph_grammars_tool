module test_final(IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_5_r,blif_reset_net_5_r,N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r);
input IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_5_r,blif_reset_net_5_r;
output N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r;
wire N6147_2_l,n5_2_l,n6_2_l,N6138_2_l,n7_2_l,N1507_6_l,N1508_6_l,n6_6_l,n7_6_l,n8_6_l,n9_6_l,N6150_9_l,N6147_9_l,N6134_9_l,n3_9_l,I_BUFF_1_9_l,n4_1_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n_431_5_r,n2_5_r,n11_5_r,n12_5_r,n13_5_r,n14_5_r,n15_5_r,n16_5_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n5_10_r,n6_10_r;
nor I_0(N6147_2_l,n5_2_l,n6_2_l);
nor I_1(n5_2_l,IN_5_2_l,n7_2_l);
not I_2(n6_2_l,N6138_2_l);
nor I_3(N6138_2_l,IN_1_2_l,IN_2_2_l);
nor I_4(n7_2_l,IN_3_2_l,IN_4_2_l);
nor I_5(N1507_6_l,n8_6_l,n9_6_l);
and I_6(N1508_6_l,IN_2_6_l,n6_6_l);
nor I_7(n6_6_l,n7_6_l,n8_6_l);
not I_8(n7_6_l,IN_1_6_l);
nor I_9(n8_6_l,IN_5_6_l,n9_6_l);
and I_10(n9_6_l,IN_3_6_l,IN_4_6_l);
not I_11(N6150_9_l,IN_2_9_l);
nor I_12(N6147_9_l,N6150_9_l,n3_9_l);
nor I_13(N6134_9_l,IN_5_9_l,n3_9_l);
nor I_14(n3_9_l,IN_3_9_l,IN_4_9_l);
buf I_15(I_BUFF_1_9_l,IN_1_9_l);
not I_16(N1372_1_r,n4_1_r);
nor I_17(N1508_1_r,n4_1_r,N6134_9_l);
nand I_18(n4_1_r,I_BUFF_1_9_l,N6147_2_l);
nor I_19(N6147_2_r,n5_2_r,n6_2_r);
nor I_20(n5_2_r,n7_2_r,N1507_6_l);
not I_21(n6_2_r,N6138_2_r);
nor I_22(N6138_2_r,N1507_6_l,N1508_6_l);
nor I_23(n7_2_r,N6147_9_l,N1508_6_l);
nor I_24(N6147_3_r,n3_3_r,N6147_9_l);
not I_25(n3_3_r,N6138_3_r);
nor I_26(N6138_3_r,N6134_9_l,I_BUFF_1_9_l);
nand I_27(n_429_or_0_5_r,n12_5_r,N6147_9_l);
DFFARX1 I_28(n_431_5_r,blif_clk_net_5_r,n2_5_r,G78_5_r,);
nand I_29(n_576_5_r,n11_5_r,N1508_6_l);
not I_30(n_102_5_r,N6147_9_l);
nand I_31(n_547_5_r,n13_5_r,I_BUFF_1_9_l);
or I_32(n_431_5_r,n14_5_r,N6147_2_l);
not I_33(n2_5_r,blif_reset_net_5_r);
nor I_34(n11_5_r,n12_5_r,N6147_9_l);
not I_35(n12_5_r,I_BUFF_1_9_l);
nor I_36(n13_5_r,N6147_9_l,N6147_2_l);
and I_37(n14_5_r,n15_5_r,N6147_2_l);
nor I_38(n15_5_r,n16_5_r,N1507_6_l);
not I_39(n16_5_r,N6147_9_l);
nor I_40(N1507_6_r,n8_6_r,n9_6_r);
and I_41(N1508_6_r,n6_6_r,N6134_9_l);
nor I_42(n6_6_r,n7_6_r,n8_6_r);
not I_43(n7_6_r,N6147_2_l);
nor I_44(n8_6_r,n9_6_r,N1508_6_l);
and I_45(n9_6_r,N6147_2_l,N6134_9_l);
not I_46(N1372_10_r,n6_10_r);
nor I_47(N1508_10_r,n5_10_r,n6_10_r);
nor I_48(n5_10_r,N1507_6_l,N1508_6_l);
nand I_49(n6_10_r,N6134_9_l,N6147_9_l);
endmodule


