module test_I16835(I14982,I1477,I1470,I16835);
input I14982,I1477,I1470;
output I16835;
wire I12619,I12670,I14948,I12584,I15485,I15047,I15064,I14936,I15406,I12587,I15519,I14965,I15372,I15423,I15502;
not I_0(I12619,I1477);
DFFARX1 I_1(I1470,I12619,,,I12670,);
DFFARX1 I_2(I15519,I1470,I14965,,,I14948,);
and I_3(I12584,I12670);
DFFARX1 I_4(I1470,I14965,,,I15485,);
nor I_5(I15047,I14982,I12584);
nand I_6(I15064,I15047,I12587);
DFFARX1 I_7(I15064,I1470,I14965,,,I14936,);
nand I_8(I16835,I14936,I14948);
nor I_9(I15406,I15064);
DFFARX1 I_10(I12670,I1470,I12619,,,I12587,);
or I_11(I15519,I15502,I15423);
not I_12(I14965,I1477);
DFFARX1 I_13(I1470,I14965,,,I15372,);
and I_14(I15423,I15372,I15406);
not I_15(I15502,I15485);
endmodule


