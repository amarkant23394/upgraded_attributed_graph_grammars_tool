module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_8_r_6,n9_6,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_6,n30_6,n33_6);
nor I_43(N1508_0_r_6,n33_6,n44_6);
not I_44(N1372_1_r_6,n41_6);
nor I_45(N1508_1_r_6,n40_6,n41_6);
nor I_46(N1507_6_r_6,n39_6,n45_6);
nor I_47(N1508_6_r_6,n37_6,n38_6);
nor I_48(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_49(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_50(N6147_9_r_6,n32_6,n33_6);
nor I_51(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_52(I_BUFF_1_9_r_6,n37_6);
not I_53(N1372_10_r_6,n43_6);
nor I_54(N1508_10_r_6,n42_6,n43_6);
nor I_55(N3_8_r_6,n36_6,n_429_or_0_5_r_11);
not I_56(n9_6,blif_reset_net_8_r_6);
nor I_57(n30_6,n53_6,N6147_2_r_11);
not I_58(n31_6,n36_6);
nor I_59(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_60(n33_6,n_429_or_0_5_r_11);
not I_61(n34_6,n35_6);
nand I_62(n35_6,n49_6,n_547_5_r_11);
nand I_63(n36_6,n51_6,G78_5_r_11);
nand I_64(n37_6,n54_6,N1507_6_r_11);
or I_65(n38_6,n35_6,n39_6);
nor I_66(n39_6,n40_6,n45_6);
and I_67(n40_6,n46_6,n47_6);
nand I_68(n41_6,n30_6,n31_6);
nor I_69(n42_6,n34_6,n40_6);
nand I_70(n43_6,n30_6,n_429_or_0_5_r_11);
nor I_71(n44_6,n31_6,n40_6);
nor I_72(n45_6,n35_6,n36_6);
nor I_73(n46_6,N1508_1_r_11,N6147_2_r_11);
or I_74(n47_6,n48_6,N1372_1_r_11);
nor I_75(n48_6,N6147_3_r_11,n_576_5_r_11);
and I_76(n49_6,n50_6,N1508_6_r_11);
nand I_77(n50_6,n51_6,n52_6);
nand I_78(n51_6,N1372_1_r_11,n_429_or_0_5_r_11);
not I_79(n52_6,G78_5_r_11);
nor I_80(n53_6,N1508_10_r_11,N6147_3_r_11);
or I_81(n54_6,N1508_10_r_11,N6147_3_r_11);
endmodule


