module test_I17998(I1477,I15579,I17498,I16069,I1470,I17645,I17998);
input I1477,I15579,I17498,I16069,I1470,I17645;
output I17998;
wire I17413,I16007,I17744,I17515,I17679,I15611,I15928,I17727,I17662,I17916,I17430,I15576,I15603,I17933;
not I_0(I17413,I1477);
or I_1(I17998,I17933,I17744);
or I_2(I16007,I15928);
and I_3(I17744,I17727,I17679);
not I_4(I17515,I17498);
nor I_5(I17679,I17662,I17515);
not I_6(I15611,I1477);
DFFARX1 I_7(I1470,I15611,,,I15928,);
nand I_8(I17727,I17430,I15576);
DFFARX1 I_9(I17645,I1470,I17413,,,I17662,);
DFFARX1 I_10(I15603,I1470,I17413,,,I17916,);
not I_11(I17430,I15579);
DFFARX1 I_12(I16007,I1470,I15611,,,I15576,);
nor I_13(I15603,I15928,I16069);
not I_14(I17933,I17916);
endmodule


