module test_I15880(I13908,I1477,I15764,I1470,I13755,I14196,I15880);
input I13908,I1477,I15764,I1470,I13755,I14196;
output I15880;
wire I14162,I13767,I13743,I15832,I15815,I15628,I13749,I15863,I15611,I13775,I15781,I15798;
DFFARX1 I_0(I1470,I13775,,,I14162,);
DFFARX1 I_1(I14196,I1470,I13775,,,I13767,);
DFFARX1 I_2(I1470,I13775,,,I13743,);
nand I_3(I15832,I15628,I13749);
DFFARX1 I_4(I15798,I1470,I15611,,,I15815,);
nor I_5(I15880,I15815,I15863);
not I_6(I15628,I13743);
nand I_7(I13749,I14162,I13908);
not I_8(I15863,I15832);
not I_9(I15611,I1477);
not I_10(I13775,I1477);
and I_11(I15781,I15764,I13755);
or I_12(I15798,I15781,I13767);
endmodule


