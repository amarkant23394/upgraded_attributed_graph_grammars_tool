module test_I14179(I1477,I11953,I1470,I11990,I12106,I12524,I14179);
input I1477,I11953,I1470,I11990,I12106,I12524;
output I14179;
wire I13826,I12270,I11947,I12239,I14162,I10014,I11938,I12208,I13792,I13775,I13809,I11973,I11965;
DFFARX1 I_0(I13809,I1470,I13775,,,I13826,);
nand I_1(I12270,I11990,I10014);
nand I_2(I11947,I12106,I12524);
nand I_3(I14179,I14162,I13826);
DFFARX1 I_4(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_5(I11938,I1470,I13775,,,I14162,);
DFFARX1 I_6(I1470,,,I10014,);
and I_7(I11938,I12270,I12239);
DFFARX1 I_8(I1470,I11973,,,I12208,);
nand I_9(I13792,I11953,I11965);
not I_10(I13775,I1477);
and I_11(I13809,I13792,I11947);
not I_12(I11973,I1477);
DFFARX1 I_13(I1470,I11973,,,I11965,);
endmodule


