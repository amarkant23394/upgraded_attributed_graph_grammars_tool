module test_I2406(I1207,I1294,I1301,I2406);
input I1207,I1294,I1301;
output I2406;
wire I1328,I1622,I1937,I1393,I1828,I2389,I1639,I1780;
nand I_0(I1328,I1639,I1828);
DFFARX1 I_1(I1294,,,I1622,);
not I_2(I1937,I1301);
DFFARX1 I_3(I1294,,,I1393,);
nor I_4(I1828,I1780,I1393);
DFFARX1 I_5(I1328,I1294,I1937,,,I2389,);
and I_6(I1639,I1622,I1207);
not I_7(I2406,I2389);
DFFARX1 I_8(I1294,,,I1780,);
endmodule


