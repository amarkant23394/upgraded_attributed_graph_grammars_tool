module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l;
output N1372_1_r,N1508_1_r,N6147_2_r,N6147_3_r,N1372_4_r,N1508_4_r,N1507_6_r,N1508_6_r,N1372_10_r,N1508_10_r;
wire N1372_1_l,N1508_1_l,n4_1_l,N6147_3_l,n3_3_l,N6138_3_l,N1372_4_l,N1508_4_l,n6_4_l,n7_4_l,n8_4_l,n4_1_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n6_4_r,n7_4_r,n8_4_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n5_10_r,n6_10_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
nor I_3(N6147_3_l,IN_3_3_l,n3_3_l);
not I_4(n3_3_l,N6138_3_l);
nor I_5(N6138_3_l,IN_1_3_l,IN_2_3_l);
not I_6(N1372_4_l,n7_4_l);
nor I_7(N1508_4_l,n6_4_l,n7_4_l);
nor I_8(n6_4_l,IN_5_4_l,n8_4_l);
nand I_9(n7_4_l,IN_1_4_l,IN_2_4_l);
and I_10(n8_4_l,IN_3_4_l,IN_4_4_l);
not I_11(N1372_1_r,n4_1_r);
nor I_12(N1508_1_r,n4_1_r,N1508_4_l);
nand I_13(n4_1_r,N1372_4_l,N1372_1_l);
nor I_14(N6147_2_r,n5_2_r,n6_2_r);
nor I_15(n5_2_r,n7_2_r,N1508_1_l);
not I_16(n6_2_r,N6138_2_r);
nor I_17(N6138_2_r,N1508_1_l,N6147_3_l);
nor I_18(n7_2_r,N6147_3_l,N1508_4_l);
nor I_19(N6147_3_r,n3_3_r,N6147_3_l);
not I_20(n3_3_r,N6138_3_r);
nor I_21(N6138_3_r,N6147_3_l,N1372_4_l);
not I_22(N1372_4_r,n7_4_r);
nor I_23(N1508_4_r,n6_4_r,n7_4_r);
nor I_24(n6_4_r,n8_4_r,N1508_1_l);
nand I_25(n7_4_r,N1508_4_l,N1372_4_l);
and I_26(n8_4_r,N1508_1_l,N1372_1_l);
nor I_27(N1507_6_r,n8_6_r,n9_6_r);
and I_28(N1508_6_r,n6_6_r,N1372_1_l);
nor I_29(n6_6_r,n7_6_r,n8_6_r);
not I_30(n7_6_r,N1508_4_l);
nor I_31(n8_6_r,n9_6_r,N1372_4_l);
and I_32(n9_6_r,N1372_1_l,N1508_4_l);
not I_33(N1372_10_r,n6_10_r);
nor I_34(N1508_10_r,n5_10_r,n6_10_r);
nor I_35(n5_10_r,N1508_1_l,N1372_1_l);
nand I_36(n6_10_r,N6147_3_l,N1372_4_l);
endmodule


