module test_I4544_rst(I1477_rst,I4544_rst);
,I4544_rst);
input I1477_rst;
output I4544_rst;
wire ;
not I_0(I4544_rst,I1477_rst);
endmodule


