module test_I4886(I1477,I4561,I1470,I2678,I4886);
input I1477,I4561,I1470,I2678;
output I4886;
wire I2181,I4544,I4595,I4869,I2149,I4578,I2345,I2161,I2695,I4612;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
DFFARX1 I_2(I4578,I1470,I4544,,,I4595,);
DFFARX1 I_3(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_4(I2695,I1470,I2181,,,I2149,);
and I_5(I4886,I4869,I4612);
and I_6(I4578,I4561,I2161);
DFFARX1 I_7(I1470,I2181,,,I2345,);
nand I_8(I2161,I2345);
and I_9(I2695,I2345,I2678);
not I_10(I4612,I4595);
endmodule


