module test_I13680(I13231,I8851,I1477,I13392,I11281,I1470,I8848,I13680);
input I13231,I8851,I1477,I13392,I11281,I1470,I8848;
output I13680;
wire I11378,I13601,I11429,I13197,I11299,I13265,I13426,I11395,I13248,I13443,I13409;
nor I_0(I11378,I8848);
DFFARX1 I_1(I11299,I1470,I13197,,,I13601,);
and I_2(I13680,I13601,I13443);
not I_3(I11429,I8848);
not I_4(I13197,I1477);
nor I_5(I11299,I11395,I11429);
not I_6(I13265,I13248);
DFFARX1 I_7(I13409,I1470,I13197,,,I13426,);
nand I_8(I11395,I11378,I8851);
DFFARX1 I_9(I13231,I1470,I13197,,,I13248,);
nor I_10(I13443,I13426,I13265);
and I_11(I13409,I13392,I11281);
endmodule


