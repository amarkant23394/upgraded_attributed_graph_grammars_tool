module Benchmark_testing1000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1539,I1546,I4918,I4942,I4924,I4927,I4915,I4933,I4936,I4921,I4930,I4939,I21463,I21442,I21445,I21460,I21457,I21454,I21451,I21439,I21448);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1539,I1546;
output I4918,I4942,I4924,I4927,I4915,I4933,I4936,I4921,I4930,I4939,I21463,I21442,I21445,I21460,I21457,I21454,I21451,I21439,I21448;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1539,I1546,I1581,I5996,I1607,I1624,I1632,I1649,I5993,I5987,I1666,I5981,I1692,I1573,I1564,I5969,I1737,I1745,I5978,I1762,I1561,I5975,I1802,I1810,I1567,I1555,I1855,I5972,I5990,I1872,I1898,I1906,I1549,I1937,I1954,I5984,I1971,I1988,I2005,I1570,I2036,I1558,I1552,I2108,I4326,I2134,I2151,I2159,I2176,I4344,I4329,I2193,I4332,I2219,I2100,I2091,I4320,I2264,I2272,I4323,I2289,I2088,I4335,I2329,I2337,I2094,I2082,I2382,I4341,I4338,I2399,I2425,I2433,I2076,I2464,I2481,I2498,I2515,I2532,I2097,I2563,I2085,I2079,I2635,I3737,I2661,I2669,I2686,I3731,I3725,I2703,I3746,I2729,I3743,I2746,I2754,I3740,I2771,I2603,I2802,I2819,I2615,I2859,I2624,I2881,I3728,I2898,I3749,I2924,I2941,I2627,I2963,I2612,I2994,I3734,I3011,I3028,I3045,I2621,I3076,I2609,I2618,I2606,I3162,I9163,I3188,I3205,I3154,I3227,I9154,I3253,I3261,I3278,I9172,I3295,I9169,I3312,I3329,I9148,I3346,I9151,I3363,I9160,I3380,I3130,I3411,I3428,I3445,I3462,I3142,I3136,I3507,I9166,I3151,I3145,I3552,I3569,I3586,I9157,I3603,I3629,I3637,I3139,I3133,I3691,I3699,I3148,I3757,I17357,I3783,I3800,I3822,I17366,I3848,I3856,I3873,I17354,I3890,I17345,I3907,I3924,I17351,I3941,I17369,I3958,I17342,I3975,I4006,I4023,I4040,I4057,I4102,I17348,I4147,I4164,I17360,I4181,I4198,I17363,I4224,I4232,I4286,I4294,I4352,I14356,I4378,I4395,I4417,I14350,I4443,I4451,I4468,I14368,I4485,I4502,I4519,I4536,I14362,I4553,I14353,I4570,I4601,I4618,I4635,I4652,I4697,I14365,I4742,I4759,I14371,I4776,I4793,I14359,I4819,I4827,I4881,I4889,I4950,I17991,I4976,I4984,I17988,I5001,I18000,I5027,I5049,I5075,I5083,I18006,I5100,I5126,I5148,I17994,I5188,I5205,I5213,I5230,I5261,I18003,I18009,I5278,I5304,I5312,I5357,I17997,I5374,I5477,I18549,I5503,I5511,I18564,I5528,I18567,I5554,I5445,I5576,I18573,I5602,I5610,I18555,I5627,I5653,I5469,I5675,I5451,I18552,I5715,I5732,I5740,I5757,I5454,I5788,I18558,I5805,I18570,I5831,I5839,I5442,I5460,I5884,I18561,I5901,I5463,I5448,I5457,I5466,I6004,I13784,I6030,I6038,I13775,I13790,I6055,I13796,I6081,I6103,I13781,I6129,I6137,I6154,I6180,I6202,I13778,I6242,I6259,I6267,I6284,I6315,I13772,I13787,I6332,I6358,I6366,I6411,I13793,I6428,I6531,I16699,I6557,I6565,I16696,I16714,I6582,I16705,I6608,I6499,I6630,I16720,I6656,I6664,I16702,I6681,I6707,I6523,I6729,I6505,I16708,I6769,I6786,I6794,I6811,I6508,I6842,I16723,I6859,I16711,I6885,I6893,I6496,I6514,I6938,I16717,I6955,I6517,I6502,I6511,I6520,I7058,I7084,I7092,I7109,I7135,I7026,I7157,I7183,I7191,I7208,I7234,I7050,I7256,I7032,I7296,I7313,I7321,I7338,I7035,I7369,I7386,I7412,I7420,I7023,I7041,I7465,I7482,I7044,I7029,I7038,I7047,I7585,I15407,I7611,I7619,I15404,I15422,I7636,I15413,I7662,I7553,I7684,I15428,I7710,I7718,I15410,I7735,I7761,I7577,I7783,I7559,I15416,I7823,I7840,I7848,I7865,I7562,I7896,I15431,I7913,I15419,I7939,I7947,I7550,I7568,I7992,I15425,I8009,I7571,I7556,I7565,I7574,I8112,I20283,I8138,I8146,I20298,I8163,I20301,I8189,I8080,I8211,I20307,I8237,I8245,I20289,I8262,I8288,I8104,I8310,I8086,I20286,I8350,I8367,I8375,I8392,I8089,I8423,I20292,I8440,I20304,I8466,I8474,I8077,I8095,I8519,I20295,I8536,I8098,I8083,I8092,I8101,I8639,I8665,I8682,I8631,I8704,I8721,I8738,I8764,I8772,I8798,I8806,I8823,I8610,I8863,I8871,I8604,I8619,I8916,I8933,I8959,I8607,I8981,I8998,I9015,I8622,I9046,I9063,I8613,I9094,I8616,I8628,I8625,I9180,I9206,I9214,I9240,I9248,I9265,I9282,I9299,I9316,I9347,I9364,I9381,I9398,I9443,I9488,I9505,I9522,I9553,I9570,I9587,I9613,I9621,I9666,I9683,I9700,I9758,I22001,I9784,I9792,I21995,I9818,I9826,I22004,I9843,I21983,I9860,I9877,I21992,I9894,I9744,I9925,I9942,I9959,I22007,I9976,I21986,I9741,I9732,I10021,I9735,I9729,I10066,I21989,I10083,I10100,I9738,I10131,I21998,I10148,I10165,I10191,I10199,I9726,I9750,I10244,I10261,I10278,I9747,I10336,I19127,I10362,I10370,I19133,I10396,I10404,I10421,I19130,I10438,I10455,I19148,I10472,I10322,I10503,I10520,I10537,I19151,I10554,I10319,I10310,I10599,I10313,I10307,I10644,I19136,I10661,I10678,I10316,I10709,I19142,I10726,I19139,I10743,I19145,I10769,I10777,I10304,I10328,I10822,I10839,I10856,I10325,I10914,I10940,I10948,I10974,I10982,I10999,I11016,I11033,I11050,I10900,I11081,I11098,I11115,I11132,I10897,I10888,I11177,I10891,I10885,I11222,I11239,I11256,I10894,I11287,I11304,I11321,I11347,I11355,I10882,I10906,I11400,I11417,I11434,I10903,I11492,I12038,I11518,I11526,I12050,I11552,I11560,I12041,I11577,I12044,I11594,I11611,I12047,I11628,I11478,I11659,I11676,I11693,I11710,I12053,I11475,I11466,I11755,I11469,I11463,I11800,I12059,I11817,I11834,I11472,I11865,I11882,I12056,I11899,I12062,I11925,I11933,I11460,I11484,I11978,I11995,I12012,I11481,I12070,I12096,I12104,I12121,I12138,I12164,I12172,I12198,I12206,I12223,I12240,I12257,I12297,I12305,I12322,I12339,I12356,I12387,I12404,I12430,I12438,I12469,I12500,I12517,I12548,I12648,I12674,I12682,I12699,I12716,I12742,I12750,I12776,I12784,I12801,I12818,I12835,I12631,I12875,I12883,I12900,I12917,I12934,I12634,I12965,I12982,I13008,I13016,I12616,I13047,I12625,I13078,I13095,I12637,I13126,I12628,I12619,I12622,I12640,I13226,I22542,I13252,I13260,I13277,I22530,I22548,I13294,I22539,I13320,I13328,I22554,I22551,I13354,I13362,I13379,I13396,I13413,I13209,I22533,I13453,I13461,I13478,I13495,I13512,I13212,I13543,I22527,I13560,I22536,I13586,I13594,I13194,I13625,I13203,I13656,I13673,I13215,I13704,I22545,I13206,I13197,I13200,I13218,I13804,I13830,I13838,I13855,I13872,I13898,I13906,I13932,I13940,I13957,I13974,I13991,I14031,I14039,I14056,I14073,I14090,I14121,I14138,I14164,I14172,I14203,I14234,I14251,I14282,I14379,I20879,I14405,I14413,I14430,I20861,I14447,I20867,I14473,I20864,I14504,I14512,I20873,I14529,I14555,I14563,I20885,I14603,I14639,I20876,I20870,I14656,I14682,I14690,I14707,I14738,I20882,I14755,I14772,I14803,I14834,I14851,I14906,I14932,I14940,I14957,I14974,I15000,I14895,I15031,I15039,I15056,I15082,I15090,I14898,I15130,I14889,I14880,I15166,I15183,I15209,I15217,I15234,I14883,I15265,I15282,I15299,I14892,I15330,I14877,I15361,I15378,I14886,I15439,I15465,I15482,I15490,I15507,I15524,I15541,I15558,I15575,I15606,I15623,I15654,I15671,I15688,I15719,I15759,I15767,I15784,I15801,I15818,I15849,I15866,I15883,I15909,I15931,I15948,I15979,I16024,I16085,I16111,I16128,I16136,I16153,I16170,I16187,I16204,I16221,I16071,I16252,I16269,I16074,I16300,I16317,I16334,I16050,I16365,I16062,I16405,I16413,I16430,I16447,I16464,I16077,I16495,I16512,I16529,I16555,I16065,I16577,I16594,I16059,I16625,I16053,I16056,I16670,I16068,I16731,I16757,I16774,I16782,I16799,I16816,I16833,I16850,I16867,I16898,I16915,I16946,I16963,I16980,I17011,I17051,I17059,I17076,I17093,I17110,I17141,I17158,I17175,I17201,I17223,I17240,I17271,I17316,I17377,I17403,I17420,I17428,I17445,I17462,I17479,I17496,I17513,I17544,I17561,I17592,I17609,I17626,I17657,I17697,I17705,I17722,I17739,I17756,I17787,I17804,I17821,I17847,I17869,I17886,I17917,I17962,I18017,I18043,I18060,I18082,I18108,I18116,I18133,I18150,I18167,I18184,I18201,I18218,I18249,I18280,I18297,I18314,I18331,I18362,I18407,I18424,I18441,I18467,I18475,I18506,I18523,I18581,I18607,I18615,I18655,I18663,I18680,I18697,I18737,I18759,I18776,I18802,I18810,I18827,I18844,I18861,I18878,I18923,I18954,I18971,I18997,I19005,I19036,I19053,I19070,I19087,I19159,I19185,I19193,I19233,I19241,I19258,I19275,I19315,I19337,I19354,I19380,I19388,I19405,I19422,I19439,I19456,I19501,I19532,I19549,I19575,I19583,I19614,I19631,I19648,I19665,I19737,I19763,I19771,I19720,I19811,I19819,I19836,I19853,I19708,I19893,I19729,I19915,I19932,I19958,I19966,I19983,I20000,I20017,I20034,I19705,I19726,I20079,I19717,I20110,I20127,I20153,I20161,I19723,I20192,I20209,I20226,I20243,I19714,I19711,I20315,I20341,I20349,I20389,I20397,I20414,I20431,I20471,I20493,I20510,I20536,I20544,I20561,I20578,I20595,I20612,I20657,I20688,I20705,I20731,I20739,I20770,I20787,I20804,I20821,I20893,I20919,I20927,I20967,I20975,I20992,I21009,I21049,I21071,I21088,I21114,I21122,I21139,I21156,I21173,I21190,I21235,I21266,I21283,I21309,I21317,I21348,I21365,I21382,I21399,I21471,I21497,I21505,I21531,I21548,I21570,I21587,I21604,I21621,I21638,I21669,I21686,I21703,I21720,I21765,I21782,I21799,I21858,I21884,I21892,I21909,I21926,I21957,I22015,I22041,I22049,I22075,I22092,I22114,I22131,I22148,I22165,I22182,I22213,I22230,I22247,I22264,I22309,I22326,I22343,I22402,I22428,I22436,I22453,I22470,I22501,I22562,I22588,I22596,I22613,I22639,I22647,I22664,I22681,I22712,I22743,I22760,I22777,I22794,I22811,I22842,I22901,I22918,I22944,I22966,I22992,I23000,I23017,I23048;
not I_0 (I1581,I1546);
DFFARX1 I_1 (I5996,I1539,I1581,I1607,);
DFFARX1 I_2 (I1607,I1539,I1581,I1624,);
not I_3 (I1632,I1624);
nand I_4 (I1649,I5993,I5987);
and I_5 (I1666,I1649,I5981);
DFFARX1 I_6 (I1666,I1539,I1581,I1692,);
DFFARX1 I_7 (I1692,I1539,I1581,I1573,);
DFFARX1 I_8 (I1692,I1539,I1581,I1564,);
DFFARX1 I_9 (I5969,I1539,I1581,I1737,);
nand I_10 (I1745,I1737,I5978);
not I_11 (I1762,I1745);
nor I_12 (I1561,I1607,I1762);
DFFARX1 I_13 (I5975,I1539,I1581,I1802,);
not I_14 (I1810,I1802);
nor I_15 (I1567,I1810,I1632);
nand I_16 (I1555,I1810,I1745);
nand I_17 (I1855,I5972,I5990);
and I_18 (I1872,I1855,I5969);
DFFARX1 I_19 (I1872,I1539,I1581,I1898,);
nor I_20 (I1906,I1898,I1607);
DFFARX1 I_21 (I1906,I1539,I1581,I1549,);
not I_22 (I1937,I1898);
nor I_23 (I1954,I5984,I5990);
not I_24 (I1971,I1954);
nor I_25 (I1988,I1745,I1971);
nor I_26 (I2005,I1937,I1988);
DFFARX1 I_27 (I2005,I1539,I1581,I1570,);
nor I_28 (I2036,I1898,I1971);
nor I_29 (I1558,I1762,I2036);
nor I_30 (I1552,I1898,I1954);
not I_31 (I2108,I1546);
DFFARX1 I_32 (I4326,I1539,I2108,I2134,);
DFFARX1 I_33 (I2134,I1539,I2108,I2151,);
not I_34 (I2159,I2151);
nand I_35 (I2176,I4344,I4329);
and I_36 (I2193,I2176,I4332);
DFFARX1 I_37 (I2193,I1539,I2108,I2219,);
DFFARX1 I_38 (I2219,I1539,I2108,I2100,);
DFFARX1 I_39 (I2219,I1539,I2108,I2091,);
DFFARX1 I_40 (I4320,I1539,I2108,I2264,);
nand I_41 (I2272,I2264,I4323);
not I_42 (I2289,I2272);
nor I_43 (I2088,I2134,I2289);
DFFARX1 I_44 (I4335,I1539,I2108,I2329,);
not I_45 (I2337,I2329);
nor I_46 (I2094,I2337,I2159);
nand I_47 (I2082,I2337,I2272);
nand I_48 (I2382,I4341,I4338);
and I_49 (I2399,I2382,I4323);
DFFARX1 I_50 (I2399,I1539,I2108,I2425,);
nor I_51 (I2433,I2425,I2134);
DFFARX1 I_52 (I2433,I1539,I2108,I2076,);
not I_53 (I2464,I2425);
nor I_54 (I2481,I4320,I4338);
not I_55 (I2498,I2481);
nor I_56 (I2515,I2272,I2498);
nor I_57 (I2532,I2464,I2515);
DFFARX1 I_58 (I2532,I1539,I2108,I2097,);
nor I_59 (I2563,I2425,I2498);
nor I_60 (I2085,I2289,I2563);
nor I_61 (I2079,I2425,I2481);
not I_62 (I2635,I1546);
DFFARX1 I_63 (I3737,I1539,I2635,I2661,);
not I_64 (I2669,I2661);
nand I_65 (I2686,I3731,I3725);
and I_66 (I2703,I2686,I3746);
DFFARX1 I_67 (I2703,I1539,I2635,I2729,);
DFFARX1 I_68 (I3743,I1539,I2635,I2746,);
and I_69 (I2754,I2746,I3740);
nor I_70 (I2771,I2729,I2754);
DFFARX1 I_71 (I2771,I1539,I2635,I2603,);
nand I_72 (I2802,I2746,I3740);
nand I_73 (I2819,I2669,I2802);
not I_74 (I2615,I2819);
DFFARX1 I_75 (I3725,I1539,I2635,I2859,);
DFFARX1 I_76 (I2859,I1539,I2635,I2624,);
nand I_77 (I2881,I3728,I3728);
and I_78 (I2898,I2881,I3749);
DFFARX1 I_79 (I2898,I1539,I2635,I2924,);
DFFARX1 I_80 (I2924,I1539,I2635,I2941,);
not I_81 (I2627,I2941);
not I_82 (I2963,I2924);
nand I_83 (I2612,I2963,I2802);
nor I_84 (I2994,I3734,I3728);
not I_85 (I3011,I2994);
nor I_86 (I3028,I2963,I3011);
nor I_87 (I3045,I2669,I3028);
DFFARX1 I_88 (I3045,I1539,I2635,I2621,);
nor I_89 (I3076,I2729,I3011);
nor I_90 (I2609,I2924,I3076);
nor I_91 (I2618,I2859,I2994);
nor I_92 (I2606,I2729,I2994);
not I_93 (I3162,I1546);
DFFARX1 I_94 (I9163,I1539,I3162,I3188,);
DFFARX1 I_95 (I3188,I1539,I3162,I3205,);
not I_96 (I3154,I3205);
not I_97 (I3227,I3188);
DFFARX1 I_98 (I9154,I1539,I3162,I3253,);
not I_99 (I3261,I3253);
and I_100 (I3278,I3227,I9172);
not I_101 (I3295,I9169);
nand I_102 (I3312,I3295,I9172);
not I_103 (I3329,I9148);
nor I_104 (I3346,I3329,I9151);
nand I_105 (I3363,I3346,I9160);
nor I_106 (I3380,I3363,I3312);
DFFARX1 I_107 (I3380,I1539,I3162,I3130,);
not I_108 (I3411,I3363);
not I_109 (I3428,I9151);
nand I_110 (I3445,I3428,I9172);
nor I_111 (I3462,I9151,I9169);
nand I_112 (I3142,I3278,I3462);
nand I_113 (I3136,I3227,I9151);
nand I_114 (I3507,I3329,I9166);
DFFARX1 I_115 (I3507,I1539,I3162,I3151,);
DFFARX1 I_116 (I3507,I1539,I3162,I3145,);
not I_117 (I3552,I9166);
nor I_118 (I3569,I3552,I9148);
and I_119 (I3586,I3569,I9157);
or I_120 (I3603,I3586,I9151);
DFFARX1 I_121 (I3603,I1539,I3162,I3629,);
nand I_122 (I3637,I3629,I3295);
nor I_123 (I3139,I3637,I3445);
nor I_124 (I3133,I3629,I3261);
DFFARX1 I_125 (I3629,I1539,I3162,I3691,);
not I_126 (I3699,I3691);
nor I_127 (I3148,I3699,I3411);
not I_128 (I3757,I1546);
DFFARX1 I_129 (I17357,I1539,I3757,I3783,);
DFFARX1 I_130 (I3783,I1539,I3757,I3800,);
not I_131 (I3749,I3800);
not I_132 (I3822,I3783);
DFFARX1 I_133 (I17366,I1539,I3757,I3848,);
not I_134 (I3856,I3848);
and I_135 (I3873,I3822,I17354);
not I_136 (I3890,I17345);
nand I_137 (I3907,I3890,I17354);
not I_138 (I3924,I17351);
nor I_139 (I3941,I3924,I17369);
nand I_140 (I3958,I3941,I17342);
nor I_141 (I3975,I3958,I3907);
DFFARX1 I_142 (I3975,I1539,I3757,I3725,);
not I_143 (I4006,I3958);
not I_144 (I4023,I17369);
nand I_145 (I4040,I4023,I17354);
nor I_146 (I4057,I17369,I17345);
nand I_147 (I3737,I3873,I4057);
nand I_148 (I3731,I3822,I17369);
nand I_149 (I4102,I3924,I17348);
DFFARX1 I_150 (I4102,I1539,I3757,I3746,);
DFFARX1 I_151 (I4102,I1539,I3757,I3740,);
not I_152 (I4147,I17348);
nor I_153 (I4164,I4147,I17360);
and I_154 (I4181,I4164,I17342);
or I_155 (I4198,I4181,I17363);
DFFARX1 I_156 (I4198,I1539,I3757,I4224,);
nand I_157 (I4232,I4224,I3890);
nor I_158 (I3734,I4232,I4040);
nor I_159 (I3728,I4224,I3856);
DFFARX1 I_160 (I4224,I1539,I3757,I4286,);
not I_161 (I4294,I4286);
nor I_162 (I3743,I4294,I4006);
not I_163 (I4352,I1546);
DFFARX1 I_164 (I14356,I1539,I4352,I4378,);
DFFARX1 I_165 (I4378,I1539,I4352,I4395,);
not I_166 (I4344,I4395);
not I_167 (I4417,I4378);
DFFARX1 I_168 (I14350,I1539,I4352,I4443,);
not I_169 (I4451,I4443);
and I_170 (I4468,I4417,I14368);
not I_171 (I4485,I14356);
nand I_172 (I4502,I4485,I14368);
not I_173 (I4519,I14350);
nor I_174 (I4536,I4519,I14362);
nand I_175 (I4553,I4536,I14353);
nor I_176 (I4570,I4553,I4502);
DFFARX1 I_177 (I4570,I1539,I4352,I4320,);
not I_178 (I4601,I4553);
not I_179 (I4618,I14362);
nand I_180 (I4635,I4618,I14368);
nor I_181 (I4652,I14362,I14356);
nand I_182 (I4332,I4468,I4652);
nand I_183 (I4326,I4417,I14362);
nand I_184 (I4697,I4519,I14365);
DFFARX1 I_185 (I4697,I1539,I4352,I4341,);
DFFARX1 I_186 (I4697,I1539,I4352,I4335,);
not I_187 (I4742,I14365);
nor I_188 (I4759,I4742,I14371);
and I_189 (I4776,I4759,I14353);
or I_190 (I4793,I4776,I14359);
DFFARX1 I_191 (I4793,I1539,I4352,I4819,);
nand I_192 (I4827,I4819,I4485);
nor I_193 (I4329,I4827,I4635);
nor I_194 (I4323,I4819,I4451);
DFFARX1 I_195 (I4819,I1539,I4352,I4881,);
not I_196 (I4889,I4881);
nor I_197 (I4338,I4889,I4601);
not I_198 (I4950,I1546);
DFFARX1 I_199 (I17991,I1539,I4950,I4976,);
nand I_200 (I4984,I17988,I17991);
and I_201 (I5001,I4984,I18000);
DFFARX1 I_202 (I5001,I1539,I4950,I5027,);
nor I_203 (I4918,I5027,I4976);
not I_204 (I5049,I5027);
DFFARX1 I_205 (I17988,I1539,I4950,I5075,);
nand I_206 (I5083,I5075,I18006);
not I_207 (I5100,I5083);
DFFARX1 I_208 (I5100,I1539,I4950,I5126,);
not I_209 (I4942,I5126);
nor I_210 (I5148,I4976,I5083);
nor I_211 (I4924,I5027,I5148);
DFFARX1 I_212 (I17994,I1539,I4950,I5188,);
DFFARX1 I_213 (I5188,I1539,I4950,I5205,);
not I_214 (I5213,I5205);
not I_215 (I5230,I5188);
nand I_216 (I4927,I5230,I5049);
nand I_217 (I5261,I18003,I18009);
and I_218 (I5278,I5261,I17994);
DFFARX1 I_219 (I5278,I1539,I4950,I5304,);
nor I_220 (I5312,I5304,I4976);
DFFARX1 I_221 (I5312,I1539,I4950,I4915,);
DFFARX1 I_222 (I5304,I1539,I4950,I4933,);
nor I_223 (I5357,I17997,I18009);
not I_224 (I5374,I5357);
nor I_225 (I4936,I5213,I5374);
nand I_226 (I4921,I5230,I5374);
nor I_227 (I4930,I4976,I5357);
DFFARX1 I_228 (I5357,I1539,I4950,I4939,);
not I_229 (I5477,I1546);
DFFARX1 I_230 (I18549,I1539,I5477,I5503,);
nand I_231 (I5511,I18564,I18549);
and I_232 (I5528,I5511,I18567);
DFFARX1 I_233 (I5528,I1539,I5477,I5554,);
nor I_234 (I5445,I5554,I5503);
not I_235 (I5576,I5554);
DFFARX1 I_236 (I18573,I1539,I5477,I5602,);
nand I_237 (I5610,I5602,I18555);
not I_238 (I5627,I5610);
DFFARX1 I_239 (I5627,I1539,I5477,I5653,);
not I_240 (I5469,I5653);
nor I_241 (I5675,I5503,I5610);
nor I_242 (I5451,I5554,I5675);
DFFARX1 I_243 (I18552,I1539,I5477,I5715,);
DFFARX1 I_244 (I5715,I1539,I5477,I5732,);
not I_245 (I5740,I5732);
not I_246 (I5757,I5715);
nand I_247 (I5454,I5757,I5576);
nand I_248 (I5788,I18552,I18558);
and I_249 (I5805,I5788,I18570);
DFFARX1 I_250 (I5805,I1539,I5477,I5831,);
nor I_251 (I5839,I5831,I5503);
DFFARX1 I_252 (I5839,I1539,I5477,I5442,);
DFFARX1 I_253 (I5831,I1539,I5477,I5460,);
nor I_254 (I5884,I18561,I18558);
not I_255 (I5901,I5884);
nor I_256 (I5463,I5740,I5901);
nand I_257 (I5448,I5757,I5901);
nor I_258 (I5457,I5503,I5884);
DFFARX1 I_259 (I5884,I1539,I5477,I5466,);
not I_260 (I6004,I1546);
DFFARX1 I_261 (I13784,I1539,I6004,I6030,);
nand I_262 (I6038,I13775,I13790);
and I_263 (I6055,I6038,I13796);
DFFARX1 I_264 (I6055,I1539,I6004,I6081,);
nor I_265 (I5972,I6081,I6030);
not I_266 (I6103,I6081);
DFFARX1 I_267 (I13781,I1539,I6004,I6129,);
nand I_268 (I6137,I6129,I13775);
not I_269 (I6154,I6137);
DFFARX1 I_270 (I6154,I1539,I6004,I6180,);
not I_271 (I5996,I6180);
nor I_272 (I6202,I6030,I6137);
nor I_273 (I5978,I6081,I6202);
DFFARX1 I_274 (I13778,I1539,I6004,I6242,);
DFFARX1 I_275 (I6242,I1539,I6004,I6259,);
not I_276 (I6267,I6259);
not I_277 (I6284,I6242);
nand I_278 (I5981,I6284,I6103);
nand I_279 (I6315,I13772,I13787);
and I_280 (I6332,I6315,I13772);
DFFARX1 I_281 (I6332,I1539,I6004,I6358,);
nor I_282 (I6366,I6358,I6030);
DFFARX1 I_283 (I6366,I1539,I6004,I5969,);
DFFARX1 I_284 (I6358,I1539,I6004,I5987,);
nor I_285 (I6411,I13793,I13787);
not I_286 (I6428,I6411);
nor I_287 (I5990,I6267,I6428);
nand I_288 (I5975,I6284,I6428);
nor I_289 (I5984,I6030,I6411);
DFFARX1 I_290 (I6411,I1539,I6004,I5993,);
not I_291 (I6531,I1546);
DFFARX1 I_292 (I16699,I1539,I6531,I6557,);
nand I_293 (I6565,I16696,I16714);
and I_294 (I6582,I6565,I16705);
DFFARX1 I_295 (I6582,I1539,I6531,I6608,);
nor I_296 (I6499,I6608,I6557);
not I_297 (I6630,I6608);
DFFARX1 I_298 (I16720,I1539,I6531,I6656,);
nand I_299 (I6664,I6656,I16702);
not I_300 (I6681,I6664);
DFFARX1 I_301 (I6681,I1539,I6531,I6707,);
not I_302 (I6523,I6707);
nor I_303 (I6729,I6557,I6664);
nor I_304 (I6505,I6608,I6729);
DFFARX1 I_305 (I16708,I1539,I6531,I6769,);
DFFARX1 I_306 (I6769,I1539,I6531,I6786,);
not I_307 (I6794,I6786);
not I_308 (I6811,I6769);
nand I_309 (I6508,I6811,I6630);
nand I_310 (I6842,I16696,I16723);
and I_311 (I6859,I6842,I16711);
DFFARX1 I_312 (I6859,I1539,I6531,I6885,);
nor I_313 (I6893,I6885,I6557);
DFFARX1 I_314 (I6893,I1539,I6531,I6496,);
DFFARX1 I_315 (I6885,I1539,I6531,I6514,);
nor I_316 (I6938,I16717,I16723);
not I_317 (I6955,I6938);
nor I_318 (I6517,I6794,I6955);
nand I_319 (I6502,I6811,I6955);
nor I_320 (I6511,I6557,I6938);
DFFARX1 I_321 (I6938,I1539,I6531,I6520,);
not I_322 (I7058,I1546);
DFFARX1 I_323 (I1549,I1539,I7058,I7084,);
nand I_324 (I7092,I1573,I1552);
and I_325 (I7109,I7092,I1549);
DFFARX1 I_326 (I7109,I1539,I7058,I7135,);
nor I_327 (I7026,I7135,I7084);
not I_328 (I7157,I7135);
DFFARX1 I_329 (I1555,I1539,I7058,I7183,);
nand I_330 (I7191,I7183,I1564);
not I_331 (I7208,I7191);
DFFARX1 I_332 (I7208,I1539,I7058,I7234,);
not I_333 (I7050,I7234);
nor I_334 (I7256,I7084,I7191);
nor I_335 (I7032,I7135,I7256);
DFFARX1 I_336 (I1558,I1539,I7058,I7296,);
DFFARX1 I_337 (I7296,I1539,I7058,I7313,);
not I_338 (I7321,I7313);
not I_339 (I7338,I7296);
nand I_340 (I7035,I7338,I7157);
nand I_341 (I7369,I1570,I1552);
and I_342 (I7386,I7369,I1561);
DFFARX1 I_343 (I7386,I1539,I7058,I7412,);
nor I_344 (I7420,I7412,I7084);
DFFARX1 I_345 (I7420,I1539,I7058,I7023,);
DFFARX1 I_346 (I7412,I1539,I7058,I7041,);
nor I_347 (I7465,I1567,I1552);
not I_348 (I7482,I7465);
nor I_349 (I7044,I7321,I7482);
nand I_350 (I7029,I7338,I7482);
nor I_351 (I7038,I7084,I7465);
DFFARX1 I_352 (I7465,I1539,I7058,I7047,);
not I_353 (I7585,I1546);
DFFARX1 I_354 (I15407,I1539,I7585,I7611,);
nand I_355 (I7619,I15404,I15422);
and I_356 (I7636,I7619,I15413);
DFFARX1 I_357 (I7636,I1539,I7585,I7662,);
nor I_358 (I7553,I7662,I7611);
not I_359 (I7684,I7662);
DFFARX1 I_360 (I15428,I1539,I7585,I7710,);
nand I_361 (I7718,I7710,I15410);
not I_362 (I7735,I7718);
DFFARX1 I_363 (I7735,I1539,I7585,I7761,);
not I_364 (I7577,I7761);
nor I_365 (I7783,I7611,I7718);
nor I_366 (I7559,I7662,I7783);
DFFARX1 I_367 (I15416,I1539,I7585,I7823,);
DFFARX1 I_368 (I7823,I1539,I7585,I7840,);
not I_369 (I7848,I7840);
not I_370 (I7865,I7823);
nand I_371 (I7562,I7865,I7684);
nand I_372 (I7896,I15404,I15431);
and I_373 (I7913,I7896,I15419);
DFFARX1 I_374 (I7913,I1539,I7585,I7939,);
nor I_375 (I7947,I7939,I7611);
DFFARX1 I_376 (I7947,I1539,I7585,I7550,);
DFFARX1 I_377 (I7939,I1539,I7585,I7568,);
nor I_378 (I7992,I15425,I15431);
not I_379 (I8009,I7992);
nor I_380 (I7571,I7848,I8009);
nand I_381 (I7556,I7865,I8009);
nor I_382 (I7565,I7611,I7992);
DFFARX1 I_383 (I7992,I1539,I7585,I7574,);
not I_384 (I8112,I1546);
DFFARX1 I_385 (I20283,I1539,I8112,I8138,);
nand I_386 (I8146,I20298,I20283);
and I_387 (I8163,I8146,I20301);
DFFARX1 I_388 (I8163,I1539,I8112,I8189,);
nor I_389 (I8080,I8189,I8138);
not I_390 (I8211,I8189);
DFFARX1 I_391 (I20307,I1539,I8112,I8237,);
nand I_392 (I8245,I8237,I20289);
not I_393 (I8262,I8245);
DFFARX1 I_394 (I8262,I1539,I8112,I8288,);
not I_395 (I8104,I8288);
nor I_396 (I8310,I8138,I8245);
nor I_397 (I8086,I8189,I8310);
DFFARX1 I_398 (I20286,I1539,I8112,I8350,);
DFFARX1 I_399 (I8350,I1539,I8112,I8367,);
not I_400 (I8375,I8367);
not I_401 (I8392,I8350);
nand I_402 (I8089,I8392,I8211);
nand I_403 (I8423,I20286,I20292);
and I_404 (I8440,I8423,I20304);
DFFARX1 I_405 (I8440,I1539,I8112,I8466,);
nor I_406 (I8474,I8466,I8138);
DFFARX1 I_407 (I8474,I1539,I8112,I8077,);
DFFARX1 I_408 (I8466,I1539,I8112,I8095,);
nor I_409 (I8519,I20295,I20292);
not I_410 (I8536,I8519);
nor I_411 (I8098,I8375,I8536);
nand I_412 (I8083,I8392,I8536);
nor I_413 (I8092,I8138,I8519);
DFFARX1 I_414 (I8519,I1539,I8112,I8101,);
not I_415 (I8639,I1546);
DFFARX1 I_416 (I1396,I1539,I8639,I8665,);
DFFARX1 I_417 (I8665,I1539,I8639,I8682,);
not I_418 (I8631,I8682);
not I_419 (I8704,I8665);
nand I_420 (I8721,I1364,I1484);
and I_421 (I8738,I8721,I1412);
DFFARX1 I_422 (I8738,I1539,I8639,I8764,);
not I_423 (I8772,I8764);
DFFARX1 I_424 (I1380,I1539,I8639,I8798,);
and I_425 (I8806,I8798,I1428);
nand I_426 (I8823,I8798,I1428);
nand I_427 (I8610,I8772,I8823);
DFFARX1 I_428 (I1420,I1539,I8639,I8863,);
nor I_429 (I8871,I8863,I8806);
DFFARX1 I_430 (I8871,I1539,I8639,I8604,);
nor I_431 (I8619,I8863,I8764);
nand I_432 (I8916,I1444,I1452);
and I_433 (I8933,I8916,I1492);
DFFARX1 I_434 (I8933,I1539,I8639,I8959,);
nor I_435 (I8607,I8959,I8863);
not I_436 (I8981,I8959);
nor I_437 (I8998,I8981,I8772);
nor I_438 (I9015,I8704,I8998);
DFFARX1 I_439 (I9015,I1539,I8639,I8622,);
nor I_440 (I9046,I8981,I8863);
nor I_441 (I9063,I1532,I1452);
nor I_442 (I8613,I9063,I9046);
not I_443 (I9094,I9063);
nand I_444 (I8616,I8823,I9094);
DFFARX1 I_445 (I9063,I1539,I8639,I8628,);
DFFARX1 I_446 (I9063,I1539,I8639,I8625,);
not I_447 (I9180,I1546);
DFFARX1 I_448 (I8083,I1539,I9180,I9206,);
not I_449 (I9214,I9206);
DFFARX1 I_450 (I8098,I1539,I9180,I9240,);
not I_451 (I9248,I8101);
nand I_452 (I9265,I9248,I8080);
not I_453 (I9282,I9265);
nor I_454 (I9299,I9282,I8104);
nor I_455 (I9316,I9214,I9299);
DFFARX1 I_456 (I9316,I1539,I9180,I9166,);
not I_457 (I9347,I8104);
nand I_458 (I9364,I9347,I9282);
and I_459 (I9381,I9347,I8086);
nand I_460 (I9398,I9381,I8077);
nor I_461 (I9163,I9398,I9347);
and I_462 (I9154,I9240,I9398);
not I_463 (I9443,I9398);
nand I_464 (I9157,I9240,I9443);
nor I_465 (I9151,I9206,I9398);
not I_466 (I9488,I8077);
nor I_467 (I9505,I9488,I8086);
nand I_468 (I9522,I9505,I9347);
nor I_469 (I9160,I9265,I9522);
nor I_470 (I9553,I9488,I8092);
and I_471 (I9570,I9553,I8095);
or I_472 (I9587,I9570,I8089);
DFFARX1 I_473 (I9587,I1539,I9180,I9613,);
nor I_474 (I9621,I9613,I9364);
DFFARX1 I_475 (I9621,I1539,I9180,I9148,);
DFFARX1 I_476 (I9613,I1539,I9180,I9172,);
not I_477 (I9666,I9613);
nor I_478 (I9683,I9666,I9240);
nor I_479 (I9700,I9505,I9683);
DFFARX1 I_480 (I9700,I1539,I9180,I9169,);
not I_481 (I9758,I1546);
DFFARX1 I_482 (I22001,I1539,I9758,I9784,);
not I_483 (I9792,I9784);
DFFARX1 I_484 (I21995,I1539,I9758,I9818,);
not I_485 (I9826,I22004);
nand I_486 (I9843,I9826,I21983);
not I_487 (I9860,I9843);
nor I_488 (I9877,I9860,I21992);
nor I_489 (I9894,I9792,I9877);
DFFARX1 I_490 (I9894,I1539,I9758,I9744,);
not I_491 (I9925,I21992);
nand I_492 (I9942,I9925,I9860);
and I_493 (I9959,I9925,I22007);
nand I_494 (I9976,I9959,I21986);
nor I_495 (I9741,I9976,I9925);
and I_496 (I9732,I9818,I9976);
not I_497 (I10021,I9976);
nand I_498 (I9735,I9818,I10021);
nor I_499 (I9729,I9784,I9976);
not I_500 (I10066,I21989);
nor I_501 (I10083,I10066,I22007);
nand I_502 (I10100,I10083,I9925);
nor I_503 (I9738,I9843,I10100);
nor I_504 (I10131,I10066,I21998);
and I_505 (I10148,I10131,I21986);
or I_506 (I10165,I10148,I21983);
DFFARX1 I_507 (I10165,I1539,I9758,I10191,);
nor I_508 (I10199,I10191,I9942);
DFFARX1 I_509 (I10199,I1539,I9758,I9726,);
DFFARX1 I_510 (I10191,I1539,I9758,I9750,);
not I_511 (I10244,I10191);
nor I_512 (I10261,I10244,I9818);
nor I_513 (I10278,I10083,I10261);
DFFARX1 I_514 (I10278,I1539,I9758,I9747,);
not I_515 (I10336,I1546);
DFFARX1 I_516 (I19127,I1539,I10336,I10362,);
not I_517 (I10370,I10362);
DFFARX1 I_518 (I19133,I1539,I10336,I10396,);
not I_519 (I10404,I19127);
nand I_520 (I10421,I10404,I19130);
not I_521 (I10438,I10421);
nor I_522 (I10455,I10438,I19148);
nor I_523 (I10472,I10370,I10455);
DFFARX1 I_524 (I10472,I1539,I10336,I10322,);
not I_525 (I10503,I19148);
nand I_526 (I10520,I10503,I10438);
and I_527 (I10537,I10503,I19151);
nand I_528 (I10554,I10537,I19130);
nor I_529 (I10319,I10554,I10503);
and I_530 (I10310,I10396,I10554);
not I_531 (I10599,I10554);
nand I_532 (I10313,I10396,I10599);
nor I_533 (I10307,I10362,I10554);
not I_534 (I10644,I19136);
nor I_535 (I10661,I10644,I19151);
nand I_536 (I10678,I10661,I10503);
nor I_537 (I10316,I10421,I10678);
nor I_538 (I10709,I10644,I19142);
and I_539 (I10726,I10709,I19139);
or I_540 (I10743,I10726,I19145);
DFFARX1 I_541 (I10743,I1539,I10336,I10769,);
nor I_542 (I10777,I10769,I10520);
DFFARX1 I_543 (I10777,I1539,I10336,I10304,);
DFFARX1 I_544 (I10769,I1539,I10336,I10328,);
not I_545 (I10822,I10769);
nor I_546 (I10839,I10822,I10396);
nor I_547 (I10856,I10661,I10839);
DFFARX1 I_548 (I10856,I1539,I10336,I10325,);
not I_549 (I10914,I1546);
DFFARX1 I_550 (I8616,I1539,I10914,I10940,);
not I_551 (I10948,I10940);
DFFARX1 I_552 (I8628,I1539,I10914,I10974,);
not I_553 (I10982,I8604);
nand I_554 (I10999,I10982,I8631);
not I_555 (I11016,I10999);
nor I_556 (I11033,I11016,I8619);
nor I_557 (I11050,I10948,I11033);
DFFARX1 I_558 (I11050,I1539,I10914,I10900,);
not I_559 (I11081,I8619);
nand I_560 (I11098,I11081,I11016);
and I_561 (I11115,I11081,I8604);
nand I_562 (I11132,I11115,I8607);
nor I_563 (I10897,I11132,I11081);
and I_564 (I10888,I10974,I11132);
not I_565 (I11177,I11132);
nand I_566 (I10891,I10974,I11177);
nor I_567 (I10885,I10940,I11132);
not I_568 (I11222,I8613);
nor I_569 (I11239,I11222,I8604);
nand I_570 (I11256,I11239,I11081);
nor I_571 (I10894,I10999,I11256);
nor I_572 (I11287,I11222,I8622);
and I_573 (I11304,I11287,I8610);
or I_574 (I11321,I11304,I8625);
DFFARX1 I_575 (I11321,I1539,I10914,I11347,);
nor I_576 (I11355,I11347,I11098);
DFFARX1 I_577 (I11355,I1539,I10914,I10882,);
DFFARX1 I_578 (I11347,I1539,I10914,I10906,);
not I_579 (I11400,I11347);
nor I_580 (I11417,I11400,I10974);
nor I_581 (I11434,I11239,I11417);
DFFARX1 I_582 (I11434,I1539,I10914,I10903,);
not I_583 (I11492,I1546);
DFFARX1 I_584 (I12038,I1539,I11492,I11518,);
not I_585 (I11526,I11518);
DFFARX1 I_586 (I12050,I1539,I11492,I11552,);
not I_587 (I11560,I12041);
nand I_588 (I11577,I11560,I12044);
not I_589 (I11594,I11577);
nor I_590 (I11611,I11594,I12047);
nor I_591 (I11628,I11526,I11611);
DFFARX1 I_592 (I11628,I1539,I11492,I11478,);
not I_593 (I11659,I12047);
nand I_594 (I11676,I11659,I11594);
and I_595 (I11693,I11659,I12041);
nand I_596 (I11710,I11693,I12053);
nor I_597 (I11475,I11710,I11659);
and I_598 (I11466,I11552,I11710);
not I_599 (I11755,I11710);
nand I_600 (I11469,I11552,I11755);
nor I_601 (I11463,I11518,I11710);
not I_602 (I11800,I12059);
nor I_603 (I11817,I11800,I12041);
nand I_604 (I11834,I11817,I11659);
nor I_605 (I11472,I11577,I11834);
nor I_606 (I11865,I11800,I12038);
and I_607 (I11882,I11865,I12056);
or I_608 (I11899,I11882,I12062);
DFFARX1 I_609 (I11899,I1539,I11492,I11925,);
nor I_610 (I11933,I11925,I11676);
DFFARX1 I_611 (I11933,I1539,I11492,I11460,);
DFFARX1 I_612 (I11925,I1539,I11492,I11484,);
not I_613 (I11978,I11925);
nor I_614 (I11995,I11978,I11552);
nor I_615 (I12012,I11817,I11995);
DFFARX1 I_616 (I12012,I1539,I11492,I11481,);
not I_617 (I12070,I1546);
DFFARX1 I_618 (I10304,I1539,I12070,I12096,);
not I_619 (I12104,I12096);
nand I_620 (I12121,I10313,I10322);
and I_621 (I12138,I12121,I10328);
DFFARX1 I_622 (I12138,I1539,I12070,I12164,);
not I_623 (I12172,I10325);
DFFARX1 I_624 (I10310,I1539,I12070,I12198,);
not I_625 (I12206,I12198);
nor I_626 (I12223,I12206,I12104);
and I_627 (I12240,I12223,I10325);
nor I_628 (I12257,I12206,I12172);
nor I_629 (I12053,I12164,I12257);
DFFARX1 I_630 (I10319,I1539,I12070,I12297,);
nor I_631 (I12305,I12297,I12164);
not I_632 (I12322,I12305);
not I_633 (I12339,I12297);
nor I_634 (I12356,I12339,I12240);
DFFARX1 I_635 (I12356,I1539,I12070,I12056,);
nand I_636 (I12387,I10316,I10307);
and I_637 (I12404,I12387,I10304);
DFFARX1 I_638 (I12404,I1539,I12070,I12430,);
nor I_639 (I12438,I12430,I12297);
DFFARX1 I_640 (I12438,I1539,I12070,I12038,);
nand I_641 (I12469,I12430,I12339);
nand I_642 (I12047,I12322,I12469);
not I_643 (I12500,I12430);
nor I_644 (I12517,I12500,I12240);
DFFARX1 I_645 (I12517,I1539,I12070,I12059,);
nor I_646 (I12548,I10307,I10307);
or I_647 (I12050,I12297,I12548);
nor I_648 (I12041,I12430,I12548);
or I_649 (I12044,I12164,I12548);
DFFARX1 I_650 (I12548,I1539,I12070,I12062,);
not I_651 (I12648,I1546);
DFFARX1 I_652 (I7047,I1539,I12648,I12674,);
not I_653 (I12682,I12674);
nand I_654 (I12699,I7050,I7026);
and I_655 (I12716,I12699,I7023);
DFFARX1 I_656 (I12716,I1539,I12648,I12742,);
not I_657 (I12750,I7029);
DFFARX1 I_658 (I7023,I1539,I12648,I12776,);
not I_659 (I12784,I12776);
nor I_660 (I12801,I12784,I12682);
and I_661 (I12818,I12801,I7029);
nor I_662 (I12835,I12784,I12750);
nor I_663 (I12631,I12742,I12835);
DFFARX1 I_664 (I7032,I1539,I12648,I12875,);
nor I_665 (I12883,I12875,I12742);
not I_666 (I12900,I12883);
not I_667 (I12917,I12875);
nor I_668 (I12934,I12917,I12818);
DFFARX1 I_669 (I12934,I1539,I12648,I12634,);
nand I_670 (I12965,I7035,I7044);
and I_671 (I12982,I12965,I7041);
DFFARX1 I_672 (I12982,I1539,I12648,I13008,);
nor I_673 (I13016,I13008,I12875);
DFFARX1 I_674 (I13016,I1539,I12648,I12616,);
nand I_675 (I13047,I13008,I12917);
nand I_676 (I12625,I12900,I13047);
not I_677 (I13078,I13008);
nor I_678 (I13095,I13078,I12818);
DFFARX1 I_679 (I13095,I1539,I12648,I12637,);
nor I_680 (I13126,I7038,I7044);
or I_681 (I12628,I12875,I13126);
nor I_682 (I12619,I13008,I13126);
or I_683 (I12622,I12742,I13126);
DFFARX1 I_684 (I13126,I1539,I12648,I12640,);
not I_685 (I13226,I1546);
DFFARX1 I_686 (I22542,I1539,I13226,I13252,);
not I_687 (I13260,I13252);
nand I_688 (I13277,I22530,I22548);
and I_689 (I13294,I13277,I22539);
DFFARX1 I_690 (I13294,I1539,I13226,I13320,);
not I_691 (I13328,I22554);
DFFARX1 I_692 (I22551,I1539,I13226,I13354,);
not I_693 (I13362,I13354);
nor I_694 (I13379,I13362,I13260);
and I_695 (I13396,I13379,I22554);
nor I_696 (I13413,I13362,I13328);
nor I_697 (I13209,I13320,I13413);
DFFARX1 I_698 (I22533,I1539,I13226,I13453,);
nor I_699 (I13461,I13453,I13320);
not I_700 (I13478,I13461);
not I_701 (I13495,I13453);
nor I_702 (I13512,I13495,I13396);
DFFARX1 I_703 (I13512,I1539,I13226,I13212,);
nand I_704 (I13543,I22527,I22527);
and I_705 (I13560,I13543,I22536);
DFFARX1 I_706 (I13560,I1539,I13226,I13586,);
nor I_707 (I13594,I13586,I13453);
DFFARX1 I_708 (I13594,I1539,I13226,I13194,);
nand I_709 (I13625,I13586,I13495);
nand I_710 (I13203,I13478,I13625);
not I_711 (I13656,I13586);
nor I_712 (I13673,I13656,I13396);
DFFARX1 I_713 (I13673,I1539,I13226,I13215,);
nor I_714 (I13704,I22545,I22527);
or I_715 (I13206,I13453,I13704);
nor I_716 (I13197,I13586,I13704);
or I_717 (I13200,I13320,I13704);
DFFARX1 I_718 (I13704,I1539,I13226,I13218,);
not I_719 (I13804,I1546);
DFFARX1 I_720 (I6520,I1539,I13804,I13830,);
not I_721 (I13838,I13830);
nand I_722 (I13855,I6523,I6499);
and I_723 (I13872,I13855,I6496);
DFFARX1 I_724 (I13872,I1539,I13804,I13898,);
not I_725 (I13906,I6502);
DFFARX1 I_726 (I6496,I1539,I13804,I13932,);
not I_727 (I13940,I13932);
nor I_728 (I13957,I13940,I13838);
and I_729 (I13974,I13957,I6502);
nor I_730 (I13991,I13940,I13906);
nor I_731 (I13787,I13898,I13991);
DFFARX1 I_732 (I6505,I1539,I13804,I14031,);
nor I_733 (I14039,I14031,I13898);
not I_734 (I14056,I14039);
not I_735 (I14073,I14031);
nor I_736 (I14090,I14073,I13974);
DFFARX1 I_737 (I14090,I1539,I13804,I13790,);
nand I_738 (I14121,I6508,I6517);
and I_739 (I14138,I14121,I6514);
DFFARX1 I_740 (I14138,I1539,I13804,I14164,);
nor I_741 (I14172,I14164,I14031);
DFFARX1 I_742 (I14172,I1539,I13804,I13772,);
nand I_743 (I14203,I14164,I14073);
nand I_744 (I13781,I14056,I14203);
not I_745 (I14234,I14164);
nor I_746 (I14251,I14234,I13974);
DFFARX1 I_747 (I14251,I1539,I13804,I13793,);
nor I_748 (I14282,I6511,I6517);
or I_749 (I13784,I14031,I14282);
nor I_750 (I13775,I14164,I14282);
or I_751 (I13778,I13898,I14282);
DFFARX1 I_752 (I14282,I1539,I13804,I13796,);
not I_753 (I14379,I1546);
DFFARX1 I_754 (I20879,I1539,I14379,I14405,);
not I_755 (I14413,I14405);
nand I_756 (I14430,I20861,I20861);
and I_757 (I14447,I14430,I20867);
DFFARX1 I_758 (I14447,I1539,I14379,I14473,);
DFFARX1 I_759 (I14473,I1539,I14379,I14368,);
DFFARX1 I_760 (I20864,I1539,I14379,I14504,);
nand I_761 (I14512,I14504,I20873);
not I_762 (I14529,I14512);
DFFARX1 I_763 (I14529,I1539,I14379,I14555,);
not I_764 (I14563,I14555);
nor I_765 (I14371,I14413,I14563);
DFFARX1 I_766 (I20885,I1539,I14379,I14603,);
nor I_767 (I14362,I14603,I14473);
nor I_768 (I14353,I14603,I14529);
nand I_769 (I14639,I20876,I20870);
and I_770 (I14656,I14639,I20864);
DFFARX1 I_771 (I14656,I1539,I14379,I14682,);
not I_772 (I14690,I14682);
nand I_773 (I14707,I14690,I14603);
nand I_774 (I14356,I14690,I14512);
nor I_775 (I14738,I20882,I20870);
and I_776 (I14755,I14603,I14738);
nor I_777 (I14772,I14690,I14755);
DFFARX1 I_778 (I14772,I1539,I14379,I14365,);
nor I_779 (I14803,I14405,I14738);
DFFARX1 I_780 (I14803,I1539,I14379,I14350,);
nor I_781 (I14834,I14682,I14738);
not I_782 (I14851,I14834);
nand I_783 (I14359,I14851,I14707);
not I_784 (I14906,I1546);
DFFARX1 I_785 (I13194,I1539,I14906,I14932,);
not I_786 (I14940,I14932);
nand I_787 (I14957,I13197,I13194);
and I_788 (I14974,I14957,I13206);
DFFARX1 I_789 (I14974,I1539,I14906,I15000,);
DFFARX1 I_790 (I15000,I1539,I14906,I14895,);
DFFARX1 I_791 (I13203,I1539,I14906,I15031,);
nand I_792 (I15039,I15031,I13209);
not I_793 (I15056,I15039);
DFFARX1 I_794 (I15056,I1539,I14906,I15082,);
not I_795 (I15090,I15082);
nor I_796 (I14898,I14940,I15090);
DFFARX1 I_797 (I13218,I1539,I14906,I15130,);
nor I_798 (I14889,I15130,I15000);
nor I_799 (I14880,I15130,I15056);
nand I_800 (I15166,I13212,I13200);
and I_801 (I15183,I15166,I13197);
DFFARX1 I_802 (I15183,I1539,I14906,I15209,);
not I_803 (I15217,I15209);
nand I_804 (I15234,I15217,I15130);
nand I_805 (I14883,I15217,I15039);
nor I_806 (I15265,I13215,I13200);
and I_807 (I15282,I15130,I15265);
nor I_808 (I15299,I15217,I15282);
DFFARX1 I_809 (I15299,I1539,I14906,I14892,);
nor I_810 (I15330,I14932,I15265);
DFFARX1 I_811 (I15330,I1539,I14906,I14877,);
nor I_812 (I15361,I15209,I15265);
not I_813 (I15378,I15361);
nand I_814 (I14886,I15378,I15234);
not I_815 (I15439,I1546);
DFFARX1 I_816 (I14883,I1539,I15439,I15465,);
DFFARX1 I_817 (I14880,I1539,I15439,I15482,);
not I_818 (I15490,I15482);
not I_819 (I15507,I14880);
nor I_820 (I15524,I15507,I14883);
not I_821 (I15541,I14895);
nor I_822 (I15558,I15524,I14889);
nor I_823 (I15575,I15482,I15558);
DFFARX1 I_824 (I15575,I1539,I15439,I15425,);
nor I_825 (I15606,I14889,I14883);
nand I_826 (I15623,I15606,I14880);
DFFARX1 I_827 (I15623,I1539,I15439,I15428,);
nor I_828 (I15654,I15541,I14889);
nand I_829 (I15671,I15654,I14877);
nor I_830 (I15688,I15465,I15671);
DFFARX1 I_831 (I15688,I1539,I15439,I15404,);
not I_832 (I15719,I15671);
nand I_833 (I15416,I15482,I15719);
DFFARX1 I_834 (I15671,I1539,I15439,I15759,);
not I_835 (I15767,I15759);
not I_836 (I15784,I14889);
not I_837 (I15801,I14886);
nor I_838 (I15818,I15801,I14895);
nor I_839 (I15431,I15767,I15818);
nor I_840 (I15849,I15801,I14892);
and I_841 (I15866,I15849,I14898);
or I_842 (I15883,I15866,I14877);
DFFARX1 I_843 (I15883,I1539,I15439,I15909,);
nor I_844 (I15419,I15909,I15465);
not I_845 (I15931,I15909);
and I_846 (I15948,I15931,I15465);
nor I_847 (I15413,I15490,I15948);
nand I_848 (I15979,I15931,I15541);
nor I_849 (I15407,I15801,I15979);
nand I_850 (I15410,I15931,I15719);
nand I_851 (I16024,I15541,I14886);
nor I_852 (I15422,I15784,I16024);
not I_853 (I16085,I1546);
DFFARX1 I_854 (I10885,I1539,I16085,I16111,);
DFFARX1 I_855 (I10897,I1539,I16085,I16128,);
not I_856 (I16136,I16128);
not I_857 (I16153,I10906);
nor I_858 (I16170,I16153,I10882);
not I_859 (I16187,I10900);
nor I_860 (I16204,I16170,I10894);
nor I_861 (I16221,I16128,I16204);
DFFARX1 I_862 (I16221,I1539,I16085,I16071,);
nor I_863 (I16252,I10894,I10882);
nand I_864 (I16269,I16252,I10906);
DFFARX1 I_865 (I16269,I1539,I16085,I16074,);
nor I_866 (I16300,I16187,I10894);
nand I_867 (I16317,I16300,I10888);
nor I_868 (I16334,I16111,I16317);
DFFARX1 I_869 (I16334,I1539,I16085,I16050,);
not I_870 (I16365,I16317);
nand I_871 (I16062,I16128,I16365);
DFFARX1 I_872 (I16317,I1539,I16085,I16405,);
not I_873 (I16413,I16405);
not I_874 (I16430,I10894);
not I_875 (I16447,I10903);
nor I_876 (I16464,I16447,I10900);
nor I_877 (I16077,I16413,I16464);
nor I_878 (I16495,I16447,I10885);
and I_879 (I16512,I16495,I10882);
or I_880 (I16529,I16512,I10891);
DFFARX1 I_881 (I16529,I1539,I16085,I16555,);
nor I_882 (I16065,I16555,I16111);
not I_883 (I16577,I16555);
and I_884 (I16594,I16577,I16111);
nor I_885 (I16059,I16136,I16594);
nand I_886 (I16625,I16577,I16187);
nor I_887 (I16053,I16447,I16625);
nand I_888 (I16056,I16577,I16365);
nand I_889 (I16670,I16187,I10903);
nor I_890 (I16068,I16430,I16670);
not I_891 (I16731,I1546);
DFFARX1 I_892 (I5442,I1539,I16731,I16757,);
DFFARX1 I_893 (I5448,I1539,I16731,I16774,);
not I_894 (I16782,I16774);
not I_895 (I16799,I5469);
nor I_896 (I16816,I16799,I5457);
not I_897 (I16833,I5466);
nor I_898 (I16850,I16816,I5451);
nor I_899 (I16867,I16774,I16850);
DFFARX1 I_900 (I16867,I1539,I16731,I16717,);
nor I_901 (I16898,I5451,I5457);
nand I_902 (I16915,I16898,I5469);
DFFARX1 I_903 (I16915,I1539,I16731,I16720,);
nor I_904 (I16946,I16833,I5451);
nand I_905 (I16963,I16946,I5442);
nor I_906 (I16980,I16757,I16963);
DFFARX1 I_907 (I16980,I1539,I16731,I16696,);
not I_908 (I17011,I16963);
nand I_909 (I16708,I16774,I17011);
DFFARX1 I_910 (I16963,I1539,I16731,I17051,);
not I_911 (I17059,I17051);
not I_912 (I17076,I5451);
not I_913 (I17093,I5454);
nor I_914 (I17110,I17093,I5466);
nor I_915 (I16723,I17059,I17110);
nor I_916 (I17141,I17093,I5463);
and I_917 (I17158,I17141,I5445);
or I_918 (I17175,I17158,I5460);
DFFARX1 I_919 (I17175,I1539,I16731,I17201,);
nor I_920 (I16711,I17201,I16757);
not I_921 (I17223,I17201);
and I_922 (I17240,I17223,I16757);
nor I_923 (I16705,I16782,I17240);
nand I_924 (I17271,I17223,I16833);
nor I_925 (I16699,I17093,I17271);
nand I_926 (I16702,I17223,I17011);
nand I_927 (I17316,I16833,I5454);
nor I_928 (I16714,I17076,I17316);
not I_929 (I17377,I1546);
DFFARX1 I_930 (I9729,I1539,I17377,I17403,);
DFFARX1 I_931 (I9741,I1539,I17377,I17420,);
not I_932 (I17428,I17420);
not I_933 (I17445,I9750);
nor I_934 (I17462,I17445,I9726);
not I_935 (I17479,I9744);
nor I_936 (I17496,I17462,I9738);
nor I_937 (I17513,I17420,I17496);
DFFARX1 I_938 (I17513,I1539,I17377,I17363,);
nor I_939 (I17544,I9738,I9726);
nand I_940 (I17561,I17544,I9750);
DFFARX1 I_941 (I17561,I1539,I17377,I17366,);
nor I_942 (I17592,I17479,I9738);
nand I_943 (I17609,I17592,I9732);
nor I_944 (I17626,I17403,I17609);
DFFARX1 I_945 (I17626,I1539,I17377,I17342,);
not I_946 (I17657,I17609);
nand I_947 (I17354,I17420,I17657);
DFFARX1 I_948 (I17609,I1539,I17377,I17697,);
not I_949 (I17705,I17697);
not I_950 (I17722,I9738);
not I_951 (I17739,I9747);
nor I_952 (I17756,I17739,I9744);
nor I_953 (I17369,I17705,I17756);
nor I_954 (I17787,I17739,I9729);
and I_955 (I17804,I17787,I9726);
or I_956 (I17821,I17804,I9735);
DFFARX1 I_957 (I17821,I1539,I17377,I17847,);
nor I_958 (I17357,I17847,I17403);
not I_959 (I17869,I17847);
and I_960 (I17886,I17869,I17403);
nor I_961 (I17351,I17428,I17886);
nand I_962 (I17917,I17869,I17479);
nor I_963 (I17345,I17739,I17917);
nand I_964 (I17348,I17869,I17657);
nand I_965 (I17962,I17479,I9747);
nor I_966 (I17360,I17722,I17962);
not I_967 (I18017,I1546);
DFFARX1 I_968 (I12619,I1539,I18017,I18043,);
DFFARX1 I_969 (I18043,I1539,I18017,I18060,);
not I_970 (I18009,I18060);
not I_971 (I18082,I18043);
DFFARX1 I_972 (I12631,I1539,I18017,I18108,);
nand I_973 (I18116,I18108,I12640);
not I_974 (I18133,I12640);
not I_975 (I18150,I12622);
nand I_976 (I18167,I12625,I12616);
and I_977 (I18184,I12625,I12616);
not I_978 (I18201,I12634);
nand I_979 (I18218,I18201,I18150);
nor I_980 (I17991,I18218,I18116);
nor I_981 (I18249,I18133,I18218);
nand I_982 (I17994,I18184,I18249);
not I_983 (I18280,I12637);
nor I_984 (I18297,I18280,I12625);
nor I_985 (I18314,I18297,I12634);
nor I_986 (I18331,I18082,I18314);
DFFARX1 I_987 (I18331,I1539,I18017,I18003,);
not I_988 (I18362,I18297);
DFFARX1 I_989 (I18362,I1539,I18017,I18006,);
and I_990 (I18000,I18108,I18297);
nor I_991 (I18407,I18280,I12616);
and I_992 (I18424,I18407,I12628);
or I_993 (I18441,I18424,I12619);
DFFARX1 I_994 (I18441,I1539,I18017,I18467,);
nor I_995 (I18475,I18467,I18201);
DFFARX1 I_996 (I18475,I1539,I18017,I17988,);
nand I_997 (I18506,I18467,I18108);
nand I_998 (I18523,I18201,I18506);
nor I_999 (I17997,I18523,I18167);
not I_1000 (I18581,I1546);
DFFARX1 I_1001 (I2076,I1539,I18581,I18607,);
and I_1002 (I18615,I18607,I2079);
DFFARX1 I_1003 (I18615,I1539,I18581,I18564,);
DFFARX1 I_1004 (I2079,I1539,I18581,I18655,);
not I_1005 (I18663,I2082);
not I_1006 (I18680,I2097);
nand I_1007 (I18697,I18680,I18663);
nor I_1008 (I18552,I18655,I18697);
DFFARX1 I_1009 (I18697,I1539,I18581,I18737,);
not I_1010 (I18573,I18737);
not I_1011 (I18759,I2091);
nand I_1012 (I18776,I18680,I18759);
DFFARX1 I_1013 (I18776,I1539,I18581,I18802,);
not I_1014 (I18810,I18802);
not I_1015 (I18827,I2094);
nand I_1016 (I18844,I18827,I2076);
and I_1017 (I18861,I18663,I18844);
nor I_1018 (I18878,I18776,I18861);
DFFARX1 I_1019 (I18878,I1539,I18581,I18549,);
DFFARX1 I_1020 (I18861,I1539,I18581,I18570,);
nor I_1021 (I18923,I2094,I2088);
nor I_1022 (I18561,I18776,I18923);
or I_1023 (I18954,I2094,I2088);
nor I_1024 (I18971,I2085,I2100);
DFFARX1 I_1025 (I18971,I1539,I18581,I18997,);
not I_1026 (I19005,I18997);
nor I_1027 (I18567,I19005,I18810);
nand I_1028 (I19036,I19005,I18655);
not I_1029 (I19053,I2085);
nand I_1030 (I19070,I19053,I18759);
nand I_1031 (I19087,I19005,I19070);
nand I_1032 (I18558,I19087,I19036);
nand I_1033 (I18555,I19070,I18954);
not I_1034 (I19159,I1546);
DFFARX1 I_1035 (I16056,I1539,I19159,I19185,);
and I_1036 (I19193,I19185,I16050);
DFFARX1 I_1037 (I19193,I1539,I19159,I19142,);
DFFARX1 I_1038 (I16068,I1539,I19159,I19233,);
not I_1039 (I19241,I16059);
not I_1040 (I19258,I16071);
nand I_1041 (I19275,I19258,I19241);
nor I_1042 (I19130,I19233,I19275);
DFFARX1 I_1043 (I19275,I1539,I19159,I19315,);
not I_1044 (I19151,I19315);
not I_1045 (I19337,I16077);
nand I_1046 (I19354,I19258,I19337);
DFFARX1 I_1047 (I19354,I1539,I19159,I19380,);
not I_1048 (I19388,I19380);
not I_1049 (I19405,I16053);
nand I_1050 (I19422,I19405,I16074);
and I_1051 (I19439,I19241,I19422);
nor I_1052 (I19456,I19354,I19439);
DFFARX1 I_1053 (I19456,I1539,I19159,I19127,);
DFFARX1 I_1054 (I19439,I1539,I19159,I19148,);
nor I_1055 (I19501,I16053,I16065);
nor I_1056 (I19139,I19354,I19501);
or I_1057 (I19532,I16053,I16065);
nor I_1058 (I19549,I16050,I16062);
DFFARX1 I_1059 (I19549,I1539,I19159,I19575,);
not I_1060 (I19583,I19575);
nor I_1061 (I19145,I19583,I19388);
nand I_1062 (I19614,I19583,I19233);
not I_1063 (I19631,I16050);
nand I_1064 (I19648,I19631,I19337);
nand I_1065 (I19665,I19583,I19648);
nand I_1066 (I19136,I19665,I19614);
nand I_1067 (I19133,I19648,I19532);
not I_1068 (I19737,I1546);
DFFARX1 I_1069 (I2627,I1539,I19737,I19763,);
and I_1070 (I19771,I19763,I2603);
DFFARX1 I_1071 (I19771,I1539,I19737,I19720,);
DFFARX1 I_1072 (I2621,I1539,I19737,I19811,);
not I_1073 (I19819,I2609);
not I_1074 (I19836,I2606);
nand I_1075 (I19853,I19836,I19819);
nor I_1076 (I19708,I19811,I19853);
DFFARX1 I_1077 (I19853,I1539,I19737,I19893,);
not I_1078 (I19729,I19893);
not I_1079 (I19915,I2615);
nand I_1080 (I19932,I19836,I19915);
DFFARX1 I_1081 (I19932,I1539,I19737,I19958,);
not I_1082 (I19966,I19958);
not I_1083 (I19983,I2606);
nand I_1084 (I20000,I19983,I2624);
and I_1085 (I20017,I19819,I20000);
nor I_1086 (I20034,I19932,I20017);
DFFARX1 I_1087 (I20034,I1539,I19737,I19705,);
DFFARX1 I_1088 (I20017,I1539,I19737,I19726,);
nor I_1089 (I20079,I2606,I2618);
nor I_1090 (I19717,I19932,I20079);
or I_1091 (I20110,I2606,I2618);
nor I_1092 (I20127,I2612,I2603);
DFFARX1 I_1093 (I20127,I1539,I19737,I20153,);
not I_1094 (I20161,I20153);
nor I_1095 (I19723,I20161,I19966);
nand I_1096 (I20192,I20161,I19811);
not I_1097 (I20209,I2612);
nand I_1098 (I20226,I20209,I19915);
nand I_1099 (I20243,I20161,I20226);
nand I_1100 (I19714,I20243,I20192);
nand I_1101 (I19711,I20226,I20110);
not I_1102 (I20315,I1546);
DFFARX1 I_1103 (I1508,I1539,I20315,I20341,);
and I_1104 (I20349,I20341,I1404);
DFFARX1 I_1105 (I20349,I1539,I20315,I20298,);
DFFARX1 I_1106 (I1460,I1539,I20315,I20389,);
not I_1107 (I20397,I1372);
not I_1108 (I20414,I1468);
nand I_1109 (I20431,I20414,I20397);
nor I_1110 (I20286,I20389,I20431);
DFFARX1 I_1111 (I20431,I1539,I20315,I20471,);
not I_1112 (I20307,I20471);
not I_1113 (I20493,I1516);
nand I_1114 (I20510,I20414,I20493);
DFFARX1 I_1115 (I20510,I1539,I20315,I20536,);
not I_1116 (I20544,I20536);
not I_1117 (I20561,I1524);
nand I_1118 (I20578,I20561,I1500);
and I_1119 (I20595,I20397,I20578);
nor I_1120 (I20612,I20510,I20595);
DFFARX1 I_1121 (I20612,I1539,I20315,I20283,);
DFFARX1 I_1122 (I20595,I1539,I20315,I20304,);
nor I_1123 (I20657,I1524,I1388);
nor I_1124 (I20295,I20510,I20657);
or I_1125 (I20688,I1524,I1388);
nor I_1126 (I20705,I1436,I1476);
DFFARX1 I_1127 (I20705,I1539,I20315,I20731,);
not I_1128 (I20739,I20731);
nor I_1129 (I20301,I20739,I20544);
nand I_1130 (I20770,I20739,I20389);
not I_1131 (I20787,I1436);
nand I_1132 (I20804,I20787,I20493);
nand I_1133 (I20821,I20739,I20804);
nand I_1134 (I20292,I20821,I20770);
nand I_1135 (I20289,I20804,I20688);
not I_1136 (I20893,I1546);
DFFARX1 I_1137 (I3130,I1539,I20893,I20919,);
and I_1138 (I20927,I20919,I3133);
DFFARX1 I_1139 (I20927,I1539,I20893,I20876,);
DFFARX1 I_1140 (I3133,I1539,I20893,I20967,);
not I_1141 (I20975,I3148);
not I_1142 (I20992,I3154);
nand I_1143 (I21009,I20992,I20975);
nor I_1144 (I20864,I20967,I21009);
DFFARX1 I_1145 (I21009,I1539,I20893,I21049,);
not I_1146 (I20885,I21049);
not I_1147 (I21071,I3142);
nand I_1148 (I21088,I20992,I21071);
DFFARX1 I_1149 (I21088,I1539,I20893,I21114,);
not I_1150 (I21122,I21114);
not I_1151 (I21139,I3139);
nand I_1152 (I21156,I21139,I3136);
and I_1153 (I21173,I20975,I21156);
nor I_1154 (I21190,I21088,I21173);
DFFARX1 I_1155 (I21190,I1539,I20893,I20861,);
DFFARX1 I_1156 (I21173,I1539,I20893,I20882,);
nor I_1157 (I21235,I3139,I3130);
nor I_1158 (I20873,I21088,I21235);
or I_1159 (I21266,I3139,I3130);
nor I_1160 (I21283,I3145,I3151);
DFFARX1 I_1161 (I21283,I1539,I20893,I21309,);
not I_1162 (I21317,I21309);
nor I_1163 (I20879,I21317,I21122);
nand I_1164 (I21348,I21317,I20967);
not I_1165 (I21365,I3145);
nand I_1166 (I21382,I21365,I21071);
nand I_1167 (I21399,I21317,I21382);
nand I_1168 (I20870,I21399,I21348);
nand I_1169 (I20867,I21382,I21266);
not I_1170 (I21471,I1546);
DFFARX1 I_1171 (I19729,I1539,I21471,I21497,);
nand I_1172 (I21505,I21497,I19708);
DFFARX1 I_1173 (I19705,I1539,I21471,I21531,);
DFFARX1 I_1174 (I21531,I1539,I21471,I21548,);
not I_1175 (I21463,I21548);
not I_1176 (I21570,I19717);
nor I_1177 (I21587,I19717,I19726);
not I_1178 (I21604,I19714);
nand I_1179 (I21621,I21570,I21604);
nor I_1180 (I21638,I19714,I19717);
and I_1181 (I21442,I21638,I21505);
not I_1182 (I21669,I19723);
nand I_1183 (I21686,I21669,I19720);
nor I_1184 (I21703,I19723,I19705);
not I_1185 (I21720,I21703);
nand I_1186 (I21445,I21587,I21720);
DFFARX1 I_1187 (I21703,I1539,I21471,I21460,);
nor I_1188 (I21765,I19708,I19714);
nor I_1189 (I21782,I21765,I19726);
and I_1190 (I21799,I21782,I21686);
DFFARX1 I_1191 (I21799,I1539,I21471,I21457,);
nor I_1192 (I21454,I21765,I21621);
or I_1193 (I21451,I21703,I21765);
nor I_1194 (I21858,I19708,I19711);
DFFARX1 I_1195 (I21858,I1539,I21471,I21884,);
not I_1196 (I21892,I21884);
nand I_1197 (I21909,I21892,I21570);
nor I_1198 (I21926,I21909,I19726);
DFFARX1 I_1199 (I21926,I1539,I21471,I21439,);
nor I_1200 (I21957,I21892,I21621);
nor I_1201 (I21448,I21765,I21957);
not I_1202 (I22015,I1546);
DFFARX1 I_1203 (I7562,I1539,I22015,I22041,);
nand I_1204 (I22049,I22041,I7565);
DFFARX1 I_1205 (I7559,I1539,I22015,I22075,);
DFFARX1 I_1206 (I22075,I1539,I22015,I22092,);
not I_1207 (I22007,I22092);
not I_1208 (I22114,I7568);
nor I_1209 (I22131,I7568,I7553);
not I_1210 (I22148,I7577);
nand I_1211 (I22165,I22114,I22148);
nor I_1212 (I22182,I7577,I7568);
and I_1213 (I21986,I22182,I22049);
not I_1214 (I22213,I7556);
nand I_1215 (I22230,I22213,I7574);
nor I_1216 (I22247,I7556,I7550);
not I_1217 (I22264,I22247);
nand I_1218 (I21989,I22131,I22264);
DFFARX1 I_1219 (I22247,I1539,I22015,I22004,);
nor I_1220 (I22309,I7571,I7577);
nor I_1221 (I22326,I22309,I7553);
and I_1222 (I22343,I22326,I22230);
DFFARX1 I_1223 (I22343,I1539,I22015,I22001,);
nor I_1224 (I21998,I22309,I22165);
or I_1225 (I21995,I22247,I22309);
nor I_1226 (I22402,I7571,I7550);
DFFARX1 I_1227 (I22402,I1539,I22015,I22428,);
not I_1228 (I22436,I22428);
nand I_1229 (I22453,I22436,I22114);
nor I_1230 (I22470,I22453,I7553);
DFFARX1 I_1231 (I22470,I1539,I22015,I21983,);
nor I_1232 (I22501,I22436,I22165);
nor I_1233 (I21992,I22309,I22501);
not I_1234 (I22562,I1546);
DFFARX1 I_1235 (I11484,I1539,I22562,I22588,);
nand I_1236 (I22596,I22588,I11463);
not I_1237 (I22613,I22596);
DFFARX1 I_1238 (I11475,I1539,I22562,I22639,);
not I_1239 (I22647,I22639);
nor I_1240 (I22664,I11463,I11472);
not I_1241 (I22681,I22664);
DFFARX1 I_1242 (I22681,I1539,I22562,I22548,);
or I_1243 (I22712,I11466,I11463);
DFFARX1 I_1244 (I22712,I1539,I22562,I22551,);
not I_1245 (I22743,I11469);
nor I_1246 (I22760,I22743,I11460);
nor I_1247 (I22777,I22760,I11472);
nor I_1248 (I22794,I11460,I11478);
nor I_1249 (I22811,I22647,I22794);
nor I_1250 (I22536,I22613,I22811);
not I_1251 (I22842,I22794);
nand I_1252 (I22539,I22842,I22596);
nand I_1253 (I22533,I22842,I22664);
nor I_1254 (I22530,I22794,I22777);
nor I_1255 (I22901,I11481,I11466);
not I_1256 (I22918,I22901);
DFFARX1 I_1257 (I22901,I1539,I22562,I22944,);
not I_1258 (I22554,I22944);
nor I_1259 (I22966,I11481,I11460);
DFFARX1 I_1260 (I22966,I1539,I22562,I22992,);
and I_1261 (I23000,I22992,I11463);
nor I_1262 (I23017,I23000,I22918);
DFFARX1 I_1263 (I23017,I1539,I22562,I22545,);
nor I_1264 (I23048,I22992,I22777);
DFFARX1 I_1265 (I23048,I1539,I22562,I22527,);
nor I_1266 (I22542,I22992,I22681);
endmodule


