module test_I4708(I1303,I2475,I1477,I2294,I1470,I2198,I1375,I1271,I4708);
input I1303,I2475,I1477,I2294,I1470,I2198,I1375,I1271;
output I4708;
wire I2215,I2492,I2540,I2181,I2232,I2557,I2574,I2164,I2345,I2393,I2146;
and I_0(I2215,I2198,I1271);
and I_1(I2492,I2294,I2475);
DFFARX1 I_2(I1470,I2181,,,I2540,);
not I_3(I2181,I1477);
DFFARX1 I_4(I2215,I1470,I2181,,,I2232,);
and I_5(I2557,I2540,I1303);
or I_6(I2574,I2557,I2492);
nand I_7(I4708,I2146,I2164);
DFFARX1 I_8(I2574,I1470,I2181,,,I2164,);
DFFARX1 I_9(I1375,I1470,I2181,,,I2345,);
DFFARX1 I_10(I2345,I1470,I2181,,,I2393,);
and I_11(I2146,I2232,I2393);
endmodule


