module test_final(G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_13,blif_reset_net_1_r_13,G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13);
input G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_13,blif_reset_net_1_r_13;
output G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13;
wire G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12,n_431_0_l_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n_569_1_r_13,n4_1_l_13,n7_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13;
DFFARX1 I_0(n4_1_r_12,blif_clk_net_1_r_13,n7_13,G42_1_r_12,);
nor I_1(n_572_1_r_12,n29_12,n30_12);
nand I_2(n_573_1_r_12,n26_12,n27_12);
nor I_3(n_549_1_r_12,n33_12,n34_12);
and I_4(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_5(N3_2_r_12,blif_clk_net_1_r_13,n7_13,G199_2_r_12,);
DFFARX1 I_6(n3_12,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_12,);
not I_7(P6_5_r_12,P6_5_r_internal_12);
or I_8(n_431_0_l_12,IN_8_0_l_12,n36_12);
DFFARX1 I_9(n_431_0_l_12,blif_clk_net_1_r_13,n7_13,n41_12,);
DFFARX1 I_10(IN_2_5_l_12,blif_clk_net_1_r_13,n7_13,ACVQN1_5_l_12,);
not I_11(n22_12,ACVQN1_5_l_12);
DFFARX1 I_12(IN_1_5_l_12,blif_clk_net_1_r_13,n7_13,n42_12,);
nor I_13(n4_1_r_12,n41_12,n31_12);
nor I_14(N3_2_r_12,n22_12,n40_12);
not I_15(n3_12,n39_12);
DFFARX1 I_16(ACVQN1_5_l_12,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_12,);
and I_17(n26_12,IN_5_0_l_12,IN_7_0_l_12);
nor I_18(n27_12,n28_12,n29_12);
not I_19(n28_12,IN_11_0_l_12);
nand I_20(n29_12,n31_12,n32_12);
nand I_21(n30_12,IN_11_0_l_12,n42_12);
not I_22(n31_12,G2_0_l_12);
not I_23(n32_12,IN_10_0_l_12);
nand I_24(n33_12,n31_12,n35_12);
nand I_25(n34_12,IN_5_0_l_12,IN_7_0_l_12);
nand I_26(n35_12,n41_12,n42_12);
and I_27(n36_12,IN_2_0_l_12,n37_12);
nor I_28(n37_12,IN_4_0_l_12,n38_12);
not I_29(n38_12,G1_0_l_12);
nor I_30(n39_12,IN_5_0_l_12,n38_12);
nor I_31(n40_12,G2_0_l_12,n39_12);
DFFARX1 I_32(n4_1_r_13,blif_clk_net_1_r_13,n7_13,G42_1_r_13,);
nor I_33(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_34(n_573_1_r_13,n18_13,n19_13);
nand I_35(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_36(n_569_1_r_13,n17_13,n18_13);
nor I_37(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_38(n_266_and_0_3_l_13,blif_clk_net_1_r_13,n7_13,ACVQN2_3_r_13,);
nor I_39(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_40(n_549_1_l_13,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_13,);
not I_41(P6_5_r_13,P6_5_r_internal_13);
nor I_42(n4_1_l_13,G42_1_r_12,n_573_1_r_12);
not I_43(n7_13,blif_reset_net_1_r_13);
DFFARX1 I_44(n4_1_l_13,blif_clk_net_1_r_13,n7_13,n17_internal_13,);
not I_45(n17_13,n17_internal_13);
DFFARX1 I_46(n_549_1_r_12,blif_clk_net_1_r_13,n7_13,n28_13,);
DFFARX1 I_47(G42_1_r_12,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_13,);
nor I_48(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_49(n_266_and_0_3_l_13,ACVQN1_3_l_13,n_572_1_r_12);
nand I_50(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_51(n_573_1_l_13,blif_clk_net_1_r_13,n7_13,n14_internal_13,);
not I_52(n14_13,n14_internal_13);
and I_53(n_549_1_l_13,n21_13,n26_13);
nand I_54(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_55(n_569_1_l_13,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_13,);
nand I_56(n18_13,n23_13,n24_13);
or I_57(n19_13,n_42_2_r_12,ACVQN1_5_r_12);
not I_58(n20_13,n_573_1_r_12);
not I_59(n21_13,P6_5_r_12);
nand I_60(n22_13,n17_13,n28_13);
not I_61(n23_13,G42_1_r_12);
not I_62(n24_13,G199_2_r_12);
nor I_63(n25_13,n_42_2_r_12,ACVQN1_5_r_12);
nand I_64(n26_13,n27_13,n_572_1_r_12);
not I_65(n27_13,ACVQN1_5_r_12);
endmodule


