module test_I7562(I1477,I7587,I1470,I7782,I6459,I6306,I7562);
input I1477,I7587,I1470,I7782,I6459,I6306;
output I7562;
wire I8107,I6297,I8090,I7816,I6309,I7570,I7799,I7652,I6493,I6380,I6318,I7833,I7669;
not I_0(I8107,I8090);
DFFARX1 I_1(I1470,,,I6297,);
DFFARX1 I_2(I6309,I1470,I7570,,,I8090,);
DFFARX1 I_3(I7799,I1470,I7570,,,I7816,);
nand I_4(I7562,I8107,I7833);
nand I_5(I6309,I6493,I6459);
not I_6(I7570,I1477);
or I_7(I7799,I7782,I6306);
nor I_8(I7652,I7587,I6297);
DFFARX1 I_9(I1470,,,I6493,);
DFFARX1 I_10(I1470,,,I6380,);
not I_11(I6318,I6380);
nor I_12(I7833,I7816,I7669);
nand I_13(I7669,I7652,I6318);
endmodule


