module test_I14083(I12270,I1477,I10041,I1470,I14083);
input I12270,I1477,I10041,I1470;
output I14083;
wire I11956,I12349,I14049,I13775,I11973,I11962,I14066;
DFFARX1 I_0(I14066,I1470,I13775,,,I14083,);
not I_1(I11956,I12349);
DFFARX1 I_2(I10041,I1470,I11973,,,I12349,);
DFFARX1 I_3(I11962,I1470,I13775,,,I14049,);
not I_4(I13775,I1477);
not I_5(I11973,I1477);
nor I_6(I11962,I12349,I12270);
and I_7(I14066,I14049,I11956);
endmodule


