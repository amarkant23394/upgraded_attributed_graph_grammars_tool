module test_final(G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12,n_431_0_l_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_12,blif_clk_net_1_r_9,n5_9,G42_1_r_12,);
nor I_1(n_572_1_r_12,n29_12,n30_12);
nand I_2(n_573_1_r_12,n26_12,n27_12);
nor I_3(n_549_1_r_12,n33_12,n34_12);
and I_4(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_5(N3_2_r_12,blif_clk_net_1_r_9,n5_9,G199_2_r_12,);
DFFARX1 I_6(n3_12,blif_clk_net_1_r_9,n5_9,ACVQN1_5_r_12,);
not I_7(P6_5_r_12,P6_5_r_internal_12);
or I_8(n_431_0_l_12,IN_8_0_l_12,n36_12);
DFFARX1 I_9(n_431_0_l_12,blif_clk_net_1_r_9,n5_9,n41_12,);
DFFARX1 I_10(IN_2_5_l_12,blif_clk_net_1_r_9,n5_9,ACVQN1_5_l_12,);
not I_11(n22_12,ACVQN1_5_l_12);
DFFARX1 I_12(IN_1_5_l_12,blif_clk_net_1_r_9,n5_9,n42_12,);
nor I_13(n4_1_r_12,n41_12,n31_12);
nor I_14(N3_2_r_12,n22_12,n40_12);
not I_15(n3_12,n39_12);
DFFARX1 I_16(ACVQN1_5_l_12,blif_clk_net_1_r_9,n5_9,P6_5_r_internal_12,);
and I_17(n26_12,IN_5_0_l_12,IN_7_0_l_12);
nor I_18(n27_12,n28_12,n29_12);
not I_19(n28_12,IN_11_0_l_12);
nand I_20(n29_12,n31_12,n32_12);
nand I_21(n30_12,IN_11_0_l_12,n42_12);
not I_22(n31_12,G2_0_l_12);
not I_23(n32_12,IN_10_0_l_12);
nand I_24(n33_12,n31_12,n35_12);
nand I_25(n34_12,IN_5_0_l_12,IN_7_0_l_12);
nand I_26(n35_12,n41_12,n42_12);
and I_27(n36_12,IN_2_0_l_12,n37_12);
nor I_28(n37_12,IN_4_0_l_12,n38_12);
not I_29(n38_12,G1_0_l_12);
nor I_30(n39_12,IN_5_0_l_12,n38_12);
nor I_31(n40_12,G2_0_l_12,n39_12);
DFFARX1 I_32(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_33(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_34(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_35(n_549_1_r_9,n17_9,n18_9);
or I_36(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_37(n_452_1_r_9,n26_9,n25_9);
nor I_38(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_39(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_40(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_41(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_42(N3_2_l_9,n22_9,n_573_1_r_12);
not I_43(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_44(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_45(n16_9,n27_9);
DFFARX1 I_46(n_42_2_r_12,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_47(n15_9,n26_9);
DFFARX1 I_48(n_572_1_r_12,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_49(n29_9,n29_internal_9);
and I_50(N1_4_l_9,n24_9,ACVQN1_5_r_12);
DFFARX1 I_51(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_52(n_573_1_r_12,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_53(n28_9,n28_internal_9);
nor I_54(n4_1_r_9,n27_9,n26_9);
nor I_55(N3_2_r_9,n15_9,n21_9);
nor I_56(N1_4_r_9,n16_9,n21_9);
nor I_57(n_42_2_l_9,G42_1_r_12,n_549_1_r_12);
not I_58(n17_9,n_452_1_r_9);
nand I_59(n18_9,n27_9,n15_9);
nor I_60(n19_9,n29_9,n20_9);
not I_61(n20_9,G42_1_r_12);
and I_62(n21_9,n23_9,G42_1_r_12);
nand I_63(n22_9,G42_1_r_12,G199_2_r_12);
nor I_64(n23_9,n29_9,n28_9);
nand I_65(n24_9,n_572_1_r_12,P6_5_r_12);
endmodule


