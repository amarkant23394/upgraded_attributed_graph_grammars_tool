module test_I3972(I1477,I2980,I1447,I3045,I2946,I1470,I2844,I3972);
input I1477,I2980,I1447,I3045,I2946,I1470,I2844;
output I3972;
wire I2733,I3107,I3076,I3983,I2742,I3155,I3200,I4068,I4263,I2724,I3310,I2963,I2745,I3217,I2759,I4246;
nand I_0(I2733,I3217,I3107);
nor I_1(I3107,I3076,I2844);
DFFARX1 I_2(I1447,I1470,I2759,,,I3076,);
or I_3(I3972,I4263,I4068);
not I_4(I3983,I1477);
or I_5(I2742,I3076,I2963);
or I_6(I3155,I3076,I3045);
DFFARX1 I_7(I1470,I2759,,,I3200,);
nor I_8(I4068,I2742,I2724);
and I_9(I4263,I4246,I2733);
DFFARX1 I_10(I3155,I1470,I2759,,,I2724,);
and I_11(I3310,I2844);
DFFARX1 I_12(I2946,I1470,I2759,,,I2963,);
nor I_13(I2745,I2980,I3310);
not I_14(I3217,I3200);
not I_15(I2759,I1477);
DFFARX1 I_16(I2745,I1470,I3983,,,I4246,);
endmodule


