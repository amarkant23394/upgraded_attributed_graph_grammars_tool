module test_I11310(I1477,I11310);
input I1477;
output I11310;
wire ;
not I_0(I11310,I1477);
endmodule


