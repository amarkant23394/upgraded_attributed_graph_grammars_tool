module test_I12599(I11105,I10633,I10664,I1477,I12831,I11184,I9459,I1470,I12599);
input I11105,I10633,I10664,I1477,I12831,I11184,I9459,I1470;
output I12599;
wire I10647,I12930,I10961,I10639,I12848,I12718,I12964,I12619,I12913,I12882,I10615,I11201,I10609;
not I_0(I10647,I1477);
and I_1(I12930,I12913,I10609);
nand I_2(I10961,I10664,I9459);
DFFARX1 I_3(I11201,I1470,I10647,,,I10639,);
DFFARX1 I_4(I12831,I1470,I12619,,,I12848,);
nor I_5(I12718,I10615,I10639);
nor I_6(I12964,I12930,I12882);
not I_7(I12619,I1477);
DFFARX1 I_8(I10633,I1470,I12619,,,I12913,);
nand I_9(I12599,I12718,I12964);
not I_10(I12882,I12848);
DFFARX1 I_11(I10961,I1470,I10647,,,I10615,);
and I_12(I11201,I10961,I11184);
DFFARX1 I_13(I11105,I1470,I10647,,,I10609,);
endmodule


