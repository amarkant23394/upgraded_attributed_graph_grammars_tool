module test_I15573(I13860,I11938,I1470,I13775,I15573);
input I13860,I11938,I1470,I13775;
output I15573;
wire I13908,I13761,I15713,I13743,I15730,I15832,I14162,I15628,I13749,I13891;
not I_0(I13908,I13891);
nand I_1(I13761,I13891,I13860);
not I_2(I15713,I13761);
DFFARX1 I_3(I13891,I1470,I13775,,,I13743,);
not I_4(I15730,I15713);
nand I_5(I15832,I15628,I13749);
DFFARX1 I_6(I11938,I1470,I13775,,,I14162,);
not I_7(I15628,I13743);
nand I_8(I13749,I14162,I13908);
DFFARX1 I_9(I1470,I13775,,,I13891,);
nand I_10(I15573,I15832,I15730);
endmodule


