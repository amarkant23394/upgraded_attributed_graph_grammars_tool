module test_I17222(I1477,I1470,I15228,I17222);
input I1477,I1470,I15228;
output I17222;
wire I14927,I14948,I14936,I17205,I16835,I16869,I16818,I16852,I14957,I14965,I15485,I15502;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
DFFARX1 I_1(I1470,I14965,,,I14948,);
nand I_2(I17222,I17205,I16869);
DFFARX1 I_3(I1470,I14965,,,I14936,);
DFFARX1 I_4(I14927,I1470,I16818,,,I17205,);
nand I_5(I16835,I14936,I14948);
DFFARX1 I_6(I16852,I1470,I16818,,,I16869,);
not I_7(I16818,I1477);
and I_8(I16852,I16835,I14957);
nand I_9(I14957,I15502,I15228);
not I_10(I14965,I1477);
DFFARX1 I_11(I1470,I14965,,,I15485,);
not I_12(I15502,I15485);
endmodule


