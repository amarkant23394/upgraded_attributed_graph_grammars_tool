module test_I14825(I1477,I14503,I13635,I13231,I1470,I14825);
input I1477,I14503,I13635,I13231,I1470;
output I14825;
wire I14667,I14684,I14650,I13165,I14537,I14808,I14370,I13313,I13162,I13197,I14520,I13248,I13361,I13189,I13174;
and I_0(I14667,I14650,I13189);
nand I_1(I14684,I14667,I14537);
DFFARX1 I_2(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_3(I13248,I1470,I13197,,,I13165,);
DFFARX1 I_4(I14520,I1470,I14370,,,I14537,);
DFFARX1 I_5(I13162,I1470,I14370,,,I14808,);
not I_6(I14370,I1477);
DFFARX1 I_7(I1470,I13197,,,I13313,);
and I_8(I13162,I13248,I13361);
not I_9(I13197,I1477);
and I_10(I14520,I14503,I13174);
and I_11(I14825,I14808,I14684);
DFFARX1 I_12(I13231,I1470,I13197,,,I13248,);
DFFARX1 I_13(I13313,I1470,I13197,,,I13361,);
DFFARX1 I_14(I13635,I1470,I13197,,,I13189,);
DFFARX1 I_15(I1470,I13197,,,I13174,);
endmodule


