module test_I10698(I9926,I8202,I8181,I1477,I9559,I1470,I10698);
input I9926,I8202,I8181,I1477,I9559,I1470;
output I10698;
wire I9477,I9576,I9754,I9816,I9480,I9960,I9771,I8178,I10681,I9943,I9833,I9456,I9491;
nor I_0(I9477,I9771,I9833);
nor I_1(I9576,I8181,I8202);
nand I_2(I10698,I10681,I9456);
DFFARX1 I_3(I1470,I9491,,,I9754,);
DFFARX1 I_4(I1470,I9491,,,I9816,);
or I_5(I9480,I9771,I9576);
or I_6(I9960,I9771,I9943);
and I_7(I9771,I9754,I8178);
DFFARX1 I_8(I1470,,,I8178,);
nor I_9(I10681,I9477,I9480);
and I_10(I9943,I9576,I9926);
and I_11(I9833,I9816,I9559);
DFFARX1 I_12(I9960,I1470,I9491,,,I9456,);
not I_13(I9491,I1477);
endmodule


