module test_I14261(I12380,I12304,I1477,I1470,I11990,I12058,I14261);
input I12380,I12304,I1477,I1470,I11990,I12058;
output I14261;
wire I12270,I11959,I12239,I14162,I14244,I11938,I14227,I10014,I12208,I13775,I11973,I13843,I11965;
nand I_0(I12270,I11990,I10014);
nand I_1(I11959,I12058,I12380);
DFFARX1 I_2(I12208,I1470,I11973,,,I12239,);
DFFARX1 I_3(I11938,I1470,I13775,,,I14162,);
nor I_4(I14244,I13843,I14227);
and I_5(I11938,I12270,I12239);
not I_6(I14227,I14162);
DFFARX1 I_7(I1470,,,I10014,);
DFFARX1 I_8(I1470,I11973,,,I12208,);
not I_9(I13775,I1477);
not I_10(I11973,I1477);
nor I_11(I13843,I11959,I11965);
and I_12(I14261,I14162,I14244);
DFFARX1 I_13(I12304,I1470,I11973,,,I11965,);
endmodule


