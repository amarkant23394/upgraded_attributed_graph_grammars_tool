module test_I9179(I1477,I5368,I1470,I5249,I5642,I6924,I9179);
input I1477,I5368,I1470,I5249,I5642,I6924;
output I9179;
wire I6992,I6975,I5070,I7026,I5481,I8862,I5097,I6896;
nand I_0(I6992,I6975,I5097);
nor I_1(I6975,I6924,I5070);
and I_2(I5070,I5249,I5481);
not I_3(I7026,I5070);
DFFARX1 I_4(I1470,,,I5481,);
not I_5(I8862,I1477);
DFFARX1 I_6(I6896,I1470,I8862,,,I9179,);
nand I_7(I5097,I5642,I5368);
nor I_8(I6896,I6992,I7026);
endmodule


