module test_I4308(I1351,I1319,I1447,I1477,I1470,I1335,I4308);
input I1351,I1319,I1447,I1477,I1470,I1335;
output I4308;
wire I2878,I2810,I2759,I3124,I2727,I3076,I2861,I2793,I3983;
not I_0(I2878,I2861);
nand I_1(I2810,I2793,I1335);
not I_2(I2759,I1477);
nor I_3(I3124,I3076,I2878);
nand I_4(I2727,I2810,I3124);
DFFARX1 I_5(I1447,I1470,I2759,,,I3076,);
DFFARX1 I_6(I2727,I1470,I3983,,,I4308,);
not I_7(I2861,I1351);
nor I_8(I2793,I1351,I1319);
not I_9(I3983,I1477);
endmodule


