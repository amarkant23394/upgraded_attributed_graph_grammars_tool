module test_I4962(I1477,I1470,I2678,I4962);
input I1477,I1470,I2678;
output I4962;
wire I2181,I4544,I4869,I2149,I2345,I2695;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
DFFARX1 I_2(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_3(I2695,I1470,I2181,,,I2149,);
not I_4(I4962,I4869);
DFFARX1 I_5(I1470,I2181,,,I2345,);
and I_6(I2695,I2345,I2678);
endmodule


