module Benchmark_testing1000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1627,I1634,I5418,I5415,I5400,I5412,I5406,I5394,I5403,I5409,I5397,I10651,I10654,I10630,I10642,I10657,I10645,I10639,I10633,I10636,I10648,I15941,I15920,I15926,I15935,I15938,I15917,I15932,I15929,I15923);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1627,I1634;
output I5418,I5415,I5400,I5412,I5406,I5394,I5403,I5409,I5397,I10651,I10654,I10630,I10642,I10657,I10645,I10639,I10633,I10636,I10648,I15941,I15920,I15926,I15935,I15938,I15917,I15932,I15929,I15923;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1627,I1634,I1666,I15397,I1692,I1700,I15385,I1717,I1658,I15373,I1757,I1765,I1782,I1799,I15379,I1816,I1833,I1637,I1864,I1881,I1898,I15376,I15391,I1640,I1929,I1946,I15382,I1963,I15394,I1980,I1997,I2014,I1649,I2045,I15388,I2062,I2079,I1655,I2110,I1652,I2141,I2167,I2175,I2192,I1646,I1643,I2264,I13663,I2290,I2307,I2315,I2332,I13651,I13642,I2349,I13639,I2375,I2256,I2247,I13645,I2420,I2428,I13657,I2445,I2244,I13654,I2485,I2493,I2250,I2238,I2538,I13648,I2555,I13660,I2581,I2589,I2232,I2620,I2637,I2654,I2671,I2688,I2253,I2719,I2241,I2235,I2791,I2817,I2825,I2842,I2859,I2885,I2902,I2910,I2927,I2759,I2958,I2975,I2771,I3015,I2780,I3037,I3054,I3080,I3097,I2783,I3119,I2768,I3150,I3167,I3184,I3201,I2777,I3232,I2765,I2774,I2762,I3318,I16507,I3344,I3352,I3369,I16501,I16522,I3386,I16498,I3412,I16519,I3429,I3437,I16516,I3454,I3286,I3485,I3502,I3298,I16504,I3542,I3307,I3564,I16513,I16510,I3581,I16495,I3607,I3624,I3310,I3646,I3295,I3677,I3694,I3711,I3728,I3304,I3759,I3292,I3301,I3289,I3848,I3874,I3882,I3899,I3925,I3816,I3947,I3973,I3981,I3998,I4024,I3840,I4046,I3822,I4086,I4103,I4111,I4128,I3825,I4159,I4176,I4202,I4210,I3813,I3831,I4255,I4272,I3834,I3819,I3828,I3837,I4375,I4401,I4409,I4426,I4452,I4343,I4474,I4500,I4508,I4525,I4551,I4367,I4573,I4349,I4613,I4630,I4638,I4655,I4352,I4686,I4703,I4729,I4737,I4340,I4358,I4782,I4799,I4361,I4346,I4355,I4364,I4902,I13061,I4928,I4936,I13076,I4953,I13079,I4979,I4870,I5001,I13085,I5027,I5035,I13067,I5052,I5078,I4894,I5100,I4876,I13064,I5140,I5157,I5165,I5182,I4879,I5213,I13070,I5230,I13082,I5256,I5264,I4867,I4885,I5309,I13073,I5326,I4888,I4873,I4882,I4891,I5426,I5452,I5469,I5500,I5508,I5525,I5542,I5559,I5576,I5593,I5610,I5641,I5658,I5675,I5720,I5737,I5768,I5785,I5816,I5833,I5850,I5876,I5884,I5915,I5932,I5963,I6021,I6047,I6055,I6081,I6089,I6106,I6123,I6140,I6157,I6007,I6188,I6205,I6222,I6239,I6004,I5995,I6284,I5998,I5992,I6329,I6346,I6363,I6001,I6394,I6411,I6428,I6454,I6462,I5989,I6013,I6507,I6524,I6541,I6010,I6599,I8879,I6625,I6633,I8891,I6659,I6667,I8882,I6684,I8885,I6701,I6718,I8888,I6735,I6585,I6766,I6783,I6800,I6817,I8894,I6582,I6573,I6862,I6576,I6570,I6907,I8900,I6924,I6941,I6579,I6972,I6989,I8897,I7006,I8903,I7032,I7040,I6567,I6591,I7085,I7102,I7119,I6588,I7177,I11282,I7203,I7211,I11279,I7237,I7245,I11276,I7262,I11303,I7279,I7296,I11291,I7313,I7163,I7344,I7361,I7378,I11297,I7395,I11288,I7160,I7151,I7440,I7154,I7148,I7485,I11285,I7502,I7519,I7157,I7550,I11300,I7567,I11294,I7584,I7610,I7618,I7145,I7169,I7663,I7680,I7697,I7166,I7755,I11928,I7781,I7789,I7806,I11925,I11943,I7823,I11940,I7849,I7857,I11922,I7883,I7891,I7908,I7925,I7942,I7738,I11934,I7982,I7990,I8007,I8024,I8041,I7741,I8072,I11937,I8089,I8115,I8123,I7723,I8154,I7732,I8185,I8202,I7744,I8233,I11931,I7735,I7726,I7729,I7747,I8333,I14235,I8359,I8367,I8384,I14217,I14229,I8401,I14232,I8427,I8435,I14226,I14223,I8461,I8469,I8486,I8503,I8520,I8316,I14241,I8560,I8568,I8585,I8602,I8619,I8319,I8650,I14220,I8667,I8693,I8701,I8301,I8732,I8310,I8763,I8780,I8322,I8811,I14238,I8313,I8304,I8307,I8325,I8911,I8937,I8945,I8962,I8979,I9005,I9013,I9039,I9047,I9064,I9081,I9098,I9138,I9146,I9163,I9180,I9197,I9228,I9245,I9271,I9279,I9310,I9341,I9358,I9389,I9486,I9512,I9520,I9537,I9554,I9580,I9475,I9611,I9619,I9636,I9662,I9670,I9478,I9710,I9469,I9460,I9746,I9763,I9789,I9797,I9814,I9463,I9845,I9862,I9879,I9472,I9910,I9457,I9941,I9958,I9466,I10019,I10045,I10062,I10070,I10087,I10104,I10121,I10138,I10155,I10005,I10186,I10203,I10008,I10234,I10251,I10268,I9984,I10299,I9996,I10339,I10347,I10364,I10381,I10398,I10011,I10429,I10446,I10463,I10489,I9999,I10511,I10528,I9993,I10559,I9987,I9990,I10604,I10002,I10665,I12501,I10691,I12483,I10708,I10716,I10733,I12492,I10750,I12504,I10767,I12486,I10784,I12495,I10801,I10832,I10849,I10880,I10897,I12507,I10914,I10945,I10985,I10993,I11010,I11027,I11044,I11075,I12489,I11092,I12498,I11109,I11135,I11157,I11174,I11205,I11250,I11311,I11337,I11354,I11362,I11379,I11396,I11413,I11430,I11447,I11478,I11495,I11526,I11543,I11560,I11591,I11631,I11639,I11656,I11673,I11690,I11721,I11738,I11755,I11781,I11803,I11820,I11851,I11896,I11951,I11977,I11994,I12016,I12042,I12050,I12067,I12084,I12101,I12118,I12135,I12152,I12183,I12214,I12231,I12248,I12265,I12296,I12341,I12358,I12375,I12401,I12409,I12440,I12457,I12515,I12541,I12549,I12589,I12597,I12614,I12631,I12671,I12693,I12710,I12736,I12744,I12761,I12778,I12795,I12812,I12857,I12888,I12905,I12931,I12939,I12970,I12987,I13004,I13021,I13093,I13119,I13127,I13167,I13175,I13192,I13209,I13249,I13271,I13288,I13314,I13322,I13339,I13356,I13373,I13390,I13435,I13466,I13483,I13509,I13517,I13548,I13565,I13582,I13599,I13671,I13697,I13705,I13745,I13753,I13770,I13787,I13827,I13849,I13866,I13892,I13900,I13917,I13934,I13951,I13968,I14013,I14044,I14061,I14087,I14095,I14126,I14143,I14160,I14177,I14249,I14275,I14283,I14323,I14331,I14348,I14365,I14405,I14427,I14444,I14470,I14478,I14495,I14512,I14529,I14546,I14591,I14622,I14639,I14665,I14673,I14704,I14721,I14738,I14755,I14827,I14853,I14861,I14810,I14901,I14909,I14926,I14943,I14798,I14983,I14819,I15005,I15022,I15048,I15056,I15073,I15090,I15107,I15124,I14795,I14816,I15169,I14807,I15200,I15217,I15243,I15251,I14813,I15282,I15299,I15316,I15333,I14804,I14801,I15405,I15431,I15439,I15465,I15482,I15504,I15521,I15538,I15555,I15572,I15603,I15620,I15637,I15654,I15699,I15716,I15733,I15792,I15818,I15826,I15843,I15860,I15891,I15949,I15975,I15983,I16000,I16026,I16034,I16051,I16068,I16085,I16102,I16133,I16150,I16167,I16198,I16215,I16255,I16263,I16294,I16311,I16328,I16345,I16376,I16407,I16433,I16455,I16530,I16556,I16573,I16581,I16626,I16643,I16660,I16677,I16694,I16711,I16728,I16759,I16776,I16821,I16838,I16855,I16886,I16912,I16920,I16951,I16968,I16985,I17011,I17019,I17036;
not I_0 (I1666,I1634);
DFFARX1 I_1 (I15397,I1627,I1666,I1692,);
nand I_2 (I1700,I1692,I15385);
not I_3 (I1717,I1700);
DFFARX1 I_4 (I1717,I1627,I1666,I1658,);
DFFARX1 I_5 (I15373,I1627,I1666,I1757,);
not I_6 (I1765,I1757);
not I_7 (I1782,I15373);
not I_8 (I1799,I15379);
nand I_9 (I1816,I1765,I1799);
nor I_10 (I1833,I1816,I15373);
DFFARX1 I_11 (I1833,I1627,I1666,I1637,);
nor I_12 (I1864,I15379,I15373);
nand I_13 (I1881,I1757,I1864);
nor I_14 (I1898,I15376,I15391);
nor I_15 (I1640,I1816,I15376);
not I_16 (I1929,I15376);
not I_17 (I1946,I15382);
nand I_18 (I1963,I1946,I15394);
nand I_19 (I1980,I1782,I1963);
not I_20 (I1997,I1980);
nor I_21 (I2014,I15382,I15391);
nor I_22 (I1649,I1997,I2014);
nor I_23 (I2045,I15388,I15382);
and I_24 (I2062,I2045,I1898);
nor I_25 (I2079,I1980,I2062);
DFFARX1 I_26 (I2079,I1627,I1666,I1655,);
nor I_27 (I2110,I1700,I2062);
DFFARX1 I_28 (I2110,I1627,I1666,I1652,);
nor I_29 (I2141,I15388,I15376);
DFFARX1 I_30 (I2141,I1627,I1666,I2167,);
nor I_31 (I2175,I2167,I15379);
nand I_32 (I2192,I2175,I1782);
nand I_33 (I1646,I2192,I1881);
nand I_34 (I1643,I2175,I1929);
not I_35 (I2264,I1634);
DFFARX1 I_36 (I13663,I1627,I2264,I2290,);
DFFARX1 I_37 (I2290,I1627,I2264,I2307,);
not I_38 (I2315,I2307);
nand I_39 (I2332,I13651,I13642);
and I_40 (I2349,I2332,I13639);
DFFARX1 I_41 (I2349,I1627,I2264,I2375,);
DFFARX1 I_42 (I2375,I1627,I2264,I2256,);
DFFARX1 I_43 (I2375,I1627,I2264,I2247,);
DFFARX1 I_44 (I13645,I1627,I2264,I2420,);
nand I_45 (I2428,I2420,I13657);
not I_46 (I2445,I2428);
nor I_47 (I2244,I2290,I2445);
DFFARX1 I_48 (I13654,I1627,I2264,I2485,);
not I_49 (I2493,I2485);
nor I_50 (I2250,I2493,I2315);
nand I_51 (I2238,I2493,I2428);
nand I_52 (I2538,I13648,I13642);
and I_53 (I2555,I2538,I13660);
DFFARX1 I_54 (I2555,I1627,I2264,I2581,);
nor I_55 (I2589,I2581,I2290);
DFFARX1 I_56 (I2589,I1627,I2264,I2232,);
not I_57 (I2620,I2581);
nor I_58 (I2637,I13639,I13642);
not I_59 (I2654,I2637);
nor I_60 (I2671,I2428,I2654);
nor I_61 (I2688,I2620,I2671);
DFFARX1 I_62 (I2688,I1627,I2264,I2253,);
nor I_63 (I2719,I2581,I2654);
nor I_64 (I2241,I2445,I2719);
nor I_65 (I2235,I2581,I2637);
not I_66 (I2791,I1634);
DFFARX1 I_67 (I1564,I1627,I2791,I2817,);
not I_68 (I2825,I2817);
nand I_69 (I2842,I1604,I1492);
and I_70 (I2859,I2842,I1508);
DFFARX1 I_71 (I2859,I1627,I2791,I2885,);
DFFARX1 I_72 (I1500,I1627,I2791,I2902,);
and I_73 (I2910,I2902,I1596);
nor I_74 (I2927,I2885,I2910);
DFFARX1 I_75 (I2927,I1627,I2791,I2759,);
nand I_76 (I2958,I2902,I1596);
nand I_77 (I2975,I2825,I2958);
not I_78 (I2771,I2975);
DFFARX1 I_79 (I1468,I1627,I2791,I3015,);
DFFARX1 I_80 (I3015,I1627,I2791,I2780,);
nand I_81 (I3037,I1388,I1412);
and I_82 (I3054,I3037,I1556);
DFFARX1 I_83 (I3054,I1627,I2791,I3080,);
DFFARX1 I_84 (I3080,I1627,I2791,I3097,);
not I_85 (I2783,I3097);
not I_86 (I3119,I3080);
nand I_87 (I2768,I3119,I2958);
nor I_88 (I3150,I1404,I1412);
not I_89 (I3167,I3150);
nor I_90 (I3184,I3119,I3167);
nor I_91 (I3201,I2825,I3184);
DFFARX1 I_92 (I3201,I1627,I2791,I2777,);
nor I_93 (I3232,I2885,I3167);
nor I_94 (I2765,I3080,I3232);
nor I_95 (I2774,I3015,I3150);
nor I_96 (I2762,I2885,I3150);
not I_97 (I3318,I1634);
DFFARX1 I_98 (I16507,I1627,I3318,I3344,);
not I_99 (I3352,I3344);
nand I_100 (I3369,I16501,I16522);
and I_101 (I3386,I3369,I16498);
DFFARX1 I_102 (I3386,I1627,I3318,I3412,);
DFFARX1 I_103 (I16519,I1627,I3318,I3429,);
and I_104 (I3437,I3429,I16516);
nor I_105 (I3454,I3412,I3437);
DFFARX1 I_106 (I3454,I1627,I3318,I3286,);
nand I_107 (I3485,I3429,I16516);
nand I_108 (I3502,I3352,I3485);
not I_109 (I3298,I3502);
DFFARX1 I_110 (I16504,I1627,I3318,I3542,);
DFFARX1 I_111 (I3542,I1627,I3318,I3307,);
nand I_112 (I3564,I16513,I16510);
and I_113 (I3581,I3564,I16495);
DFFARX1 I_114 (I3581,I1627,I3318,I3607,);
DFFARX1 I_115 (I3607,I1627,I3318,I3624,);
not I_116 (I3310,I3624);
not I_117 (I3646,I3607);
nand I_118 (I3295,I3646,I3485);
nor I_119 (I3677,I16495,I16510);
not I_120 (I3694,I3677);
nor I_121 (I3711,I3646,I3694);
nor I_122 (I3728,I3352,I3711);
DFFARX1 I_123 (I3728,I1627,I3318,I3304,);
nor I_124 (I3759,I3412,I3694);
nor I_125 (I3292,I3607,I3759);
nor I_126 (I3301,I3542,I3677);
nor I_127 (I3289,I3412,I3677);
not I_128 (I3848,I1634);
DFFARX1 I_129 (I2232,I1627,I3848,I3874,);
nand I_130 (I3882,I2256,I2235);
and I_131 (I3899,I3882,I2232);
DFFARX1 I_132 (I3899,I1627,I3848,I3925,);
nor I_133 (I3816,I3925,I3874);
not I_134 (I3947,I3925);
DFFARX1 I_135 (I2238,I1627,I3848,I3973,);
nand I_136 (I3981,I3973,I2247);
not I_137 (I3998,I3981);
DFFARX1 I_138 (I3998,I1627,I3848,I4024,);
not I_139 (I3840,I4024);
nor I_140 (I4046,I3874,I3981);
nor I_141 (I3822,I3925,I4046);
DFFARX1 I_142 (I2241,I1627,I3848,I4086,);
DFFARX1 I_143 (I4086,I1627,I3848,I4103,);
not I_144 (I4111,I4103);
not I_145 (I4128,I4086);
nand I_146 (I3825,I4128,I3947);
nand I_147 (I4159,I2253,I2235);
and I_148 (I4176,I4159,I2244);
DFFARX1 I_149 (I4176,I1627,I3848,I4202,);
nor I_150 (I4210,I4202,I3874);
DFFARX1 I_151 (I4210,I1627,I3848,I3813,);
DFFARX1 I_152 (I4202,I1627,I3848,I3831,);
nor I_153 (I4255,I2250,I2235);
not I_154 (I4272,I4255);
nor I_155 (I3834,I4111,I4272);
nand I_156 (I3819,I4128,I4272);
nor I_157 (I3828,I3874,I4255);
DFFARX1 I_158 (I4255,I1627,I3848,I3837,);
not I_159 (I4375,I1634);
DFFARX1 I_160 (I2762,I1627,I4375,I4401,);
nand I_161 (I4409,I2774,I2783);
and I_162 (I4426,I4409,I2762);
DFFARX1 I_163 (I4426,I1627,I4375,I4452,);
nor I_164 (I4343,I4452,I4401);
not I_165 (I4474,I4452);
DFFARX1 I_166 (I2777,I1627,I4375,I4500,);
nand I_167 (I4508,I4500,I2765);
not I_168 (I4525,I4508);
DFFARX1 I_169 (I4525,I1627,I4375,I4551,);
not I_170 (I4367,I4551);
nor I_171 (I4573,I4401,I4508);
nor I_172 (I4349,I4452,I4573);
DFFARX1 I_173 (I2768,I1627,I4375,I4613,);
DFFARX1 I_174 (I4613,I1627,I4375,I4630,);
not I_175 (I4638,I4630);
not I_176 (I4655,I4613);
nand I_177 (I4352,I4655,I4474);
nand I_178 (I4686,I2759,I2759);
and I_179 (I4703,I4686,I2771);
DFFARX1 I_180 (I4703,I1627,I4375,I4729,);
nor I_181 (I4737,I4729,I4401);
DFFARX1 I_182 (I4737,I1627,I4375,I4340,);
DFFARX1 I_183 (I4729,I1627,I4375,I4358,);
nor I_184 (I4782,I2780,I2759);
not I_185 (I4799,I4782);
nor I_186 (I4361,I4638,I4799);
nand I_187 (I4346,I4655,I4799);
nor I_188 (I4355,I4401,I4782);
DFFARX1 I_189 (I4782,I1627,I4375,I4364,);
not I_190 (I4902,I1634);
DFFARX1 I_191 (I13061,I1627,I4902,I4928,);
nand I_192 (I4936,I13076,I13061);
and I_193 (I4953,I4936,I13079);
DFFARX1 I_194 (I4953,I1627,I4902,I4979,);
nor I_195 (I4870,I4979,I4928);
not I_196 (I5001,I4979);
DFFARX1 I_197 (I13085,I1627,I4902,I5027,);
nand I_198 (I5035,I5027,I13067);
not I_199 (I5052,I5035);
DFFARX1 I_200 (I5052,I1627,I4902,I5078,);
not I_201 (I4894,I5078);
nor I_202 (I5100,I4928,I5035);
nor I_203 (I4876,I4979,I5100);
DFFARX1 I_204 (I13064,I1627,I4902,I5140,);
DFFARX1 I_205 (I5140,I1627,I4902,I5157,);
not I_206 (I5165,I5157);
not I_207 (I5182,I5140);
nand I_208 (I4879,I5182,I5001);
nand I_209 (I5213,I13064,I13070);
and I_210 (I5230,I5213,I13082);
DFFARX1 I_211 (I5230,I1627,I4902,I5256,);
nor I_212 (I5264,I5256,I4928);
DFFARX1 I_213 (I5264,I1627,I4902,I4867,);
DFFARX1 I_214 (I5256,I1627,I4902,I4885,);
nor I_215 (I5309,I13073,I13070);
not I_216 (I5326,I5309);
nor I_217 (I4888,I5165,I5326);
nand I_218 (I4873,I5182,I5326);
nor I_219 (I4882,I4928,I5309);
DFFARX1 I_220 (I5309,I1627,I4902,I4891,);
not I_221 (I5426,I1634);
DFFARX1 I_222 (I4882,I1627,I5426,I5452,);
DFFARX1 I_223 (I5452,I1627,I5426,I5469,);
not I_224 (I5418,I5469);
DFFARX1 I_225 (I4870,I1627,I5426,I5500,);
not I_226 (I5508,I4873);
nor I_227 (I5525,I5452,I5508);
not I_228 (I5542,I4876);
not I_229 (I5559,I4888);
nand I_230 (I5576,I5559,I4876);
nor I_231 (I5593,I5508,I5576);
nor I_232 (I5610,I5500,I5593);
DFFARX1 I_233 (I5559,I1627,I5426,I5415,);
nor I_234 (I5641,I4888,I4879);
nand I_235 (I5658,I5641,I4867);
nor I_236 (I5675,I5658,I5542);
nand I_237 (I5400,I5675,I4873);
DFFARX1 I_238 (I5658,I1627,I5426,I5412,);
nand I_239 (I5720,I5542,I4888);
nor I_240 (I5737,I5542,I4888);
nand I_241 (I5406,I5525,I5737);
not I_242 (I5768,I4885);
nor I_243 (I5785,I5768,I5720);
DFFARX1 I_244 (I5785,I1627,I5426,I5394,);
nor I_245 (I5816,I5768,I4891);
and I_246 (I5833,I5816,I4894);
or I_247 (I5850,I5833,I4867);
DFFARX1 I_248 (I5850,I1627,I5426,I5876,);
nor I_249 (I5884,I5876,I5500);
nor I_250 (I5403,I5452,I5884);
not I_251 (I5915,I5876);
nor I_252 (I5932,I5915,I5610);
DFFARX1 I_253 (I5932,I1627,I5426,I5409,);
nand I_254 (I5963,I5915,I5542);
nor I_255 (I5397,I5768,I5963);
not I_256 (I6021,I1634);
DFFARX1 I_257 (I1444,I1627,I6021,I6047,);
not I_258 (I6055,I6047);
DFFARX1 I_259 (I1532,I1627,I6021,I6081,);
not I_260 (I6089,I1484);
nand I_261 (I6106,I6089,I1588);
not I_262 (I6123,I6106);
nor I_263 (I6140,I6123,I1524);
nor I_264 (I6157,I6055,I6140);
DFFARX1 I_265 (I6157,I1627,I6021,I6007,);
not I_266 (I6188,I1524);
nand I_267 (I6205,I6188,I6123);
and I_268 (I6222,I6188,I1580);
nand I_269 (I6239,I6222,I1420);
nor I_270 (I6004,I6239,I6188);
and I_271 (I5995,I6081,I6239);
not I_272 (I6284,I6239);
nand I_273 (I5998,I6081,I6284);
nor I_274 (I5992,I6047,I6239);
not I_275 (I6329,I1372);
nor I_276 (I6346,I6329,I1580);
nand I_277 (I6363,I6346,I6188);
nor I_278 (I6001,I6106,I6363);
nor I_279 (I6394,I6329,I1380);
and I_280 (I6411,I6394,I1428);
or I_281 (I6428,I6411,I1436);
DFFARX1 I_282 (I6428,I1627,I6021,I6454,);
nor I_283 (I6462,I6454,I6205);
DFFARX1 I_284 (I6462,I1627,I6021,I5989,);
DFFARX1 I_285 (I6454,I1627,I6021,I6013,);
not I_286 (I6507,I6454);
nor I_287 (I6524,I6507,I6081);
nor I_288 (I6541,I6346,I6524);
DFFARX1 I_289 (I6541,I1627,I6021,I6010,);
not I_290 (I6599,I1634);
DFFARX1 I_291 (I8879,I1627,I6599,I6625,);
not I_292 (I6633,I6625);
DFFARX1 I_293 (I8891,I1627,I6599,I6659,);
not I_294 (I6667,I8882);
nand I_295 (I6684,I6667,I8885);
not I_296 (I6701,I6684);
nor I_297 (I6718,I6701,I8888);
nor I_298 (I6735,I6633,I6718);
DFFARX1 I_299 (I6735,I1627,I6599,I6585,);
not I_300 (I6766,I8888);
nand I_301 (I6783,I6766,I6701);
and I_302 (I6800,I6766,I8882);
nand I_303 (I6817,I6800,I8894);
nor I_304 (I6582,I6817,I6766);
and I_305 (I6573,I6659,I6817);
not I_306 (I6862,I6817);
nand I_307 (I6576,I6659,I6862);
nor I_308 (I6570,I6625,I6817);
not I_309 (I6907,I8900);
nor I_310 (I6924,I6907,I8882);
nand I_311 (I6941,I6924,I6766);
nor I_312 (I6579,I6684,I6941);
nor I_313 (I6972,I6907,I8879);
and I_314 (I6989,I6972,I8897);
or I_315 (I7006,I6989,I8903);
DFFARX1 I_316 (I7006,I1627,I6599,I7032,);
nor I_317 (I7040,I7032,I6783);
DFFARX1 I_318 (I7040,I1627,I6599,I6567,);
DFFARX1 I_319 (I7032,I1627,I6599,I6591,);
not I_320 (I7085,I7032);
nor I_321 (I7102,I7085,I6659);
nor I_322 (I7119,I6924,I7102);
DFFARX1 I_323 (I7119,I1627,I6599,I6588,);
not I_324 (I7177,I1634);
DFFARX1 I_325 (I11282,I1627,I7177,I7203,);
not I_326 (I7211,I7203);
DFFARX1 I_327 (I11279,I1627,I7177,I7237,);
not I_328 (I7245,I11276);
nand I_329 (I7262,I7245,I11303);
not I_330 (I7279,I7262);
nor I_331 (I7296,I7279,I11291);
nor I_332 (I7313,I7211,I7296);
DFFARX1 I_333 (I7313,I1627,I7177,I7163,);
not I_334 (I7344,I11291);
nand I_335 (I7361,I7344,I7279);
and I_336 (I7378,I7344,I11297);
nand I_337 (I7395,I7378,I11288);
nor I_338 (I7160,I7395,I7344);
and I_339 (I7151,I7237,I7395);
not I_340 (I7440,I7395);
nand I_341 (I7154,I7237,I7440);
nor I_342 (I7148,I7203,I7395);
not I_343 (I7485,I11285);
nor I_344 (I7502,I7485,I11297);
nand I_345 (I7519,I7502,I7344);
nor I_346 (I7157,I7262,I7519);
nor I_347 (I7550,I7485,I11300);
and I_348 (I7567,I7550,I11294);
or I_349 (I7584,I7567,I11276);
DFFARX1 I_350 (I7584,I1627,I7177,I7610,);
nor I_351 (I7618,I7610,I7361);
DFFARX1 I_352 (I7618,I1627,I7177,I7145,);
DFFARX1 I_353 (I7610,I1627,I7177,I7169,);
not I_354 (I7663,I7610);
nor I_355 (I7680,I7663,I7237);
nor I_356 (I7697,I7502,I7680);
DFFARX1 I_357 (I7697,I1627,I7177,I7166,);
not I_358 (I7755,I1634);
DFFARX1 I_359 (I11928,I1627,I7755,I7781,);
not I_360 (I7789,I7781);
nand I_361 (I7806,I11925,I11943);
and I_362 (I7823,I7806,I11940);
DFFARX1 I_363 (I7823,I1627,I7755,I7849,);
not I_364 (I7857,I11922);
DFFARX1 I_365 (I11925,I1627,I7755,I7883,);
not I_366 (I7891,I7883);
nor I_367 (I7908,I7891,I7789);
and I_368 (I7925,I7908,I11922);
nor I_369 (I7942,I7891,I7857);
nor I_370 (I7738,I7849,I7942);
DFFARX1 I_371 (I11934,I1627,I7755,I7982,);
nor I_372 (I7990,I7982,I7849);
not I_373 (I8007,I7990);
not I_374 (I8024,I7982);
nor I_375 (I8041,I8024,I7925);
DFFARX1 I_376 (I8041,I1627,I7755,I7741,);
nand I_377 (I8072,I11937,I11922);
and I_378 (I8089,I8072,I11928);
DFFARX1 I_379 (I8089,I1627,I7755,I8115,);
nor I_380 (I8123,I8115,I7982);
DFFARX1 I_381 (I8123,I1627,I7755,I7723,);
nand I_382 (I8154,I8115,I8024);
nand I_383 (I7732,I8007,I8154);
not I_384 (I8185,I8115);
nor I_385 (I8202,I8185,I7925);
DFFARX1 I_386 (I8202,I1627,I7755,I7744,);
nor I_387 (I8233,I11931,I11922);
or I_388 (I7735,I7982,I8233);
nor I_389 (I7726,I8115,I8233);
or I_390 (I7729,I7849,I8233);
DFFARX1 I_391 (I8233,I1627,I7755,I7747,);
not I_392 (I8333,I1634);
DFFARX1 I_393 (I14235,I1627,I8333,I8359,);
not I_394 (I8367,I8359);
nand I_395 (I8384,I14217,I14229);
and I_396 (I8401,I8384,I14232);
DFFARX1 I_397 (I8401,I1627,I8333,I8427,);
not I_398 (I8435,I14226);
DFFARX1 I_399 (I14223,I1627,I8333,I8461,);
not I_400 (I8469,I8461);
nor I_401 (I8486,I8469,I8367);
and I_402 (I8503,I8486,I14226);
nor I_403 (I8520,I8469,I8435);
nor I_404 (I8316,I8427,I8520);
DFFARX1 I_405 (I14241,I1627,I8333,I8560,);
nor I_406 (I8568,I8560,I8427);
not I_407 (I8585,I8568);
not I_408 (I8602,I8560);
nor I_409 (I8619,I8602,I8503);
DFFARX1 I_410 (I8619,I1627,I8333,I8319,);
nand I_411 (I8650,I14220,I14220);
and I_412 (I8667,I8650,I14217);
DFFARX1 I_413 (I8667,I1627,I8333,I8693,);
nor I_414 (I8701,I8693,I8560);
DFFARX1 I_415 (I8701,I1627,I8333,I8301,);
nand I_416 (I8732,I8693,I8602);
nand I_417 (I8310,I8585,I8732);
not I_418 (I8763,I8693);
nor I_419 (I8780,I8763,I8503);
DFFARX1 I_420 (I8780,I1627,I8333,I8322,);
nor I_421 (I8811,I14238,I14220);
or I_422 (I8313,I8560,I8811);
nor I_423 (I8304,I8693,I8811);
or I_424 (I8307,I8427,I8811);
DFFARX1 I_425 (I8811,I1627,I8333,I8325,);
not I_426 (I8911,I1634);
DFFARX1 I_427 (I1460,I1627,I8911,I8937,);
not I_428 (I8945,I8937);
nand I_429 (I8962,I1612,I1516);
and I_430 (I8979,I8962,I1476);
DFFARX1 I_431 (I8979,I1627,I8911,I9005,);
not I_432 (I9013,I1540);
DFFARX1 I_433 (I1364,I1627,I8911,I9039,);
not I_434 (I9047,I9039);
nor I_435 (I9064,I9047,I8945);
and I_436 (I9081,I9064,I1540);
nor I_437 (I9098,I9047,I9013);
nor I_438 (I8894,I9005,I9098);
DFFARX1 I_439 (I1396,I1627,I8911,I9138,);
nor I_440 (I9146,I9138,I9005);
not I_441 (I9163,I9146);
not I_442 (I9180,I9138);
nor I_443 (I9197,I9180,I9081);
DFFARX1 I_444 (I9197,I1627,I8911,I8897,);
nand I_445 (I9228,I1548,I1620);
and I_446 (I9245,I9228,I1572);
DFFARX1 I_447 (I9245,I1627,I8911,I9271,);
nor I_448 (I9279,I9271,I9138);
DFFARX1 I_449 (I9279,I1627,I8911,I8879,);
nand I_450 (I9310,I9271,I9180);
nand I_451 (I8888,I9163,I9310);
not I_452 (I9341,I9271);
nor I_453 (I9358,I9341,I9081);
DFFARX1 I_454 (I9358,I1627,I8911,I8900,);
nor I_455 (I9389,I1452,I1620);
or I_456 (I8891,I9138,I9389);
nor I_457 (I8882,I9271,I9389);
or I_458 (I8885,I9005,I9389);
DFFARX1 I_459 (I9389,I1627,I8911,I8903,);
not I_460 (I9486,I1634);
DFFARX1 I_461 (I3310,I1627,I9486,I9512,);
not I_462 (I9520,I9512);
nand I_463 (I9537,I3286,I3295);
and I_464 (I9554,I9537,I3289);
DFFARX1 I_465 (I9554,I1627,I9486,I9580,);
DFFARX1 I_466 (I9580,I1627,I9486,I9475,);
DFFARX1 I_467 (I3307,I1627,I9486,I9611,);
nand I_468 (I9619,I9611,I3298);
not I_469 (I9636,I9619);
DFFARX1 I_470 (I9636,I1627,I9486,I9662,);
not I_471 (I9670,I9662);
nor I_472 (I9478,I9520,I9670);
DFFARX1 I_473 (I3292,I1627,I9486,I9710,);
nor I_474 (I9469,I9710,I9580);
nor I_475 (I9460,I9710,I9636);
nand I_476 (I9746,I3304,I3301);
and I_477 (I9763,I9746,I3289);
DFFARX1 I_478 (I9763,I1627,I9486,I9789,);
not I_479 (I9797,I9789);
nand I_480 (I9814,I9797,I9710);
nand I_481 (I9463,I9797,I9619);
nor I_482 (I9845,I3286,I3301);
and I_483 (I9862,I9710,I9845);
nor I_484 (I9879,I9797,I9862);
DFFARX1 I_485 (I9879,I1627,I9486,I9472,);
nor I_486 (I9910,I9512,I9845);
DFFARX1 I_487 (I9910,I1627,I9486,I9457,);
nor I_488 (I9941,I9789,I9845);
not I_489 (I9958,I9941);
nand I_490 (I9466,I9958,I9814);
not I_491 (I10019,I1634);
DFFARX1 I_492 (I8307,I1627,I10019,I10045,);
DFFARX1 I_493 (I8301,I1627,I10019,I10062,);
not I_494 (I10070,I10062);
not I_495 (I10087,I8316);
nor I_496 (I10104,I10087,I8301);
not I_497 (I10121,I8310);
nor I_498 (I10138,I10104,I8319);
nor I_499 (I10155,I10062,I10138);
DFFARX1 I_500 (I10155,I1627,I10019,I10005,);
nor I_501 (I10186,I8319,I8301);
nand I_502 (I10203,I10186,I8316);
DFFARX1 I_503 (I10203,I1627,I10019,I10008,);
nor I_504 (I10234,I10121,I8319);
nand I_505 (I10251,I10234,I8304);
nor I_506 (I10268,I10045,I10251);
DFFARX1 I_507 (I10268,I1627,I10019,I9984,);
not I_508 (I10299,I10251);
nand I_509 (I9996,I10062,I10299);
DFFARX1 I_510 (I10251,I1627,I10019,I10339,);
not I_511 (I10347,I10339);
not I_512 (I10364,I8319);
not I_513 (I10381,I8313);
nor I_514 (I10398,I10381,I8310);
nor I_515 (I10011,I10347,I10398);
nor I_516 (I10429,I10381,I8322);
and I_517 (I10446,I10429,I8325);
or I_518 (I10463,I10446,I8304);
DFFARX1 I_519 (I10463,I1627,I10019,I10489,);
nor I_520 (I9999,I10489,I10045);
not I_521 (I10511,I10489);
and I_522 (I10528,I10511,I10045);
nor I_523 (I9993,I10070,I10528);
nand I_524 (I10559,I10511,I10121);
nor I_525 (I9987,I10381,I10559);
nand I_526 (I9990,I10511,I10299);
nand I_527 (I10604,I10121,I8313);
nor I_528 (I10002,I10364,I10604);
not I_529 (I10665,I1634);
DFFARX1 I_530 (I12501,I1627,I10665,I10691,);
DFFARX1 I_531 (I12483,I1627,I10665,I10708,);
not I_532 (I10716,I10708);
not I_533 (I10733,I12492);
nor I_534 (I10750,I10733,I12504);
not I_535 (I10767,I12486);
nor I_536 (I10784,I10750,I12495);
nor I_537 (I10801,I10708,I10784);
DFFARX1 I_538 (I10801,I1627,I10665,I10651,);
nor I_539 (I10832,I12495,I12504);
nand I_540 (I10849,I10832,I12492);
DFFARX1 I_541 (I10849,I1627,I10665,I10654,);
nor I_542 (I10880,I10767,I12495);
nand I_543 (I10897,I10880,I12507);
nor I_544 (I10914,I10691,I10897);
DFFARX1 I_545 (I10914,I1627,I10665,I10630,);
not I_546 (I10945,I10897);
nand I_547 (I10642,I10708,I10945);
DFFARX1 I_548 (I10897,I1627,I10665,I10985,);
not I_549 (I10993,I10985);
not I_550 (I11010,I12495);
not I_551 (I11027,I12483);
nor I_552 (I11044,I11027,I12486);
nor I_553 (I10657,I10993,I11044);
nor I_554 (I11075,I11027,I12489);
and I_555 (I11092,I11075,I12498);
or I_556 (I11109,I11092,I12486);
DFFARX1 I_557 (I11109,I1627,I10665,I11135,);
nor I_558 (I10645,I11135,I10691);
not I_559 (I11157,I11135);
and I_560 (I11174,I11157,I10691);
nor I_561 (I10639,I10716,I11174);
nand I_562 (I11205,I11157,I10767);
nor I_563 (I10633,I11027,I11205);
nand I_564 (I10636,I11157,I10945);
nand I_565 (I11250,I10767,I12483);
nor I_566 (I10648,I11010,I11250);
not I_567 (I11311,I1634);
DFFARX1 I_568 (I3813,I1627,I11311,I11337,);
DFFARX1 I_569 (I3819,I1627,I11311,I11354,);
not I_570 (I11362,I11354);
not I_571 (I11379,I3840);
nor I_572 (I11396,I11379,I3828);
not I_573 (I11413,I3837);
nor I_574 (I11430,I11396,I3822);
nor I_575 (I11447,I11354,I11430);
DFFARX1 I_576 (I11447,I1627,I11311,I11297,);
nor I_577 (I11478,I3822,I3828);
nand I_578 (I11495,I11478,I3840);
DFFARX1 I_579 (I11495,I1627,I11311,I11300,);
nor I_580 (I11526,I11413,I3822);
nand I_581 (I11543,I11526,I3813);
nor I_582 (I11560,I11337,I11543);
DFFARX1 I_583 (I11560,I1627,I11311,I11276,);
not I_584 (I11591,I11543);
nand I_585 (I11288,I11354,I11591);
DFFARX1 I_586 (I11543,I1627,I11311,I11631,);
not I_587 (I11639,I11631);
not I_588 (I11656,I3822);
not I_589 (I11673,I3825);
nor I_590 (I11690,I11673,I3837);
nor I_591 (I11303,I11639,I11690);
nor I_592 (I11721,I11673,I3834);
and I_593 (I11738,I11721,I3816);
or I_594 (I11755,I11738,I3831);
DFFARX1 I_595 (I11755,I1627,I11311,I11781,);
nor I_596 (I11291,I11781,I11337);
not I_597 (I11803,I11781);
and I_598 (I11820,I11803,I11337);
nor I_599 (I11285,I11362,I11820);
nand I_600 (I11851,I11803,I11413);
nor I_601 (I11279,I11673,I11851);
nand I_602 (I11282,I11803,I11591);
nand I_603 (I11896,I11413,I3825);
nor I_604 (I11294,I11656,I11896);
not I_605 (I11951,I1634);
DFFARX1 I_606 (I5989,I1627,I11951,I11977,);
DFFARX1 I_607 (I11977,I1627,I11951,I11994,);
not I_608 (I11943,I11994);
not I_609 (I12016,I11977);
DFFARX1 I_610 (I6004,I1627,I11951,I12042,);
nand I_611 (I12050,I12042,I5995);
not I_612 (I12067,I5995);
not I_613 (I12084,I6001);
nand I_614 (I12101,I5998,I6007);
and I_615 (I12118,I5998,I6007);
not I_616 (I12135,I5992);
nand I_617 (I12152,I12135,I12084);
nor I_618 (I11925,I12152,I12050);
nor I_619 (I12183,I12067,I12152);
nand I_620 (I11928,I12118,I12183);
not I_621 (I12214,I5989);
nor I_622 (I12231,I12214,I5998);
nor I_623 (I12248,I12231,I5992);
nor I_624 (I12265,I12016,I12248);
DFFARX1 I_625 (I12265,I1627,I11951,I11937,);
not I_626 (I12296,I12231);
DFFARX1 I_627 (I12296,I1627,I11951,I11940,);
and I_628 (I11934,I12042,I12231);
nor I_629 (I12341,I12214,I6013);
and I_630 (I12358,I12341,I5992);
or I_631 (I12375,I12358,I6010);
DFFARX1 I_632 (I12375,I1627,I11951,I12401,);
nor I_633 (I12409,I12401,I12135);
DFFARX1 I_634 (I12409,I1627,I11951,I11922,);
nand I_635 (I12440,I12401,I12042);
nand I_636 (I12457,I12135,I12440);
nor I_637 (I11931,I12457,I12101);
not I_638 (I12515,I1634);
DFFARX1 I_639 (I1652,I1627,I12515,I12541,);
and I_640 (I12549,I12541,I1658);
DFFARX1 I_641 (I12549,I1627,I12515,I12498,);
DFFARX1 I_642 (I1637,I1627,I12515,I12589,);
not I_643 (I12597,I1643);
not I_644 (I12614,I1649);
nand I_645 (I12631,I12614,I12597);
nor I_646 (I12486,I12589,I12631);
DFFARX1 I_647 (I12631,I1627,I12515,I12671,);
not I_648 (I12507,I12671);
not I_649 (I12693,I1640);
nand I_650 (I12710,I12614,I12693);
DFFARX1 I_651 (I12710,I1627,I12515,I12736,);
not I_652 (I12744,I12736);
not I_653 (I12761,I1655);
nand I_654 (I12778,I12761,I1640);
and I_655 (I12795,I12597,I12778);
nor I_656 (I12812,I12710,I12795);
DFFARX1 I_657 (I12812,I1627,I12515,I12483,);
DFFARX1 I_658 (I12795,I1627,I12515,I12504,);
nor I_659 (I12857,I1655,I1643);
nor I_660 (I12495,I12710,I12857);
or I_661 (I12888,I1655,I1643);
nor I_662 (I12905,I1646,I1637);
DFFARX1 I_663 (I12905,I1627,I12515,I12931,);
not I_664 (I12939,I12931);
nor I_665 (I12501,I12939,I12744);
nand I_666 (I12970,I12939,I12589);
not I_667 (I12987,I1646);
nand I_668 (I13004,I12987,I12693);
nand I_669 (I13021,I12939,I13004);
nand I_670 (I12492,I13021,I12970);
nand I_671 (I12489,I13004,I12888);
not I_672 (I13093,I1634);
DFFARX1 I_673 (I9460,I1627,I13093,I13119,);
and I_674 (I13127,I13119,I9466);
DFFARX1 I_675 (I13127,I1627,I13093,I13076,);
DFFARX1 I_676 (I9472,I1627,I13093,I13167,);
not I_677 (I13175,I9457);
not I_678 (I13192,I9457);
nand I_679 (I13209,I13192,I13175);
nor I_680 (I13064,I13167,I13209);
DFFARX1 I_681 (I13209,I1627,I13093,I13249,);
not I_682 (I13085,I13249);
not I_683 (I13271,I9475);
nand I_684 (I13288,I13192,I13271);
DFFARX1 I_685 (I13288,I1627,I13093,I13314,);
not I_686 (I13322,I13314);
not I_687 (I13339,I9469);
nand I_688 (I13356,I13339,I9460);
and I_689 (I13373,I13175,I13356);
nor I_690 (I13390,I13288,I13373);
DFFARX1 I_691 (I13390,I1627,I13093,I13061,);
DFFARX1 I_692 (I13373,I1627,I13093,I13082,);
nor I_693 (I13435,I9469,I9478);
nor I_694 (I13073,I13288,I13435);
or I_695 (I13466,I9469,I9478);
nor I_696 (I13483,I9463,I9463);
DFFARX1 I_697 (I13483,I1627,I13093,I13509,);
not I_698 (I13517,I13509);
nor I_699 (I13079,I13517,I13322);
nand I_700 (I13548,I13517,I13167);
not I_701 (I13565,I9463);
nand I_702 (I13582,I13565,I13271);
nand I_703 (I13599,I13517,I13582);
nand I_704 (I13070,I13599,I13548);
nand I_705 (I13067,I13582,I13466);
not I_706 (I13671,I1634);
DFFARX1 I_707 (I6582,I1627,I13671,I13697,);
and I_708 (I13705,I13697,I6570);
DFFARX1 I_709 (I13705,I1627,I13671,I13654,);
DFFARX1 I_710 (I6585,I1627,I13671,I13745,);
not I_711 (I13753,I6576);
not I_712 (I13770,I6567);
nand I_713 (I13787,I13770,I13753);
nor I_714 (I13642,I13745,I13787);
DFFARX1 I_715 (I13787,I1627,I13671,I13827,);
not I_716 (I13663,I13827);
not I_717 (I13849,I6573);
nand I_718 (I13866,I13770,I13849);
DFFARX1 I_719 (I13866,I1627,I13671,I13892,);
not I_720 (I13900,I13892);
not I_721 (I13917,I6588);
nand I_722 (I13934,I13917,I6591);
and I_723 (I13951,I13753,I13934);
nor I_724 (I13968,I13866,I13951);
DFFARX1 I_725 (I13968,I1627,I13671,I13639,);
DFFARX1 I_726 (I13951,I1627,I13671,I13660,);
nor I_727 (I14013,I6588,I6567);
nor I_728 (I13651,I13866,I14013);
or I_729 (I14044,I6588,I6567);
nor I_730 (I14061,I6579,I6570);
DFFARX1 I_731 (I14061,I1627,I13671,I14087,);
not I_732 (I14095,I14087);
nor I_733 (I13657,I14095,I13900);
nand I_734 (I14126,I14095,I13745);
not I_735 (I14143,I6579);
nand I_736 (I14160,I14143,I13849);
nand I_737 (I14177,I14095,I14160);
nand I_738 (I13648,I14177,I14126);
nand I_739 (I13645,I14160,I14044);
not I_740 (I14249,I1634);
DFFARX1 I_741 (I4367,I1627,I14249,I14275,);
and I_742 (I14283,I14275,I4352);
DFFARX1 I_743 (I14283,I1627,I14249,I14232,);
DFFARX1 I_744 (I4358,I1627,I14249,I14323,);
not I_745 (I14331,I4340);
not I_746 (I14348,I4361);
nand I_747 (I14365,I14348,I14331);
nor I_748 (I14220,I14323,I14365);
DFFARX1 I_749 (I14365,I1627,I14249,I14405,);
not I_750 (I14241,I14405);
not I_751 (I14427,I4364);
nand I_752 (I14444,I14348,I14427);
DFFARX1 I_753 (I14444,I1627,I14249,I14470,);
not I_754 (I14478,I14470);
not I_755 (I14495,I4355);
nand I_756 (I14512,I14495,I4343);
and I_757 (I14529,I14331,I14512);
nor I_758 (I14546,I14444,I14529);
DFFARX1 I_759 (I14546,I1627,I14249,I14217,);
DFFARX1 I_760 (I14529,I1627,I14249,I14238,);
nor I_761 (I14591,I4355,I4349);
nor I_762 (I14229,I14444,I14591);
or I_763 (I14622,I4355,I4349);
nor I_764 (I14639,I4346,I4340);
DFFARX1 I_765 (I14639,I1627,I14249,I14665,);
not I_766 (I14673,I14665);
nor I_767 (I14235,I14673,I14478);
nand I_768 (I14704,I14673,I14323);
not I_769 (I14721,I4346);
nand I_770 (I14738,I14721,I14427);
nand I_771 (I14755,I14673,I14738);
nand I_772 (I14226,I14755,I14704);
nand I_773 (I14223,I14738,I14622);
not I_774 (I14827,I1634);
DFFARX1 I_775 (I7160,I1627,I14827,I14853,);
and I_776 (I14861,I14853,I7148);
DFFARX1 I_777 (I14861,I1627,I14827,I14810,);
DFFARX1 I_778 (I7163,I1627,I14827,I14901,);
not I_779 (I14909,I7154);
not I_780 (I14926,I7145);
nand I_781 (I14943,I14926,I14909);
nor I_782 (I14798,I14901,I14943);
DFFARX1 I_783 (I14943,I1627,I14827,I14983,);
not I_784 (I14819,I14983);
not I_785 (I15005,I7151);
nand I_786 (I15022,I14926,I15005);
DFFARX1 I_787 (I15022,I1627,I14827,I15048,);
not I_788 (I15056,I15048);
not I_789 (I15073,I7166);
nand I_790 (I15090,I15073,I7169);
and I_791 (I15107,I14909,I15090);
nor I_792 (I15124,I15022,I15107);
DFFARX1 I_793 (I15124,I1627,I14827,I14795,);
DFFARX1 I_794 (I15107,I1627,I14827,I14816,);
nor I_795 (I15169,I7166,I7145);
nor I_796 (I14807,I15022,I15169);
or I_797 (I15200,I7166,I7145);
nor I_798 (I15217,I7157,I7148);
DFFARX1 I_799 (I15217,I1627,I14827,I15243,);
not I_800 (I15251,I15243);
nor I_801 (I14813,I15251,I15056);
nand I_802 (I15282,I15251,I14901);
not I_803 (I15299,I7157);
nand I_804 (I15316,I15299,I15005);
nand I_805 (I15333,I15251,I15316);
nand I_806 (I14804,I15333,I15282);
nand I_807 (I14801,I15316,I15200);
not I_808 (I15405,I1634);
DFFARX1 I_809 (I9984,I1627,I15405,I15431,);
nand I_810 (I15439,I15431,I9984);
DFFARX1 I_811 (I9996,I1627,I15405,I15465,);
DFFARX1 I_812 (I15465,I1627,I15405,I15482,);
not I_813 (I15397,I15482);
not I_814 (I15504,I9990);
nor I_815 (I15521,I9990,I10011);
not I_816 (I15538,I9999);
nand I_817 (I15555,I15504,I15538);
nor I_818 (I15572,I9999,I9990);
and I_819 (I15376,I15572,I15439);
not I_820 (I15603,I9993);
nand I_821 (I15620,I15603,I10008);
nor I_822 (I15637,I9993,I10002);
not I_823 (I15654,I15637);
nand I_824 (I15379,I15521,I15654);
DFFARX1 I_825 (I15637,I1627,I15405,I15394,);
nor I_826 (I15699,I10005,I9999);
nor I_827 (I15716,I15699,I10011);
and I_828 (I15733,I15716,I15620);
DFFARX1 I_829 (I15733,I1627,I15405,I15391,);
nor I_830 (I15388,I15699,I15555);
or I_831 (I15385,I15637,I15699);
nor I_832 (I15792,I10005,I9987);
DFFARX1 I_833 (I15792,I1627,I15405,I15818,);
not I_834 (I15826,I15818);
nand I_835 (I15843,I15826,I15504);
nor I_836 (I15860,I15843,I10011);
DFFARX1 I_837 (I15860,I1627,I15405,I15373,);
nor I_838 (I15891,I15826,I15555);
nor I_839 (I15382,I15699,I15891);
not I_840 (I15949,I1634);
DFFARX1 I_841 (I14813,I1627,I15949,I15975,);
nand I_842 (I15983,I15975,I14798);
not I_843 (I16000,I15983);
DFFARX1 I_844 (I14801,I1627,I15949,I16026,);
not I_845 (I16034,I16026);
not I_846 (I16051,I14816);
or I_847 (I16068,I14819,I14816);
nor I_848 (I16085,I14819,I14816);
or I_849 (I16102,I14795,I14819);
DFFARX1 I_850 (I16102,I1627,I15949,I15941,);
not I_851 (I16133,I14807);
nand I_852 (I16150,I16133,I14810);
nand I_853 (I16167,I16051,I16150);
and I_854 (I15920,I16034,I16167);
nor I_855 (I16198,I14807,I14804);
and I_856 (I16215,I16034,I16198);
nor I_857 (I15926,I16000,I16215);
DFFARX1 I_858 (I16198,I1627,I15949,I16255,);
not I_859 (I16263,I16255);
nor I_860 (I15935,I16034,I16263);
or I_861 (I16294,I16102,I14795);
nor I_862 (I16311,I14795,I14795);
nand I_863 (I16328,I16167,I16311);
nand I_864 (I16345,I16294,I16328);
DFFARX1 I_865 (I16345,I1627,I15949,I15938,);
nor I_866 (I16376,I16311,I16068);
DFFARX1 I_867 (I16376,I1627,I15949,I15917,);
nor I_868 (I16407,I14795,I14798);
DFFARX1 I_869 (I16407,I1627,I15949,I16433,);
DFFARX1 I_870 (I16433,I1627,I15949,I15932,);
not I_871 (I16455,I16433);
nand I_872 (I15929,I16455,I15983);
nand I_873 (I15923,I16455,I16085);
not I_874 (I16530,I1634);
DFFARX1 I_875 (I7744,I1627,I16530,I16556,);
DFFARX1 I_876 (I7726,I1627,I16530,I16573,);
not I_877 (I16581,I16573);
nor I_878 (I16498,I16556,I16581);
DFFARX1 I_879 (I16581,I1627,I16530,I16513,);
nor I_880 (I16626,I7732,I7735);
and I_881 (I16643,I16626,I7723);
nor I_882 (I16660,I16643,I7732);
not I_883 (I16677,I7732);
and I_884 (I16694,I16677,I7741);
nand I_885 (I16711,I16694,I7729);
nor I_886 (I16728,I16677,I16711);
DFFARX1 I_887 (I16728,I1627,I16530,I16495,);
not I_888 (I16759,I16711);
nand I_889 (I16776,I16581,I16759);
nand I_890 (I16507,I16643,I16759);
DFFARX1 I_891 (I16677,I1627,I16530,I16522,);
not I_892 (I16821,I7726);
nor I_893 (I16838,I16821,I7741);
nor I_894 (I16855,I16838,I16660);
DFFARX1 I_895 (I16855,I1627,I16530,I16519,);
not I_896 (I16886,I16838);
DFFARX1 I_897 (I16886,I1627,I16530,I16912,);
not I_898 (I16920,I16912);
nor I_899 (I16516,I16920,I16838);
nor I_900 (I16951,I16821,I7738);
and I_901 (I16968,I16951,I7747);
or I_902 (I16985,I16968,I7723);
DFFARX1 I_903 (I16985,I1627,I16530,I17011,);
not I_904 (I17019,I17011);
nand I_905 (I17036,I17019,I16759);
not I_906 (I16510,I17036);
nand I_907 (I16504,I17036,I16776);
nand I_908 (I16501,I17019,I16643);
endmodule


