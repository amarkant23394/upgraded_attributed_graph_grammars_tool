module test_final(G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input G1_0_l_8,G2_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_5_0_l_8,IN_7_0_l_8,IN_8_0_l_8,IN_10_0_l_8,IN_11_0_l_8,IN_1_5_l_8,IN_2_5_l_8,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8,n_431_0_l_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n4_1_r_8,blif_clk_net_1_r_1,n5_1,G42_1_r_8,);
nor I_1(n_572_1_r_8,n39_8,n23_8);
and I_2(n_549_1_r_8,n38_8,n23_8);
nand I_3(n_569_1_r_8,n38_8,n24_8);
nor I_4(n_452_1_r_8,n25_8,n26_8);
nor I_5(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_6(N3_2_r_8,blif_clk_net_1_r_1,n5_1,G199_2_r_8,);
DFFARX1 I_7(N1_4_r_8,blif_clk_net_1_r_1,n5_1,G199_4_r_8,);
DFFARX1 I_8(G78_0_l_8,blif_clk_net_1_r_1,n5_1,G214_4_r_8,);
or I_9(n_431_0_l_8,IN_8_0_l_8,n29_8);
DFFARX1 I_10(n_431_0_l_8,blif_clk_net_1_r_1,n5_1,G78_0_l_8,);
not I_11(n19_8,G78_0_l_8);
DFFARX1 I_12(IN_2_5_l_8,blif_clk_net_1_r_1,n5_1,n39_8,);
not I_13(n22_8,n39_8);
DFFARX1 I_14(IN_1_5_l_8,blif_clk_net_1_r_1,n5_1,n38_8,);
nor I_15(n4_1_r_8,G78_0_l_8,n33_8);
nor I_16(N3_2_r_8,n22_8,n35_8);
nor I_17(N1_4_r_8,n27_8,n37_8);
nand I_18(n23_8,IN_7_0_l_8,n32_8);
not I_19(n24_8,n23_8);
nand I_20(n25_8,IN_11_0_l_8,n36_8);
nand I_21(n26_8,n27_8,n28_8);
nor I_22(n27_8,IN_5_0_l_8,n31_8);
not I_23(n28_8,G2_0_l_8);
and I_24(n29_8,IN_2_0_l_8,n30_8);
nor I_25(n30_8,IN_4_0_l_8,n31_8);
not I_26(n31_8,G1_0_l_8);
and I_27(n32_8,IN_5_0_l_8,n28_8);
nand I_28(n33_8,n28_8,n34_8);
not I_29(n34_8,n25_8);
nor I_30(n35_8,G2_0_l_8,n34_8);
not I_31(n36_8,IN_10_0_l_8);
nor I_32(n37_8,n19_8,n38_8);
DFFARX1 I_33(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_34(n_572_1_r_1,n26_1,n19_1);
nand I_35(n_573_1_r_1,n16_1,n18_1);
nor I_36(n_549_1_r_1,n20_1,n21_1);
nor I_37(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_38(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_39(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_40(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_41(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_42(N3_2_l_1,n23_1,n_549_1_r_8);
not I_43(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_44(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_45(n17_1,n26_1);
DFFARX1 I_46(n_452_1_r_8,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_47(n16_1,n16_internal_1);
DFFARX1 I_48(G199_2_r_8,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_49(N1_4_l_1,n25_1,G42_1_r_8);
DFFARX1 I_50(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_51(G214_4_r_8,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_52(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_53(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_54(n14_1,n14_internal_1);
nor I_55(N1_4_r_1,n17_1,n24_1);
nand I_56(n18_1,ACVQN1_3_l_1,G199_4_r_8);
nor I_57(n19_1,n_572_1_r_8,n_42_2_r_8);
not I_58(n20_1,n18_1);
nor I_59(n21_1,n26_1,n22_1);
not I_60(n22_1,n19_1);
nand I_61(n23_1,n_572_1_r_8,n_569_1_r_8);
nor I_62(n24_1,n18_1,n22_1);
nand I_63(n25_1,G42_1_r_8,n_572_1_r_8);
endmodule


