module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_7_r_12,n8_12,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_7_r_12,n8_12,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
nor I_37(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_38(N1508_0_r_12,n30_12,n37_12);
nor I_39(N1507_6_r_12,n25_12,n39_12);
nor I_40(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_41(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_42(n_572_7_r_12,n23_12,n24_12);
nand I_43(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_44(n_549_7_r_12,n27_12,n28_12);
nand I_45(n_569_7_r_12,n25_12,n26_12);
nand I_46(n_452_7_r_12,n_572_7_r_14,n_452_7_r_14);
nand I_47(N6147_9_r_12,n30_12,n31_12);
nor I_48(N6134_9_r_12,n35_12,n36_12);
not I_49(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_50(n1_12,n_573_7_r_12);
not I_51(n8_12,blif_reset_net_7_r_12);
not I_52(n23_12,n36_12);
nor I_53(n24_12,n_452_7_r_12,n_573_7_r_14);
nand I_54(n25_12,n23_12,n40_12);
not I_55(n26_12,n35_12);
not I_56(n27_12,N6134_9_r_12);
nand I_57(n28_12,n26_12,n29_12);
not I_58(n29_12,n24_12);
nand I_59(n30_12,n33_12,n41_12);
nand I_60(n31_12,n32_12,n33_12);
nor I_61(n32_12,n26_12,n34_12);
nor I_62(n33_12,N1508_0_r_14,N1507_6_r_14);
nor I_63(n34_12,n42_12,n_549_7_r_14);
nor I_64(n35_12,n38_12,N6134_9_r_14);
nand I_65(n36_12,N6147_9_r_14,N1371_0_r_14);
nand I_66(n37_12,n23_12,n35_12);
or I_67(n38_12,N1371_0_r_14,N1507_6_r_14);
not I_68(n39_12,n30_12);
or I_69(n40_12,N1508_6_r_14,n_569_7_r_14);
nor I_70(n41_12,n34_12,n36_12);
nor I_71(n42_12,N1508_0_r_14,G42_7_r_14);
endmodule


