module test_I11864(I1477,I9148,I8913,I9083,I1470,I11864);
input I1477,I9148,I8913,I9083,I1470;
output I11864;
wire I8830,I9179,I8827,I8854,I11830,I11847,I11395,I11624,I8862,I9258,I8848,I11378,I9066,I11813,I9227,I11310,I11327,I8851;
nand I_0(I8830,I8913,I9227);
DFFARX1 I_1(I1470,I8862,,,I9179,);
DFFARX1 I_2(I9258,I1470,I8862,,,I8827,);
nor I_3(I8854,I9179);
not I_4(I11830,I11813);
nand I_5(I11847,I11830,I11395);
nand I_6(I11395,I11378,I8851);
nand I_7(I11624,I11327,I8827);
not I_8(I8862,I1477);
or I_9(I9258,I9179,I9148);
nor I_10(I8848,I9083);
nor I_11(I11378,I11327,I8848);
DFFARX1 I_12(I1470,I8862,,,I9066,);
DFFARX1 I_13(I8854,I1470,I11310,,,I11813,);
nor I_14(I9227,I9179);
not I_15(I11310,I1477);
not I_16(I11327,I8830);
or I_17(I8851,I9083,I9066);
and I_18(I11864,I11624,I11847);
endmodule


