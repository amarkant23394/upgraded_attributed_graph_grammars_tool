module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_7_r_4,n6_4,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_7_r_4,n6_4,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_7_r_4,n6_4,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_7_r_4,n6_4,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
nor I_43(N1371_0_r_4,n25_4,G78_5_r_9);
not I_44(N1508_0_r_4,n25_4);
nor I_45(N1507_6_r_4,n32_4,n33_4);
nor I_46(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_47(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_48(n_572_7_r_4,n_573_7_r_4);
nand I_49(n_573_7_r_4,n21_4,n22_4);
nor I_50(n_549_7_r_4,n24_4,G78_5_r_9);
nand I_51(n_569_7_r_4,n22_4,n23_4);
nor I_52(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_53(N6147_9_r_4,n28_4);
nor I_54(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_55(I_BUFF_1_9_r_4,n21_4);
nor I_56(n4_7_r_4,N6147_9_r_4,G78_5_r_9);
not I_57(n6_4,blif_reset_net_7_r_4);
nand I_58(n21_4,n39_4,n40_4);
or I_59(n22_4,n31_4,N1372_4_r_9);
not I_60(n23_4,G78_5_r_9);
nor I_61(n24_4,n25_4,n26_4);
nand I_62(n25_4,n_42_8_r_9,N6147_9_r_9);
nand I_63(n26_4,n21_4,n27_4);
nand I_64(n27_4,n36_4,n37_4);
nand I_65(n28_4,n38_4,N6147_2_r_9);
nand I_66(n29_4,N1508_0_r_4,n30_4);
nand I_67(n30_4,n34_4,n35_4);
nor I_68(n31_4,n_576_5_r_9,n_547_5_r_9);
not I_69(n32_4,n30_4);
nor I_70(n33_4,n21_4,n28_4);
nand I_71(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_72(n35_4,N1508_0_r_4,n27_4);
not I_73(n36_4,N6147_2_r_9);
nand I_74(n37_4,G199_8_r_9,N6134_9_r_9);
or I_75(n38_4,n_576_5_r_9,n_547_5_r_9);
nor I_76(n39_4,N1372_4_r_9,n_576_5_r_9);
or I_77(n40_4,n41_4,N1508_4_r_9);
nor I_78(n41_4,N1508_4_r_9,G78_5_r_9);
endmodule


