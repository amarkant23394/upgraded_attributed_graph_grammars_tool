module test_I4725(I2215,I2492,I2557,I1477,I1470,I4725);
input I2215,I2492,I2557,I1477,I1470;
output I4725;
wire I2181,I2232,I2574,I4708,I2164,I2345,I2393,I2263,I2158,I2146;
not I_0(I2181,I1477);
DFFARX1 I_1(I2215,I1470,I2181,,,I2232,);
or I_2(I2574,I2557,I2492);
nand I_3(I4708,I2146,I2164);
and I_4(I4725,I4708,I2158);
DFFARX1 I_5(I2574,I1470,I2181,,,I2164,);
DFFARX1 I_6(I1470,I2181,,,I2345,);
DFFARX1 I_7(I2345,I1470,I2181,,,I2393,);
DFFARX1 I_8(I2232,I1470,I2181,,,I2263,);
not I_9(I2158,I2263);
and I_10(I2146,I2232,I2393);
endmodule


