module test_I2103(I1750,I1477,I1295,I1603,I1470,I1207,I1455,I2103);
input I1750,I1477,I1295,I1603,I1470,I1207,I1455;
output I2103;
wire I1518,I1784,I2038,I2021,I1535,I1832,I1849,I1620,I1767;
not I_0(I1518,I1477);
nor I_1(I1784,I1767,I1620);
not I_2(I2038,I2021);
DFFARX1 I_3(I1295,I1470,I1518,,,I2021,);
or I_4(I2103,I2038,I1849);
not I_5(I1535,I1455);
nand I_6(I1832,I1535,I1207);
and I_7(I1849,I1832,I1784);
not I_8(I1620,I1603);
DFFARX1 I_9(I1750,I1470,I1518,,,I1767,);
endmodule


