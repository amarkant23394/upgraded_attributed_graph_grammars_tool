module test_final(IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_clk_net_3_r_10,blif_reset_net_3_r_10,n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10);
input IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_clk_net_3_r_10,blif_reset_net_3_r_10;
output n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10;
wire ACVQN2_0_r_8,n_266_and_0_0_r_8,ACVQN1_2_r_8,P6_2_r_8,n_429_or_0_3_r_8,G78_3_r_8,n_576_3_r_8,n_102_3_r_8,n_547_3_r_8,n_42_5_r_8,G199_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8,ACVQN1_0_l_8,N1_1_l_8,G199_1_l_8,G214_1_l_8,n3_1_l_8,n_42_5_l_8,N3_5_l_8,G199_5_l_8,n3_5_l_8,ACVQN1_0_r_8,P6_internal_2_r_8,n12_3_r_8,n_431_3_r_8,n11_3_r_8,n13_3_r_8,n14_3_r_8,n15_3_r_8,n16_3_r_8,N3_5_r_8,n3_5_r_8,n2_3_r_10,ACVQN2_0_l_10,n_266_and_0_0_l_10,ACVQN1_0_l_10,n4_4_l_10,G42_4_l_10,n_87_4_l_10,n_572_4_l_10,n_573_4_l_10,n_549_4_l_10,n7_4_l_10,n_569_4_l_10,n_452_4_l_10,n12_3_r_10,n_431_3_r_10,n11_3_r_10,n13_3_r_10,n14_3_r_10,n15_3_r_10,n16_3_r_10,n4_4_r_10,n_87_4_r_10,n7_4_r_10;
DFFARX1 I_0(n_266_and_0_0_l_8,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_r_8,);
and I_1(n_266_and_0_0_r_8,G199_5_l_8,ACVQN1_0_r_8);
DFFARX1 I_2(G199_5_l_8,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_2_r_8,);
not I_3(P6_2_r_8,P6_internal_2_r_8);
nand I_4(n_429_or_0_3_r_8,G199_5_l_8,n12_3_r_8);
DFFARX1 I_5(n_431_3_r_8,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_8,);
nand I_6(n_576_3_r_8,n_42_5_l_8,n11_3_r_8);
not I_7(n_102_3_r_8,n_266_and_0_0_l_8);
nand I_8(n_547_3_r_8,ACVQN2_0_l_8,n13_3_r_8);
nor I_9(n_42_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8);
DFFARX1 I_10(N3_5_r_8,blif_clk_net_3_r_10,n2_3_r_10,G199_5_r_8,);
DFFARX1 I_11(IN_1_0_l_8,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_8,);
and I_12(n_266_and_0_0_l_8,IN_4_0_l_8,ACVQN1_0_l_8);
DFFARX1 I_13(IN_2_0_l_8,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_8,);
and I_14(N1_1_l_8,IN_6_1_l_8,n3_1_l_8);
DFFARX1 I_15(N1_1_l_8,blif_clk_net_3_r_10,n2_3_r_10,G199_1_l_8,);
DFFARX1 I_16(IN_3_1_l_8,blif_clk_net_3_r_10,n2_3_r_10,G214_1_l_8,);
nand I_17(n3_1_l_8,IN_1_1_l_8,IN_2_1_l_8);
nor I_18(n_42_5_l_8,IN_1_5_l_8,IN_3_5_l_8);
and I_19(N3_5_l_8,IN_6_5_l_8,n3_5_l_8);
DFFARX1 I_20(N3_5_l_8,blif_clk_net_3_r_10,n2_3_r_10,G199_5_l_8,);
nand I_21(n3_5_l_8,IN_2_5_l_8,IN_3_5_l_8);
DFFARX1 I_22(G214_1_l_8,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_r_8,);
DFFARX1 I_23(G214_1_l_8,blif_clk_net_3_r_10,n2_3_r_10,P6_internal_2_r_8,);
not I_24(n12_3_r_8,G199_1_l_8);
or I_25(n_431_3_r_8,n_42_5_l_8,n14_3_r_8);
nor I_26(n11_3_r_8,n_266_and_0_0_l_8,n12_3_r_8);
nor I_27(n13_3_r_8,n_266_and_0_0_l_8,G199_1_l_8);
and I_28(n14_3_r_8,ACVQN2_0_l_8,n15_3_r_8);
nor I_29(n15_3_r_8,G199_1_l_8,n16_3_r_8);
not I_30(n16_3_r_8,G199_5_l_8);
and I_31(N3_5_r_8,n_42_5_l_8,n3_5_r_8);
nand I_32(n3_5_r_8,ACVQN2_0_l_8,G214_1_l_8);
nand I_33(n_429_or_0_3_r_10,n_266_and_0_0_l_10,n12_3_r_10);
DFFARX1 I_34(n_431_3_r_10,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_10,);
nand I_35(n_576_3_r_10,ACVQN2_0_l_10,n11_3_r_10);
not I_36(n_102_3_r_10,G42_4_l_10);
nand I_37(n_547_3_r_10,n_569_4_l_10,n13_3_r_10);
DFFARX1 I_38(n4_4_r_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_10,);
nor I_39(n_572_4_r_10,ACVQN2_0_l_10,n_573_4_l_10);
or I_40(n_573_4_r_10,n_569_4_l_10,n_452_4_l_10);
nor I_41(n_549_4_r_10,n_572_4_l_10,n7_4_r_10);
or I_42(n_569_4_r_10,n_572_4_l_10,n_569_4_l_10);
nor I_43(n_452_4_r_10,n_266_and_0_0_l_10,n_452_4_l_10);
not I_44(n2_3_r_10,blif_reset_net_3_r_10);
DFFARX1 I_45(G78_3_r_8,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_10,);
and I_46(n_266_and_0_0_l_10,ACVQN1_0_l_10,P6_2_r_8);
DFFARX1 I_47(n_102_3_r_8,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_10,);
nor I_48(n4_4_l_10,ACVQN1_2_r_8,n_42_5_r_8);
DFFARX1 I_49(n4_4_l_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_l_10,);
not I_50(n_87_4_l_10,n_429_or_0_3_r_8);
nor I_51(n_572_4_l_10,n_429_or_0_3_r_8,n_547_3_r_8);
or I_52(n_573_4_l_10,ACVQN2_0_r_8,G199_5_r_8);
nor I_53(n_549_4_l_10,n7_4_l_10,n_266_and_0_0_r_8);
and I_54(n7_4_l_10,n_87_4_l_10,n_576_3_r_8);
or I_55(n_569_4_l_10,n_266_and_0_0_r_8,G199_5_r_8);
nor I_56(n_452_4_l_10,ACVQN2_0_r_8,ACVQN1_2_r_8);
not I_57(n12_3_r_10,n_549_4_l_10);
or I_58(n_431_3_r_10,n_572_4_l_10,n14_3_r_10);
nor I_59(n11_3_r_10,G42_4_l_10,n12_3_r_10);
nor I_60(n13_3_r_10,G42_4_l_10,n_549_4_l_10);
and I_61(n14_3_r_10,ACVQN2_0_l_10,n15_3_r_10);
nor I_62(n15_3_r_10,n_573_4_l_10,n16_3_r_10);
not I_63(n16_3_r_10,n_266_and_0_0_l_10);
nor I_64(n4_4_r_10,n_266_and_0_0_l_10,G42_4_l_10);
not I_65(n_87_4_r_10,ACVQN2_0_l_10);
and I_66(n7_4_r_10,n_452_4_l_10,n_87_4_r_10);
endmodule


