module test_I13248(I1477,I1470,I11460,I11864,I13248);
input I1477,I1470,I11460,I11864;
output I13248;
wire I13214,I11672,I13231,I11290,I11720,I13197,I11813,I11830,I11275,I11302,I11310;
nand I_0(I13214,I11275,I11302);
DFFARX1 I_1(I1470,I11310,,,I11672,);
and I_2(I13231,I13214,I11290);
nand I_3(I11290,I11830,I11720);
nor I_4(I11720,I11672,I11460);
not I_5(I13197,I1477);
DFFARX1 I_6(I1470,I11310,,,I11813,);
not I_7(I11830,I11813);
DFFARX1 I_8(I11672,I1470,I11310,,,I11275,);
DFFARX1 I_9(I11864,I1470,I11310,,,I11302,);
DFFARX1 I_10(I13231,I1470,I13197,,,I13248,);
not I_11(I11310,I1477);
endmodule


