module test_I3348(I1294,I2569,I2702,I1301,I3348);
input I1294,I2569,I2702,I1301;
output I3348;
wire I3263,I3314,I2548,I2583,I3024,I3041,I3331,I2545,I3246,I2945;
not I_0(I3263,I2569);
nor I_1(I3314,I3263,I2548);
DFFARX1 I_2(I2945,I1294,I2583,,,I2548,);
not I_3(I2583,I1301);
nand I_4(I3024,I2945);
and I_5(I3041,I2702,I3024);
nand I_6(I3331,I3314,I2545);
DFFARX1 I_7(I3041,I1294,I2583,,,I2545,);
not I_8(I3246,I1301);
DFFARX1 I_9(I3331,I1294,I3246,,,I3348,);
DFFARX1 I_10(I1294,I2583,,,I2945,);
endmodule


