module test_I2167(I1231,I1477,I1470,I1239,I1271,I1287,I2167);
input I1231,I1477,I1470,I1239,I1271,I1287;
output I2167;
wire I2181,I2328,I2232,I2294,I2311,I2198,I2633,I2215;
nand I_0(I2167,I2633,I2328);
not I_1(I2181,I1477);
nor I_2(I2328,I2232,I2311);
DFFARX1 I_3(I2215,I1470,I2181,,,I2232,);
nor I_4(I2294,I1287,I1231);
not I_5(I2311,I2294);
nand I_6(I2198,I1231);
DFFARX1 I_7(I1239,I1470,I2181,,,I2633,);
and I_8(I2215,I2198,I1271);
endmodule


