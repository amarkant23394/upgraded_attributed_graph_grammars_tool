module test_I4051(I2721,I1477,I1470,I4051);
input I2721,I1477,I1470;
output I4051;
wire I2730,I4017,I4000,I3076,I4034,I2724,I3983;
not I_0(I2730,I3076);
and I_1(I4017,I4000,I2730);
nand I_2(I4000,I2721,I2724);
DFFARX1 I_3(I1470,,,I3076,);
DFFARX1 I_4(I4017,I1470,I3983,,,I4034,);
not I_5(I4051,I4034);
DFFARX1 I_6(I1470,,,I2724,);
not I_7(I3983,I1477);
endmodule


