module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2,n4_7_l_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_2,n32_2,n35_2);
nor I_1(N1508_0_r_2,n32_2,n55_2);
not I_2(N1372_1_r_2,n54_2);
nor I_3(N1508_1_r_2,n59_2,n54_2);
nor I_4(N6147_2_r_2,n42_2,n43_2);
nor I_5(N1507_6_r_2,n40_2,n53_2);
nor I_6(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_7(n4_7_r_2,blif_clk_net_8_r_6,n9_6,G42_7_r_2,);
nor I_8(n_572_7_r_2,n36_2,n37_2);
or I_9(n_573_7_r_2,n34_2,n35_2);
nor I_10(n_549_7_r_2,n40_2,n41_2);
nand I_11(n_569_7_r_2,n38_2,n39_2);
nor I_12(n_452_7_r_2,n59_2,n35_2);
nor I_13(n4_7_l_2,G18_7_l_2,IN_1_7_l_2);
DFFARX1 I_14(n4_7_l_2,blif_clk_net_8_r_6,n9_6,n59_2,);
not I_15(n33_2,n59_2);
and I_16(N3_8_l_2,IN_6_8_l_2,n49_2);
DFFARX1 I_17(N3_8_l_2,blif_clk_net_8_r_6,n9_6,n32_internal_2,);
not I_18(n32_2,n32_internal_2);
nor I_19(n4_7_r_2,n59_2,n36_2);
not I_20(n34_2,n39_2);
nor I_21(n35_2,IN_1_8_l_2,IN_3_8_l_2);
nor I_22(n36_2,G18_7_l_2,IN_5_7_l_2);
or I_23(n37_2,IN_9_7_l_2,IN_10_7_l_2);
not I_24(n38_2,n40_2);
nand I_25(n39_2,n45_2,n57_2);
nor I_26(n40_2,IN_3_1_l_2,n47_2);
nor I_27(n41_2,n32_2,n36_2);
not I_28(n42_2,n53_2);
nand I_29(n43_2,n44_2,n45_2);
nand I_30(n44_2,n38_2,n46_2);
not I_31(n45_2,IN_10_7_l_2);
nand I_32(n46_2,n47_2,n48_2);
nand I_33(n47_2,IN_1_1_l_2,IN_2_1_l_2);
or I_34(n48_2,G15_7_l_2,IN_7_7_l_2);
nand I_35(n49_2,IN_2_8_l_2,IN_3_8_l_2);
nand I_36(n50_2,n51_2,n52_2);
not I_37(n51_2,n47_2);
nand I_38(n52_2,n38_2,n53_2);
nor I_39(n53_2,IN_5_7_l_2,IN_9_7_l_2);
nand I_40(n54_2,n42_2,n56_2);
nor I_41(n55_2,n34_2,n56_2);
nor I_42(n56_2,G15_7_l_2,IN_7_7_l_2);
nand I_43(n57_2,IN_4_7_l_2,n58_2);
not I_44(n58_2,G15_7_l_2);
nor I_45(N1371_0_r_6,n30_6,n33_6);
nor I_46(N1508_0_r_6,n33_6,n44_6);
not I_47(N1372_1_r_6,n41_6);
nor I_48(N1508_1_r_6,n40_6,n41_6);
nor I_49(N1507_6_r_6,n39_6,n45_6);
nor I_50(N1508_6_r_6,n37_6,n38_6);
nor I_51(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_52(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_53(N6147_9_r_6,n32_6,n33_6);
nor I_54(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_55(I_BUFF_1_9_r_6,n37_6);
not I_56(N1372_10_r_6,n43_6);
nor I_57(N1508_10_r_6,n42_6,n43_6);
nor I_58(N3_8_r_6,n36_6,N1372_1_r_2);
not I_59(n9_6,blif_reset_net_8_r_6);
nor I_60(n30_6,n53_6,n_569_7_r_2);
not I_61(n31_6,n36_6);
nor I_62(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_63(n33_6,N1372_1_r_2);
not I_64(n34_6,n35_6);
nand I_65(n35_6,n49_6,n_572_7_r_2);
nand I_66(n36_6,n51_6,N1371_0_r_2);
nand I_67(n37_6,n54_6,n_452_7_r_2);
or I_68(n38_6,n35_6,n39_6);
nor I_69(n39_6,n40_6,n45_6);
and I_70(n40_6,n46_6,n47_6);
nand I_71(n41_6,n30_6,n31_6);
nor I_72(n42_6,n34_6,n40_6);
nand I_73(n43_6,n30_6,N1372_1_r_2);
nor I_74(n44_6,n31_6,n40_6);
nor I_75(n45_6,n35_6,n36_6);
nor I_76(n46_6,N1508_6_r_2,n_573_7_r_2);
or I_77(n47_6,n48_6,N6147_2_r_2);
nor I_78(n48_6,N1508_1_r_2,N1508_0_r_2);
and I_79(n49_6,n50_6,N1508_0_r_2);
nand I_80(n50_6,n51_6,n52_6);
nand I_81(n51_6,G42_7_r_2,N1371_0_r_2);
not I_82(n52_6,N1371_0_r_2);
nor I_83(n53_6,N1507_6_r_2,n_549_7_r_2);
or I_84(n54_6,N1507_6_r_2,n_549_7_r_2);
endmodule


