module test_I10366(I8107,I1477,I7547,I7669,I6321,I7714,I1470,I10366);
input I8107,I1477,I7547,I7669,I6321,I7714,I1470;
output I10366;
wire I10185,I10202,I10219,I7731,I10052,I7977,I10349,I7541,I10332,I7550,I7562,I7570,I7532;
nand I_0(I10185,I7547,I7562);
and I_1(I10202,I10185,I7541);
DFFARX1 I_2(I10202,I1470,I10052,,,I10219,);
not I_3(I7731,I7714);
not I_4(I10052,I1477);
DFFARX1 I_5(I6321,I1470,I7570,,,I7977,);
nand I_6(I10366,I10349,I10219);
and I_7(I10349,I10332,I7550);
DFFARX1 I_8(I7669,I1470,I7570,,,I7541,);
DFFARX1 I_9(I7532,I1470,I10052,,,I10332,);
nand I_10(I7550,I7977,I7731);
nand I_11(I7562,I8107);
not I_12(I7570,I1477);
DFFARX1 I_13(I8107,I1470,I7570,,,I7532,);
endmodule


