module test_I1699(I1207,I1699);
input I1207;
output I1699;
wire ;
not I_0(I1699,I1207);
endmodule


