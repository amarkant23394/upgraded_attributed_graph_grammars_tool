module test_I14948(I12602,I12605,I15064,I1477,I1470,I14948);
input I12602,I12605,I15064,I1477,I1470;
output I14948;
wire I15485,I15389,I15406,I15519,I14965,I15372,I15423,I15502;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
DFFARX1 I_1(I12605,I1470,I14965,,,I15485,);
not I_2(I15389,I15372);
nor I_3(I15406,I15064,I15389);
or I_4(I15519,I15502,I15423);
not I_5(I14965,I1477);
DFFARX1 I_6(I12602,I1470,I14965,,,I15372,);
and I_7(I15423,I15372,I15406);
not I_8(I15502,I15485);
endmodule


