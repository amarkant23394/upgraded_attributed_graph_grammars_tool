module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_12,n8_12,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_12,n8_12,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_12,n8_12,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_12,n8_12,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_12,n8_12,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_12,n8_12,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_33(n_572_1_r_12,n29_12,n30_12);
nand I_34(n_573_1_r_12,n26_12,n27_12);
nor I_35(n_549_1_r_12,n33_12,n34_12);
and I_36(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_37(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_38(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_39(P6_5_r_12,P6_5_r_internal_12);
or I_40(n_431_0_l_12,n36_12,n_569_1_r_16);
not I_41(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_42(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_43(G214_4_r_16,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_44(n22_12,ACVQN1_5_l_12);
DFFARX1 I_45(n_573_1_r_16,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_46(n4_1_r_12,n41_12,n31_12);
nor I_47(N3_2_r_12,n22_12,n40_12);
not I_48(n3_12,n39_12);
DFFARX1 I_49(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_50(n26_12,ACVQN1_5_r_16,P6_5_r_16);
nor I_51(n27_12,n28_12,n29_12);
not I_52(n28_12,n_452_1_r_16);
nand I_53(n29_12,n31_12,n32_12);
nand I_54(n30_12,n42_12,n_452_1_r_16);
not I_55(n31_12,G42_1_r_16);
not I_56(n32_12,n_549_1_r_16);
nand I_57(n33_12,n31_12,n35_12);
nand I_58(n34_12,ACVQN1_5_r_16,P6_5_r_16);
nand I_59(n35_12,n41_12,n42_12);
and I_60(n36_12,n37_12,G199_4_r_16);
nor I_61(n37_12,n38_12,G42_1_r_16);
not I_62(n38_12,n_572_1_r_16);
nor I_63(n39_12,n38_12,P6_5_r_16);
nor I_64(n40_12,n39_12,G42_1_r_16);
endmodule


