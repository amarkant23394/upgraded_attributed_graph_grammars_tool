module test_I1316(I1255,I1247,I1279,I1294,I1271,I1207,I1301,I1316);
input I1255,I1247,I1279,I1294,I1271,I1207,I1301;
output I1316;
wire I1622,I1342,I1475,I1509,I1492,I1687,I1639;
nand I_0(I1316,I1509,I1687);
DFFARX1 I_1(I1255,I1294,I1342,,,I1622,);
not I_2(I1342,I1301);
nand I_3(I1475,I1247,I1271);
DFFARX1 I_4(I1492,I1294,I1342,,,I1509,);
and I_5(I1492,I1475,I1279);
not I_6(I1687,I1639);
and I_7(I1639,I1622,I1207);
endmodule


