module test_I11232(I10879,I1477,I9737,I9771,I10732,I9576,I1470,I11232);
input I10879,I1477,I9737,I9771,I10732,I9576,I1470;
output I11232;
wire I10647,I10961,I10978,I10664,I9474,I9471,I9542,I11167,I9459,I10896,I10749,I11150,I10913;
not I_0(I10647,I1477);
nand I_1(I10961,I10664,I9459);
and I_2(I10978,I10961,I10913);
not I_3(I10664,I9471);
or I_4(I9474,I9576,I9542);
nor I_5(I9471,I9542);
DFFARX1 I_6(I1470,,,I9542,);
not I_7(I11167,I11150);
nand I_8(I9459,I9771,I9737);
DFFARX1 I_9(I10879,I1470,I10647,,,I10896,);
not I_10(I10749,I10732);
DFFARX1 I_11(I9474,I1470,I10647,,,I11150,);
nor I_12(I10913,I10896,I10749);
or I_13(I11232,I11167,I10978);
endmodule


