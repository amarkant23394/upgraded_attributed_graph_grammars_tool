module test_I13174(I1477,I11299,I13265,I1470,I11624,I13174);
input I1477,I11299,I13265,I1470,I11624;
output I13174;
wire I13697,I13680,I13601,I13197,I13426,I11302,I11278,I11310,I13296,I13443,I11864;
or I_0(I13697,I13296,I13680);
and I_1(I13680,I13601,I13443);
DFFARX1 I_2(I11299,I1470,I13197,,,I13601,);
not I_3(I13197,I1477);
DFFARX1 I_4(I1470,I13197,,,I13426,);
DFFARX1 I_5(I13697,I1470,I13197,,,I13174,);
DFFARX1 I_6(I11864,I1470,I11310,,,I11302,);
DFFARX1 I_7(I11624,I1470,I11310,,,I11278,);
not I_8(I11310,I1477);
nor I_9(I13296,I11278,I11302);
nor I_10(I13443,I13426,I13265);
and I_11(I11864,I11624);
endmodule


