module Benchmark_testing10000(I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I252,I260,I268,I276,I284,I292,I300,I308,I316,I324,I332,I340,I348,I356,I364,I372,I380,I388,I396,I404,I412,I420,I428,I436,I444,I452,I460,I468,I476,I484,I492,I500,I508,I516,I524,I532,I540,I548,I556,I564,I572,I580,I588,I596,I604,I612,I620,I628,I636,I644,I652,I660,I668,I676,I684,I691,I698,I23855,I24026,I24089,I24116,I24161,I24224,I24323,I24386,I24413,I47327,I47498,I47561,I47588,I47633,I47696,I47795,I47858,I47885,I71024,I71087,I71141,I71195,I71294,I71330,I71384,I71411,I71429,I94343,I94460,I94550,I94577,I94640,I94667,I94685,I94703,I94730,I117878,I117959,I117995,I118166,I118184,I118211,I118301,I118391,I118409,I141062,I141125,I141179,I141233,I141332,I141368,I141422,I141449,I141467,I164381,I164498,I164588,I164615,I164678,I164705,I164723,I164741,I164768);
input I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I252,I260,I268,I276,I284,I292,I300,I308,I316,I324,I332,I340,I348,I356,I364,I372,I380,I388,I396,I404,I412,I420,I428,I436,I444,I452,I460,I468,I476,I484,I492,I500,I508,I516,I524,I532,I540,I548,I556,I564,I572,I580,I588,I596,I604,I612,I620,I628,I636,I644,I652,I660,I668,I676,I684,I691,I698;
output I23855,I24026,I24089,I24116,I24161,I24224,I24323,I24386,I24413,I47327,I47498,I47561,I47588,I47633,I47696,I47795,I47858,I47885,I71024,I71087,I71141,I71195,I71294,I71330,I71384,I71411,I71429,I94343,I94460,I94550,I94577,I94640,I94667,I94685,I94703,I94730,I117878,I117959,I117995,I118166,I118184,I118211,I118301,I118391,I118409,I141062,I141125,I141179,I141233,I141332,I141368,I141422,I141449,I141467,I164381,I164498,I164588,I164615,I164678,I164705,I164723,I164741,I164768;
wire I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I252,I260,I268,I276,I284,I292,I300,I308,I316,I324,I332,I340,I348,I356,I364,I372,I380,I388,I396,I404,I412,I420,I428,I436,I444,I452,I460,I468,I476,I484,I492,I500,I508,I516,I524,I532,I540,I548,I556,I564,I572,I580,I588,I596,I604,I612,I620,I628,I636,I644,I652,I660,I668,I676,I684,I691,I698,I707,I734,I752,I761,I779,I806,I815,I833,I851,I869,I887,I905,I923,I941,I968,I977,I995,I1013,I1031,I1049,I1067,I1085,I1112,I1130,I1139,I1157,I1175,I1193,I1220,I1229,I1247,I1265,I1292,I1301,I1319,I1337,I1364,I1373,I1391,I1409,I1436,I1454,I1463,I1481,I1508,I1517,I1535,I1553,I1580,I1598,I1607,I1625,I1652,I1670,I1679,I1697,I1715,I1733,I1751,I1769,I1787,I1814,I1823,I1841,I1859,I1877,I1895,I1922,I1940,I1949,I1967,I1994,I2003,I2021,I2039,I2057,I2075,I2093,I2111,I2138,I2147,I2165,I2183,I2210,I2219,I2237,I2255,I2282,I2291,I2318,I2327,I2345,I2363,I2381,I2399,I2426,I2435,I2453,I2471,I2489,I2507,I2525,I2552,I2561,I2588,I2606,I2615,I2633,I2651,I2669,I2696,I2705,I2723,I2741,I2768,I2777,I2795,I2813,I2831,I2849,I2876,I2894,I2903,I2921,I2939,I2957,I2984,I2993,I3011,I3029,I3047,I3065,I3083,I3101,I3119,I3137,I3164,I3173,I3191,I3218,I3227,I3245,I3272,I3281,I3299,I3326,I3335,I3353,I3371,I3398,I3416,I3425,I3443,I3461,I3479,I3497,I3524,I3533,I3560,I3578,I3587,I3605,I3623,I3641,I3659,I3686,I3695,I3722,I3740,I3749,I3767,I3794,I3803,I3821,I3839,I3857,I3875,I3893,I3911,I3929,I3947,I3965,I3983,I4001,I4019,I4037,I4064,I4073,I4100,I4109,I4127,I4145,I4163,I4190,I4199,I4226,I4235,I4253,I4271,I4289,I4316,I4325,I4343,I4361,I4388,I4406,I4424,I4433,I4451,I4478,I4487,I4505,I4532,I4541,I4559,I4577,I4595,I4622,I4631,I4649,I4667,I4685,I4703,I4721,I4748,I4757,I4784,I4793,I4811,I4829,I4847,I4874,I4883,I4901,I4919,I4946,I4955,I4982,I4991,I5009,I5027,I5045,I5063,I5090,I5099,I5117,I5135,I5153,I5180,I5189,I5207,I5234,I5243,I5270,I5279,I5297,I5315,I5333,I5360,I5369,I5387,I5405,I5423,I5450,I5459,I5486,I5495,I5522,I5531,I5549,I5567,I5585,I5603,I5630,I5639,I5657,I5675,I5693,I5711,I5729,I5747,I5765,I5783,I5801,I5819,I5837,I5855,I5873,I5891,I5909,I5936,I5945,I5972,I5990,I5999,I6017,I6035,I6062,I6071,I6098,I6116,I6125,I6143,I6161,I6179,I6206,I6215,I6242,I6251,I6269,I6287,I6314,I6323,I6350,I6359,I6377,I6395,I6422,I6431,I6449,I6467,I6485,I6512,I6521,I6539,I6557,I6575,I6593,I6620,I6638,I6647,I6674,I6683,I6701,I6719,I6746,I6755,I6782,I6791,I6809,I6827,I6845,I6863,I6890,I6899,I6917,I6935,I6953,I6980,I6989,I7007,I7034,I7043,I7070,I7079,I7097,I7115,I7133,I7160,I7169,I7187,I7205,I7223,I7250,I7259,I7286,I7304,I7313,I7331,I7349,I7376,I7394,I7412,I7430,I7439,I7457,I7475,I7502,I7511,I7529,I7547,I7565,I7583,I7610,I7619,I7646,I7655,I7673,I7691,I7709,I7727,I7754,I7763,I7781,I7799,I7817,I7844,I7853,I7871,I7889,I7916,I7925,I7952,I7961,I7979,I7997,I8015,I8033,I8060,I8069,I8087,I8105,I8123,I8150,I8159,I8177,I8204,I8213,I8240,I8249,I8267,I8285,I8303,I8330,I8339,I8357,I8375,I8393,I8420,I8429,I8456,I8474,I8483,I8501,I8519,I8537,I8555,I8573,I8600,I8609,I8627,I8654,I8663,I8681,I8699,I8726,I8735,I8753,I8780,I8789,I8807,I8825,I8843,I8861,I8879,I8897,I8915,I8942,I8951,I8969,I8987,I9005,I9023,I9041,I9059,I9077,I9095,I9113,I9140,I9158,I9167,I9185,I9203,I9230,I9248,I9266,I9284,I9293,I9311,I9329,I9356,I9365,I9383,I9401,I9419,I9437,I9464,I9473,I9500,I9509,I9527,I9545,I9563,I9581,I9608,I9617,I9635,I9653,I9671,I9698,I9707,I9734,I9743,I9761,I9779,I9797,I9815,I9842,I9851,I9869,I9887,I9905,I9923,I9941,I9959,I9977,I9995,I10013,I10031,I10049,I10067,I10085,I10103,I10121,I10148,I10157,I10184,I10202,I10211,I10229,I10247,I10274,I10283,I10310,I10328,I10337,I10355,I10382,I10391,I10409,I10427,I10445,I10463,I10481,I10499,I10517,I10544,I10553,I10571,I10589,I10607,I10625,I10643,I10661,I10688,I10706,I10715,I10733,I10751,I10769,I10796,I10805,I10823,I10841,I10868,I10877,I10895,I10913,I10940,I10949,I10976,I10994,I11003,I11021,I11039,I11057,I11084,I11093,I11111,I11129,I11156,I11165,I11183,I11201,I11219,I11237,I11264,I11282,I11291,I11309,I11327,I11345,I11372,I11381,I11399,I11417,I11435,I11453,I11471,I11489,I11507,I11525,I11552,I11561,I11588,I11597,I11615,I11633,I11651,I11669,I11696,I11705,I11723,I11741,I11759,I11777,I11795,I11813,I11831,I11849,I11867,I11885,I11903,I11921,I11939,I11957,I11975,I12002,I12011,I12038,I12056,I12065,I12083,I12101,I12128,I12137,I12164,I12182,I12191,I12209,I12236,I12245,I12263,I12281,I12299,I12317,I12335,I12353,I12371,I12398,I12407,I12425,I12443,I12461,I12479,I12497,I12515,I12542,I12560,I12569,I12587,I12605,I12623,I12650,I12659,I12677,I12695,I12722,I12731,I12749,I12767,I12794,I12812,I12821,I12839,I12857,I12875,I12893,I12911,I12938,I12947,I12965,I12992,I13001,I13019,I13037,I13064,I13073,I13091,I13118,I13127,I13145,I13163,I13181,I13199,I13217,I13235,I13253,I13280,I13289,I13307,I13325,I13343,I13361,I13379,I13397,I13415,I13433,I13451,I13478,I13496,I13505,I13523,I13541,I13568,I13586,I13604,I13622,I13631,I13649,I13667,I13694,I13703,I13721,I13739,I13757,I13775,I13802,I13811,I13838,I13847,I13865,I13883,I13901,I13919,I13946,I13955,I13973,I13991,I14009,I14036,I14054,I14063,I14081,I14108,I14117,I14135,I14153,I14171,I14189,I14207,I14225,I14252,I14261,I14279,I14297,I14324,I14333,I14351,I14369,I14396,I14405,I14432,I14441,I14459,I14477,I14495,I14513,I14540,I14549,I14567,I14585,I14603,I14621,I14639,I14666,I14684,I14693,I14711,I14729,I14747,I14774,I14783,I14810,I14819,I14837,I14855,I14882,I14891,I14918,I14927,I14945,I14963,I14990,I14999,I15017,I15035,I15053,I15080,I15089,I15107,I15125,I15143,I15161,I15188,I15206,I15215,I15242,I15251,I15269,I15287,I15314,I15332,I15341,I15359,I15386,I15395,I15413,I15431,I15458,I15476,I15485,I15503,I15530,I15548,I15557,I15575,I15593,I15611,I15629,I15647,I15665,I15692,I15701,I15719,I15737,I15755,I15773,I15800,I15818,I15827,I15845,I15872,I15881,I15899,I15917,I15935,I15953,I15971,I15989,I16016,I16025,I16043,I16061,I16088,I16097,I16115,I16133,I16160,I16169,I16196,I16205,I16223,I16241,I16259,I16277,I16304,I16313,I16331,I16349,I16367,I16385,I16403,I16430,I16439,I16457,I16475,I16502,I16511,I16538,I16547,I16565,I16583,I16601,I16619,I16646,I16655,I16673,I16691,I16709,I16736,I16745,I16763,I16790,I16799,I16826,I16835,I16853,I16871,I16889,I16916,I16925,I16943,I16961,I16979,I17006,I17015,I17042,I17051,I17078,I17096,I17105,I17123,I17141,I17159,I17186,I17195,I17213,I17231,I17258,I17267,I17285,I17303,I17321,I17339,I17366,I17384,I17393,I17411,I17429,I17447,I17474,I17483,I17501,I17519,I17537,I17555,I17573,I17591,I17609,I17627,I17654,I17663,I17690,I17699,I17717,I17735,I17753,I17771,I17798,I17807,I17825,I17843,I17861,I17879,I17897,I17915,I17933,I17951,I17969,I17987,I18005,I18023,I18041,I18059,I18077,I18104,I18113,I18140,I18158,I18167,I18185,I18203,I18230,I18239,I18266,I18284,I18293,I18320,I18329,I18347,I18365,I18383,I18401,I18419,I18437,I18464,I18473,I18491,I18509,I18527,I18554,I18563,I18581,I18599,I18617,I18635,I18662,I18671,I18689,I18707,I18734,I18743,I18761,I18779,I18797,I18824,I18833,I18851,I18869,I18896,I18905,I18923,I18941,I18968,I18977,I19004,I19013,I19031,I19049,I19067,I19085,I19112,I19121,I19139,I19157,I19175,I19202,I19211,I19229,I19256,I19265,I19292,I19301,I19319,I19337,I19355,I19382,I19391,I19409,I19427,I19445,I19472,I19481,I19508,I19517,I19544,I19562,I19571,I19589,I19607,I19625,I19643,I19661,I19679,I19697,I19715,I19733,I19751,I19769,I19796,I19805,I19823,I19841,I19868,I19877,I19895,I19913,I19940,I19949,I19967,I19985,I20012,I20021,I20039,I20057,I20084,I20093,I20120,I20138,I20147,I20165,I20183,I20201,I20228,I20237,I20255,I20273,I20300,I20309,I20327,I20345,I20363,I20381,I20408,I20426,I20435,I20453,I20471,I20489,I20516,I20525,I20543,I20561,I20579,I20597,I20615,I20633,I20651,I20669,I20696,I20705,I20723,I20741,I20768,I20777,I20804,I20813,I20831,I20849,I20867,I20885,I20912,I20921,I20939,I20957,I20975,I21002,I21011,I21029,I21056,I21065,I21092,I21101,I21119,I21137,I21155,I21182,I21191,I21209,I21227,I21245,I21272,I21281,I21308,I21326,I21335,I21353,I21380,I21389,I21407,I21425,I21443,I21461,I21479,I21497,I21515,I21533,I21551,I21569,I21587,I21605,I21623,I21650,I21659,I21686,I21695,I21713,I21731,I21749,I21776,I21785,I21812,I21821,I21839,I21857,I21875,I21902,I21911,I21929,I21947,I21974,I21983,I22010,I22019,I22037,I22055,I22073,I22091,I22118,I22127,I22145,I22163,I22181,I22208,I22217,I22235,I22262,I22271,I22298,I22307,I22325,I22343,I22361,I22388,I22397,I22415,I22433,I22451,I22478,I22487,I22514,I22532,I22541,I22568,I22577,I22595,I22613,I22631,I22649,I22667,I22685,I22712,I22721,I22739,I22757,I22775,I22802,I22811,I22829,I22847,I22865,I22883,I22910,I22919,I22937,I22955,I22982,I22991,I23009,I23027,I23045,I23072,I23081,I23099,I23117,I23144,I23162,I23171,I23189,I23207,I23225,I23243,I23261,I23288,I23297,I23315,I23342,I23351,I23369,I23387,I23414,I23423,I23441,I23468,I23477,I23495,I23513,I23531,I23549,I23567,I23585,I23603,I23630,I23639,I23657,I23675,I23693,I23711,I23729,I23747,I23765,I23783,I23801,I23828,I23846,I23882,I23891,I23909,I23927,I23945,I23963,I23981,I23999,I24035,I24053,I24071,I24125,I24143,I24179,I24197,I24233,I24251,I24269,I24296,I24305,I24341,I24359,I24395,I24431,I24458,I24476,I24485,I24503,I24530,I24539,I24557,I24575,I24593,I24611,I24629,I24647,I24665,I24683,I24701,I24719,I24737,I24755,I24773,I24800,I24809,I24836,I24845,I24863,I24881,I24899,I24926,I24935,I24962,I24971,I24989,I25007,I25025,I25052,I25061,I25079,I25106,I25115,I25133,I25151,I25169,I25187,I25214,I25223,I25241,I25259,I25277,I25295,I25313,I25331,I25358,I25367,I25385,I25403,I25421,I25439,I25457,I25484,I25493,I25520,I25529,I25556,I25574,I25583,I25601,I25619,I25637,I25664,I25673,I25691,I25709,I25736,I25754,I25772,I25781,I25799,I25826,I25835,I25853,I25880,I25889,I25907,I25925,I25943,I25970,I25979,I25997,I26015,I26033,I26051,I26069,I26096,I26105,I26132,I26141,I26159,I26177,I26195,I26222,I26240,I26249,I26267,I26294,I26303,I26321,I26339,I26357,I26375,I26393,I26411,I26438,I26447,I26465,I26483,I26510,I26519,I26537,I26555,I26582,I26591,I26618,I26627,I26645,I26663,I26681,I26699,I26726,I26735,I26753,I26771,I26789,I26807,I26825,I26852,I26870,I26879,I26897,I26924,I26933,I26951,I26969,I26987,I27005,I27023,I27041,I27059,I27086,I27095,I27113,I27131,I27149,I27167,I27185,I27203,I27230,I27248,I27257,I27275,I27293,I27311,I27338,I27347,I27365,I27383,I27410,I27419,I27437,I27455,I27482,I27491,I27509,I27527,I27554,I27563,I27590,I27599,I27617,I27635,I27653,I27671,I27698,I27707,I27725,I27743,I27761,I27788,I27797,I27815,I27842,I27851,I27878,I27887,I27905,I27923,I27941,I27968,I27977,I27995,I28013,I28031,I28058,I28067,I28094,I28112,I28121,I28139,I28157,I28184,I28202,I28220,I28238,I28247,I28265,I28283,I28310,I28319,I28337,I28355,I28373,I28391,I28418,I28427,I28454,I28463,I28481,I28499,I28517,I28535,I28562,I28571,I28589,I28607,I28625,I28652,I28670,I28679,I28706,I28715,I28733,I28751,I28769,I28787,I28805,I28823,I28850,I28859,I28877,I28895,I28913,I28940,I28949,I28967,I28985,I29003,I29021,I29048,I29057,I29075,I29093,I29120,I29129,I29147,I29165,I29183,I29210,I29219,I29237,I29255,I29282,I29291,I29318,I29327,I29345,I29363,I29381,I29399,I29426,I29435,I29453,I29471,I29489,I29507,I29525,I29543,I29561,I29579,I29597,I29615,I29633,I29651,I29669,I29687,I29705,I29732,I29741,I29768,I29786,I29795,I29813,I29831,I29858,I29867,I29894,I29912,I29921,I29939,I29966,I29975,I29993,I30011,I30029,I30047,I30065,I30083,I30110,I30119,I30137,I30155,I30182,I30191,I30209,I30227,I30254,I30263,I30290,I30299,I30317,I30335,I30353,I30371,I30398,I30407,I30425,I30443,I30461,I30479,I30497,I30524,I30533,I30551,I30569,I30596,I30605,I30632,I30641,I30659,I30677,I30695,I30713,I30740,I30749,I30767,I30785,I30803,I30830,I30839,I30857,I30884,I30893,I30920,I30929,I30947,I30965,I30983,I31010,I31019,I31037,I31055,I31073,I31100,I31109,I31136,I31154,I31163,I31181,I31208,I31217,I31235,I31253,I31271,I31289,I31307,I31325,I31352,I31361,I31379,I31397,I31424,I31433,I31451,I31469,I31496,I31505,I31532,I31541,I31559,I31577,I31595,I31613,I31640,I31649,I31667,I31685,I31703,I31721,I31739,I31766,I31775,I31793,I31811,I31838,I31856,I31874,I31883,I31901,I31928,I31937,I31955,I31982,I31991,I32009,I32027,I32045,I32072,I32081,I32099,I32117,I32135,I32153,I32171,I32198,I32207,I32234,I32243,I32261,I32279,I32297,I32324,I32342,I32351,I32369,I32396,I32405,I32423,I32441,I32459,I32477,I32495,I32513,I32531,I32558,I32567,I32585,I32603,I32621,I32639,I32657,I32675,I32702,I32720,I32729,I32747,I32765,I32783,I32810,I32819,I32837,I32855,I32882,I32891,I32909,I32927,I32954,I32963,I32981,I32999,I33026,I33044,I33053,I33071,I33098,I33107,I33125,I33143,I33170,I33188,I33197,I33215,I33242,I33260,I33269,I33287,I33305,I33323,I33341,I33359,I33377,I33404,I33413,I33431,I33449,I33467,I33485,I33512,I33521,I33539,I33566,I33575,I33593,I33620,I33629,I33647,I33674,I33683,I33701,I33719,I33746,I33764,I33773,I33791,I33809,I33827,I33845,I33872,I33881,I33908,I33926,I33935,I33953,I33971,I33989,I34007,I34034,I34043,I34070,I34079,I34097,I34124,I34133,I34151,I34169,I34187,I34205,I34232,I34241,I34259,I34277,I34295,I34313,I34331,I34349,I34376,I34385,I34403,I34421,I34439,I34457,I34475,I34502,I34511,I34538,I34547,I34574,I34592,I34601,I34619,I34637,I34655,I34682,I34691,I34709,I34727,I34754,I34772,I34781,I34799,I34826,I34835,I34853,I34871,I34898,I34916,I34925,I34943,I34970,I34988,I34997,I35015,I35033,I35051,I35069,I35087,I35105,I35132,I35141,I35159,I35177,I35195,I35213,I35240,I35258,I35267,I35285,I35303,I35321,I35339,I35357,I35384,I35393,I35411,I35438,I35447,I35465,I35483,I35510,I35519,I35537,I35564,I35573,I35591,I35609,I35627,I35645,I35663,I35681,I35699,I35726,I35735,I35753,I35771,I35789,I35807,I35825,I35843,I35861,I35879,I35897,I35924,I35933,I35951,I35969,I35996,I36005,I36032,I36041,I36059,I36077,I36095,I36113,I36140,I36149,I36167,I36185,I36203,I36230,I36239,I36257,I36284,I36293,I36320,I36329,I36347,I36365,I36383,I36410,I36419,I36437,I36455,I36473,I36500,I36509,I36536,I36545,I36572,I36581,I36599,I36617,I36635,I36653,I36680,I36689,I36707,I36725,I36743,I36761,I36779,I36797,I36815,I36833,I36851,I36869,I36887,I36905,I36923,I36941,I36959,I36986,I36995,I37022,I37040,I37049,I37067,I37085,I37112,I37121,I37148,I37166,I37175,I37193,I37220,I37229,I37247,I37265,I37283,I37301,I37319,I37337,I37355,I37382,I37391,I37409,I37427,I37445,I37463,I37481,I37499,I37526,I37544,I37553,I37571,I37589,I37607,I37634,I37643,I37661,I37679,I37706,I37715,I37733,I37751,I37778,I37787,I37805,I37823,I37850,I37868,I37886,I37895,I37913,I37940,I37949,I37967,I37994,I38003,I38021,I38039,I38057,I38084,I38093,I38111,I38129,I38147,I38165,I38183,I38210,I38219,I38246,I38255,I38273,I38291,I38309,I38336,I38354,I38363,I38381,I38408,I38417,I38435,I38453,I38471,I38489,I38507,I38525,I38552,I38561,I38579,I38597,I38624,I38633,I38651,I38669,I38696,I38705,I38732,I38741,I38759,I38777,I38795,I38813,I38840,I38849,I38867,I38885,I38903,I38921,I38939,I38966,I38975,I38993,I39011,I39038,I39056,I39074,I39083,I39101,I39128,I39137,I39155,I39182,I39191,I39209,I39227,I39245,I39272,I39281,I39299,I39317,I39335,I39353,I39371,I39398,I39407,I39434,I39443,I39461,I39479,I39497,I39524,I39542,I39551,I39569,I39587,I39605,I39632,I39641,I39668,I39677,I39695,I39713,I39740,I39749,I39776,I39785,I39803,I39821,I39848,I39857,I39875,I39893,I39911,I39938,I39947,I39965,I39983,I40001,I40019,I40046,I40064,I40073,I40100,I40118,I40127,I40145,I40172,I40181,I40199,I40217,I40235,I40253,I40271,I40289,I40307,I40334,I40343,I40361,I40379,I40397,I40415,I40433,I40451,I40478,I40496,I40505,I40523,I40541,I40559,I40586,I40595,I40613,I40631,I40658,I40667,I40685,I40703,I40730,I40739,I40757,I40775,I40802,I40820,I40829,I40847,I40874,I40883,I40901,I40919,I40946,I40964,I40973,I40991,I41018,I41036,I41045,I41063,I41081,I41099,I41117,I41135,I41153,I41180,I41189,I41207,I41225,I41243,I41261,I41288,I41297,I41324,I41342,I41351,I41369,I41387,I41405,I41432,I41441,I41459,I41477,I41504,I41513,I41531,I41549,I41567,I41585,I41612,I41630,I41639,I41657,I41675,I41693,I41720,I41729,I41747,I41765,I41783,I41801,I41819,I41837,I41855,I41873,I41900,I41918,I41927,I41945,I41963,I41990,I42008,I42026,I42044,I42053,I42071,I42089,I42116,I42125,I42143,I42161,I42179,I42197,I42224,I42233,I42260,I42269,I42287,I42305,I42323,I42341,I42368,I42377,I42395,I42413,I42431,I42458,I42476,I42485,I42503,I42521,I42539,I42557,I42575,I42602,I42611,I42629,I42656,I42665,I42683,I42701,I42728,I42737,I42755,I42782,I42791,I42809,I42827,I42845,I42863,I42881,I42899,I42917,I42944,I42953,I42971,I42989,I43007,I43025,I43043,I43061,I43079,I43097,I43115,I43142,I43160,I43169,I43187,I43214,I43223,I43241,I43259,I43277,I43295,I43313,I43331,I43358,I43367,I43385,I43403,I43430,I43439,I43457,I43475,I43502,I43511,I43538,I43547,I43565,I43583,I43601,I43619,I43646,I43655,I43673,I43691,I43709,I43727,I43745,I43772,I43781,I43808,I43826,I43835,I43853,I43871,I43889,I43916,I43925,I43943,I43961,I43988,I43997,I44015,I44033,I44051,I44069,I44096,I44114,I44123,I44141,I44159,I44177,I44204,I44213,I44231,I44249,I44267,I44285,I44303,I44321,I44339,I44357,I44384,I44393,I44411,I44429,I44456,I44474,I44483,I44501,I44528,I44537,I44555,I44573,I44600,I44618,I44627,I44645,I44672,I44690,I44699,I44717,I44735,I44753,I44771,I44789,I44807,I44834,I44843,I44861,I44879,I44897,I44915,I44942,I44951,I44969,I44987,I45014,I45023,I45050,I45059,I45077,I45095,I45113,I45131,I45158,I45167,I45185,I45203,I45221,I45248,I45257,I45275,I45302,I45311,I45338,I45347,I45365,I45383,I45401,I45428,I45437,I45455,I45473,I45491,I45518,I45527,I45554,I45572,I45581,I45599,I45626,I45635,I45653,I45671,I45689,I45707,I45725,I45743,I45770,I45779,I45797,I45815,I45842,I45851,I45869,I45887,I45914,I45923,I45950,I45959,I45977,I45995,I46013,I46031,I46058,I46067,I46085,I46103,I46121,I46139,I46157,I46184,I46202,I46211,I46229,I46247,I46274,I46292,I46310,I46328,I46337,I46355,I46373,I46400,I46409,I46427,I46445,I46463,I46481,I46508,I46517,I46544,I46553,I46571,I46589,I46607,I46625,I46652,I46661,I46679,I46697,I46715,I46742,I46751,I46769,I46796,I46805,I46823,I46850,I46859,I46877,I46904,I46913,I46931,I46949,I46976,I46994,I47003,I47021,I47039,I47057,I47075,I47102,I47111,I47138,I47156,I47165,I47183,I47201,I47219,I47237,I47264,I47273,I47300,I47318,I47354,I47363,I47381,I47399,I47417,I47435,I47453,I47471,I47507,I47525,I47543,I47597,I47615,I47651,I47669,I47705,I47723,I47741,I47768,I47777,I47813,I47831,I47867,I47903,I47930,I47939,I47957,I47984,I47993,I48011,I48029,I48047,I48065,I48092,I48101,I48119,I48137,I48155,I48173,I48191,I48209,I48236,I48245,I48263,I48281,I48299,I48317,I48335,I48362,I48371,I48398,I48407,I48434,I48452,I48461,I48479,I48497,I48515,I48542,I48551,I48569,I48587,I48614,I48623,I48650,I48659,I48677,I48695,I48713,I48731,I48758,I48767,I48785,I48803,I48821,I48848,I48857,I48875,I48902,I48911,I48938,I48947,I48965,I48983,I49001,I49028,I49037,I49055,I49073,I49091,I49118,I49127,I49154,I49163,I49190,I49208,I49217,I49235,I49253,I49271,I49298,I49307,I49325,I49343,I49370,I49379,I49397,I49415,I49433,I49451,I49478,I49496,I49505,I49523,I49541,I49559,I49586,I49595,I49613,I49631,I49649,I49667,I49685,I49703,I49721,I49739,I49766,I49784,I49793,I49811,I49829,I49856,I49874,I49892,I49910,I49919,I49937,I49955,I49982,I49991,I50009,I50027,I50045,I50063,I50090,I50099,I50126,I50135,I50153,I50171,I50189,I50207,I50234,I50243,I50261,I50279,I50297,I50324,I50333,I50360,I50378,I50387,I50405,I50423,I50441,I50468,I50477,I50495,I50513,I50540,I50549,I50567,I50585,I50603,I50621,I50648,I50666,I50675,I50693,I50711,I50729,I50756,I50765,I50783,I50801,I50819,I50837,I50855,I50873,I50891,I50909,I50936,I50954,I50963,I50981,I51008,I51017,I51035,I51053,I51071,I51089,I51107,I51125,I51143,I51170,I51179,I51197,I51215,I51233,I51251,I51269,I51287,I51314,I51332,I51341,I51359,I51377,I51395,I51422,I51431,I51449,I51467,I51494,I51503,I51521,I51539,I51566,I51575,I51602,I51620,I51629,I51647,I51665,I51683,I51710,I51719,I51737,I51755,I51782,I51791,I51809,I51827,I51845,I51863,I51890,I51908,I51917,I51935,I51953,I51971,I51998,I52007,I52025,I52043,I52061,I52079,I52097,I52115,I52133,I52151,I52178,I52196,I52205,I52223,I52250,I52259,I52277,I52295,I52313,I52331,I52349,I52367,I52385,I52412,I52421,I52439,I52457,I52475,I52493,I52511,I52529,I52556,I52574,I52583,I52601,I52619,I52637,I52664,I52673,I52691,I52709,I52736,I52745,I52763,I52781,I52808,I52817,I52844,I52853,I52871,I52889,I52907,I52925,I52952,I52961,I52979,I52997,I53015,I53033,I53051,I53069,I53087,I53105,I53123,I53141,I53159,I53177,I53195,I53213,I53231,I53258,I53267,I53294,I53312,I53321,I53339,I53357,I53384,I53393,I53420,I53429,I53456,I53474,I53483,I53501,I53519,I53537,I53564,I53573,I53591,I53609,I53636,I53645,I53663,I53681,I53699,I53717,I53744,I53762,I53771,I53789,I53807,I53825,I53852,I53861,I53879,I53897,I53915,I53933,I53951,I53969,I53987,I54005,I54032,I54050,I54059,I54077,I54104,I54113,I54131,I54149,I54167,I54185,I54203,I54221,I54239,I54257,I54275,I54293,I54311,I54329,I54347,I54374,I54383,I54410,I54419,I54437,I54455,I54473,I54500,I54509,I54536,I54545,I54563,I54581,I54599,I54626,I54635,I54653,I54680,I54689,I54707,I54734,I54743,I54761,I54788,I54797,I54815,I54833,I54860,I54878,I54887,I54905,I54923,I54941,I54959,I54986,I54995,I55022,I55040,I55049,I55067,I55085,I55103,I55121,I55148,I55157,I55184,I55193,I55220,I55238,I55247,I55265,I55283,I55301,I55328,I55337,I55355,I55373,I55400,I55409,I55427,I55445,I55463,I55481,I55508,I55526,I55535,I55553,I55571,I55589,I55616,I55625,I55643,I55661,I55679,I55697,I55715,I55733,I55751,I55769,I55796,I55814,I55823,I55841,I55868,I55877,I55895,I55913,I55931,I55949,I55967,I55985,I56012,I56021,I56039,I56057,I56084,I56093,I56111,I56129,I56156,I56165,I56192,I56201,I56219,I56237,I56255,I56273,I56300,I56309,I56327,I56345,I56363,I56381,I56399,I56426,I56435,I56453,I56471,I56498,I56507,I56534,I56543,I56561,I56579,I56597,I56615,I56642,I56651,I56669,I56687,I56705,I56732,I56741,I56759,I56786,I56795,I56822,I56831,I56849,I56867,I56885,I56912,I56921,I56939,I56957,I56975,I57002,I57011,I57038,I57056,I57065,I57083,I57101,I57119,I57146,I57155,I57182,I57191,I57209,I57227,I57254,I57263,I57290,I57299,I57317,I57335,I57362,I57371,I57389,I57407,I57425,I57452,I57461,I57479,I57497,I57515,I57533,I57560,I57578,I57587,I57614,I57623,I57641,I57659,I57686,I57704,I57713,I57731,I57758,I57767,I57785,I57803,I57830,I57848,I57857,I57875,I57902,I57920,I57929,I57947,I57965,I57983,I58001,I58019,I58037,I58064,I58073,I58091,I58109,I58127,I58145,I58172,I58181,I58199,I58226,I58235,I58253,I58280,I58289,I58307,I58334,I58343,I58361,I58379,I58406,I58424,I58433,I58451,I58469,I58487,I58505,I58532,I58541,I58568,I58586,I58595,I58613,I58631,I58649,I58667,I58694,I58703,I58730,I58748,I58757,I58775,I58793,I58820,I58838,I58856,I58874,I58883,I58901,I58919,I58946,I58955,I58973,I58991,I59009,I59027,I59054,I59063,I59090,I59099,I59117,I59135,I59153,I59171,I59198,I59207,I59225,I59243,I59261,I59288,I59306,I59315,I59333,I59360,I59369,I59387,I59405,I59423,I59441,I59459,I59477,I59495,I59522,I59531,I59549,I59567,I59585,I59603,I59621,I59639,I59666,I59684,I59693,I59711,I59729,I59747,I59774,I59783,I59801,I59819,I59846,I59855,I59873,I59891,I59918,I59927,I59954,I59972,I59981,I59999,I60017,I60035,I60062,I60071,I60089,I60107,I60134,I60143,I60161,I60179,I60197,I60215,I60242,I60260,I60269,I60287,I60305,I60323,I60350,I60359,I60377,I60395,I60413,I60431,I60449,I60467,I60485,I60503,I60530,I60548,I60557,I60584,I60593,I60611,I60629,I60647,I60665,I60683,I60701,I60728,I60737,I60755,I60773,I60791,I60818,I60827,I60845,I60863,I60881,I60899,I60926,I60935,I60953,I60971,I60998,I61007,I61025,I61043,I61061,I61088,I61097,I61115,I61133,I61160,I61178,I61187,I61205,I61223,I61241,I61259,I61277,I61304,I61313,I61331,I61358,I61367,I61385,I61403,I61430,I61439,I61457,I61484,I61493,I61511,I61529,I61547,I61565,I61583,I61601,I61619,I61646,I61655,I61673,I61691,I61709,I61727,I61745,I61763,I61781,I61799,I61817,I61844,I61853,I61880,I61889,I61907,I61925,I61943,I61961,I61988,I61997,I62015,I62033,I62051,I62069,I62087,I62105,I62123,I62141,I62159,I62177,I62195,I62213,I62231,I62249,I62267,I62294,I62303,I62330,I62348,I62357,I62375,I62393,I62420,I62429,I62456,I62465,I62492,I62510,I62519,I62537,I62555,I62573,I62600,I62609,I62627,I62645,I62672,I62681,I62699,I62717,I62735,I62753,I62780,I62798,I62807,I62825,I62843,I62861,I62888,I62897,I62915,I62933,I62951,I62969,I62987,I63005,I63023,I63041,I63068,I63077,I63095,I63113,I63140,I63158,I63176,I63185,I63203,I63230,I63239,I63257,I63284,I63293,I63311,I63329,I63347,I63374,I63383,I63401,I63419,I63437,I63455,I63473,I63500,I63509,I63536,I63545,I63563,I63581,I63599,I63626,I63635,I63662,I63680,I63689,I63707,I63725,I63743,I63770,I63779,I63797,I63815,I63842,I63851,I63869,I63887,I63905,I63923,I63950,I63968,I63977,I63995,I64013,I64031,I64058,I64067,I64085,I64103,I64121,I64139,I64157,I64175,I64193,I64211,I64238,I64247,I64265,I64283,I64310,I64328,I64337,I64355,I64382,I64391,I64409,I64427,I64454,I64472,I64481,I64499,I64526,I64544,I64553,I64571,I64589,I64607,I64625,I64643,I64661,I64688,I64697,I64715,I64733,I64751,I64769,I64796,I64805,I64823,I64841,I64868,I64877,I64904,I64913,I64931,I64949,I64967,I64985,I65012,I65021,I65039,I65057,I65075,I65102,I65111,I65129,I65156,I65165,I65192,I65201,I65219,I65237,I65255,I65282,I65291,I65309,I65327,I65345,I65372,I65381,I65408,I65426,I65435,I65453,I65471,I65489,I65507,I65525,I65552,I65561,I65579,I65606,I65615,I65633,I65651,I65678,I65687,I65705,I65732,I65741,I65759,I65777,I65795,I65813,I65831,I65849,I65867,I65894,I65903,I65921,I65939,I65957,I65975,I65993,I66011,I66029,I66047,I66065,I66092,I66101,I66119,I66137,I66164,I66182,I66191,I66209,I66236,I66245,I66263,I66281,I66308,I66326,I66335,I66353,I66380,I66398,I66407,I66425,I66443,I66461,I66479,I66497,I66515,I66542,I66551,I66569,I66587,I66605,I66623,I66650,I66668,I66677,I66695,I66722,I66731,I66749,I66767,I66785,I66803,I66821,I66839,I66857,I66875,I66893,I66911,I66929,I66947,I66965,I66992,I67001,I67028,I67037,I67055,I67073,I67091,I67118,I67127,I67154,I67163,I67181,I67199,I67217,I67244,I67262,I67271,I67289,I67316,I67325,I67343,I67361,I67379,I67397,I67415,I67433,I67451,I67478,I67487,I67505,I67523,I67541,I67559,I67577,I67595,I67622,I67640,I67649,I67667,I67685,I67703,I67730,I67739,I67757,I67775,I67802,I67811,I67829,I67847,I67874,I67883,I67910,I67919,I67937,I67955,I67973,I67991,I68018,I68027,I68045,I68063,I68081,I68099,I68117,I68135,I68153,I68171,I68189,I68207,I68225,I68243,I68261,I68279,I68297,I68324,I68333,I68360,I68378,I68387,I68405,I68423,I68450,I68459,I68486,I68504,I68513,I68531,I68558,I68567,I68585,I68603,I68621,I68639,I68657,I68675,I68693,I68720,I68729,I68747,I68765,I68783,I68801,I68819,I68837,I68864,I68882,I68891,I68909,I68927,I68945,I68972,I68981,I68999,I69017,I69044,I69053,I69071,I69089,I69116,I69125,I69143,I69170,I69179,I69197,I69224,I69233,I69251,I69278,I69287,I69305,I69323,I69350,I69368,I69377,I69395,I69413,I69431,I69449,I69476,I69485,I69512,I69530,I69539,I69557,I69575,I69593,I69611,I69638,I69647,I69674,I69683,I69710,I69728,I69737,I69755,I69773,I69791,I69818,I69827,I69845,I69863,I69890,I69899,I69917,I69935,I69953,I69971,I69998,I70016,I70025,I70043,I70061,I70079,I70106,I70115,I70133,I70151,I70169,I70187,I70205,I70223,I70241,I70259,I70286,I70304,I70313,I70331,I70349,I70367,I70394,I70403,I70430,I70439,I70457,I70475,I70502,I70511,I70538,I70547,I70565,I70583,I70610,I70619,I70637,I70655,I70673,I70700,I70709,I70727,I70745,I70763,I70781,I70808,I70826,I70835,I70862,I70871,I70889,I70916,I70925,I70943,I70961,I70979,I70997,I71033,I71051,I71069,I71105,I71123,I71168,I71177,I71213,I71231,I71249,I71267,I71303,I71339,I71366,I71393,I71447,I71474,I71492,I71501,I71519,I71546,I71555,I71573,I71591,I71609,I71627,I71645,I71663,I71681,I71708,I71717,I71735,I71753,I71771,I71789,I71807,I71825,I71852,I71870,I71879,I71897,I71915,I71933,I71960,I71969,I71987,I72005,I72032,I72041,I72059,I72077,I72104,I72113,I72140,I72158,I72167,I72185,I72203,I72221,I72248,I72257,I72275,I72293,I72320,I72329,I72347,I72365,I72383,I72401,I72428,I72446,I72455,I72473,I72491,I72509,I72536,I72545,I72563,I72581,I72599,I72617,I72635,I72653,I72671,I72689,I72716,I72725,I72743,I72761,I72788,I72806,I72815,I72833,I72860,I72869,I72887,I72905,I72932,I72950,I72959,I72977,I73004,I73022,I73031,I73049,I73067,I73085,I73103,I73121,I73139,I73166,I73175,I73193,I73211,I73229,I73247,I73274,I73292,I73301,I73319,I73346,I73355,I73373,I73391,I73409,I73427,I73445,I73463,I73481,I73508,I73517,I73535,I73553,I73571,I73589,I73607,I73625,I73652,I73670,I73679,I73697,I73715,I73733,I73760,I73769,I73787,I73805,I73832,I73841,I73859,I73877,I73904,I73913,I73931,I73949,I73976,I73994,I74012,I74021,I74039,I74066,I74075,I74093,I74120,I74129,I74147,I74165,I74183,I74210,I74219,I74237,I74255,I74273,I74291,I74309,I74336,I74345,I74372,I74381,I74399,I74417,I74435,I74462,I74471,I74498,I74516,I74525,I74543,I74561,I74579,I74606,I74615,I74633,I74651,I74678,I74687,I74705,I74723,I74741,I74759,I74786,I74804,I74813,I74831,I74849,I74867,I74894,I74903,I74921,I74939,I74957,I74975,I74993,I75011,I75029,I75047,I75074,I75083,I75101,I75128,I75137,I75155,I75182,I75191,I75209,I75236,I75245,I75263,I75281,I75308,I75326,I75335,I75353,I75371,I75389,I75407,I75434,I75443,I75470,I75488,I75497,I75515,I75533,I75551,I75569,I75596,I75605,I75632,I75641,I75659,I75686,I75695,I75713,I75731,I75749,I75767,I75794,I75803,I75821,I75839,I75857,I75875,I75893,I75911,I75938,I75947,I75965,I75983,I76001,I76019,I76037,I76064,I76073,I76100,I76109,I76136,I76154,I76163,I76181,I76199,I76217,I76244,I76253,I76271,I76298,I76307,I76325,I76352,I76361,I76379,I76406,I76415,I76433,I76451,I76478,I76496,I76505,I76523,I76541,I76559,I76577,I76604,I76613,I76640,I76658,I76667,I76685,I76703,I76721,I76739,I76766,I76775,I76802,I76811,I76829,I76847,I76874,I76892,I76910,I76919,I76937,I76964,I76973,I76991,I77018,I77027,I77045,I77063,I77081,I77108,I77117,I77135,I77153,I77171,I77189,I77207,I77234,I77243,I77270,I77279,I77297,I77315,I77333,I77360,I77378,I77387,I77405,I77432,I77441,I77459,I77477,I77495,I77513,I77531,I77549,I77567,I77594,I77603,I77621,I77639,I77657,I77675,I77693,I77711,I77738,I77756,I77765,I77783,I77801,I77819,I77846,I77855,I77873,I77891,I77918,I77927,I77945,I77963,I77990,I78008,I78017,I78044,I78053,I78071,I78089,I78107,I78125,I78143,I78161,I78188,I78197,I78215,I78233,I78251,I78278,I78287,I78305,I78323,I78341,I78359,I78386,I78395,I78413,I78431,I78458,I78467,I78485,I78503,I78521,I78548,I78557,I78575,I78593,I78620,I78638,I78647,I78665,I78692,I78701,I78719,I78737,I78755,I78773,I78791,I78809,I78827,I78854,I78863,I78881,I78899,I78917,I78935,I78953,I78971,I78998,I79016,I79025,I79043,I79061,I79079,I79106,I79115,I79133,I79151,I79178,I79187,I79205,I79223,I79250,I79259,I79286,I79295,I79313,I79331,I79349,I79367,I79394,I79403,I79421,I79439,I79457,I79475,I79493,I79511,I79529,I79547,I79565,I79583,I79601,I79619,I79637,I79655,I79673,I79700,I79709,I79736,I79754,I79763,I79781,I79799,I79826,I79835,I79862,I79871,I79889,I79907,I79934,I79943,I79970,I79979,I79997,I80015,I80033,I80051,I80078,I80087,I80105,I80123,I80141,I80168,I80177,I80195,I80222,I80231,I80258,I80267,I80285,I80303,I80321,I80348,I80357,I80375,I80393,I80411,I80438,I80447,I80474,I80483,I80501,I80528,I80537,I80555,I80582,I80591,I80609,I80636,I80645,I80663,I80681,I80708,I80726,I80735,I80753,I80771,I80789,I80807,I80834,I80843,I80870,I80888,I80897,I80915,I80933,I80951,I80969,I80996,I81005,I81032,I81041,I81059,I81077,I81104,I81122,I81131,I81149,I81176,I81185,I81203,I81221,I81248,I81266,I81275,I81293,I81320,I81338,I81347,I81365,I81383,I81401,I81419,I81437,I81455,I81482,I81491,I81509,I81527,I81545,I81563,I81590,I81608,I81617,I81635,I81653,I81671,I81698,I81707,I81734,I81743,I81761,I81779,I81806,I81815,I81842,I81851,I81869,I81887,I81914,I81923,I81941,I81959,I81977,I82004,I82013,I82031,I82049,I82067,I82085,I82112,I82130,I82139,I82166,I82175,I82193,I82211,I82238,I82247,I82274,I82283,I82301,I82319,I82337,I82355,I82382,I82391,I82409,I82427,I82445,I82472,I82481,I82499,I82526,I82535,I82562,I82571,I82589,I82607,I82625,I82652,I82661,I82679,I82697,I82715,I82742,I82751,I82778,I82787,I82814,I82832,I82841,I82859,I82877,I82895,I82922,I82931,I82949,I82967,I82994,I83003,I83021,I83039,I83057,I83075,I83102,I83120,I83129,I83147,I83165,I83183,I83210,I83219,I83237,I83255,I83273,I83291,I83309,I83327,I83345,I83363,I83390,I83399,I83417,I83444,I83453,I83471,I83498,I83507,I83525,I83552,I83561,I83579,I83597,I83624,I83642,I83651,I83669,I83687,I83705,I83723,I83750,I83759,I83786,I83804,I83813,I83831,I83849,I83867,I83885,I83912,I83921,I83948,I83957,I83984,I84002,I84011,I84029,I84047,I84065,I84083,I84101,I84119,I84137,I84155,I84173,I84191,I84209,I84236,I84245,I84263,I84281,I84308,I84317,I84335,I84353,I84380,I84389,I84407,I84425,I84452,I84461,I84479,I84497,I84524,I84542,I84551,I84569,I84596,I84605,I84623,I84641,I84659,I84677,I84695,I84713,I84731,I84758,I84767,I84785,I84803,I84821,I84839,I84857,I84875,I84902,I84920,I84929,I84947,I84965,I84983,I85010,I85019,I85037,I85055,I85082,I85091,I85109,I85127,I85154,I85163,I85190,I85208,I85217,I85235,I85253,I85271,I85298,I85307,I85325,I85343,I85370,I85379,I85397,I85415,I85433,I85451,I85478,I85496,I85505,I85523,I85541,I85559,I85586,I85595,I85613,I85631,I85649,I85667,I85685,I85703,I85721,I85739,I85766,I85775,I85793,I85811,I85838,I85847,I85874,I85883,I85901,I85919,I85937,I85955,I85982,I85991,I86009,I86027,I86045,I86072,I86081,I86099,I86126,I86135,I86162,I86171,I86189,I86207,I86225,I86252,I86261,I86279,I86297,I86315,I86342,I86351,I86378,I86387,I86405,I86423,I86450,I86468,I86486,I86495,I86513,I86540,I86549,I86567,I86594,I86603,I86621,I86639,I86657,I86684,I86693,I86711,I86729,I86747,I86765,I86783,I86810,I86819,I86846,I86855,I86873,I86891,I86909,I86936,I86954,I86963,I86981,I87008,I87017,I87035,I87053,I87071,I87089,I87107,I87125,I87143,I87170,I87179,I87197,I87215,I87233,I87251,I87269,I87287,I87314,I87332,I87341,I87359,I87377,I87395,I87422,I87431,I87449,I87467,I87494,I87503,I87521,I87539,I87566,I87575,I87593,I87620,I87629,I87647,I87674,I87683,I87701,I87728,I87737,I87755,I87773,I87800,I87818,I87827,I87845,I87863,I87881,I87899,I87926,I87935,I87962,I87980,I87989,I88007,I88025,I88043,I88061,I88088,I88097,I88124,I88133,I88151,I88169,I88196,I88214,I88232,I88241,I88259,I88286,I88295,I88313,I88340,I88349,I88367,I88385,I88403,I88430,I88439,I88457,I88475,I88493,I88511,I88529,I88556,I88565,I88592,I88601,I88619,I88637,I88655,I88682,I88691,I88718,I88736,I88745,I88763,I88781,I88799,I88826,I88835,I88853,I88871,I88898,I88907,I88925,I88943,I88961,I88979,I89006,I89024,I89033,I89051,I89069,I89087,I89114,I89123,I89141,I89159,I89177,I89195,I89213,I89231,I89249,I89267,I89294,I89303,I89330,I89339,I89357,I89375,I89393,I89411,I89438,I89447,I89465,I89483,I89501,I89519,I89537,I89555,I89573,I89591,I89609,I89627,I89645,I89663,I89681,I89699,I89717,I89744,I89753,I89780,I89798,I89807,I89825,I89843,I89870,I89879,I89906,I89915,I89933,I89951,I89978,I89987,I90014,I90023,I90041,I90059,I90077,I90095,I90122,I90131,I90149,I90167,I90185,I90212,I90221,I90239,I90266,I90275,I90302,I90311,I90329,I90347,I90365,I90392,I90401,I90419,I90437,I90455,I90482,I90491,I90518,I90536,I90545,I90563,I90590,I90599,I90617,I90635,I90653,I90671,I90689,I90707,I90725,I90752,I90761,I90779,I90797,I90815,I90833,I90851,I90869,I90896,I90914,I90923,I90941,I90959,I90977,I91004,I91013,I91031,I91049,I91076,I91085,I91103,I91121,I91148,I91157,I91184,I91193,I91211,I91229,I91247,I91265,I91292,I91301,I91319,I91337,I91355,I91373,I91391,I91409,I91427,I91445,I91463,I91481,I91499,I91517,I91535,I91553,I91571,I91598,I91607,I91634,I91652,I91661,I91679,I91697,I91724,I91733,I91760,I91778,I91787,I91805,I91823,I91841,I91868,I91877,I91904,I91913,I91931,I91949,I91976,I91985,I92012,I92021,I92039,I92057,I92084,I92093,I92111,I92129,I92147,I92174,I92183,I92201,I92219,I92237,I92255,I92282,I92300,I92309,I92336,I92345,I92363,I92381,I92408,I92426,I92444,I92453,I92471,I92498,I92507,I92525,I92552,I92561,I92579,I92597,I92615,I92642,I92651,I92669,I92687,I92705,I92723,I92741,I92768,I92777,I92804,I92813,I92831,I92849,I92867,I92894,I92912,I92921,I92939,I92966,I92975,I92993,I93011,I93029,I93047,I93065,I93083,I93110,I93119,I93137,I93155,I93182,I93191,I93209,I93227,I93254,I93263,I93290,I93299,I93317,I93335,I93353,I93371,I93398,I93407,I93425,I93443,I93461,I93479,I93497,I93524,I93542,I93551,I93569,I93596,I93605,I93623,I93641,I93659,I93677,I93695,I93713,I93731,I93758,I93767,I93785,I93803,I93821,I93839,I93857,I93875,I93902,I93920,I93929,I93947,I93965,I93983,I94010,I94019,I94037,I94055,I94082,I94091,I94109,I94127,I94154,I94163,I94181,I94199,I94226,I94235,I94262,I94271,I94289,I94307,I94325,I94370,I94379,I94397,I94415,I94433,I94469,I94487,I94514,I94523,I94559,I94595,I94613,I94649,I94739,I94766,I94775,I94793,I94811,I94838,I94847,I94874,I94883,I94901,I94919,I94937,I94955,I94982,I94991,I95009,I95027,I95045,I95072,I95081,I95099,I95126,I95135,I95162,I95171,I95189,I95207,I95225,I95252,I95261,I95279,I95297,I95315,I95342,I95351,I95378,I95396,I95405,I95423,I95441,I95459,I95486,I95495,I95522,I95531,I95549,I95567,I95594,I95603,I95630,I95639,I95657,I95675,I95702,I95711,I95729,I95747,I95765,I95792,I95801,I95819,I95837,I95855,I95873,I95900,I95918,I95927,I95954,I95963,I95981,I95999,I96026,I96044,I96062,I96071,I96089,I96116,I96125,I96143,I96170,I96179,I96197,I96215,I96233,I96260,I96269,I96287,I96305,I96323,I96341,I96359,I96386,I96395,I96422,I96431,I96449,I96467,I96485,I96512,I96521,I96548,I96557,I96575,I96593,I96611,I96629,I96656,I96665,I96683,I96701,I96719,I96737,I96755,I96773,I96791,I96809,I96827,I96845,I96863,I96881,I96899,I96917,I96935,I96962,I96971,I96998,I97016,I97025,I97043,I97061,I97088,I97097,I97124,I97142,I97151,I97169,I97187,I97205,I97223,I97241,I97268,I97277,I97295,I97322,I97331,I97349,I97367,I97394,I97403,I97421,I97448,I97457,I97475,I97493,I97511,I97529,I97547,I97565,I97583,I97610,I97619,I97637,I97655,I97673,I97691,I97709,I97727,I97745,I97763,I97781,I97808,I97817,I97835,I97853,I97880,I97889,I97916,I97925,I97943,I97961,I97979,I97997,I98024,I98033,I98051,I98069,I98087,I98114,I98123,I98141,I98168,I98177,I98204,I98213,I98231,I98249,I98267,I98294,I98303,I98321,I98339,I98357,I98384,I98393,I98420,I98438,I98447,I98465,I98492,I98501,I98519,I98537,I98555,I98573,I98591,I98609,I98627,I98654,I98663,I98681,I98699,I98717,I98735,I98753,I98771,I98798,I98816,I98825,I98843,I98861,I98879,I98906,I98915,I98933,I98951,I98978,I98987,I99005,I99023,I99050,I99059,I99077,I99095,I99122,I99140,I99158,I99167,I99185,I99212,I99221,I99239,I99266,I99275,I99293,I99311,I99329,I99356,I99365,I99383,I99401,I99419,I99437,I99455,I99482,I99491,I99518,I99527,I99545,I99563,I99581,I99608,I99617,I99635,I99653,I99680,I99689,I99716,I99725,I99743,I99761,I99779,I99797,I99824,I99833,I99851,I99869,I99887,I99914,I99923,I99941,I99968,I99977,I100004,I100013,I100031,I100049,I100067,I100094,I100103,I100121,I100139,I100157,I100184,I100193,I100220,I100238,I100247,I100265,I100292,I100301,I100319,I100337,I100355,I100373,I100391,I100409,I100427,I100445,I100463,I100481,I100499,I100517,I100535,I100562,I100571,I100598,I100607,I100625,I100643,I100661,I100688,I100697,I100724,I100733,I100751,I100769,I100787,I100814,I100823,I100841,I100868,I100877,I100895,I100913,I100940,I100949,I100976,I100985,I101003,I101021,I101039,I101057,I101075,I101093,I101111,I101129,I101147,I101165,I101183,I101210,I101219,I101237,I101264,I101273,I101291,I101318,I101327,I101354,I101363,I101381,I101408,I101417,I101435,I101453,I101480,I101498,I101516,I101525,I101543,I101570,I101579,I101597,I101624,I101633,I101651,I101669,I101687,I101714,I101723,I101741,I101759,I101777,I101795,I101813,I101840,I101849,I101876,I101885,I101903,I101921,I101939,I101966,I101984,I101993,I102011,I102029,I102047,I102065,I102083,I102110,I102119,I102137,I102164,I102173,I102191,I102209,I102236,I102245,I102263,I102290,I102299,I102317,I102335,I102353,I102371,I102389,I102407,I102425,I102452,I102461,I102479,I102497,I102515,I102533,I102551,I102569,I102587,I102605,I102623,I102650,I102659,I102677,I102695,I102722,I102731,I102758,I102767,I102785,I102803,I102821,I102839,I102866,I102875,I102893,I102911,I102929,I102956,I102965,I102983,I103010,I103019,I103046,I103055,I103073,I103091,I103109,I103136,I103145,I103163,I103181,I103199,I103226,I103235,I103262,I103271,I103298,I103316,I103325,I103343,I103361,I103379,I103406,I103415,I103433,I103451,I103478,I103487,I103505,I103523,I103541,I103559,I103586,I103604,I103613,I103631,I103649,I103667,I103694,I103703,I103721,I103739,I103757,I103775,I103793,I103811,I103829,I103847,I103874,I103892,I103901,I103928,I103937,I103955,I103973,I103991,I104009,I104027,I104045,I104072,I104081,I104099,I104117,I104135,I104162,I104171,I104189,I104207,I104225,I104243,I104270,I104279,I104297,I104315,I104342,I104351,I104369,I104387,I104405,I104432,I104441,I104459,I104477,I104504,I104513,I104531,I104549,I104576,I104585,I104612,I104621,I104639,I104657,I104675,I104693,I104720,I104729,I104747,I104765,I104783,I104810,I104819,I104837,I104864,I104873,I104900,I104909,I104927,I104945,I104963,I104990,I104999,I105017,I105035,I105053,I105080,I105089,I105116,I105125,I105143,I105170,I105179,I105197,I105215,I105233,I105251,I105278,I105287,I105305,I105323,I105341,I105359,I105377,I105395,I105422,I105431,I105449,I105467,I105485,I105503,I105521,I105548,I105557,I105584,I105593,I105620,I105638,I105647,I105665,I105683,I105701,I105728,I105746,I105755,I105782,I105791,I105809,I105827,I105845,I105863,I105881,I105899,I105926,I105935,I105953,I105971,I105989,I106016,I106025,I106043,I106061,I106079,I106097,I106124,I106133,I106151,I106169,I106196,I106205,I106223,I106241,I106259,I106286,I106295,I106313,I106331,I106358,I106367,I106385,I106403,I106430,I106439,I106466,I106475,I106493,I106511,I106529,I106547,I106574,I106583,I106601,I106619,I106637,I106664,I106673,I106691,I106718,I106727,I106754,I106763,I106781,I106799,I106817,I106844,I106853,I106871,I106889,I106907,I106934,I106943,I106970,I106979,I107006,I107024,I107033,I107051,I107069,I107087,I107114,I107123,I107141,I107159,I107186,I107195,I107213,I107231,I107249,I107267,I107294,I107312,I107321,I107339,I107357,I107375,I107402,I107411,I107429,I107447,I107465,I107483,I107501,I107519,I107537,I107555,I107582,I107600,I107609,I107636,I107645,I107663,I107681,I107699,I107717,I107735,I107753,I107780,I107789,I107807,I107825,I107843,I107870,I107879,I107897,I107915,I107933,I107951,I107978,I107987,I108005,I108023,I108050,I108059,I108077,I108095,I108113,I108140,I108149,I108167,I108185,I108212,I108230,I108239,I108257,I108275,I108293,I108311,I108329,I108356,I108365,I108383,I108410,I108419,I108437,I108455,I108482,I108491,I108509,I108536,I108545,I108563,I108581,I108599,I108617,I108635,I108653,I108671,I108698,I108707,I108725,I108743,I108761,I108779,I108797,I108815,I108833,I108851,I108869,I108896,I108905,I108923,I108941,I108968,I108977,I109004,I109013,I109031,I109049,I109067,I109085,I109112,I109121,I109139,I109157,I109175,I109202,I109211,I109229,I109256,I109265,I109292,I109301,I109319,I109337,I109355,I109382,I109391,I109409,I109427,I109445,I109472,I109481,I109508,I109517,I109544,I109562,I109571,I109589,I109607,I109625,I109652,I109661,I109679,I109697,I109724,I109733,I109751,I109769,I109787,I109805,I109832,I109850,I109859,I109877,I109895,I109913,I109940,I109949,I109967,I109985,I110003,I110021,I110039,I110057,I110075,I110093,I110120,I110129,I110147,I110165,I110192,I110210,I110219,I110237,I110264,I110273,I110291,I110309,I110336,I110354,I110363,I110381,I110408,I110426,I110435,I110453,I110471,I110489,I110507,I110525,I110543,I110570,I110579,I110597,I110615,I110633,I110651,I110678,I110687,I110705,I110723,I110750,I110759,I110786,I110795,I110813,I110831,I110849,I110867,I110894,I110903,I110921,I110939,I110957,I110984,I110993,I111011,I111038,I111047,I111074,I111083,I111101,I111119,I111137,I111164,I111173,I111191,I111209,I111227,I111254,I111263,I111290,I111299,I111326,I111344,I111353,I111371,I111389,I111407,I111434,I111443,I111461,I111479,I111506,I111515,I111533,I111551,I111569,I111587,I111614,I111632,I111641,I111659,I111677,I111695,I111722,I111731,I111749,I111767,I111785,I111803,I111821,I111839,I111857,I111875,I111902,I111920,I111929,I111947,I111965,I111983,I112010,I112019,I112046,I112055,I112073,I112091,I112118,I112127,I112154,I112163,I112181,I112199,I112226,I112235,I112253,I112271,I112289,I112316,I112325,I112343,I112361,I112379,I112397,I112424,I112442,I112451,I112478,I112487,I112505,I112532,I112541,I112559,I112586,I112595,I112613,I112640,I112649,I112667,I112685,I112712,I112730,I112739,I112757,I112775,I112793,I112811,I112838,I112847,I112874,I112892,I112901,I112919,I112937,I112955,I112973,I113000,I113009,I113036,I113045,I113072,I113081,I113099,I113117,I113135,I113153,I113180,I113189,I113207,I113225,I113243,I113261,I113279,I113297,I113315,I113333,I113351,I113369,I113387,I113405,I113423,I113441,I113459,I113486,I113495,I113522,I113540,I113549,I113567,I113585,I113612,I113621,I113648,I113657,I113684,I113702,I113711,I113729,I113747,I113765,I113792,I113801,I113819,I113837,I113864,I113873,I113891,I113909,I113927,I113945,I113972,I113990,I113999,I114017,I114035,I114053,I114080,I114089,I114107,I114125,I114143,I114161,I114179,I114197,I114215,I114233,I114260,I114278,I114287,I114305,I114323,I114341,I114359,I114377,I114404,I114413,I114431,I114458,I114467,I114485,I114503,I114530,I114539,I114557,I114584,I114593,I114611,I114629,I114647,I114665,I114683,I114701,I114719,I114746,I114755,I114773,I114791,I114809,I114827,I114845,I114863,I114881,I114899,I114917,I114944,I114953,I114971,I114989,I115016,I115034,I115052,I115061,I115079,I115106,I115115,I115133,I115160,I115169,I115187,I115205,I115223,I115250,I115259,I115277,I115295,I115313,I115331,I115349,I115376,I115385,I115412,I115421,I115439,I115457,I115475,I115502,I115511,I115538,I115556,I115565,I115583,I115601,I115619,I115646,I115655,I115673,I115691,I115718,I115727,I115745,I115763,I115781,I115799,I115826,I115844,I115853,I115871,I115889,I115907,I115934,I115943,I115961,I115979,I115997,I116015,I116033,I116051,I116069,I116087,I116114,I116123,I116141,I116168,I116177,I116195,I116213,I116231,I116249,I116276,I116285,I116303,I116321,I116339,I116357,I116375,I116393,I116420,I116429,I116447,I116465,I116483,I116501,I116519,I116546,I116555,I116582,I116591,I116618,I116636,I116645,I116663,I116681,I116699,I116726,I116735,I116753,I116771,I116798,I116816,I116825,I116843,I116870,I116879,I116897,I116915,I116942,I116960,I116969,I116987,I117014,I117032,I117041,I117059,I117077,I117095,I117113,I117131,I117149,I117176,I117185,I117203,I117221,I117239,I117257,I117284,I117293,I117311,I117329,I117356,I117374,I117392,I117401,I117419,I117446,I117455,I117473,I117500,I117509,I117527,I117545,I117563,I117590,I117599,I117617,I117635,I117653,I117671,I117689,I117716,I117725,I117752,I117761,I117779,I117797,I117815,I117842,I117851,I117896,I117905,I117923,I117941,I117986,I118013,I118031,I118058,I118067,I118085,I118103,I118121,I118139,I118193,I118229,I118247,I118274,I118283,I118319,I118337,I118355,I118373,I118427,I118454,I118472,I118481,I118499,I118517,I118544,I118562,I118580,I118598,I118607,I118625,I118643,I118670,I118679,I118697,I118715,I118733,I118751,I118778,I118787,I118814,I118823,I118841,I118859,I118877,I118895,I118922,I118931,I118949,I118967,I118985,I119012,I119030,I119039,I119057,I119075,I119093,I119120,I119129,I119156,I119165,I119183,I119201,I119228,I119237,I119264,I119273,I119291,I119309,I119336,I119345,I119363,I119381,I119399,I119426,I119435,I119453,I119471,I119489,I119507,I119534,I119552,I119561,I119588,I119597,I119615,I119633,I119660,I119669,I119696,I119705,I119723,I119741,I119759,I119777,I119804,I119813,I119831,I119849,I119867,I119894,I119903,I119921,I119948,I119957,I119984,I119993,I120011,I120029,I120047,I120074,I120083,I120101,I120119,I120137,I120164,I120173,I120200,I120218,I120227,I120245,I120263,I120281,I120308,I120317,I120344,I120353,I120371,I120389,I120416,I120425,I120452,I120461,I120479,I120497,I120524,I120533,I120551,I120569,I120587,I120614,I120623,I120641,I120659,I120677,I120695,I120722,I120740,I120749,I120776,I120785,I120803,I120821,I120848,I120866,I120875,I120893,I120920,I120929,I120947,I120965,I120992,I121010,I121019,I121037,I121064,I121082,I121091,I121109,I121127,I121145,I121163,I121181,I121199,I121226,I121235,I121253,I121271,I121289,I121307,I121334,I121343,I121361,I121388,I121397,I121415,I121442,I121451,I121469,I121496,I121505,I121523,I121541,I121568,I121586,I121595,I121613,I121631,I121649,I121667,I121694,I121703,I121730,I121748,I121757,I121775,I121793,I121811,I121829,I121856,I121865,I121892,I121901,I121928,I121946,I121955,I121973,I121991,I122009,I122036,I122045,I122063,I122081,I122108,I122117,I122135,I122153,I122171,I122189,I122216,I122234,I122243,I122261,I122279,I122297,I122324,I122333,I122351,I122369,I122387,I122405,I122423,I122441,I122459,I122477,I122504,I122522,I122531,I122549,I122567,I122585,I122612,I122621,I122648,I122657,I122675,I122693,I122720,I122729,I122756,I122765,I122783,I122801,I122828,I122837,I122855,I122873,I122891,I122918,I122927,I122945,I122963,I122981,I122999,I123026,I123044,I123053,I123080,I123089,I123107,I123125,I123152,I123161,I123188,I123197,I123215,I123233,I123251,I123269,I123296,I123305,I123323,I123341,I123359,I123386,I123395,I123413,I123440,I123449,I123476,I123485,I123503,I123521,I123539,I123566,I123575,I123593,I123611,I123629,I123656,I123665,I123692,I123701,I123728,I123737,I123755,I123773,I123791,I123809,I123827,I123845,I123863,I123881,I123899,I123917,I123935,I123962,I123971,I123998,I124007,I124025,I124043,I124070,I124079,I124106,I124115,I124133,I124151,I124169,I124187,I124205,I124223,I124241,I124268,I124277,I124295,I124322,I124340,I124349,I124367,I124385,I124412,I124430,I124448,I124466,I124475,I124493,I124511,I124538,I124547,I124565,I124583,I124601,I124619,I124646,I124655,I124682,I124691,I124709,I124727,I124745,I124763,I124790,I124799,I124817,I124835,I124853,I124880,I124889,I124907,I124934,I124943,I124961,I124988,I124997,I125015,I125042,I125051,I125069,I125087,I125114,I125132,I125141,I125159,I125177,I125195,I125213,I125240,I125249,I125276,I125294,I125303,I125321,I125339,I125357,I125375,I125402,I125411,I125438,I125456,I125465,I125483,I125501,I125519,I125537,I125555,I125582,I125591,I125609,I125636,I125645,I125663,I125681,I125708,I125717,I125735,I125762,I125771,I125789,I125807,I125825,I125843,I125861,I125879,I125897,I125924,I125933,I125951,I125969,I125987,I126005,I126023,I126041,I126059,I126077,I126095,I126122,I126131,I126149,I126167,I126194,I126203,I126230,I126239,I126257,I126275,I126293,I126311,I126338,I126347,I126365,I126383,I126401,I126428,I126437,I126455,I126482,I126491,I126518,I126527,I126545,I126563,I126581,I126608,I126617,I126635,I126653,I126671,I126698,I126707,I126734,I126743,I126770,I126788,I126797,I126815,I126833,I126851,I126878,I126887,I126905,I126923,I126950,I126959,I126977,I126995,I127013,I127031,I127058,I127076,I127085,I127103,I127121,I127139,I127166,I127175,I127193,I127211,I127229,I127247,I127265,I127283,I127301,I127319,I127346,I127355,I127373,I127400,I127409,I127427,I127454,I127463,I127481,I127508,I127517,I127535,I127553,I127580,I127598,I127607,I127625,I127643,I127661,I127679,I127706,I127715,I127742,I127760,I127769,I127787,I127805,I127823,I127841,I127868,I127877,I127904,I127922,I127931,I127949,I127967,I127985,I128012,I128021,I128048,I128057,I128075,I128093,I128120,I128129,I128156,I128165,I128183,I128201,I128228,I128237,I128255,I128273,I128291,I128318,I128327,I128345,I128363,I128381,I128399,I128426,I128444,I128453,I128480,I128498,I128507,I128525,I128543,I128561,I128579,I128597,I128624,I128633,I128651,I128678,I128687,I128705,I128723,I128750,I128759,I128777,I128804,I128813,I128831,I128849,I128867,I128885,I128903,I128921,I128939,I128966,I128975,I128993,I129011,I129029,I129047,I129065,I129083,I129101,I129119,I129137,I129164,I129173,I129191,I129209,I129236,I129254,I129272,I129281,I129299,I129326,I129335,I129353,I129380,I129389,I129407,I129425,I129443,I129470,I129479,I129497,I129515,I129533,I129551,I129569,I129596,I129605,I129632,I129641,I129659,I129677,I129695,I129722,I129740,I129749,I129767,I129785,I129812,I129830,I129848,I129866,I129875,I129893,I129911,I129938,I129947,I129965,I129983,I130001,I130019,I130046,I130055,I130082,I130091,I130109,I130127,I130145,I130163,I130190,I130199,I130217,I130235,I130253,I130280,I130289,I130307,I130325,I130352,I130361,I130388,I130397,I130415,I130433,I130451,I130469,I130496,I130505,I130523,I130541,I130559,I130586,I130595,I130613,I130640,I130649,I130676,I130685,I130703,I130721,I130739,I130766,I130775,I130793,I130811,I130829,I130856,I130865,I130892,I130901,I130919,I130946,I130955,I130973,I130991,I131009,I131027,I131054,I131063,I131081,I131099,I131117,I131135,I131153,I131171,I131198,I131207,I131225,I131243,I131261,I131279,I131297,I131324,I131333,I131360,I131369,I131396,I131414,I131423,I131441,I131459,I131477,I131504,I131513,I131540,I131558,I131567,I131585,I131603,I131621,I131648,I131657,I131675,I131693,I131720,I131729,I131747,I131765,I131783,I131801,I131828,I131846,I131855,I131873,I131891,I131909,I131936,I131945,I131963,I131981,I131999,I132017,I132035,I132053,I132071,I132089,I132116,I132125,I132143,I132170,I132179,I132197,I132224,I132233,I132251,I132278,I132287,I132305,I132323,I132350,I132368,I132377,I132395,I132413,I132431,I132449,I132476,I132485,I132512,I132530,I132539,I132557,I132575,I132593,I132611,I132638,I132647,I132674,I132683,I132701,I132719,I132746,I132755,I132782,I132791,I132809,I132827,I132845,I132863,I132890,I132899,I132917,I132935,I132953,I132980,I132989,I133007,I133034,I133043,I133070,I133079,I133097,I133115,I133133,I133160,I133169,I133187,I133205,I133223,I133250,I133259,I133286,I133295,I133322,I133331,I133349,I133367,I133385,I133403,I133430,I133439,I133457,I133475,I133493,I133511,I133529,I133547,I133565,I133583,I133601,I133619,I133637,I133655,I133673,I133691,I133709,I133736,I133745,I133772,I133790,I133799,I133817,I133835,I133862,I133871,I133898,I133907,I133925,I133943,I133970,I133988,I133997,I134015,I134042,I134051,I134069,I134087,I134114,I134132,I134141,I134159,I134186,I134204,I134213,I134231,I134249,I134267,I134285,I134303,I134321,I134348,I134357,I134375,I134393,I134411,I134429,I134456,I134474,I134483,I134501,I134519,I134537,I134564,I134573,I134600,I134609,I134627,I134645,I134672,I134681,I134708,I134717,I134735,I134753,I134780,I134789,I134807,I134825,I134843,I134870,I134879,I134897,I134915,I134933,I134951,I134978,I134996,I135005,I135032,I135041,I135059,I135086,I135095,I135113,I135131,I135149,I135167,I135194,I135203,I135221,I135239,I135257,I135275,I135293,I135311,I135338,I135347,I135365,I135383,I135401,I135419,I135437,I135464,I135473,I135500,I135509,I135536,I135554,I135563,I135581,I135599,I135617,I135644,I135653,I135680,I135698,I135707,I135725,I135743,I135761,I135788,I135797,I135815,I135833,I135860,I135869,I135887,I135905,I135923,I135941,I135968,I135986,I135995,I136013,I136031,I136049,I136076,I136085,I136103,I136121,I136139,I136157,I136175,I136193,I136211,I136229,I136256,I136265,I136283,I136301,I136328,I136346,I136364,I136373,I136391,I136418,I136427,I136445,I136472,I136481,I136499,I136517,I136535,I136562,I136571,I136589,I136607,I136625,I136643,I136661,I136688,I136697,I136724,I136733,I136751,I136769,I136787,I136814,I136823,I136841,I136868,I136877,I136895,I136913,I136931,I136949,I136976,I136985,I137003,I137021,I137039,I137057,I137075,I137093,I137120,I137129,I137147,I137165,I137183,I137201,I137219,I137246,I137255,I137282,I137291,I137318,I137336,I137345,I137363,I137381,I137399,I137426,I137435,I137453,I137471,I137498,I137507,I137534,I137543,I137561,I137579,I137597,I137615,I137642,I137651,I137669,I137687,I137705,I137732,I137741,I137759,I137786,I137795,I137822,I137831,I137849,I137867,I137885,I137912,I137921,I137939,I137957,I137975,I138002,I138011,I138038,I138047,I138074,I138083,I138101,I138119,I138137,I138155,I138182,I138191,I138209,I138227,I138245,I138263,I138281,I138299,I138317,I138335,I138353,I138371,I138389,I138407,I138425,I138443,I138461,I138488,I138497,I138524,I138542,I138551,I138569,I138587,I138614,I138623,I138650,I138659,I138677,I138695,I138722,I138740,I138758,I138767,I138785,I138812,I138821,I138839,I138866,I138875,I138893,I138911,I138929,I138956,I138965,I138983,I139001,I139019,I139037,I139055,I139082,I139091,I139118,I139127,I139145,I139163,I139181,I139208,I139217,I139235,I139262,I139271,I139289,I139316,I139325,I139343,I139370,I139379,I139397,I139415,I139442,I139460,I139469,I139487,I139505,I139523,I139541,I139568,I139577,I139604,I139622,I139631,I139649,I139667,I139685,I139703,I139730,I139739,I139766,I139775,I139793,I139811,I139838,I139856,I139865,I139883,I139910,I139919,I139937,I139955,I139982,I140000,I140009,I140027,I140054,I140072,I140081,I140099,I140117,I140135,I140153,I140171,I140189,I140216,I140225,I140243,I140261,I140279,I140297,I140324,I140333,I140360,I140378,I140387,I140405,I140423,I140441,I140459,I140477,I140495,I140513,I140531,I140549,I140567,I140585,I140612,I140621,I140639,I140657,I140684,I140693,I140711,I140729,I140756,I140765,I140783,I140801,I140828,I140837,I140855,I140873,I140900,I140909,I140927,I140954,I140963,I140981,I140999,I141017,I141035,I141071,I141089,I141107,I141143,I141161,I141206,I141215,I141251,I141269,I141287,I141305,I141341,I141377,I141404,I141431,I141485,I141512,I141521,I141548,I141557,I141575,I141593,I141611,I141629,I141656,I141665,I141683,I141701,I141719,I141737,I141755,I141773,I141791,I141809,I141827,I141845,I141863,I141881,I141899,I141917,I141935,I141962,I141971,I141998,I142016,I142025,I142043,I142061,I142088,I142097,I142124,I142142,I142151,I142169,I142187,I142214,I142232,I142250,I142268,I142277,I142295,I142313,I142340,I142349,I142367,I142385,I142403,I142421,I142448,I142457,I142484,I142493,I142511,I142529,I142547,I142565,I142592,I142601,I142619,I142637,I142655,I142682,I142691,I142709,I142736,I142745,I142763,I142781,I142799,I142817,I142844,I142853,I142871,I142889,I142907,I142925,I142943,I142961,I142988,I142997,I143015,I143033,I143051,I143069,I143087,I143114,I143123,I143150,I143159,I143186,I143204,I143213,I143231,I143249,I143267,I143294,I143303,I143330,I143348,I143357,I143375,I143393,I143411,I143429,I143447,I143465,I143483,I143501,I143519,I143537,I143555,I143582,I143591,I143609,I143627,I143654,I143663,I143681,I143699,I143726,I143735,I143753,I143771,I143798,I143807,I143825,I143843,I143870,I143888,I143897,I143915,I143942,I143951,I143969,I143987,I144005,I144023,I144041,I144059,I144077,I144104,I144113,I144131,I144149,I144167,I144185,I144203,I144221,I144248,I144266,I144275,I144293,I144311,I144329,I144356,I144365,I144383,I144401,I144428,I144437,I144455,I144473,I144500,I144509,I144527,I144554,I144563,I144581,I144608,I144617,I144635,I144662,I144671,I144689,I144707,I144734,I144752,I144761,I144779,I144797,I144815,I144833,I144860,I144869,I144896,I144914,I144923,I144941,I144959,I144977,I144995,I145022,I145031,I145058,I145067,I145085,I145103,I145130,I145148,I145157,I145175,I145202,I145211,I145229,I145247,I145274,I145292,I145301,I145319,I145346,I145364,I145373,I145391,I145409,I145427,I145445,I145463,I145481,I145508,I145517,I145535,I145553,I145571,I145589,I145616,I145625,I145643,I145661,I145688,I145706,I145724,I145733,I145751,I145778,I145787,I145805,I145832,I145841,I145859,I145877,I145895,I145922,I145931,I145949,I145967,I145985,I146003,I146021,I146048,I146057,I146084,I146093,I146111,I146129,I146147,I146174,I146183,I146201,I146219,I146246,I146255,I146282,I146291,I146309,I146327,I146345,I146363,I146390,I146399,I146417,I146435,I146453,I146480,I146489,I146507,I146534,I146543,I146570,I146579,I146597,I146615,I146633,I146660,I146669,I146687,I146705,I146723,I146750,I146759,I146786,I146795,I146822,I146840,I146849,I146867,I146885,I146903,I146930,I146939,I146957,I146975,I147002,I147011,I147029,I147047,I147065,I147083,I147110,I147128,I147137,I147155,I147173,I147191,I147218,I147227,I147245,I147263,I147281,I147299,I147317,I147335,I147353,I147371,I147398,I147407,I147425,I147443,I147470,I147488,I147506,I147515,I147533,I147560,I147569,I147587,I147614,I147623,I147641,I147659,I147677,I147704,I147713,I147731,I147749,I147767,I147785,I147803,I147830,I147839,I147866,I147875,I147893,I147911,I147929,I147956,I147965,I147992,I148010,I148019,I148037,I148055,I148073,I148100,I148109,I148127,I148145,I148172,I148181,I148199,I148217,I148235,I148253,I148280,I148298,I148307,I148325,I148343,I148361,I148388,I148397,I148415,I148433,I148451,I148469,I148487,I148505,I148523,I148541,I148568,I148577,I148595,I148622,I148631,I148649,I148676,I148685,I148703,I148730,I148739,I148757,I148775,I148802,I148820,I148829,I148847,I148865,I148883,I148901,I148928,I148937,I148964,I148982,I148991,I149009,I149027,I149045,I149063,I149090,I149099,I149126,I149144,I149153,I149171,I149189,I149207,I149225,I149243,I149270,I149279,I149297,I149324,I149333,I149351,I149369,I149396,I149405,I149423,I149450,I149459,I149477,I149495,I149513,I149531,I149549,I149567,I149585,I149612,I149621,I149639,I149657,I149675,I149693,I149711,I149729,I149747,I149765,I149783,I149810,I149819,I149837,I149855,I149882,I149900,I149909,I149927,I149954,I149963,I149981,I149999,I150026,I150044,I150053,I150071,I150098,I150116,I150125,I150143,I150161,I150179,I150197,I150215,I150233,I150260,I150269,I150287,I150305,I150323,I150341,I150368,I150377,I150395,I150413,I150440,I150449,I150476,I150485,I150503,I150521,I150539,I150557,I150584,I150593,I150611,I150629,I150647,I150674,I150683,I150701,I150728,I150737,I150764,I150773,I150791,I150809,I150827,I150854,I150863,I150881,I150899,I150917,I150944,I150953,I150980,I150998,I151007,I151025,I151043,I151061,I151088,I151097,I151124,I151133,I151151,I151169,I151196,I151205,I151232,I151241,I151259,I151277,I151304,I151313,I151331,I151349,I151367,I151394,I151403,I151421,I151439,I151457,I151475,I151502,I151520,I151529,I151556,I151565,I151583,I151601,I151628,I151646,I151664,I151673,I151691,I151718,I151727,I151745,I151772,I151781,I151799,I151817,I151835,I151862,I151871,I151889,I151907,I151925,I151943,I151961,I151988,I151997,I152024,I152033,I152051,I152069,I152087,I152114,I152132,I152141,I152159,I152186,I152195,I152213,I152231,I152249,I152267,I152285,I152303,I152330,I152339,I152357,I152375,I152402,I152411,I152429,I152447,I152474,I152483,I152510,I152519,I152537,I152555,I152573,I152591,I152618,I152627,I152645,I152663,I152681,I152699,I152717,I152744,I152753,I152771,I152798,I152807,I152825,I152852,I152861,I152879,I152906,I152915,I152933,I152951,I152978,I152996,I153005,I153023,I153041,I153059,I153077,I153104,I153113,I153140,I153158,I153167,I153185,I153203,I153221,I153239,I153266,I153275,I153302,I153311,I153338,I153347,I153365,I153383,I153401,I153419,I153446,I153455,I153473,I153491,I153509,I153527,I153545,I153563,I153581,I153599,I153617,I153635,I153653,I153671,I153689,I153707,I153725,I153752,I153761,I153788,I153806,I153815,I153833,I153851,I153878,I153887,I153914,I153932,I153941,I153959,I153986,I153995,I154013,I154031,I154049,I154067,I154085,I154103,I154121,I154148,I154157,I154175,I154193,I154211,I154229,I154247,I154265,I154292,I154310,I154319,I154337,I154355,I154373,I154400,I154409,I154427,I154445,I154472,I154481,I154499,I154517,I154544,I154553,I154571,I154589,I154616,I154634,I154652,I154661,I154679,I154706,I154715,I154733,I154760,I154769,I154787,I154805,I154823,I154850,I154859,I154877,I154895,I154913,I154931,I154949,I154976,I154985,I155012,I155021,I155039,I155057,I155075,I155102,I155111,I155129,I155147,I155174,I155183,I155210,I155219,I155237,I155255,I155273,I155291,I155318,I155327,I155345,I155363,I155381,I155408,I155417,I155435,I155462,I155471,I155498,I155507,I155525,I155543,I155561,I155588,I155597,I155615,I155633,I155651,I155678,I155687,I155714,I155732,I155741,I155759,I155786,I155795,I155813,I155831,I155849,I155867,I155885,I155903,I155930,I155939,I155957,I155975,I156002,I156011,I156029,I156047,I156074,I156083,I156110,I156119,I156137,I156155,I156173,I156191,I156218,I156227,I156245,I156263,I156281,I156299,I156317,I156344,I156353,I156371,I156389,I156416,I156425,I156452,I156461,I156479,I156497,I156515,I156533,I156560,I156569,I156587,I156605,I156623,I156650,I156659,I156677,I156704,I156713,I156740,I156749,I156767,I156785,I156803,I156830,I156839,I156857,I156875,I156893,I156920,I156929,I156956,I156974,I156983,I157001,I157028,I157037,I157055,I157073,I157091,I157109,I157127,I157145,I157163,I157190,I157199,I157217,I157235,I157253,I157271,I157289,I157307,I157334,I157352,I157361,I157379,I157397,I157415,I157442,I157451,I157469,I157487,I157514,I157523,I157541,I157559,I157586,I157595,I157622,I157631,I157649,I157667,I157685,I157703,I157730,I157739,I157757,I157775,I157793,I157811,I157829,I157847,I157865,I157883,I157901,I157919,I157937,I157955,I157973,I157991,I158009,I158036,I158045,I158072,I158090,I158099,I158117,I158135,I158162,I158171,I158198,I158207,I158225,I158243,I158270,I158279,I158306,I158315,I158333,I158351,I158369,I158387,I158414,I158423,I158441,I158459,I158477,I158504,I158513,I158531,I158558,I158567,I158594,I158603,I158621,I158639,I158657,I158684,I158693,I158711,I158729,I158747,I158774,I158783,I158810,I158828,I158837,I158855,I158882,I158891,I158909,I158927,I158945,I158963,I158981,I158999,I159026,I159035,I159053,I159071,I159098,I159107,I159125,I159143,I159170,I159179,I159206,I159215,I159233,I159251,I159269,I159287,I159314,I159323,I159341,I159359,I159377,I159395,I159413,I159440,I159449,I159467,I159485,I159512,I159530,I159539,I159557,I159584,I159593,I159611,I159629,I159656,I159674,I159683,I159701,I159728,I159746,I159755,I159773,I159791,I159809,I159827,I159845,I159863,I159890,I159899,I159917,I159935,I159953,I159971,I159998,I160007,I160034,I160052,I160061,I160079,I160097,I160115,I160142,I160151,I160169,I160187,I160214,I160223,I160241,I160259,I160277,I160295,I160322,I160340,I160349,I160367,I160385,I160403,I160430,I160439,I160457,I160475,I160493,I160511,I160529,I160547,I160565,I160583,I160610,I160628,I160637,I160655,I160682,I160691,I160709,I160727,I160745,I160763,I160781,I160799,I160826,I160835,I160853,I160871,I160898,I160907,I160925,I160943,I160970,I160979,I161006,I161015,I161033,I161051,I161069,I161087,I161114,I161123,I161141,I161159,I161177,I161195,I161213,I161240,I161249,I161267,I161294,I161312,I161321,I161339,I161357,I161375,I161393,I161420,I161429,I161447,I161465,I161483,I161501,I161519,I161537,I161555,I161573,I161591,I161609,I161627,I161645,I161663,I161690,I161699,I161726,I161735,I161762,I161771,I161789,I161807,I161825,I161843,I161870,I161879,I161897,I161915,I161942,I161951,I161978,I161987,I162005,I162023,I162041,I162059,I162086,I162095,I162113,I162131,I162149,I162176,I162185,I162203,I162230,I162239,I162266,I162275,I162293,I162311,I162329,I162356,I162365,I162383,I162401,I162419,I162446,I162455,I162482,I162500,I162509,I162527,I162545,I162563,I162590,I162599,I162626,I162635,I162653,I162671,I162698,I162707,I162734,I162743,I162761,I162779,I162806,I162815,I162833,I162851,I162869,I162896,I162905,I162923,I162941,I162959,I162977,I163004,I163022,I163031,I163058,I163067,I163085,I163103,I163130,I163148,I163157,I163175,I163202,I163211,I163229,I163247,I163274,I163292,I163301,I163319,I163346,I163364,I163373,I163391,I163409,I163427,I163445,I163463,I163481,I163508,I163517,I163535,I163553,I163571,I163589,I163616,I163625,I163652,I163670,I163679,I163697,I163715,I163733,I163751,I163769,I163787,I163805,I163823,I163841,I163859,I163877,I163904,I163913,I163931,I163949,I163976,I163985,I164003,I164021,I164048,I164057,I164075,I164093,I164120,I164129,I164147,I164165,I164192,I164201,I164219,I164237,I164264,I164273,I164300,I164309,I164327,I164345,I164363,I164408,I164417,I164435,I164453,I164471,I164507,I164525,I164552,I164561,I164597,I164633,I164651,I164687;
not I_0 (I707,I698);
DFFARX1 I_1 (I116,I691,I707,I734,);
DFFARX1 I_2 (I734,I691,I707,I752,);
not I_3 (I761,I752);
not I_4 (I779,I734);
DFFARX1 I_5 (I108,I691,I707,I806,);
not I_6 (I815,I806);
and I_7 (I833,I779,I500);
not I_8 (I851,I164);
nand I_9 (I869,I851,I500);
not I_10 (I887,I468);
nor I_11 (I905,I887,I348);
nand I_12 (I923,I905,I516);
nor I_13 (I941,I923,I869);
DFFARX1 I_14 (I941,I691,I707,I968,);
not I_15 (I977,I923);
not I_16 (I995,I348);
nand I_17 (I1013,I995,I500);
nor I_18 (I1031,I348,I164);
nand I_19 (I1049,I833,I1031);
nand I_20 (I1067,I779,I348);
nand I_21 (I1085,I887,I508);
DFFARX1 I_22 (I1085,I691,I707,I1112,);
DFFARX1 I_23 (I1085,I691,I707,I1130,);
not I_24 (I1139,I508);
nor I_25 (I1157,I1139,I132);
and I_26 (I1175,I1157,I492);
or I_27 (I1193,I1175,I332);
DFFARX1 I_28 (I1193,I691,I707,I1220,);
nand I_29 (I1229,I1220,I851);
nor I_30 (I1247,I1229,I1013);
nor I_31 (I1265,I1220,I815);
DFFARX1 I_32 (I1220,I691,I707,I1292,);
not I_33 (I1301,I1292);
nor I_34 (I1319,I1301,I977);
not I_35 (I1337,I698);
DFFARX1 I_36 (I1049,I691,I1337,I1364,);
not I_37 (I1373,I1364);
nand I_38 (I1391,I1067,I968);
and I_39 (I1409,I1391,I1112);
DFFARX1 I_40 (I1409,I691,I1337,I1436,);
DFFARX1 I_41 (I1319,I691,I1337,I1454,);
and I_42 (I1463,I1454,I1130);
nor I_43 (I1481,I1436,I1463);
DFFARX1 I_44 (I1481,I691,I1337,I1508,);
nand I_45 (I1517,I1454,I1130);
nand I_46 (I1535,I1373,I1517);
not I_47 (I1553,I1535);
DFFARX1 I_48 (I968,I691,I1337,I1580,);
DFFARX1 I_49 (I1580,I691,I1337,I1598,);
nand I_50 (I1607,I1265,I1265);
and I_51 (I1625,I1607,I761);
DFFARX1 I_52 (I1625,I691,I1337,I1652,);
DFFARX1 I_53 (I1652,I691,I1337,I1670,);
not I_54 (I1679,I1670);
not I_55 (I1697,I1652);
nand I_56 (I1715,I1697,I1517);
nor I_57 (I1733,I1247,I1265);
not I_58 (I1751,I1733);
nor I_59 (I1769,I1697,I1751);
nor I_60 (I1787,I1373,I1769);
DFFARX1 I_61 (I1787,I691,I1337,I1814,);
nor I_62 (I1823,I1436,I1751);
nor I_63 (I1841,I1652,I1823);
nor I_64 (I1859,I1580,I1733);
nor I_65 (I1877,I1436,I1733);
not I_66 (I1895,I698);
DFFARX1 I_67 (I1598,I691,I1895,I1922,);
DFFARX1 I_68 (I1715,I691,I1895,I1940,);
not I_69 (I1949,I1940);
nor I_70 (I1967,I1922,I1949);
DFFARX1 I_71 (I1949,I691,I1895,I1994,);
nor I_72 (I2003,I1508,I1679);
and I_73 (I2021,I2003,I1877);
nor I_74 (I2039,I2021,I1508);
not I_75 (I2057,I1508);
and I_76 (I2075,I2057,I1841);
nand I_77 (I2093,I2075,I1814);
nor I_78 (I2111,I2057,I2093);
DFFARX1 I_79 (I2111,I691,I1895,I2138,);
not I_80 (I2147,I2093);
nand I_81 (I2165,I1949,I2147);
nand I_82 (I2183,I2021,I2147);
DFFARX1 I_83 (I2057,I691,I1895,I2210,);
not I_84 (I2219,I1508);
nor I_85 (I2237,I2219,I1841);
nor I_86 (I2255,I2237,I2039);
DFFARX1 I_87 (I2255,I691,I1895,I2282,);
not I_88 (I2291,I2237);
DFFARX1 I_89 (I2291,I691,I1895,I2318,);
not I_90 (I2327,I2318);
nor I_91 (I2345,I2327,I2237);
nor I_92 (I2363,I2219,I1877);
and I_93 (I2381,I2363,I1553);
or I_94 (I2399,I2381,I1859);
DFFARX1 I_95 (I2399,I691,I1895,I2426,);
not I_96 (I2435,I2426);
nand I_97 (I2453,I2435,I2147);
not I_98 (I2471,I2453);
nand I_99 (I2489,I2453,I2165);
nand I_100 (I2507,I2435,I2021);
not I_101 (I2525,I698);
DFFARX1 I_102 (I2210,I691,I2525,I2552,);
and I_103 (I2561,I2552,I2489);
DFFARX1 I_104 (I2561,I691,I2525,I2588,);
DFFARX1 I_105 (I2138,I691,I2525,I2606,);
not I_106 (I2615,I2471);
not I_107 (I2633,I1967);
nand I_108 (I2651,I2633,I2615);
nor I_109 (I2669,I2606,I2651);
DFFARX1 I_110 (I2651,I691,I2525,I2696,);
not I_111 (I2705,I2696);
not I_112 (I2723,I2183);
nand I_113 (I2741,I2633,I2723);
DFFARX1 I_114 (I2741,I691,I2525,I2768,);
not I_115 (I2777,I2768);
not I_116 (I2795,I2345);
nand I_117 (I2813,I2795,I2138);
and I_118 (I2831,I2615,I2813);
nor I_119 (I2849,I2741,I2831);
DFFARX1 I_120 (I2849,I691,I2525,I2876,);
DFFARX1 I_121 (I2831,I691,I2525,I2894,);
nor I_122 (I2903,I2345,I2282);
nor I_123 (I2921,I2741,I2903);
or I_124 (I2939,I2345,I2282);
nor I_125 (I2957,I1994,I2507);
DFFARX1 I_126 (I2957,I691,I2525,I2984,);
not I_127 (I2993,I2984);
nor I_128 (I3011,I2993,I2777);
nand I_129 (I3029,I2993,I2606);
not I_130 (I3047,I1994);
nand I_131 (I3065,I3047,I2723);
nand I_132 (I3083,I2993,I3065);
nand I_133 (I3101,I3083,I3029);
nand I_134 (I3119,I3065,I2939);
not I_135 (I3137,I698);
DFFARX1 I_136 (I2876,I691,I3137,I3164,);
nand I_137 (I3173,I2588,I2876);
and I_138 (I3191,I3173,I3011);
DFFARX1 I_139 (I3191,I691,I3137,I3218,);
nor I_140 (I3227,I3218,I3164);
not I_141 (I3245,I3218);
DFFARX1 I_142 (I2705,I691,I3137,I3272,);
nand I_143 (I3281,I3272,I3119);
not I_144 (I3299,I3281);
DFFARX1 I_145 (I3299,I691,I3137,I3326,);
not I_146 (I3335,I3326);
nor I_147 (I3353,I3164,I3281);
nor I_148 (I3371,I3218,I3353);
DFFARX1 I_149 (I2669,I691,I3137,I3398,);
DFFARX1 I_150 (I3398,I691,I3137,I3416,);
not I_151 (I3425,I3416);
not I_152 (I3443,I3398);
nand I_153 (I3461,I3443,I3245);
nand I_154 (I3479,I2669,I3101);
and I_155 (I3497,I3479,I2894);
DFFARX1 I_156 (I3497,I691,I3137,I3524,);
nor I_157 (I3533,I3524,I3164);
DFFARX1 I_158 (I3533,I691,I3137,I3560,);
DFFARX1 I_159 (I3524,I691,I3137,I3578,);
nor I_160 (I3587,I2921,I3101);
not I_161 (I3605,I3587);
nor I_162 (I3623,I3425,I3605);
nand I_163 (I3641,I3443,I3605);
nor I_164 (I3659,I3164,I3587);
DFFARX1 I_165 (I3587,I691,I3137,I3686,);
not I_166 (I3695,I698);
DFFARX1 I_167 (I3623,I691,I3695,I3722,);
DFFARX1 I_168 (I3722,I691,I3695,I3740,);
not I_169 (I3749,I3740);
not I_170 (I3767,I3722);
DFFARX1 I_171 (I3578,I691,I3695,I3794,);
nand I_172 (I3803,I3794,I3461);
not I_173 (I3821,I3461);
not I_174 (I3839,I3371);
nand I_175 (I3857,I3227,I3560);
and I_176 (I3875,I3227,I3560);
not I_177 (I3893,I3659);
nand I_178 (I3911,I3893,I3839);
nor I_179 (I3929,I3911,I3803);
nor I_180 (I3947,I3821,I3911);
nand I_181 (I3965,I3875,I3947);
not I_182 (I3983,I3335);
nor I_183 (I4001,I3983,I3227);
nor I_184 (I4019,I4001,I3659);
nor I_185 (I4037,I3767,I4019);
DFFARX1 I_186 (I4037,I691,I3695,I4064,);
not I_187 (I4073,I4001);
DFFARX1 I_188 (I4073,I691,I3695,I4100,);
and I_189 (I4109,I3794,I4001);
nor I_190 (I4127,I3983,I3686);
and I_191 (I4145,I4127,I3560);
or I_192 (I4163,I4145,I3641);
DFFARX1 I_193 (I4163,I691,I3695,I4190,);
nor I_194 (I4199,I4190,I3893);
DFFARX1 I_195 (I4199,I691,I3695,I4226,);
nand I_196 (I4235,I4190,I3794);
nand I_197 (I4253,I3893,I4235);
nor I_198 (I4271,I4253,I3857);
not I_199 (I4289,I698);
DFFARX1 I_200 (I4271,I691,I4289,I4316,);
not I_201 (I4325,I4316);
nand I_202 (I4343,I4100,I3965);
and I_203 (I4361,I4343,I3929);
DFFARX1 I_204 (I4361,I691,I4289,I4388,);
DFFARX1 I_205 (I4388,I691,I4289,I4406,);
DFFARX1 I_206 (I3929,I691,I4289,I4424,);
nand I_207 (I4433,I4424,I4226);
not I_208 (I4451,I4433);
DFFARX1 I_209 (I4451,I691,I4289,I4478,);
not I_210 (I4487,I4478);
nor I_211 (I4505,I4325,I4487);
DFFARX1 I_212 (I3965,I691,I4289,I4532,);
nor I_213 (I4541,I4532,I4388);
nor I_214 (I4559,I4532,I4451);
nand I_215 (I4577,I3749,I4109);
and I_216 (I4595,I4577,I4064);
DFFARX1 I_217 (I4595,I691,I4289,I4622,);
not I_218 (I4631,I4622);
nand I_219 (I4649,I4631,I4532);
nand I_220 (I4667,I4631,I4433);
nor I_221 (I4685,I4226,I4109);
and I_222 (I4703,I4532,I4685);
nor I_223 (I4721,I4631,I4703);
DFFARX1 I_224 (I4721,I691,I4289,I4748,);
nor I_225 (I4757,I4316,I4685);
DFFARX1 I_226 (I4757,I691,I4289,I4784,);
nor I_227 (I4793,I4622,I4685);
not I_228 (I4811,I4793);
nand I_229 (I4829,I4811,I4649);
not I_230 (I4847,I698);
DFFARX1 I_231 (I4748,I691,I4847,I4874,);
not I_232 (I4883,I4874);
nand I_233 (I4901,I4559,I4505);
and I_234 (I4919,I4901,I4406);
DFFARX1 I_235 (I4919,I691,I4847,I4946,);
not I_236 (I4955,I4829);
DFFARX1 I_237 (I4667,I691,I4847,I4982,);
not I_238 (I4991,I4982);
nor I_239 (I5009,I4991,I4883);
and I_240 (I5027,I5009,I4829);
nor I_241 (I5045,I4991,I4955);
nor I_242 (I5063,I4946,I5045);
DFFARX1 I_243 (I4784,I691,I4847,I5090,);
nor I_244 (I5099,I5090,I4946);
not I_245 (I5117,I5099);
not I_246 (I5135,I5090);
nor I_247 (I5153,I5135,I5027);
DFFARX1 I_248 (I5153,I691,I4847,I5180,);
nand I_249 (I5189,I4784,I4559);
and I_250 (I5207,I5189,I4667);
DFFARX1 I_251 (I5207,I691,I4847,I5234,);
nor I_252 (I5243,I5234,I5090);
DFFARX1 I_253 (I5243,I691,I4847,I5270,);
nand I_254 (I5279,I5234,I5135);
nand I_255 (I5297,I5117,I5279);
not I_256 (I5315,I5234);
nor I_257 (I5333,I5315,I5027);
DFFARX1 I_258 (I5333,I691,I4847,I5360,);
nor I_259 (I5369,I4541,I4559);
or I_260 (I5387,I5090,I5369);
nor I_261 (I5405,I5234,I5369);
or I_262 (I5423,I4946,I5369);
DFFARX1 I_263 (I5369,I691,I4847,I5450,);
not I_264 (I5459,I698);
DFFARX1 I_265 (I5270,I691,I5459,I5486,);
not I_266 (I5495,I5486);
DFFARX1 I_267 (I5387,I691,I5459,I5522,);
not I_268 (I5531,I5405);
nand I_269 (I5549,I5531,I5423);
not I_270 (I5567,I5549);
nor I_271 (I5585,I5567,I5297);
nor I_272 (I5603,I5495,I5585);
DFFARX1 I_273 (I5603,I691,I5459,I5630,);
not I_274 (I5639,I5297);
nand I_275 (I5657,I5639,I5567);
and I_276 (I5675,I5639,I5405);
nand I_277 (I5693,I5675,I5063);
nor I_278 (I5711,I5693,I5639);
and I_279 (I5729,I5522,I5693);
not I_280 (I5747,I5693);
nand I_281 (I5765,I5522,I5747);
nor I_282 (I5783,I5486,I5693);
not I_283 (I5801,I5360);
nor I_284 (I5819,I5801,I5405);
nand I_285 (I5837,I5819,I5639);
nor I_286 (I5855,I5549,I5837);
nor I_287 (I5873,I5801,I5270);
and I_288 (I5891,I5873,I5180);
or I_289 (I5909,I5891,I5450);
DFFARX1 I_290 (I5909,I691,I5459,I5936,);
nor I_291 (I5945,I5936,I5657);
DFFARX1 I_292 (I5945,I691,I5459,I5972,);
DFFARX1 I_293 (I5936,I691,I5459,I5990,);
not I_294 (I5999,I5936);
nor I_295 (I6017,I5999,I5522);
nor I_296 (I6035,I5819,I6017);
DFFARX1 I_297 (I6035,I691,I5459,I6062,);
not I_298 (I6071,I698);
DFFARX1 I_299 (I5783,I691,I6071,I6098,);
DFFARX1 I_300 (I6098,I691,I6071,I6116,);
not I_301 (I6125,I6116);
not I_302 (I6143,I6098);
nand I_303 (I6161,I5972,I6062);
and I_304 (I6179,I6161,I5990);
DFFARX1 I_305 (I6179,I691,I6071,I6206,);
not I_306 (I6215,I6206);
DFFARX1 I_307 (I5765,I691,I6071,I6242,);
and I_308 (I6251,I6242,I5855);
nand I_309 (I6269,I6242,I5855);
nand I_310 (I6287,I6215,I6269);
DFFARX1 I_311 (I5711,I691,I6071,I6314,);
nor I_312 (I6323,I6314,I6251);
DFFARX1 I_313 (I6323,I691,I6071,I6350,);
nor I_314 (I6359,I6314,I6206);
nand I_315 (I6377,I5972,I5729);
and I_316 (I6395,I6377,I5630);
DFFARX1 I_317 (I6395,I691,I6071,I6422,);
nor I_318 (I6431,I6422,I6314);
not I_319 (I6449,I6422);
nor I_320 (I6467,I6449,I6215);
nor I_321 (I6485,I6143,I6467);
DFFARX1 I_322 (I6485,I691,I6071,I6512,);
nor I_323 (I6521,I6449,I6314);
nor I_324 (I6539,I5783,I5729);
nor I_325 (I6557,I6539,I6521);
not I_326 (I6575,I6539);
nand I_327 (I6593,I6269,I6575);
DFFARX1 I_328 (I6539,I691,I6071,I6620,);
DFFARX1 I_329 (I6539,I691,I6071,I6638,);
not I_330 (I6647,I698);
DFFARX1 I_331 (I6557,I691,I6647,I6674,);
not I_332 (I6683,I6674);
nand I_333 (I6701,I6350,I6512);
and I_334 (I6719,I6701,I6638);
DFFARX1 I_335 (I6719,I691,I6647,I6746,);
not I_336 (I6755,I6359);
DFFARX1 I_337 (I6431,I691,I6647,I6782,);
not I_338 (I6791,I6782);
nor I_339 (I6809,I6791,I6683);
and I_340 (I6827,I6809,I6359);
nor I_341 (I6845,I6791,I6755);
nor I_342 (I6863,I6746,I6845);
DFFARX1 I_343 (I6593,I691,I6647,I6890,);
nor I_344 (I6899,I6890,I6746);
not I_345 (I6917,I6899);
not I_346 (I6935,I6890);
nor I_347 (I6953,I6935,I6827);
DFFARX1 I_348 (I6953,I691,I6647,I6980,);
nand I_349 (I6989,I6125,I6620);
and I_350 (I7007,I6989,I6287);
DFFARX1 I_351 (I7007,I691,I6647,I7034,);
nor I_352 (I7043,I7034,I6890);
DFFARX1 I_353 (I7043,I691,I6647,I7070,);
nand I_354 (I7079,I7034,I6935);
nand I_355 (I7097,I6917,I7079);
not I_356 (I7115,I7034);
nor I_357 (I7133,I7115,I6827);
DFFARX1 I_358 (I7133,I691,I6647,I7160,);
nor I_359 (I7169,I6350,I6620);
or I_360 (I7187,I6890,I7169);
nor I_361 (I7205,I7034,I7169);
or I_362 (I7223,I6746,I7169);
DFFARX1 I_363 (I7169,I691,I6647,I7250,);
not I_364 (I7259,I698);
DFFARX1 I_365 (I7223,I691,I7259,I7286,);
DFFARX1 I_366 (I7286,I691,I7259,I7304,);
not I_367 (I7313,I7304);
nand I_368 (I7331,I7160,I7250);
and I_369 (I7349,I7331,I7205);
DFFARX1 I_370 (I7349,I691,I7259,I7376,);
DFFARX1 I_371 (I7376,I691,I7259,I7394,);
DFFARX1 I_372 (I7376,I691,I7259,I7412,);
DFFARX1 I_373 (I7097,I691,I7259,I7430,);
nand I_374 (I7439,I7430,I6863);
not I_375 (I7457,I7439);
nor I_376 (I7475,I7286,I7457);
DFFARX1 I_377 (I7205,I691,I7259,I7502,);
not I_378 (I7511,I7502);
nor I_379 (I7529,I7511,I7313);
nand I_380 (I7547,I7511,I7439);
nand I_381 (I7565,I6980,I7070);
and I_382 (I7583,I7565,I7187);
DFFARX1 I_383 (I7583,I691,I7259,I7610,);
nor I_384 (I7619,I7610,I7286);
DFFARX1 I_385 (I7619,I691,I7259,I7646,);
not I_386 (I7655,I7610);
nor I_387 (I7673,I7070,I7070);
not I_388 (I7691,I7673);
nor I_389 (I7709,I7439,I7691);
nor I_390 (I7727,I7655,I7709);
DFFARX1 I_391 (I7727,I691,I7259,I7754,);
nor I_392 (I7763,I7610,I7691);
nor I_393 (I7781,I7457,I7763);
nor I_394 (I7799,I7610,I7673);
not I_395 (I7817,I698);
DFFARX1 I_396 (I7475,I691,I7817,I7844,);
not I_397 (I7853,I7844);
nand I_398 (I7871,I7781,I7646);
and I_399 (I7889,I7871,I7646);
DFFARX1 I_400 (I7889,I691,I7817,I7916,);
not I_401 (I7925,I7799);
DFFARX1 I_402 (I7529,I691,I7817,I7952,);
not I_403 (I7961,I7952);
nor I_404 (I7979,I7961,I7853);
and I_405 (I7997,I7979,I7799);
nor I_406 (I8015,I7961,I7925);
nor I_407 (I8033,I7916,I8015);
DFFARX1 I_408 (I7799,I691,I7817,I8060,);
nor I_409 (I8069,I8060,I7916);
not I_410 (I8087,I8069);
not I_411 (I8105,I8060);
nor I_412 (I8123,I8105,I7997);
DFFARX1 I_413 (I8123,I691,I7817,I8150,);
nand I_414 (I8159,I7754,I7547);
and I_415 (I8177,I8159,I7412);
DFFARX1 I_416 (I8177,I691,I7817,I8204,);
nor I_417 (I8213,I8204,I8060);
DFFARX1 I_418 (I8213,I691,I7817,I8240,);
nand I_419 (I8249,I8204,I8105);
nand I_420 (I8267,I8087,I8249);
not I_421 (I8285,I8204);
nor I_422 (I8303,I8285,I7997);
DFFARX1 I_423 (I8303,I691,I7817,I8330,);
nor I_424 (I8339,I7394,I7547);
or I_425 (I8357,I8060,I8339);
nor I_426 (I8375,I8204,I8339);
or I_427 (I8393,I7916,I8339);
DFFARX1 I_428 (I8339,I691,I7817,I8420,);
not I_429 (I8429,I698);
DFFARX1 I_430 (I8393,I691,I8429,I8456,);
DFFARX1 I_431 (I8240,I691,I8429,I8474,);
not I_432 (I8483,I8474);
not I_433 (I8501,I8033);
nor I_434 (I8519,I8501,I8240);
not I_435 (I8537,I8267);
nor I_436 (I8555,I8519,I8150);
nor I_437 (I8573,I8474,I8555);
DFFARX1 I_438 (I8573,I691,I8429,I8600,);
nor I_439 (I8609,I8150,I8240);
nand I_440 (I8627,I8609,I8033);
DFFARX1 I_441 (I8627,I691,I8429,I8654,);
nor I_442 (I8663,I8537,I8150);
nand I_443 (I8681,I8663,I8375);
nor I_444 (I8699,I8456,I8681);
DFFARX1 I_445 (I8699,I691,I8429,I8726,);
not I_446 (I8735,I8681);
nand I_447 (I8753,I8474,I8735);
DFFARX1 I_448 (I8681,I691,I8429,I8780,);
not I_449 (I8789,I8780);
not I_450 (I8807,I8150);
not I_451 (I8825,I8357);
nor I_452 (I8843,I8825,I8267);
nor I_453 (I8861,I8789,I8843);
nor I_454 (I8879,I8825,I8330);
and I_455 (I8897,I8879,I8420);
or I_456 (I8915,I8897,I8375);
DFFARX1 I_457 (I8915,I691,I8429,I8942,);
nor I_458 (I8951,I8942,I8456);
not I_459 (I8969,I8942);
and I_460 (I8987,I8969,I8456);
nor I_461 (I9005,I8483,I8987);
nand I_462 (I9023,I8969,I8537);
nor I_463 (I9041,I8825,I9023);
nand I_464 (I9059,I8969,I8735);
nand I_465 (I9077,I8537,I8357);
nor I_466 (I9095,I8807,I9077);
not I_467 (I9113,I698);
DFFARX1 I_468 (I8654,I691,I9113,I9140,);
DFFARX1 I_469 (I9140,I691,I9113,I9158,);
not I_470 (I9167,I9158);
nand I_471 (I9185,I8726,I8861);
and I_472 (I9203,I9185,I8753);
DFFARX1 I_473 (I9203,I691,I9113,I9230,);
DFFARX1 I_474 (I9230,I691,I9113,I9248,);
DFFARX1 I_475 (I9230,I691,I9113,I9266,);
DFFARX1 I_476 (I9095,I691,I9113,I9284,);
nand I_477 (I9293,I9284,I9041);
not I_478 (I9311,I9293);
nor I_479 (I9329,I9140,I9311);
DFFARX1 I_480 (I8600,I691,I9113,I9356,);
not I_481 (I9365,I9356);
nor I_482 (I9383,I9365,I9167);
nand I_483 (I9401,I9365,I9293);
nand I_484 (I9419,I9059,I9005);
and I_485 (I9437,I9419,I8726);
DFFARX1 I_486 (I9437,I691,I9113,I9464,);
nor I_487 (I9473,I9464,I9140);
DFFARX1 I_488 (I9473,I691,I9113,I9500,);
not I_489 (I9509,I9464);
nor I_490 (I9527,I8951,I9005);
not I_491 (I9545,I9527);
nor I_492 (I9563,I9293,I9545);
nor I_493 (I9581,I9509,I9563);
DFFARX1 I_494 (I9581,I691,I9113,I9608,);
nor I_495 (I9617,I9464,I9545);
nor I_496 (I9635,I9311,I9617);
nor I_497 (I9653,I9464,I9527);
not I_498 (I9671,I698);
DFFARX1 I_499 (I9653,I691,I9671,I9698,);
not I_500 (I9707,I9698);
DFFARX1 I_501 (I9401,I691,I9671,I9734,);
not I_502 (I9743,I9500);
nand I_503 (I9761,I9743,I9248);
not I_504 (I9779,I9761);
nor I_505 (I9797,I9779,I9653);
nor I_506 (I9815,I9707,I9797);
DFFARX1 I_507 (I9815,I691,I9671,I9842,);
not I_508 (I9851,I9653);
nand I_509 (I9869,I9851,I9779);
and I_510 (I9887,I9851,I9383);
nand I_511 (I9905,I9887,I9329);
nor I_512 (I9923,I9905,I9851);
and I_513 (I9941,I9734,I9905);
not I_514 (I9959,I9905);
nand I_515 (I9977,I9734,I9959);
nor I_516 (I9995,I9698,I9905);
not I_517 (I10013,I9608);
nor I_518 (I10031,I10013,I9383);
nand I_519 (I10049,I10031,I9851);
nor I_520 (I10067,I9761,I10049);
nor I_521 (I10085,I10013,I9500);
and I_522 (I10103,I10085,I9635);
or I_523 (I10121,I10103,I9266);
DFFARX1 I_524 (I10121,I691,I9671,I10148,);
nor I_525 (I10157,I10148,I9869);
DFFARX1 I_526 (I10157,I691,I9671,I10184,);
DFFARX1 I_527 (I10148,I691,I9671,I10202,);
not I_528 (I10211,I10148);
nor I_529 (I10229,I10211,I9734);
nor I_530 (I10247,I10031,I10229);
DFFARX1 I_531 (I10247,I691,I9671,I10274,);
not I_532 (I10283,I698);
DFFARX1 I_533 (I9923,I691,I10283,I10310,);
DFFARX1 I_534 (I10310,I691,I10283,I10328,);
not I_535 (I10337,I10328);
not I_536 (I10355,I10310);
DFFARX1 I_537 (I9941,I691,I10283,I10382,);
not I_538 (I10391,I10382);
and I_539 (I10409,I10355,I10202);
not I_540 (I10427,I10274);
nand I_541 (I10445,I10427,I10202);
not I_542 (I10463,I10184);
nor I_543 (I10481,I10463,I9995);
nand I_544 (I10499,I10481,I10067);
nor I_545 (I10517,I10499,I10445);
DFFARX1 I_546 (I10517,I691,I10283,I10544,);
not I_547 (I10553,I10499);
not I_548 (I10571,I9995);
nand I_549 (I10589,I10571,I10202);
nor I_550 (I10607,I9995,I10274);
nand I_551 (I10625,I10409,I10607);
nand I_552 (I10643,I10355,I9995);
nand I_553 (I10661,I10463,I9842);
DFFARX1 I_554 (I10661,I691,I10283,I10688,);
DFFARX1 I_555 (I10661,I691,I10283,I10706,);
not I_556 (I10715,I9842);
nor I_557 (I10733,I10715,I10184);
and I_558 (I10751,I10733,I9977);
or I_559 (I10769,I10751,I9995);
DFFARX1 I_560 (I10769,I691,I10283,I10796,);
nand I_561 (I10805,I10796,I10427);
nor I_562 (I10823,I10805,I10589);
nor I_563 (I10841,I10796,I10391);
DFFARX1 I_564 (I10796,I691,I10283,I10868,);
not I_565 (I10877,I10868);
nor I_566 (I10895,I10877,I10553);
not I_567 (I10913,I698);
DFFARX1 I_568 (I10544,I691,I10913,I10940,);
and I_569 (I10949,I10940,I10841);
DFFARX1 I_570 (I10949,I691,I10913,I10976,);
DFFARX1 I_571 (I10841,I691,I10913,I10994,);
not I_572 (I11003,I10895);
not I_573 (I11021,I10337);
nand I_574 (I11039,I11021,I11003);
nor I_575 (I11057,I10994,I11039);
DFFARX1 I_576 (I11039,I691,I10913,I11084,);
not I_577 (I11093,I11084);
not I_578 (I11111,I10625);
nand I_579 (I11129,I11021,I11111);
DFFARX1 I_580 (I11129,I691,I10913,I11156,);
not I_581 (I11165,I11156);
not I_582 (I11183,I10823);
nand I_583 (I11201,I11183,I10643);
and I_584 (I11219,I11003,I11201);
nor I_585 (I11237,I11129,I11219);
DFFARX1 I_586 (I11237,I691,I10913,I11264,);
DFFARX1 I_587 (I11219,I691,I10913,I11282,);
nor I_588 (I11291,I10823,I10544);
nor I_589 (I11309,I11129,I11291);
or I_590 (I11327,I10823,I10544);
nor I_591 (I11345,I10706,I10688);
DFFARX1 I_592 (I11345,I691,I10913,I11372,);
not I_593 (I11381,I11372);
nor I_594 (I11399,I11381,I11165);
nand I_595 (I11417,I11381,I10994);
not I_596 (I11435,I10706);
nand I_597 (I11453,I11435,I11111);
nand I_598 (I11471,I11381,I11453);
nand I_599 (I11489,I11471,I11417);
nand I_600 (I11507,I11453,I11327);
not I_601 (I11525,I698);
DFFARX1 I_602 (I11264,I691,I11525,I11552,);
not I_603 (I11561,I11552);
DFFARX1 I_604 (I11507,I691,I11525,I11588,);
not I_605 (I11597,I11264);
nand I_606 (I11615,I11597,I11057);
not I_607 (I11633,I11615);
nor I_608 (I11651,I11633,I11282);
nor I_609 (I11669,I11561,I11651);
DFFARX1 I_610 (I11669,I691,I11525,I11696,);
not I_611 (I11705,I11282);
nand I_612 (I11723,I11705,I11633);
and I_613 (I11741,I11705,I11093);
nand I_614 (I11759,I11741,I11057);
nor I_615 (I11777,I11759,I11705);
and I_616 (I11795,I11588,I11759);
not I_617 (I11813,I11759);
nand I_618 (I11831,I11588,I11813);
nor I_619 (I11849,I11552,I11759);
not I_620 (I11867,I11489);
nor I_621 (I11885,I11867,I11093);
nand I_622 (I11903,I11885,I11705);
nor I_623 (I11921,I11615,I11903);
nor I_624 (I11939,I11867,I10976);
and I_625 (I11957,I11939,I11309);
or I_626 (I11975,I11957,I11399);
DFFARX1 I_627 (I11975,I691,I11525,I12002,);
nor I_628 (I12011,I12002,I11723);
DFFARX1 I_629 (I12011,I691,I11525,I12038,);
DFFARX1 I_630 (I12002,I691,I11525,I12056,);
not I_631 (I12065,I12002);
nor I_632 (I12083,I12065,I11588);
nor I_633 (I12101,I11885,I12083);
DFFARX1 I_634 (I12101,I691,I11525,I12128,);
not I_635 (I12137,I698);
DFFARX1 I_636 (I11777,I691,I12137,I12164,);
DFFARX1 I_637 (I12164,I691,I12137,I12182,);
not I_638 (I12191,I12182);
not I_639 (I12209,I12164);
DFFARX1 I_640 (I11795,I691,I12137,I12236,);
not I_641 (I12245,I12236);
and I_642 (I12263,I12209,I12056);
not I_643 (I12281,I12128);
nand I_644 (I12299,I12281,I12056);
not I_645 (I12317,I12038);
nor I_646 (I12335,I12317,I11849);
nand I_647 (I12353,I12335,I11921);
nor I_648 (I12371,I12353,I12299);
DFFARX1 I_649 (I12371,I691,I12137,I12398,);
not I_650 (I12407,I12353);
not I_651 (I12425,I11849);
nand I_652 (I12443,I12425,I12056);
nor I_653 (I12461,I11849,I12128);
nand I_654 (I12479,I12263,I12461);
nand I_655 (I12497,I12209,I11849);
nand I_656 (I12515,I12317,I11696);
DFFARX1 I_657 (I12515,I691,I12137,I12542,);
DFFARX1 I_658 (I12515,I691,I12137,I12560,);
not I_659 (I12569,I11696);
nor I_660 (I12587,I12569,I12038);
and I_661 (I12605,I12587,I11831);
or I_662 (I12623,I12605,I11849);
DFFARX1 I_663 (I12623,I691,I12137,I12650,);
nand I_664 (I12659,I12650,I12281);
nor I_665 (I12677,I12659,I12443);
nor I_666 (I12695,I12650,I12245);
DFFARX1 I_667 (I12650,I691,I12137,I12722,);
not I_668 (I12731,I12722);
nor I_669 (I12749,I12731,I12407);
not I_670 (I12767,I698);
DFFARX1 I_671 (I12497,I691,I12767,I12794,);
DFFARX1 I_672 (I12749,I691,I12767,I12812,);
not I_673 (I12821,I12812);
not I_674 (I12839,I12191);
nor I_675 (I12857,I12839,I12677);
not I_676 (I12875,I12398);
nor I_677 (I12893,I12857,I12542);
nor I_678 (I12911,I12812,I12893);
DFFARX1 I_679 (I12911,I691,I12767,I12938,);
nor I_680 (I12947,I12542,I12677);
nand I_681 (I12965,I12947,I12191);
DFFARX1 I_682 (I12965,I691,I12767,I12992,);
nor I_683 (I13001,I12875,I12542);
nand I_684 (I13019,I13001,I12695);
nor I_685 (I13037,I12794,I13019);
DFFARX1 I_686 (I13037,I691,I12767,I13064,);
not I_687 (I13073,I13019);
nand I_688 (I13091,I12812,I13073);
DFFARX1 I_689 (I13019,I691,I12767,I13118,);
not I_690 (I13127,I13118);
not I_691 (I13145,I12542);
not I_692 (I13163,I12479);
nor I_693 (I13181,I13163,I12398);
nor I_694 (I13199,I13127,I13181);
nor I_695 (I13217,I13163,I12560);
and I_696 (I13235,I13217,I12695);
or I_697 (I13253,I13235,I12398);
DFFARX1 I_698 (I13253,I691,I12767,I13280,);
nor I_699 (I13289,I13280,I12794);
not I_700 (I13307,I13280);
and I_701 (I13325,I13307,I12794);
nor I_702 (I13343,I12821,I13325);
nand I_703 (I13361,I13307,I12875);
nor I_704 (I13379,I13163,I13361);
nand I_705 (I13397,I13307,I13073);
nand I_706 (I13415,I12875,I12479);
nor I_707 (I13433,I13145,I13415);
not I_708 (I13451,I698);
DFFARX1 I_709 (I12992,I691,I13451,I13478,);
DFFARX1 I_710 (I13478,I691,I13451,I13496,);
not I_711 (I13505,I13496);
nand I_712 (I13523,I13064,I13199);
and I_713 (I13541,I13523,I13091);
DFFARX1 I_714 (I13541,I691,I13451,I13568,);
DFFARX1 I_715 (I13568,I691,I13451,I13586,);
DFFARX1 I_716 (I13568,I691,I13451,I13604,);
DFFARX1 I_717 (I13433,I691,I13451,I13622,);
nand I_718 (I13631,I13622,I13379);
not I_719 (I13649,I13631);
nor I_720 (I13667,I13478,I13649);
DFFARX1 I_721 (I12938,I691,I13451,I13694,);
not I_722 (I13703,I13694);
nor I_723 (I13721,I13703,I13505);
nand I_724 (I13739,I13703,I13631);
nand I_725 (I13757,I13397,I13343);
and I_726 (I13775,I13757,I13064);
DFFARX1 I_727 (I13775,I691,I13451,I13802,);
nor I_728 (I13811,I13802,I13478);
DFFARX1 I_729 (I13811,I691,I13451,I13838,);
not I_730 (I13847,I13802);
nor I_731 (I13865,I13289,I13343);
not I_732 (I13883,I13865);
nor I_733 (I13901,I13631,I13883);
nor I_734 (I13919,I13847,I13901);
DFFARX1 I_735 (I13919,I691,I13451,I13946,);
nor I_736 (I13955,I13802,I13883);
nor I_737 (I13973,I13649,I13955);
nor I_738 (I13991,I13802,I13865);
not I_739 (I14009,I698);
DFFARX1 I_740 (I13721,I691,I14009,I14036,);
DFFARX1 I_741 (I13838,I691,I14009,I14054,);
not I_742 (I14063,I14054);
nor I_743 (I14081,I14036,I14063);
DFFARX1 I_744 (I14063,I691,I14009,I14108,);
nor I_745 (I14117,I13838,I13604);
and I_746 (I14135,I14117,I13973);
nor I_747 (I14153,I14135,I13838);
not I_748 (I14171,I13838);
and I_749 (I14189,I14171,I13991);
nand I_750 (I14207,I14189,I13739);
nor I_751 (I14225,I14171,I14207);
DFFARX1 I_752 (I14225,I691,I14009,I14252,);
not I_753 (I14261,I14207);
nand I_754 (I14279,I14063,I14261);
nand I_755 (I14297,I14135,I14261);
DFFARX1 I_756 (I14171,I691,I14009,I14324,);
not I_757 (I14333,I13667);
nor I_758 (I14351,I14333,I13991);
nor I_759 (I14369,I14351,I14153);
DFFARX1 I_760 (I14369,I691,I14009,I14396,);
not I_761 (I14405,I14351);
DFFARX1 I_762 (I14405,I691,I14009,I14432,);
not I_763 (I14441,I14432);
nor I_764 (I14459,I14441,I14351);
nor I_765 (I14477,I14333,I13586);
and I_766 (I14495,I14477,I13946);
or I_767 (I14513,I14495,I13991);
DFFARX1 I_768 (I14513,I691,I14009,I14540,);
not I_769 (I14549,I14540);
nand I_770 (I14567,I14549,I14261);
not I_771 (I14585,I14567);
nand I_772 (I14603,I14567,I14279);
nand I_773 (I14621,I14549,I14135);
not I_774 (I14639,I698);
DFFARX1 I_775 (I14324,I691,I14639,I14666,);
DFFARX1 I_776 (I14666,I691,I14639,I14684,);
not I_777 (I14693,I14684);
not I_778 (I14711,I14666);
nand I_779 (I14729,I14081,I14396);
and I_780 (I14747,I14729,I14459);
DFFARX1 I_781 (I14747,I691,I14639,I14774,);
not I_782 (I14783,I14774);
DFFARX1 I_783 (I14252,I691,I14639,I14810,);
and I_784 (I14819,I14810,I14297);
nand I_785 (I14837,I14810,I14297);
nand I_786 (I14855,I14783,I14837);
DFFARX1 I_787 (I14585,I691,I14639,I14882,);
nor I_788 (I14891,I14882,I14819);
DFFARX1 I_789 (I14891,I691,I14639,I14918,);
nor I_790 (I14927,I14882,I14774);
nand I_791 (I14945,I14108,I14621);
and I_792 (I14963,I14945,I14603);
DFFARX1 I_793 (I14963,I691,I14639,I14990,);
nor I_794 (I14999,I14990,I14882);
not I_795 (I15017,I14990);
nor I_796 (I15035,I15017,I14783);
nor I_797 (I15053,I14711,I15035);
DFFARX1 I_798 (I15053,I691,I14639,I15080,);
nor I_799 (I15089,I15017,I14882);
nor I_800 (I15107,I14252,I14621);
nor I_801 (I15125,I15107,I15089);
not I_802 (I15143,I15107);
nand I_803 (I15161,I14837,I15143);
DFFARX1 I_804 (I15107,I691,I14639,I15188,);
DFFARX1 I_805 (I15107,I691,I14639,I15206,);
not I_806 (I15215,I698);
DFFARX1 I_807 (I15080,I691,I15215,I15242,);
not I_808 (I15251,I15242);
nand I_809 (I15269,I15161,I14999);
and I_810 (I15287,I15269,I15188);
DFFARX1 I_811 (I15287,I691,I15215,I15314,);
DFFARX1 I_812 (I14855,I691,I15215,I15332,);
and I_813 (I15341,I15332,I14918);
nor I_814 (I15359,I15314,I15341);
DFFARX1 I_815 (I15359,I691,I15215,I15386,);
nand I_816 (I15395,I15332,I14918);
nand I_817 (I15413,I15251,I15395);
not I_818 (I15431,I15413);
DFFARX1 I_819 (I14918,I691,I15215,I15458,);
DFFARX1 I_820 (I15458,I691,I15215,I15476,);
nand I_821 (I15485,I14693,I15125);
and I_822 (I15503,I15485,I14927);
DFFARX1 I_823 (I15503,I691,I15215,I15530,);
DFFARX1 I_824 (I15530,I691,I15215,I15548,);
not I_825 (I15557,I15548);
not I_826 (I15575,I15530);
nand I_827 (I15593,I15575,I15395);
nor I_828 (I15611,I15206,I15125);
not I_829 (I15629,I15611);
nor I_830 (I15647,I15575,I15629);
nor I_831 (I15665,I15251,I15647);
DFFARX1 I_832 (I15665,I691,I15215,I15692,);
nor I_833 (I15701,I15314,I15629);
nor I_834 (I15719,I15530,I15701);
nor I_835 (I15737,I15458,I15611);
nor I_836 (I15755,I15314,I15611);
not I_837 (I15773,I698);
DFFARX1 I_838 (I15476,I691,I15773,I15800,);
DFFARX1 I_839 (I15593,I691,I15773,I15818,);
not I_840 (I15827,I15818);
nor I_841 (I15845,I15800,I15827);
DFFARX1 I_842 (I15827,I691,I15773,I15872,);
nor I_843 (I15881,I15386,I15557);
and I_844 (I15899,I15881,I15755);
nor I_845 (I15917,I15899,I15386);
not I_846 (I15935,I15386);
and I_847 (I15953,I15935,I15719);
nand I_848 (I15971,I15953,I15692);
nor I_849 (I15989,I15935,I15971);
DFFARX1 I_850 (I15989,I691,I15773,I16016,);
not I_851 (I16025,I15971);
nand I_852 (I16043,I15827,I16025);
nand I_853 (I16061,I15899,I16025);
DFFARX1 I_854 (I15935,I691,I15773,I16088,);
not I_855 (I16097,I15386);
nor I_856 (I16115,I16097,I15719);
nor I_857 (I16133,I16115,I15917);
DFFARX1 I_858 (I16133,I691,I15773,I16160,);
not I_859 (I16169,I16115);
DFFARX1 I_860 (I16169,I691,I15773,I16196,);
not I_861 (I16205,I16196);
nor I_862 (I16223,I16205,I16115);
nor I_863 (I16241,I16097,I15755);
and I_864 (I16259,I16241,I15431);
or I_865 (I16277,I16259,I15737);
DFFARX1 I_866 (I16277,I691,I15773,I16304,);
not I_867 (I16313,I16304);
nand I_868 (I16331,I16313,I16025);
not I_869 (I16349,I16331);
nand I_870 (I16367,I16331,I16043);
nand I_871 (I16385,I16313,I15899);
not I_872 (I16403,I698);
DFFARX1 I_873 (I16088,I691,I16403,I16430,);
not I_874 (I16439,I16430);
nand I_875 (I16457,I16061,I16016);
and I_876 (I16475,I16457,I16349);
DFFARX1 I_877 (I16475,I691,I16403,I16502,);
not I_878 (I16511,I16016);
DFFARX1 I_879 (I15872,I691,I16403,I16538,);
not I_880 (I16547,I16538);
nor I_881 (I16565,I16547,I16439);
and I_882 (I16583,I16565,I16016);
nor I_883 (I16601,I16547,I16511);
nor I_884 (I16619,I16502,I16601);
DFFARX1 I_885 (I16385,I691,I16403,I16646,);
nor I_886 (I16655,I16646,I16502);
not I_887 (I16673,I16655);
not I_888 (I16691,I16646);
nor I_889 (I16709,I16691,I16583);
DFFARX1 I_890 (I16709,I691,I16403,I16736,);
nand I_891 (I16745,I15845,I16367);
and I_892 (I16763,I16745,I16160);
DFFARX1 I_893 (I16763,I691,I16403,I16790,);
nor I_894 (I16799,I16790,I16646);
DFFARX1 I_895 (I16799,I691,I16403,I16826,);
nand I_896 (I16835,I16790,I16691);
nand I_897 (I16853,I16673,I16835);
not I_898 (I16871,I16790);
nor I_899 (I16889,I16871,I16583);
DFFARX1 I_900 (I16889,I691,I16403,I16916,);
nor I_901 (I16925,I16223,I16367);
or I_902 (I16943,I16646,I16925);
nor I_903 (I16961,I16790,I16925);
or I_904 (I16979,I16502,I16925);
DFFARX1 I_905 (I16925,I691,I16403,I17006,);
not I_906 (I17015,I698);
DFFARX1 I_907 (I16619,I691,I17015,I17042,);
and I_908 (I17051,I17042,I16961);
DFFARX1 I_909 (I17051,I691,I17015,I17078,);
DFFARX1 I_910 (I16979,I691,I17015,I17096,);
not I_911 (I17105,I16826);
not I_912 (I17123,I17006);
nand I_913 (I17141,I17123,I17105);
nor I_914 (I17159,I17096,I17141);
DFFARX1 I_915 (I17141,I691,I17015,I17186,);
not I_916 (I17195,I17186);
not I_917 (I17213,I16943);
nand I_918 (I17231,I17123,I17213);
DFFARX1 I_919 (I17231,I691,I17015,I17258,);
not I_920 (I17267,I17258);
not I_921 (I17285,I16916);
nand I_922 (I17303,I17285,I16736);
and I_923 (I17321,I17105,I17303);
nor I_924 (I17339,I17231,I17321);
DFFARX1 I_925 (I17339,I691,I17015,I17366,);
DFFARX1 I_926 (I17321,I691,I17015,I17384,);
nor I_927 (I17393,I16916,I16853);
nor I_928 (I17411,I17231,I17393);
or I_929 (I17429,I16916,I16853);
nor I_930 (I17447,I16826,I16961);
DFFARX1 I_931 (I17447,I691,I17015,I17474,);
not I_932 (I17483,I17474);
nor I_933 (I17501,I17483,I17267);
nand I_934 (I17519,I17483,I17096);
not I_935 (I17537,I16826);
nand I_936 (I17555,I17537,I17213);
nand I_937 (I17573,I17483,I17555);
nand I_938 (I17591,I17573,I17519);
nand I_939 (I17609,I17555,I17429);
not I_940 (I17627,I698);
DFFARX1 I_941 (I17366,I691,I17627,I17654,);
not I_942 (I17663,I17654);
DFFARX1 I_943 (I17609,I691,I17627,I17690,);
not I_944 (I17699,I17366);
nand I_945 (I17717,I17699,I17159);
not I_946 (I17735,I17717);
nor I_947 (I17753,I17735,I17384);
nor I_948 (I17771,I17663,I17753);
DFFARX1 I_949 (I17771,I691,I17627,I17798,);
not I_950 (I17807,I17384);
nand I_951 (I17825,I17807,I17735);
and I_952 (I17843,I17807,I17195);
nand I_953 (I17861,I17843,I17159);
nor I_954 (I17879,I17861,I17807);
and I_955 (I17897,I17690,I17861);
not I_956 (I17915,I17861);
nand I_957 (I17933,I17690,I17915);
nor I_958 (I17951,I17654,I17861);
not I_959 (I17969,I17591);
nor I_960 (I17987,I17969,I17195);
nand I_961 (I18005,I17987,I17807);
nor I_962 (I18023,I17717,I18005);
nor I_963 (I18041,I17969,I17078);
and I_964 (I18059,I18041,I17411);
or I_965 (I18077,I18059,I17501);
DFFARX1 I_966 (I18077,I691,I17627,I18104,);
nor I_967 (I18113,I18104,I17825);
DFFARX1 I_968 (I18113,I691,I17627,I18140,);
DFFARX1 I_969 (I18104,I691,I17627,I18158,);
not I_970 (I18167,I18104);
nor I_971 (I18185,I18167,I17690);
nor I_972 (I18203,I17987,I18185);
DFFARX1 I_973 (I18203,I691,I17627,I18230,);
not I_974 (I18239,I698);
DFFARX1 I_975 (I17951,I691,I18239,I18266,);
DFFARX1 I_976 (I18266,I691,I18239,I18284,);
not I_977 (I18293,I18284);
DFFARX1 I_978 (I17879,I691,I18239,I18320,);
not I_979 (I18329,I18140);
nor I_980 (I18347,I18266,I18329);
not I_981 (I18365,I17798);
not I_982 (I18383,I17933);
nand I_983 (I18401,I18383,I17798);
nor I_984 (I18419,I18329,I18401);
nor I_985 (I18437,I18320,I18419);
DFFARX1 I_986 (I18383,I691,I18239,I18464,);
nor I_987 (I18473,I17933,I18230);
nand I_988 (I18491,I18473,I18158);
nor I_989 (I18509,I18491,I18365);
nand I_990 (I18527,I18509,I18140);
DFFARX1 I_991 (I18491,I691,I18239,I18554,);
nand I_992 (I18563,I18365,I17933);
nor I_993 (I18581,I18365,I17933);
nand I_994 (I18599,I18347,I18581);
not I_995 (I18617,I18140);
nor I_996 (I18635,I18617,I18563);
DFFARX1 I_997 (I18635,I691,I18239,I18662,);
nor I_998 (I18671,I18617,I18023);
and I_999 (I18689,I18671,I17897);
or I_1000 (I18707,I18689,I17951);
DFFARX1 I_1001 (I18707,I691,I18239,I18734,);
nor I_1002 (I18743,I18734,I18320);
nor I_1003 (I18761,I18266,I18743);
not I_1004 (I18779,I18734);
nor I_1005 (I18797,I18779,I18437);
DFFARX1 I_1006 (I18797,I691,I18239,I18824,);
nand I_1007 (I18833,I18779,I18365);
nor I_1008 (I18851,I18617,I18833);
not I_1009 (I18869,I698);
DFFARX1 I_1010 (I18662,I691,I18869,I18896,);
not I_1011 (I18905,I18896);
nand I_1012 (I18923,I18824,I18662);
and I_1013 (I18941,I18923,I18851);
DFFARX1 I_1014 (I18941,I691,I18869,I18968,);
not I_1015 (I18977,I18851);
DFFARX1 I_1016 (I18599,I691,I18869,I19004,);
not I_1017 (I19013,I19004);
nor I_1018 (I19031,I19013,I18905);
and I_1019 (I19049,I19031,I18851);
nor I_1020 (I19067,I19013,I18977);
nor I_1021 (I19085,I18968,I19067);
DFFARX1 I_1022 (I18527,I691,I18869,I19112,);
nor I_1023 (I19121,I19112,I18968);
not I_1024 (I19139,I19121);
not I_1025 (I19157,I19112);
nor I_1026 (I19175,I19157,I19049);
DFFARX1 I_1027 (I19175,I691,I18869,I19202,);
nand I_1028 (I19211,I18761,I18554);
and I_1029 (I19229,I19211,I18293);
DFFARX1 I_1030 (I19229,I691,I18869,I19256,);
nor I_1031 (I19265,I19256,I19112);
DFFARX1 I_1032 (I19265,I691,I18869,I19292,);
nand I_1033 (I19301,I19256,I19157);
nand I_1034 (I19319,I19139,I19301);
not I_1035 (I19337,I19256);
nor I_1036 (I19355,I19337,I19049);
DFFARX1 I_1037 (I19355,I691,I18869,I19382,);
nor I_1038 (I19391,I18464,I18554);
or I_1039 (I19409,I19112,I19391);
nor I_1040 (I19427,I19256,I19391);
or I_1041 (I19445,I18968,I19391);
DFFARX1 I_1042 (I19391,I691,I18869,I19472,);
not I_1043 (I19481,I698);
DFFARX1 I_1044 (I19427,I691,I19481,I19508,);
nand I_1045 (I19517,I19508,I19202);
DFFARX1 I_1046 (I19409,I691,I19481,I19544,);
DFFARX1 I_1047 (I19544,I691,I19481,I19562,);
not I_1048 (I19571,I19562);
not I_1049 (I19589,I19085);
nor I_1050 (I19607,I19085,I19382);
not I_1051 (I19625,I19427);
nand I_1052 (I19643,I19589,I19625);
nor I_1053 (I19661,I19427,I19085);
and I_1054 (I19679,I19661,I19517);
not I_1055 (I19697,I19292);
nand I_1056 (I19715,I19697,I19445);
nor I_1057 (I19733,I19292,I19292);
not I_1058 (I19751,I19733);
nand I_1059 (I19769,I19607,I19751);
DFFARX1 I_1060 (I19733,I691,I19481,I19796,);
nor I_1061 (I19805,I19319,I19427);
nor I_1062 (I19823,I19805,I19382);
and I_1063 (I19841,I19823,I19715);
DFFARX1 I_1064 (I19841,I691,I19481,I19868,);
nor I_1065 (I19877,I19805,I19643);
or I_1066 (I19895,I19733,I19805);
nor I_1067 (I19913,I19319,I19472);
DFFARX1 I_1068 (I19913,I691,I19481,I19940,);
not I_1069 (I19949,I19940);
nand I_1070 (I19967,I19949,I19589);
nor I_1071 (I19985,I19967,I19382);
DFFARX1 I_1072 (I19985,I691,I19481,I20012,);
nor I_1073 (I20021,I19949,I19643);
nor I_1074 (I20039,I19805,I20021);
not I_1075 (I20057,I698);
DFFARX1 I_1076 (I19796,I691,I20057,I20084,);
and I_1077 (I20093,I20084,I19877);
DFFARX1 I_1078 (I20093,I691,I20057,I20120,);
DFFARX1 I_1079 (I20012,I691,I20057,I20138,);
not I_1080 (I20147,I19769);
not I_1081 (I20165,I19868);
nand I_1082 (I20183,I20165,I20147);
nor I_1083 (I20201,I20138,I20183);
DFFARX1 I_1084 (I20183,I691,I20057,I20228,);
not I_1085 (I20237,I20228);
not I_1086 (I20255,I20012);
nand I_1087 (I20273,I20165,I20255);
DFFARX1 I_1088 (I20273,I691,I20057,I20300,);
not I_1089 (I20309,I20300);
not I_1090 (I20327,I19571);
nand I_1091 (I20345,I20327,I19895);
and I_1092 (I20363,I20147,I20345);
nor I_1093 (I20381,I20273,I20363);
DFFARX1 I_1094 (I20381,I691,I20057,I20408,);
DFFARX1 I_1095 (I20363,I691,I20057,I20426,);
nor I_1096 (I20435,I19571,I19679);
nor I_1097 (I20453,I20273,I20435);
or I_1098 (I20471,I19571,I19679);
nor I_1099 (I20489,I20039,I19679);
DFFARX1 I_1100 (I20489,I691,I20057,I20516,);
not I_1101 (I20525,I20516);
nor I_1102 (I20543,I20525,I20309);
nand I_1103 (I20561,I20525,I20138);
not I_1104 (I20579,I20039);
nand I_1105 (I20597,I20579,I20255);
nand I_1106 (I20615,I20525,I20597);
nand I_1107 (I20633,I20615,I20561);
nand I_1108 (I20651,I20597,I20471);
not I_1109 (I20669,I698);
DFFARX1 I_1110 (I20543,I691,I20669,I20696,);
not I_1111 (I20705,I20696);
nand I_1112 (I20723,I20408,I20453);
and I_1113 (I20741,I20723,I20120);
DFFARX1 I_1114 (I20741,I691,I20669,I20768,);
not I_1115 (I20777,I20633);
DFFARX1 I_1116 (I20651,I691,I20669,I20804,);
not I_1117 (I20813,I20804);
nor I_1118 (I20831,I20813,I20705);
and I_1119 (I20849,I20831,I20633);
nor I_1120 (I20867,I20813,I20777);
nor I_1121 (I20885,I20768,I20867);
DFFARX1 I_1122 (I20237,I691,I20669,I20912,);
nor I_1123 (I20921,I20912,I20768);
not I_1124 (I20939,I20921);
not I_1125 (I20957,I20912);
nor I_1126 (I20975,I20957,I20849);
DFFARX1 I_1127 (I20975,I691,I20669,I21002,);
nand I_1128 (I21011,I20201,I20201);
and I_1129 (I21029,I21011,I20408);
DFFARX1 I_1130 (I21029,I691,I20669,I21056,);
nor I_1131 (I21065,I21056,I20912);
DFFARX1 I_1132 (I21065,I691,I20669,I21092,);
nand I_1133 (I21101,I21056,I20957);
nand I_1134 (I21119,I20939,I21101);
not I_1135 (I21137,I21056);
nor I_1136 (I21155,I21137,I20849);
DFFARX1 I_1137 (I21155,I691,I20669,I21182,);
nor I_1138 (I21191,I20426,I20201);
or I_1139 (I21209,I20912,I21191);
nor I_1140 (I21227,I21056,I21191);
or I_1141 (I21245,I20768,I21191);
DFFARX1 I_1142 (I21191,I691,I20669,I21272,);
not I_1143 (I21281,I698);
DFFARX1 I_1144 (I21227,I691,I21281,I21308,);
DFFARX1 I_1145 (I21308,I691,I21281,I21326,);
not I_1146 (I21335,I21326);
not I_1147 (I21353,I21308);
DFFARX1 I_1148 (I20885,I691,I21281,I21380,);
nand I_1149 (I21389,I21380,I21272);
not I_1150 (I21407,I21272);
not I_1151 (I21425,I21245);
nand I_1152 (I21443,I21119,I21092);
and I_1153 (I21461,I21119,I21092);
not I_1154 (I21479,I21002);
nand I_1155 (I21497,I21479,I21425);
nor I_1156 (I21515,I21497,I21389);
nor I_1157 (I21533,I21407,I21497);
nand I_1158 (I21551,I21461,I21533);
not I_1159 (I21569,I21182);
nor I_1160 (I21587,I21569,I21119);
nor I_1161 (I21605,I21587,I21002);
nor I_1162 (I21623,I21353,I21605);
DFFARX1 I_1163 (I21623,I691,I21281,I21650,);
not I_1164 (I21659,I21587);
DFFARX1 I_1165 (I21659,I691,I21281,I21686,);
and I_1166 (I21695,I21380,I21587);
nor I_1167 (I21713,I21569,I21092);
and I_1168 (I21731,I21713,I21209);
or I_1169 (I21749,I21731,I21227);
DFFARX1 I_1170 (I21749,I691,I21281,I21776,);
nor I_1171 (I21785,I21776,I21479);
DFFARX1 I_1172 (I21785,I691,I21281,I21812,);
nand I_1173 (I21821,I21776,I21380);
nand I_1174 (I21839,I21479,I21821);
nor I_1175 (I21857,I21839,I21443);
not I_1176 (I21875,I698);
DFFARX1 I_1177 (I21551,I691,I21875,I21902,);
not I_1178 (I21911,I21902);
nand I_1179 (I21929,I21515,I21335);
and I_1180 (I21947,I21929,I21686);
DFFARX1 I_1181 (I21947,I691,I21875,I21974,);
not I_1182 (I21983,I21812);
DFFARX1 I_1183 (I21515,I691,I21875,I22010,);
not I_1184 (I22019,I22010);
nor I_1185 (I22037,I22019,I21911);
and I_1186 (I22055,I22037,I21812);
nor I_1187 (I22073,I22019,I21983);
nor I_1188 (I22091,I21974,I22073);
DFFARX1 I_1189 (I21695,I691,I21875,I22118,);
nor I_1190 (I22127,I22118,I21974);
not I_1191 (I22145,I22127);
not I_1192 (I22163,I22118);
nor I_1193 (I22181,I22163,I22055);
DFFARX1 I_1194 (I22181,I691,I21875,I22208,);
nand I_1195 (I22217,I21650,I21812);
and I_1196 (I22235,I22217,I21551);
DFFARX1 I_1197 (I22235,I691,I21875,I22262,);
nor I_1198 (I22271,I22262,I22118);
DFFARX1 I_1199 (I22271,I691,I21875,I22298,);
nand I_1200 (I22307,I22262,I22163);
nand I_1201 (I22325,I22145,I22307);
not I_1202 (I22343,I22262);
nor I_1203 (I22361,I22343,I22055);
DFFARX1 I_1204 (I22361,I691,I21875,I22388,);
nor I_1205 (I22397,I21857,I21812);
or I_1206 (I22415,I22118,I22397);
nor I_1207 (I22433,I22262,I22397);
or I_1208 (I22451,I21974,I22397);
DFFARX1 I_1209 (I22397,I691,I21875,I22478,);
not I_1210 (I22487,I698);
DFFARX1 I_1211 (I22325,I691,I22487,I22514,);
DFFARX1 I_1212 (I22514,I691,I22487,I22532,);
not I_1213 (I22541,I22532);
DFFARX1 I_1214 (I22433,I691,I22487,I22568,);
not I_1215 (I22577,I22298);
nor I_1216 (I22595,I22514,I22577);
not I_1217 (I22613,I22415);
not I_1218 (I22631,I22091);
nand I_1219 (I22649,I22631,I22415);
nor I_1220 (I22667,I22577,I22649);
nor I_1221 (I22685,I22568,I22667);
DFFARX1 I_1222 (I22631,I691,I22487,I22712,);
nor I_1223 (I22721,I22091,I22478);
nand I_1224 (I22739,I22721,I22208);
nor I_1225 (I22757,I22739,I22613);
nand I_1226 (I22775,I22757,I22298);
DFFARX1 I_1227 (I22739,I691,I22487,I22802,);
nand I_1228 (I22811,I22613,I22091);
nor I_1229 (I22829,I22613,I22091);
nand I_1230 (I22847,I22595,I22829);
not I_1231 (I22865,I22451);
nor I_1232 (I22883,I22865,I22811);
DFFARX1 I_1233 (I22883,I691,I22487,I22910,);
nor I_1234 (I22919,I22865,I22388);
and I_1235 (I22937,I22919,I22298);
or I_1236 (I22955,I22937,I22433);
DFFARX1 I_1237 (I22955,I691,I22487,I22982,);
nor I_1238 (I22991,I22982,I22568);
nor I_1239 (I23009,I22514,I22991);
not I_1240 (I23027,I22982);
nor I_1241 (I23045,I23027,I22685);
DFFARX1 I_1242 (I23045,I691,I22487,I23072,);
nand I_1243 (I23081,I23027,I22613);
nor I_1244 (I23099,I22865,I23081);
not I_1245 (I23117,I698);
DFFARX1 I_1246 (I23099,I691,I23117,I23144,);
DFFARX1 I_1247 (I23072,I691,I23117,I23162,);
not I_1248 (I23171,I23162);
not I_1249 (I23189,I22910);
nor I_1250 (I23207,I23189,I22802);
not I_1251 (I23225,I22541);
nor I_1252 (I23243,I23207,I22775);
nor I_1253 (I23261,I23162,I23243);
DFFARX1 I_1254 (I23261,I691,I23117,I23288,);
nor I_1255 (I23297,I22775,I22802);
nand I_1256 (I23315,I23297,I22910);
DFFARX1 I_1257 (I23315,I691,I23117,I23342,);
nor I_1258 (I23351,I23225,I22775);
nand I_1259 (I23369,I23351,I23009);
nor I_1260 (I23387,I23144,I23369);
DFFARX1 I_1261 (I23387,I691,I23117,I23414,);
not I_1262 (I23423,I23369);
nand I_1263 (I23441,I23162,I23423);
DFFARX1 I_1264 (I23369,I691,I23117,I23468,);
not I_1265 (I23477,I23468);
not I_1266 (I23495,I22775);
not I_1267 (I23513,I22847);
nor I_1268 (I23531,I23513,I22541);
nor I_1269 (I23549,I23477,I23531);
nor I_1270 (I23567,I23513,I22712);
and I_1271 (I23585,I23567,I22910);
or I_1272 (I23603,I23585,I23099);
DFFARX1 I_1273 (I23603,I691,I23117,I23630,);
nor I_1274 (I23639,I23630,I23144);
not I_1275 (I23657,I23630);
and I_1276 (I23675,I23657,I23144);
nor I_1277 (I23693,I23171,I23675);
nand I_1278 (I23711,I23657,I23225);
nor I_1279 (I23729,I23513,I23711);
nand I_1280 (I23747,I23657,I23423);
nand I_1281 (I23765,I23225,I22847);
nor I_1282 (I23783,I23495,I23765);
not I_1283 (I23801,I698);
DFFARX1 I_1284 (I23639,I691,I23801,I23828,);
DFFARX1 I_1285 (I23828,I691,I23801,I23846,);
not I_1286 (I23855,I23846);
DFFARX1 I_1287 (I23729,I691,I23801,I23882,);
not I_1288 (I23891,I23414);
nor I_1289 (I23909,I23828,I23891);
not I_1290 (I23927,I23441);
not I_1291 (I23945,I23693);
nand I_1292 (I23963,I23945,I23441);
nor I_1293 (I23981,I23891,I23963);
nor I_1294 (I23999,I23882,I23981);
DFFARX1 I_1295 (I23945,I691,I23801,I24026,);
nor I_1296 (I24035,I23693,I23783);
nand I_1297 (I24053,I24035,I23288);
nor I_1298 (I24071,I24053,I23927);
nand I_1299 (I24089,I24071,I23414);
DFFARX1 I_1300 (I24053,I691,I23801,I24116,);
nand I_1301 (I24125,I23927,I23693);
nor I_1302 (I24143,I23927,I23693);
nand I_1303 (I24161,I23909,I24143);
not I_1304 (I24179,I23342);
nor I_1305 (I24197,I24179,I24125);
DFFARX1 I_1306 (I24197,I691,I23801,I24224,);
nor I_1307 (I24233,I24179,I23549);
and I_1308 (I24251,I24233,I23747);
or I_1309 (I24269,I24251,I23414);
DFFARX1 I_1310 (I24269,I691,I23801,I24296,);
nor I_1311 (I24305,I24296,I23882);
nor I_1312 (I24323,I23828,I24305);
not I_1313 (I24341,I24296);
nor I_1314 (I24359,I24341,I23999);
DFFARX1 I_1315 (I24359,I691,I23801,I24386,);
nand I_1316 (I24395,I24341,I23927);
nor I_1317 (I24413,I24179,I24395);
not I_1318 (I24431,I698);
DFFARX1 I_1319 (I380,I691,I24431,I24458,);
DFFARX1 I_1320 (I24458,I691,I24431,I24476,);
not I_1321 (I24485,I24476);
not I_1322 (I24503,I24458);
DFFARX1 I_1323 (I436,I691,I24431,I24530,);
nand I_1324 (I24539,I24530,I572);
not I_1325 (I24557,I572);
not I_1326 (I24575,I684);
nand I_1327 (I24593,I476,I100);
and I_1328 (I24611,I476,I100);
not I_1329 (I24629,I276);
nand I_1330 (I24647,I24629,I24575);
nor I_1331 (I24665,I24647,I24539);
nor I_1332 (I24683,I24557,I24647);
nand I_1333 (I24701,I24611,I24683);
not I_1334 (I24719,I588);
nor I_1335 (I24737,I24719,I476);
nor I_1336 (I24755,I24737,I276);
nor I_1337 (I24773,I24503,I24755);
DFFARX1 I_1338 (I24773,I691,I24431,I24800,);
not I_1339 (I24809,I24737);
DFFARX1 I_1340 (I24809,I691,I24431,I24836,);
and I_1341 (I24845,I24530,I24737);
nor I_1342 (I24863,I24719,I228);
and I_1343 (I24881,I24863,I444);
or I_1344 (I24899,I24881,I300);
DFFARX1 I_1345 (I24899,I691,I24431,I24926,);
nor I_1346 (I24935,I24926,I24629);
DFFARX1 I_1347 (I24935,I691,I24431,I24962,);
nand I_1348 (I24971,I24926,I24530);
nand I_1349 (I24989,I24629,I24971);
nor I_1350 (I25007,I24989,I24593);
not I_1351 (I25025,I698);
DFFARX1 I_1352 (I25007,I691,I25025,I25052,);
nand I_1353 (I25061,I25052,I24701);
not I_1354 (I25079,I25061);
DFFARX1 I_1355 (I24701,I691,I25025,I25106,);
not I_1356 (I25115,I25106);
not I_1357 (I25133,I24665);
or I_1358 (I25151,I24845,I24665);
nor I_1359 (I25169,I24845,I24665);
or I_1360 (I25187,I24800,I24845);
DFFARX1 I_1361 (I25187,I691,I25025,I25214,);
not I_1362 (I25223,I24665);
nand I_1363 (I25241,I25223,I24962);
nand I_1364 (I25259,I25133,I25241);
and I_1365 (I25277,I25115,I25259);
nor I_1366 (I25295,I24665,I24836);
and I_1367 (I25313,I25115,I25295);
nor I_1368 (I25331,I25079,I25313);
DFFARX1 I_1369 (I25295,I691,I25025,I25358,);
not I_1370 (I25367,I25358);
nor I_1371 (I25385,I25115,I25367);
or I_1372 (I25403,I25187,I24485);
nor I_1373 (I25421,I24485,I24800);
nand I_1374 (I25439,I25259,I25421);
nand I_1375 (I25457,I25403,I25439);
DFFARX1 I_1376 (I25457,I691,I25025,I25484,);
nor I_1377 (I25493,I25421,I25151);
DFFARX1 I_1378 (I25493,I691,I25025,I25520,);
nor I_1379 (I25529,I24485,I24962);
DFFARX1 I_1380 (I25529,I691,I25025,I25556,);
DFFARX1 I_1381 (I25556,I691,I25025,I25574,);
not I_1382 (I25583,I25556);
nand I_1383 (I25601,I25583,I25061);
nand I_1384 (I25619,I25583,I25169);
not I_1385 (I25637,I698);
DFFARX1 I_1386 (I25385,I691,I25637,I25664,);
not I_1387 (I25673,I25664);
nand I_1388 (I25691,I25520,I25277);
and I_1389 (I25709,I25691,I25574);
DFFARX1 I_1390 (I25709,I691,I25637,I25736,);
DFFARX1 I_1391 (I25736,I691,I25637,I25754,);
DFFARX1 I_1392 (I25214,I691,I25637,I25772,);
nand I_1393 (I25781,I25772,I25331);
not I_1394 (I25799,I25781);
DFFARX1 I_1395 (I25799,I691,I25637,I25826,);
not I_1396 (I25835,I25826);
nor I_1397 (I25853,I25673,I25835);
DFFARX1 I_1398 (I25484,I691,I25637,I25880,);
nor I_1399 (I25889,I25880,I25736);
nor I_1400 (I25907,I25880,I25799);
nand I_1401 (I25925,I25601,I25619);
and I_1402 (I25943,I25925,I25520);
DFFARX1 I_1403 (I25943,I691,I25637,I25970,);
not I_1404 (I25979,I25970);
nand I_1405 (I25997,I25979,I25880);
nand I_1406 (I26015,I25979,I25781);
nor I_1407 (I26033,I25277,I25619);
and I_1408 (I26051,I25880,I26033);
nor I_1409 (I26069,I25979,I26051);
DFFARX1 I_1410 (I26069,I691,I25637,I26096,);
nor I_1411 (I26105,I25664,I26033);
DFFARX1 I_1412 (I26105,I691,I25637,I26132,);
nor I_1413 (I26141,I25970,I26033);
not I_1414 (I26159,I26141);
nand I_1415 (I26177,I26159,I25997);
not I_1416 (I26195,I698);
DFFARX1 I_1417 (I26177,I691,I26195,I26222,);
DFFARX1 I_1418 (I26015,I691,I26195,I26240,);
not I_1419 (I26249,I26240);
nor I_1420 (I26267,I26222,I26249);
DFFARX1 I_1421 (I26249,I691,I26195,I26294,);
nor I_1422 (I26303,I25853,I25907);
and I_1423 (I26321,I26303,I26132);
nor I_1424 (I26339,I26321,I25853);
not I_1425 (I26357,I25853);
and I_1426 (I26375,I26357,I26015);
nand I_1427 (I26393,I26375,I25754);
nor I_1428 (I26411,I26357,I26393);
DFFARX1 I_1429 (I26411,I691,I26195,I26438,);
not I_1430 (I26447,I26393);
nand I_1431 (I26465,I26249,I26447);
nand I_1432 (I26483,I26321,I26447);
DFFARX1 I_1433 (I26357,I691,I26195,I26510,);
not I_1434 (I26519,I25889);
nor I_1435 (I26537,I26519,I26015);
nor I_1436 (I26555,I26537,I26339);
DFFARX1 I_1437 (I26555,I691,I26195,I26582,);
not I_1438 (I26591,I26537);
DFFARX1 I_1439 (I26591,I691,I26195,I26618,);
not I_1440 (I26627,I26618);
nor I_1441 (I26645,I26627,I26537);
nor I_1442 (I26663,I26519,I26132);
and I_1443 (I26681,I26663,I26096);
or I_1444 (I26699,I26681,I25907);
DFFARX1 I_1445 (I26699,I691,I26195,I26726,);
not I_1446 (I26735,I26726);
nand I_1447 (I26753,I26735,I26447);
not I_1448 (I26771,I26753);
nand I_1449 (I26789,I26753,I26465);
nand I_1450 (I26807,I26735,I26321);
not I_1451 (I26825,I698);
DFFARX1 I_1452 (I26645,I691,I26825,I26852,);
DFFARX1 I_1453 (I26852,I691,I26825,I26870,);
not I_1454 (I26879,I26870);
not I_1455 (I26897,I26852);
DFFARX1 I_1456 (I26483,I691,I26825,I26924,);
not I_1457 (I26933,I26924);
and I_1458 (I26951,I26897,I26807);
not I_1459 (I26969,I26438);
nand I_1460 (I26987,I26969,I26807);
not I_1461 (I27005,I26510);
nor I_1462 (I27023,I27005,I26438);
nand I_1463 (I27041,I27023,I26582);
nor I_1464 (I27059,I27041,I26987);
DFFARX1 I_1465 (I27059,I691,I26825,I27086,);
not I_1466 (I27095,I27041);
not I_1467 (I27113,I26438);
nand I_1468 (I27131,I27113,I26807);
nor I_1469 (I27149,I26438,I26438);
nand I_1470 (I27167,I26951,I27149);
nand I_1471 (I27185,I26897,I26438);
nand I_1472 (I27203,I27005,I26789);
DFFARX1 I_1473 (I27203,I691,I26825,I27230,);
DFFARX1 I_1474 (I27203,I691,I26825,I27248,);
not I_1475 (I27257,I26789);
nor I_1476 (I27275,I27257,I26771);
and I_1477 (I27293,I27275,I26294);
or I_1478 (I27311,I27293,I26267);
DFFARX1 I_1479 (I27311,I691,I26825,I27338,);
nand I_1480 (I27347,I27338,I26969);
nor I_1481 (I27365,I27347,I27131);
nor I_1482 (I27383,I27338,I26933);
DFFARX1 I_1483 (I27338,I691,I26825,I27410,);
not I_1484 (I27419,I27410);
nor I_1485 (I27437,I27419,I27095);
not I_1486 (I27455,I698);
DFFARX1 I_1487 (I27086,I691,I27455,I27482,);
not I_1488 (I27491,I27482);
nand I_1489 (I27509,I27383,I26879);
and I_1490 (I27527,I27509,I27167);
DFFARX1 I_1491 (I27527,I691,I27455,I27554,);
not I_1492 (I27563,I27365);
DFFARX1 I_1493 (I27086,I691,I27455,I27590,);
not I_1494 (I27599,I27590);
nor I_1495 (I27617,I27599,I27491);
and I_1496 (I27635,I27617,I27365);
nor I_1497 (I27653,I27599,I27563);
nor I_1498 (I27671,I27554,I27653);
DFFARX1 I_1499 (I27437,I691,I27455,I27698,);
nor I_1500 (I27707,I27698,I27554);
not I_1501 (I27725,I27707);
not I_1502 (I27743,I27698);
nor I_1503 (I27761,I27743,I27635);
DFFARX1 I_1504 (I27761,I691,I27455,I27788,);
nand I_1505 (I27797,I27383,I27185);
and I_1506 (I27815,I27797,I27248);
DFFARX1 I_1507 (I27815,I691,I27455,I27842,);
nor I_1508 (I27851,I27842,I27698);
DFFARX1 I_1509 (I27851,I691,I27455,I27878,);
nand I_1510 (I27887,I27842,I27743);
nand I_1511 (I27905,I27725,I27887);
not I_1512 (I27923,I27842);
nor I_1513 (I27941,I27923,I27635);
DFFARX1 I_1514 (I27941,I691,I27455,I27968,);
nor I_1515 (I27977,I27230,I27185);
or I_1516 (I27995,I27698,I27977);
nor I_1517 (I28013,I27842,I27977);
or I_1518 (I28031,I27554,I27977);
DFFARX1 I_1519 (I27977,I691,I27455,I28058,);
not I_1520 (I28067,I698);
DFFARX1 I_1521 (I28031,I691,I28067,I28094,);
DFFARX1 I_1522 (I28094,I691,I28067,I28112,);
not I_1523 (I28121,I28112);
nand I_1524 (I28139,I27968,I28058);
and I_1525 (I28157,I28139,I28013);
DFFARX1 I_1526 (I28157,I691,I28067,I28184,);
DFFARX1 I_1527 (I28184,I691,I28067,I28202,);
DFFARX1 I_1528 (I28184,I691,I28067,I28220,);
DFFARX1 I_1529 (I27905,I691,I28067,I28238,);
nand I_1530 (I28247,I28238,I27671);
not I_1531 (I28265,I28247);
nor I_1532 (I28283,I28094,I28265);
DFFARX1 I_1533 (I28013,I691,I28067,I28310,);
not I_1534 (I28319,I28310);
nor I_1535 (I28337,I28319,I28121);
nand I_1536 (I28355,I28319,I28247);
nand I_1537 (I28373,I27788,I27878);
and I_1538 (I28391,I28373,I27995);
DFFARX1 I_1539 (I28391,I691,I28067,I28418,);
nor I_1540 (I28427,I28418,I28094);
DFFARX1 I_1541 (I28427,I691,I28067,I28454,);
not I_1542 (I28463,I28418);
nor I_1543 (I28481,I27878,I27878);
not I_1544 (I28499,I28481);
nor I_1545 (I28517,I28247,I28499);
nor I_1546 (I28535,I28463,I28517);
DFFARX1 I_1547 (I28535,I691,I28067,I28562,);
nor I_1548 (I28571,I28418,I28499);
nor I_1549 (I28589,I28265,I28571);
nor I_1550 (I28607,I28418,I28481);
not I_1551 (I28625,I698);
DFFARX1 I_1552 (I28454,I691,I28625,I28652,);
DFFARX1 I_1553 (I28652,I691,I28625,I28670,);
not I_1554 (I28679,I28670);
DFFARX1 I_1555 (I28454,I691,I28625,I28706,);
not I_1556 (I28715,I28202);
nor I_1557 (I28733,I28652,I28715);
not I_1558 (I28751,I28337);
not I_1559 (I28769,I28589);
nand I_1560 (I28787,I28769,I28337);
nor I_1561 (I28805,I28715,I28787);
nor I_1562 (I28823,I28706,I28805);
DFFARX1 I_1563 (I28769,I691,I28625,I28850,);
nor I_1564 (I28859,I28589,I28562);
nand I_1565 (I28877,I28859,I28607);
nor I_1566 (I28895,I28877,I28751);
nand I_1567 (I28913,I28895,I28202);
DFFARX1 I_1568 (I28877,I691,I28625,I28940,);
nand I_1569 (I28949,I28751,I28589);
nor I_1570 (I28967,I28751,I28589);
nand I_1571 (I28985,I28733,I28967);
not I_1572 (I29003,I28607);
nor I_1573 (I29021,I29003,I28949);
DFFARX1 I_1574 (I29021,I691,I28625,I29048,);
nor I_1575 (I29057,I29003,I28283);
and I_1576 (I29075,I29057,I28355);
or I_1577 (I29093,I29075,I28220);
DFFARX1 I_1578 (I29093,I691,I28625,I29120,);
nor I_1579 (I29129,I29120,I28706);
nor I_1580 (I29147,I28652,I29129);
not I_1581 (I29165,I29120);
nor I_1582 (I29183,I29165,I28823);
DFFARX1 I_1583 (I29183,I691,I28625,I29210,);
nand I_1584 (I29219,I29165,I28751);
nor I_1585 (I29237,I29003,I29219);
not I_1586 (I29255,I698);
DFFARX1 I_1587 (I29237,I691,I29255,I29282,);
not I_1588 (I29291,I29282);
DFFARX1 I_1589 (I29210,I691,I29255,I29318,);
not I_1590 (I29327,I28850);
nand I_1591 (I29345,I29327,I28985);
not I_1592 (I29363,I29345);
nor I_1593 (I29381,I29363,I28940);
nor I_1594 (I29399,I29291,I29381);
DFFARX1 I_1595 (I29399,I691,I29255,I29426,);
not I_1596 (I29435,I28940);
nand I_1597 (I29453,I29435,I29363);
and I_1598 (I29471,I29435,I29147);
nand I_1599 (I29489,I29471,I29048);
nor I_1600 (I29507,I29489,I29435);
and I_1601 (I29525,I29318,I29489);
not I_1602 (I29543,I29489);
nand I_1603 (I29561,I29318,I29543);
nor I_1604 (I29579,I29282,I29489);
not I_1605 (I29597,I28913);
nor I_1606 (I29615,I29597,I29147);
nand I_1607 (I29633,I29615,I29435);
nor I_1608 (I29651,I29345,I29633);
nor I_1609 (I29669,I29597,I29237);
and I_1610 (I29687,I29669,I29048);
or I_1611 (I29705,I29687,I28679);
DFFARX1 I_1612 (I29705,I691,I29255,I29732,);
nor I_1613 (I29741,I29732,I29453);
DFFARX1 I_1614 (I29741,I691,I29255,I29768,);
DFFARX1 I_1615 (I29732,I691,I29255,I29786,);
not I_1616 (I29795,I29732);
nor I_1617 (I29813,I29795,I29318);
nor I_1618 (I29831,I29615,I29813);
DFFARX1 I_1619 (I29831,I691,I29255,I29858,);
not I_1620 (I29867,I698);
DFFARX1 I_1621 (I29858,I691,I29867,I29894,);
DFFARX1 I_1622 (I29507,I691,I29867,I29912,);
not I_1623 (I29921,I29912);
nor I_1624 (I29939,I29894,I29921);
DFFARX1 I_1625 (I29921,I691,I29867,I29966,);
nor I_1626 (I29975,I29651,I29579);
and I_1627 (I29993,I29975,I29768);
nor I_1628 (I30011,I29993,I29651);
not I_1629 (I30029,I29651);
and I_1630 (I30047,I30029,I29525);
nand I_1631 (I30065,I30047,I29426);
nor I_1632 (I30083,I30029,I30065);
DFFARX1 I_1633 (I30083,I691,I29867,I30110,);
not I_1634 (I30119,I30065);
nand I_1635 (I30137,I29921,I30119);
nand I_1636 (I30155,I29993,I30119);
DFFARX1 I_1637 (I30029,I691,I29867,I30182,);
not I_1638 (I30191,I29786);
nor I_1639 (I30209,I30191,I29525);
nor I_1640 (I30227,I30209,I30011);
DFFARX1 I_1641 (I30227,I691,I29867,I30254,);
not I_1642 (I30263,I30209);
DFFARX1 I_1643 (I30263,I691,I29867,I30290,);
not I_1644 (I30299,I30290);
nor I_1645 (I30317,I30299,I30209);
nor I_1646 (I30335,I30191,I29579);
and I_1647 (I30353,I30335,I29561);
or I_1648 (I30371,I30353,I29768);
DFFARX1 I_1649 (I30371,I691,I29867,I30398,);
not I_1650 (I30407,I30398);
nand I_1651 (I30425,I30407,I30119);
not I_1652 (I30443,I30425);
nand I_1653 (I30461,I30425,I30137);
nand I_1654 (I30479,I30407,I29993);
not I_1655 (I30497,I698);
DFFARX1 I_1656 (I30182,I691,I30497,I30524,);
not I_1657 (I30533,I30524);
nand I_1658 (I30551,I30155,I30110);
and I_1659 (I30569,I30551,I30443);
DFFARX1 I_1660 (I30569,I691,I30497,I30596,);
not I_1661 (I30605,I30110);
DFFARX1 I_1662 (I29966,I691,I30497,I30632,);
not I_1663 (I30641,I30632);
nor I_1664 (I30659,I30641,I30533);
and I_1665 (I30677,I30659,I30110);
nor I_1666 (I30695,I30641,I30605);
nor I_1667 (I30713,I30596,I30695);
DFFARX1 I_1668 (I30479,I691,I30497,I30740,);
nor I_1669 (I30749,I30740,I30596);
not I_1670 (I30767,I30749);
not I_1671 (I30785,I30740);
nor I_1672 (I30803,I30785,I30677);
DFFARX1 I_1673 (I30803,I691,I30497,I30830,);
nand I_1674 (I30839,I29939,I30461);
and I_1675 (I30857,I30839,I30254);
DFFARX1 I_1676 (I30857,I691,I30497,I30884,);
nor I_1677 (I30893,I30884,I30740);
DFFARX1 I_1678 (I30893,I691,I30497,I30920,);
nand I_1679 (I30929,I30884,I30785);
nand I_1680 (I30947,I30767,I30929);
not I_1681 (I30965,I30884);
nor I_1682 (I30983,I30965,I30677);
DFFARX1 I_1683 (I30983,I691,I30497,I31010,);
nor I_1684 (I31019,I30317,I30461);
or I_1685 (I31037,I30740,I31019);
nor I_1686 (I31055,I30884,I31019);
or I_1687 (I31073,I30596,I31019);
DFFARX1 I_1688 (I31019,I691,I30497,I31100,);
not I_1689 (I31109,I698);
DFFARX1 I_1690 (I31010,I691,I31109,I31136,);
DFFARX1 I_1691 (I31055,I691,I31109,I31154,);
not I_1692 (I31163,I31154);
nor I_1693 (I31181,I31136,I31163);
DFFARX1 I_1694 (I31163,I691,I31109,I31208,);
nor I_1695 (I31217,I30947,I31037);
and I_1696 (I31235,I31217,I30920);
nor I_1697 (I31253,I31235,I30947);
not I_1698 (I31271,I30947);
and I_1699 (I31289,I31271,I30830);
nand I_1700 (I31307,I31289,I31073);
nor I_1701 (I31325,I31271,I31307);
DFFARX1 I_1702 (I31325,I691,I31109,I31352,);
not I_1703 (I31361,I31307);
nand I_1704 (I31379,I31163,I31361);
nand I_1705 (I31397,I31235,I31361);
DFFARX1 I_1706 (I31271,I691,I31109,I31424,);
not I_1707 (I31433,I31055);
nor I_1708 (I31451,I31433,I30830);
nor I_1709 (I31469,I31451,I31253);
DFFARX1 I_1710 (I31469,I691,I31109,I31496,);
not I_1711 (I31505,I31451);
DFFARX1 I_1712 (I31505,I691,I31109,I31532,);
not I_1713 (I31541,I31532);
nor I_1714 (I31559,I31541,I31451);
nor I_1715 (I31577,I31433,I30713);
and I_1716 (I31595,I31577,I31100);
or I_1717 (I31613,I31595,I30920);
DFFARX1 I_1718 (I31613,I691,I31109,I31640,);
not I_1719 (I31649,I31640);
nand I_1720 (I31667,I31649,I31361);
not I_1721 (I31685,I31667);
nand I_1722 (I31703,I31667,I31379);
nand I_1723 (I31721,I31649,I31235);
not I_1724 (I31739,I698);
DFFARX1 I_1725 (I31685,I691,I31739,I31766,);
not I_1726 (I31775,I31766);
nand I_1727 (I31793,I31397,I31559);
and I_1728 (I31811,I31793,I31352);
DFFARX1 I_1729 (I31811,I691,I31739,I31838,);
DFFARX1 I_1730 (I31838,I691,I31739,I31856,);
DFFARX1 I_1731 (I31181,I691,I31739,I31874,);
nand I_1732 (I31883,I31874,I31208);
not I_1733 (I31901,I31883);
DFFARX1 I_1734 (I31901,I691,I31739,I31928,);
not I_1735 (I31937,I31928);
nor I_1736 (I31955,I31775,I31937);
DFFARX1 I_1737 (I31496,I691,I31739,I31982,);
nor I_1738 (I31991,I31982,I31838);
nor I_1739 (I32009,I31982,I31901);
nand I_1740 (I32027,I31721,I31424);
and I_1741 (I32045,I32027,I31703);
DFFARX1 I_1742 (I32045,I691,I31739,I32072,);
not I_1743 (I32081,I32072);
nand I_1744 (I32099,I32081,I31982);
nand I_1745 (I32117,I32081,I31883);
nor I_1746 (I32135,I31352,I31424);
and I_1747 (I32153,I31982,I32135);
nor I_1748 (I32171,I32081,I32153);
DFFARX1 I_1749 (I32171,I691,I31739,I32198,);
nor I_1750 (I32207,I31766,I32135);
DFFARX1 I_1751 (I32207,I691,I31739,I32234,);
nor I_1752 (I32243,I32072,I32135);
not I_1753 (I32261,I32243);
nand I_1754 (I32279,I32261,I32099);
not I_1755 (I32297,I698);
DFFARX1 I_1756 (I32117,I691,I32297,I32324,);
DFFARX1 I_1757 (I32324,I691,I32297,I32342,);
not I_1758 (I32351,I32342);
not I_1759 (I32369,I32324);
DFFARX1 I_1760 (I32234,I691,I32297,I32396,);
not I_1761 (I32405,I32396);
and I_1762 (I32423,I32369,I31856);
not I_1763 (I32441,I32117);
nand I_1764 (I32459,I32441,I31856);
not I_1765 (I32477,I32234);
nor I_1766 (I32495,I32477,I31991);
nand I_1767 (I32513,I32495,I32009);
nor I_1768 (I32531,I32513,I32459);
DFFARX1 I_1769 (I32531,I691,I32297,I32558,);
not I_1770 (I32567,I32513);
not I_1771 (I32585,I31991);
nand I_1772 (I32603,I32585,I31856);
nor I_1773 (I32621,I31991,I32117);
nand I_1774 (I32639,I32423,I32621);
nand I_1775 (I32657,I32369,I31991);
nand I_1776 (I32675,I32477,I32198);
DFFARX1 I_1777 (I32675,I691,I32297,I32702,);
DFFARX1 I_1778 (I32675,I691,I32297,I32720,);
not I_1779 (I32729,I32198);
nor I_1780 (I32747,I32729,I31955);
and I_1781 (I32765,I32747,I32009);
or I_1782 (I32783,I32765,I32279);
DFFARX1 I_1783 (I32783,I691,I32297,I32810,);
nand I_1784 (I32819,I32810,I32441);
nor I_1785 (I32837,I32819,I32603);
nor I_1786 (I32855,I32810,I32405);
DFFARX1 I_1787 (I32810,I691,I32297,I32882,);
not I_1788 (I32891,I32882);
nor I_1789 (I32909,I32891,I32567);
not I_1790 (I32927,I698);
DFFARX1 I_1791 (I32639,I691,I32927,I32954,);
not I_1792 (I32963,I32954);
nand I_1793 (I32981,I32657,I32558);
and I_1794 (I32999,I32981,I32702);
DFFARX1 I_1795 (I32999,I691,I32927,I33026,);
DFFARX1 I_1796 (I32909,I691,I32927,I33044,);
and I_1797 (I33053,I33044,I32720);
nor I_1798 (I33071,I33026,I33053);
DFFARX1 I_1799 (I33071,I691,I32927,I33098,);
nand I_1800 (I33107,I33044,I32720);
nand I_1801 (I33125,I32963,I33107);
not I_1802 (I33143,I33125);
DFFARX1 I_1803 (I32558,I691,I32927,I33170,);
DFFARX1 I_1804 (I33170,I691,I32927,I33188,);
nand I_1805 (I33197,I32855,I32855);
and I_1806 (I33215,I33197,I32351);
DFFARX1 I_1807 (I33215,I691,I32927,I33242,);
DFFARX1 I_1808 (I33242,I691,I32927,I33260,);
not I_1809 (I33269,I33260);
not I_1810 (I33287,I33242);
nand I_1811 (I33305,I33287,I33107);
nor I_1812 (I33323,I32837,I32855);
not I_1813 (I33341,I33323);
nor I_1814 (I33359,I33287,I33341);
nor I_1815 (I33377,I32963,I33359);
DFFARX1 I_1816 (I33377,I691,I32927,I33404,);
nor I_1817 (I33413,I33026,I33341);
nor I_1818 (I33431,I33242,I33413);
nor I_1819 (I33449,I33170,I33323);
nor I_1820 (I33467,I33026,I33323);
not I_1821 (I33485,I698);
DFFARX1 I_1822 (I33467,I691,I33485,I33512,);
nand I_1823 (I33521,I33449,I33269);
and I_1824 (I33539,I33521,I33467);
DFFARX1 I_1825 (I33539,I691,I33485,I33566,);
nor I_1826 (I33575,I33566,I33512);
not I_1827 (I33593,I33566);
DFFARX1 I_1828 (I33404,I691,I33485,I33620,);
nand I_1829 (I33629,I33620,I33431);
not I_1830 (I33647,I33629);
DFFARX1 I_1831 (I33647,I691,I33485,I33674,);
not I_1832 (I33683,I33674);
nor I_1833 (I33701,I33512,I33629);
nor I_1834 (I33719,I33566,I33701);
DFFARX1 I_1835 (I33305,I691,I33485,I33746,);
DFFARX1 I_1836 (I33746,I691,I33485,I33764,);
not I_1837 (I33773,I33764);
not I_1838 (I33791,I33746);
nand I_1839 (I33809,I33791,I33593);
nand I_1840 (I33827,I33098,I33098);
and I_1841 (I33845,I33827,I33143);
DFFARX1 I_1842 (I33845,I691,I33485,I33872,);
nor I_1843 (I33881,I33872,I33512);
DFFARX1 I_1844 (I33881,I691,I33485,I33908,);
DFFARX1 I_1845 (I33872,I691,I33485,I33926,);
nor I_1846 (I33935,I33188,I33098);
not I_1847 (I33953,I33935);
nor I_1848 (I33971,I33773,I33953);
nand I_1849 (I33989,I33791,I33953);
nor I_1850 (I34007,I33512,I33935);
DFFARX1 I_1851 (I33935,I691,I33485,I34034,);
not I_1852 (I34043,I698);
DFFARX1 I_1853 (I33989,I691,I34043,I34070,);
nand I_1854 (I34079,I34070,I33683);
not I_1855 (I34097,I34079);
DFFARX1 I_1856 (I33971,I691,I34043,I34124,);
not I_1857 (I34133,I34124);
not I_1858 (I34151,I33719);
or I_1859 (I34169,I34034,I33719);
nor I_1860 (I34187,I34034,I33719);
or I_1861 (I34205,I34007,I34034);
DFFARX1 I_1862 (I34205,I691,I34043,I34232,);
not I_1863 (I34241,I33575);
nand I_1864 (I34259,I34241,I33908);
nand I_1865 (I34277,I34151,I34259);
and I_1866 (I34295,I34133,I34277);
nor I_1867 (I34313,I33575,I33809);
and I_1868 (I34331,I34133,I34313);
nor I_1869 (I34349,I34097,I34331);
DFFARX1 I_1870 (I34313,I691,I34043,I34376,);
not I_1871 (I34385,I34376);
nor I_1872 (I34403,I34133,I34385);
or I_1873 (I34421,I34205,I33926);
nor I_1874 (I34439,I33926,I34007);
nand I_1875 (I34457,I34277,I34439);
nand I_1876 (I34475,I34421,I34457);
DFFARX1 I_1877 (I34475,I691,I34043,I34502,);
nor I_1878 (I34511,I34439,I34169);
DFFARX1 I_1879 (I34511,I691,I34043,I34538,);
nor I_1880 (I34547,I33926,I33908);
DFFARX1 I_1881 (I34547,I691,I34043,I34574,);
DFFARX1 I_1882 (I34574,I691,I34043,I34592,);
not I_1883 (I34601,I34574);
nand I_1884 (I34619,I34601,I34079);
nand I_1885 (I34637,I34601,I34187);
not I_1886 (I34655,I698);
DFFARX1 I_1887 (I34502,I691,I34655,I34682,);
not I_1888 (I34691,I34682);
nand I_1889 (I34709,I34232,I34403);
and I_1890 (I34727,I34709,I34592);
DFFARX1 I_1891 (I34727,I691,I34655,I34754,);
DFFARX1 I_1892 (I34538,I691,I34655,I34772,);
and I_1893 (I34781,I34772,I34349);
nor I_1894 (I34799,I34754,I34781);
DFFARX1 I_1895 (I34799,I691,I34655,I34826,);
nand I_1896 (I34835,I34772,I34349);
nand I_1897 (I34853,I34691,I34835);
not I_1898 (I34871,I34853);
DFFARX1 I_1899 (I34538,I691,I34655,I34898,);
DFFARX1 I_1900 (I34898,I691,I34655,I34916,);
nand I_1901 (I34925,I34295,I34637);
and I_1902 (I34943,I34925,I34619);
DFFARX1 I_1903 (I34943,I691,I34655,I34970,);
DFFARX1 I_1904 (I34970,I691,I34655,I34988,);
not I_1905 (I34997,I34988);
not I_1906 (I35015,I34970);
nand I_1907 (I35033,I35015,I34835);
nor I_1908 (I35051,I34295,I34637);
not I_1909 (I35069,I35051);
nor I_1910 (I35087,I35015,I35069);
nor I_1911 (I35105,I34691,I35087);
DFFARX1 I_1912 (I35105,I691,I34655,I35132,);
nor I_1913 (I35141,I34754,I35069);
nor I_1914 (I35159,I34970,I35141);
nor I_1915 (I35177,I34898,I35051);
nor I_1916 (I35195,I34754,I35051);
not I_1917 (I35213,I698);
DFFARX1 I_1918 (I34826,I691,I35213,I35240,);
DFFARX1 I_1919 (I35159,I691,I35213,I35258,);
not I_1920 (I35267,I35258);
not I_1921 (I35285,I34997);
nor I_1922 (I35303,I35285,I35195);
not I_1923 (I35321,I35033);
nor I_1924 (I35339,I35303,I35177);
nor I_1925 (I35357,I35258,I35339);
DFFARX1 I_1926 (I35357,I691,I35213,I35384,);
nor I_1927 (I35393,I35177,I35195);
nand I_1928 (I35411,I35393,I34997);
DFFARX1 I_1929 (I35411,I691,I35213,I35438,);
nor I_1930 (I35447,I35321,I35177);
nand I_1931 (I35465,I35447,I34916);
nor I_1932 (I35483,I35240,I35465);
DFFARX1 I_1933 (I35483,I691,I35213,I35510,);
not I_1934 (I35519,I35465);
nand I_1935 (I35537,I35258,I35519);
DFFARX1 I_1936 (I35465,I691,I35213,I35564,);
not I_1937 (I35573,I35564);
not I_1938 (I35591,I35177);
not I_1939 (I35609,I35195);
nor I_1940 (I35627,I35609,I35033);
nor I_1941 (I35645,I35573,I35627);
nor I_1942 (I35663,I35609,I34871);
and I_1943 (I35681,I35663,I34826);
or I_1944 (I35699,I35681,I35132);
DFFARX1 I_1945 (I35699,I691,I35213,I35726,);
nor I_1946 (I35735,I35726,I35240);
not I_1947 (I35753,I35726);
and I_1948 (I35771,I35753,I35240);
nor I_1949 (I35789,I35267,I35771);
nand I_1950 (I35807,I35753,I35321);
nor I_1951 (I35825,I35609,I35807);
nand I_1952 (I35843,I35753,I35519);
nand I_1953 (I35861,I35321,I35195);
nor I_1954 (I35879,I35591,I35861);
not I_1955 (I35897,I698);
DFFARX1 I_1956 (I35438,I691,I35897,I35924,);
not I_1957 (I35933,I35924);
nand I_1958 (I35951,I35510,I35735);
and I_1959 (I35969,I35951,I35645);
DFFARX1 I_1960 (I35969,I691,I35897,I35996,);
not I_1961 (I36005,I35537);
DFFARX1 I_1962 (I35825,I691,I35897,I36032,);
not I_1963 (I36041,I36032);
nor I_1964 (I36059,I36041,I35933);
and I_1965 (I36077,I36059,I35537);
nor I_1966 (I36095,I36041,I36005);
nor I_1967 (I36113,I35996,I36095);
DFFARX1 I_1968 (I35510,I691,I35897,I36140,);
nor I_1969 (I36149,I36140,I35996);
not I_1970 (I36167,I36149);
not I_1971 (I36185,I36140);
nor I_1972 (I36203,I36185,I36077);
DFFARX1 I_1973 (I36203,I691,I35897,I36230,);
nand I_1974 (I36239,I35879,I35789);
and I_1975 (I36257,I36239,I35384);
DFFARX1 I_1976 (I36257,I691,I35897,I36284,);
nor I_1977 (I36293,I36284,I36140);
DFFARX1 I_1978 (I36293,I691,I35897,I36320,);
nand I_1979 (I36329,I36284,I36185);
nand I_1980 (I36347,I36167,I36329);
not I_1981 (I36365,I36284);
nor I_1982 (I36383,I36365,I36077);
DFFARX1 I_1983 (I36383,I691,I35897,I36410,);
nor I_1984 (I36419,I35843,I35789);
or I_1985 (I36437,I36140,I36419);
nor I_1986 (I36455,I36284,I36419);
or I_1987 (I36473,I35996,I36419);
DFFARX1 I_1988 (I36419,I691,I35897,I36500,);
not I_1989 (I36509,I698);
DFFARX1 I_1990 (I36320,I691,I36509,I36536,);
not I_1991 (I36545,I36536);
DFFARX1 I_1992 (I36437,I691,I36509,I36572,);
not I_1993 (I36581,I36455);
nand I_1994 (I36599,I36581,I36473);
not I_1995 (I36617,I36599);
nor I_1996 (I36635,I36617,I36347);
nor I_1997 (I36653,I36545,I36635);
DFFARX1 I_1998 (I36653,I691,I36509,I36680,);
not I_1999 (I36689,I36347);
nand I_2000 (I36707,I36689,I36617);
and I_2001 (I36725,I36689,I36455);
nand I_2002 (I36743,I36725,I36113);
nor I_2003 (I36761,I36743,I36689);
and I_2004 (I36779,I36572,I36743);
not I_2005 (I36797,I36743);
nand I_2006 (I36815,I36572,I36797);
nor I_2007 (I36833,I36536,I36743);
not I_2008 (I36851,I36410);
nor I_2009 (I36869,I36851,I36455);
nand I_2010 (I36887,I36869,I36689);
nor I_2011 (I36905,I36599,I36887);
nor I_2012 (I36923,I36851,I36320);
and I_2013 (I36941,I36923,I36230);
or I_2014 (I36959,I36941,I36500);
DFFARX1 I_2015 (I36959,I691,I36509,I36986,);
nor I_2016 (I36995,I36986,I36707);
DFFARX1 I_2017 (I36995,I691,I36509,I37022,);
DFFARX1 I_2018 (I36986,I691,I36509,I37040,);
not I_2019 (I37049,I36986);
nor I_2020 (I37067,I37049,I36572);
nor I_2021 (I37085,I36869,I37067);
DFFARX1 I_2022 (I37085,I691,I36509,I37112,);
not I_2023 (I37121,I698);
DFFARX1 I_2024 (I36761,I691,I37121,I37148,);
DFFARX1 I_2025 (I37148,I691,I37121,I37166,);
not I_2026 (I37175,I37166);
not I_2027 (I37193,I37148);
DFFARX1 I_2028 (I36779,I691,I37121,I37220,);
not I_2029 (I37229,I37220);
and I_2030 (I37247,I37193,I37040);
not I_2031 (I37265,I37112);
nand I_2032 (I37283,I37265,I37040);
not I_2033 (I37301,I37022);
nor I_2034 (I37319,I37301,I36833);
nand I_2035 (I37337,I37319,I36905);
nor I_2036 (I37355,I37337,I37283);
DFFARX1 I_2037 (I37355,I691,I37121,I37382,);
not I_2038 (I37391,I37337);
not I_2039 (I37409,I36833);
nand I_2040 (I37427,I37409,I37040);
nor I_2041 (I37445,I36833,I37112);
nand I_2042 (I37463,I37247,I37445);
nand I_2043 (I37481,I37193,I36833);
nand I_2044 (I37499,I37301,I36680);
DFFARX1 I_2045 (I37499,I691,I37121,I37526,);
DFFARX1 I_2046 (I37499,I691,I37121,I37544,);
not I_2047 (I37553,I36680);
nor I_2048 (I37571,I37553,I37022);
and I_2049 (I37589,I37571,I36815);
or I_2050 (I37607,I37589,I36833);
DFFARX1 I_2051 (I37607,I691,I37121,I37634,);
nand I_2052 (I37643,I37634,I37265);
nor I_2053 (I37661,I37643,I37427);
nor I_2054 (I37679,I37634,I37229);
DFFARX1 I_2055 (I37634,I691,I37121,I37706,);
not I_2056 (I37715,I37706);
nor I_2057 (I37733,I37715,I37391);
not I_2058 (I37751,I698);
DFFARX1 I_2059 (I37481,I691,I37751,I37778,);
not I_2060 (I37787,I37778);
nand I_2061 (I37805,I37679,I37526);
and I_2062 (I37823,I37805,I37463);
DFFARX1 I_2063 (I37823,I691,I37751,I37850,);
DFFARX1 I_2064 (I37850,I691,I37751,I37868,);
DFFARX1 I_2065 (I37733,I691,I37751,I37886,);
nand I_2066 (I37895,I37886,I37544);
not I_2067 (I37913,I37895);
DFFARX1 I_2068 (I37913,I691,I37751,I37940,);
not I_2069 (I37949,I37940);
nor I_2070 (I37967,I37787,I37949);
DFFARX1 I_2071 (I37661,I691,I37751,I37994,);
nor I_2072 (I38003,I37994,I37850);
nor I_2073 (I38021,I37994,I37913);
nand I_2074 (I38039,I37382,I37175);
and I_2075 (I38057,I38039,I37679);
DFFARX1 I_2076 (I38057,I691,I37751,I38084,);
not I_2077 (I38093,I38084);
nand I_2078 (I38111,I38093,I37994);
nand I_2079 (I38129,I38093,I37895);
nor I_2080 (I38147,I37382,I37175);
and I_2081 (I38165,I37994,I38147);
nor I_2082 (I38183,I38093,I38165);
DFFARX1 I_2083 (I38183,I691,I37751,I38210,);
nor I_2084 (I38219,I37778,I38147);
DFFARX1 I_2085 (I38219,I691,I37751,I38246,);
nor I_2086 (I38255,I38084,I38147);
not I_2087 (I38273,I38255);
nand I_2088 (I38291,I38273,I38111);
not I_2089 (I38309,I698);
DFFARX1 I_2090 (I38291,I691,I38309,I38336,);
DFFARX1 I_2091 (I38129,I691,I38309,I38354,);
not I_2092 (I38363,I38354);
nor I_2093 (I38381,I38336,I38363);
DFFARX1 I_2094 (I38363,I691,I38309,I38408,);
nor I_2095 (I38417,I37967,I38021);
and I_2096 (I38435,I38417,I38246);
nor I_2097 (I38453,I38435,I37967);
not I_2098 (I38471,I37967);
and I_2099 (I38489,I38471,I38129);
nand I_2100 (I38507,I38489,I37868);
nor I_2101 (I38525,I38471,I38507);
DFFARX1 I_2102 (I38525,I691,I38309,I38552,);
not I_2103 (I38561,I38507);
nand I_2104 (I38579,I38363,I38561);
nand I_2105 (I38597,I38435,I38561);
DFFARX1 I_2106 (I38471,I691,I38309,I38624,);
not I_2107 (I38633,I38003);
nor I_2108 (I38651,I38633,I38129);
nor I_2109 (I38669,I38651,I38453);
DFFARX1 I_2110 (I38669,I691,I38309,I38696,);
not I_2111 (I38705,I38651);
DFFARX1 I_2112 (I38705,I691,I38309,I38732,);
not I_2113 (I38741,I38732);
nor I_2114 (I38759,I38741,I38651);
nor I_2115 (I38777,I38633,I38246);
and I_2116 (I38795,I38777,I38210);
or I_2117 (I38813,I38795,I38021);
DFFARX1 I_2118 (I38813,I691,I38309,I38840,);
not I_2119 (I38849,I38840);
nand I_2120 (I38867,I38849,I38561);
not I_2121 (I38885,I38867);
nand I_2122 (I38903,I38867,I38579);
nand I_2123 (I38921,I38849,I38435);
not I_2124 (I38939,I698);
DFFARX1 I_2125 (I38885,I691,I38939,I38966,);
not I_2126 (I38975,I38966);
nand I_2127 (I38993,I38597,I38759);
and I_2128 (I39011,I38993,I38552);
DFFARX1 I_2129 (I39011,I691,I38939,I39038,);
DFFARX1 I_2130 (I39038,I691,I38939,I39056,);
DFFARX1 I_2131 (I38381,I691,I38939,I39074,);
nand I_2132 (I39083,I39074,I38408);
not I_2133 (I39101,I39083);
DFFARX1 I_2134 (I39101,I691,I38939,I39128,);
not I_2135 (I39137,I39128);
nor I_2136 (I39155,I38975,I39137);
DFFARX1 I_2137 (I38696,I691,I38939,I39182,);
nor I_2138 (I39191,I39182,I39038);
nor I_2139 (I39209,I39182,I39101);
nand I_2140 (I39227,I38921,I38624);
and I_2141 (I39245,I39227,I38903);
DFFARX1 I_2142 (I39245,I691,I38939,I39272,);
not I_2143 (I39281,I39272);
nand I_2144 (I39299,I39281,I39182);
nand I_2145 (I39317,I39281,I39083);
nor I_2146 (I39335,I38552,I38624);
and I_2147 (I39353,I39182,I39335);
nor I_2148 (I39371,I39281,I39353);
DFFARX1 I_2149 (I39371,I691,I38939,I39398,);
nor I_2150 (I39407,I38966,I39335);
DFFARX1 I_2151 (I39407,I691,I38939,I39434,);
nor I_2152 (I39443,I39272,I39335);
not I_2153 (I39461,I39443);
nand I_2154 (I39479,I39461,I39299);
not I_2155 (I39497,I698);
DFFARX1 I_2156 (I39191,I691,I39497,I39524,);
DFFARX1 I_2157 (I39524,I691,I39497,I39542,);
not I_2158 (I39551,I39542);
not I_2159 (I39569,I39524);
nand I_2160 (I39587,I39317,I39209);
and I_2161 (I39605,I39587,I39056);
DFFARX1 I_2162 (I39605,I691,I39497,I39632,);
not I_2163 (I39641,I39632);
DFFARX1 I_2164 (I39317,I691,I39497,I39668,);
and I_2165 (I39677,I39668,I39434);
nand I_2166 (I39695,I39668,I39434);
nand I_2167 (I39713,I39641,I39695);
DFFARX1 I_2168 (I39434,I691,I39497,I39740,);
nor I_2169 (I39749,I39740,I39677);
DFFARX1 I_2170 (I39749,I691,I39497,I39776,);
nor I_2171 (I39785,I39740,I39632);
nand I_2172 (I39803,I39398,I39479);
and I_2173 (I39821,I39803,I39209);
DFFARX1 I_2174 (I39821,I691,I39497,I39848,);
nor I_2175 (I39857,I39848,I39740);
not I_2176 (I39875,I39848);
nor I_2177 (I39893,I39875,I39641);
nor I_2178 (I39911,I39569,I39893);
DFFARX1 I_2179 (I39911,I691,I39497,I39938,);
nor I_2180 (I39947,I39875,I39740);
nor I_2181 (I39965,I39155,I39479);
nor I_2182 (I39983,I39965,I39947);
not I_2183 (I40001,I39965);
nand I_2184 (I40019,I39695,I40001);
DFFARX1 I_2185 (I39965,I691,I39497,I40046,);
DFFARX1 I_2186 (I39965,I691,I39497,I40064,);
not I_2187 (I40073,I698);
DFFARX1 I_2188 (I40064,I691,I40073,I40100,);
DFFARX1 I_2189 (I40100,I691,I40073,I40118,);
not I_2190 (I40127,I40118);
not I_2191 (I40145,I40100);
DFFARX1 I_2192 (I40019,I691,I40073,I40172,);
not I_2193 (I40181,I40172);
and I_2194 (I40199,I40145,I40046);
not I_2195 (I40217,I39938);
nand I_2196 (I40235,I40217,I40046);
not I_2197 (I40253,I39983);
nor I_2198 (I40271,I40253,I39785);
nand I_2199 (I40289,I40271,I39776);
nor I_2200 (I40307,I40289,I40235);
DFFARX1 I_2201 (I40307,I691,I40073,I40334,);
not I_2202 (I40343,I40289);
not I_2203 (I40361,I39785);
nand I_2204 (I40379,I40361,I40046);
nor I_2205 (I40397,I39785,I39938);
nand I_2206 (I40415,I40199,I40397);
nand I_2207 (I40433,I40145,I39785);
nand I_2208 (I40451,I40253,I39776);
DFFARX1 I_2209 (I40451,I691,I40073,I40478,);
DFFARX1 I_2210 (I40451,I691,I40073,I40496,);
not I_2211 (I40505,I39776);
nor I_2212 (I40523,I40505,I39713);
and I_2213 (I40541,I40523,I39857);
or I_2214 (I40559,I40541,I39551);
DFFARX1 I_2215 (I40559,I691,I40073,I40586,);
nand I_2216 (I40595,I40586,I40217);
nor I_2217 (I40613,I40595,I40379);
nor I_2218 (I40631,I40586,I40181);
DFFARX1 I_2219 (I40586,I691,I40073,I40658,);
not I_2220 (I40667,I40658);
nor I_2221 (I40685,I40667,I40343);
not I_2222 (I40703,I698);
DFFARX1 I_2223 (I40415,I691,I40703,I40730,);
not I_2224 (I40739,I40730);
nand I_2225 (I40757,I40433,I40334);
and I_2226 (I40775,I40757,I40478);
DFFARX1 I_2227 (I40775,I691,I40703,I40802,);
DFFARX1 I_2228 (I40685,I691,I40703,I40820,);
and I_2229 (I40829,I40820,I40496);
nor I_2230 (I40847,I40802,I40829);
DFFARX1 I_2231 (I40847,I691,I40703,I40874,);
nand I_2232 (I40883,I40820,I40496);
nand I_2233 (I40901,I40739,I40883);
not I_2234 (I40919,I40901);
DFFARX1 I_2235 (I40334,I691,I40703,I40946,);
DFFARX1 I_2236 (I40946,I691,I40703,I40964,);
nand I_2237 (I40973,I40631,I40631);
and I_2238 (I40991,I40973,I40127);
DFFARX1 I_2239 (I40991,I691,I40703,I41018,);
DFFARX1 I_2240 (I41018,I691,I40703,I41036,);
not I_2241 (I41045,I41036);
not I_2242 (I41063,I41018);
nand I_2243 (I41081,I41063,I40883);
nor I_2244 (I41099,I40613,I40631);
not I_2245 (I41117,I41099);
nor I_2246 (I41135,I41063,I41117);
nor I_2247 (I41153,I40739,I41135);
DFFARX1 I_2248 (I41153,I691,I40703,I41180,);
nor I_2249 (I41189,I40802,I41117);
nor I_2250 (I41207,I41018,I41189);
nor I_2251 (I41225,I40946,I41099);
nor I_2252 (I41243,I40802,I41099);
not I_2253 (I41261,I698);
DFFARX1 I_2254 (I41045,I691,I41261,I41288,);
and I_2255 (I41297,I41288,I40874);
DFFARX1 I_2256 (I41297,I691,I41261,I41324,);
DFFARX1 I_2257 (I41180,I691,I41261,I41342,);
not I_2258 (I41351,I41207);
not I_2259 (I41369,I41243);
nand I_2260 (I41387,I41369,I41351);
nor I_2261 (I41405,I41342,I41387);
DFFARX1 I_2262 (I41387,I691,I41261,I41432,);
not I_2263 (I41441,I41432);
not I_2264 (I41459,I40919);
nand I_2265 (I41477,I41369,I41459);
DFFARX1 I_2266 (I41477,I691,I41261,I41504,);
not I_2267 (I41513,I41504);
not I_2268 (I41531,I41243);
nand I_2269 (I41549,I41531,I40964);
and I_2270 (I41567,I41351,I41549);
nor I_2271 (I41585,I41477,I41567);
DFFARX1 I_2272 (I41585,I691,I41261,I41612,);
DFFARX1 I_2273 (I41567,I691,I41261,I41630,);
nor I_2274 (I41639,I41243,I41225);
nor I_2275 (I41657,I41477,I41639);
or I_2276 (I41675,I41243,I41225);
nor I_2277 (I41693,I41081,I40874);
DFFARX1 I_2278 (I41693,I691,I41261,I41720,);
not I_2279 (I41729,I41720);
nor I_2280 (I41747,I41729,I41513);
nand I_2281 (I41765,I41729,I41342);
not I_2282 (I41783,I41081);
nand I_2283 (I41801,I41783,I41459);
nand I_2284 (I41819,I41729,I41801);
nand I_2285 (I41837,I41819,I41765);
nand I_2286 (I41855,I41801,I41675);
not I_2287 (I41873,I698);
DFFARX1 I_2288 (I41441,I691,I41873,I41900,);
DFFARX1 I_2289 (I41900,I691,I41873,I41918,);
not I_2290 (I41927,I41918);
nand I_2291 (I41945,I41657,I41405);
and I_2292 (I41963,I41945,I41612);
DFFARX1 I_2293 (I41963,I691,I41873,I41990,);
DFFARX1 I_2294 (I41990,I691,I41873,I42008,);
DFFARX1 I_2295 (I41990,I691,I41873,I42026,);
DFFARX1 I_2296 (I41855,I691,I41873,I42044,);
nand I_2297 (I42053,I42044,I41747);
not I_2298 (I42071,I42053);
nor I_2299 (I42089,I41900,I42071);
DFFARX1 I_2300 (I41324,I691,I41873,I42116,);
not I_2301 (I42125,I42116);
nor I_2302 (I42143,I42125,I41927);
nand I_2303 (I42161,I42125,I42053);
nand I_2304 (I42179,I41837,I41405);
and I_2305 (I42197,I42179,I41630);
DFFARX1 I_2306 (I42197,I691,I41873,I42224,);
nor I_2307 (I42233,I42224,I41900);
DFFARX1 I_2308 (I42233,I691,I41873,I42260,);
not I_2309 (I42269,I42224);
nor I_2310 (I42287,I41612,I41405);
not I_2311 (I42305,I42287);
nor I_2312 (I42323,I42053,I42305);
nor I_2313 (I42341,I42269,I42323);
DFFARX1 I_2314 (I42341,I691,I41873,I42368,);
nor I_2315 (I42377,I42224,I42305);
nor I_2316 (I42395,I42071,I42377);
nor I_2317 (I42413,I42224,I42287);
not I_2318 (I42431,I698);
DFFARX1 I_2319 (I42260,I691,I42431,I42458,);
DFFARX1 I_2320 (I42161,I691,I42431,I42476,);
not I_2321 (I42485,I42476);
not I_2322 (I42503,I42260);
nor I_2323 (I42521,I42503,I42089);
not I_2324 (I42539,I42026);
nor I_2325 (I42557,I42521,I42143);
nor I_2326 (I42575,I42476,I42557);
DFFARX1 I_2327 (I42575,I691,I42431,I42602,);
nor I_2328 (I42611,I42143,I42089);
nand I_2329 (I42629,I42611,I42260);
DFFARX1 I_2330 (I42629,I691,I42431,I42656,);
nor I_2331 (I42665,I42539,I42143);
nand I_2332 (I42683,I42665,I42413);
nor I_2333 (I42701,I42458,I42683);
DFFARX1 I_2334 (I42701,I691,I42431,I42728,);
not I_2335 (I42737,I42683);
nand I_2336 (I42755,I42476,I42737);
DFFARX1 I_2337 (I42683,I691,I42431,I42782,);
not I_2338 (I42791,I42782);
not I_2339 (I42809,I42143);
not I_2340 (I42827,I42413);
nor I_2341 (I42845,I42827,I42026);
nor I_2342 (I42863,I42791,I42845);
nor I_2343 (I42881,I42827,I42368);
and I_2344 (I42899,I42881,I42008);
or I_2345 (I42917,I42899,I42395);
DFFARX1 I_2346 (I42917,I691,I42431,I42944,);
nor I_2347 (I42953,I42944,I42458);
not I_2348 (I42971,I42944);
and I_2349 (I42989,I42971,I42458);
nor I_2350 (I43007,I42485,I42989);
nand I_2351 (I43025,I42971,I42539);
nor I_2352 (I43043,I42827,I43025);
nand I_2353 (I43061,I42971,I42737);
nand I_2354 (I43079,I42539,I42413);
nor I_2355 (I43097,I42809,I43079);
not I_2356 (I43115,I698);
DFFARX1 I_2357 (I43061,I691,I43115,I43142,);
DFFARX1 I_2358 (I42656,I691,I43115,I43160,);
not I_2359 (I43169,I43160);
nor I_2360 (I43187,I43142,I43169);
DFFARX1 I_2361 (I43169,I691,I43115,I43214,);
nor I_2362 (I43223,I43043,I42953);
and I_2363 (I43241,I43223,I42728);
nor I_2364 (I43259,I43241,I43043);
not I_2365 (I43277,I43043);
and I_2366 (I43295,I43277,I43007);
nand I_2367 (I43313,I43295,I42602);
nor I_2368 (I43331,I43277,I43313);
DFFARX1 I_2369 (I43331,I691,I43115,I43358,);
not I_2370 (I43367,I43313);
nand I_2371 (I43385,I43169,I43367);
nand I_2372 (I43403,I43241,I43367);
DFFARX1 I_2373 (I43277,I691,I43115,I43430,);
not I_2374 (I43439,I42755);
nor I_2375 (I43457,I43439,I43007);
nor I_2376 (I43475,I43457,I43259);
DFFARX1 I_2377 (I43475,I691,I43115,I43502,);
not I_2378 (I43511,I43457);
DFFARX1 I_2379 (I43511,I691,I43115,I43538,);
not I_2380 (I43547,I43538);
nor I_2381 (I43565,I43547,I43457);
nor I_2382 (I43583,I43439,I42728);
and I_2383 (I43601,I43583,I42863);
or I_2384 (I43619,I43601,I43097);
DFFARX1 I_2385 (I43619,I691,I43115,I43646,);
not I_2386 (I43655,I43646);
nand I_2387 (I43673,I43655,I43367);
not I_2388 (I43691,I43673);
nand I_2389 (I43709,I43673,I43385);
nand I_2390 (I43727,I43655,I43241);
not I_2391 (I43745,I698);
DFFARX1 I_2392 (I43430,I691,I43745,I43772,);
and I_2393 (I43781,I43772,I43709);
DFFARX1 I_2394 (I43781,I691,I43745,I43808,);
DFFARX1 I_2395 (I43358,I691,I43745,I43826,);
not I_2396 (I43835,I43691);
not I_2397 (I43853,I43187);
nand I_2398 (I43871,I43853,I43835);
nor I_2399 (I43889,I43826,I43871);
DFFARX1 I_2400 (I43871,I691,I43745,I43916,);
not I_2401 (I43925,I43916);
not I_2402 (I43943,I43403);
nand I_2403 (I43961,I43853,I43943);
DFFARX1 I_2404 (I43961,I691,I43745,I43988,);
not I_2405 (I43997,I43988);
not I_2406 (I44015,I43565);
nand I_2407 (I44033,I44015,I43358);
and I_2408 (I44051,I43835,I44033);
nor I_2409 (I44069,I43961,I44051);
DFFARX1 I_2410 (I44069,I691,I43745,I44096,);
DFFARX1 I_2411 (I44051,I691,I43745,I44114,);
nor I_2412 (I44123,I43565,I43502);
nor I_2413 (I44141,I43961,I44123);
or I_2414 (I44159,I43565,I43502);
nor I_2415 (I44177,I43214,I43727);
DFFARX1 I_2416 (I44177,I691,I43745,I44204,);
not I_2417 (I44213,I44204);
nor I_2418 (I44231,I44213,I43997);
nand I_2419 (I44249,I44213,I43826);
not I_2420 (I44267,I43214);
nand I_2421 (I44285,I44267,I43943);
nand I_2422 (I44303,I44213,I44285);
nand I_2423 (I44321,I44303,I44249);
nand I_2424 (I44339,I44285,I44159);
not I_2425 (I44357,I698);
DFFARX1 I_2426 (I44339,I691,I44357,I44384,);
not I_2427 (I44393,I44384);
nand I_2428 (I44411,I44114,I44096);
and I_2429 (I44429,I44411,I43889);
DFFARX1 I_2430 (I44429,I691,I44357,I44456,);
DFFARX1 I_2431 (I43925,I691,I44357,I44474,);
and I_2432 (I44483,I44474,I43889);
nor I_2433 (I44501,I44456,I44483);
DFFARX1 I_2434 (I44501,I691,I44357,I44528,);
nand I_2435 (I44537,I44474,I43889);
nand I_2436 (I44555,I44393,I44537);
not I_2437 (I44573,I44555);
DFFARX1 I_2438 (I44096,I691,I44357,I44600,);
DFFARX1 I_2439 (I44600,I691,I44357,I44618,);
nand I_2440 (I44627,I44141,I44321);
and I_2441 (I44645,I44627,I43808);
DFFARX1 I_2442 (I44645,I691,I44357,I44672,);
DFFARX1 I_2443 (I44672,I691,I44357,I44690,);
not I_2444 (I44699,I44690);
not I_2445 (I44717,I44672);
nand I_2446 (I44735,I44717,I44537);
nor I_2447 (I44753,I44231,I44321);
not I_2448 (I44771,I44753);
nor I_2449 (I44789,I44717,I44771);
nor I_2450 (I44807,I44393,I44789);
DFFARX1 I_2451 (I44807,I691,I44357,I44834,);
nor I_2452 (I44843,I44456,I44771);
nor I_2453 (I44861,I44672,I44843);
nor I_2454 (I44879,I44600,I44753);
nor I_2455 (I44897,I44456,I44753);
not I_2456 (I44915,I698);
DFFARX1 I_2457 (I44897,I691,I44915,I44942,);
not I_2458 (I44951,I44942);
nand I_2459 (I44969,I44573,I44618);
and I_2460 (I44987,I44969,I44528);
DFFARX1 I_2461 (I44987,I691,I44915,I45014,);
not I_2462 (I45023,I44897);
DFFARX1 I_2463 (I44834,I691,I44915,I45050,);
not I_2464 (I45059,I45050);
nor I_2465 (I45077,I45059,I44951);
and I_2466 (I45095,I45077,I44897);
nor I_2467 (I45113,I45059,I45023);
nor I_2468 (I45131,I45014,I45113);
DFFARX1 I_2469 (I44735,I691,I44915,I45158,);
nor I_2470 (I45167,I45158,I45014);
not I_2471 (I45185,I45167);
not I_2472 (I45203,I45158);
nor I_2473 (I45221,I45203,I45095);
DFFARX1 I_2474 (I45221,I691,I44915,I45248,);
nand I_2475 (I45257,I44699,I44528);
and I_2476 (I45275,I45257,I44861);
DFFARX1 I_2477 (I45275,I691,I44915,I45302,);
nor I_2478 (I45311,I45302,I45158);
DFFARX1 I_2479 (I45311,I691,I44915,I45338,);
nand I_2480 (I45347,I45302,I45203);
nand I_2481 (I45365,I45185,I45347);
not I_2482 (I45383,I45302);
nor I_2483 (I45401,I45383,I45095);
DFFARX1 I_2484 (I45401,I691,I44915,I45428,);
nor I_2485 (I45437,I44879,I44528);
or I_2486 (I45455,I45158,I45437);
nor I_2487 (I45473,I45302,I45437);
or I_2488 (I45491,I45014,I45437);
DFFARX1 I_2489 (I45437,I691,I44915,I45518,);
not I_2490 (I45527,I698);
DFFARX1 I_2491 (I45428,I691,I45527,I45554,);
DFFARX1 I_2492 (I45473,I691,I45527,I45572,);
not I_2493 (I45581,I45572);
nor I_2494 (I45599,I45554,I45581);
DFFARX1 I_2495 (I45581,I691,I45527,I45626,);
nor I_2496 (I45635,I45365,I45455);
and I_2497 (I45653,I45635,I45338);
nor I_2498 (I45671,I45653,I45365);
not I_2499 (I45689,I45365);
and I_2500 (I45707,I45689,I45248);
nand I_2501 (I45725,I45707,I45491);
nor I_2502 (I45743,I45689,I45725);
DFFARX1 I_2503 (I45743,I691,I45527,I45770,);
not I_2504 (I45779,I45725);
nand I_2505 (I45797,I45581,I45779);
nand I_2506 (I45815,I45653,I45779);
DFFARX1 I_2507 (I45689,I691,I45527,I45842,);
not I_2508 (I45851,I45473);
nor I_2509 (I45869,I45851,I45248);
nor I_2510 (I45887,I45869,I45671);
DFFARX1 I_2511 (I45887,I691,I45527,I45914,);
not I_2512 (I45923,I45869);
DFFARX1 I_2513 (I45923,I691,I45527,I45950,);
not I_2514 (I45959,I45950);
nor I_2515 (I45977,I45959,I45869);
nor I_2516 (I45995,I45851,I45131);
and I_2517 (I46013,I45995,I45518);
or I_2518 (I46031,I46013,I45338);
DFFARX1 I_2519 (I46031,I691,I45527,I46058,);
not I_2520 (I46067,I46058);
nand I_2521 (I46085,I46067,I45779);
not I_2522 (I46103,I46085);
nand I_2523 (I46121,I46085,I45797);
nand I_2524 (I46139,I46067,I45653);
not I_2525 (I46157,I698);
DFFARX1 I_2526 (I45770,I691,I46157,I46184,);
DFFARX1 I_2527 (I46184,I691,I46157,I46202,);
not I_2528 (I46211,I46202);
nand I_2529 (I46229,I45599,I46121);
and I_2530 (I46247,I46229,I45626);
DFFARX1 I_2531 (I46247,I691,I46157,I46274,);
DFFARX1 I_2532 (I46274,I691,I46157,I46292,);
DFFARX1 I_2533 (I46274,I691,I46157,I46310,);
DFFARX1 I_2534 (I45977,I691,I46157,I46328,);
nand I_2535 (I46337,I46328,I45815);
not I_2536 (I46355,I46337);
nor I_2537 (I46373,I46184,I46355);
DFFARX1 I_2538 (I45770,I691,I46157,I46400,);
not I_2539 (I46409,I46400);
nor I_2540 (I46427,I46409,I46211);
nand I_2541 (I46445,I46409,I46337);
nand I_2542 (I46463,I45842,I46139);
and I_2543 (I46481,I46463,I46103);
DFFARX1 I_2544 (I46481,I691,I46157,I46508,);
nor I_2545 (I46517,I46508,I46184);
DFFARX1 I_2546 (I46517,I691,I46157,I46544,);
not I_2547 (I46553,I46508);
nor I_2548 (I46571,I45914,I46139);
not I_2549 (I46589,I46571);
nor I_2550 (I46607,I46337,I46589);
nor I_2551 (I46625,I46553,I46607);
DFFARX1 I_2552 (I46625,I691,I46157,I46652,);
nor I_2553 (I46661,I46508,I46589);
nor I_2554 (I46679,I46355,I46661);
nor I_2555 (I46697,I46508,I46571);
not I_2556 (I46715,I698);
DFFARX1 I_2557 (I46544,I691,I46715,I46742,);
nand I_2558 (I46751,I46310,I46697);
and I_2559 (I46769,I46751,I46544);
DFFARX1 I_2560 (I46769,I691,I46715,I46796,);
nor I_2561 (I46805,I46796,I46742);
not I_2562 (I46823,I46796);
DFFARX1 I_2563 (I46445,I691,I46715,I46850,);
nand I_2564 (I46859,I46850,I46292);
not I_2565 (I46877,I46859);
DFFARX1 I_2566 (I46877,I691,I46715,I46904,);
not I_2567 (I46913,I46904);
nor I_2568 (I46931,I46742,I46859);
nor I_2569 (I46949,I46796,I46931);
DFFARX1 I_2570 (I46679,I691,I46715,I46976,);
DFFARX1 I_2571 (I46976,I691,I46715,I46994,);
not I_2572 (I47003,I46994);
not I_2573 (I47021,I46976);
nand I_2574 (I47039,I47021,I46823);
nand I_2575 (I47057,I46652,I46697);
and I_2576 (I47075,I47057,I46373);
DFFARX1 I_2577 (I47075,I691,I46715,I47102,);
nor I_2578 (I47111,I47102,I46742);
DFFARX1 I_2579 (I47111,I691,I46715,I47138,);
DFFARX1 I_2580 (I47102,I691,I46715,I47156,);
nor I_2581 (I47165,I46427,I46697);
not I_2582 (I47183,I47165);
nor I_2583 (I47201,I47003,I47183);
nand I_2584 (I47219,I47021,I47183);
nor I_2585 (I47237,I46742,I47165);
DFFARX1 I_2586 (I47165,I691,I46715,I47264,);
not I_2587 (I47273,I698);
DFFARX1 I_2588 (I47237,I691,I47273,I47300,);
DFFARX1 I_2589 (I47300,I691,I47273,I47318,);
not I_2590 (I47327,I47318);
DFFARX1 I_2591 (I46805,I691,I47273,I47354,);
not I_2592 (I47363,I47219);
nor I_2593 (I47381,I47300,I47363);
not I_2594 (I47399,I46949);
not I_2595 (I47417,I47201);
nand I_2596 (I47435,I47417,I46949);
nor I_2597 (I47453,I47363,I47435);
nor I_2598 (I47471,I47354,I47453);
DFFARX1 I_2599 (I47417,I691,I47273,I47498,);
nor I_2600 (I47507,I47201,I47039);
nand I_2601 (I47525,I47507,I47138);
nor I_2602 (I47543,I47525,I47399);
nand I_2603 (I47561,I47543,I47219);
DFFARX1 I_2604 (I47525,I691,I47273,I47588,);
nand I_2605 (I47597,I47399,I47201);
nor I_2606 (I47615,I47399,I47201);
nand I_2607 (I47633,I47381,I47615);
not I_2608 (I47651,I47156);
nor I_2609 (I47669,I47651,I47597);
DFFARX1 I_2610 (I47669,I691,I47273,I47696,);
nor I_2611 (I47705,I47651,I47264);
and I_2612 (I47723,I47705,I46913);
or I_2613 (I47741,I47723,I47138);
DFFARX1 I_2614 (I47741,I691,I47273,I47768,);
nor I_2615 (I47777,I47768,I47354);
nor I_2616 (I47795,I47300,I47777);
not I_2617 (I47813,I47768);
nor I_2618 (I47831,I47813,I47471);
DFFARX1 I_2619 (I47831,I691,I47273,I47858,);
nand I_2620 (I47867,I47813,I47399);
nor I_2621 (I47885,I47651,I47867);
not I_2622 (I47903,I698);
DFFARX1 I_2623 (I452,I691,I47903,I47930,);
nand I_2624 (I47939,I47930,I260);
not I_2625 (I47957,I47939);
DFFARX1 I_2626 (I188,I691,I47903,I47984,);
not I_2627 (I47993,I47984);
not I_2628 (I48011,I284);
or I_2629 (I48029,I324,I284);
nor I_2630 (I48047,I324,I284);
or I_2631 (I48065,I236,I324);
DFFARX1 I_2632 (I48065,I691,I47903,I48092,);
not I_2633 (I48101,I532);
nand I_2634 (I48119,I48101,I404);
nand I_2635 (I48137,I48011,I48119);
and I_2636 (I48155,I47993,I48137);
nor I_2637 (I48173,I532,I636);
and I_2638 (I48191,I47993,I48173);
nor I_2639 (I48209,I47957,I48191);
DFFARX1 I_2640 (I48173,I691,I47903,I48236,);
not I_2641 (I48245,I48236);
nor I_2642 (I48263,I47993,I48245);
or I_2643 (I48281,I48065,I148);
nor I_2644 (I48299,I148,I236);
nand I_2645 (I48317,I48137,I48299);
nand I_2646 (I48335,I48281,I48317);
DFFARX1 I_2647 (I48335,I691,I47903,I48362,);
nor I_2648 (I48371,I48299,I48029);
DFFARX1 I_2649 (I48371,I691,I47903,I48398,);
nor I_2650 (I48407,I148,I220);
DFFARX1 I_2651 (I48407,I691,I47903,I48434,);
DFFARX1 I_2652 (I48434,I691,I47903,I48452,);
not I_2653 (I48461,I48434);
nand I_2654 (I48479,I48461,I47939);
nand I_2655 (I48497,I48461,I48047);
not I_2656 (I48515,I698);
DFFARX1 I_2657 (I48398,I691,I48515,I48542,);
not I_2658 (I48551,I48542);
nand I_2659 (I48569,I48092,I48497);
and I_2660 (I48587,I48569,I48479);
DFFARX1 I_2661 (I48587,I691,I48515,I48614,);
not I_2662 (I48623,I48263);
DFFARX1 I_2663 (I48155,I691,I48515,I48650,);
not I_2664 (I48659,I48650);
nor I_2665 (I48677,I48659,I48551);
and I_2666 (I48695,I48677,I48263);
nor I_2667 (I48713,I48659,I48623);
nor I_2668 (I48731,I48614,I48713);
DFFARX1 I_2669 (I48452,I691,I48515,I48758,);
nor I_2670 (I48767,I48758,I48614);
not I_2671 (I48785,I48767);
not I_2672 (I48803,I48758);
nor I_2673 (I48821,I48803,I48695);
DFFARX1 I_2674 (I48821,I691,I48515,I48848,);
nand I_2675 (I48857,I48362,I48209);
and I_2676 (I48875,I48857,I48155);
DFFARX1 I_2677 (I48875,I691,I48515,I48902,);
nor I_2678 (I48911,I48902,I48758);
DFFARX1 I_2679 (I48911,I691,I48515,I48938,);
nand I_2680 (I48947,I48902,I48803);
nand I_2681 (I48965,I48785,I48947);
not I_2682 (I48983,I48902);
nor I_2683 (I49001,I48983,I48695);
DFFARX1 I_2684 (I49001,I691,I48515,I49028,);
nor I_2685 (I49037,I48398,I48209);
or I_2686 (I49055,I48758,I49037);
nor I_2687 (I49073,I48902,I49037);
or I_2688 (I49091,I48614,I49037);
DFFARX1 I_2689 (I49037,I691,I48515,I49118,);
not I_2690 (I49127,I698);
DFFARX1 I_2691 (I48731,I691,I49127,I49154,);
and I_2692 (I49163,I49154,I49073);
DFFARX1 I_2693 (I49163,I691,I49127,I49190,);
DFFARX1 I_2694 (I49091,I691,I49127,I49208,);
not I_2695 (I49217,I48938);
not I_2696 (I49235,I49118);
nand I_2697 (I49253,I49235,I49217);
nor I_2698 (I49271,I49208,I49253);
DFFARX1 I_2699 (I49253,I691,I49127,I49298,);
not I_2700 (I49307,I49298);
not I_2701 (I49325,I49055);
nand I_2702 (I49343,I49235,I49325);
DFFARX1 I_2703 (I49343,I691,I49127,I49370,);
not I_2704 (I49379,I49370);
not I_2705 (I49397,I49028);
nand I_2706 (I49415,I49397,I48848);
and I_2707 (I49433,I49217,I49415);
nor I_2708 (I49451,I49343,I49433);
DFFARX1 I_2709 (I49451,I691,I49127,I49478,);
DFFARX1 I_2710 (I49433,I691,I49127,I49496,);
nor I_2711 (I49505,I49028,I48965);
nor I_2712 (I49523,I49343,I49505);
or I_2713 (I49541,I49028,I48965);
nor I_2714 (I49559,I48938,I49073);
DFFARX1 I_2715 (I49559,I691,I49127,I49586,);
not I_2716 (I49595,I49586);
nor I_2717 (I49613,I49595,I49379);
nand I_2718 (I49631,I49595,I49208);
not I_2719 (I49649,I48938);
nand I_2720 (I49667,I49649,I49325);
nand I_2721 (I49685,I49595,I49667);
nand I_2722 (I49703,I49685,I49631);
nand I_2723 (I49721,I49667,I49541);
not I_2724 (I49739,I698);
DFFARX1 I_2725 (I49307,I691,I49739,I49766,);
DFFARX1 I_2726 (I49766,I691,I49739,I49784,);
not I_2727 (I49793,I49784);
nand I_2728 (I49811,I49523,I49271);
and I_2729 (I49829,I49811,I49478);
DFFARX1 I_2730 (I49829,I691,I49739,I49856,);
DFFARX1 I_2731 (I49856,I691,I49739,I49874,);
DFFARX1 I_2732 (I49856,I691,I49739,I49892,);
DFFARX1 I_2733 (I49721,I691,I49739,I49910,);
nand I_2734 (I49919,I49910,I49613);
not I_2735 (I49937,I49919);
nor I_2736 (I49955,I49766,I49937);
DFFARX1 I_2737 (I49190,I691,I49739,I49982,);
not I_2738 (I49991,I49982);
nor I_2739 (I50009,I49991,I49793);
nand I_2740 (I50027,I49991,I49919);
nand I_2741 (I50045,I49703,I49271);
and I_2742 (I50063,I50045,I49496);
DFFARX1 I_2743 (I50063,I691,I49739,I50090,);
nor I_2744 (I50099,I50090,I49766);
DFFARX1 I_2745 (I50099,I691,I49739,I50126,);
not I_2746 (I50135,I50090);
nor I_2747 (I50153,I49478,I49271);
not I_2748 (I50171,I50153);
nor I_2749 (I50189,I49919,I50171);
nor I_2750 (I50207,I50135,I50189);
DFFARX1 I_2751 (I50207,I691,I49739,I50234,);
nor I_2752 (I50243,I50090,I50171);
nor I_2753 (I50261,I49937,I50243);
nor I_2754 (I50279,I50090,I50153);
not I_2755 (I50297,I698);
DFFARX1 I_2756 (I50126,I691,I50297,I50324,);
and I_2757 (I50333,I50324,I50279);
DFFARX1 I_2758 (I50333,I691,I50297,I50360,);
DFFARX1 I_2759 (I50279,I691,I50297,I50378,);
not I_2760 (I50387,I50027);
not I_2761 (I50405,I50234);
nand I_2762 (I50423,I50405,I50387);
nor I_2763 (I50441,I50378,I50423);
DFFARX1 I_2764 (I50423,I691,I50297,I50468,);
not I_2765 (I50477,I50468);
not I_2766 (I50495,I49892);
nand I_2767 (I50513,I50405,I50495);
DFFARX1 I_2768 (I50513,I691,I50297,I50540,);
not I_2769 (I50549,I50540);
not I_2770 (I50567,I50009);
nand I_2771 (I50585,I50567,I50126);
and I_2772 (I50603,I50387,I50585);
nor I_2773 (I50621,I50513,I50603);
DFFARX1 I_2774 (I50621,I691,I50297,I50648,);
DFFARX1 I_2775 (I50603,I691,I50297,I50666,);
nor I_2776 (I50675,I50009,I49955);
nor I_2777 (I50693,I50513,I50675);
or I_2778 (I50711,I50009,I49955);
nor I_2779 (I50729,I50261,I49874);
DFFARX1 I_2780 (I50729,I691,I50297,I50756,);
not I_2781 (I50765,I50756);
nor I_2782 (I50783,I50765,I50549);
nand I_2783 (I50801,I50765,I50378);
not I_2784 (I50819,I50261);
nand I_2785 (I50837,I50819,I50495);
nand I_2786 (I50855,I50765,I50837);
nand I_2787 (I50873,I50855,I50801);
nand I_2788 (I50891,I50837,I50711);
not I_2789 (I50909,I698);
DFFARX1 I_2790 (I50648,I691,I50909,I50936,);
DFFARX1 I_2791 (I50936,I691,I50909,I50954,);
not I_2792 (I50963,I50954);
not I_2793 (I50981,I50936);
DFFARX1 I_2794 (I50648,I691,I50909,I51008,);
not I_2795 (I51017,I51008);
and I_2796 (I51035,I50981,I50441);
not I_2797 (I51053,I50360);
nand I_2798 (I51071,I51053,I50441);
not I_2799 (I51089,I50666);
nor I_2800 (I51107,I51089,I50693);
nand I_2801 (I51125,I51107,I50783);
nor I_2802 (I51143,I51125,I51071);
DFFARX1 I_2803 (I51143,I691,I50909,I51170,);
not I_2804 (I51179,I51125);
not I_2805 (I51197,I50693);
nand I_2806 (I51215,I51197,I50441);
nor I_2807 (I51233,I50693,I50360);
nand I_2808 (I51251,I51035,I51233);
nand I_2809 (I51269,I50981,I50693);
nand I_2810 (I51287,I51089,I50873);
DFFARX1 I_2811 (I51287,I691,I50909,I51314,);
DFFARX1 I_2812 (I51287,I691,I50909,I51332,);
not I_2813 (I51341,I50873);
nor I_2814 (I51359,I51341,I50891);
and I_2815 (I51377,I51359,I50477);
or I_2816 (I51395,I51377,I50441);
DFFARX1 I_2817 (I51395,I691,I50909,I51422,);
nand I_2818 (I51431,I51422,I51053);
nor I_2819 (I51449,I51431,I51215);
nor I_2820 (I51467,I51422,I51017);
DFFARX1 I_2821 (I51422,I691,I50909,I51494,);
not I_2822 (I51503,I51494);
nor I_2823 (I51521,I51503,I51179);
not I_2824 (I51539,I698);
DFFARX1 I_2825 (I51170,I691,I51539,I51566,);
and I_2826 (I51575,I51566,I51467);
DFFARX1 I_2827 (I51575,I691,I51539,I51602,);
DFFARX1 I_2828 (I51467,I691,I51539,I51620,);
not I_2829 (I51629,I51521);
not I_2830 (I51647,I50963);
nand I_2831 (I51665,I51647,I51629);
nor I_2832 (I51683,I51620,I51665);
DFFARX1 I_2833 (I51665,I691,I51539,I51710,);
not I_2834 (I51719,I51710);
not I_2835 (I51737,I51251);
nand I_2836 (I51755,I51647,I51737);
DFFARX1 I_2837 (I51755,I691,I51539,I51782,);
not I_2838 (I51791,I51782);
not I_2839 (I51809,I51449);
nand I_2840 (I51827,I51809,I51269);
and I_2841 (I51845,I51629,I51827);
nor I_2842 (I51863,I51755,I51845);
DFFARX1 I_2843 (I51863,I691,I51539,I51890,);
DFFARX1 I_2844 (I51845,I691,I51539,I51908,);
nor I_2845 (I51917,I51449,I51170);
nor I_2846 (I51935,I51755,I51917);
or I_2847 (I51953,I51449,I51170);
nor I_2848 (I51971,I51332,I51314);
DFFARX1 I_2849 (I51971,I691,I51539,I51998,);
not I_2850 (I52007,I51998);
nor I_2851 (I52025,I52007,I51791);
nand I_2852 (I52043,I52007,I51620);
not I_2853 (I52061,I51332);
nand I_2854 (I52079,I52061,I51737);
nand I_2855 (I52097,I52007,I52079);
nand I_2856 (I52115,I52097,I52043);
nand I_2857 (I52133,I52079,I51953);
not I_2858 (I52151,I698);
DFFARX1 I_2859 (I51890,I691,I52151,I52178,);
DFFARX1 I_2860 (I52178,I691,I52151,I52196,);
not I_2861 (I52205,I52196);
not I_2862 (I52223,I52178);
DFFARX1 I_2863 (I51890,I691,I52151,I52250,);
not I_2864 (I52259,I52250);
and I_2865 (I52277,I52223,I51683);
not I_2866 (I52295,I51602);
nand I_2867 (I52313,I52295,I51683);
not I_2868 (I52331,I51908);
nor I_2869 (I52349,I52331,I51935);
nand I_2870 (I52367,I52349,I52025);
nor I_2871 (I52385,I52367,I52313);
DFFARX1 I_2872 (I52385,I691,I52151,I52412,);
not I_2873 (I52421,I52367);
not I_2874 (I52439,I51935);
nand I_2875 (I52457,I52439,I51683);
nor I_2876 (I52475,I51935,I51602);
nand I_2877 (I52493,I52277,I52475);
nand I_2878 (I52511,I52223,I51935);
nand I_2879 (I52529,I52331,I52115);
DFFARX1 I_2880 (I52529,I691,I52151,I52556,);
DFFARX1 I_2881 (I52529,I691,I52151,I52574,);
not I_2882 (I52583,I52115);
nor I_2883 (I52601,I52583,I52133);
and I_2884 (I52619,I52601,I51719);
or I_2885 (I52637,I52619,I51683);
DFFARX1 I_2886 (I52637,I691,I52151,I52664,);
nand I_2887 (I52673,I52664,I52295);
nor I_2888 (I52691,I52673,I52457);
nor I_2889 (I52709,I52664,I52259);
DFFARX1 I_2890 (I52664,I691,I52151,I52736,);
not I_2891 (I52745,I52736);
nor I_2892 (I52763,I52745,I52421);
not I_2893 (I52781,I698);
DFFARX1 I_2894 (I52574,I691,I52781,I52808,);
not I_2895 (I52817,I52808);
DFFARX1 I_2896 (I52412,I691,I52781,I52844,);
not I_2897 (I52853,I52763);
nand I_2898 (I52871,I52853,I52709);
not I_2899 (I52889,I52871);
nor I_2900 (I52907,I52889,I52412);
nor I_2901 (I52925,I52817,I52907);
DFFARX1 I_2902 (I52925,I691,I52781,I52952,);
not I_2903 (I52961,I52412);
nand I_2904 (I52979,I52961,I52889);
and I_2905 (I52997,I52961,I52709);
nand I_2906 (I53015,I52997,I52205);
nor I_2907 (I53033,I53015,I52961);
and I_2908 (I53051,I52844,I53015);
not I_2909 (I53069,I53015);
nand I_2910 (I53087,I52844,I53069);
nor I_2911 (I53105,I52808,I53015);
not I_2912 (I53123,I52493);
nor I_2913 (I53141,I53123,I52709);
nand I_2914 (I53159,I53141,I52961);
nor I_2915 (I53177,I52871,I53159);
nor I_2916 (I53195,I53123,I52511);
and I_2917 (I53213,I53195,I52556);
or I_2918 (I53231,I53213,I52691);
DFFARX1 I_2919 (I53231,I691,I52781,I53258,);
nor I_2920 (I53267,I53258,I52979);
DFFARX1 I_2921 (I53267,I691,I52781,I53294,);
DFFARX1 I_2922 (I53258,I691,I52781,I53312,);
not I_2923 (I53321,I53258);
nor I_2924 (I53339,I53321,I52844);
nor I_2925 (I53357,I53141,I53339);
DFFARX1 I_2926 (I53357,I691,I52781,I53384,);
not I_2927 (I53393,I698);
DFFARX1 I_2928 (I53033,I691,I53393,I53420,);
and I_2929 (I53429,I53420,I53105);
DFFARX1 I_2930 (I53429,I691,I53393,I53456,);
DFFARX1 I_2931 (I52952,I691,I53393,I53474,);
not I_2932 (I53483,I53087);
not I_2933 (I53501,I53294);
nand I_2934 (I53519,I53501,I53483);
nor I_2935 (I53537,I53474,I53519);
DFFARX1 I_2936 (I53519,I691,I53393,I53564,);
not I_2937 (I53573,I53564);
not I_2938 (I53591,I53051);
nand I_2939 (I53609,I53501,I53591);
DFFARX1 I_2940 (I53609,I691,I53393,I53636,);
not I_2941 (I53645,I53636);
not I_2942 (I53663,I53384);
nand I_2943 (I53681,I53663,I53312);
and I_2944 (I53699,I53483,I53681);
nor I_2945 (I53717,I53609,I53699);
DFFARX1 I_2946 (I53717,I691,I53393,I53744,);
DFFARX1 I_2947 (I53699,I691,I53393,I53762,);
nor I_2948 (I53771,I53384,I53294);
nor I_2949 (I53789,I53609,I53771);
or I_2950 (I53807,I53384,I53294);
nor I_2951 (I53825,I53177,I53105);
DFFARX1 I_2952 (I53825,I691,I53393,I53852,);
not I_2953 (I53861,I53852);
nor I_2954 (I53879,I53861,I53645);
nand I_2955 (I53897,I53861,I53474);
not I_2956 (I53915,I53177);
nand I_2957 (I53933,I53915,I53591);
nand I_2958 (I53951,I53861,I53933);
nand I_2959 (I53969,I53951,I53897);
nand I_2960 (I53987,I53933,I53807);
not I_2961 (I54005,I698);
DFFARX1 I_2962 (I53456,I691,I54005,I54032,);
DFFARX1 I_2963 (I54032,I691,I54005,I54050,);
not I_2964 (I54059,I54050);
not I_2965 (I54077,I54032);
DFFARX1 I_2966 (I53987,I691,I54005,I54104,);
nand I_2967 (I54113,I54104,I53537);
not I_2968 (I54131,I53537);
not I_2969 (I54149,I53789);
nand I_2970 (I54167,I53762,I53537);
and I_2971 (I54185,I53762,I53537);
not I_2972 (I54203,I53744);
nand I_2973 (I54221,I54203,I54149);
nor I_2974 (I54239,I54221,I54113);
nor I_2975 (I54257,I54131,I54221);
nand I_2976 (I54275,I54185,I54257);
not I_2977 (I54293,I53969);
nor I_2978 (I54311,I54293,I53762);
nor I_2979 (I54329,I54311,I53744);
nor I_2980 (I54347,I54077,I54329);
DFFARX1 I_2981 (I54347,I691,I54005,I54374,);
not I_2982 (I54383,I54311);
DFFARX1 I_2983 (I54383,I691,I54005,I54410,);
and I_2984 (I54419,I54104,I54311);
nor I_2985 (I54437,I54293,I53573);
and I_2986 (I54455,I54437,I53744);
or I_2987 (I54473,I54455,I53879);
DFFARX1 I_2988 (I54473,I691,I54005,I54500,);
nor I_2989 (I54509,I54500,I54203);
DFFARX1 I_2990 (I54509,I691,I54005,I54536,);
nand I_2991 (I54545,I54500,I54104);
nand I_2992 (I54563,I54203,I54545);
nor I_2993 (I54581,I54563,I54167);
not I_2994 (I54599,I698);
DFFARX1 I_2995 (I54239,I691,I54599,I54626,);
nand I_2996 (I54635,I54536,I54239);
and I_2997 (I54653,I54635,I54419);
DFFARX1 I_2998 (I54653,I691,I54599,I54680,);
nor I_2999 (I54689,I54680,I54626);
not I_3000 (I54707,I54680);
DFFARX1 I_3001 (I54536,I691,I54599,I54734,);
nand I_3002 (I54743,I54734,I54410);
not I_3003 (I54761,I54743);
DFFARX1 I_3004 (I54761,I691,I54599,I54788,);
not I_3005 (I54797,I54788);
nor I_3006 (I54815,I54626,I54743);
nor I_3007 (I54833,I54680,I54815);
DFFARX1 I_3008 (I54275,I691,I54599,I54860,);
DFFARX1 I_3009 (I54860,I691,I54599,I54878,);
not I_3010 (I54887,I54878);
not I_3011 (I54905,I54860);
nand I_3012 (I54923,I54905,I54707);
nand I_3013 (I54941,I54374,I54059);
and I_3014 (I54959,I54941,I54275);
DFFARX1 I_3015 (I54959,I691,I54599,I54986,);
nor I_3016 (I54995,I54986,I54626);
DFFARX1 I_3017 (I54995,I691,I54599,I55022,);
DFFARX1 I_3018 (I54986,I691,I54599,I55040,);
nor I_3019 (I55049,I54581,I54059);
not I_3020 (I55067,I55049);
nor I_3021 (I55085,I54887,I55067);
nand I_3022 (I55103,I54905,I55067);
nor I_3023 (I55121,I54626,I55049);
DFFARX1 I_3024 (I55049,I691,I54599,I55148,);
not I_3025 (I55157,I698);
DFFARX1 I_3026 (I54797,I691,I55157,I55184,);
and I_3027 (I55193,I55184,I54923);
DFFARX1 I_3028 (I55193,I691,I55157,I55220,);
DFFARX1 I_3029 (I55040,I691,I55157,I55238,);
not I_3030 (I55247,I55022);
not I_3031 (I55265,I55085);
nand I_3032 (I55283,I55265,I55247);
nor I_3033 (I55301,I55238,I55283);
DFFARX1 I_3034 (I55283,I691,I55157,I55328,);
not I_3035 (I55337,I55328);
not I_3036 (I55355,I55148);
nand I_3037 (I55373,I55265,I55355);
DFFARX1 I_3038 (I55373,I691,I55157,I55400,);
not I_3039 (I55409,I55400);
not I_3040 (I55427,I55121);
nand I_3041 (I55445,I55427,I54689);
and I_3042 (I55463,I55247,I55445);
nor I_3043 (I55481,I55373,I55463);
DFFARX1 I_3044 (I55481,I691,I55157,I55508,);
DFFARX1 I_3045 (I55463,I691,I55157,I55526,);
nor I_3046 (I55535,I55121,I54833);
nor I_3047 (I55553,I55373,I55535);
or I_3048 (I55571,I55121,I54833);
nor I_3049 (I55589,I55103,I55022);
DFFARX1 I_3050 (I55589,I691,I55157,I55616,);
not I_3051 (I55625,I55616);
nor I_3052 (I55643,I55625,I55409);
nand I_3053 (I55661,I55625,I55238);
not I_3054 (I55679,I55103);
nand I_3055 (I55697,I55679,I55355);
nand I_3056 (I55715,I55625,I55697);
nand I_3057 (I55733,I55715,I55661);
nand I_3058 (I55751,I55697,I55571);
not I_3059 (I55769,I698);
DFFARX1 I_3060 (I55301,I691,I55769,I55796,);
DFFARX1 I_3061 (I55220,I691,I55769,I55814,);
not I_3062 (I55823,I55814);
nor I_3063 (I55841,I55796,I55823);
DFFARX1 I_3064 (I55823,I691,I55769,I55868,);
nor I_3065 (I55877,I55553,I55751);
and I_3066 (I55895,I55877,I55508);
nor I_3067 (I55913,I55895,I55553);
not I_3068 (I55931,I55553);
and I_3069 (I55949,I55931,I55733);
nand I_3070 (I55967,I55949,I55508);
nor I_3071 (I55985,I55931,I55967);
DFFARX1 I_3072 (I55985,I691,I55769,I56012,);
not I_3073 (I56021,I55967);
nand I_3074 (I56039,I55823,I56021);
nand I_3075 (I56057,I55895,I56021);
DFFARX1 I_3076 (I55931,I691,I55769,I56084,);
not I_3077 (I56093,I55337);
nor I_3078 (I56111,I56093,I55733);
nor I_3079 (I56129,I56111,I55913);
DFFARX1 I_3080 (I56129,I691,I55769,I56156,);
not I_3081 (I56165,I56111);
DFFARX1 I_3082 (I56165,I691,I55769,I56192,);
not I_3083 (I56201,I56192);
nor I_3084 (I56219,I56201,I56111);
nor I_3085 (I56237,I56093,I55643);
and I_3086 (I56255,I56237,I55526);
or I_3087 (I56273,I56255,I55301);
DFFARX1 I_3088 (I56273,I691,I55769,I56300,);
not I_3089 (I56309,I56300);
nand I_3090 (I56327,I56309,I56021);
not I_3091 (I56345,I56327);
nand I_3092 (I56363,I56327,I56039);
nand I_3093 (I56381,I56309,I55895);
not I_3094 (I56399,I698);
DFFARX1 I_3095 (I56084,I691,I56399,I56426,);
not I_3096 (I56435,I56426);
nand I_3097 (I56453,I56057,I56012);
and I_3098 (I56471,I56453,I56345);
DFFARX1 I_3099 (I56471,I691,I56399,I56498,);
not I_3100 (I56507,I56012);
DFFARX1 I_3101 (I55868,I691,I56399,I56534,);
not I_3102 (I56543,I56534);
nor I_3103 (I56561,I56543,I56435);
and I_3104 (I56579,I56561,I56012);
nor I_3105 (I56597,I56543,I56507);
nor I_3106 (I56615,I56498,I56597);
DFFARX1 I_3107 (I56381,I691,I56399,I56642,);
nor I_3108 (I56651,I56642,I56498);
not I_3109 (I56669,I56651);
not I_3110 (I56687,I56642);
nor I_3111 (I56705,I56687,I56579);
DFFARX1 I_3112 (I56705,I691,I56399,I56732,);
nand I_3113 (I56741,I55841,I56363);
and I_3114 (I56759,I56741,I56156);
DFFARX1 I_3115 (I56759,I691,I56399,I56786,);
nor I_3116 (I56795,I56786,I56642);
DFFARX1 I_3117 (I56795,I691,I56399,I56822,);
nand I_3118 (I56831,I56786,I56687);
nand I_3119 (I56849,I56669,I56831);
not I_3120 (I56867,I56786);
nor I_3121 (I56885,I56867,I56579);
DFFARX1 I_3122 (I56885,I691,I56399,I56912,);
nor I_3123 (I56921,I56219,I56363);
or I_3124 (I56939,I56642,I56921);
nor I_3125 (I56957,I56786,I56921);
or I_3126 (I56975,I56498,I56921);
DFFARX1 I_3127 (I56921,I691,I56399,I57002,);
not I_3128 (I57011,I698);
DFFARX1 I_3129 (I56957,I691,I57011,I57038,);
DFFARX1 I_3130 (I57038,I691,I57011,I57056,);
not I_3131 (I57065,I57056);
not I_3132 (I57083,I57038);
nand I_3133 (I57101,I57002,I56615);
and I_3134 (I57119,I57101,I56957);
DFFARX1 I_3135 (I57119,I691,I57011,I57146,);
not I_3136 (I57155,I57146);
DFFARX1 I_3137 (I56849,I691,I57011,I57182,);
and I_3138 (I57191,I57182,I56975);
nand I_3139 (I57209,I57182,I56975);
nand I_3140 (I57227,I57155,I57209);
DFFARX1 I_3141 (I56822,I691,I57011,I57254,);
nor I_3142 (I57263,I57254,I57191);
DFFARX1 I_3143 (I57263,I691,I57011,I57290,);
nor I_3144 (I57299,I57254,I57146);
nand I_3145 (I57317,I56822,I56939);
and I_3146 (I57335,I57317,I56912);
DFFARX1 I_3147 (I57335,I691,I57011,I57362,);
nor I_3148 (I57371,I57362,I57254);
not I_3149 (I57389,I57362);
nor I_3150 (I57407,I57389,I57155);
nor I_3151 (I57425,I57083,I57407);
DFFARX1 I_3152 (I57425,I691,I57011,I57452,);
nor I_3153 (I57461,I57389,I57254);
nor I_3154 (I57479,I56732,I56939);
nor I_3155 (I57497,I57479,I57461);
not I_3156 (I57515,I57479);
nand I_3157 (I57533,I57209,I57515);
DFFARX1 I_3158 (I57479,I691,I57011,I57560,);
DFFARX1 I_3159 (I57479,I691,I57011,I57578,);
not I_3160 (I57587,I698);
DFFARX1 I_3161 (I57452,I691,I57587,I57614,);
not I_3162 (I57623,I57614);
nand I_3163 (I57641,I57533,I57371);
and I_3164 (I57659,I57641,I57560);
DFFARX1 I_3165 (I57659,I691,I57587,I57686,);
DFFARX1 I_3166 (I57227,I691,I57587,I57704,);
and I_3167 (I57713,I57704,I57290);
nor I_3168 (I57731,I57686,I57713);
DFFARX1 I_3169 (I57731,I691,I57587,I57758,);
nand I_3170 (I57767,I57704,I57290);
nand I_3171 (I57785,I57623,I57767);
not I_3172 (I57803,I57785);
DFFARX1 I_3173 (I57290,I691,I57587,I57830,);
DFFARX1 I_3174 (I57830,I691,I57587,I57848,);
nand I_3175 (I57857,I57065,I57497);
and I_3176 (I57875,I57857,I57299);
DFFARX1 I_3177 (I57875,I691,I57587,I57902,);
DFFARX1 I_3178 (I57902,I691,I57587,I57920,);
not I_3179 (I57929,I57920);
not I_3180 (I57947,I57902);
nand I_3181 (I57965,I57947,I57767);
nor I_3182 (I57983,I57578,I57497);
not I_3183 (I58001,I57983);
nor I_3184 (I58019,I57947,I58001);
nor I_3185 (I58037,I57623,I58019);
DFFARX1 I_3186 (I58037,I691,I57587,I58064,);
nor I_3187 (I58073,I57686,I58001);
nor I_3188 (I58091,I57902,I58073);
nor I_3189 (I58109,I57830,I57983);
nor I_3190 (I58127,I57686,I57983);
not I_3191 (I58145,I698);
DFFARX1 I_3192 (I58127,I691,I58145,I58172,);
nand I_3193 (I58181,I58109,I57929);
and I_3194 (I58199,I58181,I58127);
DFFARX1 I_3195 (I58199,I691,I58145,I58226,);
nor I_3196 (I58235,I58226,I58172);
not I_3197 (I58253,I58226);
DFFARX1 I_3198 (I58064,I691,I58145,I58280,);
nand I_3199 (I58289,I58280,I58091);
not I_3200 (I58307,I58289);
DFFARX1 I_3201 (I58307,I691,I58145,I58334,);
not I_3202 (I58343,I58334);
nor I_3203 (I58361,I58172,I58289);
nor I_3204 (I58379,I58226,I58361);
DFFARX1 I_3205 (I57965,I691,I58145,I58406,);
DFFARX1 I_3206 (I58406,I691,I58145,I58424,);
not I_3207 (I58433,I58424);
not I_3208 (I58451,I58406);
nand I_3209 (I58469,I58451,I58253);
nand I_3210 (I58487,I57758,I57758);
and I_3211 (I58505,I58487,I57803);
DFFARX1 I_3212 (I58505,I691,I58145,I58532,);
nor I_3213 (I58541,I58532,I58172);
DFFARX1 I_3214 (I58541,I691,I58145,I58568,);
DFFARX1 I_3215 (I58532,I691,I58145,I58586,);
nor I_3216 (I58595,I57848,I57758);
not I_3217 (I58613,I58595);
nor I_3218 (I58631,I58433,I58613);
nand I_3219 (I58649,I58451,I58613);
nor I_3220 (I58667,I58172,I58595);
DFFARX1 I_3221 (I58595,I691,I58145,I58694,);
not I_3222 (I58703,I698);
DFFARX1 I_3223 (I58343,I691,I58703,I58730,);
DFFARX1 I_3224 (I58730,I691,I58703,I58748,);
not I_3225 (I58757,I58748);
nand I_3226 (I58775,I58694,I58586);
and I_3227 (I58793,I58775,I58469);
DFFARX1 I_3228 (I58793,I691,I58703,I58820,);
DFFARX1 I_3229 (I58820,I691,I58703,I58838,);
DFFARX1 I_3230 (I58820,I691,I58703,I58856,);
DFFARX1 I_3231 (I58568,I691,I58703,I58874,);
nand I_3232 (I58883,I58874,I58379);
not I_3233 (I58901,I58883);
nor I_3234 (I58919,I58730,I58901);
DFFARX1 I_3235 (I58649,I691,I58703,I58946,);
not I_3236 (I58955,I58946);
nor I_3237 (I58973,I58955,I58757);
nand I_3238 (I58991,I58955,I58883);
nand I_3239 (I59009,I58235,I58631);
and I_3240 (I59027,I59009,I58568);
DFFARX1 I_3241 (I59027,I691,I58703,I59054,);
nor I_3242 (I59063,I59054,I58730);
DFFARX1 I_3243 (I59063,I691,I58703,I59090,);
not I_3244 (I59099,I59054);
nor I_3245 (I59117,I58667,I58631);
not I_3246 (I59135,I59117);
nor I_3247 (I59153,I58883,I59135);
nor I_3248 (I59171,I59099,I59153);
DFFARX1 I_3249 (I59171,I691,I58703,I59198,);
nor I_3250 (I59207,I59054,I59135);
nor I_3251 (I59225,I58901,I59207);
nor I_3252 (I59243,I59054,I59117);
not I_3253 (I59261,I698);
DFFARX1 I_3254 (I58856,I691,I59261,I59288,);
DFFARX1 I_3255 (I59288,I691,I59261,I59306,);
not I_3256 (I59315,I59306);
not I_3257 (I59333,I59288);
DFFARX1 I_3258 (I59090,I691,I59261,I59360,);
not I_3259 (I59369,I59360);
and I_3260 (I59387,I59333,I58838);
not I_3261 (I59405,I59243);
nand I_3262 (I59423,I59405,I58838);
not I_3263 (I59441,I58991);
nor I_3264 (I59459,I59441,I58973);
nand I_3265 (I59477,I59459,I59225);
nor I_3266 (I59495,I59477,I59423);
DFFARX1 I_3267 (I59495,I691,I59261,I59522,);
not I_3268 (I59531,I59477);
not I_3269 (I59549,I58973);
nand I_3270 (I59567,I59549,I58838);
nor I_3271 (I59585,I58973,I59243);
nand I_3272 (I59603,I59387,I59585);
nand I_3273 (I59621,I59333,I58973);
nand I_3274 (I59639,I59441,I58919);
DFFARX1 I_3275 (I59639,I691,I59261,I59666,);
DFFARX1 I_3276 (I59639,I691,I59261,I59684,);
not I_3277 (I59693,I58919);
nor I_3278 (I59711,I59693,I59243);
and I_3279 (I59729,I59711,I59090);
or I_3280 (I59747,I59729,I59198);
DFFARX1 I_3281 (I59747,I691,I59261,I59774,);
nand I_3282 (I59783,I59774,I59405);
nor I_3283 (I59801,I59783,I59567);
nor I_3284 (I59819,I59774,I59369);
DFFARX1 I_3285 (I59774,I691,I59261,I59846,);
not I_3286 (I59855,I59846);
nor I_3287 (I59873,I59855,I59531);
not I_3288 (I59891,I698);
DFFARX1 I_3289 (I59522,I691,I59891,I59918,);
and I_3290 (I59927,I59918,I59819);
DFFARX1 I_3291 (I59927,I691,I59891,I59954,);
DFFARX1 I_3292 (I59819,I691,I59891,I59972,);
not I_3293 (I59981,I59873);
not I_3294 (I59999,I59315);
nand I_3295 (I60017,I59999,I59981);
nor I_3296 (I60035,I59972,I60017);
DFFARX1 I_3297 (I60017,I691,I59891,I60062,);
not I_3298 (I60071,I60062);
not I_3299 (I60089,I59603);
nand I_3300 (I60107,I59999,I60089);
DFFARX1 I_3301 (I60107,I691,I59891,I60134,);
not I_3302 (I60143,I60134);
not I_3303 (I60161,I59801);
nand I_3304 (I60179,I60161,I59621);
and I_3305 (I60197,I59981,I60179);
nor I_3306 (I60215,I60107,I60197);
DFFARX1 I_3307 (I60215,I691,I59891,I60242,);
DFFARX1 I_3308 (I60197,I691,I59891,I60260,);
nor I_3309 (I60269,I59801,I59522);
nor I_3310 (I60287,I60107,I60269);
or I_3311 (I60305,I59801,I59522);
nor I_3312 (I60323,I59684,I59666);
DFFARX1 I_3313 (I60323,I691,I59891,I60350,);
not I_3314 (I60359,I60350);
nor I_3315 (I60377,I60359,I60143);
nand I_3316 (I60395,I60359,I59972);
not I_3317 (I60413,I59684);
nand I_3318 (I60431,I60413,I60089);
nand I_3319 (I60449,I60359,I60431);
nand I_3320 (I60467,I60449,I60395);
nand I_3321 (I60485,I60431,I60305);
not I_3322 (I60503,I698);
DFFARX1 I_3323 (I60377,I691,I60503,I60530,);
DFFARX1 I_3324 (I60530,I691,I60503,I60548,);
not I_3325 (I60557,I60548);
DFFARX1 I_3326 (I60242,I691,I60503,I60584,);
not I_3327 (I60593,I60485);
nor I_3328 (I60611,I60530,I60593);
not I_3329 (I60629,I60260);
not I_3330 (I60647,I60287);
nand I_3331 (I60665,I60647,I60260);
nor I_3332 (I60683,I60593,I60665);
nor I_3333 (I60701,I60584,I60683);
DFFARX1 I_3334 (I60647,I691,I60503,I60728,);
nor I_3335 (I60737,I60287,I60071);
nand I_3336 (I60755,I60737,I60035);
nor I_3337 (I60773,I60755,I60629);
nand I_3338 (I60791,I60773,I60485);
DFFARX1 I_3339 (I60755,I691,I60503,I60818,);
nand I_3340 (I60827,I60629,I60287);
nor I_3341 (I60845,I60629,I60287);
nand I_3342 (I60863,I60611,I60845);
not I_3343 (I60881,I60467);
nor I_3344 (I60899,I60881,I60827);
DFFARX1 I_3345 (I60899,I691,I60503,I60926,);
nor I_3346 (I60935,I60881,I59954);
and I_3347 (I60953,I60935,I60242);
or I_3348 (I60971,I60953,I60035);
DFFARX1 I_3349 (I60971,I691,I60503,I60998,);
nor I_3350 (I61007,I60998,I60584);
nor I_3351 (I61025,I60530,I61007);
not I_3352 (I61043,I60998);
nor I_3353 (I61061,I61043,I60701);
DFFARX1 I_3354 (I61061,I691,I60503,I61088,);
nand I_3355 (I61097,I61043,I60629);
nor I_3356 (I61115,I60881,I61097);
not I_3357 (I61133,I698);
DFFARX1 I_3358 (I61115,I691,I61133,I61160,);
DFFARX1 I_3359 (I61088,I691,I61133,I61178,);
not I_3360 (I61187,I61178);
not I_3361 (I61205,I60926);
nor I_3362 (I61223,I61205,I60818);
not I_3363 (I61241,I60557);
nor I_3364 (I61259,I61223,I60791);
nor I_3365 (I61277,I61178,I61259);
DFFARX1 I_3366 (I61277,I691,I61133,I61304,);
nor I_3367 (I61313,I60791,I60818);
nand I_3368 (I61331,I61313,I60926);
DFFARX1 I_3369 (I61331,I691,I61133,I61358,);
nor I_3370 (I61367,I61241,I60791);
nand I_3371 (I61385,I61367,I61025);
nor I_3372 (I61403,I61160,I61385);
DFFARX1 I_3373 (I61403,I691,I61133,I61430,);
not I_3374 (I61439,I61385);
nand I_3375 (I61457,I61178,I61439);
DFFARX1 I_3376 (I61385,I691,I61133,I61484,);
not I_3377 (I61493,I61484);
not I_3378 (I61511,I60791);
not I_3379 (I61529,I60863);
nor I_3380 (I61547,I61529,I60557);
nor I_3381 (I61565,I61493,I61547);
nor I_3382 (I61583,I61529,I60728);
and I_3383 (I61601,I61583,I60926);
or I_3384 (I61619,I61601,I61115);
DFFARX1 I_3385 (I61619,I691,I61133,I61646,);
nor I_3386 (I61655,I61646,I61160);
not I_3387 (I61673,I61646);
and I_3388 (I61691,I61673,I61160);
nor I_3389 (I61709,I61187,I61691);
nand I_3390 (I61727,I61673,I61241);
nor I_3391 (I61745,I61529,I61727);
nand I_3392 (I61763,I61673,I61439);
nand I_3393 (I61781,I61241,I60863);
nor I_3394 (I61799,I61511,I61781);
not I_3395 (I61817,I698);
DFFARX1 I_3396 (I61763,I691,I61817,I61844,);
not I_3397 (I61853,I61844);
DFFARX1 I_3398 (I61745,I691,I61817,I61880,);
not I_3399 (I61889,I61430);
nand I_3400 (I61907,I61889,I61565);
not I_3401 (I61925,I61907);
nor I_3402 (I61943,I61925,I61655);
nor I_3403 (I61961,I61853,I61943);
DFFARX1 I_3404 (I61961,I691,I61817,I61988,);
not I_3405 (I61997,I61655);
nand I_3406 (I62015,I61997,I61925);
and I_3407 (I62033,I61997,I61304);
nand I_3408 (I62051,I62033,I61457);
nor I_3409 (I62069,I62051,I61997);
and I_3410 (I62087,I61880,I62051);
not I_3411 (I62105,I62051);
nand I_3412 (I62123,I61880,I62105);
nor I_3413 (I62141,I61844,I62051);
not I_3414 (I62159,I61709);
nor I_3415 (I62177,I62159,I61304);
nand I_3416 (I62195,I62177,I61997);
nor I_3417 (I62213,I61907,I62195);
nor I_3418 (I62231,I62159,I61358);
and I_3419 (I62249,I62231,I61799);
or I_3420 (I62267,I62249,I61430);
DFFARX1 I_3421 (I62267,I691,I61817,I62294,);
nor I_3422 (I62303,I62294,I62015);
DFFARX1 I_3423 (I62303,I691,I61817,I62330,);
DFFARX1 I_3424 (I62294,I691,I61817,I62348,);
not I_3425 (I62357,I62294);
nor I_3426 (I62375,I62357,I61880);
nor I_3427 (I62393,I62177,I62375);
DFFARX1 I_3428 (I62393,I691,I61817,I62420,);
not I_3429 (I62429,I698);
DFFARX1 I_3430 (I62069,I691,I62429,I62456,);
and I_3431 (I62465,I62456,I62141);
DFFARX1 I_3432 (I62465,I691,I62429,I62492,);
DFFARX1 I_3433 (I61988,I691,I62429,I62510,);
not I_3434 (I62519,I62123);
not I_3435 (I62537,I62330);
nand I_3436 (I62555,I62537,I62519);
nor I_3437 (I62573,I62510,I62555);
DFFARX1 I_3438 (I62555,I691,I62429,I62600,);
not I_3439 (I62609,I62600);
not I_3440 (I62627,I62087);
nand I_3441 (I62645,I62537,I62627);
DFFARX1 I_3442 (I62645,I691,I62429,I62672,);
not I_3443 (I62681,I62672);
not I_3444 (I62699,I62420);
nand I_3445 (I62717,I62699,I62348);
and I_3446 (I62735,I62519,I62717);
nor I_3447 (I62753,I62645,I62735);
DFFARX1 I_3448 (I62753,I691,I62429,I62780,);
DFFARX1 I_3449 (I62735,I691,I62429,I62798,);
nor I_3450 (I62807,I62420,I62330);
nor I_3451 (I62825,I62645,I62807);
or I_3452 (I62843,I62420,I62330);
nor I_3453 (I62861,I62213,I62141);
DFFARX1 I_3454 (I62861,I691,I62429,I62888,);
not I_3455 (I62897,I62888);
nor I_3456 (I62915,I62897,I62681);
nand I_3457 (I62933,I62897,I62510);
not I_3458 (I62951,I62213);
nand I_3459 (I62969,I62951,I62627);
nand I_3460 (I62987,I62897,I62969);
nand I_3461 (I63005,I62987,I62933);
nand I_3462 (I63023,I62969,I62843);
not I_3463 (I63041,I698);
DFFARX1 I_3464 (I62915,I691,I63041,I63068,);
not I_3465 (I63077,I63068);
nand I_3466 (I63095,I62780,I62780);
and I_3467 (I63113,I63095,I63023);
DFFARX1 I_3468 (I63113,I691,I63041,I63140,);
DFFARX1 I_3469 (I63140,I691,I63041,I63158,);
DFFARX1 I_3470 (I62573,I691,I63041,I63176,);
nand I_3471 (I63185,I63176,I62825);
not I_3472 (I63203,I63185);
DFFARX1 I_3473 (I63203,I691,I63041,I63230,);
not I_3474 (I63239,I63230);
nor I_3475 (I63257,I63077,I63239);
DFFARX1 I_3476 (I62609,I691,I63041,I63284,);
nor I_3477 (I63293,I63284,I63140);
nor I_3478 (I63311,I63284,I63203);
nand I_3479 (I63329,I62492,I63005);
and I_3480 (I63347,I63329,I62573);
DFFARX1 I_3481 (I63347,I691,I63041,I63374,);
not I_3482 (I63383,I63374);
nand I_3483 (I63401,I63383,I63284);
nand I_3484 (I63419,I63383,I63185);
nor I_3485 (I63437,I62798,I63005);
and I_3486 (I63455,I63284,I63437);
nor I_3487 (I63473,I63383,I63455);
DFFARX1 I_3488 (I63473,I691,I63041,I63500,);
nor I_3489 (I63509,I63068,I63437);
DFFARX1 I_3490 (I63509,I691,I63041,I63536,);
nor I_3491 (I63545,I63374,I63437);
not I_3492 (I63563,I63545);
nand I_3493 (I63581,I63563,I63401);
not I_3494 (I63599,I698);
DFFARX1 I_3495 (I63311,I691,I63599,I63626,);
and I_3496 (I63635,I63626,I63581);
DFFARX1 I_3497 (I63635,I691,I63599,I63662,);
DFFARX1 I_3498 (I63500,I691,I63599,I63680,);
not I_3499 (I63689,I63536);
not I_3500 (I63707,I63536);
nand I_3501 (I63725,I63707,I63689);
nor I_3502 (I63743,I63680,I63725);
DFFARX1 I_3503 (I63725,I691,I63599,I63770,);
not I_3504 (I63779,I63770);
not I_3505 (I63797,I63158);
nand I_3506 (I63815,I63707,I63797);
DFFARX1 I_3507 (I63815,I691,I63599,I63842,);
not I_3508 (I63851,I63842);
not I_3509 (I63869,I63293);
nand I_3510 (I63887,I63869,I63311);
and I_3511 (I63905,I63689,I63887);
nor I_3512 (I63923,I63815,I63905);
DFFARX1 I_3513 (I63923,I691,I63599,I63950,);
DFFARX1 I_3514 (I63905,I691,I63599,I63968,);
nor I_3515 (I63977,I63293,I63257);
nor I_3516 (I63995,I63815,I63977);
or I_3517 (I64013,I63293,I63257);
nor I_3518 (I64031,I63419,I63419);
DFFARX1 I_3519 (I64031,I691,I63599,I64058,);
not I_3520 (I64067,I64058);
nor I_3521 (I64085,I64067,I63851);
nand I_3522 (I64103,I64067,I63680);
not I_3523 (I64121,I63419);
nand I_3524 (I64139,I64121,I63797);
nand I_3525 (I64157,I64067,I64139);
nand I_3526 (I64175,I64157,I64103);
nand I_3527 (I64193,I64139,I64013);
not I_3528 (I64211,I698);
DFFARX1 I_3529 (I64193,I691,I64211,I64238,);
not I_3530 (I64247,I64238);
nand I_3531 (I64265,I63968,I63950);
and I_3532 (I64283,I64265,I63743);
DFFARX1 I_3533 (I64283,I691,I64211,I64310,);
DFFARX1 I_3534 (I63779,I691,I64211,I64328,);
and I_3535 (I64337,I64328,I63743);
nor I_3536 (I64355,I64310,I64337);
DFFARX1 I_3537 (I64355,I691,I64211,I64382,);
nand I_3538 (I64391,I64328,I63743);
nand I_3539 (I64409,I64247,I64391);
not I_3540 (I64427,I64409);
DFFARX1 I_3541 (I63950,I691,I64211,I64454,);
DFFARX1 I_3542 (I64454,I691,I64211,I64472,);
nand I_3543 (I64481,I63995,I64175);
and I_3544 (I64499,I64481,I63662);
DFFARX1 I_3545 (I64499,I691,I64211,I64526,);
DFFARX1 I_3546 (I64526,I691,I64211,I64544,);
not I_3547 (I64553,I64544);
not I_3548 (I64571,I64526);
nand I_3549 (I64589,I64571,I64391);
nor I_3550 (I64607,I64085,I64175);
not I_3551 (I64625,I64607);
nor I_3552 (I64643,I64571,I64625);
nor I_3553 (I64661,I64247,I64643);
DFFARX1 I_3554 (I64661,I691,I64211,I64688,);
nor I_3555 (I64697,I64310,I64625);
nor I_3556 (I64715,I64526,I64697);
nor I_3557 (I64733,I64454,I64607);
nor I_3558 (I64751,I64310,I64607);
not I_3559 (I64769,I698);
DFFARX1 I_3560 (I64751,I691,I64769,I64796,);
not I_3561 (I64805,I64796);
nand I_3562 (I64823,I64427,I64472);
and I_3563 (I64841,I64823,I64382);
DFFARX1 I_3564 (I64841,I691,I64769,I64868,);
not I_3565 (I64877,I64751);
DFFARX1 I_3566 (I64688,I691,I64769,I64904,);
not I_3567 (I64913,I64904);
nor I_3568 (I64931,I64913,I64805);
and I_3569 (I64949,I64931,I64751);
nor I_3570 (I64967,I64913,I64877);
nor I_3571 (I64985,I64868,I64967);
DFFARX1 I_3572 (I64589,I691,I64769,I65012,);
nor I_3573 (I65021,I65012,I64868);
not I_3574 (I65039,I65021);
not I_3575 (I65057,I65012);
nor I_3576 (I65075,I65057,I64949);
DFFARX1 I_3577 (I65075,I691,I64769,I65102,);
nand I_3578 (I65111,I64553,I64382);
and I_3579 (I65129,I65111,I64715);
DFFARX1 I_3580 (I65129,I691,I64769,I65156,);
nor I_3581 (I65165,I65156,I65012);
DFFARX1 I_3582 (I65165,I691,I64769,I65192,);
nand I_3583 (I65201,I65156,I65057);
nand I_3584 (I65219,I65039,I65201);
not I_3585 (I65237,I65156);
nor I_3586 (I65255,I65237,I64949);
DFFARX1 I_3587 (I65255,I691,I64769,I65282,);
nor I_3588 (I65291,I64733,I64382);
or I_3589 (I65309,I65012,I65291);
nor I_3590 (I65327,I65156,I65291);
or I_3591 (I65345,I64868,I65291);
DFFARX1 I_3592 (I65291,I691,I64769,I65372,);
not I_3593 (I65381,I698);
DFFARX1 I_3594 (I65345,I691,I65381,I65408,);
DFFARX1 I_3595 (I65192,I691,I65381,I65426,);
not I_3596 (I65435,I65426);
not I_3597 (I65453,I64985);
nor I_3598 (I65471,I65453,I65192);
not I_3599 (I65489,I65219);
nor I_3600 (I65507,I65471,I65102);
nor I_3601 (I65525,I65426,I65507);
DFFARX1 I_3602 (I65525,I691,I65381,I65552,);
nor I_3603 (I65561,I65102,I65192);
nand I_3604 (I65579,I65561,I64985);
DFFARX1 I_3605 (I65579,I691,I65381,I65606,);
nor I_3606 (I65615,I65489,I65102);
nand I_3607 (I65633,I65615,I65327);
nor I_3608 (I65651,I65408,I65633);
DFFARX1 I_3609 (I65651,I691,I65381,I65678,);
not I_3610 (I65687,I65633);
nand I_3611 (I65705,I65426,I65687);
DFFARX1 I_3612 (I65633,I691,I65381,I65732,);
not I_3613 (I65741,I65732);
not I_3614 (I65759,I65102);
not I_3615 (I65777,I65309);
nor I_3616 (I65795,I65777,I65219);
nor I_3617 (I65813,I65741,I65795);
nor I_3618 (I65831,I65777,I65282);
and I_3619 (I65849,I65831,I65372);
or I_3620 (I65867,I65849,I65327);
DFFARX1 I_3621 (I65867,I691,I65381,I65894,);
nor I_3622 (I65903,I65894,I65408);
not I_3623 (I65921,I65894);
and I_3624 (I65939,I65921,I65408);
nor I_3625 (I65957,I65435,I65939);
nand I_3626 (I65975,I65921,I65489);
nor I_3627 (I65993,I65777,I65975);
nand I_3628 (I66011,I65921,I65687);
nand I_3629 (I66029,I65489,I65309);
nor I_3630 (I66047,I65759,I66029);
not I_3631 (I66065,I698);
DFFARX1 I_3632 (I65957,I691,I66065,I66092,);
not I_3633 (I66101,I66092);
nand I_3634 (I66119,I65813,I65552);
and I_3635 (I66137,I66119,I65678);
DFFARX1 I_3636 (I66137,I691,I66065,I66164,);
DFFARX1 I_3637 (I66047,I691,I66065,I66182,);
and I_3638 (I66191,I66182,I65993);
nor I_3639 (I66209,I66164,I66191);
DFFARX1 I_3640 (I66209,I691,I66065,I66236,);
nand I_3641 (I66245,I66182,I65993);
nand I_3642 (I66263,I66101,I66245);
not I_3643 (I66281,I66263);
DFFARX1 I_3644 (I65903,I691,I66065,I66308,);
DFFARX1 I_3645 (I66308,I691,I66065,I66326,);
nand I_3646 (I66335,I65606,I65705);
and I_3647 (I66353,I66335,I66011);
DFFARX1 I_3648 (I66353,I691,I66065,I66380,);
DFFARX1 I_3649 (I66380,I691,I66065,I66398,);
not I_3650 (I66407,I66398);
not I_3651 (I66425,I66380);
nand I_3652 (I66443,I66425,I66245);
nor I_3653 (I66461,I65678,I65705);
not I_3654 (I66479,I66461);
nor I_3655 (I66497,I66425,I66479);
nor I_3656 (I66515,I66101,I66497);
DFFARX1 I_3657 (I66515,I691,I66065,I66542,);
nor I_3658 (I66551,I66164,I66479);
nor I_3659 (I66569,I66380,I66551);
nor I_3660 (I66587,I66308,I66461);
nor I_3661 (I66605,I66164,I66461);
not I_3662 (I66623,I698);
DFFARX1 I_3663 (I66281,I691,I66623,I66650,);
DFFARX1 I_3664 (I66650,I691,I66623,I66668,);
not I_3665 (I66677,I66668);
not I_3666 (I66695,I66650);
DFFARX1 I_3667 (I66236,I691,I66623,I66722,);
nand I_3668 (I66731,I66722,I66587);
not I_3669 (I66749,I66587);
not I_3670 (I66767,I66605);
nand I_3671 (I66785,I66407,I66542);
and I_3672 (I66803,I66407,I66542);
not I_3673 (I66821,I66569);
nand I_3674 (I66839,I66821,I66767);
nor I_3675 (I66857,I66839,I66731);
nor I_3676 (I66875,I66749,I66839);
nand I_3677 (I66893,I66803,I66875);
not I_3678 (I66911,I66443);
nor I_3679 (I66929,I66911,I66407);
nor I_3680 (I66947,I66929,I66569);
nor I_3681 (I66965,I66695,I66947);
DFFARX1 I_3682 (I66965,I691,I66623,I66992,);
not I_3683 (I67001,I66929);
DFFARX1 I_3684 (I67001,I691,I66623,I67028,);
and I_3685 (I67037,I66722,I66929);
nor I_3686 (I67055,I66911,I66605);
and I_3687 (I67073,I67055,I66236);
or I_3688 (I67091,I67073,I66326);
DFFARX1 I_3689 (I67091,I691,I66623,I67118,);
nor I_3690 (I67127,I67118,I66821);
DFFARX1 I_3691 (I67127,I691,I66623,I67154,);
nand I_3692 (I67163,I67118,I66722);
nand I_3693 (I67181,I66821,I67163);
nor I_3694 (I67199,I67181,I66785);
not I_3695 (I67217,I698);
DFFARX1 I_3696 (I66857,I691,I67217,I67244,);
DFFARX1 I_3697 (I67244,I691,I67217,I67262,);
not I_3698 (I67271,I67262);
not I_3699 (I67289,I67244);
DFFARX1 I_3700 (I67037,I691,I67217,I67316,);
not I_3701 (I67325,I67316);
and I_3702 (I67343,I67289,I66893);
not I_3703 (I67361,I67154);
nand I_3704 (I67379,I67361,I66893);
not I_3705 (I67397,I66992);
nor I_3706 (I67415,I67397,I66857);
nand I_3707 (I67433,I67415,I67199);
nor I_3708 (I67451,I67433,I67379);
DFFARX1 I_3709 (I67451,I691,I67217,I67478,);
not I_3710 (I67487,I67433);
not I_3711 (I67505,I66857);
nand I_3712 (I67523,I67505,I66893);
nor I_3713 (I67541,I66857,I67154);
nand I_3714 (I67559,I67343,I67541);
nand I_3715 (I67577,I67289,I66857);
nand I_3716 (I67595,I67397,I66893);
DFFARX1 I_3717 (I67595,I691,I67217,I67622,);
DFFARX1 I_3718 (I67595,I691,I67217,I67640,);
not I_3719 (I67649,I66893);
nor I_3720 (I67667,I67649,I66677);
and I_3721 (I67685,I67667,I67028);
or I_3722 (I67703,I67685,I67154);
DFFARX1 I_3723 (I67703,I691,I67217,I67730,);
nand I_3724 (I67739,I67730,I67361);
nor I_3725 (I67757,I67739,I67523);
nor I_3726 (I67775,I67730,I67325);
DFFARX1 I_3727 (I67730,I691,I67217,I67802,);
not I_3728 (I67811,I67802);
nor I_3729 (I67829,I67811,I67487);
not I_3730 (I67847,I698);
DFFARX1 I_3731 (I67640,I691,I67847,I67874,);
not I_3732 (I67883,I67874);
DFFARX1 I_3733 (I67478,I691,I67847,I67910,);
not I_3734 (I67919,I67829);
nand I_3735 (I67937,I67919,I67775);
not I_3736 (I67955,I67937);
nor I_3737 (I67973,I67955,I67478);
nor I_3738 (I67991,I67883,I67973);
DFFARX1 I_3739 (I67991,I691,I67847,I68018,);
not I_3740 (I68027,I67478);
nand I_3741 (I68045,I68027,I67955);
and I_3742 (I68063,I68027,I67775);
nand I_3743 (I68081,I68063,I67271);
nor I_3744 (I68099,I68081,I68027);
and I_3745 (I68117,I67910,I68081);
not I_3746 (I68135,I68081);
nand I_3747 (I68153,I67910,I68135);
nor I_3748 (I68171,I67874,I68081);
not I_3749 (I68189,I67559);
nor I_3750 (I68207,I68189,I67775);
nand I_3751 (I68225,I68207,I68027);
nor I_3752 (I68243,I67937,I68225);
nor I_3753 (I68261,I68189,I67577);
and I_3754 (I68279,I68261,I67622);
or I_3755 (I68297,I68279,I67757);
DFFARX1 I_3756 (I68297,I691,I67847,I68324,);
nor I_3757 (I68333,I68324,I68045);
DFFARX1 I_3758 (I68333,I691,I67847,I68360,);
DFFARX1 I_3759 (I68324,I691,I67847,I68378,);
not I_3760 (I68387,I68324);
nor I_3761 (I68405,I68387,I67910);
nor I_3762 (I68423,I68207,I68405);
DFFARX1 I_3763 (I68423,I691,I67847,I68450,);
not I_3764 (I68459,I698);
DFFARX1 I_3765 (I68099,I691,I68459,I68486,);
DFFARX1 I_3766 (I68486,I691,I68459,I68504,);
not I_3767 (I68513,I68504);
not I_3768 (I68531,I68486);
DFFARX1 I_3769 (I68117,I691,I68459,I68558,);
not I_3770 (I68567,I68558);
and I_3771 (I68585,I68531,I68378);
not I_3772 (I68603,I68450);
nand I_3773 (I68621,I68603,I68378);
not I_3774 (I68639,I68360);
nor I_3775 (I68657,I68639,I68171);
nand I_3776 (I68675,I68657,I68243);
nor I_3777 (I68693,I68675,I68621);
DFFARX1 I_3778 (I68693,I691,I68459,I68720,);
not I_3779 (I68729,I68675);
not I_3780 (I68747,I68171);
nand I_3781 (I68765,I68747,I68378);
nor I_3782 (I68783,I68171,I68450);
nand I_3783 (I68801,I68585,I68783);
nand I_3784 (I68819,I68531,I68171);
nand I_3785 (I68837,I68639,I68018);
DFFARX1 I_3786 (I68837,I691,I68459,I68864,);
DFFARX1 I_3787 (I68837,I691,I68459,I68882,);
not I_3788 (I68891,I68018);
nor I_3789 (I68909,I68891,I68360);
and I_3790 (I68927,I68909,I68153);
or I_3791 (I68945,I68927,I68171);
DFFARX1 I_3792 (I68945,I691,I68459,I68972,);
nand I_3793 (I68981,I68972,I68603);
nor I_3794 (I68999,I68981,I68765);
nor I_3795 (I69017,I68972,I68567);
DFFARX1 I_3796 (I68972,I691,I68459,I69044,);
not I_3797 (I69053,I69044);
nor I_3798 (I69071,I69053,I68729);
not I_3799 (I69089,I698);
DFFARX1 I_3800 (I68720,I691,I69089,I69116,);
nand I_3801 (I69125,I68720,I68819);
and I_3802 (I69143,I69125,I68513);
DFFARX1 I_3803 (I69143,I691,I69089,I69170,);
nor I_3804 (I69179,I69170,I69116);
not I_3805 (I69197,I69170);
DFFARX1 I_3806 (I68801,I691,I69089,I69224,);
nand I_3807 (I69233,I69224,I68999);
not I_3808 (I69251,I69233);
DFFARX1 I_3809 (I69251,I691,I69089,I69278,);
not I_3810 (I69287,I69278);
nor I_3811 (I69305,I69116,I69233);
nor I_3812 (I69323,I69170,I69305);
DFFARX1 I_3813 (I69071,I691,I69089,I69350,);
DFFARX1 I_3814 (I69350,I691,I69089,I69368,);
not I_3815 (I69377,I69368);
not I_3816 (I69395,I69350);
nand I_3817 (I69413,I69395,I69197);
nand I_3818 (I69431,I69017,I69017);
and I_3819 (I69449,I69431,I68864);
DFFARX1 I_3820 (I69449,I691,I69089,I69476,);
nor I_3821 (I69485,I69476,I69116);
DFFARX1 I_3822 (I69485,I691,I69089,I69512,);
DFFARX1 I_3823 (I69476,I691,I69089,I69530,);
nor I_3824 (I69539,I68882,I69017);
not I_3825 (I69557,I69539);
nor I_3826 (I69575,I69377,I69557);
nand I_3827 (I69593,I69395,I69557);
nor I_3828 (I69611,I69116,I69539);
DFFARX1 I_3829 (I69539,I691,I69089,I69638,);
not I_3830 (I69647,I698);
DFFARX1 I_3831 (I69287,I691,I69647,I69674,);
and I_3832 (I69683,I69674,I69413);
DFFARX1 I_3833 (I69683,I691,I69647,I69710,);
DFFARX1 I_3834 (I69530,I691,I69647,I69728,);
not I_3835 (I69737,I69512);
not I_3836 (I69755,I69575);
nand I_3837 (I69773,I69755,I69737);
nor I_3838 (I69791,I69728,I69773);
DFFARX1 I_3839 (I69773,I691,I69647,I69818,);
not I_3840 (I69827,I69818);
not I_3841 (I69845,I69638);
nand I_3842 (I69863,I69755,I69845);
DFFARX1 I_3843 (I69863,I691,I69647,I69890,);
not I_3844 (I69899,I69890);
not I_3845 (I69917,I69611);
nand I_3846 (I69935,I69917,I69179);
and I_3847 (I69953,I69737,I69935);
nor I_3848 (I69971,I69863,I69953);
DFFARX1 I_3849 (I69971,I691,I69647,I69998,);
DFFARX1 I_3850 (I69953,I691,I69647,I70016,);
nor I_3851 (I70025,I69611,I69323);
nor I_3852 (I70043,I69863,I70025);
or I_3853 (I70061,I69611,I69323);
nor I_3854 (I70079,I69593,I69512);
DFFARX1 I_3855 (I70079,I691,I69647,I70106,);
not I_3856 (I70115,I70106);
nor I_3857 (I70133,I70115,I69899);
nand I_3858 (I70151,I70115,I69728);
not I_3859 (I70169,I69593);
nand I_3860 (I70187,I70169,I69845);
nand I_3861 (I70205,I70115,I70187);
nand I_3862 (I70223,I70205,I70151);
nand I_3863 (I70241,I70187,I70061);
not I_3864 (I70259,I698);
DFFARX1 I_3865 (I69791,I691,I70259,I70286,);
DFFARX1 I_3866 (I70286,I691,I70259,I70304,);
not I_3867 (I70313,I70304);
not I_3868 (I70331,I70286);
nand I_3869 (I70349,I69710,I69791);
and I_3870 (I70367,I70349,I70241);
DFFARX1 I_3871 (I70367,I691,I70259,I70394,);
not I_3872 (I70403,I70394);
DFFARX1 I_3873 (I69827,I691,I70259,I70430,);
and I_3874 (I70439,I70430,I69998);
nand I_3875 (I70457,I70430,I69998);
nand I_3876 (I70475,I70403,I70457);
DFFARX1 I_3877 (I70133,I691,I70259,I70502,);
nor I_3878 (I70511,I70502,I70439);
DFFARX1 I_3879 (I70511,I691,I70259,I70538,);
nor I_3880 (I70547,I70502,I70394);
nand I_3881 (I70565,I70043,I70223);
and I_3882 (I70583,I70565,I70016);
DFFARX1 I_3883 (I70583,I691,I70259,I70610,);
nor I_3884 (I70619,I70610,I70502);
not I_3885 (I70637,I70610);
nor I_3886 (I70655,I70637,I70403);
nor I_3887 (I70673,I70331,I70655);
DFFARX1 I_3888 (I70673,I691,I70259,I70700,);
nor I_3889 (I70709,I70637,I70502);
nor I_3890 (I70727,I69998,I70223);
nor I_3891 (I70745,I70727,I70709);
not I_3892 (I70763,I70727);
nand I_3893 (I70781,I70457,I70763);
DFFARX1 I_3894 (I70727,I691,I70259,I70808,);
DFFARX1 I_3895 (I70727,I691,I70259,I70826,);
not I_3896 (I70835,I698);
DFFARX1 I_3897 (I70619,I691,I70835,I70862,);
nand I_3898 (I70871,I70862,I70781);
not I_3899 (I70889,I70871);
DFFARX1 I_3900 (I70538,I691,I70835,I70916,);
not I_3901 (I70925,I70916);
not I_3902 (I70943,I70475);
or I_3903 (I70961,I70538,I70475);
nor I_3904 (I70979,I70538,I70475);
or I_3905 (I70997,I70547,I70538);
DFFARX1 I_3906 (I70997,I691,I70835,I71024,);
not I_3907 (I71033,I70745);
nand I_3908 (I71051,I71033,I70826);
nand I_3909 (I71069,I70943,I71051);
and I_3910 (I71087,I70925,I71069);
nor I_3911 (I71105,I70745,I70313);
and I_3912 (I71123,I70925,I71105);
nor I_3913 (I71141,I70889,I71123);
DFFARX1 I_3914 (I71105,I691,I70835,I71168,);
not I_3915 (I71177,I71168);
nor I_3916 (I71195,I70925,I71177);
or I_3917 (I71213,I70997,I70700);
nor I_3918 (I71231,I70700,I70547);
nand I_3919 (I71249,I71069,I71231);
nand I_3920 (I71267,I71213,I71249);
DFFARX1 I_3921 (I71267,I691,I70835,I71294,);
nor I_3922 (I71303,I71231,I70961);
DFFARX1 I_3923 (I71303,I691,I70835,I71330,);
nor I_3924 (I71339,I70700,I70808);
DFFARX1 I_3925 (I71339,I691,I70835,I71366,);
DFFARX1 I_3926 (I71366,I691,I70835,I71384,);
not I_3927 (I71393,I71366);
nand I_3928 (I71411,I71393,I70871);
nand I_3929 (I71429,I71393,I70979);
not I_3930 (I71447,I698);
DFFARX1 I_3931 (I156,I691,I71447,I71474,);
DFFARX1 I_3932 (I71474,I691,I71447,I71492,);
not I_3933 (I71501,I71492);
not I_3934 (I71519,I71474);
DFFARX1 I_3935 (I252,I691,I71447,I71546,);
not I_3936 (I71555,I71546);
and I_3937 (I71573,I71519,I580);
not I_3938 (I71591,I268);
nand I_3939 (I71609,I71591,I580);
not I_3940 (I71627,I84);
nor I_3941 (I71645,I71627,I540);
nand I_3942 (I71663,I71645,I316);
nor I_3943 (I71681,I71663,I71609);
DFFARX1 I_3944 (I71681,I691,I71447,I71708,);
not I_3945 (I71717,I71663);
not I_3946 (I71735,I540);
nand I_3947 (I71753,I71735,I580);
nor I_3948 (I71771,I540,I268);
nand I_3949 (I71789,I71573,I71771);
nand I_3950 (I71807,I71519,I540);
nand I_3951 (I71825,I71627,I460);
DFFARX1 I_3952 (I71825,I691,I71447,I71852,);
DFFARX1 I_3953 (I71825,I691,I71447,I71870,);
not I_3954 (I71879,I460);
nor I_3955 (I71897,I71879,I212);
and I_3956 (I71915,I71897,I652);
or I_3957 (I71933,I71915,I596);
DFFARX1 I_3958 (I71933,I691,I71447,I71960,);
nand I_3959 (I71969,I71960,I71591);
nor I_3960 (I71987,I71969,I71753);
nor I_3961 (I72005,I71960,I71555);
DFFARX1 I_3962 (I71960,I691,I71447,I72032,);
not I_3963 (I72041,I72032);
nor I_3964 (I72059,I72041,I71717);
not I_3965 (I72077,I698);
DFFARX1 I_3966 (I71708,I691,I72077,I72104,);
and I_3967 (I72113,I72104,I72005);
DFFARX1 I_3968 (I72113,I691,I72077,I72140,);
DFFARX1 I_3969 (I72005,I691,I72077,I72158,);
not I_3970 (I72167,I72059);
not I_3971 (I72185,I71501);
nand I_3972 (I72203,I72185,I72167);
nor I_3973 (I72221,I72158,I72203);
DFFARX1 I_3974 (I72203,I691,I72077,I72248,);
not I_3975 (I72257,I72248);
not I_3976 (I72275,I71789);
nand I_3977 (I72293,I72185,I72275);
DFFARX1 I_3978 (I72293,I691,I72077,I72320,);
not I_3979 (I72329,I72320);
not I_3980 (I72347,I71987);
nand I_3981 (I72365,I72347,I71807);
and I_3982 (I72383,I72167,I72365);
nor I_3983 (I72401,I72293,I72383);
DFFARX1 I_3984 (I72401,I691,I72077,I72428,);
DFFARX1 I_3985 (I72383,I691,I72077,I72446,);
nor I_3986 (I72455,I71987,I71708);
nor I_3987 (I72473,I72293,I72455);
or I_3988 (I72491,I71987,I71708);
nor I_3989 (I72509,I71870,I71852);
DFFARX1 I_3990 (I72509,I691,I72077,I72536,);
not I_3991 (I72545,I72536);
nor I_3992 (I72563,I72545,I72329);
nand I_3993 (I72581,I72545,I72158);
not I_3994 (I72599,I71870);
nand I_3995 (I72617,I72599,I72275);
nand I_3996 (I72635,I72545,I72617);
nand I_3997 (I72653,I72635,I72581);
nand I_3998 (I72671,I72617,I72491);
not I_3999 (I72689,I698);
DFFARX1 I_4000 (I72671,I691,I72689,I72716,);
not I_4001 (I72725,I72716);
nand I_4002 (I72743,I72446,I72428);
and I_4003 (I72761,I72743,I72221);
DFFARX1 I_4004 (I72761,I691,I72689,I72788,);
DFFARX1 I_4005 (I72257,I691,I72689,I72806,);
and I_4006 (I72815,I72806,I72221);
nor I_4007 (I72833,I72788,I72815);
DFFARX1 I_4008 (I72833,I691,I72689,I72860,);
nand I_4009 (I72869,I72806,I72221);
nand I_4010 (I72887,I72725,I72869);
not I_4011 (I72905,I72887);
DFFARX1 I_4012 (I72428,I691,I72689,I72932,);
DFFARX1 I_4013 (I72932,I691,I72689,I72950,);
nand I_4014 (I72959,I72473,I72653);
and I_4015 (I72977,I72959,I72140);
DFFARX1 I_4016 (I72977,I691,I72689,I73004,);
DFFARX1 I_4017 (I73004,I691,I72689,I73022,);
not I_4018 (I73031,I73022);
not I_4019 (I73049,I73004);
nand I_4020 (I73067,I73049,I72869);
nor I_4021 (I73085,I72563,I72653);
not I_4022 (I73103,I73085);
nor I_4023 (I73121,I73049,I73103);
nor I_4024 (I73139,I72725,I73121);
DFFARX1 I_4025 (I73139,I691,I72689,I73166,);
nor I_4026 (I73175,I72788,I73103);
nor I_4027 (I73193,I73004,I73175);
nor I_4028 (I73211,I72932,I73085);
nor I_4029 (I73229,I72788,I73085);
not I_4030 (I73247,I698);
DFFARX1 I_4031 (I73067,I691,I73247,I73274,);
DFFARX1 I_4032 (I73274,I691,I73247,I73292,);
not I_4033 (I73301,I73292);
not I_4034 (I73319,I73274);
DFFARX1 I_4035 (I73229,I691,I73247,I73346,);
not I_4036 (I73355,I73346);
and I_4037 (I73373,I73319,I72860);
not I_4038 (I73391,I72950);
nand I_4039 (I73409,I73391,I72860);
not I_4040 (I73427,I73211);
nor I_4041 (I73445,I73427,I73193);
nand I_4042 (I73463,I73445,I72905);
nor I_4043 (I73481,I73463,I73409);
DFFARX1 I_4044 (I73481,I691,I73247,I73508,);
not I_4045 (I73517,I73463);
not I_4046 (I73535,I73193);
nand I_4047 (I73553,I73535,I72860);
nor I_4048 (I73571,I73193,I72950);
nand I_4049 (I73589,I73373,I73571);
nand I_4050 (I73607,I73319,I73193);
nand I_4051 (I73625,I73427,I72860);
DFFARX1 I_4052 (I73625,I691,I73247,I73652,);
DFFARX1 I_4053 (I73625,I691,I73247,I73670,);
not I_4054 (I73679,I72860);
nor I_4055 (I73697,I73679,I73166);
and I_4056 (I73715,I73697,I73031);
or I_4057 (I73733,I73715,I73229);
DFFARX1 I_4058 (I73733,I691,I73247,I73760,);
nand I_4059 (I73769,I73760,I73391);
nor I_4060 (I73787,I73769,I73553);
nor I_4061 (I73805,I73760,I73355);
DFFARX1 I_4062 (I73760,I691,I73247,I73832,);
not I_4063 (I73841,I73832);
nor I_4064 (I73859,I73841,I73517);
not I_4065 (I73877,I698);
DFFARX1 I_4066 (I73607,I691,I73877,I73904,);
not I_4067 (I73913,I73904);
nand I_4068 (I73931,I73805,I73652);
and I_4069 (I73949,I73931,I73589);
DFFARX1 I_4070 (I73949,I691,I73877,I73976,);
DFFARX1 I_4071 (I73976,I691,I73877,I73994,);
DFFARX1 I_4072 (I73859,I691,I73877,I74012,);
nand I_4073 (I74021,I74012,I73670);
not I_4074 (I74039,I74021);
DFFARX1 I_4075 (I74039,I691,I73877,I74066,);
not I_4076 (I74075,I74066);
nor I_4077 (I74093,I73913,I74075);
DFFARX1 I_4078 (I73787,I691,I73877,I74120,);
nor I_4079 (I74129,I74120,I73976);
nor I_4080 (I74147,I74120,I74039);
nand I_4081 (I74165,I73508,I73301);
and I_4082 (I74183,I74165,I73805);
DFFARX1 I_4083 (I74183,I691,I73877,I74210,);
not I_4084 (I74219,I74210);
nand I_4085 (I74237,I74219,I74120);
nand I_4086 (I74255,I74219,I74021);
nor I_4087 (I74273,I73508,I73301);
and I_4088 (I74291,I74120,I74273);
nor I_4089 (I74309,I74219,I74291);
DFFARX1 I_4090 (I74309,I691,I73877,I74336,);
nor I_4091 (I74345,I73904,I74273);
DFFARX1 I_4092 (I74345,I691,I73877,I74372,);
nor I_4093 (I74381,I74210,I74273);
not I_4094 (I74399,I74381);
nand I_4095 (I74417,I74399,I74237);
not I_4096 (I74435,I698);
DFFARX1 I_4097 (I74147,I691,I74435,I74462,);
and I_4098 (I74471,I74462,I74417);
DFFARX1 I_4099 (I74471,I691,I74435,I74498,);
DFFARX1 I_4100 (I74336,I691,I74435,I74516,);
not I_4101 (I74525,I74372);
not I_4102 (I74543,I74372);
nand I_4103 (I74561,I74543,I74525);
nor I_4104 (I74579,I74516,I74561);
DFFARX1 I_4105 (I74561,I691,I74435,I74606,);
not I_4106 (I74615,I74606);
not I_4107 (I74633,I73994);
nand I_4108 (I74651,I74543,I74633);
DFFARX1 I_4109 (I74651,I691,I74435,I74678,);
not I_4110 (I74687,I74678);
not I_4111 (I74705,I74129);
nand I_4112 (I74723,I74705,I74147);
and I_4113 (I74741,I74525,I74723);
nor I_4114 (I74759,I74651,I74741);
DFFARX1 I_4115 (I74759,I691,I74435,I74786,);
DFFARX1 I_4116 (I74741,I691,I74435,I74804,);
nor I_4117 (I74813,I74129,I74093);
nor I_4118 (I74831,I74651,I74813);
or I_4119 (I74849,I74129,I74093);
nor I_4120 (I74867,I74255,I74255);
DFFARX1 I_4121 (I74867,I691,I74435,I74894,);
not I_4122 (I74903,I74894);
nor I_4123 (I74921,I74903,I74687);
nand I_4124 (I74939,I74903,I74516);
not I_4125 (I74957,I74255);
nand I_4126 (I74975,I74957,I74633);
nand I_4127 (I74993,I74903,I74975);
nand I_4128 (I75011,I74993,I74939);
nand I_4129 (I75029,I74975,I74849);
not I_4130 (I75047,I698);
DFFARX1 I_4131 (I74786,I691,I75047,I75074,);
nand I_4132 (I75083,I74498,I74786);
and I_4133 (I75101,I75083,I74921);
DFFARX1 I_4134 (I75101,I691,I75047,I75128,);
nor I_4135 (I75137,I75128,I75074);
not I_4136 (I75155,I75128);
DFFARX1 I_4137 (I74615,I691,I75047,I75182,);
nand I_4138 (I75191,I75182,I75029);
not I_4139 (I75209,I75191);
DFFARX1 I_4140 (I75209,I691,I75047,I75236,);
not I_4141 (I75245,I75236);
nor I_4142 (I75263,I75074,I75191);
nor I_4143 (I75281,I75128,I75263);
DFFARX1 I_4144 (I74579,I691,I75047,I75308,);
DFFARX1 I_4145 (I75308,I691,I75047,I75326,);
not I_4146 (I75335,I75326);
not I_4147 (I75353,I75308);
nand I_4148 (I75371,I75353,I75155);
nand I_4149 (I75389,I74579,I75011);
and I_4150 (I75407,I75389,I74804);
DFFARX1 I_4151 (I75407,I691,I75047,I75434,);
nor I_4152 (I75443,I75434,I75074);
DFFARX1 I_4153 (I75443,I691,I75047,I75470,);
DFFARX1 I_4154 (I75434,I691,I75047,I75488,);
nor I_4155 (I75497,I74831,I75011);
not I_4156 (I75515,I75497);
nor I_4157 (I75533,I75335,I75515);
nand I_4158 (I75551,I75353,I75515);
nor I_4159 (I75569,I75074,I75497);
DFFARX1 I_4160 (I75497,I691,I75047,I75596,);
not I_4161 (I75605,I698);
DFFARX1 I_4162 (I75551,I691,I75605,I75632,);
nand I_4163 (I75641,I75632,I75245);
not I_4164 (I75659,I75641);
DFFARX1 I_4165 (I75533,I691,I75605,I75686,);
not I_4166 (I75695,I75686);
not I_4167 (I75713,I75281);
or I_4168 (I75731,I75596,I75281);
nor I_4169 (I75749,I75596,I75281);
or I_4170 (I75767,I75569,I75596);
DFFARX1 I_4171 (I75767,I691,I75605,I75794,);
not I_4172 (I75803,I75137);
nand I_4173 (I75821,I75803,I75470);
nand I_4174 (I75839,I75713,I75821);
and I_4175 (I75857,I75695,I75839);
nor I_4176 (I75875,I75137,I75371);
and I_4177 (I75893,I75695,I75875);
nor I_4178 (I75911,I75659,I75893);
DFFARX1 I_4179 (I75875,I691,I75605,I75938,);
not I_4180 (I75947,I75938);
nor I_4181 (I75965,I75695,I75947);
or I_4182 (I75983,I75767,I75488);
nor I_4183 (I76001,I75488,I75569);
nand I_4184 (I76019,I75839,I76001);
nand I_4185 (I76037,I75983,I76019);
DFFARX1 I_4186 (I76037,I691,I75605,I76064,);
nor I_4187 (I76073,I76001,I75731);
DFFARX1 I_4188 (I76073,I691,I75605,I76100,);
nor I_4189 (I76109,I75488,I75470);
DFFARX1 I_4190 (I76109,I691,I75605,I76136,);
DFFARX1 I_4191 (I76136,I691,I75605,I76154,);
not I_4192 (I76163,I76136);
nand I_4193 (I76181,I76163,I75641);
nand I_4194 (I76199,I76163,I75749);
not I_4195 (I76217,I698);
DFFARX1 I_4196 (I76154,I691,I76217,I76244,);
nand I_4197 (I76253,I76181,I75857);
and I_4198 (I76271,I76253,I76100);
DFFARX1 I_4199 (I76271,I691,I76217,I76298,);
nor I_4200 (I76307,I76298,I76244);
not I_4201 (I76325,I76298);
DFFARX1 I_4202 (I75911,I691,I76217,I76352,);
nand I_4203 (I76361,I76352,I75965);
not I_4204 (I76379,I76361);
DFFARX1 I_4205 (I76379,I691,I76217,I76406,);
not I_4206 (I76415,I76406);
nor I_4207 (I76433,I76244,I76361);
nor I_4208 (I76451,I76298,I76433);
DFFARX1 I_4209 (I76064,I691,I76217,I76478,);
DFFARX1 I_4210 (I76478,I691,I76217,I76496,);
not I_4211 (I76505,I76496);
not I_4212 (I76523,I76478);
nand I_4213 (I76541,I76523,I76325);
nand I_4214 (I76559,I76100,I76199);
and I_4215 (I76577,I76559,I75794);
DFFARX1 I_4216 (I76577,I691,I76217,I76604,);
nor I_4217 (I76613,I76604,I76244);
DFFARX1 I_4218 (I76613,I691,I76217,I76640,);
DFFARX1 I_4219 (I76604,I691,I76217,I76658,);
nor I_4220 (I76667,I75857,I76199);
not I_4221 (I76685,I76667);
nor I_4222 (I76703,I76505,I76685);
nand I_4223 (I76721,I76523,I76685);
nor I_4224 (I76739,I76244,I76667);
DFFARX1 I_4225 (I76667,I691,I76217,I76766,);
not I_4226 (I76775,I698);
DFFARX1 I_4227 (I76451,I691,I76775,I76802,);
not I_4228 (I76811,I76802);
nand I_4229 (I76829,I76640,I76640);
and I_4230 (I76847,I76829,I76658);
DFFARX1 I_4231 (I76847,I691,I76775,I76874,);
DFFARX1 I_4232 (I76874,I691,I76775,I76892,);
DFFARX1 I_4233 (I76703,I691,I76775,I76910,);
nand I_4234 (I76919,I76910,I76307);
not I_4235 (I76937,I76919);
DFFARX1 I_4236 (I76937,I691,I76775,I76964,);
not I_4237 (I76973,I76964);
nor I_4238 (I76991,I76811,I76973);
DFFARX1 I_4239 (I76739,I691,I76775,I77018,);
nor I_4240 (I77027,I77018,I76874);
nor I_4241 (I77045,I77018,I76937);
nand I_4242 (I77063,I76415,I76721);
and I_4243 (I77081,I77063,I76541);
DFFARX1 I_4244 (I77081,I691,I76775,I77108,);
not I_4245 (I77117,I77108);
nand I_4246 (I77135,I77117,I77018);
nand I_4247 (I77153,I77117,I76919);
nor I_4248 (I77171,I76766,I76721);
and I_4249 (I77189,I77018,I77171);
nor I_4250 (I77207,I77117,I77189);
DFFARX1 I_4251 (I77207,I691,I76775,I77234,);
nor I_4252 (I77243,I76802,I77171);
DFFARX1 I_4253 (I77243,I691,I76775,I77270,);
nor I_4254 (I77279,I77108,I77171);
not I_4255 (I77297,I77279);
nand I_4256 (I77315,I77297,I77135);
not I_4257 (I77333,I698);
DFFARX1 I_4258 (I77153,I691,I77333,I77360,);
DFFARX1 I_4259 (I77360,I691,I77333,I77378,);
not I_4260 (I77387,I77378);
not I_4261 (I77405,I77360);
DFFARX1 I_4262 (I77270,I691,I77333,I77432,);
not I_4263 (I77441,I77432);
and I_4264 (I77459,I77405,I76892);
not I_4265 (I77477,I77153);
nand I_4266 (I77495,I77477,I76892);
not I_4267 (I77513,I77270);
nor I_4268 (I77531,I77513,I77027);
nand I_4269 (I77549,I77531,I77045);
nor I_4270 (I77567,I77549,I77495);
DFFARX1 I_4271 (I77567,I691,I77333,I77594,);
not I_4272 (I77603,I77549);
not I_4273 (I77621,I77027);
nand I_4274 (I77639,I77621,I76892);
nor I_4275 (I77657,I77027,I77153);
nand I_4276 (I77675,I77459,I77657);
nand I_4277 (I77693,I77405,I77027);
nand I_4278 (I77711,I77513,I77234);
DFFARX1 I_4279 (I77711,I691,I77333,I77738,);
DFFARX1 I_4280 (I77711,I691,I77333,I77756,);
not I_4281 (I77765,I77234);
nor I_4282 (I77783,I77765,I76991);
and I_4283 (I77801,I77783,I77045);
or I_4284 (I77819,I77801,I77315);
DFFARX1 I_4285 (I77819,I691,I77333,I77846,);
nand I_4286 (I77855,I77846,I77477);
nor I_4287 (I77873,I77855,I77639);
nor I_4288 (I77891,I77846,I77441);
DFFARX1 I_4289 (I77846,I691,I77333,I77918,);
not I_4290 (I77927,I77918);
nor I_4291 (I77945,I77927,I77603);
not I_4292 (I77963,I698);
DFFARX1 I_4293 (I77594,I691,I77963,I77990,);
DFFARX1 I_4294 (I77990,I691,I77963,I78008,);
not I_4295 (I78017,I78008);
DFFARX1 I_4296 (I77387,I691,I77963,I78044,);
not I_4297 (I78053,I77945);
nor I_4298 (I78071,I77990,I78053);
not I_4299 (I78089,I77675);
not I_4300 (I78107,I77873);
nand I_4301 (I78125,I78107,I77675);
nor I_4302 (I78143,I78053,I78125);
nor I_4303 (I78161,I78044,I78143);
DFFARX1 I_4304 (I78107,I691,I77963,I78188,);
nor I_4305 (I78197,I77873,I77891);
nand I_4306 (I78215,I78197,I77738);
nor I_4307 (I78233,I78215,I78089);
nand I_4308 (I78251,I78233,I77945);
DFFARX1 I_4309 (I78215,I691,I77963,I78278,);
nand I_4310 (I78287,I78089,I77873);
nor I_4311 (I78305,I78089,I77873);
nand I_4312 (I78323,I78071,I78305);
not I_4313 (I78341,I77756);
nor I_4314 (I78359,I78341,I78287);
DFFARX1 I_4315 (I78359,I691,I77963,I78386,);
nor I_4316 (I78395,I78341,I77594);
and I_4317 (I78413,I78395,I77693);
or I_4318 (I78431,I78413,I77891);
DFFARX1 I_4319 (I78431,I691,I77963,I78458,);
nor I_4320 (I78467,I78458,I78044);
nor I_4321 (I78485,I77990,I78467);
not I_4322 (I78503,I78458);
nor I_4323 (I78521,I78503,I78161);
DFFARX1 I_4324 (I78521,I691,I77963,I78548,);
nand I_4325 (I78557,I78503,I78089);
nor I_4326 (I78575,I78341,I78557);
not I_4327 (I78593,I698);
DFFARX1 I_4328 (I78323,I691,I78593,I78620,);
DFFARX1 I_4329 (I78620,I691,I78593,I78638,);
not I_4330 (I78647,I78638);
not I_4331 (I78665,I78620);
DFFARX1 I_4332 (I78251,I691,I78593,I78692,);
not I_4333 (I78701,I78692);
and I_4334 (I78719,I78665,I78188);
not I_4335 (I78737,I78278);
nand I_4336 (I78755,I78737,I78188);
not I_4337 (I78773,I78485);
nor I_4338 (I78791,I78773,I78386);
nand I_4339 (I78809,I78791,I78575);
nor I_4340 (I78827,I78809,I78755);
DFFARX1 I_4341 (I78827,I691,I78593,I78854,);
not I_4342 (I78863,I78809);
not I_4343 (I78881,I78386);
nand I_4344 (I78899,I78881,I78188);
nor I_4345 (I78917,I78386,I78278);
nand I_4346 (I78935,I78719,I78917);
nand I_4347 (I78953,I78665,I78386);
nand I_4348 (I78971,I78773,I78017);
DFFARX1 I_4349 (I78971,I691,I78593,I78998,);
DFFARX1 I_4350 (I78971,I691,I78593,I79016,);
not I_4351 (I79025,I78017);
nor I_4352 (I79043,I79025,I78548);
and I_4353 (I79061,I79043,I78386);
or I_4354 (I79079,I79061,I78575);
DFFARX1 I_4355 (I79079,I691,I78593,I79106,);
nand I_4356 (I79115,I79106,I78737);
nor I_4357 (I79133,I79115,I78899);
nor I_4358 (I79151,I79106,I78701);
DFFARX1 I_4359 (I79106,I691,I78593,I79178,);
not I_4360 (I79187,I79178);
nor I_4361 (I79205,I79187,I78863);
not I_4362 (I79223,I698);
DFFARX1 I_4363 (I79016,I691,I79223,I79250,);
not I_4364 (I79259,I79250);
DFFARX1 I_4365 (I78854,I691,I79223,I79286,);
not I_4366 (I79295,I79205);
nand I_4367 (I79313,I79295,I79151);
not I_4368 (I79331,I79313);
nor I_4369 (I79349,I79331,I78854);
nor I_4370 (I79367,I79259,I79349);
DFFARX1 I_4371 (I79367,I691,I79223,I79394,);
not I_4372 (I79403,I78854);
nand I_4373 (I79421,I79403,I79331);
and I_4374 (I79439,I79403,I79151);
nand I_4375 (I79457,I79439,I78647);
nor I_4376 (I79475,I79457,I79403);
and I_4377 (I79493,I79286,I79457);
not I_4378 (I79511,I79457);
nand I_4379 (I79529,I79286,I79511);
nor I_4380 (I79547,I79250,I79457);
not I_4381 (I79565,I78935);
nor I_4382 (I79583,I79565,I79151);
nand I_4383 (I79601,I79583,I79403);
nor I_4384 (I79619,I79313,I79601);
nor I_4385 (I79637,I79565,I78953);
and I_4386 (I79655,I79637,I78998);
or I_4387 (I79673,I79655,I79133);
DFFARX1 I_4388 (I79673,I691,I79223,I79700,);
nor I_4389 (I79709,I79700,I79421);
DFFARX1 I_4390 (I79709,I691,I79223,I79736,);
DFFARX1 I_4391 (I79700,I691,I79223,I79754,);
not I_4392 (I79763,I79700);
nor I_4393 (I79781,I79763,I79286);
nor I_4394 (I79799,I79583,I79781);
DFFARX1 I_4395 (I79799,I691,I79223,I79826,);
not I_4396 (I79835,I698);
DFFARX1 I_4397 (I79736,I691,I79835,I79862,);
not I_4398 (I79871,I79862);
nand I_4399 (I79889,I79529,I79394);
and I_4400 (I79907,I79889,I79754);
DFFARX1 I_4401 (I79907,I691,I79835,I79934,);
not I_4402 (I79943,I79826);
DFFARX1 I_4403 (I79493,I691,I79835,I79970,);
not I_4404 (I79979,I79970);
nor I_4405 (I79997,I79979,I79871);
and I_4406 (I80015,I79997,I79826);
nor I_4407 (I80033,I79979,I79943);
nor I_4408 (I80051,I79934,I80033);
DFFARX1 I_4409 (I79475,I691,I79835,I80078,);
nor I_4410 (I80087,I80078,I79934);
not I_4411 (I80105,I80087);
not I_4412 (I80123,I80078);
nor I_4413 (I80141,I80123,I80015);
DFFARX1 I_4414 (I80141,I691,I79835,I80168,);
nand I_4415 (I80177,I79619,I79547);
and I_4416 (I80195,I80177,I79736);
DFFARX1 I_4417 (I80195,I691,I79835,I80222,);
nor I_4418 (I80231,I80222,I80078);
DFFARX1 I_4419 (I80231,I691,I79835,I80258,);
nand I_4420 (I80267,I80222,I80123);
nand I_4421 (I80285,I80105,I80267);
not I_4422 (I80303,I80222);
nor I_4423 (I80321,I80303,I80015);
DFFARX1 I_4424 (I80321,I691,I79835,I80348,);
nor I_4425 (I80357,I79547,I79547);
or I_4426 (I80375,I80078,I80357);
nor I_4427 (I80393,I80222,I80357);
or I_4428 (I80411,I79934,I80357);
DFFARX1 I_4429 (I80357,I691,I79835,I80438,);
not I_4430 (I80447,I698);
DFFARX1 I_4431 (I80375,I691,I80447,I80474,);
nand I_4432 (I80483,I80393,I80168);
and I_4433 (I80501,I80483,I80438);
DFFARX1 I_4434 (I80501,I691,I80447,I80528,);
nor I_4435 (I80537,I80528,I80474);
not I_4436 (I80555,I80528);
DFFARX1 I_4437 (I80285,I691,I80447,I80582,);
nand I_4438 (I80591,I80582,I80393);
not I_4439 (I80609,I80591);
DFFARX1 I_4440 (I80609,I691,I80447,I80636,);
not I_4441 (I80645,I80636);
nor I_4442 (I80663,I80474,I80591);
nor I_4443 (I80681,I80528,I80663);
DFFARX1 I_4444 (I80411,I691,I80447,I80708,);
DFFARX1 I_4445 (I80708,I691,I80447,I80726,);
not I_4446 (I80735,I80726);
not I_4447 (I80753,I80708);
nand I_4448 (I80771,I80753,I80555);
nand I_4449 (I80789,I80258,I80051);
and I_4450 (I80807,I80789,I80258);
DFFARX1 I_4451 (I80807,I691,I80447,I80834,);
nor I_4452 (I80843,I80834,I80474);
DFFARX1 I_4453 (I80843,I691,I80447,I80870,);
DFFARX1 I_4454 (I80834,I691,I80447,I80888,);
nor I_4455 (I80897,I80348,I80051);
not I_4456 (I80915,I80897);
nor I_4457 (I80933,I80735,I80915);
nand I_4458 (I80951,I80753,I80915);
nor I_4459 (I80969,I80474,I80897);
DFFARX1 I_4460 (I80897,I691,I80447,I80996,);
not I_4461 (I81005,I698);
DFFARX1 I_4462 (I80645,I691,I81005,I81032,);
not I_4463 (I81041,I81032);
nand I_4464 (I81059,I80681,I80996);
and I_4465 (I81077,I81059,I80870);
DFFARX1 I_4466 (I81077,I691,I81005,I81104,);
DFFARX1 I_4467 (I80537,I691,I81005,I81122,);
and I_4468 (I81131,I81122,I80888);
nor I_4469 (I81149,I81104,I81131);
DFFARX1 I_4470 (I81149,I691,I81005,I81176,);
nand I_4471 (I81185,I81122,I80888);
nand I_4472 (I81203,I81041,I81185);
not I_4473 (I81221,I81203);
DFFARX1 I_4474 (I80933,I691,I81005,I81248,);
DFFARX1 I_4475 (I81248,I691,I81005,I81266,);
nand I_4476 (I81275,I80870,I80771);
and I_4477 (I81293,I81275,I80951);
DFFARX1 I_4478 (I81293,I691,I81005,I81320,);
DFFARX1 I_4479 (I81320,I691,I81005,I81338,);
not I_4480 (I81347,I81338);
not I_4481 (I81365,I81320);
nand I_4482 (I81383,I81365,I81185);
nor I_4483 (I81401,I80969,I80771);
not I_4484 (I81419,I81401);
nor I_4485 (I81437,I81365,I81419);
nor I_4486 (I81455,I81041,I81437);
DFFARX1 I_4487 (I81455,I691,I81005,I81482,);
nor I_4488 (I81491,I81104,I81419);
nor I_4489 (I81509,I81320,I81491);
nor I_4490 (I81527,I81248,I81401);
nor I_4491 (I81545,I81104,I81401);
not I_4492 (I81563,I698);
DFFARX1 I_4493 (I81509,I691,I81563,I81590,);
DFFARX1 I_4494 (I81590,I691,I81563,I81608,);
not I_4495 (I81617,I81608);
not I_4496 (I81635,I81590);
nand I_4497 (I81653,I81266,I81176);
and I_4498 (I81671,I81653,I81545);
DFFARX1 I_4499 (I81671,I691,I81563,I81698,);
not I_4500 (I81707,I81698);
DFFARX1 I_4501 (I81383,I691,I81563,I81734,);
and I_4502 (I81743,I81734,I81545);
nand I_4503 (I81761,I81734,I81545);
nand I_4504 (I81779,I81707,I81761);
DFFARX1 I_4505 (I81482,I691,I81563,I81806,);
nor I_4506 (I81815,I81806,I81743);
DFFARX1 I_4507 (I81815,I691,I81563,I81842,);
nor I_4508 (I81851,I81806,I81698);
nand I_4509 (I81869,I81176,I81527);
and I_4510 (I81887,I81869,I81221);
DFFARX1 I_4511 (I81887,I691,I81563,I81914,);
nor I_4512 (I81923,I81914,I81806);
not I_4513 (I81941,I81914);
nor I_4514 (I81959,I81941,I81707);
nor I_4515 (I81977,I81635,I81959);
DFFARX1 I_4516 (I81977,I691,I81563,I82004,);
nor I_4517 (I82013,I81941,I81806);
nor I_4518 (I82031,I81347,I81527);
nor I_4519 (I82049,I82031,I82013);
not I_4520 (I82067,I82031);
nand I_4521 (I82085,I81761,I82067);
DFFARX1 I_4522 (I82031,I691,I81563,I82112,);
DFFARX1 I_4523 (I82031,I691,I81563,I82130,);
not I_4524 (I82139,I698);
DFFARX1 I_4525 (I82049,I691,I82139,I82166,);
not I_4526 (I82175,I82166);
nand I_4527 (I82193,I81842,I82004);
and I_4528 (I82211,I82193,I82130);
DFFARX1 I_4529 (I82211,I691,I82139,I82238,);
not I_4530 (I82247,I81851);
DFFARX1 I_4531 (I81923,I691,I82139,I82274,);
not I_4532 (I82283,I82274);
nor I_4533 (I82301,I82283,I82175);
and I_4534 (I82319,I82301,I81851);
nor I_4535 (I82337,I82283,I82247);
nor I_4536 (I82355,I82238,I82337);
DFFARX1 I_4537 (I82085,I691,I82139,I82382,);
nor I_4538 (I82391,I82382,I82238);
not I_4539 (I82409,I82391);
not I_4540 (I82427,I82382);
nor I_4541 (I82445,I82427,I82319);
DFFARX1 I_4542 (I82445,I691,I82139,I82472,);
nand I_4543 (I82481,I81617,I82112);
and I_4544 (I82499,I82481,I81779);
DFFARX1 I_4545 (I82499,I691,I82139,I82526,);
nor I_4546 (I82535,I82526,I82382);
DFFARX1 I_4547 (I82535,I691,I82139,I82562,);
nand I_4548 (I82571,I82526,I82427);
nand I_4549 (I82589,I82409,I82571);
not I_4550 (I82607,I82526);
nor I_4551 (I82625,I82607,I82319);
DFFARX1 I_4552 (I82625,I691,I82139,I82652,);
nor I_4553 (I82661,I81842,I82112);
or I_4554 (I82679,I82382,I82661);
nor I_4555 (I82697,I82526,I82661);
or I_4556 (I82715,I82238,I82661);
DFFARX1 I_4557 (I82661,I691,I82139,I82742,);
not I_4558 (I82751,I698);
DFFARX1 I_4559 (I82355,I691,I82751,I82778,);
and I_4560 (I82787,I82778,I82697);
DFFARX1 I_4561 (I82787,I691,I82751,I82814,);
DFFARX1 I_4562 (I82715,I691,I82751,I82832,);
not I_4563 (I82841,I82562);
not I_4564 (I82859,I82742);
nand I_4565 (I82877,I82859,I82841);
nor I_4566 (I82895,I82832,I82877);
DFFARX1 I_4567 (I82877,I691,I82751,I82922,);
not I_4568 (I82931,I82922);
not I_4569 (I82949,I82679);
nand I_4570 (I82967,I82859,I82949);
DFFARX1 I_4571 (I82967,I691,I82751,I82994,);
not I_4572 (I83003,I82994);
not I_4573 (I83021,I82652);
nand I_4574 (I83039,I83021,I82472);
and I_4575 (I83057,I82841,I83039);
nor I_4576 (I83075,I82967,I83057);
DFFARX1 I_4577 (I83075,I691,I82751,I83102,);
DFFARX1 I_4578 (I83057,I691,I82751,I83120,);
nor I_4579 (I83129,I82652,I82589);
nor I_4580 (I83147,I82967,I83129);
or I_4581 (I83165,I82652,I82589);
nor I_4582 (I83183,I82562,I82697);
DFFARX1 I_4583 (I83183,I691,I82751,I83210,);
not I_4584 (I83219,I83210);
nor I_4585 (I83237,I83219,I83003);
nand I_4586 (I83255,I83219,I82832);
not I_4587 (I83273,I82562);
nand I_4588 (I83291,I83273,I82949);
nand I_4589 (I83309,I83219,I83291);
nand I_4590 (I83327,I83309,I83255);
nand I_4591 (I83345,I83291,I83165);
not I_4592 (I83363,I698);
DFFARX1 I_4593 (I83102,I691,I83363,I83390,);
nand I_4594 (I83399,I82814,I83102);
and I_4595 (I83417,I83399,I83237);
DFFARX1 I_4596 (I83417,I691,I83363,I83444,);
nor I_4597 (I83453,I83444,I83390);
not I_4598 (I83471,I83444);
DFFARX1 I_4599 (I82931,I691,I83363,I83498,);
nand I_4600 (I83507,I83498,I83345);
not I_4601 (I83525,I83507);
DFFARX1 I_4602 (I83525,I691,I83363,I83552,);
not I_4603 (I83561,I83552);
nor I_4604 (I83579,I83390,I83507);
nor I_4605 (I83597,I83444,I83579);
DFFARX1 I_4606 (I82895,I691,I83363,I83624,);
DFFARX1 I_4607 (I83624,I691,I83363,I83642,);
not I_4608 (I83651,I83642);
not I_4609 (I83669,I83624);
nand I_4610 (I83687,I83669,I83471);
nand I_4611 (I83705,I82895,I83327);
and I_4612 (I83723,I83705,I83120);
DFFARX1 I_4613 (I83723,I691,I83363,I83750,);
nor I_4614 (I83759,I83750,I83390);
DFFARX1 I_4615 (I83759,I691,I83363,I83786,);
DFFARX1 I_4616 (I83750,I691,I83363,I83804,);
nor I_4617 (I83813,I83147,I83327);
not I_4618 (I83831,I83813);
nor I_4619 (I83849,I83651,I83831);
nand I_4620 (I83867,I83669,I83831);
nor I_4621 (I83885,I83390,I83813);
DFFARX1 I_4622 (I83813,I691,I83363,I83912,);
not I_4623 (I83921,I698);
DFFARX1 I_4624 (I83687,I691,I83921,I83948,);
nand I_4625 (I83957,I83948,I83885);
DFFARX1 I_4626 (I83597,I691,I83921,I83984,);
DFFARX1 I_4627 (I83984,I691,I83921,I84002,);
not I_4628 (I84011,I84002);
not I_4629 (I84029,I83804);
nor I_4630 (I84047,I83804,I83453);
not I_4631 (I84065,I83561);
nand I_4632 (I84083,I84029,I84065);
nor I_4633 (I84101,I83561,I83804);
and I_4634 (I84119,I84101,I83957);
not I_4635 (I84137,I83867);
nand I_4636 (I84155,I84137,I83912);
nor I_4637 (I84173,I83867,I83786);
not I_4638 (I84191,I84173);
nand I_4639 (I84209,I84047,I84191);
DFFARX1 I_4640 (I84173,I691,I83921,I84236,);
nor I_4641 (I84245,I83849,I83561);
nor I_4642 (I84263,I84245,I83453);
and I_4643 (I84281,I84263,I84155);
DFFARX1 I_4644 (I84281,I691,I83921,I84308,);
nor I_4645 (I84317,I84245,I84083);
or I_4646 (I84335,I84173,I84245);
nor I_4647 (I84353,I83849,I83786);
DFFARX1 I_4648 (I84353,I691,I83921,I84380,);
not I_4649 (I84389,I84380);
nand I_4650 (I84407,I84389,I84029);
nor I_4651 (I84425,I84407,I83453);
DFFARX1 I_4652 (I84425,I691,I83921,I84452,);
nor I_4653 (I84461,I84389,I84083);
nor I_4654 (I84479,I84245,I84461);
not I_4655 (I84497,I698);
DFFARX1 I_4656 (I84308,I691,I84497,I84524,);
DFFARX1 I_4657 (I84524,I691,I84497,I84542,);
not I_4658 (I84551,I84542);
not I_4659 (I84569,I84524);
DFFARX1 I_4660 (I84119,I691,I84497,I84596,);
not I_4661 (I84605,I84596);
and I_4662 (I84623,I84569,I84236);
not I_4663 (I84641,I84119);
nand I_4664 (I84659,I84641,I84236);
not I_4665 (I84677,I84011);
nor I_4666 (I84695,I84677,I84317);
nand I_4667 (I84713,I84695,I84335);
nor I_4668 (I84731,I84713,I84659);
DFFARX1 I_4669 (I84731,I691,I84497,I84758,);
not I_4670 (I84767,I84713);
not I_4671 (I84785,I84317);
nand I_4672 (I84803,I84785,I84236);
nor I_4673 (I84821,I84317,I84119);
nand I_4674 (I84839,I84623,I84821);
nand I_4675 (I84857,I84569,I84317);
nand I_4676 (I84875,I84677,I84479);
DFFARX1 I_4677 (I84875,I691,I84497,I84902,);
DFFARX1 I_4678 (I84875,I691,I84497,I84920,);
not I_4679 (I84929,I84479);
nor I_4680 (I84947,I84929,I84452);
and I_4681 (I84965,I84947,I84209);
or I_4682 (I84983,I84965,I84452);
DFFARX1 I_4683 (I84983,I691,I84497,I85010,);
nand I_4684 (I85019,I85010,I84641);
nor I_4685 (I85037,I85019,I84803);
nor I_4686 (I85055,I85010,I84605);
DFFARX1 I_4687 (I85010,I691,I84497,I85082,);
not I_4688 (I85091,I85082);
nor I_4689 (I85109,I85091,I84767);
not I_4690 (I85127,I698);
DFFARX1 I_4691 (I84758,I691,I85127,I85154,);
and I_4692 (I85163,I85154,I85055);
DFFARX1 I_4693 (I85163,I691,I85127,I85190,);
DFFARX1 I_4694 (I85055,I691,I85127,I85208,);
not I_4695 (I85217,I85109);
not I_4696 (I85235,I84551);
nand I_4697 (I85253,I85235,I85217);
nor I_4698 (I85271,I85208,I85253);
DFFARX1 I_4699 (I85253,I691,I85127,I85298,);
not I_4700 (I85307,I85298);
not I_4701 (I85325,I84839);
nand I_4702 (I85343,I85235,I85325);
DFFARX1 I_4703 (I85343,I691,I85127,I85370,);
not I_4704 (I85379,I85370);
not I_4705 (I85397,I85037);
nand I_4706 (I85415,I85397,I84857);
and I_4707 (I85433,I85217,I85415);
nor I_4708 (I85451,I85343,I85433);
DFFARX1 I_4709 (I85451,I691,I85127,I85478,);
DFFARX1 I_4710 (I85433,I691,I85127,I85496,);
nor I_4711 (I85505,I85037,I84758);
nor I_4712 (I85523,I85343,I85505);
or I_4713 (I85541,I85037,I84758);
nor I_4714 (I85559,I84920,I84902);
DFFARX1 I_4715 (I85559,I691,I85127,I85586,);
not I_4716 (I85595,I85586);
nor I_4717 (I85613,I85595,I85379);
nand I_4718 (I85631,I85595,I85208);
not I_4719 (I85649,I84920);
nand I_4720 (I85667,I85649,I85325);
nand I_4721 (I85685,I85595,I85667);
nand I_4722 (I85703,I85685,I85631);
nand I_4723 (I85721,I85667,I85541);
not I_4724 (I85739,I698);
DFFARX1 I_4725 (I85613,I691,I85739,I85766,);
not I_4726 (I85775,I85766);
nand I_4727 (I85793,I85478,I85523);
and I_4728 (I85811,I85793,I85190);
DFFARX1 I_4729 (I85811,I691,I85739,I85838,);
not I_4730 (I85847,I85703);
DFFARX1 I_4731 (I85721,I691,I85739,I85874,);
not I_4732 (I85883,I85874);
nor I_4733 (I85901,I85883,I85775);
and I_4734 (I85919,I85901,I85703);
nor I_4735 (I85937,I85883,I85847);
nor I_4736 (I85955,I85838,I85937);
DFFARX1 I_4737 (I85307,I691,I85739,I85982,);
nor I_4738 (I85991,I85982,I85838);
not I_4739 (I86009,I85991);
not I_4740 (I86027,I85982);
nor I_4741 (I86045,I86027,I85919);
DFFARX1 I_4742 (I86045,I691,I85739,I86072,);
nand I_4743 (I86081,I85271,I85271);
and I_4744 (I86099,I86081,I85478);
DFFARX1 I_4745 (I86099,I691,I85739,I86126,);
nor I_4746 (I86135,I86126,I85982);
DFFARX1 I_4747 (I86135,I691,I85739,I86162,);
nand I_4748 (I86171,I86126,I86027);
nand I_4749 (I86189,I86009,I86171);
not I_4750 (I86207,I86126);
nor I_4751 (I86225,I86207,I85919);
DFFARX1 I_4752 (I86225,I691,I85739,I86252,);
nor I_4753 (I86261,I85496,I85271);
or I_4754 (I86279,I85982,I86261);
nor I_4755 (I86297,I86126,I86261);
or I_4756 (I86315,I85838,I86261);
DFFARX1 I_4757 (I86261,I691,I85739,I86342,);
not I_4758 (I86351,I698);
DFFARX1 I_4759 (I86162,I691,I86351,I86378,);
not I_4760 (I86387,I86378);
nand I_4761 (I86405,I86297,I86162);
and I_4762 (I86423,I86405,I86279);
DFFARX1 I_4763 (I86423,I691,I86351,I86450,);
DFFARX1 I_4764 (I86450,I691,I86351,I86468,);
DFFARX1 I_4765 (I86189,I691,I86351,I86486,);
nand I_4766 (I86495,I86486,I85955);
not I_4767 (I86513,I86495);
DFFARX1 I_4768 (I86513,I691,I86351,I86540,);
not I_4769 (I86549,I86540);
nor I_4770 (I86567,I86387,I86549);
DFFARX1 I_4771 (I86342,I691,I86351,I86594,);
nor I_4772 (I86603,I86594,I86450);
nor I_4773 (I86621,I86594,I86513);
nand I_4774 (I86639,I86072,I86315);
and I_4775 (I86657,I86639,I86297);
DFFARX1 I_4776 (I86657,I691,I86351,I86684,);
not I_4777 (I86693,I86684);
nand I_4778 (I86711,I86693,I86594);
nand I_4779 (I86729,I86693,I86495);
nor I_4780 (I86747,I86252,I86315);
and I_4781 (I86765,I86594,I86747);
nor I_4782 (I86783,I86693,I86765);
DFFARX1 I_4783 (I86783,I691,I86351,I86810,);
nor I_4784 (I86819,I86378,I86747);
DFFARX1 I_4785 (I86819,I691,I86351,I86846,);
nor I_4786 (I86855,I86684,I86747);
not I_4787 (I86873,I86855);
nand I_4788 (I86891,I86873,I86711);
not I_4789 (I86909,I698);
DFFARX1 I_4790 (I86729,I691,I86909,I86936,);
DFFARX1 I_4791 (I86936,I691,I86909,I86954,);
not I_4792 (I86963,I86954);
not I_4793 (I86981,I86936);
DFFARX1 I_4794 (I86846,I691,I86909,I87008,);
not I_4795 (I87017,I87008);
and I_4796 (I87035,I86981,I86468);
not I_4797 (I87053,I86729);
nand I_4798 (I87071,I87053,I86468);
not I_4799 (I87089,I86846);
nor I_4800 (I87107,I87089,I86603);
nand I_4801 (I87125,I87107,I86621);
nor I_4802 (I87143,I87125,I87071);
DFFARX1 I_4803 (I87143,I691,I86909,I87170,);
not I_4804 (I87179,I87125);
not I_4805 (I87197,I86603);
nand I_4806 (I87215,I87197,I86468);
nor I_4807 (I87233,I86603,I86729);
nand I_4808 (I87251,I87035,I87233);
nand I_4809 (I87269,I86981,I86603);
nand I_4810 (I87287,I87089,I86810);
DFFARX1 I_4811 (I87287,I691,I86909,I87314,);
DFFARX1 I_4812 (I87287,I691,I86909,I87332,);
not I_4813 (I87341,I86810);
nor I_4814 (I87359,I87341,I86567);
and I_4815 (I87377,I87359,I86621);
or I_4816 (I87395,I87377,I86891);
DFFARX1 I_4817 (I87395,I691,I86909,I87422,);
nand I_4818 (I87431,I87422,I87053);
nor I_4819 (I87449,I87431,I87215);
nor I_4820 (I87467,I87422,I87017);
DFFARX1 I_4821 (I87422,I691,I86909,I87494,);
not I_4822 (I87503,I87494);
nor I_4823 (I87521,I87503,I87179);
not I_4824 (I87539,I698);
DFFARX1 I_4825 (I87170,I691,I87539,I87566,);
nand I_4826 (I87575,I87170,I87269);
and I_4827 (I87593,I87575,I86963);
DFFARX1 I_4828 (I87593,I691,I87539,I87620,);
nor I_4829 (I87629,I87620,I87566);
not I_4830 (I87647,I87620);
DFFARX1 I_4831 (I87251,I691,I87539,I87674,);
nand I_4832 (I87683,I87674,I87449);
not I_4833 (I87701,I87683);
DFFARX1 I_4834 (I87701,I691,I87539,I87728,);
not I_4835 (I87737,I87728);
nor I_4836 (I87755,I87566,I87683);
nor I_4837 (I87773,I87620,I87755);
DFFARX1 I_4838 (I87521,I691,I87539,I87800,);
DFFARX1 I_4839 (I87800,I691,I87539,I87818,);
not I_4840 (I87827,I87818);
not I_4841 (I87845,I87800);
nand I_4842 (I87863,I87845,I87647);
nand I_4843 (I87881,I87467,I87467);
and I_4844 (I87899,I87881,I87314);
DFFARX1 I_4845 (I87899,I691,I87539,I87926,);
nor I_4846 (I87935,I87926,I87566);
DFFARX1 I_4847 (I87935,I691,I87539,I87962,);
DFFARX1 I_4848 (I87926,I691,I87539,I87980,);
nor I_4849 (I87989,I87332,I87467);
not I_4850 (I88007,I87989);
nor I_4851 (I88025,I87827,I88007);
nand I_4852 (I88043,I87845,I88007);
nor I_4853 (I88061,I87566,I87989);
DFFARX1 I_4854 (I87989,I691,I87539,I88088,);
not I_4855 (I88097,I698);
DFFARX1 I_4856 (I87773,I691,I88097,I88124,);
not I_4857 (I88133,I88124);
nand I_4858 (I88151,I87962,I87962);
and I_4859 (I88169,I88151,I87980);
DFFARX1 I_4860 (I88169,I691,I88097,I88196,);
DFFARX1 I_4861 (I88196,I691,I88097,I88214,);
DFFARX1 I_4862 (I88025,I691,I88097,I88232,);
nand I_4863 (I88241,I88232,I87629);
not I_4864 (I88259,I88241);
DFFARX1 I_4865 (I88259,I691,I88097,I88286,);
not I_4866 (I88295,I88286);
nor I_4867 (I88313,I88133,I88295);
DFFARX1 I_4868 (I88061,I691,I88097,I88340,);
nor I_4869 (I88349,I88340,I88196);
nor I_4870 (I88367,I88340,I88259);
nand I_4871 (I88385,I87737,I88043);
and I_4872 (I88403,I88385,I87863);
DFFARX1 I_4873 (I88403,I691,I88097,I88430,);
not I_4874 (I88439,I88430);
nand I_4875 (I88457,I88439,I88340);
nand I_4876 (I88475,I88439,I88241);
nor I_4877 (I88493,I88088,I88043);
and I_4878 (I88511,I88340,I88493);
nor I_4879 (I88529,I88439,I88511);
DFFARX1 I_4880 (I88529,I691,I88097,I88556,);
nor I_4881 (I88565,I88124,I88493);
DFFARX1 I_4882 (I88565,I691,I88097,I88592,);
nor I_4883 (I88601,I88430,I88493);
not I_4884 (I88619,I88601);
nand I_4885 (I88637,I88619,I88457);
not I_4886 (I88655,I698);
DFFARX1 I_4887 (I88367,I691,I88655,I88682,);
and I_4888 (I88691,I88682,I88637);
DFFARX1 I_4889 (I88691,I691,I88655,I88718,);
DFFARX1 I_4890 (I88556,I691,I88655,I88736,);
not I_4891 (I88745,I88592);
not I_4892 (I88763,I88592);
nand I_4893 (I88781,I88763,I88745);
nor I_4894 (I88799,I88736,I88781);
DFFARX1 I_4895 (I88781,I691,I88655,I88826,);
not I_4896 (I88835,I88826);
not I_4897 (I88853,I88214);
nand I_4898 (I88871,I88763,I88853);
DFFARX1 I_4899 (I88871,I691,I88655,I88898,);
not I_4900 (I88907,I88898);
not I_4901 (I88925,I88349);
nand I_4902 (I88943,I88925,I88367);
and I_4903 (I88961,I88745,I88943);
nor I_4904 (I88979,I88871,I88961);
DFFARX1 I_4905 (I88979,I691,I88655,I89006,);
DFFARX1 I_4906 (I88961,I691,I88655,I89024,);
nor I_4907 (I89033,I88349,I88313);
nor I_4908 (I89051,I88871,I89033);
or I_4909 (I89069,I88349,I88313);
nor I_4910 (I89087,I88475,I88475);
DFFARX1 I_4911 (I89087,I691,I88655,I89114,);
not I_4912 (I89123,I89114);
nor I_4913 (I89141,I89123,I88907);
nand I_4914 (I89159,I89123,I88736);
not I_4915 (I89177,I88475);
nand I_4916 (I89195,I89177,I88853);
nand I_4917 (I89213,I89123,I89195);
nand I_4918 (I89231,I89213,I89159);
nand I_4919 (I89249,I89195,I89069);
not I_4920 (I89267,I698);
DFFARX1 I_4921 (I89006,I691,I89267,I89294,);
not I_4922 (I89303,I89294);
DFFARX1 I_4923 (I89249,I691,I89267,I89330,);
not I_4924 (I89339,I89006);
nand I_4925 (I89357,I89339,I88799);
not I_4926 (I89375,I89357);
nor I_4927 (I89393,I89375,I89024);
nor I_4928 (I89411,I89303,I89393);
DFFARX1 I_4929 (I89411,I691,I89267,I89438,);
not I_4930 (I89447,I89024);
nand I_4931 (I89465,I89447,I89375);
and I_4932 (I89483,I89447,I88835);
nand I_4933 (I89501,I89483,I88799);
nor I_4934 (I89519,I89501,I89447);
and I_4935 (I89537,I89330,I89501);
not I_4936 (I89555,I89501);
nand I_4937 (I89573,I89330,I89555);
nor I_4938 (I89591,I89294,I89501);
not I_4939 (I89609,I89231);
nor I_4940 (I89627,I89609,I88835);
nand I_4941 (I89645,I89627,I89447);
nor I_4942 (I89663,I89357,I89645);
nor I_4943 (I89681,I89609,I88718);
and I_4944 (I89699,I89681,I89051);
or I_4945 (I89717,I89699,I89141);
DFFARX1 I_4946 (I89717,I691,I89267,I89744,);
nor I_4947 (I89753,I89744,I89465);
DFFARX1 I_4948 (I89753,I691,I89267,I89780,);
DFFARX1 I_4949 (I89744,I691,I89267,I89798,);
not I_4950 (I89807,I89744);
nor I_4951 (I89825,I89807,I89330);
nor I_4952 (I89843,I89627,I89825);
DFFARX1 I_4953 (I89843,I691,I89267,I89870,);
not I_4954 (I89879,I698);
DFFARX1 I_4955 (I89780,I691,I89879,I89906,);
not I_4956 (I89915,I89906);
nand I_4957 (I89933,I89573,I89438);
and I_4958 (I89951,I89933,I89798);
DFFARX1 I_4959 (I89951,I691,I89879,I89978,);
not I_4960 (I89987,I89870);
DFFARX1 I_4961 (I89537,I691,I89879,I90014,);
not I_4962 (I90023,I90014);
nor I_4963 (I90041,I90023,I89915);
and I_4964 (I90059,I90041,I89870);
nor I_4965 (I90077,I90023,I89987);
nor I_4966 (I90095,I89978,I90077);
DFFARX1 I_4967 (I89519,I691,I89879,I90122,);
nor I_4968 (I90131,I90122,I89978);
not I_4969 (I90149,I90131);
not I_4970 (I90167,I90122);
nor I_4971 (I90185,I90167,I90059);
DFFARX1 I_4972 (I90185,I691,I89879,I90212,);
nand I_4973 (I90221,I89663,I89591);
and I_4974 (I90239,I90221,I89780);
DFFARX1 I_4975 (I90239,I691,I89879,I90266,);
nor I_4976 (I90275,I90266,I90122);
DFFARX1 I_4977 (I90275,I691,I89879,I90302,);
nand I_4978 (I90311,I90266,I90167);
nand I_4979 (I90329,I90149,I90311);
not I_4980 (I90347,I90266);
nor I_4981 (I90365,I90347,I90059);
DFFARX1 I_4982 (I90365,I691,I89879,I90392,);
nor I_4983 (I90401,I89591,I89591);
or I_4984 (I90419,I90122,I90401);
nor I_4985 (I90437,I90266,I90401);
or I_4986 (I90455,I89978,I90401);
DFFARX1 I_4987 (I90401,I691,I89879,I90482,);
not I_4988 (I90491,I698);
DFFARX1 I_4989 (I90419,I691,I90491,I90518,);
DFFARX1 I_4990 (I90518,I691,I90491,I90536,);
not I_4991 (I90545,I90536);
not I_4992 (I90563,I90518);
DFFARX1 I_4993 (I90329,I691,I90491,I90590,);
not I_4994 (I90599,I90590);
and I_4995 (I90617,I90563,I90095);
not I_4996 (I90635,I90302);
nand I_4997 (I90653,I90635,I90095);
not I_4998 (I90671,I90437);
nor I_4999 (I90689,I90671,I90482);
nand I_5000 (I90707,I90689,I90392);
nor I_5001 (I90725,I90707,I90653);
DFFARX1 I_5002 (I90725,I691,I90491,I90752,);
not I_5003 (I90761,I90707);
not I_5004 (I90779,I90482);
nand I_5005 (I90797,I90779,I90095);
nor I_5006 (I90815,I90482,I90302);
nand I_5007 (I90833,I90617,I90815);
nand I_5008 (I90851,I90563,I90482);
nand I_5009 (I90869,I90671,I90302);
DFFARX1 I_5010 (I90869,I691,I90491,I90896,);
DFFARX1 I_5011 (I90869,I691,I90491,I90914,);
not I_5012 (I90923,I90302);
nor I_5013 (I90941,I90923,I90455);
and I_5014 (I90959,I90941,I90212);
or I_5015 (I90977,I90959,I90437);
DFFARX1 I_5016 (I90977,I691,I90491,I91004,);
nand I_5017 (I91013,I91004,I90635);
nor I_5018 (I91031,I91013,I90797);
nor I_5019 (I91049,I91004,I90599);
DFFARX1 I_5020 (I91004,I691,I90491,I91076,);
not I_5021 (I91085,I91076);
nor I_5022 (I91103,I91085,I90761);
not I_5023 (I91121,I698);
DFFARX1 I_5024 (I90914,I691,I91121,I91148,);
not I_5025 (I91157,I91148);
DFFARX1 I_5026 (I90752,I691,I91121,I91184,);
not I_5027 (I91193,I91103);
nand I_5028 (I91211,I91193,I91049);
not I_5029 (I91229,I91211);
nor I_5030 (I91247,I91229,I90752);
nor I_5031 (I91265,I91157,I91247);
DFFARX1 I_5032 (I91265,I691,I91121,I91292,);
not I_5033 (I91301,I90752);
nand I_5034 (I91319,I91301,I91229);
and I_5035 (I91337,I91301,I91049);
nand I_5036 (I91355,I91337,I90545);
nor I_5037 (I91373,I91355,I91301);
and I_5038 (I91391,I91184,I91355);
not I_5039 (I91409,I91355);
nand I_5040 (I91427,I91184,I91409);
nor I_5041 (I91445,I91148,I91355);
not I_5042 (I91463,I90833);
nor I_5043 (I91481,I91463,I91049);
nand I_5044 (I91499,I91481,I91301);
nor I_5045 (I91517,I91211,I91499);
nor I_5046 (I91535,I91463,I90851);
and I_5047 (I91553,I91535,I90896);
or I_5048 (I91571,I91553,I91031);
DFFARX1 I_5049 (I91571,I691,I91121,I91598,);
nor I_5050 (I91607,I91598,I91319);
DFFARX1 I_5051 (I91607,I691,I91121,I91634,);
DFFARX1 I_5052 (I91598,I691,I91121,I91652,);
not I_5053 (I91661,I91598);
nor I_5054 (I91679,I91661,I91184);
nor I_5055 (I91697,I91481,I91679);
DFFARX1 I_5056 (I91697,I691,I91121,I91724,);
not I_5057 (I91733,I698);
DFFARX1 I_5058 (I91445,I691,I91733,I91760,);
DFFARX1 I_5059 (I91760,I691,I91733,I91778,);
not I_5060 (I91787,I91778);
not I_5061 (I91805,I91760);
nand I_5062 (I91823,I91634,I91724);
and I_5063 (I91841,I91823,I91652);
DFFARX1 I_5064 (I91841,I691,I91733,I91868,);
not I_5065 (I91877,I91868);
DFFARX1 I_5066 (I91427,I691,I91733,I91904,);
and I_5067 (I91913,I91904,I91517);
nand I_5068 (I91931,I91904,I91517);
nand I_5069 (I91949,I91877,I91931);
DFFARX1 I_5070 (I91373,I691,I91733,I91976,);
nor I_5071 (I91985,I91976,I91913);
DFFARX1 I_5072 (I91985,I691,I91733,I92012,);
nor I_5073 (I92021,I91976,I91868);
nand I_5074 (I92039,I91634,I91391);
and I_5075 (I92057,I92039,I91292);
DFFARX1 I_5076 (I92057,I691,I91733,I92084,);
nor I_5077 (I92093,I92084,I91976);
not I_5078 (I92111,I92084);
nor I_5079 (I92129,I92111,I91877);
nor I_5080 (I92147,I91805,I92129);
DFFARX1 I_5081 (I92147,I691,I91733,I92174,);
nor I_5082 (I92183,I92111,I91976);
nor I_5083 (I92201,I91445,I91391);
nor I_5084 (I92219,I92201,I92183);
not I_5085 (I92237,I92201);
nand I_5086 (I92255,I91931,I92237);
DFFARX1 I_5087 (I92201,I691,I91733,I92282,);
DFFARX1 I_5088 (I92201,I691,I91733,I92300,);
not I_5089 (I92309,I698);
DFFARX1 I_5090 (I91949,I691,I92309,I92336,);
not I_5091 (I92345,I92336);
nand I_5092 (I92363,I92093,I92255);
and I_5093 (I92381,I92363,I92300);
DFFARX1 I_5094 (I92381,I691,I92309,I92408,);
DFFARX1 I_5095 (I92408,I691,I92309,I92426,);
DFFARX1 I_5096 (I92282,I691,I92309,I92444,);
nand I_5097 (I92453,I92444,I91787);
not I_5098 (I92471,I92453);
DFFARX1 I_5099 (I92471,I691,I92309,I92498,);
not I_5100 (I92507,I92498);
nor I_5101 (I92525,I92345,I92507);
DFFARX1 I_5102 (I92012,I691,I92309,I92552,);
nor I_5103 (I92561,I92552,I92408);
nor I_5104 (I92579,I92552,I92471);
nand I_5105 (I92597,I92021,I92174);
and I_5106 (I92615,I92597,I92219);
DFFARX1 I_5107 (I92615,I691,I92309,I92642,);
not I_5108 (I92651,I92642);
nand I_5109 (I92669,I92651,I92552);
nand I_5110 (I92687,I92651,I92453);
nor I_5111 (I92705,I92012,I92174);
and I_5112 (I92723,I92552,I92705);
nor I_5113 (I92741,I92651,I92723);
DFFARX1 I_5114 (I92741,I691,I92309,I92768,);
nor I_5115 (I92777,I92336,I92705);
DFFARX1 I_5116 (I92777,I691,I92309,I92804,);
nor I_5117 (I92813,I92642,I92705);
not I_5118 (I92831,I92813);
nand I_5119 (I92849,I92831,I92669);
not I_5120 (I92867,I698);
DFFARX1 I_5121 (I92849,I691,I92867,I92894,);
DFFARX1 I_5122 (I92687,I691,I92867,I92912,);
not I_5123 (I92921,I92912);
nor I_5124 (I92939,I92894,I92921);
DFFARX1 I_5125 (I92921,I691,I92867,I92966,);
nor I_5126 (I92975,I92525,I92579);
and I_5127 (I92993,I92975,I92804);
nor I_5128 (I93011,I92993,I92525);
not I_5129 (I93029,I92525);
and I_5130 (I93047,I93029,I92687);
nand I_5131 (I93065,I93047,I92426);
nor I_5132 (I93083,I93029,I93065);
DFFARX1 I_5133 (I93083,I691,I92867,I93110,);
not I_5134 (I93119,I93065);
nand I_5135 (I93137,I92921,I93119);
nand I_5136 (I93155,I92993,I93119);
DFFARX1 I_5137 (I93029,I691,I92867,I93182,);
not I_5138 (I93191,I92561);
nor I_5139 (I93209,I93191,I92687);
nor I_5140 (I93227,I93209,I93011);
DFFARX1 I_5141 (I93227,I691,I92867,I93254,);
not I_5142 (I93263,I93209);
DFFARX1 I_5143 (I93263,I691,I92867,I93290,);
not I_5144 (I93299,I93290);
nor I_5145 (I93317,I93299,I93209);
nor I_5146 (I93335,I93191,I92804);
and I_5147 (I93353,I93335,I92768);
or I_5148 (I93371,I93353,I92579);
DFFARX1 I_5149 (I93371,I691,I92867,I93398,);
not I_5150 (I93407,I93398);
nand I_5151 (I93425,I93407,I93119);
not I_5152 (I93443,I93425);
nand I_5153 (I93461,I93425,I93137);
nand I_5154 (I93479,I93407,I92993);
not I_5155 (I93497,I698);
DFFARX1 I_5156 (I93317,I691,I93497,I93524,);
DFFARX1 I_5157 (I93524,I691,I93497,I93542,);
not I_5158 (I93551,I93542);
not I_5159 (I93569,I93524);
DFFARX1 I_5160 (I93155,I691,I93497,I93596,);
not I_5161 (I93605,I93596);
and I_5162 (I93623,I93569,I93479);
not I_5163 (I93641,I93110);
nand I_5164 (I93659,I93641,I93479);
not I_5165 (I93677,I93182);
nor I_5166 (I93695,I93677,I93110);
nand I_5167 (I93713,I93695,I93254);
nor I_5168 (I93731,I93713,I93659);
DFFARX1 I_5169 (I93731,I691,I93497,I93758,);
not I_5170 (I93767,I93713);
not I_5171 (I93785,I93110);
nand I_5172 (I93803,I93785,I93479);
nor I_5173 (I93821,I93110,I93110);
nand I_5174 (I93839,I93623,I93821);
nand I_5175 (I93857,I93569,I93110);
nand I_5176 (I93875,I93677,I93461);
DFFARX1 I_5177 (I93875,I691,I93497,I93902,);
DFFARX1 I_5178 (I93875,I691,I93497,I93920,);
not I_5179 (I93929,I93461);
nor I_5180 (I93947,I93929,I93443);
and I_5181 (I93965,I93947,I92966);
or I_5182 (I93983,I93965,I92939);
DFFARX1 I_5183 (I93983,I691,I93497,I94010,);
nand I_5184 (I94019,I94010,I93641);
nor I_5185 (I94037,I94019,I93803);
nor I_5186 (I94055,I94010,I93605);
DFFARX1 I_5187 (I94010,I691,I93497,I94082,);
not I_5188 (I94091,I94082);
nor I_5189 (I94109,I94091,I93767);
not I_5190 (I94127,I698);
DFFARX1 I_5191 (I93758,I691,I94127,I94154,);
not I_5192 (I94163,I94154);
nand I_5193 (I94181,I94055,I93551);
and I_5194 (I94199,I94181,I93839);
DFFARX1 I_5195 (I94199,I691,I94127,I94226,);
not I_5196 (I94235,I94037);
DFFARX1 I_5197 (I93758,I691,I94127,I94262,);
not I_5198 (I94271,I94262);
nor I_5199 (I94289,I94271,I94163);
and I_5200 (I94307,I94289,I94037);
nor I_5201 (I94325,I94271,I94235);
nor I_5202 (I94343,I94226,I94325);
DFFARX1 I_5203 (I94109,I691,I94127,I94370,);
nor I_5204 (I94379,I94370,I94226);
not I_5205 (I94397,I94379);
not I_5206 (I94415,I94370);
nor I_5207 (I94433,I94415,I94307);
DFFARX1 I_5208 (I94433,I691,I94127,I94460,);
nand I_5209 (I94469,I94055,I93857);
and I_5210 (I94487,I94469,I93920);
DFFARX1 I_5211 (I94487,I691,I94127,I94514,);
nor I_5212 (I94523,I94514,I94370);
DFFARX1 I_5213 (I94523,I691,I94127,I94550,);
nand I_5214 (I94559,I94514,I94415);
nand I_5215 (I94577,I94397,I94559);
not I_5216 (I94595,I94514);
nor I_5217 (I94613,I94595,I94307);
DFFARX1 I_5218 (I94613,I691,I94127,I94640,);
nor I_5219 (I94649,I93902,I93857);
or I_5220 (I94667,I94370,I94649);
nor I_5221 (I94685,I94514,I94649);
or I_5222 (I94703,I94226,I94649);
DFFARX1 I_5223 (I94649,I691,I94127,I94730,);
not I_5224 (I94739,I698);
DFFARX1 I_5225 (I620,I691,I94739,I94766,);
not I_5226 (I94775,I94766);
nand I_5227 (I94793,I292,I484);
and I_5228 (I94811,I94793,I412);
DFFARX1 I_5229 (I94811,I691,I94739,I94838,);
not I_5230 (I94847,I172);
DFFARX1 I_5231 (I356,I691,I94739,I94874,);
not I_5232 (I94883,I94874);
nor I_5233 (I94901,I94883,I94775);
and I_5234 (I94919,I94901,I172);
nor I_5235 (I94937,I94883,I94847);
nor I_5236 (I94955,I94838,I94937);
DFFARX1 I_5237 (I196,I691,I94739,I94982,);
nor I_5238 (I94991,I94982,I94838);
not I_5239 (I95009,I94991);
not I_5240 (I95027,I94982);
nor I_5241 (I95045,I95027,I94919);
DFFARX1 I_5242 (I95045,I691,I94739,I95072,);
nand I_5243 (I95081,I76,I644);
and I_5244 (I95099,I95081,I204);
DFFARX1 I_5245 (I95099,I691,I94739,I95126,);
nor I_5246 (I95135,I95126,I94982);
DFFARX1 I_5247 (I95135,I691,I94739,I95162,);
nand I_5248 (I95171,I95126,I95027);
nand I_5249 (I95189,I95009,I95171);
not I_5250 (I95207,I95126);
nor I_5251 (I95225,I95207,I94919);
DFFARX1 I_5252 (I95225,I691,I94739,I95252,);
nor I_5253 (I95261,I548,I644);
or I_5254 (I95279,I94982,I95261);
nor I_5255 (I95297,I95126,I95261);
or I_5256 (I95315,I94838,I95261);
DFFARX1 I_5257 (I95261,I691,I94739,I95342,);
not I_5258 (I95351,I698);
DFFARX1 I_5259 (I95297,I691,I95351,I95378,);
DFFARX1 I_5260 (I95378,I691,I95351,I95396,);
not I_5261 (I95405,I95396);
not I_5262 (I95423,I95378);
nand I_5263 (I95441,I95342,I94955);
and I_5264 (I95459,I95441,I95297);
DFFARX1 I_5265 (I95459,I691,I95351,I95486,);
not I_5266 (I95495,I95486);
DFFARX1 I_5267 (I95189,I691,I95351,I95522,);
and I_5268 (I95531,I95522,I95315);
nand I_5269 (I95549,I95522,I95315);
nand I_5270 (I95567,I95495,I95549);
DFFARX1 I_5271 (I95162,I691,I95351,I95594,);
nor I_5272 (I95603,I95594,I95531);
DFFARX1 I_5273 (I95603,I691,I95351,I95630,);
nor I_5274 (I95639,I95594,I95486);
nand I_5275 (I95657,I95162,I95279);
and I_5276 (I95675,I95657,I95252);
DFFARX1 I_5277 (I95675,I691,I95351,I95702,);
nor I_5278 (I95711,I95702,I95594);
not I_5279 (I95729,I95702);
nor I_5280 (I95747,I95729,I95495);
nor I_5281 (I95765,I95423,I95747);
DFFARX1 I_5282 (I95765,I691,I95351,I95792,);
nor I_5283 (I95801,I95729,I95594);
nor I_5284 (I95819,I95072,I95279);
nor I_5285 (I95837,I95819,I95801);
not I_5286 (I95855,I95819);
nand I_5287 (I95873,I95549,I95855);
DFFARX1 I_5288 (I95819,I691,I95351,I95900,);
DFFARX1 I_5289 (I95819,I691,I95351,I95918,);
not I_5290 (I95927,I698);
DFFARX1 I_5291 (I95567,I691,I95927,I95954,);
not I_5292 (I95963,I95954);
nand I_5293 (I95981,I95711,I95873);
and I_5294 (I95999,I95981,I95918);
DFFARX1 I_5295 (I95999,I691,I95927,I96026,);
DFFARX1 I_5296 (I96026,I691,I95927,I96044,);
DFFARX1 I_5297 (I95900,I691,I95927,I96062,);
nand I_5298 (I96071,I96062,I95405);
not I_5299 (I96089,I96071);
DFFARX1 I_5300 (I96089,I691,I95927,I96116,);
not I_5301 (I96125,I96116);
nor I_5302 (I96143,I95963,I96125);
DFFARX1 I_5303 (I95630,I691,I95927,I96170,);
nor I_5304 (I96179,I96170,I96026);
nor I_5305 (I96197,I96170,I96089);
nand I_5306 (I96215,I95639,I95792);
and I_5307 (I96233,I96215,I95837);
DFFARX1 I_5308 (I96233,I691,I95927,I96260,);
not I_5309 (I96269,I96260);
nand I_5310 (I96287,I96269,I96170);
nand I_5311 (I96305,I96269,I96071);
nor I_5312 (I96323,I95630,I95792);
and I_5313 (I96341,I96170,I96323);
nor I_5314 (I96359,I96269,I96341);
DFFARX1 I_5315 (I96359,I691,I95927,I96386,);
nor I_5316 (I96395,I95954,I96323);
DFFARX1 I_5317 (I96395,I691,I95927,I96422,);
nor I_5318 (I96431,I96260,I96323);
not I_5319 (I96449,I96431);
nand I_5320 (I96467,I96449,I96287);
not I_5321 (I96485,I698);
DFFARX1 I_5322 (I96305,I691,I96485,I96512,);
not I_5323 (I96521,I96512);
DFFARX1 I_5324 (I96305,I691,I96485,I96548,);
not I_5325 (I96557,I96197);
nand I_5326 (I96575,I96557,I96044);
not I_5327 (I96593,I96575);
nor I_5328 (I96611,I96593,I96179);
nor I_5329 (I96629,I96521,I96611);
DFFARX1 I_5330 (I96629,I691,I96485,I96656,);
not I_5331 (I96665,I96179);
nand I_5332 (I96683,I96665,I96593);
and I_5333 (I96701,I96665,I96467);
nand I_5334 (I96719,I96701,I96422);
nor I_5335 (I96737,I96719,I96665);
and I_5336 (I96755,I96548,I96719);
not I_5337 (I96773,I96719);
nand I_5338 (I96791,I96548,I96773);
nor I_5339 (I96809,I96512,I96719);
not I_5340 (I96827,I96143);
nor I_5341 (I96845,I96827,I96467);
nand I_5342 (I96863,I96845,I96665);
nor I_5343 (I96881,I96575,I96863);
nor I_5344 (I96899,I96827,I96422);
and I_5345 (I96917,I96899,I96197);
or I_5346 (I96935,I96917,I96386);
DFFARX1 I_5347 (I96935,I691,I96485,I96962,);
nor I_5348 (I96971,I96962,I96683);
DFFARX1 I_5349 (I96971,I691,I96485,I96998,);
DFFARX1 I_5350 (I96962,I691,I96485,I97016,);
not I_5351 (I97025,I96962);
nor I_5352 (I97043,I97025,I96548);
nor I_5353 (I97061,I96845,I97043);
DFFARX1 I_5354 (I97061,I691,I96485,I97088,);
not I_5355 (I97097,I698);
DFFARX1 I_5356 (I96809,I691,I97097,I97124,);
DFFARX1 I_5357 (I96737,I691,I97097,I97142,);
not I_5358 (I97151,I97142);
not I_5359 (I97169,I97016);
nor I_5360 (I97187,I97169,I96998);
not I_5361 (I97205,I96656);
nor I_5362 (I97223,I97187,I96881);
nor I_5363 (I97241,I97142,I97223);
DFFARX1 I_5364 (I97241,I691,I97097,I97268,);
nor I_5365 (I97277,I96881,I96998);
nand I_5366 (I97295,I97277,I97016);
DFFARX1 I_5367 (I97295,I691,I97097,I97322,);
nor I_5368 (I97331,I97205,I96881);
nand I_5369 (I97349,I97331,I96755);
nor I_5370 (I97367,I97124,I97349);
DFFARX1 I_5371 (I97367,I691,I97097,I97394,);
not I_5372 (I97403,I97349);
nand I_5373 (I97421,I97142,I97403);
DFFARX1 I_5374 (I97349,I691,I97097,I97448,);
not I_5375 (I97457,I97448);
not I_5376 (I97475,I96881);
not I_5377 (I97493,I97088);
nor I_5378 (I97511,I97493,I96656);
nor I_5379 (I97529,I97457,I97511);
nor I_5380 (I97547,I97493,I96809);
and I_5381 (I97565,I97547,I96998);
or I_5382 (I97583,I97565,I96791);
DFFARX1 I_5383 (I97583,I691,I97097,I97610,);
nor I_5384 (I97619,I97610,I97124);
not I_5385 (I97637,I97610);
and I_5386 (I97655,I97637,I97124);
nor I_5387 (I97673,I97151,I97655);
nand I_5388 (I97691,I97637,I97205);
nor I_5389 (I97709,I97493,I97691);
nand I_5390 (I97727,I97637,I97403);
nand I_5391 (I97745,I97205,I97088);
nor I_5392 (I97763,I97475,I97745);
not I_5393 (I97781,I698);
DFFARX1 I_5394 (I97322,I691,I97781,I97808,);
not I_5395 (I97817,I97808);
nand I_5396 (I97835,I97394,I97619);
and I_5397 (I97853,I97835,I97529);
DFFARX1 I_5398 (I97853,I691,I97781,I97880,);
not I_5399 (I97889,I97421);
DFFARX1 I_5400 (I97709,I691,I97781,I97916,);
not I_5401 (I97925,I97916);
nor I_5402 (I97943,I97925,I97817);
and I_5403 (I97961,I97943,I97421);
nor I_5404 (I97979,I97925,I97889);
nor I_5405 (I97997,I97880,I97979);
DFFARX1 I_5406 (I97394,I691,I97781,I98024,);
nor I_5407 (I98033,I98024,I97880);
not I_5408 (I98051,I98033);
not I_5409 (I98069,I98024);
nor I_5410 (I98087,I98069,I97961);
DFFARX1 I_5411 (I98087,I691,I97781,I98114,);
nand I_5412 (I98123,I97763,I97673);
and I_5413 (I98141,I98123,I97268);
DFFARX1 I_5414 (I98141,I691,I97781,I98168,);
nor I_5415 (I98177,I98168,I98024);
DFFARX1 I_5416 (I98177,I691,I97781,I98204,);
nand I_5417 (I98213,I98168,I98069);
nand I_5418 (I98231,I98051,I98213);
not I_5419 (I98249,I98168);
nor I_5420 (I98267,I98249,I97961);
DFFARX1 I_5421 (I98267,I691,I97781,I98294,);
nor I_5422 (I98303,I97727,I97673);
or I_5423 (I98321,I98024,I98303);
nor I_5424 (I98339,I98168,I98303);
or I_5425 (I98357,I97880,I98303);
DFFARX1 I_5426 (I98303,I691,I97781,I98384,);
not I_5427 (I98393,I698);
DFFARX1 I_5428 (I98321,I691,I98393,I98420,);
DFFARX1 I_5429 (I98420,I691,I98393,I98438,);
not I_5430 (I98447,I98438);
not I_5431 (I98465,I98420);
DFFARX1 I_5432 (I98231,I691,I98393,I98492,);
not I_5433 (I98501,I98492);
and I_5434 (I98519,I98465,I97997);
not I_5435 (I98537,I98204);
nand I_5436 (I98555,I98537,I97997);
not I_5437 (I98573,I98339);
nor I_5438 (I98591,I98573,I98384);
nand I_5439 (I98609,I98591,I98294);
nor I_5440 (I98627,I98609,I98555);
DFFARX1 I_5441 (I98627,I691,I98393,I98654,);
not I_5442 (I98663,I98609);
not I_5443 (I98681,I98384);
nand I_5444 (I98699,I98681,I97997);
nor I_5445 (I98717,I98384,I98204);
nand I_5446 (I98735,I98519,I98717);
nand I_5447 (I98753,I98465,I98384);
nand I_5448 (I98771,I98573,I98204);
DFFARX1 I_5449 (I98771,I691,I98393,I98798,);
DFFARX1 I_5450 (I98771,I691,I98393,I98816,);
not I_5451 (I98825,I98204);
nor I_5452 (I98843,I98825,I98357);
and I_5453 (I98861,I98843,I98114);
or I_5454 (I98879,I98861,I98339);
DFFARX1 I_5455 (I98879,I691,I98393,I98906,);
nand I_5456 (I98915,I98906,I98537);
nor I_5457 (I98933,I98915,I98699);
nor I_5458 (I98951,I98906,I98501);
DFFARX1 I_5459 (I98906,I691,I98393,I98978,);
not I_5460 (I98987,I98978);
nor I_5461 (I99005,I98987,I98663);
not I_5462 (I99023,I698);
DFFARX1 I_5463 (I98753,I691,I99023,I99050,);
not I_5464 (I99059,I99050);
nand I_5465 (I99077,I98951,I98798);
and I_5466 (I99095,I99077,I98735);
DFFARX1 I_5467 (I99095,I691,I99023,I99122,);
DFFARX1 I_5468 (I99122,I691,I99023,I99140,);
DFFARX1 I_5469 (I99005,I691,I99023,I99158,);
nand I_5470 (I99167,I99158,I98816);
not I_5471 (I99185,I99167);
DFFARX1 I_5472 (I99185,I691,I99023,I99212,);
not I_5473 (I99221,I99212);
nor I_5474 (I99239,I99059,I99221);
DFFARX1 I_5475 (I98933,I691,I99023,I99266,);
nor I_5476 (I99275,I99266,I99122);
nor I_5477 (I99293,I99266,I99185);
nand I_5478 (I99311,I98654,I98447);
and I_5479 (I99329,I99311,I98951);
DFFARX1 I_5480 (I99329,I691,I99023,I99356,);
not I_5481 (I99365,I99356);
nand I_5482 (I99383,I99365,I99266);
nand I_5483 (I99401,I99365,I99167);
nor I_5484 (I99419,I98654,I98447);
and I_5485 (I99437,I99266,I99419);
nor I_5486 (I99455,I99365,I99437);
DFFARX1 I_5487 (I99455,I691,I99023,I99482,);
nor I_5488 (I99491,I99050,I99419);
DFFARX1 I_5489 (I99491,I691,I99023,I99518,);
nor I_5490 (I99527,I99356,I99419);
not I_5491 (I99545,I99527);
nand I_5492 (I99563,I99545,I99383);
not I_5493 (I99581,I698);
DFFARX1 I_5494 (I99482,I691,I99581,I99608,);
not I_5495 (I99617,I99608);
nand I_5496 (I99635,I99293,I99239);
and I_5497 (I99653,I99635,I99140);
DFFARX1 I_5498 (I99653,I691,I99581,I99680,);
not I_5499 (I99689,I99563);
DFFARX1 I_5500 (I99401,I691,I99581,I99716,);
not I_5501 (I99725,I99716);
nor I_5502 (I99743,I99725,I99617);
and I_5503 (I99761,I99743,I99563);
nor I_5504 (I99779,I99725,I99689);
nor I_5505 (I99797,I99680,I99779);
DFFARX1 I_5506 (I99518,I691,I99581,I99824,);
nor I_5507 (I99833,I99824,I99680);
not I_5508 (I99851,I99833);
not I_5509 (I99869,I99824);
nor I_5510 (I99887,I99869,I99761);
DFFARX1 I_5511 (I99887,I691,I99581,I99914,);
nand I_5512 (I99923,I99518,I99293);
and I_5513 (I99941,I99923,I99401);
DFFARX1 I_5514 (I99941,I691,I99581,I99968,);
nor I_5515 (I99977,I99968,I99824);
DFFARX1 I_5516 (I99977,I691,I99581,I100004,);
nand I_5517 (I100013,I99968,I99869);
nand I_5518 (I100031,I99851,I100013);
not I_5519 (I100049,I99968);
nor I_5520 (I100067,I100049,I99761);
DFFARX1 I_5521 (I100067,I691,I99581,I100094,);
nor I_5522 (I100103,I99275,I99293);
or I_5523 (I100121,I99824,I100103);
nor I_5524 (I100139,I99968,I100103);
or I_5525 (I100157,I99680,I100103);
DFFARX1 I_5526 (I100103,I691,I99581,I100184,);
not I_5527 (I100193,I698);
DFFARX1 I_5528 (I100139,I691,I100193,I100220,);
DFFARX1 I_5529 (I100220,I691,I100193,I100238,);
not I_5530 (I100247,I100238);
not I_5531 (I100265,I100220);
DFFARX1 I_5532 (I99797,I691,I100193,I100292,);
nand I_5533 (I100301,I100292,I100184);
not I_5534 (I100319,I100184);
not I_5535 (I100337,I100157);
nand I_5536 (I100355,I100031,I100004);
and I_5537 (I100373,I100031,I100004);
not I_5538 (I100391,I99914);
nand I_5539 (I100409,I100391,I100337);
nor I_5540 (I100427,I100409,I100301);
nor I_5541 (I100445,I100319,I100409);
nand I_5542 (I100463,I100373,I100445);
not I_5543 (I100481,I100094);
nor I_5544 (I100499,I100481,I100031);
nor I_5545 (I100517,I100499,I99914);
nor I_5546 (I100535,I100265,I100517);
DFFARX1 I_5547 (I100535,I691,I100193,I100562,);
not I_5548 (I100571,I100499);
DFFARX1 I_5549 (I100571,I691,I100193,I100598,);
and I_5550 (I100607,I100292,I100499);
nor I_5551 (I100625,I100481,I100004);
and I_5552 (I100643,I100625,I100121);
or I_5553 (I100661,I100643,I100139);
DFFARX1 I_5554 (I100661,I691,I100193,I100688,);
nor I_5555 (I100697,I100688,I100391);
DFFARX1 I_5556 (I100697,I691,I100193,I100724,);
nand I_5557 (I100733,I100688,I100292);
nand I_5558 (I100751,I100391,I100733);
nor I_5559 (I100769,I100751,I100355);
not I_5560 (I100787,I698);
DFFARX1 I_5561 (I100607,I691,I100787,I100814,);
nand I_5562 (I100823,I100814,I100562);
not I_5563 (I100841,I100823);
DFFARX1 I_5564 (I100427,I691,I100787,I100868,);
not I_5565 (I100877,I100868);
nor I_5566 (I100895,I100247,I100598);
not I_5567 (I100913,I100895);
DFFARX1 I_5568 (I100913,I691,I100787,I100940,);
or I_5569 (I100949,I100724,I100247);
DFFARX1 I_5570 (I100949,I691,I100787,I100976,);
not I_5571 (I100985,I100724);
nor I_5572 (I101003,I100985,I100427);
nor I_5573 (I101021,I101003,I100598);
nor I_5574 (I101039,I100427,I100463);
nor I_5575 (I101057,I100877,I101039);
nor I_5576 (I101075,I100841,I101057);
not I_5577 (I101093,I101039);
nand I_5578 (I101111,I101093,I100823);
nand I_5579 (I101129,I101093,I100895);
nor I_5580 (I101147,I101039,I101021);
nor I_5581 (I101165,I100769,I100724);
not I_5582 (I101183,I101165);
DFFARX1 I_5583 (I101165,I691,I100787,I101210,);
not I_5584 (I101219,I101210);
nor I_5585 (I101237,I100769,I100463);
DFFARX1 I_5586 (I101237,I691,I100787,I101264,);
and I_5587 (I101273,I101264,I100247);
nor I_5588 (I101291,I101273,I101183);
DFFARX1 I_5589 (I101291,I691,I100787,I101318,);
nor I_5590 (I101327,I101264,I101021);
DFFARX1 I_5591 (I101327,I691,I100787,I101354,);
nor I_5592 (I101363,I101264,I100913);
not I_5593 (I101381,I698);
DFFARX1 I_5594 (I101129,I691,I101381,I101408,);
not I_5595 (I101417,I101408);
nand I_5596 (I101435,I101354,I101318);
and I_5597 (I101453,I101435,I101147);
DFFARX1 I_5598 (I101453,I691,I101381,I101480,);
DFFARX1 I_5599 (I101480,I691,I101381,I101498,);
DFFARX1 I_5600 (I100976,I691,I101381,I101516,);
nand I_5601 (I101525,I101516,I101075);
not I_5602 (I101543,I101525);
DFFARX1 I_5603 (I101543,I691,I101381,I101570,);
not I_5604 (I101579,I101570);
nor I_5605 (I101597,I101417,I101579);
DFFARX1 I_5606 (I100940,I691,I101381,I101624,);
nor I_5607 (I101633,I101624,I101480);
nor I_5608 (I101651,I101624,I101543);
nand I_5609 (I101669,I101111,I101219);
and I_5610 (I101687,I101669,I101363);
DFFARX1 I_5611 (I101687,I691,I101381,I101714,);
not I_5612 (I101723,I101714);
nand I_5613 (I101741,I101723,I101624);
nand I_5614 (I101759,I101723,I101525);
nor I_5615 (I101777,I101354,I101219);
and I_5616 (I101795,I101624,I101777);
nor I_5617 (I101813,I101723,I101795);
DFFARX1 I_5618 (I101813,I691,I101381,I101840,);
nor I_5619 (I101849,I101408,I101777);
DFFARX1 I_5620 (I101849,I691,I101381,I101876,);
nor I_5621 (I101885,I101714,I101777);
not I_5622 (I101903,I101885);
nand I_5623 (I101921,I101903,I101741);
not I_5624 (I101939,I698);
DFFARX1 I_5625 (I101759,I691,I101939,I101966,);
DFFARX1 I_5626 (I101651,I691,I101939,I101984,);
not I_5627 (I101993,I101984);
not I_5628 (I102011,I101651);
nor I_5629 (I102029,I102011,I101759);
not I_5630 (I102047,I101498);
nor I_5631 (I102065,I102029,I101633);
nor I_5632 (I102083,I101984,I102065);
DFFARX1 I_5633 (I102083,I691,I101939,I102110,);
nor I_5634 (I102119,I101633,I101759);
nand I_5635 (I102137,I102119,I101651);
DFFARX1 I_5636 (I102137,I691,I101939,I102164,);
nor I_5637 (I102173,I102047,I101633);
nand I_5638 (I102191,I102173,I101876);
nor I_5639 (I102209,I101966,I102191);
DFFARX1 I_5640 (I102209,I691,I101939,I102236,);
not I_5641 (I102245,I102191);
nand I_5642 (I102263,I101984,I102245);
DFFARX1 I_5643 (I102191,I691,I101939,I102290,);
not I_5644 (I102299,I102290);
not I_5645 (I102317,I101633);
not I_5646 (I102335,I101921);
nor I_5647 (I102353,I102335,I101498);
nor I_5648 (I102371,I102299,I102353);
nor I_5649 (I102389,I102335,I101840);
and I_5650 (I102407,I102389,I101597);
or I_5651 (I102425,I102407,I101876);
DFFARX1 I_5652 (I102425,I691,I101939,I102452,);
nor I_5653 (I102461,I102452,I101966);
not I_5654 (I102479,I102452);
and I_5655 (I102497,I102479,I101966);
nor I_5656 (I102515,I101993,I102497);
nand I_5657 (I102533,I102479,I102047);
nor I_5658 (I102551,I102335,I102533);
nand I_5659 (I102569,I102479,I102245);
nand I_5660 (I102587,I102047,I101921);
nor I_5661 (I102605,I102317,I102587);
not I_5662 (I102623,I698);
DFFARX1 I_5663 (I102164,I691,I102623,I102650,);
not I_5664 (I102659,I102650);
nand I_5665 (I102677,I102236,I102461);
and I_5666 (I102695,I102677,I102371);
DFFARX1 I_5667 (I102695,I691,I102623,I102722,);
not I_5668 (I102731,I102263);
DFFARX1 I_5669 (I102551,I691,I102623,I102758,);
not I_5670 (I102767,I102758);
nor I_5671 (I102785,I102767,I102659);
and I_5672 (I102803,I102785,I102263);
nor I_5673 (I102821,I102767,I102731);
nor I_5674 (I102839,I102722,I102821);
DFFARX1 I_5675 (I102236,I691,I102623,I102866,);
nor I_5676 (I102875,I102866,I102722);
not I_5677 (I102893,I102875);
not I_5678 (I102911,I102866);
nor I_5679 (I102929,I102911,I102803);
DFFARX1 I_5680 (I102929,I691,I102623,I102956,);
nand I_5681 (I102965,I102605,I102515);
and I_5682 (I102983,I102965,I102110);
DFFARX1 I_5683 (I102983,I691,I102623,I103010,);
nor I_5684 (I103019,I103010,I102866);
DFFARX1 I_5685 (I103019,I691,I102623,I103046,);
nand I_5686 (I103055,I103010,I102911);
nand I_5687 (I103073,I102893,I103055);
not I_5688 (I103091,I103010);
nor I_5689 (I103109,I103091,I102803);
DFFARX1 I_5690 (I103109,I691,I102623,I103136,);
nor I_5691 (I103145,I102569,I102515);
or I_5692 (I103163,I102866,I103145);
nor I_5693 (I103181,I103010,I103145);
or I_5694 (I103199,I102722,I103145);
DFFARX1 I_5695 (I103145,I691,I102623,I103226,);
not I_5696 (I103235,I698);
DFFARX1 I_5697 (I102839,I691,I103235,I103262,);
and I_5698 (I103271,I103262,I103181);
DFFARX1 I_5699 (I103271,I691,I103235,I103298,);
DFFARX1 I_5700 (I103199,I691,I103235,I103316,);
not I_5701 (I103325,I103046);
not I_5702 (I103343,I103226);
nand I_5703 (I103361,I103343,I103325);
nor I_5704 (I103379,I103316,I103361);
DFFARX1 I_5705 (I103361,I691,I103235,I103406,);
not I_5706 (I103415,I103406);
not I_5707 (I103433,I103163);
nand I_5708 (I103451,I103343,I103433);
DFFARX1 I_5709 (I103451,I691,I103235,I103478,);
not I_5710 (I103487,I103478);
not I_5711 (I103505,I103136);
nand I_5712 (I103523,I103505,I102956);
and I_5713 (I103541,I103325,I103523);
nor I_5714 (I103559,I103451,I103541);
DFFARX1 I_5715 (I103559,I691,I103235,I103586,);
DFFARX1 I_5716 (I103541,I691,I103235,I103604,);
nor I_5717 (I103613,I103136,I103073);
nor I_5718 (I103631,I103451,I103613);
or I_5719 (I103649,I103136,I103073);
nor I_5720 (I103667,I103046,I103181);
DFFARX1 I_5721 (I103667,I691,I103235,I103694,);
not I_5722 (I103703,I103694);
nor I_5723 (I103721,I103703,I103487);
nand I_5724 (I103739,I103703,I103316);
not I_5725 (I103757,I103046);
nand I_5726 (I103775,I103757,I103433);
nand I_5727 (I103793,I103703,I103775);
nand I_5728 (I103811,I103793,I103739);
nand I_5729 (I103829,I103775,I103649);
not I_5730 (I103847,I698);
DFFARX1 I_5731 (I103721,I691,I103847,I103874,);
DFFARX1 I_5732 (I103874,I691,I103847,I103892,);
not I_5733 (I103901,I103892);
DFFARX1 I_5734 (I103586,I691,I103847,I103928,);
not I_5735 (I103937,I103829);
nor I_5736 (I103955,I103874,I103937);
not I_5737 (I103973,I103604);
not I_5738 (I103991,I103631);
nand I_5739 (I104009,I103991,I103604);
nor I_5740 (I104027,I103937,I104009);
nor I_5741 (I104045,I103928,I104027);
DFFARX1 I_5742 (I103991,I691,I103847,I104072,);
nor I_5743 (I104081,I103631,I103415);
nand I_5744 (I104099,I104081,I103379);
nor I_5745 (I104117,I104099,I103973);
nand I_5746 (I104135,I104117,I103829);
DFFARX1 I_5747 (I104099,I691,I103847,I104162,);
nand I_5748 (I104171,I103973,I103631);
nor I_5749 (I104189,I103973,I103631);
nand I_5750 (I104207,I103955,I104189);
not I_5751 (I104225,I103811);
nor I_5752 (I104243,I104225,I104171);
DFFARX1 I_5753 (I104243,I691,I103847,I104270,);
nor I_5754 (I104279,I104225,I103298);
and I_5755 (I104297,I104279,I103586);
or I_5756 (I104315,I104297,I103379);
DFFARX1 I_5757 (I104315,I691,I103847,I104342,);
nor I_5758 (I104351,I104342,I103928);
nor I_5759 (I104369,I103874,I104351);
not I_5760 (I104387,I104342);
nor I_5761 (I104405,I104387,I104045);
DFFARX1 I_5762 (I104405,I691,I103847,I104432,);
nand I_5763 (I104441,I104387,I103973);
nor I_5764 (I104459,I104225,I104441);
not I_5765 (I104477,I698);
DFFARX1 I_5766 (I104270,I691,I104477,I104504,);
not I_5767 (I104513,I104504);
nand I_5768 (I104531,I104432,I104270);
and I_5769 (I104549,I104531,I104459);
DFFARX1 I_5770 (I104549,I691,I104477,I104576,);
not I_5771 (I104585,I104459);
DFFARX1 I_5772 (I104207,I691,I104477,I104612,);
not I_5773 (I104621,I104612);
nor I_5774 (I104639,I104621,I104513);
and I_5775 (I104657,I104639,I104459);
nor I_5776 (I104675,I104621,I104585);
nor I_5777 (I104693,I104576,I104675);
DFFARX1 I_5778 (I104135,I691,I104477,I104720,);
nor I_5779 (I104729,I104720,I104576);
not I_5780 (I104747,I104729);
not I_5781 (I104765,I104720);
nor I_5782 (I104783,I104765,I104657);
DFFARX1 I_5783 (I104783,I691,I104477,I104810,);
nand I_5784 (I104819,I104369,I104162);
and I_5785 (I104837,I104819,I103901);
DFFARX1 I_5786 (I104837,I691,I104477,I104864,);
nor I_5787 (I104873,I104864,I104720);
DFFARX1 I_5788 (I104873,I691,I104477,I104900,);
nand I_5789 (I104909,I104864,I104765);
nand I_5790 (I104927,I104747,I104909);
not I_5791 (I104945,I104864);
nor I_5792 (I104963,I104945,I104657);
DFFARX1 I_5793 (I104963,I691,I104477,I104990,);
nor I_5794 (I104999,I104072,I104162);
or I_5795 (I105017,I104720,I104999);
nor I_5796 (I105035,I104864,I104999);
or I_5797 (I105053,I104576,I104999);
DFFARX1 I_5798 (I104999,I691,I104477,I105080,);
not I_5799 (I105089,I698);
DFFARX1 I_5800 (I104900,I691,I105089,I105116,);
nand I_5801 (I105125,I105116,I105035);
not I_5802 (I105143,I105125);
DFFARX1 I_5803 (I104693,I691,I105089,I105170,);
not I_5804 (I105179,I105170);
not I_5805 (I105197,I104900);
or I_5806 (I105215,I104927,I104900);
nor I_5807 (I105233,I104927,I104900);
or I_5808 (I105251,I104810,I104927);
DFFARX1 I_5809 (I105251,I691,I105089,I105278,);
not I_5810 (I105287,I104990);
nand I_5811 (I105305,I105287,I105035);
nand I_5812 (I105323,I105197,I105305);
and I_5813 (I105341,I105179,I105323);
nor I_5814 (I105359,I104990,I105053);
and I_5815 (I105377,I105179,I105359);
nor I_5816 (I105395,I105143,I105377);
DFFARX1 I_5817 (I105359,I691,I105089,I105422,);
not I_5818 (I105431,I105422);
nor I_5819 (I105449,I105179,I105431);
or I_5820 (I105467,I105251,I105017);
nor I_5821 (I105485,I105017,I104810);
nand I_5822 (I105503,I105323,I105485);
nand I_5823 (I105521,I105467,I105503);
DFFARX1 I_5824 (I105521,I691,I105089,I105548,);
nor I_5825 (I105557,I105485,I105215);
DFFARX1 I_5826 (I105557,I691,I105089,I105584,);
nor I_5827 (I105593,I105017,I105080);
DFFARX1 I_5828 (I105593,I691,I105089,I105620,);
DFFARX1 I_5829 (I105620,I691,I105089,I105638,);
not I_5830 (I105647,I105620);
nand I_5831 (I105665,I105647,I105125);
nand I_5832 (I105683,I105647,I105233);
not I_5833 (I105701,I698);
DFFARX1 I_5834 (I105395,I691,I105701,I105728,);
DFFARX1 I_5835 (I105728,I691,I105701,I105746,);
not I_5836 (I105755,I105746);
DFFARX1 I_5837 (I105638,I691,I105701,I105782,);
not I_5838 (I105791,I105341);
nor I_5839 (I105809,I105728,I105791);
not I_5840 (I105827,I105683);
not I_5841 (I105845,I105665);
nand I_5842 (I105863,I105845,I105683);
nor I_5843 (I105881,I105791,I105863);
nor I_5844 (I105899,I105782,I105881);
DFFARX1 I_5845 (I105845,I691,I105701,I105926,);
nor I_5846 (I105935,I105665,I105341);
nand I_5847 (I105953,I105935,I105548);
nor I_5848 (I105971,I105953,I105827);
nand I_5849 (I105989,I105971,I105341);
DFFARX1 I_5850 (I105953,I691,I105701,I106016,);
nand I_5851 (I106025,I105827,I105665);
nor I_5852 (I106043,I105827,I105665);
nand I_5853 (I106061,I105809,I106043);
not I_5854 (I106079,I105584);
nor I_5855 (I106097,I106079,I106025);
DFFARX1 I_5856 (I106097,I691,I105701,I106124,);
nor I_5857 (I106133,I106079,I105278);
and I_5858 (I106151,I106133,I105584);
or I_5859 (I106169,I106151,I105449);
DFFARX1 I_5860 (I106169,I691,I105701,I106196,);
nor I_5861 (I106205,I106196,I105782);
nor I_5862 (I106223,I105728,I106205);
not I_5863 (I106241,I106196);
nor I_5864 (I106259,I106241,I105899);
DFFARX1 I_5865 (I106259,I691,I105701,I106286,);
nand I_5866 (I106295,I106241,I105827);
nor I_5867 (I106313,I106079,I106295);
not I_5868 (I106331,I698);
DFFARX1 I_5869 (I106124,I691,I106331,I106358,);
not I_5870 (I106367,I106358);
nand I_5871 (I106385,I106286,I106124);
and I_5872 (I106403,I106385,I106313);
DFFARX1 I_5873 (I106403,I691,I106331,I106430,);
not I_5874 (I106439,I106313);
DFFARX1 I_5875 (I106061,I691,I106331,I106466,);
not I_5876 (I106475,I106466);
nor I_5877 (I106493,I106475,I106367);
and I_5878 (I106511,I106493,I106313);
nor I_5879 (I106529,I106475,I106439);
nor I_5880 (I106547,I106430,I106529);
DFFARX1 I_5881 (I105989,I691,I106331,I106574,);
nor I_5882 (I106583,I106574,I106430);
not I_5883 (I106601,I106583);
not I_5884 (I106619,I106574);
nor I_5885 (I106637,I106619,I106511);
DFFARX1 I_5886 (I106637,I691,I106331,I106664,);
nand I_5887 (I106673,I106223,I106016);
and I_5888 (I106691,I106673,I105755);
DFFARX1 I_5889 (I106691,I691,I106331,I106718,);
nor I_5890 (I106727,I106718,I106574);
DFFARX1 I_5891 (I106727,I691,I106331,I106754,);
nand I_5892 (I106763,I106718,I106619);
nand I_5893 (I106781,I106601,I106763);
not I_5894 (I106799,I106718);
nor I_5895 (I106817,I106799,I106511);
DFFARX1 I_5896 (I106817,I691,I106331,I106844,);
nor I_5897 (I106853,I105926,I106016);
or I_5898 (I106871,I106574,I106853);
nor I_5899 (I106889,I106718,I106853);
or I_5900 (I106907,I106430,I106853);
DFFARX1 I_5901 (I106853,I691,I106331,I106934,);
not I_5902 (I106943,I698);
DFFARX1 I_5903 (I106547,I691,I106943,I106970,);
and I_5904 (I106979,I106970,I106889);
DFFARX1 I_5905 (I106979,I691,I106943,I107006,);
DFFARX1 I_5906 (I106907,I691,I106943,I107024,);
not I_5907 (I107033,I106754);
not I_5908 (I107051,I106934);
nand I_5909 (I107069,I107051,I107033);
nor I_5910 (I107087,I107024,I107069);
DFFARX1 I_5911 (I107069,I691,I106943,I107114,);
not I_5912 (I107123,I107114);
not I_5913 (I107141,I106871);
nand I_5914 (I107159,I107051,I107141);
DFFARX1 I_5915 (I107159,I691,I106943,I107186,);
not I_5916 (I107195,I107186);
not I_5917 (I107213,I106844);
nand I_5918 (I107231,I107213,I106664);
and I_5919 (I107249,I107033,I107231);
nor I_5920 (I107267,I107159,I107249);
DFFARX1 I_5921 (I107267,I691,I106943,I107294,);
DFFARX1 I_5922 (I107249,I691,I106943,I107312,);
nor I_5923 (I107321,I106844,I106781);
nor I_5924 (I107339,I107159,I107321);
or I_5925 (I107357,I106844,I106781);
nor I_5926 (I107375,I106754,I106889);
DFFARX1 I_5927 (I107375,I691,I106943,I107402,);
not I_5928 (I107411,I107402);
nor I_5929 (I107429,I107411,I107195);
nand I_5930 (I107447,I107411,I107024);
not I_5931 (I107465,I106754);
nand I_5932 (I107483,I107465,I107141);
nand I_5933 (I107501,I107411,I107483);
nand I_5934 (I107519,I107501,I107447);
nand I_5935 (I107537,I107483,I107357);
not I_5936 (I107555,I698);
DFFARX1 I_5937 (I107429,I691,I107555,I107582,);
DFFARX1 I_5938 (I107582,I691,I107555,I107600,);
not I_5939 (I107609,I107600);
DFFARX1 I_5940 (I107294,I691,I107555,I107636,);
not I_5941 (I107645,I107537);
nor I_5942 (I107663,I107582,I107645);
not I_5943 (I107681,I107312);
not I_5944 (I107699,I107339);
nand I_5945 (I107717,I107699,I107312);
nor I_5946 (I107735,I107645,I107717);
nor I_5947 (I107753,I107636,I107735);
DFFARX1 I_5948 (I107699,I691,I107555,I107780,);
nor I_5949 (I107789,I107339,I107123);
nand I_5950 (I107807,I107789,I107087);
nor I_5951 (I107825,I107807,I107681);
nand I_5952 (I107843,I107825,I107537);
DFFARX1 I_5953 (I107807,I691,I107555,I107870,);
nand I_5954 (I107879,I107681,I107339);
nor I_5955 (I107897,I107681,I107339);
nand I_5956 (I107915,I107663,I107897);
not I_5957 (I107933,I107519);
nor I_5958 (I107951,I107933,I107879);
DFFARX1 I_5959 (I107951,I691,I107555,I107978,);
nor I_5960 (I107987,I107933,I107006);
and I_5961 (I108005,I107987,I107294);
or I_5962 (I108023,I108005,I107087);
DFFARX1 I_5963 (I108023,I691,I107555,I108050,);
nor I_5964 (I108059,I108050,I107636);
nor I_5965 (I108077,I107582,I108059);
not I_5966 (I108095,I108050);
nor I_5967 (I108113,I108095,I107753);
DFFARX1 I_5968 (I108113,I691,I107555,I108140,);
nand I_5969 (I108149,I108095,I107681);
nor I_5970 (I108167,I107933,I108149);
not I_5971 (I108185,I698);
DFFARX1 I_5972 (I108167,I691,I108185,I108212,);
DFFARX1 I_5973 (I108140,I691,I108185,I108230,);
not I_5974 (I108239,I108230);
not I_5975 (I108257,I107978);
nor I_5976 (I108275,I108257,I107870);
not I_5977 (I108293,I107609);
nor I_5978 (I108311,I108275,I107843);
nor I_5979 (I108329,I108230,I108311);
DFFARX1 I_5980 (I108329,I691,I108185,I108356,);
nor I_5981 (I108365,I107843,I107870);
nand I_5982 (I108383,I108365,I107978);
DFFARX1 I_5983 (I108383,I691,I108185,I108410,);
nor I_5984 (I108419,I108293,I107843);
nand I_5985 (I108437,I108419,I108077);
nor I_5986 (I108455,I108212,I108437);
DFFARX1 I_5987 (I108455,I691,I108185,I108482,);
not I_5988 (I108491,I108437);
nand I_5989 (I108509,I108230,I108491);
DFFARX1 I_5990 (I108437,I691,I108185,I108536,);
not I_5991 (I108545,I108536);
not I_5992 (I108563,I107843);
not I_5993 (I108581,I107915);
nor I_5994 (I108599,I108581,I107609);
nor I_5995 (I108617,I108545,I108599);
nor I_5996 (I108635,I108581,I107780);
and I_5997 (I108653,I108635,I107978);
or I_5998 (I108671,I108653,I108167);
DFFARX1 I_5999 (I108671,I691,I108185,I108698,);
nor I_6000 (I108707,I108698,I108212);
not I_6001 (I108725,I108698);
and I_6002 (I108743,I108725,I108212);
nor I_6003 (I108761,I108239,I108743);
nand I_6004 (I108779,I108725,I108293);
nor I_6005 (I108797,I108581,I108779);
nand I_6006 (I108815,I108725,I108491);
nand I_6007 (I108833,I108293,I107915);
nor I_6008 (I108851,I108563,I108833);
not I_6009 (I108869,I698);
DFFARX1 I_6010 (I108410,I691,I108869,I108896,);
not I_6011 (I108905,I108896);
nand I_6012 (I108923,I108482,I108707);
and I_6013 (I108941,I108923,I108617);
DFFARX1 I_6014 (I108941,I691,I108869,I108968,);
not I_6015 (I108977,I108509);
DFFARX1 I_6016 (I108797,I691,I108869,I109004,);
not I_6017 (I109013,I109004);
nor I_6018 (I109031,I109013,I108905);
and I_6019 (I109049,I109031,I108509);
nor I_6020 (I109067,I109013,I108977);
nor I_6021 (I109085,I108968,I109067);
DFFARX1 I_6022 (I108482,I691,I108869,I109112,);
nor I_6023 (I109121,I109112,I108968);
not I_6024 (I109139,I109121);
not I_6025 (I109157,I109112);
nor I_6026 (I109175,I109157,I109049);
DFFARX1 I_6027 (I109175,I691,I108869,I109202,);
nand I_6028 (I109211,I108851,I108761);
and I_6029 (I109229,I109211,I108356);
DFFARX1 I_6030 (I109229,I691,I108869,I109256,);
nor I_6031 (I109265,I109256,I109112);
DFFARX1 I_6032 (I109265,I691,I108869,I109292,);
nand I_6033 (I109301,I109256,I109157);
nand I_6034 (I109319,I109139,I109301);
not I_6035 (I109337,I109256);
nor I_6036 (I109355,I109337,I109049);
DFFARX1 I_6037 (I109355,I691,I108869,I109382,);
nor I_6038 (I109391,I108815,I108761);
or I_6039 (I109409,I109112,I109391);
nor I_6040 (I109427,I109256,I109391);
or I_6041 (I109445,I108968,I109391);
DFFARX1 I_6042 (I109391,I691,I108869,I109472,);
not I_6043 (I109481,I698);
DFFARX1 I_6044 (I109085,I691,I109481,I109508,);
and I_6045 (I109517,I109508,I109427);
DFFARX1 I_6046 (I109517,I691,I109481,I109544,);
DFFARX1 I_6047 (I109445,I691,I109481,I109562,);
not I_6048 (I109571,I109292);
not I_6049 (I109589,I109472);
nand I_6050 (I109607,I109589,I109571);
nor I_6051 (I109625,I109562,I109607);
DFFARX1 I_6052 (I109607,I691,I109481,I109652,);
not I_6053 (I109661,I109652);
not I_6054 (I109679,I109409);
nand I_6055 (I109697,I109589,I109679);
DFFARX1 I_6056 (I109697,I691,I109481,I109724,);
not I_6057 (I109733,I109724);
not I_6058 (I109751,I109382);
nand I_6059 (I109769,I109751,I109202);
and I_6060 (I109787,I109571,I109769);
nor I_6061 (I109805,I109697,I109787);
DFFARX1 I_6062 (I109805,I691,I109481,I109832,);
DFFARX1 I_6063 (I109787,I691,I109481,I109850,);
nor I_6064 (I109859,I109382,I109319);
nor I_6065 (I109877,I109697,I109859);
or I_6066 (I109895,I109382,I109319);
nor I_6067 (I109913,I109292,I109427);
DFFARX1 I_6068 (I109913,I691,I109481,I109940,);
not I_6069 (I109949,I109940);
nor I_6070 (I109967,I109949,I109733);
nand I_6071 (I109985,I109949,I109562);
not I_6072 (I110003,I109292);
nand I_6073 (I110021,I110003,I109679);
nand I_6074 (I110039,I109949,I110021);
nand I_6075 (I110057,I110039,I109985);
nand I_6076 (I110075,I110021,I109895);
not I_6077 (I110093,I698);
DFFARX1 I_6078 (I110075,I691,I110093,I110120,);
not I_6079 (I110129,I110120);
nand I_6080 (I110147,I109850,I109832);
and I_6081 (I110165,I110147,I109625);
DFFARX1 I_6082 (I110165,I691,I110093,I110192,);
DFFARX1 I_6083 (I109661,I691,I110093,I110210,);
and I_6084 (I110219,I110210,I109625);
nor I_6085 (I110237,I110192,I110219);
DFFARX1 I_6086 (I110237,I691,I110093,I110264,);
nand I_6087 (I110273,I110210,I109625);
nand I_6088 (I110291,I110129,I110273);
not I_6089 (I110309,I110291);
DFFARX1 I_6090 (I109832,I691,I110093,I110336,);
DFFARX1 I_6091 (I110336,I691,I110093,I110354,);
nand I_6092 (I110363,I109877,I110057);
and I_6093 (I110381,I110363,I109544);
DFFARX1 I_6094 (I110381,I691,I110093,I110408,);
DFFARX1 I_6095 (I110408,I691,I110093,I110426,);
not I_6096 (I110435,I110426);
not I_6097 (I110453,I110408);
nand I_6098 (I110471,I110453,I110273);
nor I_6099 (I110489,I109967,I110057);
not I_6100 (I110507,I110489);
nor I_6101 (I110525,I110453,I110507);
nor I_6102 (I110543,I110129,I110525);
DFFARX1 I_6103 (I110543,I691,I110093,I110570,);
nor I_6104 (I110579,I110192,I110507);
nor I_6105 (I110597,I110408,I110579);
nor I_6106 (I110615,I110336,I110489);
nor I_6107 (I110633,I110192,I110489);
not I_6108 (I110651,I698);
DFFARX1 I_6109 (I110633,I691,I110651,I110678,);
not I_6110 (I110687,I110678);
nand I_6111 (I110705,I110309,I110354);
and I_6112 (I110723,I110705,I110264);
DFFARX1 I_6113 (I110723,I691,I110651,I110750,);
not I_6114 (I110759,I110633);
DFFARX1 I_6115 (I110570,I691,I110651,I110786,);
not I_6116 (I110795,I110786);
nor I_6117 (I110813,I110795,I110687);
and I_6118 (I110831,I110813,I110633);
nor I_6119 (I110849,I110795,I110759);
nor I_6120 (I110867,I110750,I110849);
DFFARX1 I_6121 (I110471,I691,I110651,I110894,);
nor I_6122 (I110903,I110894,I110750);
not I_6123 (I110921,I110903);
not I_6124 (I110939,I110894);
nor I_6125 (I110957,I110939,I110831);
DFFARX1 I_6126 (I110957,I691,I110651,I110984,);
nand I_6127 (I110993,I110435,I110264);
and I_6128 (I111011,I110993,I110597);
DFFARX1 I_6129 (I111011,I691,I110651,I111038,);
nor I_6130 (I111047,I111038,I110894);
DFFARX1 I_6131 (I111047,I691,I110651,I111074,);
nand I_6132 (I111083,I111038,I110939);
nand I_6133 (I111101,I110921,I111083);
not I_6134 (I111119,I111038);
nor I_6135 (I111137,I111119,I110831);
DFFARX1 I_6136 (I111137,I691,I110651,I111164,);
nor I_6137 (I111173,I110615,I110264);
or I_6138 (I111191,I110894,I111173);
nor I_6139 (I111209,I111038,I111173);
or I_6140 (I111227,I110750,I111173);
DFFARX1 I_6141 (I111173,I691,I110651,I111254,);
not I_6142 (I111263,I698);
DFFARX1 I_6143 (I110867,I691,I111263,I111290,);
and I_6144 (I111299,I111290,I111209);
DFFARX1 I_6145 (I111299,I691,I111263,I111326,);
DFFARX1 I_6146 (I111227,I691,I111263,I111344,);
not I_6147 (I111353,I111074);
not I_6148 (I111371,I111254);
nand I_6149 (I111389,I111371,I111353);
nor I_6150 (I111407,I111344,I111389);
DFFARX1 I_6151 (I111389,I691,I111263,I111434,);
not I_6152 (I111443,I111434);
not I_6153 (I111461,I111191);
nand I_6154 (I111479,I111371,I111461);
DFFARX1 I_6155 (I111479,I691,I111263,I111506,);
not I_6156 (I111515,I111506);
not I_6157 (I111533,I111164);
nand I_6158 (I111551,I111533,I110984);
and I_6159 (I111569,I111353,I111551);
nor I_6160 (I111587,I111479,I111569);
DFFARX1 I_6161 (I111587,I691,I111263,I111614,);
DFFARX1 I_6162 (I111569,I691,I111263,I111632,);
nor I_6163 (I111641,I111164,I111101);
nor I_6164 (I111659,I111479,I111641);
or I_6165 (I111677,I111164,I111101);
nor I_6166 (I111695,I111074,I111209);
DFFARX1 I_6167 (I111695,I691,I111263,I111722,);
not I_6168 (I111731,I111722);
nor I_6169 (I111749,I111731,I111515);
nand I_6170 (I111767,I111731,I111344);
not I_6171 (I111785,I111074);
nand I_6172 (I111803,I111785,I111461);
nand I_6173 (I111821,I111731,I111803);
nand I_6174 (I111839,I111821,I111767);
nand I_6175 (I111857,I111803,I111677);
not I_6176 (I111875,I698);
DFFARX1 I_6177 (I111407,I691,I111875,I111902,);
DFFARX1 I_6178 (I111902,I691,I111875,I111920,);
not I_6179 (I111929,I111920);
not I_6180 (I111947,I111902);
nand I_6181 (I111965,I111326,I111407);
and I_6182 (I111983,I111965,I111857);
DFFARX1 I_6183 (I111983,I691,I111875,I112010,);
not I_6184 (I112019,I112010);
DFFARX1 I_6185 (I111443,I691,I111875,I112046,);
and I_6186 (I112055,I112046,I111614);
nand I_6187 (I112073,I112046,I111614);
nand I_6188 (I112091,I112019,I112073);
DFFARX1 I_6189 (I111749,I691,I111875,I112118,);
nor I_6190 (I112127,I112118,I112055);
DFFARX1 I_6191 (I112127,I691,I111875,I112154,);
nor I_6192 (I112163,I112118,I112010);
nand I_6193 (I112181,I111659,I111839);
and I_6194 (I112199,I112181,I111632);
DFFARX1 I_6195 (I112199,I691,I111875,I112226,);
nor I_6196 (I112235,I112226,I112118);
not I_6197 (I112253,I112226);
nor I_6198 (I112271,I112253,I112019);
nor I_6199 (I112289,I111947,I112271);
DFFARX1 I_6200 (I112289,I691,I111875,I112316,);
nor I_6201 (I112325,I112253,I112118);
nor I_6202 (I112343,I111614,I111839);
nor I_6203 (I112361,I112343,I112325);
not I_6204 (I112379,I112343);
nand I_6205 (I112397,I112073,I112379);
DFFARX1 I_6206 (I112343,I691,I111875,I112424,);
DFFARX1 I_6207 (I112343,I691,I111875,I112442,);
not I_6208 (I112451,I698);
DFFARX1 I_6209 (I112397,I691,I112451,I112478,);
nand I_6210 (I112487,I112424,I112235);
and I_6211 (I112505,I112487,I111929);
DFFARX1 I_6212 (I112505,I691,I112451,I112532,);
nor I_6213 (I112541,I112532,I112478);
not I_6214 (I112559,I112532);
DFFARX1 I_6215 (I112316,I691,I112451,I112586,);
nand I_6216 (I112595,I112586,I112154);
not I_6217 (I112613,I112595);
DFFARX1 I_6218 (I112613,I691,I112451,I112640,);
not I_6219 (I112649,I112640);
nor I_6220 (I112667,I112478,I112595);
nor I_6221 (I112685,I112532,I112667);
DFFARX1 I_6222 (I112163,I691,I112451,I112712,);
DFFARX1 I_6223 (I112712,I691,I112451,I112730,);
not I_6224 (I112739,I112730);
not I_6225 (I112757,I112712);
nand I_6226 (I112775,I112757,I112559);
nand I_6227 (I112793,I112154,I112091);
and I_6228 (I112811,I112793,I112361);
DFFARX1 I_6229 (I112811,I691,I112451,I112838,);
nor I_6230 (I112847,I112838,I112478);
DFFARX1 I_6231 (I112847,I691,I112451,I112874,);
DFFARX1 I_6232 (I112838,I691,I112451,I112892,);
nor I_6233 (I112901,I112442,I112091);
not I_6234 (I112919,I112901);
nor I_6235 (I112937,I112739,I112919);
nand I_6236 (I112955,I112757,I112919);
nor I_6237 (I112973,I112478,I112901);
DFFARX1 I_6238 (I112901,I691,I112451,I113000,);
not I_6239 (I113009,I698);
DFFARX1 I_6240 (I112955,I691,I113009,I113036,);
not I_6241 (I113045,I113036);
DFFARX1 I_6242 (I112937,I691,I113009,I113072,);
not I_6243 (I113081,I113000);
nand I_6244 (I113099,I113081,I112541);
not I_6245 (I113117,I113099);
nor I_6246 (I113135,I113117,I112649);
nor I_6247 (I113153,I113045,I113135);
DFFARX1 I_6248 (I113153,I691,I113009,I113180,);
not I_6249 (I113189,I112649);
nand I_6250 (I113207,I113189,I113117);
and I_6251 (I113225,I113189,I112685);
nand I_6252 (I113243,I113225,I112874);
nor I_6253 (I113261,I113243,I113189);
and I_6254 (I113279,I113072,I113243);
not I_6255 (I113297,I113243);
nand I_6256 (I113315,I113072,I113297);
nor I_6257 (I113333,I113036,I113243);
not I_6258 (I113351,I112874);
nor I_6259 (I113369,I113351,I112685);
nand I_6260 (I113387,I113369,I113189);
nor I_6261 (I113405,I113099,I113387);
nor I_6262 (I113423,I113351,I112973);
and I_6263 (I113441,I113423,I112892);
or I_6264 (I113459,I113441,I112775);
DFFARX1 I_6265 (I113459,I691,I113009,I113486,);
nor I_6266 (I113495,I113486,I113207);
DFFARX1 I_6267 (I113495,I691,I113009,I113522,);
DFFARX1 I_6268 (I113486,I691,I113009,I113540,);
not I_6269 (I113549,I113486);
nor I_6270 (I113567,I113549,I113072);
nor I_6271 (I113585,I113369,I113567);
DFFARX1 I_6272 (I113585,I691,I113009,I113612,);
not I_6273 (I113621,I698);
DFFARX1 I_6274 (I113261,I691,I113621,I113648,);
and I_6275 (I113657,I113648,I113333);
DFFARX1 I_6276 (I113657,I691,I113621,I113684,);
DFFARX1 I_6277 (I113180,I691,I113621,I113702,);
not I_6278 (I113711,I113315);
not I_6279 (I113729,I113522);
nand I_6280 (I113747,I113729,I113711);
nor I_6281 (I113765,I113702,I113747);
DFFARX1 I_6282 (I113747,I691,I113621,I113792,);
not I_6283 (I113801,I113792);
not I_6284 (I113819,I113279);
nand I_6285 (I113837,I113729,I113819);
DFFARX1 I_6286 (I113837,I691,I113621,I113864,);
not I_6287 (I113873,I113864);
not I_6288 (I113891,I113612);
nand I_6289 (I113909,I113891,I113540);
and I_6290 (I113927,I113711,I113909);
nor I_6291 (I113945,I113837,I113927);
DFFARX1 I_6292 (I113945,I691,I113621,I113972,);
DFFARX1 I_6293 (I113927,I691,I113621,I113990,);
nor I_6294 (I113999,I113612,I113522);
nor I_6295 (I114017,I113837,I113999);
or I_6296 (I114035,I113612,I113522);
nor I_6297 (I114053,I113405,I113333);
DFFARX1 I_6298 (I114053,I691,I113621,I114080,);
not I_6299 (I114089,I114080);
nor I_6300 (I114107,I114089,I113873);
nand I_6301 (I114125,I114089,I113702);
not I_6302 (I114143,I113405);
nand I_6303 (I114161,I114143,I113819);
nand I_6304 (I114179,I114089,I114161);
nand I_6305 (I114197,I114179,I114125);
nand I_6306 (I114215,I114161,I114035);
not I_6307 (I114233,I698);
DFFARX1 I_6308 (I114107,I691,I114233,I114260,);
DFFARX1 I_6309 (I113972,I691,I114233,I114278,);
not I_6310 (I114287,I114278);
not I_6311 (I114305,I114197);
nor I_6312 (I114323,I114305,I113990);
not I_6313 (I114341,I113765);
nor I_6314 (I114359,I114323,I114017);
nor I_6315 (I114377,I114278,I114359);
DFFARX1 I_6316 (I114377,I691,I114233,I114404,);
nor I_6317 (I114413,I114017,I113990);
nand I_6318 (I114431,I114413,I114197);
DFFARX1 I_6319 (I114431,I691,I114233,I114458,);
nor I_6320 (I114467,I114341,I114017);
nand I_6321 (I114485,I114467,I113801);
nor I_6322 (I114503,I114260,I114485);
DFFARX1 I_6323 (I114503,I691,I114233,I114530,);
not I_6324 (I114539,I114485);
nand I_6325 (I114557,I114278,I114539);
DFFARX1 I_6326 (I114485,I691,I114233,I114584,);
not I_6327 (I114593,I114584);
not I_6328 (I114611,I114017);
not I_6329 (I114629,I113972);
nor I_6330 (I114647,I114629,I113765);
nor I_6331 (I114665,I114593,I114647);
nor I_6332 (I114683,I114629,I114215);
and I_6333 (I114701,I114683,I113684);
or I_6334 (I114719,I114701,I113765);
DFFARX1 I_6335 (I114719,I691,I114233,I114746,);
nor I_6336 (I114755,I114746,I114260);
not I_6337 (I114773,I114746);
and I_6338 (I114791,I114773,I114260);
nor I_6339 (I114809,I114287,I114791);
nand I_6340 (I114827,I114773,I114341);
nor I_6341 (I114845,I114629,I114827);
nand I_6342 (I114863,I114773,I114539);
nand I_6343 (I114881,I114341,I113972);
nor I_6344 (I114899,I114611,I114881);
not I_6345 (I114917,I698);
DFFARX1 I_6346 (I114845,I691,I114917,I114944,);
not I_6347 (I114953,I114944);
nand I_6348 (I114971,I114899,I114530);
and I_6349 (I114989,I114971,I114530);
DFFARX1 I_6350 (I114989,I691,I114917,I115016,);
DFFARX1 I_6351 (I115016,I691,I114917,I115034,);
DFFARX1 I_6352 (I114809,I691,I114917,I115052,);
nand I_6353 (I115061,I115052,I114665);
not I_6354 (I115079,I115061);
DFFARX1 I_6355 (I115079,I691,I114917,I115106,);
not I_6356 (I115115,I115106);
nor I_6357 (I115133,I114953,I115115);
DFFARX1 I_6358 (I114458,I691,I114917,I115160,);
nor I_6359 (I115169,I115160,I115016);
nor I_6360 (I115187,I115160,I115079);
nand I_6361 (I115205,I114404,I114557);
and I_6362 (I115223,I115205,I114863);
DFFARX1 I_6363 (I115223,I691,I114917,I115250,);
not I_6364 (I115259,I115250);
nand I_6365 (I115277,I115259,I115160);
nand I_6366 (I115295,I115259,I115061);
nor I_6367 (I115313,I114755,I114557);
and I_6368 (I115331,I115160,I115313);
nor I_6369 (I115349,I115259,I115331);
DFFARX1 I_6370 (I115349,I691,I114917,I115376,);
nor I_6371 (I115385,I114944,I115313);
DFFARX1 I_6372 (I115385,I691,I114917,I115412,);
nor I_6373 (I115421,I115250,I115313);
not I_6374 (I115439,I115421);
nand I_6375 (I115457,I115439,I115277);
not I_6376 (I115475,I698);
DFFARX1 I_6377 (I115187,I691,I115475,I115502,);
and I_6378 (I115511,I115502,I115457);
DFFARX1 I_6379 (I115511,I691,I115475,I115538,);
DFFARX1 I_6380 (I115376,I691,I115475,I115556,);
not I_6381 (I115565,I115412);
not I_6382 (I115583,I115412);
nand I_6383 (I115601,I115583,I115565);
nor I_6384 (I115619,I115556,I115601);
DFFARX1 I_6385 (I115601,I691,I115475,I115646,);
not I_6386 (I115655,I115646);
not I_6387 (I115673,I115034);
nand I_6388 (I115691,I115583,I115673);
DFFARX1 I_6389 (I115691,I691,I115475,I115718,);
not I_6390 (I115727,I115718);
not I_6391 (I115745,I115169);
nand I_6392 (I115763,I115745,I115187);
and I_6393 (I115781,I115565,I115763);
nor I_6394 (I115799,I115691,I115781);
DFFARX1 I_6395 (I115799,I691,I115475,I115826,);
DFFARX1 I_6396 (I115781,I691,I115475,I115844,);
nor I_6397 (I115853,I115169,I115133);
nor I_6398 (I115871,I115691,I115853);
or I_6399 (I115889,I115169,I115133);
nor I_6400 (I115907,I115295,I115295);
DFFARX1 I_6401 (I115907,I691,I115475,I115934,);
not I_6402 (I115943,I115934);
nor I_6403 (I115961,I115943,I115727);
nand I_6404 (I115979,I115943,I115556);
not I_6405 (I115997,I115295);
nand I_6406 (I116015,I115997,I115673);
nand I_6407 (I116033,I115943,I116015);
nand I_6408 (I116051,I116033,I115979);
nand I_6409 (I116069,I116015,I115889);
not I_6410 (I116087,I698);
DFFARX1 I_6411 (I115961,I691,I116087,I116114,);
nand I_6412 (I116123,I116114,I115619);
not I_6413 (I116141,I116123);
DFFARX1 I_6414 (I116069,I691,I116087,I116168,);
not I_6415 (I116177,I116168);
not I_6416 (I116195,I115844);
or I_6417 (I116213,I115655,I115844);
nor I_6418 (I116231,I115655,I115844);
or I_6419 (I116249,I115826,I115655);
DFFARX1 I_6420 (I116249,I691,I116087,I116276,);
not I_6421 (I116285,I115871);
nand I_6422 (I116303,I116285,I115538);
nand I_6423 (I116321,I116195,I116303);
and I_6424 (I116339,I116177,I116321);
nor I_6425 (I116357,I115871,I116051);
and I_6426 (I116375,I116177,I116357);
nor I_6427 (I116393,I116141,I116375);
DFFARX1 I_6428 (I116357,I691,I116087,I116420,);
not I_6429 (I116429,I116420);
nor I_6430 (I116447,I116177,I116429);
or I_6431 (I116465,I116249,I115826);
nor I_6432 (I116483,I115826,I115826);
nand I_6433 (I116501,I116321,I116483);
nand I_6434 (I116519,I116465,I116501);
DFFARX1 I_6435 (I116519,I691,I116087,I116546,);
nor I_6436 (I116555,I116483,I116213);
DFFARX1 I_6437 (I116555,I691,I116087,I116582,);
nor I_6438 (I116591,I115826,I115619);
DFFARX1 I_6439 (I116591,I691,I116087,I116618,);
DFFARX1 I_6440 (I116618,I691,I116087,I116636,);
not I_6441 (I116645,I116618);
nand I_6442 (I116663,I116645,I116123);
nand I_6443 (I116681,I116645,I116231);
not I_6444 (I116699,I698);
DFFARX1 I_6445 (I116546,I691,I116699,I116726,);
not I_6446 (I116735,I116726);
nand I_6447 (I116753,I116276,I116447);
and I_6448 (I116771,I116753,I116636);
DFFARX1 I_6449 (I116771,I691,I116699,I116798,);
DFFARX1 I_6450 (I116582,I691,I116699,I116816,);
and I_6451 (I116825,I116816,I116393);
nor I_6452 (I116843,I116798,I116825);
DFFARX1 I_6453 (I116843,I691,I116699,I116870,);
nand I_6454 (I116879,I116816,I116393);
nand I_6455 (I116897,I116735,I116879);
not I_6456 (I116915,I116897);
DFFARX1 I_6457 (I116582,I691,I116699,I116942,);
DFFARX1 I_6458 (I116942,I691,I116699,I116960,);
nand I_6459 (I116969,I116339,I116681);
and I_6460 (I116987,I116969,I116663);
DFFARX1 I_6461 (I116987,I691,I116699,I117014,);
DFFARX1 I_6462 (I117014,I691,I116699,I117032,);
not I_6463 (I117041,I117032);
not I_6464 (I117059,I117014);
nand I_6465 (I117077,I117059,I116879);
nor I_6466 (I117095,I116339,I116681);
not I_6467 (I117113,I117095);
nor I_6468 (I117131,I117059,I117113);
nor I_6469 (I117149,I116735,I117131);
DFFARX1 I_6470 (I117149,I691,I116699,I117176,);
nor I_6471 (I117185,I116798,I117113);
nor I_6472 (I117203,I117014,I117185);
nor I_6473 (I117221,I116942,I117095);
nor I_6474 (I117239,I116798,I117095);
not I_6475 (I117257,I698);
DFFARX1 I_6476 (I117041,I691,I117257,I117284,);
not I_6477 (I117293,I117284);
nand I_6478 (I117311,I116870,I117077);
and I_6479 (I117329,I117311,I117239);
DFFARX1 I_6480 (I117329,I691,I117257,I117356,);
DFFARX1 I_6481 (I117356,I691,I117257,I117374,);
DFFARX1 I_6482 (I116960,I691,I117257,I117392,);
nand I_6483 (I117401,I117392,I116915);
not I_6484 (I117419,I117401);
DFFARX1 I_6485 (I117419,I691,I117257,I117446,);
not I_6486 (I117455,I117446);
nor I_6487 (I117473,I117293,I117455);
DFFARX1 I_6488 (I117203,I691,I117257,I117500,);
nor I_6489 (I117509,I117500,I117356);
nor I_6490 (I117527,I117500,I117419);
nand I_6491 (I117545,I117176,I117221);
and I_6492 (I117563,I117545,I117239);
DFFARX1 I_6493 (I117563,I691,I117257,I117590,);
not I_6494 (I117599,I117590);
nand I_6495 (I117617,I117599,I117500);
nand I_6496 (I117635,I117599,I117401);
nor I_6497 (I117653,I116870,I117221);
and I_6498 (I117671,I117500,I117653);
nor I_6499 (I117689,I117599,I117671);
DFFARX1 I_6500 (I117689,I691,I117257,I117716,);
nor I_6501 (I117725,I117284,I117653);
DFFARX1 I_6502 (I117725,I691,I117257,I117752,);
nor I_6503 (I117761,I117590,I117653);
not I_6504 (I117779,I117761);
nand I_6505 (I117797,I117779,I117617);
not I_6506 (I117815,I698);
DFFARX1 I_6507 (I117527,I691,I117815,I117842,);
and I_6508 (I117851,I117842,I117797);
DFFARX1 I_6509 (I117851,I691,I117815,I117878,);
DFFARX1 I_6510 (I117716,I691,I117815,I117896,);
not I_6511 (I117905,I117752);
not I_6512 (I117923,I117752);
nand I_6513 (I117941,I117923,I117905);
nor I_6514 (I117959,I117896,I117941);
DFFARX1 I_6515 (I117941,I691,I117815,I117986,);
not I_6516 (I117995,I117986);
not I_6517 (I118013,I117374);
nand I_6518 (I118031,I117923,I118013);
DFFARX1 I_6519 (I118031,I691,I117815,I118058,);
not I_6520 (I118067,I118058);
not I_6521 (I118085,I117509);
nand I_6522 (I118103,I118085,I117527);
and I_6523 (I118121,I117905,I118103);
nor I_6524 (I118139,I118031,I118121);
DFFARX1 I_6525 (I118139,I691,I117815,I118166,);
DFFARX1 I_6526 (I118121,I691,I117815,I118184,);
nor I_6527 (I118193,I117509,I117473);
nor I_6528 (I118211,I118031,I118193);
or I_6529 (I118229,I117509,I117473);
nor I_6530 (I118247,I117635,I117635);
DFFARX1 I_6531 (I118247,I691,I117815,I118274,);
not I_6532 (I118283,I118274);
nor I_6533 (I118301,I118283,I118067);
nand I_6534 (I118319,I118283,I117896);
not I_6535 (I118337,I117635);
nand I_6536 (I118355,I118337,I118013);
nand I_6537 (I118373,I118283,I118355);
nand I_6538 (I118391,I118373,I118319);
nand I_6539 (I118409,I118355,I118229);
not I_6540 (I118427,I698);
DFFARX1 I_6541 (I124,I691,I118427,I118454,);
DFFARX1 I_6542 (I118454,I691,I118427,I118472,);
not I_6543 (I118481,I118472);
nand I_6544 (I118499,I660,I420);
and I_6545 (I118517,I118499,I564);
DFFARX1 I_6546 (I118517,I691,I118427,I118544,);
DFFARX1 I_6547 (I118544,I691,I118427,I118562,);
DFFARX1 I_6548 (I118544,I691,I118427,I118580,);
DFFARX1 I_6549 (I396,I691,I118427,I118598,);
nand I_6550 (I118607,I118598,I676);
not I_6551 (I118625,I118607);
nor I_6552 (I118643,I118454,I118625);
DFFARX1 I_6553 (I340,I691,I118427,I118670,);
not I_6554 (I118679,I118670);
nor I_6555 (I118697,I118679,I118481);
nand I_6556 (I118715,I118679,I118607);
nand I_6557 (I118733,I388,I140);
and I_6558 (I118751,I118733,I244);
DFFARX1 I_6559 (I118751,I691,I118427,I118778,);
nor I_6560 (I118787,I118778,I118454);
DFFARX1 I_6561 (I118787,I691,I118427,I118814,);
not I_6562 (I118823,I118778);
nor I_6563 (I118841,I308,I140);
not I_6564 (I118859,I118841);
nor I_6565 (I118877,I118607,I118859);
nor I_6566 (I118895,I118823,I118877);
DFFARX1 I_6567 (I118895,I691,I118427,I118922,);
nor I_6568 (I118931,I118778,I118859);
nor I_6569 (I118949,I118625,I118931);
nor I_6570 (I118967,I118778,I118841);
not I_6571 (I118985,I698);
DFFARX1 I_6572 (I118643,I691,I118985,I119012,);
DFFARX1 I_6573 (I119012,I691,I118985,I119030,);
not I_6574 (I119039,I119030);
not I_6575 (I119057,I119012);
nand I_6576 (I119075,I118814,I118580);
and I_6577 (I119093,I119075,I118967);
DFFARX1 I_6578 (I119093,I691,I118985,I119120,);
not I_6579 (I119129,I119120);
DFFARX1 I_6580 (I118562,I691,I118985,I119156,);
and I_6581 (I119165,I119156,I118697);
nand I_6582 (I119183,I119156,I118697);
nand I_6583 (I119201,I119129,I119183);
DFFARX1 I_6584 (I118922,I691,I118985,I119228,);
nor I_6585 (I119237,I119228,I119165);
DFFARX1 I_6586 (I119237,I691,I118985,I119264,);
nor I_6587 (I119273,I119228,I119120);
nand I_6588 (I119291,I118814,I118967);
and I_6589 (I119309,I119291,I118715);
DFFARX1 I_6590 (I119309,I691,I118985,I119336,);
nor I_6591 (I119345,I119336,I119228);
not I_6592 (I119363,I119336);
nor I_6593 (I119381,I119363,I119129);
nor I_6594 (I119399,I119057,I119381);
DFFARX1 I_6595 (I119399,I691,I118985,I119426,);
nor I_6596 (I119435,I119363,I119228);
nor I_6597 (I119453,I118949,I118967);
nor I_6598 (I119471,I119453,I119435);
not I_6599 (I119489,I119453);
nand I_6600 (I119507,I119183,I119489);
DFFARX1 I_6601 (I119453,I691,I118985,I119534,);
DFFARX1 I_6602 (I119453,I691,I118985,I119552,);
not I_6603 (I119561,I698);
DFFARX1 I_6604 (I119471,I691,I119561,I119588,);
not I_6605 (I119597,I119588);
nand I_6606 (I119615,I119264,I119426);
and I_6607 (I119633,I119615,I119552);
DFFARX1 I_6608 (I119633,I691,I119561,I119660,);
not I_6609 (I119669,I119273);
DFFARX1 I_6610 (I119345,I691,I119561,I119696,);
not I_6611 (I119705,I119696);
nor I_6612 (I119723,I119705,I119597);
and I_6613 (I119741,I119723,I119273);
nor I_6614 (I119759,I119705,I119669);
nor I_6615 (I119777,I119660,I119759);
DFFARX1 I_6616 (I119507,I691,I119561,I119804,);
nor I_6617 (I119813,I119804,I119660);
not I_6618 (I119831,I119813);
not I_6619 (I119849,I119804);
nor I_6620 (I119867,I119849,I119741);
DFFARX1 I_6621 (I119867,I691,I119561,I119894,);
nand I_6622 (I119903,I119039,I119534);
and I_6623 (I119921,I119903,I119201);
DFFARX1 I_6624 (I119921,I691,I119561,I119948,);
nor I_6625 (I119957,I119948,I119804);
DFFARX1 I_6626 (I119957,I691,I119561,I119984,);
nand I_6627 (I119993,I119948,I119849);
nand I_6628 (I120011,I119831,I119993);
not I_6629 (I120029,I119948);
nor I_6630 (I120047,I120029,I119741);
DFFARX1 I_6631 (I120047,I691,I119561,I120074,);
nor I_6632 (I120083,I119264,I119534);
or I_6633 (I120101,I119804,I120083);
nor I_6634 (I120119,I119948,I120083);
or I_6635 (I120137,I119660,I120083);
DFFARX1 I_6636 (I120083,I691,I119561,I120164,);
not I_6637 (I120173,I698);
DFFARX1 I_6638 (I120119,I691,I120173,I120200,);
DFFARX1 I_6639 (I120200,I691,I120173,I120218,);
not I_6640 (I120227,I120218);
not I_6641 (I120245,I120200);
nand I_6642 (I120263,I120164,I119777);
and I_6643 (I120281,I120263,I120119);
DFFARX1 I_6644 (I120281,I691,I120173,I120308,);
not I_6645 (I120317,I120308);
DFFARX1 I_6646 (I120011,I691,I120173,I120344,);
and I_6647 (I120353,I120344,I120137);
nand I_6648 (I120371,I120344,I120137);
nand I_6649 (I120389,I120317,I120371);
DFFARX1 I_6650 (I119984,I691,I120173,I120416,);
nor I_6651 (I120425,I120416,I120353);
DFFARX1 I_6652 (I120425,I691,I120173,I120452,);
nor I_6653 (I120461,I120416,I120308);
nand I_6654 (I120479,I119984,I120101);
and I_6655 (I120497,I120479,I120074);
DFFARX1 I_6656 (I120497,I691,I120173,I120524,);
nor I_6657 (I120533,I120524,I120416);
not I_6658 (I120551,I120524);
nor I_6659 (I120569,I120551,I120317);
nor I_6660 (I120587,I120245,I120569);
DFFARX1 I_6661 (I120587,I691,I120173,I120614,);
nor I_6662 (I120623,I120551,I120416);
nor I_6663 (I120641,I119894,I120101);
nor I_6664 (I120659,I120641,I120623);
not I_6665 (I120677,I120641);
nand I_6666 (I120695,I120371,I120677);
DFFARX1 I_6667 (I120641,I691,I120173,I120722,);
DFFARX1 I_6668 (I120641,I691,I120173,I120740,);
not I_6669 (I120749,I698);
DFFARX1 I_6670 (I120614,I691,I120749,I120776,);
not I_6671 (I120785,I120776);
nand I_6672 (I120803,I120695,I120533);
and I_6673 (I120821,I120803,I120722);
DFFARX1 I_6674 (I120821,I691,I120749,I120848,);
DFFARX1 I_6675 (I120389,I691,I120749,I120866,);
and I_6676 (I120875,I120866,I120452);
nor I_6677 (I120893,I120848,I120875);
DFFARX1 I_6678 (I120893,I691,I120749,I120920,);
nand I_6679 (I120929,I120866,I120452);
nand I_6680 (I120947,I120785,I120929);
not I_6681 (I120965,I120947);
DFFARX1 I_6682 (I120452,I691,I120749,I120992,);
DFFARX1 I_6683 (I120992,I691,I120749,I121010,);
nand I_6684 (I121019,I120227,I120659);
and I_6685 (I121037,I121019,I120461);
DFFARX1 I_6686 (I121037,I691,I120749,I121064,);
DFFARX1 I_6687 (I121064,I691,I120749,I121082,);
not I_6688 (I121091,I121082);
not I_6689 (I121109,I121064);
nand I_6690 (I121127,I121109,I120929);
nor I_6691 (I121145,I120740,I120659);
not I_6692 (I121163,I121145);
nor I_6693 (I121181,I121109,I121163);
nor I_6694 (I121199,I120785,I121181);
DFFARX1 I_6695 (I121199,I691,I120749,I121226,);
nor I_6696 (I121235,I120848,I121163);
nor I_6697 (I121253,I121064,I121235);
nor I_6698 (I121271,I120992,I121145);
nor I_6699 (I121289,I120848,I121145);
not I_6700 (I121307,I698);
DFFARX1 I_6701 (I121289,I691,I121307,I121334,);
nand I_6702 (I121343,I121271,I121091);
and I_6703 (I121361,I121343,I121289);
DFFARX1 I_6704 (I121361,I691,I121307,I121388,);
nor I_6705 (I121397,I121388,I121334);
not I_6706 (I121415,I121388);
DFFARX1 I_6707 (I121226,I691,I121307,I121442,);
nand I_6708 (I121451,I121442,I121253);
not I_6709 (I121469,I121451);
DFFARX1 I_6710 (I121469,I691,I121307,I121496,);
not I_6711 (I121505,I121496);
nor I_6712 (I121523,I121334,I121451);
nor I_6713 (I121541,I121388,I121523);
DFFARX1 I_6714 (I121127,I691,I121307,I121568,);
DFFARX1 I_6715 (I121568,I691,I121307,I121586,);
not I_6716 (I121595,I121586);
not I_6717 (I121613,I121568);
nand I_6718 (I121631,I121613,I121415);
nand I_6719 (I121649,I120920,I120920);
and I_6720 (I121667,I121649,I120965);
DFFARX1 I_6721 (I121667,I691,I121307,I121694,);
nor I_6722 (I121703,I121694,I121334);
DFFARX1 I_6723 (I121703,I691,I121307,I121730,);
DFFARX1 I_6724 (I121694,I691,I121307,I121748,);
nor I_6725 (I121757,I121010,I120920);
not I_6726 (I121775,I121757);
nor I_6727 (I121793,I121595,I121775);
nand I_6728 (I121811,I121613,I121775);
nor I_6729 (I121829,I121334,I121757);
DFFARX1 I_6730 (I121757,I691,I121307,I121856,);
not I_6731 (I121865,I698);
DFFARX1 I_6732 (I121505,I691,I121865,I121892,);
and I_6733 (I121901,I121892,I121631);
DFFARX1 I_6734 (I121901,I691,I121865,I121928,);
DFFARX1 I_6735 (I121748,I691,I121865,I121946,);
not I_6736 (I121955,I121730);
not I_6737 (I121973,I121793);
nand I_6738 (I121991,I121973,I121955);
nor I_6739 (I122009,I121946,I121991);
DFFARX1 I_6740 (I121991,I691,I121865,I122036,);
not I_6741 (I122045,I122036);
not I_6742 (I122063,I121856);
nand I_6743 (I122081,I121973,I122063);
DFFARX1 I_6744 (I122081,I691,I121865,I122108,);
not I_6745 (I122117,I122108);
not I_6746 (I122135,I121829);
nand I_6747 (I122153,I122135,I121397);
and I_6748 (I122171,I121955,I122153);
nor I_6749 (I122189,I122081,I122171);
DFFARX1 I_6750 (I122189,I691,I121865,I122216,);
DFFARX1 I_6751 (I122171,I691,I121865,I122234,);
nor I_6752 (I122243,I121829,I121541);
nor I_6753 (I122261,I122081,I122243);
or I_6754 (I122279,I121829,I121541);
nor I_6755 (I122297,I121811,I121730);
DFFARX1 I_6756 (I122297,I691,I121865,I122324,);
not I_6757 (I122333,I122324);
nor I_6758 (I122351,I122333,I122117);
nand I_6759 (I122369,I122333,I121946);
not I_6760 (I122387,I121811);
nand I_6761 (I122405,I122387,I122063);
nand I_6762 (I122423,I122333,I122405);
nand I_6763 (I122441,I122423,I122369);
nand I_6764 (I122459,I122405,I122279);
not I_6765 (I122477,I698);
DFFARX1 I_6766 (I122009,I691,I122477,I122504,);
DFFARX1 I_6767 (I122504,I691,I122477,I122522,);
not I_6768 (I122531,I122522);
not I_6769 (I122549,I122504);
nand I_6770 (I122567,I121928,I122009);
and I_6771 (I122585,I122567,I122459);
DFFARX1 I_6772 (I122585,I691,I122477,I122612,);
not I_6773 (I122621,I122612);
DFFARX1 I_6774 (I122045,I691,I122477,I122648,);
and I_6775 (I122657,I122648,I122216);
nand I_6776 (I122675,I122648,I122216);
nand I_6777 (I122693,I122621,I122675);
DFFARX1 I_6778 (I122351,I691,I122477,I122720,);
nor I_6779 (I122729,I122720,I122657);
DFFARX1 I_6780 (I122729,I691,I122477,I122756,);
nor I_6781 (I122765,I122720,I122612);
nand I_6782 (I122783,I122261,I122441);
and I_6783 (I122801,I122783,I122234);
DFFARX1 I_6784 (I122801,I691,I122477,I122828,);
nor I_6785 (I122837,I122828,I122720);
not I_6786 (I122855,I122828);
nor I_6787 (I122873,I122855,I122621);
nor I_6788 (I122891,I122549,I122873);
DFFARX1 I_6789 (I122891,I691,I122477,I122918,);
nor I_6790 (I122927,I122855,I122720);
nor I_6791 (I122945,I122216,I122441);
nor I_6792 (I122963,I122945,I122927);
not I_6793 (I122981,I122945);
nand I_6794 (I122999,I122675,I122981);
DFFARX1 I_6795 (I122945,I691,I122477,I123026,);
DFFARX1 I_6796 (I122945,I691,I122477,I123044,);
not I_6797 (I123053,I698);
DFFARX1 I_6798 (I122963,I691,I123053,I123080,);
not I_6799 (I123089,I123080);
nand I_6800 (I123107,I122756,I122918);
and I_6801 (I123125,I123107,I123044);
DFFARX1 I_6802 (I123125,I691,I123053,I123152,);
not I_6803 (I123161,I122765);
DFFARX1 I_6804 (I122837,I691,I123053,I123188,);
not I_6805 (I123197,I123188);
nor I_6806 (I123215,I123197,I123089);
and I_6807 (I123233,I123215,I122765);
nor I_6808 (I123251,I123197,I123161);
nor I_6809 (I123269,I123152,I123251);
DFFARX1 I_6810 (I122999,I691,I123053,I123296,);
nor I_6811 (I123305,I123296,I123152);
not I_6812 (I123323,I123305);
not I_6813 (I123341,I123296);
nor I_6814 (I123359,I123341,I123233);
DFFARX1 I_6815 (I123359,I691,I123053,I123386,);
nand I_6816 (I123395,I122531,I123026);
and I_6817 (I123413,I123395,I122693);
DFFARX1 I_6818 (I123413,I691,I123053,I123440,);
nor I_6819 (I123449,I123440,I123296);
DFFARX1 I_6820 (I123449,I691,I123053,I123476,);
nand I_6821 (I123485,I123440,I123341);
nand I_6822 (I123503,I123323,I123485);
not I_6823 (I123521,I123440);
nor I_6824 (I123539,I123521,I123233);
DFFARX1 I_6825 (I123539,I691,I123053,I123566,);
nor I_6826 (I123575,I122756,I123026);
or I_6827 (I123593,I123296,I123575);
nor I_6828 (I123611,I123440,I123575);
or I_6829 (I123629,I123152,I123575);
DFFARX1 I_6830 (I123575,I691,I123053,I123656,);
not I_6831 (I123665,I698);
DFFARX1 I_6832 (I123476,I691,I123665,I123692,);
not I_6833 (I123701,I123692);
DFFARX1 I_6834 (I123566,I691,I123665,I123728,);
not I_6835 (I123737,I123476);
or I_6836 (I123755,I123593,I123476);
nor I_6837 (I123773,I123728,I123593);
nand I_6838 (I123791,I123737,I123773);
nor I_6839 (I123809,I123503,I123593);
nand I_6840 (I123827,I123809,I123737);
not I_6841 (I123845,I123386);
nand I_6842 (I123863,I123737,I123845);
nor I_6843 (I123881,I123611,I123611);
not I_6844 (I123899,I123881);
nor I_6845 (I123917,I123899,I123863);
nor I_6846 (I123935,I123809,I123917);
DFFARX1 I_6847 (I123935,I691,I123665,I123962,);
nor I_6848 (I123971,I123881,I123755);
DFFARX1 I_6849 (I123881,I691,I123665,I123998,);
nor I_6850 (I124007,I123845,I123611);
nor I_6851 (I124025,I124007,I123476);
nor I_6852 (I124043,I123656,I123629);
DFFARX1 I_6853 (I124043,I691,I123665,I124070,);
nor I_6854 (I124079,I124070,I124025);
DFFARX1 I_6855 (I124070,I691,I123665,I124106,);
nand I_6856 (I124115,I124106,I123269);
nor I_6857 (I124133,I123701,I124115);
not I_6858 (I124151,I124070);
nand I_6859 (I124169,I124151,I123269);
nor I_6860 (I124187,I123701,I124169);
nor I_6861 (I124205,I123728,I124187);
nor I_6862 (I124223,I123656,I123503);
nor I_6863 (I124241,I123728,I124223);
DFFARX1 I_6864 (I124241,I691,I123665,I124268,);
and I_6865 (I124277,I123809,I123656);
not I_6866 (I124295,I698);
DFFARX1 I_6867 (I124277,I691,I124295,I124322,);
DFFARX1 I_6868 (I124322,I691,I124295,I124340,);
not I_6869 (I124349,I124340);
nand I_6870 (I124367,I123971,I124268);
and I_6871 (I124385,I124367,I123827);
DFFARX1 I_6872 (I124385,I691,I124295,I124412,);
DFFARX1 I_6873 (I124412,I691,I124295,I124430,);
DFFARX1 I_6874 (I124412,I691,I124295,I124448,);
DFFARX1 I_6875 (I124205,I691,I124295,I124466,);
nand I_6876 (I124475,I124466,I124268);
not I_6877 (I124493,I124475);
nor I_6878 (I124511,I124322,I124493);
DFFARX1 I_6879 (I123962,I691,I124295,I124538,);
not I_6880 (I124547,I124538);
nor I_6881 (I124565,I124547,I124349);
nand I_6882 (I124583,I124547,I124475);
nand I_6883 (I124601,I123998,I123791);
and I_6884 (I124619,I124601,I124079);
DFFARX1 I_6885 (I124619,I691,I124295,I124646,);
nor I_6886 (I124655,I124646,I124322);
DFFARX1 I_6887 (I124655,I691,I124295,I124682,);
not I_6888 (I124691,I124646);
nor I_6889 (I124709,I124133,I123791);
not I_6890 (I124727,I124709);
nor I_6891 (I124745,I124475,I124727);
nor I_6892 (I124763,I124691,I124745);
DFFARX1 I_6893 (I124763,I691,I124295,I124790,);
nor I_6894 (I124799,I124646,I124727);
nor I_6895 (I124817,I124493,I124799);
nor I_6896 (I124835,I124646,I124709);
not I_6897 (I124853,I698);
DFFARX1 I_6898 (I124682,I691,I124853,I124880,);
nand I_6899 (I124889,I124448,I124835);
and I_6900 (I124907,I124889,I124682);
DFFARX1 I_6901 (I124907,I691,I124853,I124934,);
nor I_6902 (I124943,I124934,I124880);
not I_6903 (I124961,I124934);
DFFARX1 I_6904 (I124583,I691,I124853,I124988,);
nand I_6905 (I124997,I124988,I124430);
not I_6906 (I125015,I124997);
DFFARX1 I_6907 (I125015,I691,I124853,I125042,);
not I_6908 (I125051,I125042);
nor I_6909 (I125069,I124880,I124997);
nor I_6910 (I125087,I124934,I125069);
DFFARX1 I_6911 (I124817,I691,I124853,I125114,);
DFFARX1 I_6912 (I125114,I691,I124853,I125132,);
not I_6913 (I125141,I125132);
not I_6914 (I125159,I125114);
nand I_6915 (I125177,I125159,I124961);
nand I_6916 (I125195,I124790,I124835);
and I_6917 (I125213,I125195,I124511);
DFFARX1 I_6918 (I125213,I691,I124853,I125240,);
nor I_6919 (I125249,I125240,I124880);
DFFARX1 I_6920 (I125249,I691,I124853,I125276,);
DFFARX1 I_6921 (I125240,I691,I124853,I125294,);
nor I_6922 (I125303,I124565,I124835);
not I_6923 (I125321,I125303);
nor I_6924 (I125339,I125141,I125321);
nand I_6925 (I125357,I125159,I125321);
nor I_6926 (I125375,I124880,I125303);
DFFARX1 I_6927 (I125303,I691,I124853,I125402,);
not I_6928 (I125411,I698);
DFFARX1 I_6929 (I125276,I691,I125411,I125438,);
DFFARX1 I_6930 (I125357,I691,I125411,I125456,);
not I_6931 (I125465,I125456);
not I_6932 (I125483,I125051);
nor I_6933 (I125501,I125483,I125375);
not I_6934 (I125519,I125402);
nor I_6935 (I125537,I125501,I125087);
nor I_6936 (I125555,I125456,I125537);
DFFARX1 I_6937 (I125555,I691,I125411,I125582,);
nor I_6938 (I125591,I125087,I125375);
nand I_6939 (I125609,I125591,I125051);
DFFARX1 I_6940 (I125609,I691,I125411,I125636,);
nor I_6941 (I125645,I125519,I125087);
nand I_6942 (I125663,I125645,I125276);
nor I_6943 (I125681,I125438,I125663);
DFFARX1 I_6944 (I125681,I691,I125411,I125708,);
not I_6945 (I125717,I125663);
nand I_6946 (I125735,I125456,I125717);
DFFARX1 I_6947 (I125663,I691,I125411,I125762,);
not I_6948 (I125771,I125762);
not I_6949 (I125789,I125087);
not I_6950 (I125807,I125177);
nor I_6951 (I125825,I125807,I125402);
nor I_6952 (I125843,I125771,I125825);
nor I_6953 (I125861,I125807,I125339);
and I_6954 (I125879,I125861,I124943);
or I_6955 (I125897,I125879,I125294);
DFFARX1 I_6956 (I125897,I691,I125411,I125924,);
nor I_6957 (I125933,I125924,I125438);
not I_6958 (I125951,I125924);
and I_6959 (I125969,I125951,I125438);
nor I_6960 (I125987,I125465,I125969);
nand I_6961 (I126005,I125951,I125519);
nor I_6962 (I126023,I125807,I126005);
nand I_6963 (I126041,I125951,I125717);
nand I_6964 (I126059,I125519,I125177);
nor I_6965 (I126077,I125789,I126059);
not I_6966 (I126095,I698);
DFFARX1 I_6967 (I125636,I691,I126095,I126122,);
not I_6968 (I126131,I126122);
nand I_6969 (I126149,I125708,I125933);
and I_6970 (I126167,I126149,I125843);
DFFARX1 I_6971 (I126167,I691,I126095,I126194,);
not I_6972 (I126203,I125735);
DFFARX1 I_6973 (I126023,I691,I126095,I126230,);
not I_6974 (I126239,I126230);
nor I_6975 (I126257,I126239,I126131);
and I_6976 (I126275,I126257,I125735);
nor I_6977 (I126293,I126239,I126203);
nor I_6978 (I126311,I126194,I126293);
DFFARX1 I_6979 (I125708,I691,I126095,I126338,);
nor I_6980 (I126347,I126338,I126194);
not I_6981 (I126365,I126347);
not I_6982 (I126383,I126338);
nor I_6983 (I126401,I126383,I126275);
DFFARX1 I_6984 (I126401,I691,I126095,I126428,);
nand I_6985 (I126437,I126077,I125987);
and I_6986 (I126455,I126437,I125582);
DFFARX1 I_6987 (I126455,I691,I126095,I126482,);
nor I_6988 (I126491,I126482,I126338);
DFFARX1 I_6989 (I126491,I691,I126095,I126518,);
nand I_6990 (I126527,I126482,I126383);
nand I_6991 (I126545,I126365,I126527);
not I_6992 (I126563,I126482);
nor I_6993 (I126581,I126563,I126275);
DFFARX1 I_6994 (I126581,I691,I126095,I126608,);
nor I_6995 (I126617,I126041,I125987);
or I_6996 (I126635,I126338,I126617);
nor I_6997 (I126653,I126482,I126617);
or I_6998 (I126671,I126194,I126617);
DFFARX1 I_6999 (I126617,I691,I126095,I126698,);
not I_7000 (I126707,I698);
DFFARX1 I_7001 (I126311,I691,I126707,I126734,);
and I_7002 (I126743,I126734,I126653);
DFFARX1 I_7003 (I126743,I691,I126707,I126770,);
DFFARX1 I_7004 (I126671,I691,I126707,I126788,);
not I_7005 (I126797,I126518);
not I_7006 (I126815,I126698);
nand I_7007 (I126833,I126815,I126797);
nor I_7008 (I126851,I126788,I126833);
DFFARX1 I_7009 (I126833,I691,I126707,I126878,);
not I_7010 (I126887,I126878);
not I_7011 (I126905,I126635);
nand I_7012 (I126923,I126815,I126905);
DFFARX1 I_7013 (I126923,I691,I126707,I126950,);
not I_7014 (I126959,I126950);
not I_7015 (I126977,I126608);
nand I_7016 (I126995,I126977,I126428);
and I_7017 (I127013,I126797,I126995);
nor I_7018 (I127031,I126923,I127013);
DFFARX1 I_7019 (I127031,I691,I126707,I127058,);
DFFARX1 I_7020 (I127013,I691,I126707,I127076,);
nor I_7021 (I127085,I126608,I126545);
nor I_7022 (I127103,I126923,I127085);
or I_7023 (I127121,I126608,I126545);
nor I_7024 (I127139,I126518,I126653);
DFFARX1 I_7025 (I127139,I691,I126707,I127166,);
not I_7026 (I127175,I127166);
nor I_7027 (I127193,I127175,I126959);
nand I_7028 (I127211,I127175,I126788);
not I_7029 (I127229,I126518);
nand I_7030 (I127247,I127229,I126905);
nand I_7031 (I127265,I127175,I127247);
nand I_7032 (I127283,I127265,I127211);
nand I_7033 (I127301,I127247,I127121);
not I_7034 (I127319,I698);
DFFARX1 I_7035 (I127058,I691,I127319,I127346,);
nand I_7036 (I127355,I126770,I127058);
and I_7037 (I127373,I127355,I127193);
DFFARX1 I_7038 (I127373,I691,I127319,I127400,);
nor I_7039 (I127409,I127400,I127346);
not I_7040 (I127427,I127400);
DFFARX1 I_7041 (I126887,I691,I127319,I127454,);
nand I_7042 (I127463,I127454,I127301);
not I_7043 (I127481,I127463);
DFFARX1 I_7044 (I127481,I691,I127319,I127508,);
not I_7045 (I127517,I127508);
nor I_7046 (I127535,I127346,I127463);
nor I_7047 (I127553,I127400,I127535);
DFFARX1 I_7048 (I126851,I691,I127319,I127580,);
DFFARX1 I_7049 (I127580,I691,I127319,I127598,);
not I_7050 (I127607,I127598);
not I_7051 (I127625,I127580);
nand I_7052 (I127643,I127625,I127427);
nand I_7053 (I127661,I126851,I127283);
and I_7054 (I127679,I127661,I127076);
DFFARX1 I_7055 (I127679,I691,I127319,I127706,);
nor I_7056 (I127715,I127706,I127346);
DFFARX1 I_7057 (I127715,I691,I127319,I127742,);
DFFARX1 I_7058 (I127706,I691,I127319,I127760,);
nor I_7059 (I127769,I127103,I127283);
not I_7060 (I127787,I127769);
nor I_7061 (I127805,I127607,I127787);
nand I_7062 (I127823,I127625,I127787);
nor I_7063 (I127841,I127346,I127769);
DFFARX1 I_7064 (I127769,I691,I127319,I127868,);
not I_7065 (I127877,I698);
DFFARX1 I_7066 (I127805,I691,I127877,I127904,);
DFFARX1 I_7067 (I127904,I691,I127877,I127922,);
not I_7068 (I127931,I127922);
not I_7069 (I127949,I127904);
nand I_7070 (I127967,I127742,I127868);
and I_7071 (I127985,I127967,I127517);
DFFARX1 I_7072 (I127985,I691,I127877,I128012,);
not I_7073 (I128021,I128012);
DFFARX1 I_7074 (I127553,I691,I127877,I128048,);
and I_7075 (I128057,I128048,I127841);
nand I_7076 (I128075,I128048,I127841);
nand I_7077 (I128093,I128021,I128075);
DFFARX1 I_7078 (I127409,I691,I127877,I128120,);
nor I_7079 (I128129,I128120,I128057);
DFFARX1 I_7080 (I128129,I691,I127877,I128156,);
nor I_7081 (I128165,I128120,I128012);
nand I_7082 (I128183,I127643,I127742);
and I_7083 (I128201,I128183,I127823);
DFFARX1 I_7084 (I128201,I691,I127877,I128228,);
nor I_7085 (I128237,I128228,I128120);
not I_7086 (I128255,I128228);
nor I_7087 (I128273,I128255,I128021);
nor I_7088 (I128291,I127949,I128273);
DFFARX1 I_7089 (I128291,I691,I127877,I128318,);
nor I_7090 (I128327,I128255,I128120);
nor I_7091 (I128345,I127760,I127742);
nor I_7092 (I128363,I128345,I128327);
not I_7093 (I128381,I128345);
nand I_7094 (I128399,I128075,I128381);
DFFARX1 I_7095 (I128345,I691,I127877,I128426,);
DFFARX1 I_7096 (I128345,I691,I127877,I128444,);
not I_7097 (I128453,I698);
DFFARX1 I_7098 (I128093,I691,I128453,I128480,);
DFFARX1 I_7099 (I128237,I691,I128453,I128498,);
not I_7100 (I128507,I128498);
not I_7101 (I128525,I128318);
nor I_7102 (I128543,I128525,I128444);
not I_7103 (I128561,I128363);
nor I_7104 (I128579,I128543,I128165);
nor I_7105 (I128597,I128498,I128579);
DFFARX1 I_7106 (I128597,I691,I128453,I128624,);
nor I_7107 (I128633,I128165,I128444);
nand I_7108 (I128651,I128633,I128318);
DFFARX1 I_7109 (I128651,I691,I128453,I128678,);
nor I_7110 (I128687,I128561,I128165);
nand I_7111 (I128705,I128687,I127931);
nor I_7112 (I128723,I128480,I128705);
DFFARX1 I_7113 (I128723,I691,I128453,I128750,);
not I_7114 (I128759,I128705);
nand I_7115 (I128777,I128498,I128759);
DFFARX1 I_7116 (I128705,I691,I128453,I128804,);
not I_7117 (I128813,I128804);
not I_7118 (I128831,I128165);
not I_7119 (I128849,I128156);
nor I_7120 (I128867,I128849,I128363);
nor I_7121 (I128885,I128813,I128867);
nor I_7122 (I128903,I128849,I128399);
and I_7123 (I128921,I128903,I128156);
or I_7124 (I128939,I128921,I128426);
DFFARX1 I_7125 (I128939,I691,I128453,I128966,);
nor I_7126 (I128975,I128966,I128480);
not I_7127 (I128993,I128966);
and I_7128 (I129011,I128993,I128480);
nor I_7129 (I129029,I128507,I129011);
nand I_7130 (I129047,I128993,I128561);
nor I_7131 (I129065,I128849,I129047);
nand I_7132 (I129083,I128993,I128759);
nand I_7133 (I129101,I128561,I128156);
nor I_7134 (I129119,I128831,I129101);
not I_7135 (I129137,I698);
DFFARX1 I_7136 (I129065,I691,I129137,I129164,);
not I_7137 (I129173,I129164);
nand I_7138 (I129191,I129119,I128750);
and I_7139 (I129209,I129191,I128750);
DFFARX1 I_7140 (I129209,I691,I129137,I129236,);
DFFARX1 I_7141 (I129236,I691,I129137,I129254,);
DFFARX1 I_7142 (I129029,I691,I129137,I129272,);
nand I_7143 (I129281,I129272,I128885);
not I_7144 (I129299,I129281);
DFFARX1 I_7145 (I129299,I691,I129137,I129326,);
not I_7146 (I129335,I129326);
nor I_7147 (I129353,I129173,I129335);
DFFARX1 I_7148 (I128678,I691,I129137,I129380,);
nor I_7149 (I129389,I129380,I129236);
nor I_7150 (I129407,I129380,I129299);
nand I_7151 (I129425,I128624,I128777);
and I_7152 (I129443,I129425,I129083);
DFFARX1 I_7153 (I129443,I691,I129137,I129470,);
not I_7154 (I129479,I129470);
nand I_7155 (I129497,I129479,I129380);
nand I_7156 (I129515,I129479,I129281);
nor I_7157 (I129533,I128975,I128777);
and I_7158 (I129551,I129380,I129533);
nor I_7159 (I129569,I129479,I129551);
DFFARX1 I_7160 (I129569,I691,I129137,I129596,);
nor I_7161 (I129605,I129164,I129533);
DFFARX1 I_7162 (I129605,I691,I129137,I129632,);
nor I_7163 (I129641,I129470,I129533);
not I_7164 (I129659,I129641);
nand I_7165 (I129677,I129659,I129497);
not I_7166 (I129695,I698);
DFFARX1 I_7167 (I129677,I691,I129695,I129722,);
DFFARX1 I_7168 (I129722,I691,I129695,I129740,);
not I_7169 (I129749,I129740);
nand I_7170 (I129767,I129632,I129353);
and I_7171 (I129785,I129767,I129407);
DFFARX1 I_7172 (I129785,I691,I129695,I129812,);
DFFARX1 I_7173 (I129812,I691,I129695,I129830,);
DFFARX1 I_7174 (I129812,I691,I129695,I129848,);
DFFARX1 I_7175 (I129407,I691,I129695,I129866,);
nand I_7176 (I129875,I129866,I129254);
not I_7177 (I129893,I129875);
nor I_7178 (I129911,I129722,I129893);
DFFARX1 I_7179 (I129389,I691,I129695,I129938,);
not I_7180 (I129947,I129938);
nor I_7181 (I129965,I129947,I129749);
nand I_7182 (I129983,I129947,I129875);
nand I_7183 (I130001,I129515,I129596);
and I_7184 (I130019,I130001,I129632);
DFFARX1 I_7185 (I130019,I691,I129695,I130046,);
nor I_7186 (I130055,I130046,I129722);
DFFARX1 I_7187 (I130055,I691,I129695,I130082,);
not I_7188 (I130091,I130046);
nor I_7189 (I130109,I129515,I129596);
not I_7190 (I130127,I130109);
nor I_7191 (I130145,I129875,I130127);
nor I_7192 (I130163,I130091,I130145);
DFFARX1 I_7193 (I130163,I691,I129695,I130190,);
nor I_7194 (I130199,I130046,I130127);
nor I_7195 (I130217,I129893,I130199);
nor I_7196 (I130235,I130046,I130109);
not I_7197 (I130253,I698);
DFFARX1 I_7198 (I129911,I691,I130253,I130280,);
not I_7199 (I130289,I130280);
nand I_7200 (I130307,I130217,I130082);
and I_7201 (I130325,I130307,I130082);
DFFARX1 I_7202 (I130325,I691,I130253,I130352,);
not I_7203 (I130361,I130235);
DFFARX1 I_7204 (I129965,I691,I130253,I130388,);
not I_7205 (I130397,I130388);
nor I_7206 (I130415,I130397,I130289);
and I_7207 (I130433,I130415,I130235);
nor I_7208 (I130451,I130397,I130361);
nor I_7209 (I130469,I130352,I130451);
DFFARX1 I_7210 (I130235,I691,I130253,I130496,);
nor I_7211 (I130505,I130496,I130352);
not I_7212 (I130523,I130505);
not I_7213 (I130541,I130496);
nor I_7214 (I130559,I130541,I130433);
DFFARX1 I_7215 (I130559,I691,I130253,I130586,);
nand I_7216 (I130595,I130190,I129983);
and I_7217 (I130613,I130595,I129848);
DFFARX1 I_7218 (I130613,I691,I130253,I130640,);
nor I_7219 (I130649,I130640,I130496);
DFFARX1 I_7220 (I130649,I691,I130253,I130676,);
nand I_7221 (I130685,I130640,I130541);
nand I_7222 (I130703,I130523,I130685);
not I_7223 (I130721,I130640);
nor I_7224 (I130739,I130721,I130433);
DFFARX1 I_7225 (I130739,I691,I130253,I130766,);
nor I_7226 (I130775,I129830,I129983);
or I_7227 (I130793,I130496,I130775);
nor I_7228 (I130811,I130640,I130775);
or I_7229 (I130829,I130352,I130775);
DFFARX1 I_7230 (I130775,I691,I130253,I130856,);
not I_7231 (I130865,I698);
DFFARX1 I_7232 (I130676,I691,I130865,I130892,);
nand I_7233 (I130901,I130892,I130811);
not I_7234 (I130919,I130901);
DFFARX1 I_7235 (I130469,I691,I130865,I130946,);
not I_7236 (I130955,I130946);
not I_7237 (I130973,I130676);
or I_7238 (I130991,I130703,I130676);
nor I_7239 (I131009,I130703,I130676);
or I_7240 (I131027,I130586,I130703);
DFFARX1 I_7241 (I131027,I691,I130865,I131054,);
not I_7242 (I131063,I130766);
nand I_7243 (I131081,I131063,I130811);
nand I_7244 (I131099,I130973,I131081);
and I_7245 (I131117,I130955,I131099);
nor I_7246 (I131135,I130766,I130829);
and I_7247 (I131153,I130955,I131135);
nor I_7248 (I131171,I130919,I131153);
DFFARX1 I_7249 (I131135,I691,I130865,I131198,);
not I_7250 (I131207,I131198);
nor I_7251 (I131225,I130955,I131207);
or I_7252 (I131243,I131027,I130793);
nor I_7253 (I131261,I130793,I130586);
nand I_7254 (I131279,I131099,I131261);
nand I_7255 (I131297,I131243,I131279);
DFFARX1 I_7256 (I131297,I691,I130865,I131324,);
nor I_7257 (I131333,I131261,I130991);
DFFARX1 I_7258 (I131333,I691,I130865,I131360,);
nor I_7259 (I131369,I130793,I130856);
DFFARX1 I_7260 (I131369,I691,I130865,I131396,);
DFFARX1 I_7261 (I131396,I691,I130865,I131414,);
not I_7262 (I131423,I131396);
nand I_7263 (I131441,I131423,I130901);
nand I_7264 (I131459,I131423,I131009);
not I_7265 (I131477,I698);
DFFARX1 I_7266 (I131054,I691,I131477,I131504,);
and I_7267 (I131513,I131504,I131459);
DFFARX1 I_7268 (I131513,I691,I131477,I131540,);
DFFARX1 I_7269 (I131414,I691,I131477,I131558,);
not I_7270 (I131567,I131360);
not I_7271 (I131585,I131441);
nand I_7272 (I131603,I131585,I131567);
nor I_7273 (I131621,I131558,I131603);
DFFARX1 I_7274 (I131603,I691,I131477,I131648,);
not I_7275 (I131657,I131648);
not I_7276 (I131675,I131117);
nand I_7277 (I131693,I131585,I131675);
DFFARX1 I_7278 (I131693,I691,I131477,I131720,);
not I_7279 (I131729,I131720);
not I_7280 (I131747,I131360);
nand I_7281 (I131765,I131747,I131117);
and I_7282 (I131783,I131567,I131765);
nor I_7283 (I131801,I131693,I131783);
DFFARX1 I_7284 (I131801,I691,I131477,I131828,);
DFFARX1 I_7285 (I131783,I691,I131477,I131846,);
nor I_7286 (I131855,I131360,I131324);
nor I_7287 (I131873,I131693,I131855);
or I_7288 (I131891,I131360,I131324);
nor I_7289 (I131909,I131171,I131225);
DFFARX1 I_7290 (I131909,I691,I131477,I131936,);
not I_7291 (I131945,I131936);
nor I_7292 (I131963,I131945,I131729);
nand I_7293 (I131981,I131945,I131558);
not I_7294 (I131999,I131171);
nand I_7295 (I132017,I131999,I131675);
nand I_7296 (I132035,I131945,I132017);
nand I_7297 (I132053,I132035,I131981);
nand I_7298 (I132071,I132017,I131891);
not I_7299 (I132089,I698);
DFFARX1 I_7300 (I131828,I691,I132089,I132116,);
nand I_7301 (I132125,I131540,I131828);
and I_7302 (I132143,I132125,I131963);
DFFARX1 I_7303 (I132143,I691,I132089,I132170,);
nor I_7304 (I132179,I132170,I132116);
not I_7305 (I132197,I132170);
DFFARX1 I_7306 (I131657,I691,I132089,I132224,);
nand I_7307 (I132233,I132224,I132071);
not I_7308 (I132251,I132233);
DFFARX1 I_7309 (I132251,I691,I132089,I132278,);
not I_7310 (I132287,I132278);
nor I_7311 (I132305,I132116,I132233);
nor I_7312 (I132323,I132170,I132305);
DFFARX1 I_7313 (I131621,I691,I132089,I132350,);
DFFARX1 I_7314 (I132350,I691,I132089,I132368,);
not I_7315 (I132377,I132368);
not I_7316 (I132395,I132350);
nand I_7317 (I132413,I132395,I132197);
nand I_7318 (I132431,I131621,I132053);
and I_7319 (I132449,I132431,I131846);
DFFARX1 I_7320 (I132449,I691,I132089,I132476,);
nor I_7321 (I132485,I132476,I132116);
DFFARX1 I_7322 (I132485,I691,I132089,I132512,);
DFFARX1 I_7323 (I132476,I691,I132089,I132530,);
nor I_7324 (I132539,I131873,I132053);
not I_7325 (I132557,I132539);
nor I_7326 (I132575,I132377,I132557);
nand I_7327 (I132593,I132395,I132557);
nor I_7328 (I132611,I132116,I132539);
DFFARX1 I_7329 (I132539,I691,I132089,I132638,);
not I_7330 (I132647,I698);
DFFARX1 I_7331 (I132638,I691,I132647,I132674,);
not I_7332 (I132683,I132674);
nand I_7333 (I132701,I132287,I132179);
and I_7334 (I132719,I132701,I132512);
DFFARX1 I_7335 (I132719,I691,I132647,I132746,);
not I_7336 (I132755,I132593);
DFFARX1 I_7337 (I132512,I691,I132647,I132782,);
not I_7338 (I132791,I132782);
nor I_7339 (I132809,I132791,I132683);
and I_7340 (I132827,I132809,I132593);
nor I_7341 (I132845,I132791,I132755);
nor I_7342 (I132863,I132746,I132845);
DFFARX1 I_7343 (I132323,I691,I132647,I132890,);
nor I_7344 (I132899,I132890,I132746);
not I_7345 (I132917,I132899);
not I_7346 (I132935,I132890);
nor I_7347 (I132953,I132935,I132827);
DFFARX1 I_7348 (I132953,I691,I132647,I132980,);
nand I_7349 (I132989,I132413,I132575);
and I_7350 (I133007,I132989,I132530);
DFFARX1 I_7351 (I133007,I691,I132647,I133034,);
nor I_7352 (I133043,I133034,I132890);
DFFARX1 I_7353 (I133043,I691,I132647,I133070,);
nand I_7354 (I133079,I133034,I132935);
nand I_7355 (I133097,I132917,I133079);
not I_7356 (I133115,I133034);
nor I_7357 (I133133,I133115,I132827);
DFFARX1 I_7358 (I133133,I691,I132647,I133160,);
nor I_7359 (I133169,I132611,I132575);
or I_7360 (I133187,I132890,I133169);
nor I_7361 (I133205,I133034,I133169);
or I_7362 (I133223,I132746,I133169);
DFFARX1 I_7363 (I133169,I691,I132647,I133250,);
not I_7364 (I133259,I698);
DFFARX1 I_7365 (I133070,I691,I133259,I133286,);
not I_7366 (I133295,I133286);
DFFARX1 I_7367 (I133187,I691,I133259,I133322,);
not I_7368 (I133331,I133205);
nand I_7369 (I133349,I133331,I133223);
not I_7370 (I133367,I133349);
nor I_7371 (I133385,I133367,I133097);
nor I_7372 (I133403,I133295,I133385);
DFFARX1 I_7373 (I133403,I691,I133259,I133430,);
not I_7374 (I133439,I133097);
nand I_7375 (I133457,I133439,I133367);
and I_7376 (I133475,I133439,I133205);
nand I_7377 (I133493,I133475,I132863);
nor I_7378 (I133511,I133493,I133439);
and I_7379 (I133529,I133322,I133493);
not I_7380 (I133547,I133493);
nand I_7381 (I133565,I133322,I133547);
nor I_7382 (I133583,I133286,I133493);
not I_7383 (I133601,I133160);
nor I_7384 (I133619,I133601,I133205);
nand I_7385 (I133637,I133619,I133439);
nor I_7386 (I133655,I133349,I133637);
nor I_7387 (I133673,I133601,I133070);
and I_7388 (I133691,I133673,I132980);
or I_7389 (I133709,I133691,I133250);
DFFARX1 I_7390 (I133709,I691,I133259,I133736,);
nor I_7391 (I133745,I133736,I133457);
DFFARX1 I_7392 (I133745,I691,I133259,I133772,);
DFFARX1 I_7393 (I133736,I691,I133259,I133790,);
not I_7394 (I133799,I133736);
nor I_7395 (I133817,I133799,I133322);
nor I_7396 (I133835,I133619,I133817);
DFFARX1 I_7397 (I133835,I691,I133259,I133862,);
not I_7398 (I133871,I698);
DFFARX1 I_7399 (I133565,I691,I133871,I133898,);
not I_7400 (I133907,I133898);
nand I_7401 (I133925,I133862,I133529);
and I_7402 (I133943,I133925,I133772);
DFFARX1 I_7403 (I133943,I691,I133871,I133970,);
DFFARX1 I_7404 (I133511,I691,I133871,I133988,);
and I_7405 (I133997,I133988,I133583);
nor I_7406 (I134015,I133970,I133997);
DFFARX1 I_7407 (I134015,I691,I133871,I134042,);
nand I_7408 (I134051,I133988,I133583);
nand I_7409 (I134069,I133907,I134051);
not I_7410 (I134087,I134069);
DFFARX1 I_7411 (I133655,I691,I133871,I134114,);
DFFARX1 I_7412 (I134114,I691,I133871,I134132,);
nand I_7413 (I134141,I133430,I133790);
and I_7414 (I134159,I134141,I133772);
DFFARX1 I_7415 (I134159,I691,I133871,I134186,);
DFFARX1 I_7416 (I134186,I691,I133871,I134204,);
not I_7417 (I134213,I134204);
not I_7418 (I134231,I134186);
nand I_7419 (I134249,I134231,I134051);
nor I_7420 (I134267,I133583,I133790);
not I_7421 (I134285,I134267);
nor I_7422 (I134303,I134231,I134285);
nor I_7423 (I134321,I133907,I134303);
DFFARX1 I_7424 (I134321,I691,I133871,I134348,);
nor I_7425 (I134357,I133970,I134285);
nor I_7426 (I134375,I134186,I134357);
nor I_7427 (I134393,I134114,I134267);
nor I_7428 (I134411,I133970,I134267);
not I_7429 (I134429,I698);
DFFARX1 I_7430 (I134375,I691,I134429,I134456,);
DFFARX1 I_7431 (I134456,I691,I134429,I134474,);
not I_7432 (I134483,I134474);
not I_7433 (I134501,I134456);
nand I_7434 (I134519,I134132,I134042);
and I_7435 (I134537,I134519,I134411);
DFFARX1 I_7436 (I134537,I691,I134429,I134564,);
not I_7437 (I134573,I134564);
DFFARX1 I_7438 (I134249,I691,I134429,I134600,);
and I_7439 (I134609,I134600,I134411);
nand I_7440 (I134627,I134600,I134411);
nand I_7441 (I134645,I134573,I134627);
DFFARX1 I_7442 (I134348,I691,I134429,I134672,);
nor I_7443 (I134681,I134672,I134609);
DFFARX1 I_7444 (I134681,I691,I134429,I134708,);
nor I_7445 (I134717,I134672,I134564);
nand I_7446 (I134735,I134042,I134393);
and I_7447 (I134753,I134735,I134087);
DFFARX1 I_7448 (I134753,I691,I134429,I134780,);
nor I_7449 (I134789,I134780,I134672);
not I_7450 (I134807,I134780);
nor I_7451 (I134825,I134807,I134573);
nor I_7452 (I134843,I134501,I134825);
DFFARX1 I_7453 (I134843,I691,I134429,I134870,);
nor I_7454 (I134879,I134807,I134672);
nor I_7455 (I134897,I134213,I134393);
nor I_7456 (I134915,I134897,I134879);
not I_7457 (I134933,I134897);
nand I_7458 (I134951,I134627,I134933);
DFFARX1 I_7459 (I134897,I691,I134429,I134978,);
DFFARX1 I_7460 (I134897,I691,I134429,I134996,);
not I_7461 (I135005,I698);
DFFARX1 I_7462 (I134789,I691,I135005,I135032,);
nand I_7463 (I135041,I135032,I134951);
not I_7464 (I135059,I135041);
DFFARX1 I_7465 (I134708,I691,I135005,I135086,);
not I_7466 (I135095,I135086);
not I_7467 (I135113,I134645);
or I_7468 (I135131,I134708,I134645);
nor I_7469 (I135149,I134708,I134645);
or I_7470 (I135167,I134717,I134708);
DFFARX1 I_7471 (I135167,I691,I135005,I135194,);
not I_7472 (I135203,I134915);
nand I_7473 (I135221,I135203,I134996);
nand I_7474 (I135239,I135113,I135221);
and I_7475 (I135257,I135095,I135239);
nor I_7476 (I135275,I134915,I134483);
and I_7477 (I135293,I135095,I135275);
nor I_7478 (I135311,I135059,I135293);
DFFARX1 I_7479 (I135275,I691,I135005,I135338,);
not I_7480 (I135347,I135338);
nor I_7481 (I135365,I135095,I135347);
or I_7482 (I135383,I135167,I134870);
nor I_7483 (I135401,I134870,I134717);
nand I_7484 (I135419,I135239,I135401);
nand I_7485 (I135437,I135383,I135419);
DFFARX1 I_7486 (I135437,I691,I135005,I135464,);
nor I_7487 (I135473,I135401,I135131);
DFFARX1 I_7488 (I135473,I691,I135005,I135500,);
nor I_7489 (I135509,I134870,I134978);
DFFARX1 I_7490 (I135509,I691,I135005,I135536,);
DFFARX1 I_7491 (I135536,I691,I135005,I135554,);
not I_7492 (I135563,I135536);
nand I_7493 (I135581,I135563,I135041);
nand I_7494 (I135599,I135563,I135149);
not I_7495 (I135617,I698);
DFFARX1 I_7496 (I135194,I691,I135617,I135644,);
and I_7497 (I135653,I135644,I135599);
DFFARX1 I_7498 (I135653,I691,I135617,I135680,);
DFFARX1 I_7499 (I135554,I691,I135617,I135698,);
not I_7500 (I135707,I135500);
not I_7501 (I135725,I135581);
nand I_7502 (I135743,I135725,I135707);
nor I_7503 (I135761,I135698,I135743);
DFFARX1 I_7504 (I135743,I691,I135617,I135788,);
not I_7505 (I135797,I135788);
not I_7506 (I135815,I135257);
nand I_7507 (I135833,I135725,I135815);
DFFARX1 I_7508 (I135833,I691,I135617,I135860,);
not I_7509 (I135869,I135860);
not I_7510 (I135887,I135500);
nand I_7511 (I135905,I135887,I135257);
and I_7512 (I135923,I135707,I135905);
nor I_7513 (I135941,I135833,I135923);
DFFARX1 I_7514 (I135941,I691,I135617,I135968,);
DFFARX1 I_7515 (I135923,I691,I135617,I135986,);
nor I_7516 (I135995,I135500,I135464);
nor I_7517 (I136013,I135833,I135995);
or I_7518 (I136031,I135500,I135464);
nor I_7519 (I136049,I135311,I135365);
DFFARX1 I_7520 (I136049,I691,I135617,I136076,);
not I_7521 (I136085,I136076);
nor I_7522 (I136103,I136085,I135869);
nand I_7523 (I136121,I136085,I135698);
not I_7524 (I136139,I135311);
nand I_7525 (I136157,I136139,I135815);
nand I_7526 (I136175,I136085,I136157);
nand I_7527 (I136193,I136175,I136121);
nand I_7528 (I136211,I136157,I136031);
not I_7529 (I136229,I698);
DFFARX1 I_7530 (I136103,I691,I136229,I136256,);
not I_7531 (I136265,I136256);
nand I_7532 (I136283,I135968,I135968);
and I_7533 (I136301,I136283,I136211);
DFFARX1 I_7534 (I136301,I691,I136229,I136328,);
DFFARX1 I_7535 (I136328,I691,I136229,I136346,);
DFFARX1 I_7536 (I135761,I691,I136229,I136364,);
nand I_7537 (I136373,I136364,I136013);
not I_7538 (I136391,I136373);
DFFARX1 I_7539 (I136391,I691,I136229,I136418,);
not I_7540 (I136427,I136418);
nor I_7541 (I136445,I136265,I136427);
DFFARX1 I_7542 (I135797,I691,I136229,I136472,);
nor I_7543 (I136481,I136472,I136328);
nor I_7544 (I136499,I136472,I136391);
nand I_7545 (I136517,I135680,I136193);
and I_7546 (I136535,I136517,I135761);
DFFARX1 I_7547 (I136535,I691,I136229,I136562,);
not I_7548 (I136571,I136562);
nand I_7549 (I136589,I136571,I136472);
nand I_7550 (I136607,I136571,I136373);
nor I_7551 (I136625,I135986,I136193);
and I_7552 (I136643,I136472,I136625);
nor I_7553 (I136661,I136571,I136643);
DFFARX1 I_7554 (I136661,I691,I136229,I136688,);
nor I_7555 (I136697,I136256,I136625);
DFFARX1 I_7556 (I136697,I691,I136229,I136724,);
nor I_7557 (I136733,I136562,I136625);
not I_7558 (I136751,I136733);
nand I_7559 (I136769,I136751,I136589);
not I_7560 (I136787,I698);
DFFARX1 I_7561 (I136499,I691,I136787,I136814,);
nand I_7562 (I136823,I136814,I136499);
not I_7563 (I136841,I136823);
DFFARX1 I_7564 (I136769,I691,I136787,I136868,);
not I_7565 (I136877,I136868);
not I_7566 (I136895,I136445);
or I_7567 (I136913,I136607,I136445);
nor I_7568 (I136931,I136607,I136445);
or I_7569 (I136949,I136724,I136607);
DFFARX1 I_7570 (I136949,I691,I136787,I136976,);
not I_7571 (I136985,I136346);
nand I_7572 (I137003,I136985,I136481);
nand I_7573 (I137021,I136895,I137003);
and I_7574 (I137039,I136877,I137021);
nor I_7575 (I137057,I136346,I136724);
and I_7576 (I137075,I136877,I137057);
nor I_7577 (I137093,I136841,I137075);
DFFARX1 I_7578 (I137057,I691,I136787,I137120,);
not I_7579 (I137129,I137120);
nor I_7580 (I137147,I136877,I137129);
or I_7581 (I137165,I136949,I136688);
nor I_7582 (I137183,I136688,I136724);
nand I_7583 (I137201,I137021,I137183);
nand I_7584 (I137219,I137165,I137201);
DFFARX1 I_7585 (I137219,I691,I136787,I137246,);
nor I_7586 (I137255,I137183,I136913);
DFFARX1 I_7587 (I137255,I691,I136787,I137282,);
nor I_7588 (I137291,I136688,I136607);
DFFARX1 I_7589 (I137291,I691,I136787,I137318,);
DFFARX1 I_7590 (I137318,I691,I136787,I137336,);
not I_7591 (I137345,I137318);
nand I_7592 (I137363,I137345,I136823);
nand I_7593 (I137381,I137345,I136931);
not I_7594 (I137399,I698);
DFFARX1 I_7595 (I137282,I691,I137399,I137426,);
not I_7596 (I137435,I137426);
nand I_7597 (I137453,I136976,I137381);
and I_7598 (I137471,I137453,I137363);
DFFARX1 I_7599 (I137471,I691,I137399,I137498,);
not I_7600 (I137507,I137147);
DFFARX1 I_7601 (I137039,I691,I137399,I137534,);
not I_7602 (I137543,I137534);
nor I_7603 (I137561,I137543,I137435);
and I_7604 (I137579,I137561,I137147);
nor I_7605 (I137597,I137543,I137507);
nor I_7606 (I137615,I137498,I137597);
DFFARX1 I_7607 (I137336,I691,I137399,I137642,);
nor I_7608 (I137651,I137642,I137498);
not I_7609 (I137669,I137651);
not I_7610 (I137687,I137642);
nor I_7611 (I137705,I137687,I137579);
DFFARX1 I_7612 (I137705,I691,I137399,I137732,);
nand I_7613 (I137741,I137246,I137093);
and I_7614 (I137759,I137741,I137039);
DFFARX1 I_7615 (I137759,I691,I137399,I137786,);
nor I_7616 (I137795,I137786,I137642);
DFFARX1 I_7617 (I137795,I691,I137399,I137822,);
nand I_7618 (I137831,I137786,I137687);
nand I_7619 (I137849,I137669,I137831);
not I_7620 (I137867,I137786);
nor I_7621 (I137885,I137867,I137579);
DFFARX1 I_7622 (I137885,I691,I137399,I137912,);
nor I_7623 (I137921,I137282,I137093);
or I_7624 (I137939,I137642,I137921);
nor I_7625 (I137957,I137786,I137921);
or I_7626 (I137975,I137498,I137921);
DFFARX1 I_7627 (I137921,I691,I137399,I138002,);
not I_7628 (I138011,I698);
DFFARX1 I_7629 (I137822,I691,I138011,I138038,);
not I_7630 (I138047,I138038);
DFFARX1 I_7631 (I137939,I691,I138011,I138074,);
not I_7632 (I138083,I137957);
nand I_7633 (I138101,I138083,I137975);
not I_7634 (I138119,I138101);
nor I_7635 (I138137,I138119,I137849);
nor I_7636 (I138155,I138047,I138137);
DFFARX1 I_7637 (I138155,I691,I138011,I138182,);
not I_7638 (I138191,I137849);
nand I_7639 (I138209,I138191,I138119);
and I_7640 (I138227,I138191,I137957);
nand I_7641 (I138245,I138227,I137615);
nor I_7642 (I138263,I138245,I138191);
and I_7643 (I138281,I138074,I138245);
not I_7644 (I138299,I138245);
nand I_7645 (I138317,I138074,I138299);
nor I_7646 (I138335,I138038,I138245);
not I_7647 (I138353,I137912);
nor I_7648 (I138371,I138353,I137957);
nand I_7649 (I138389,I138371,I138191);
nor I_7650 (I138407,I138101,I138389);
nor I_7651 (I138425,I138353,I137822);
and I_7652 (I138443,I138425,I137732);
or I_7653 (I138461,I138443,I138002);
DFFARX1 I_7654 (I138461,I691,I138011,I138488,);
nor I_7655 (I138497,I138488,I138209);
DFFARX1 I_7656 (I138497,I691,I138011,I138524,);
DFFARX1 I_7657 (I138488,I691,I138011,I138542,);
not I_7658 (I138551,I138488);
nor I_7659 (I138569,I138551,I138074);
nor I_7660 (I138587,I138371,I138569);
DFFARX1 I_7661 (I138587,I691,I138011,I138614,);
not I_7662 (I138623,I698);
DFFARX1 I_7663 (I138263,I691,I138623,I138650,);
not I_7664 (I138659,I138650);
nand I_7665 (I138677,I138524,I138614);
and I_7666 (I138695,I138677,I138317);
DFFARX1 I_7667 (I138695,I691,I138623,I138722,);
DFFARX1 I_7668 (I138722,I691,I138623,I138740,);
DFFARX1 I_7669 (I138335,I691,I138623,I138758,);
nand I_7670 (I138767,I138758,I138407);
not I_7671 (I138785,I138767);
DFFARX1 I_7672 (I138785,I691,I138623,I138812,);
not I_7673 (I138821,I138812);
nor I_7674 (I138839,I138659,I138821);
DFFARX1 I_7675 (I138182,I691,I138623,I138866,);
nor I_7676 (I138875,I138866,I138722);
nor I_7677 (I138893,I138866,I138785);
nand I_7678 (I138911,I138524,I138335);
and I_7679 (I138929,I138911,I138542);
DFFARX1 I_7680 (I138929,I691,I138623,I138956,);
not I_7681 (I138965,I138956);
nand I_7682 (I138983,I138965,I138866);
nand I_7683 (I139001,I138965,I138767);
nor I_7684 (I139019,I138281,I138335);
and I_7685 (I139037,I138866,I139019);
nor I_7686 (I139055,I138965,I139037);
DFFARX1 I_7687 (I139055,I691,I138623,I139082,);
nor I_7688 (I139091,I138650,I139019);
DFFARX1 I_7689 (I139091,I691,I138623,I139118,);
nor I_7690 (I139127,I138956,I139019);
not I_7691 (I139145,I139127);
nand I_7692 (I139163,I139145,I138983);
not I_7693 (I139181,I698);
DFFARX1 I_7694 (I138893,I691,I139181,I139208,);
nand I_7695 (I139217,I139001,I139118);
and I_7696 (I139235,I139217,I138875);
DFFARX1 I_7697 (I139235,I691,I139181,I139262,);
nor I_7698 (I139271,I139262,I139208);
not I_7699 (I139289,I139262);
DFFARX1 I_7700 (I139082,I691,I139181,I139316,);
nand I_7701 (I139325,I139316,I139001);
not I_7702 (I139343,I139325);
DFFARX1 I_7703 (I139343,I691,I139181,I139370,);
not I_7704 (I139379,I139370);
nor I_7705 (I139397,I139208,I139325);
nor I_7706 (I139415,I139262,I139397);
DFFARX1 I_7707 (I138740,I691,I139181,I139442,);
DFFARX1 I_7708 (I139442,I691,I139181,I139460,);
not I_7709 (I139469,I139460);
not I_7710 (I139487,I139442);
nand I_7711 (I139505,I139487,I139289);
nand I_7712 (I139523,I139118,I139163);
and I_7713 (I139541,I139523,I138893);
DFFARX1 I_7714 (I139541,I691,I139181,I139568,);
nor I_7715 (I139577,I139568,I139208);
DFFARX1 I_7716 (I139577,I691,I139181,I139604,);
DFFARX1 I_7717 (I139568,I691,I139181,I139622,);
nor I_7718 (I139631,I138839,I139163);
not I_7719 (I139649,I139631);
nor I_7720 (I139667,I139469,I139649);
nand I_7721 (I139685,I139487,I139649);
nor I_7722 (I139703,I139208,I139631);
DFFARX1 I_7723 (I139631,I691,I139181,I139730,);
not I_7724 (I139739,I698);
DFFARX1 I_7725 (I139379,I691,I139739,I139766,);
not I_7726 (I139775,I139766);
nand I_7727 (I139793,I139415,I139730);
and I_7728 (I139811,I139793,I139604);
DFFARX1 I_7729 (I139811,I691,I139739,I139838,);
DFFARX1 I_7730 (I139271,I691,I139739,I139856,);
and I_7731 (I139865,I139856,I139622);
nor I_7732 (I139883,I139838,I139865);
DFFARX1 I_7733 (I139883,I691,I139739,I139910,);
nand I_7734 (I139919,I139856,I139622);
nand I_7735 (I139937,I139775,I139919);
not I_7736 (I139955,I139937);
DFFARX1 I_7737 (I139667,I691,I139739,I139982,);
DFFARX1 I_7738 (I139982,I691,I139739,I140000,);
nand I_7739 (I140009,I139604,I139505);
and I_7740 (I140027,I140009,I139685);
DFFARX1 I_7741 (I140027,I691,I139739,I140054,);
DFFARX1 I_7742 (I140054,I691,I139739,I140072,);
not I_7743 (I140081,I140072);
not I_7744 (I140099,I140054);
nand I_7745 (I140117,I140099,I139919);
nor I_7746 (I140135,I139703,I139505);
not I_7747 (I140153,I140135);
nor I_7748 (I140171,I140099,I140153);
nor I_7749 (I140189,I139775,I140171);
DFFARX1 I_7750 (I140189,I691,I139739,I140216,);
nor I_7751 (I140225,I139838,I140153);
nor I_7752 (I140243,I140054,I140225);
nor I_7753 (I140261,I139982,I140135);
nor I_7754 (I140279,I139838,I140135);
not I_7755 (I140297,I698);
DFFARX1 I_7756 (I140000,I691,I140297,I140324,);
nand I_7757 (I140333,I140324,I140279);
DFFARX1 I_7758 (I139910,I691,I140297,I140360,);
DFFARX1 I_7759 (I140360,I691,I140297,I140378,);
not I_7760 (I140387,I140378);
not I_7761 (I140405,I140216);
nor I_7762 (I140423,I140216,I139955);
not I_7763 (I140441,I139910);
nand I_7764 (I140459,I140405,I140441);
nor I_7765 (I140477,I139910,I140216);
and I_7766 (I140495,I140477,I140333);
not I_7767 (I140513,I140117);
nand I_7768 (I140531,I140513,I140261);
nor I_7769 (I140549,I140117,I140279);
not I_7770 (I140567,I140549);
nand I_7771 (I140585,I140423,I140567);
DFFARX1 I_7772 (I140549,I691,I140297,I140612,);
nor I_7773 (I140621,I140243,I139910);
nor I_7774 (I140639,I140621,I139955);
and I_7775 (I140657,I140639,I140531);
DFFARX1 I_7776 (I140657,I691,I140297,I140684,);
nor I_7777 (I140693,I140621,I140459);
or I_7778 (I140711,I140549,I140621);
nor I_7779 (I140729,I140243,I140081);
DFFARX1 I_7780 (I140729,I691,I140297,I140756,);
not I_7781 (I140765,I140756);
nand I_7782 (I140783,I140765,I140405);
nor I_7783 (I140801,I140783,I139955);
DFFARX1 I_7784 (I140801,I691,I140297,I140828,);
nor I_7785 (I140837,I140765,I140459);
nor I_7786 (I140855,I140621,I140837);
not I_7787 (I140873,I698);
DFFARX1 I_7788 (I140693,I691,I140873,I140900,);
nand I_7789 (I140909,I140900,I140387);
not I_7790 (I140927,I140909);
DFFARX1 I_7791 (I140828,I691,I140873,I140954,);
not I_7792 (I140963,I140954);
not I_7793 (I140981,I140495);
or I_7794 (I140999,I140828,I140495);
nor I_7795 (I141017,I140828,I140495);
or I_7796 (I141035,I140684,I140828);
DFFARX1 I_7797 (I141035,I691,I140873,I141062,);
not I_7798 (I141071,I140585);
nand I_7799 (I141089,I141071,I140612);
nand I_7800 (I141107,I140981,I141089);
and I_7801 (I141125,I140963,I141107);
nor I_7802 (I141143,I140585,I140855);
and I_7803 (I141161,I140963,I141143);
nor I_7804 (I141179,I140927,I141161);
DFFARX1 I_7805 (I141143,I691,I140873,I141206,);
not I_7806 (I141215,I141206);
nor I_7807 (I141233,I140963,I141215);
or I_7808 (I141251,I141035,I140711);
nor I_7809 (I141269,I140711,I140684);
nand I_7810 (I141287,I141107,I141269);
nand I_7811 (I141305,I141251,I141287);
DFFARX1 I_7812 (I141305,I691,I140873,I141332,);
nor I_7813 (I141341,I141269,I140999);
DFFARX1 I_7814 (I141341,I691,I140873,I141368,);
nor I_7815 (I141377,I140711,I140495);
DFFARX1 I_7816 (I141377,I691,I140873,I141404,);
DFFARX1 I_7817 (I141404,I691,I140873,I141422,);
not I_7818 (I141431,I141404);
nand I_7819 (I141449,I141431,I140909);
nand I_7820 (I141467,I141431,I141017);
not I_7821 (I141485,I698);
DFFARX1 I_7822 (I92,I691,I141485,I141512,);
not I_7823 (I141521,I141512);
DFFARX1 I_7824 (I372,I691,I141485,I141548,);
not I_7825 (I141557,I604);
nand I_7826 (I141575,I141557,I428);
not I_7827 (I141593,I141575);
nor I_7828 (I141611,I141593,I556);
nor I_7829 (I141629,I141521,I141611);
DFFARX1 I_7830 (I141629,I691,I141485,I141656,);
not I_7831 (I141665,I556);
nand I_7832 (I141683,I141665,I141593);
and I_7833 (I141701,I141665,I180);
nand I_7834 (I141719,I141701,I612);
nor I_7835 (I141737,I141719,I141665);
and I_7836 (I141755,I141548,I141719);
not I_7837 (I141773,I141719);
nand I_7838 (I141791,I141548,I141773);
nor I_7839 (I141809,I141512,I141719);
not I_7840 (I141827,I668);
nor I_7841 (I141845,I141827,I180);
nand I_7842 (I141863,I141845,I141665);
nor I_7843 (I141881,I141575,I141863);
nor I_7844 (I141899,I141827,I364);
and I_7845 (I141917,I141899,I524);
or I_7846 (I141935,I141917,I628);
DFFARX1 I_7847 (I141935,I691,I141485,I141962,);
nor I_7848 (I141971,I141962,I141683);
DFFARX1 I_7849 (I141971,I691,I141485,I141998,);
DFFARX1 I_7850 (I141962,I691,I141485,I142016,);
not I_7851 (I142025,I141962);
nor I_7852 (I142043,I142025,I141548);
nor I_7853 (I142061,I141845,I142043);
DFFARX1 I_7854 (I142061,I691,I141485,I142088,);
not I_7855 (I142097,I698);
DFFARX1 I_7856 (I141737,I691,I142097,I142124,);
DFFARX1 I_7857 (I142124,I691,I142097,I142142,);
not I_7858 (I142151,I142142);
nand I_7859 (I142169,I141998,I141656);
and I_7860 (I142187,I142169,I141881);
DFFARX1 I_7861 (I142187,I691,I142097,I142214,);
DFFARX1 I_7862 (I142214,I691,I142097,I142232,);
DFFARX1 I_7863 (I142214,I691,I142097,I142250,);
DFFARX1 I_7864 (I141791,I691,I142097,I142268,);
nand I_7865 (I142277,I142268,I141998);
not I_7866 (I142295,I142277);
nor I_7867 (I142313,I142124,I142295);
DFFARX1 I_7868 (I141809,I691,I142097,I142340,);
not I_7869 (I142349,I142340);
nor I_7870 (I142367,I142349,I142151);
nand I_7871 (I142385,I142349,I142277);
nand I_7872 (I142403,I142016,I141755);
and I_7873 (I142421,I142403,I142088);
DFFARX1 I_7874 (I142421,I691,I142097,I142448,);
nor I_7875 (I142457,I142448,I142124);
DFFARX1 I_7876 (I142457,I691,I142097,I142484,);
not I_7877 (I142493,I142448);
nor I_7878 (I142511,I141809,I141755);
not I_7879 (I142529,I142511);
nor I_7880 (I142547,I142277,I142529);
nor I_7881 (I142565,I142493,I142547);
DFFARX1 I_7882 (I142565,I691,I142097,I142592,);
nor I_7883 (I142601,I142448,I142529);
nor I_7884 (I142619,I142295,I142601);
nor I_7885 (I142637,I142448,I142511);
not I_7886 (I142655,I698);
DFFARX1 I_7887 (I142385,I691,I142655,I142682,);
nand I_7888 (I142691,I142682,I142484);
not I_7889 (I142709,I142691);
DFFARX1 I_7890 (I142367,I691,I142655,I142736,);
not I_7891 (I142745,I142736);
not I_7892 (I142763,I142592);
or I_7893 (I142781,I142250,I142592);
nor I_7894 (I142799,I142250,I142592);
or I_7895 (I142817,I142619,I142250);
DFFARX1 I_7896 (I142817,I691,I142655,I142844,);
not I_7897 (I142853,I142313);
nand I_7898 (I142871,I142853,I142232);
nand I_7899 (I142889,I142763,I142871);
and I_7900 (I142907,I142745,I142889);
nor I_7901 (I142925,I142313,I142637);
and I_7902 (I142943,I142745,I142925);
nor I_7903 (I142961,I142709,I142943);
DFFARX1 I_7904 (I142925,I691,I142655,I142988,);
not I_7905 (I142997,I142988);
nor I_7906 (I143015,I142745,I142997);
or I_7907 (I143033,I142817,I142637);
nor I_7908 (I143051,I142637,I142619);
nand I_7909 (I143069,I142889,I143051);
nand I_7910 (I143087,I143033,I143069);
DFFARX1 I_7911 (I143087,I691,I142655,I143114,);
nor I_7912 (I143123,I143051,I142781);
DFFARX1 I_7913 (I143123,I691,I142655,I143150,);
nor I_7914 (I143159,I142637,I142484);
DFFARX1 I_7915 (I143159,I691,I142655,I143186,);
DFFARX1 I_7916 (I143186,I691,I142655,I143204,);
not I_7917 (I143213,I143186);
nand I_7918 (I143231,I143213,I142691);
nand I_7919 (I143249,I143213,I142799);
not I_7920 (I143267,I698);
DFFARX1 I_7921 (I142961,I691,I143267,I143294,);
nand I_7922 (I143303,I143294,I143015);
DFFARX1 I_7923 (I143114,I691,I143267,I143330,);
DFFARX1 I_7924 (I143330,I691,I143267,I143348,);
not I_7925 (I143357,I143348);
not I_7926 (I143375,I143204);
nor I_7927 (I143393,I143204,I143231);
not I_7928 (I143411,I143249);
nand I_7929 (I143429,I143375,I143411);
nor I_7930 (I143447,I143249,I143204);
and I_7931 (I143465,I143447,I143303);
not I_7932 (I143483,I142907);
nand I_7933 (I143501,I143483,I143150);
nor I_7934 (I143519,I142907,I143150);
not I_7935 (I143537,I143519);
nand I_7936 (I143555,I143393,I143537);
DFFARX1 I_7937 (I143519,I691,I143267,I143582,);
nor I_7938 (I143591,I142907,I143249);
nor I_7939 (I143609,I143591,I143231);
and I_7940 (I143627,I143609,I143501);
DFFARX1 I_7941 (I143627,I691,I143267,I143654,);
nor I_7942 (I143663,I143591,I143429);
or I_7943 (I143681,I143519,I143591);
nor I_7944 (I143699,I142907,I142844);
DFFARX1 I_7945 (I143699,I691,I143267,I143726,);
not I_7946 (I143735,I143726);
nand I_7947 (I143753,I143735,I143375);
nor I_7948 (I143771,I143753,I143231);
DFFARX1 I_7949 (I143771,I691,I143267,I143798,);
nor I_7950 (I143807,I143735,I143429);
nor I_7951 (I143825,I143591,I143807);
not I_7952 (I143843,I698);
DFFARX1 I_7953 (I143654,I691,I143843,I143870,);
DFFARX1 I_7954 (I143870,I691,I143843,I143888,);
not I_7955 (I143897,I143888);
not I_7956 (I143915,I143870);
DFFARX1 I_7957 (I143465,I691,I143843,I143942,);
not I_7958 (I143951,I143942);
and I_7959 (I143969,I143915,I143582);
not I_7960 (I143987,I143465);
nand I_7961 (I144005,I143987,I143582);
not I_7962 (I144023,I143357);
nor I_7963 (I144041,I144023,I143663);
nand I_7964 (I144059,I144041,I143681);
nor I_7965 (I144077,I144059,I144005);
DFFARX1 I_7966 (I144077,I691,I143843,I144104,);
not I_7967 (I144113,I144059);
not I_7968 (I144131,I143663);
nand I_7969 (I144149,I144131,I143582);
nor I_7970 (I144167,I143663,I143465);
nand I_7971 (I144185,I143969,I144167);
nand I_7972 (I144203,I143915,I143663);
nand I_7973 (I144221,I144023,I143825);
DFFARX1 I_7974 (I144221,I691,I143843,I144248,);
DFFARX1 I_7975 (I144221,I691,I143843,I144266,);
not I_7976 (I144275,I143825);
nor I_7977 (I144293,I144275,I143798);
and I_7978 (I144311,I144293,I143555);
or I_7979 (I144329,I144311,I143798);
DFFARX1 I_7980 (I144329,I691,I143843,I144356,);
nand I_7981 (I144365,I144356,I143987);
nor I_7982 (I144383,I144365,I144149);
nor I_7983 (I144401,I144356,I143951);
DFFARX1 I_7984 (I144356,I691,I143843,I144428,);
not I_7985 (I144437,I144428);
nor I_7986 (I144455,I144437,I144113);
not I_7987 (I144473,I698);
DFFARX1 I_7988 (I144104,I691,I144473,I144500,);
nand I_7989 (I144509,I144104,I144203);
and I_7990 (I144527,I144509,I143897);
DFFARX1 I_7991 (I144527,I691,I144473,I144554,);
nor I_7992 (I144563,I144554,I144500);
not I_7993 (I144581,I144554);
DFFARX1 I_7994 (I144185,I691,I144473,I144608,);
nand I_7995 (I144617,I144608,I144383);
not I_7996 (I144635,I144617);
DFFARX1 I_7997 (I144635,I691,I144473,I144662,);
not I_7998 (I144671,I144662);
nor I_7999 (I144689,I144500,I144617);
nor I_8000 (I144707,I144554,I144689);
DFFARX1 I_8001 (I144455,I691,I144473,I144734,);
DFFARX1 I_8002 (I144734,I691,I144473,I144752,);
not I_8003 (I144761,I144752);
not I_8004 (I144779,I144734);
nand I_8005 (I144797,I144779,I144581);
nand I_8006 (I144815,I144401,I144401);
and I_8007 (I144833,I144815,I144248);
DFFARX1 I_8008 (I144833,I691,I144473,I144860,);
nor I_8009 (I144869,I144860,I144500);
DFFARX1 I_8010 (I144869,I691,I144473,I144896,);
DFFARX1 I_8011 (I144860,I691,I144473,I144914,);
nor I_8012 (I144923,I144266,I144401);
not I_8013 (I144941,I144923);
nor I_8014 (I144959,I144761,I144941);
nand I_8015 (I144977,I144779,I144941);
nor I_8016 (I144995,I144500,I144923);
DFFARX1 I_8017 (I144923,I691,I144473,I145022,);
not I_8018 (I145031,I698);
DFFARX1 I_8019 (I144671,I691,I145031,I145058,);
not I_8020 (I145067,I145058);
nand I_8021 (I145085,I144707,I145022);
and I_8022 (I145103,I145085,I144896);
DFFARX1 I_8023 (I145103,I691,I145031,I145130,);
DFFARX1 I_8024 (I144563,I691,I145031,I145148,);
and I_8025 (I145157,I145148,I144914);
nor I_8026 (I145175,I145130,I145157);
DFFARX1 I_8027 (I145175,I691,I145031,I145202,);
nand I_8028 (I145211,I145148,I144914);
nand I_8029 (I145229,I145067,I145211);
not I_8030 (I145247,I145229);
DFFARX1 I_8031 (I144959,I691,I145031,I145274,);
DFFARX1 I_8032 (I145274,I691,I145031,I145292,);
nand I_8033 (I145301,I144896,I144797);
and I_8034 (I145319,I145301,I144977);
DFFARX1 I_8035 (I145319,I691,I145031,I145346,);
DFFARX1 I_8036 (I145346,I691,I145031,I145364,);
not I_8037 (I145373,I145364);
not I_8038 (I145391,I145346);
nand I_8039 (I145409,I145391,I145211);
nor I_8040 (I145427,I144995,I144797);
not I_8041 (I145445,I145427);
nor I_8042 (I145463,I145391,I145445);
nor I_8043 (I145481,I145067,I145463);
DFFARX1 I_8044 (I145481,I691,I145031,I145508,);
nor I_8045 (I145517,I145130,I145445);
nor I_8046 (I145535,I145346,I145517);
nor I_8047 (I145553,I145274,I145427);
nor I_8048 (I145571,I145130,I145427);
not I_8049 (I145589,I698);
DFFARX1 I_8050 (I145373,I691,I145589,I145616,);
not I_8051 (I145625,I145616);
nand I_8052 (I145643,I145202,I145409);
and I_8053 (I145661,I145643,I145571);
DFFARX1 I_8054 (I145661,I691,I145589,I145688,);
DFFARX1 I_8055 (I145688,I691,I145589,I145706,);
DFFARX1 I_8056 (I145292,I691,I145589,I145724,);
nand I_8057 (I145733,I145724,I145247);
not I_8058 (I145751,I145733);
DFFARX1 I_8059 (I145751,I691,I145589,I145778,);
not I_8060 (I145787,I145778);
nor I_8061 (I145805,I145625,I145787);
DFFARX1 I_8062 (I145535,I691,I145589,I145832,);
nor I_8063 (I145841,I145832,I145688);
nor I_8064 (I145859,I145832,I145751);
nand I_8065 (I145877,I145508,I145553);
and I_8066 (I145895,I145877,I145571);
DFFARX1 I_8067 (I145895,I691,I145589,I145922,);
not I_8068 (I145931,I145922);
nand I_8069 (I145949,I145931,I145832);
nand I_8070 (I145967,I145931,I145733);
nor I_8071 (I145985,I145202,I145553);
and I_8072 (I146003,I145832,I145985);
nor I_8073 (I146021,I145931,I146003);
DFFARX1 I_8074 (I146021,I691,I145589,I146048,);
nor I_8075 (I146057,I145616,I145985);
DFFARX1 I_8076 (I146057,I691,I145589,I146084,);
nor I_8077 (I146093,I145922,I145985);
not I_8078 (I146111,I146093);
nand I_8079 (I146129,I146111,I145949);
not I_8080 (I146147,I698);
DFFARX1 I_8081 (I146048,I691,I146147,I146174,);
not I_8082 (I146183,I146174);
nand I_8083 (I146201,I145859,I145805);
and I_8084 (I146219,I146201,I145706);
DFFARX1 I_8085 (I146219,I691,I146147,I146246,);
not I_8086 (I146255,I146129);
DFFARX1 I_8087 (I145967,I691,I146147,I146282,);
not I_8088 (I146291,I146282);
nor I_8089 (I146309,I146291,I146183);
and I_8090 (I146327,I146309,I146129);
nor I_8091 (I146345,I146291,I146255);
nor I_8092 (I146363,I146246,I146345);
DFFARX1 I_8093 (I146084,I691,I146147,I146390,);
nor I_8094 (I146399,I146390,I146246);
not I_8095 (I146417,I146399);
not I_8096 (I146435,I146390);
nor I_8097 (I146453,I146435,I146327);
DFFARX1 I_8098 (I146453,I691,I146147,I146480,);
nand I_8099 (I146489,I146084,I145859);
and I_8100 (I146507,I146489,I145967);
DFFARX1 I_8101 (I146507,I691,I146147,I146534,);
nor I_8102 (I146543,I146534,I146390);
DFFARX1 I_8103 (I146543,I691,I146147,I146570,);
nand I_8104 (I146579,I146534,I146435);
nand I_8105 (I146597,I146417,I146579);
not I_8106 (I146615,I146534);
nor I_8107 (I146633,I146615,I146327);
DFFARX1 I_8108 (I146633,I691,I146147,I146660,);
nor I_8109 (I146669,I145841,I145859);
or I_8110 (I146687,I146390,I146669);
nor I_8111 (I146705,I146534,I146669);
or I_8112 (I146723,I146246,I146669);
DFFARX1 I_8113 (I146669,I691,I146147,I146750,);
not I_8114 (I146759,I698);
DFFARX1 I_8115 (I146363,I691,I146759,I146786,);
and I_8116 (I146795,I146786,I146705);
DFFARX1 I_8117 (I146795,I691,I146759,I146822,);
DFFARX1 I_8118 (I146723,I691,I146759,I146840,);
not I_8119 (I146849,I146570);
not I_8120 (I146867,I146750);
nand I_8121 (I146885,I146867,I146849);
nor I_8122 (I146903,I146840,I146885);
DFFARX1 I_8123 (I146885,I691,I146759,I146930,);
not I_8124 (I146939,I146930);
not I_8125 (I146957,I146687);
nand I_8126 (I146975,I146867,I146957);
DFFARX1 I_8127 (I146975,I691,I146759,I147002,);
not I_8128 (I147011,I147002);
not I_8129 (I147029,I146660);
nand I_8130 (I147047,I147029,I146480);
and I_8131 (I147065,I146849,I147047);
nor I_8132 (I147083,I146975,I147065);
DFFARX1 I_8133 (I147083,I691,I146759,I147110,);
DFFARX1 I_8134 (I147065,I691,I146759,I147128,);
nor I_8135 (I147137,I146660,I146597);
nor I_8136 (I147155,I146975,I147137);
or I_8137 (I147173,I146660,I146597);
nor I_8138 (I147191,I146570,I146705);
DFFARX1 I_8139 (I147191,I691,I146759,I147218,);
not I_8140 (I147227,I147218);
nor I_8141 (I147245,I147227,I147011);
nand I_8142 (I147263,I147227,I146840);
not I_8143 (I147281,I146570);
nand I_8144 (I147299,I147281,I146957);
nand I_8145 (I147317,I147227,I147299);
nand I_8146 (I147335,I147317,I147263);
nand I_8147 (I147353,I147299,I147173);
not I_8148 (I147371,I698);
DFFARX1 I_8149 (I147245,I691,I147371,I147398,);
not I_8150 (I147407,I147398);
nand I_8151 (I147425,I147110,I147110);
and I_8152 (I147443,I147425,I147353);
DFFARX1 I_8153 (I147443,I691,I147371,I147470,);
DFFARX1 I_8154 (I147470,I691,I147371,I147488,);
DFFARX1 I_8155 (I146903,I691,I147371,I147506,);
nand I_8156 (I147515,I147506,I147155);
not I_8157 (I147533,I147515);
DFFARX1 I_8158 (I147533,I691,I147371,I147560,);
not I_8159 (I147569,I147560);
nor I_8160 (I147587,I147407,I147569);
DFFARX1 I_8161 (I146939,I691,I147371,I147614,);
nor I_8162 (I147623,I147614,I147470);
nor I_8163 (I147641,I147614,I147533);
nand I_8164 (I147659,I146822,I147335);
and I_8165 (I147677,I147659,I146903);
DFFARX1 I_8166 (I147677,I691,I147371,I147704,);
not I_8167 (I147713,I147704);
nand I_8168 (I147731,I147713,I147614);
nand I_8169 (I147749,I147713,I147515);
nor I_8170 (I147767,I147128,I147335);
and I_8171 (I147785,I147614,I147767);
nor I_8172 (I147803,I147713,I147785);
DFFARX1 I_8173 (I147803,I691,I147371,I147830,);
nor I_8174 (I147839,I147398,I147767);
DFFARX1 I_8175 (I147839,I691,I147371,I147866,);
nor I_8176 (I147875,I147704,I147767);
not I_8177 (I147893,I147875);
nand I_8178 (I147911,I147893,I147731);
not I_8179 (I147929,I698);
DFFARX1 I_8180 (I147641,I691,I147929,I147956,);
and I_8181 (I147965,I147956,I147911);
DFFARX1 I_8182 (I147965,I691,I147929,I147992,);
DFFARX1 I_8183 (I147830,I691,I147929,I148010,);
not I_8184 (I148019,I147866);
not I_8185 (I148037,I147866);
nand I_8186 (I148055,I148037,I148019);
nor I_8187 (I148073,I148010,I148055);
DFFARX1 I_8188 (I148055,I691,I147929,I148100,);
not I_8189 (I148109,I148100);
not I_8190 (I148127,I147488);
nand I_8191 (I148145,I148037,I148127);
DFFARX1 I_8192 (I148145,I691,I147929,I148172,);
not I_8193 (I148181,I148172);
not I_8194 (I148199,I147623);
nand I_8195 (I148217,I148199,I147641);
and I_8196 (I148235,I148019,I148217);
nor I_8197 (I148253,I148145,I148235);
DFFARX1 I_8198 (I148253,I691,I147929,I148280,);
DFFARX1 I_8199 (I148235,I691,I147929,I148298,);
nor I_8200 (I148307,I147623,I147587);
nor I_8201 (I148325,I148145,I148307);
or I_8202 (I148343,I147623,I147587);
nor I_8203 (I148361,I147749,I147749);
DFFARX1 I_8204 (I148361,I691,I147929,I148388,);
not I_8205 (I148397,I148388);
nor I_8206 (I148415,I148397,I148181);
nand I_8207 (I148433,I148397,I148010);
not I_8208 (I148451,I147749);
nand I_8209 (I148469,I148451,I148127);
nand I_8210 (I148487,I148397,I148469);
nand I_8211 (I148505,I148487,I148433);
nand I_8212 (I148523,I148469,I148343);
not I_8213 (I148541,I698);
DFFARX1 I_8214 (I148280,I691,I148541,I148568,);
nand I_8215 (I148577,I147992,I148280);
and I_8216 (I148595,I148577,I148415);
DFFARX1 I_8217 (I148595,I691,I148541,I148622,);
nor I_8218 (I148631,I148622,I148568);
not I_8219 (I148649,I148622);
DFFARX1 I_8220 (I148109,I691,I148541,I148676,);
nand I_8221 (I148685,I148676,I148523);
not I_8222 (I148703,I148685);
DFFARX1 I_8223 (I148703,I691,I148541,I148730,);
not I_8224 (I148739,I148730);
nor I_8225 (I148757,I148568,I148685);
nor I_8226 (I148775,I148622,I148757);
DFFARX1 I_8227 (I148073,I691,I148541,I148802,);
DFFARX1 I_8228 (I148802,I691,I148541,I148820,);
not I_8229 (I148829,I148820);
not I_8230 (I148847,I148802);
nand I_8231 (I148865,I148847,I148649);
nand I_8232 (I148883,I148073,I148505);
and I_8233 (I148901,I148883,I148298);
DFFARX1 I_8234 (I148901,I691,I148541,I148928,);
nor I_8235 (I148937,I148928,I148568);
DFFARX1 I_8236 (I148937,I691,I148541,I148964,);
DFFARX1 I_8237 (I148928,I691,I148541,I148982,);
nor I_8238 (I148991,I148325,I148505);
not I_8239 (I149009,I148991);
nor I_8240 (I149027,I148829,I149009);
nand I_8241 (I149045,I148847,I149009);
nor I_8242 (I149063,I148568,I148991);
DFFARX1 I_8243 (I148991,I691,I148541,I149090,);
not I_8244 (I149099,I698);
DFFARX1 I_8245 (I148964,I691,I149099,I149126,);
DFFARX1 I_8246 (I149045,I691,I149099,I149144,);
not I_8247 (I149153,I149144);
not I_8248 (I149171,I148739);
nor I_8249 (I149189,I149171,I149063);
not I_8250 (I149207,I149090);
nor I_8251 (I149225,I149189,I148775);
nor I_8252 (I149243,I149144,I149225);
DFFARX1 I_8253 (I149243,I691,I149099,I149270,);
nor I_8254 (I149279,I148775,I149063);
nand I_8255 (I149297,I149279,I148739);
DFFARX1 I_8256 (I149297,I691,I149099,I149324,);
nor I_8257 (I149333,I149207,I148775);
nand I_8258 (I149351,I149333,I148964);
nor I_8259 (I149369,I149126,I149351);
DFFARX1 I_8260 (I149369,I691,I149099,I149396,);
not I_8261 (I149405,I149351);
nand I_8262 (I149423,I149144,I149405);
DFFARX1 I_8263 (I149351,I691,I149099,I149450,);
not I_8264 (I149459,I149450);
not I_8265 (I149477,I148775);
not I_8266 (I149495,I148865);
nor I_8267 (I149513,I149495,I149090);
nor I_8268 (I149531,I149459,I149513);
nor I_8269 (I149549,I149495,I149027);
and I_8270 (I149567,I149549,I148631);
or I_8271 (I149585,I149567,I148982);
DFFARX1 I_8272 (I149585,I691,I149099,I149612,);
nor I_8273 (I149621,I149612,I149126);
not I_8274 (I149639,I149612);
and I_8275 (I149657,I149639,I149126);
nor I_8276 (I149675,I149153,I149657);
nand I_8277 (I149693,I149639,I149207);
nor I_8278 (I149711,I149495,I149693);
nand I_8279 (I149729,I149639,I149405);
nand I_8280 (I149747,I149207,I148865);
nor I_8281 (I149765,I149477,I149747);
not I_8282 (I149783,I698);
DFFARX1 I_8283 (I149675,I691,I149783,I149810,);
not I_8284 (I149819,I149810);
nand I_8285 (I149837,I149531,I149270);
and I_8286 (I149855,I149837,I149396);
DFFARX1 I_8287 (I149855,I691,I149783,I149882,);
DFFARX1 I_8288 (I149765,I691,I149783,I149900,);
and I_8289 (I149909,I149900,I149711);
nor I_8290 (I149927,I149882,I149909);
DFFARX1 I_8291 (I149927,I691,I149783,I149954,);
nand I_8292 (I149963,I149900,I149711);
nand I_8293 (I149981,I149819,I149963);
not I_8294 (I149999,I149981);
DFFARX1 I_8295 (I149621,I691,I149783,I150026,);
DFFARX1 I_8296 (I150026,I691,I149783,I150044,);
nand I_8297 (I150053,I149324,I149423);
and I_8298 (I150071,I150053,I149729);
DFFARX1 I_8299 (I150071,I691,I149783,I150098,);
DFFARX1 I_8300 (I150098,I691,I149783,I150116,);
not I_8301 (I150125,I150116);
not I_8302 (I150143,I150098);
nand I_8303 (I150161,I150143,I149963);
nor I_8304 (I150179,I149396,I149423);
not I_8305 (I150197,I150179);
nor I_8306 (I150215,I150143,I150197);
nor I_8307 (I150233,I149819,I150215);
DFFARX1 I_8308 (I150233,I691,I149783,I150260,);
nor I_8309 (I150269,I149882,I150197);
nor I_8310 (I150287,I150098,I150269);
nor I_8311 (I150305,I150026,I150179);
nor I_8312 (I150323,I149882,I150179);
not I_8313 (I150341,I698);
DFFARX1 I_8314 (I150323,I691,I150341,I150368,);
not I_8315 (I150377,I150368);
nand I_8316 (I150395,I149999,I150044);
and I_8317 (I150413,I150395,I149954);
DFFARX1 I_8318 (I150413,I691,I150341,I150440,);
not I_8319 (I150449,I150323);
DFFARX1 I_8320 (I150260,I691,I150341,I150476,);
not I_8321 (I150485,I150476);
nor I_8322 (I150503,I150485,I150377);
and I_8323 (I150521,I150503,I150323);
nor I_8324 (I150539,I150485,I150449);
nor I_8325 (I150557,I150440,I150539);
DFFARX1 I_8326 (I150161,I691,I150341,I150584,);
nor I_8327 (I150593,I150584,I150440);
not I_8328 (I150611,I150593);
not I_8329 (I150629,I150584);
nor I_8330 (I150647,I150629,I150521);
DFFARX1 I_8331 (I150647,I691,I150341,I150674,);
nand I_8332 (I150683,I150125,I149954);
and I_8333 (I150701,I150683,I150287);
DFFARX1 I_8334 (I150701,I691,I150341,I150728,);
nor I_8335 (I150737,I150728,I150584);
DFFARX1 I_8336 (I150737,I691,I150341,I150764,);
nand I_8337 (I150773,I150728,I150629);
nand I_8338 (I150791,I150611,I150773);
not I_8339 (I150809,I150728);
nor I_8340 (I150827,I150809,I150521);
DFFARX1 I_8341 (I150827,I691,I150341,I150854,);
nor I_8342 (I150863,I150305,I149954);
or I_8343 (I150881,I150584,I150863);
nor I_8344 (I150899,I150728,I150863);
or I_8345 (I150917,I150440,I150863);
DFFARX1 I_8346 (I150863,I691,I150341,I150944,);
not I_8347 (I150953,I698);
DFFARX1 I_8348 (I150899,I691,I150953,I150980,);
DFFARX1 I_8349 (I150980,I691,I150953,I150998,);
not I_8350 (I151007,I150998);
not I_8351 (I151025,I150980);
nand I_8352 (I151043,I150944,I150557);
and I_8353 (I151061,I151043,I150899);
DFFARX1 I_8354 (I151061,I691,I150953,I151088,);
not I_8355 (I151097,I151088);
DFFARX1 I_8356 (I150791,I691,I150953,I151124,);
and I_8357 (I151133,I151124,I150917);
nand I_8358 (I151151,I151124,I150917);
nand I_8359 (I151169,I151097,I151151);
DFFARX1 I_8360 (I150764,I691,I150953,I151196,);
nor I_8361 (I151205,I151196,I151133);
DFFARX1 I_8362 (I151205,I691,I150953,I151232,);
nor I_8363 (I151241,I151196,I151088);
nand I_8364 (I151259,I150764,I150881);
and I_8365 (I151277,I151259,I150854);
DFFARX1 I_8366 (I151277,I691,I150953,I151304,);
nor I_8367 (I151313,I151304,I151196);
not I_8368 (I151331,I151304);
nor I_8369 (I151349,I151331,I151097);
nor I_8370 (I151367,I151025,I151349);
DFFARX1 I_8371 (I151367,I691,I150953,I151394,);
nor I_8372 (I151403,I151331,I151196);
nor I_8373 (I151421,I150674,I150881);
nor I_8374 (I151439,I151421,I151403);
not I_8375 (I151457,I151421);
nand I_8376 (I151475,I151151,I151457);
DFFARX1 I_8377 (I151421,I691,I150953,I151502,);
DFFARX1 I_8378 (I151421,I691,I150953,I151520,);
not I_8379 (I151529,I698);
DFFARX1 I_8380 (I151169,I691,I151529,I151556,);
not I_8381 (I151565,I151556);
nand I_8382 (I151583,I151313,I151475);
and I_8383 (I151601,I151583,I151520);
DFFARX1 I_8384 (I151601,I691,I151529,I151628,);
DFFARX1 I_8385 (I151628,I691,I151529,I151646,);
DFFARX1 I_8386 (I151502,I691,I151529,I151664,);
nand I_8387 (I151673,I151664,I151007);
not I_8388 (I151691,I151673);
DFFARX1 I_8389 (I151691,I691,I151529,I151718,);
not I_8390 (I151727,I151718);
nor I_8391 (I151745,I151565,I151727);
DFFARX1 I_8392 (I151232,I691,I151529,I151772,);
nor I_8393 (I151781,I151772,I151628);
nor I_8394 (I151799,I151772,I151691);
nand I_8395 (I151817,I151241,I151394);
and I_8396 (I151835,I151817,I151439);
DFFARX1 I_8397 (I151835,I691,I151529,I151862,);
not I_8398 (I151871,I151862);
nand I_8399 (I151889,I151871,I151772);
nand I_8400 (I151907,I151871,I151673);
nor I_8401 (I151925,I151232,I151394);
and I_8402 (I151943,I151772,I151925);
nor I_8403 (I151961,I151871,I151943);
DFFARX1 I_8404 (I151961,I691,I151529,I151988,);
nor I_8405 (I151997,I151556,I151925);
DFFARX1 I_8406 (I151997,I691,I151529,I152024,);
nor I_8407 (I152033,I151862,I151925);
not I_8408 (I152051,I152033);
nand I_8409 (I152069,I152051,I151889);
not I_8410 (I152087,I698);
DFFARX1 I_8411 (I152069,I691,I152087,I152114,);
DFFARX1 I_8412 (I151907,I691,I152087,I152132,);
not I_8413 (I152141,I152132);
nor I_8414 (I152159,I152114,I152141);
DFFARX1 I_8415 (I152141,I691,I152087,I152186,);
nor I_8416 (I152195,I151745,I151799);
and I_8417 (I152213,I152195,I152024);
nor I_8418 (I152231,I152213,I151745);
not I_8419 (I152249,I151745);
and I_8420 (I152267,I152249,I151907);
nand I_8421 (I152285,I152267,I151646);
nor I_8422 (I152303,I152249,I152285);
DFFARX1 I_8423 (I152303,I691,I152087,I152330,);
not I_8424 (I152339,I152285);
nand I_8425 (I152357,I152141,I152339);
nand I_8426 (I152375,I152213,I152339);
DFFARX1 I_8427 (I152249,I691,I152087,I152402,);
not I_8428 (I152411,I151781);
nor I_8429 (I152429,I152411,I151907);
nor I_8430 (I152447,I152429,I152231);
DFFARX1 I_8431 (I152447,I691,I152087,I152474,);
not I_8432 (I152483,I152429);
DFFARX1 I_8433 (I152483,I691,I152087,I152510,);
not I_8434 (I152519,I152510);
nor I_8435 (I152537,I152519,I152429);
nor I_8436 (I152555,I152411,I152024);
and I_8437 (I152573,I152555,I151988);
or I_8438 (I152591,I152573,I151799);
DFFARX1 I_8439 (I152591,I691,I152087,I152618,);
not I_8440 (I152627,I152618);
nand I_8441 (I152645,I152627,I152339);
not I_8442 (I152663,I152645);
nand I_8443 (I152681,I152645,I152357);
nand I_8444 (I152699,I152627,I152213);
not I_8445 (I152717,I698);
DFFARX1 I_8446 (I152537,I691,I152717,I152744,);
nand I_8447 (I152753,I152330,I152330);
and I_8448 (I152771,I152753,I152402);
DFFARX1 I_8449 (I152771,I691,I152717,I152798,);
nor I_8450 (I152807,I152798,I152744);
not I_8451 (I152825,I152798);
DFFARX1 I_8452 (I152663,I691,I152717,I152852,);
nand I_8453 (I152861,I152852,I152186);
not I_8454 (I152879,I152861);
DFFARX1 I_8455 (I152879,I691,I152717,I152906,);
not I_8456 (I152915,I152906);
nor I_8457 (I152933,I152744,I152861);
nor I_8458 (I152951,I152798,I152933);
DFFARX1 I_8459 (I152681,I691,I152717,I152978,);
DFFARX1 I_8460 (I152978,I691,I152717,I152996,);
not I_8461 (I153005,I152996);
not I_8462 (I153023,I152978);
nand I_8463 (I153041,I153023,I152825);
nand I_8464 (I153059,I152699,I152159);
and I_8465 (I153077,I153059,I152474);
DFFARX1 I_8466 (I153077,I691,I152717,I153104,);
nor I_8467 (I153113,I153104,I152744);
DFFARX1 I_8468 (I153113,I691,I152717,I153140,);
DFFARX1 I_8469 (I153104,I691,I152717,I153158,);
nor I_8470 (I153167,I152375,I152159);
not I_8471 (I153185,I153167);
nor I_8472 (I153203,I153005,I153185);
nand I_8473 (I153221,I153023,I153185);
nor I_8474 (I153239,I152744,I153167);
DFFARX1 I_8475 (I153167,I691,I152717,I153266,);
not I_8476 (I153275,I698);
DFFARX1 I_8477 (I153221,I691,I153275,I153302,);
not I_8478 (I153311,I153302);
DFFARX1 I_8479 (I153203,I691,I153275,I153338,);
not I_8480 (I153347,I153266);
nand I_8481 (I153365,I153347,I152807);
not I_8482 (I153383,I153365);
nor I_8483 (I153401,I153383,I152915);
nor I_8484 (I153419,I153311,I153401);
DFFARX1 I_8485 (I153419,I691,I153275,I153446,);
not I_8486 (I153455,I152915);
nand I_8487 (I153473,I153455,I153383);
and I_8488 (I153491,I153455,I152951);
nand I_8489 (I153509,I153491,I153140);
nor I_8490 (I153527,I153509,I153455);
and I_8491 (I153545,I153338,I153509);
not I_8492 (I153563,I153509);
nand I_8493 (I153581,I153338,I153563);
nor I_8494 (I153599,I153302,I153509);
not I_8495 (I153617,I153140);
nor I_8496 (I153635,I153617,I152951);
nand I_8497 (I153653,I153635,I153455);
nor I_8498 (I153671,I153365,I153653);
nor I_8499 (I153689,I153617,I153239);
and I_8500 (I153707,I153689,I153158);
or I_8501 (I153725,I153707,I153041);
DFFARX1 I_8502 (I153725,I691,I153275,I153752,);
nor I_8503 (I153761,I153752,I153473);
DFFARX1 I_8504 (I153761,I691,I153275,I153788,);
DFFARX1 I_8505 (I153752,I691,I153275,I153806,);
not I_8506 (I153815,I153752);
nor I_8507 (I153833,I153815,I153338);
nor I_8508 (I153851,I153635,I153833);
DFFARX1 I_8509 (I153851,I691,I153275,I153878,);
not I_8510 (I153887,I698);
DFFARX1 I_8511 (I153527,I691,I153887,I153914,);
DFFARX1 I_8512 (I153914,I691,I153887,I153932,);
not I_8513 (I153941,I153932);
not I_8514 (I153959,I153914);
DFFARX1 I_8515 (I153545,I691,I153887,I153986,);
not I_8516 (I153995,I153986);
and I_8517 (I154013,I153959,I153806);
not I_8518 (I154031,I153878);
nand I_8519 (I154049,I154031,I153806);
not I_8520 (I154067,I153788);
nor I_8521 (I154085,I154067,I153599);
nand I_8522 (I154103,I154085,I153671);
nor I_8523 (I154121,I154103,I154049);
DFFARX1 I_8524 (I154121,I691,I153887,I154148,);
not I_8525 (I154157,I154103);
not I_8526 (I154175,I153599);
nand I_8527 (I154193,I154175,I153806);
nor I_8528 (I154211,I153599,I153878);
nand I_8529 (I154229,I154013,I154211);
nand I_8530 (I154247,I153959,I153599);
nand I_8531 (I154265,I154067,I153446);
DFFARX1 I_8532 (I154265,I691,I153887,I154292,);
DFFARX1 I_8533 (I154265,I691,I153887,I154310,);
not I_8534 (I154319,I153446);
nor I_8535 (I154337,I154319,I153788);
and I_8536 (I154355,I154337,I153581);
or I_8537 (I154373,I154355,I153599);
DFFARX1 I_8538 (I154373,I691,I153887,I154400,);
nand I_8539 (I154409,I154400,I154031);
nor I_8540 (I154427,I154409,I154193);
nor I_8541 (I154445,I154400,I153995);
DFFARX1 I_8542 (I154400,I691,I153887,I154472,);
not I_8543 (I154481,I154472);
nor I_8544 (I154499,I154481,I154157);
not I_8545 (I154517,I698);
DFFARX1 I_8546 (I154247,I691,I154517,I154544,);
not I_8547 (I154553,I154544);
nand I_8548 (I154571,I154445,I154292);
and I_8549 (I154589,I154571,I154229);
DFFARX1 I_8550 (I154589,I691,I154517,I154616,);
DFFARX1 I_8551 (I154616,I691,I154517,I154634,);
DFFARX1 I_8552 (I154499,I691,I154517,I154652,);
nand I_8553 (I154661,I154652,I154310);
not I_8554 (I154679,I154661);
DFFARX1 I_8555 (I154679,I691,I154517,I154706,);
not I_8556 (I154715,I154706);
nor I_8557 (I154733,I154553,I154715);
DFFARX1 I_8558 (I154427,I691,I154517,I154760,);
nor I_8559 (I154769,I154760,I154616);
nor I_8560 (I154787,I154760,I154679);
nand I_8561 (I154805,I154148,I153941);
and I_8562 (I154823,I154805,I154445);
DFFARX1 I_8563 (I154823,I691,I154517,I154850,);
not I_8564 (I154859,I154850);
nand I_8565 (I154877,I154859,I154760);
nand I_8566 (I154895,I154859,I154661);
nor I_8567 (I154913,I154148,I153941);
and I_8568 (I154931,I154760,I154913);
nor I_8569 (I154949,I154859,I154931);
DFFARX1 I_8570 (I154949,I691,I154517,I154976,);
nor I_8571 (I154985,I154544,I154913);
DFFARX1 I_8572 (I154985,I691,I154517,I155012,);
nor I_8573 (I155021,I154850,I154913);
not I_8574 (I155039,I155021);
nand I_8575 (I155057,I155039,I154877);
not I_8576 (I155075,I698);
DFFARX1 I_8577 (I154976,I691,I155075,I155102,);
not I_8578 (I155111,I155102);
nand I_8579 (I155129,I154787,I154733);
and I_8580 (I155147,I155129,I154634);
DFFARX1 I_8581 (I155147,I691,I155075,I155174,);
not I_8582 (I155183,I155057);
DFFARX1 I_8583 (I154895,I691,I155075,I155210,);
not I_8584 (I155219,I155210);
nor I_8585 (I155237,I155219,I155111);
and I_8586 (I155255,I155237,I155057);
nor I_8587 (I155273,I155219,I155183);
nor I_8588 (I155291,I155174,I155273);
DFFARX1 I_8589 (I155012,I691,I155075,I155318,);
nor I_8590 (I155327,I155318,I155174);
not I_8591 (I155345,I155327);
not I_8592 (I155363,I155318);
nor I_8593 (I155381,I155363,I155255);
DFFARX1 I_8594 (I155381,I691,I155075,I155408,);
nand I_8595 (I155417,I155012,I154787);
and I_8596 (I155435,I155417,I154895);
DFFARX1 I_8597 (I155435,I691,I155075,I155462,);
nor I_8598 (I155471,I155462,I155318);
DFFARX1 I_8599 (I155471,I691,I155075,I155498,);
nand I_8600 (I155507,I155462,I155363);
nand I_8601 (I155525,I155345,I155507);
not I_8602 (I155543,I155462);
nor I_8603 (I155561,I155543,I155255);
DFFARX1 I_8604 (I155561,I691,I155075,I155588,);
nor I_8605 (I155597,I154769,I154787);
or I_8606 (I155615,I155318,I155597);
nor I_8607 (I155633,I155462,I155597);
or I_8608 (I155651,I155174,I155597);
DFFARX1 I_8609 (I155597,I691,I155075,I155678,);
not I_8610 (I155687,I698);
DFFARX1 I_8611 (I155588,I691,I155687,I155714,);
DFFARX1 I_8612 (I155633,I691,I155687,I155732,);
not I_8613 (I155741,I155732);
nor I_8614 (I155759,I155714,I155741);
DFFARX1 I_8615 (I155741,I691,I155687,I155786,);
nor I_8616 (I155795,I155525,I155615);
and I_8617 (I155813,I155795,I155498);
nor I_8618 (I155831,I155813,I155525);
not I_8619 (I155849,I155525);
and I_8620 (I155867,I155849,I155408);
nand I_8621 (I155885,I155867,I155651);
nor I_8622 (I155903,I155849,I155885);
DFFARX1 I_8623 (I155903,I691,I155687,I155930,);
not I_8624 (I155939,I155885);
nand I_8625 (I155957,I155741,I155939);
nand I_8626 (I155975,I155813,I155939);
DFFARX1 I_8627 (I155849,I691,I155687,I156002,);
not I_8628 (I156011,I155633);
nor I_8629 (I156029,I156011,I155408);
nor I_8630 (I156047,I156029,I155831);
DFFARX1 I_8631 (I156047,I691,I155687,I156074,);
not I_8632 (I156083,I156029);
DFFARX1 I_8633 (I156083,I691,I155687,I156110,);
not I_8634 (I156119,I156110);
nor I_8635 (I156137,I156119,I156029);
nor I_8636 (I156155,I156011,I155291);
and I_8637 (I156173,I156155,I155678);
or I_8638 (I156191,I156173,I155498);
DFFARX1 I_8639 (I156191,I691,I155687,I156218,);
not I_8640 (I156227,I156218);
nand I_8641 (I156245,I156227,I155939);
not I_8642 (I156263,I156245);
nand I_8643 (I156281,I156245,I155957);
nand I_8644 (I156299,I156227,I155813);
not I_8645 (I156317,I698);
DFFARX1 I_8646 (I156002,I691,I156317,I156344,);
not I_8647 (I156353,I156344);
nand I_8648 (I156371,I155975,I155930);
and I_8649 (I156389,I156371,I156263);
DFFARX1 I_8650 (I156389,I691,I156317,I156416,);
not I_8651 (I156425,I155930);
DFFARX1 I_8652 (I155786,I691,I156317,I156452,);
not I_8653 (I156461,I156452);
nor I_8654 (I156479,I156461,I156353);
and I_8655 (I156497,I156479,I155930);
nor I_8656 (I156515,I156461,I156425);
nor I_8657 (I156533,I156416,I156515);
DFFARX1 I_8658 (I156299,I691,I156317,I156560,);
nor I_8659 (I156569,I156560,I156416);
not I_8660 (I156587,I156569);
not I_8661 (I156605,I156560);
nor I_8662 (I156623,I156605,I156497);
DFFARX1 I_8663 (I156623,I691,I156317,I156650,);
nand I_8664 (I156659,I155759,I156281);
and I_8665 (I156677,I156659,I156074);
DFFARX1 I_8666 (I156677,I691,I156317,I156704,);
nor I_8667 (I156713,I156704,I156560);
DFFARX1 I_8668 (I156713,I691,I156317,I156740,);
nand I_8669 (I156749,I156704,I156605);
nand I_8670 (I156767,I156587,I156749);
not I_8671 (I156785,I156704);
nor I_8672 (I156803,I156785,I156497);
DFFARX1 I_8673 (I156803,I691,I156317,I156830,);
nor I_8674 (I156839,I156137,I156281);
or I_8675 (I156857,I156560,I156839);
nor I_8676 (I156875,I156704,I156839);
or I_8677 (I156893,I156416,I156839);
DFFARX1 I_8678 (I156839,I691,I156317,I156920,);
not I_8679 (I156929,I698);
DFFARX1 I_8680 (I156857,I691,I156929,I156956,);
DFFARX1 I_8681 (I156956,I691,I156929,I156974,);
not I_8682 (I156983,I156974);
not I_8683 (I157001,I156956);
DFFARX1 I_8684 (I156767,I691,I156929,I157028,);
not I_8685 (I157037,I157028);
and I_8686 (I157055,I157001,I156533);
not I_8687 (I157073,I156740);
nand I_8688 (I157091,I157073,I156533);
not I_8689 (I157109,I156875);
nor I_8690 (I157127,I157109,I156920);
nand I_8691 (I157145,I157127,I156830);
nor I_8692 (I157163,I157145,I157091);
DFFARX1 I_8693 (I157163,I691,I156929,I157190,);
not I_8694 (I157199,I157145);
not I_8695 (I157217,I156920);
nand I_8696 (I157235,I157217,I156533);
nor I_8697 (I157253,I156920,I156740);
nand I_8698 (I157271,I157055,I157253);
nand I_8699 (I157289,I157001,I156920);
nand I_8700 (I157307,I157109,I156740);
DFFARX1 I_8701 (I157307,I691,I156929,I157334,);
DFFARX1 I_8702 (I157307,I691,I156929,I157352,);
not I_8703 (I157361,I156740);
nor I_8704 (I157379,I157361,I156893);
and I_8705 (I157397,I157379,I156650);
or I_8706 (I157415,I157397,I156875);
DFFARX1 I_8707 (I157415,I691,I156929,I157442,);
nand I_8708 (I157451,I157442,I157073);
nor I_8709 (I157469,I157451,I157235);
nor I_8710 (I157487,I157442,I157037);
DFFARX1 I_8711 (I157442,I691,I156929,I157514,);
not I_8712 (I157523,I157514);
nor I_8713 (I157541,I157523,I157199);
not I_8714 (I157559,I698);
DFFARX1 I_8715 (I157352,I691,I157559,I157586,);
not I_8716 (I157595,I157586);
DFFARX1 I_8717 (I157190,I691,I157559,I157622,);
not I_8718 (I157631,I157541);
nand I_8719 (I157649,I157631,I157487);
not I_8720 (I157667,I157649);
nor I_8721 (I157685,I157667,I157190);
nor I_8722 (I157703,I157595,I157685);
DFFARX1 I_8723 (I157703,I691,I157559,I157730,);
not I_8724 (I157739,I157190);
nand I_8725 (I157757,I157739,I157667);
and I_8726 (I157775,I157739,I157487);
nand I_8727 (I157793,I157775,I156983);
nor I_8728 (I157811,I157793,I157739);
and I_8729 (I157829,I157622,I157793);
not I_8730 (I157847,I157793);
nand I_8731 (I157865,I157622,I157847);
nor I_8732 (I157883,I157586,I157793);
not I_8733 (I157901,I157271);
nor I_8734 (I157919,I157901,I157487);
nand I_8735 (I157937,I157919,I157739);
nor I_8736 (I157955,I157649,I157937);
nor I_8737 (I157973,I157901,I157289);
and I_8738 (I157991,I157973,I157334);
or I_8739 (I158009,I157991,I157469);
DFFARX1 I_8740 (I158009,I691,I157559,I158036,);
nor I_8741 (I158045,I158036,I157757);
DFFARX1 I_8742 (I158045,I691,I157559,I158072,);
DFFARX1 I_8743 (I158036,I691,I157559,I158090,);
not I_8744 (I158099,I158036);
nor I_8745 (I158117,I158099,I157622);
nor I_8746 (I158135,I157919,I158117);
DFFARX1 I_8747 (I158135,I691,I157559,I158162,);
not I_8748 (I158171,I698);
DFFARX1 I_8749 (I158072,I691,I158171,I158198,);
not I_8750 (I158207,I158198);
nand I_8751 (I158225,I157865,I157730);
and I_8752 (I158243,I158225,I158090);
DFFARX1 I_8753 (I158243,I691,I158171,I158270,);
not I_8754 (I158279,I158162);
DFFARX1 I_8755 (I157829,I691,I158171,I158306,);
not I_8756 (I158315,I158306);
nor I_8757 (I158333,I158315,I158207);
and I_8758 (I158351,I158333,I158162);
nor I_8759 (I158369,I158315,I158279);
nor I_8760 (I158387,I158270,I158369);
DFFARX1 I_8761 (I157811,I691,I158171,I158414,);
nor I_8762 (I158423,I158414,I158270);
not I_8763 (I158441,I158423);
not I_8764 (I158459,I158414);
nor I_8765 (I158477,I158459,I158351);
DFFARX1 I_8766 (I158477,I691,I158171,I158504,);
nand I_8767 (I158513,I157955,I157883);
and I_8768 (I158531,I158513,I158072);
DFFARX1 I_8769 (I158531,I691,I158171,I158558,);
nor I_8770 (I158567,I158558,I158414);
DFFARX1 I_8771 (I158567,I691,I158171,I158594,);
nand I_8772 (I158603,I158558,I158459);
nand I_8773 (I158621,I158441,I158603);
not I_8774 (I158639,I158558);
nor I_8775 (I158657,I158639,I158351);
DFFARX1 I_8776 (I158657,I691,I158171,I158684,);
nor I_8777 (I158693,I157883,I157883);
or I_8778 (I158711,I158414,I158693);
nor I_8779 (I158729,I158558,I158693);
or I_8780 (I158747,I158270,I158693);
DFFARX1 I_8781 (I158693,I691,I158171,I158774,);
not I_8782 (I158783,I698);
DFFARX1 I_8783 (I158684,I691,I158783,I158810,);
DFFARX1 I_8784 (I158729,I691,I158783,I158828,);
not I_8785 (I158837,I158828);
nor I_8786 (I158855,I158810,I158837);
DFFARX1 I_8787 (I158837,I691,I158783,I158882,);
nor I_8788 (I158891,I158621,I158711);
and I_8789 (I158909,I158891,I158594);
nor I_8790 (I158927,I158909,I158621);
not I_8791 (I158945,I158621);
and I_8792 (I158963,I158945,I158504);
nand I_8793 (I158981,I158963,I158747);
nor I_8794 (I158999,I158945,I158981);
DFFARX1 I_8795 (I158999,I691,I158783,I159026,);
not I_8796 (I159035,I158981);
nand I_8797 (I159053,I158837,I159035);
nand I_8798 (I159071,I158909,I159035);
DFFARX1 I_8799 (I158945,I691,I158783,I159098,);
not I_8800 (I159107,I158729);
nor I_8801 (I159125,I159107,I158504);
nor I_8802 (I159143,I159125,I158927);
DFFARX1 I_8803 (I159143,I691,I158783,I159170,);
not I_8804 (I159179,I159125);
DFFARX1 I_8805 (I159179,I691,I158783,I159206,);
not I_8806 (I159215,I159206);
nor I_8807 (I159233,I159215,I159125);
nor I_8808 (I159251,I159107,I158387);
and I_8809 (I159269,I159251,I158774);
or I_8810 (I159287,I159269,I158594);
DFFARX1 I_8811 (I159287,I691,I158783,I159314,);
not I_8812 (I159323,I159314);
nand I_8813 (I159341,I159323,I159035);
not I_8814 (I159359,I159341);
nand I_8815 (I159377,I159341,I159053);
nand I_8816 (I159395,I159323,I158909);
not I_8817 (I159413,I698);
DFFARX1 I_8818 (I159071,I691,I159413,I159440,);
not I_8819 (I159449,I159440);
nand I_8820 (I159467,I159395,I159098);
and I_8821 (I159485,I159467,I158855);
DFFARX1 I_8822 (I159485,I691,I159413,I159512,);
DFFARX1 I_8823 (I159170,I691,I159413,I159530,);
and I_8824 (I159539,I159530,I159233);
nor I_8825 (I159557,I159512,I159539);
DFFARX1 I_8826 (I159557,I691,I159413,I159584,);
nand I_8827 (I159593,I159530,I159233);
nand I_8828 (I159611,I159449,I159593);
not I_8829 (I159629,I159611);
DFFARX1 I_8830 (I159377,I691,I159413,I159656,);
DFFARX1 I_8831 (I159656,I691,I159413,I159674,);
nand I_8832 (I159683,I158882,I159359);
and I_8833 (I159701,I159683,I159026);
DFFARX1 I_8834 (I159701,I691,I159413,I159728,);
DFFARX1 I_8835 (I159728,I691,I159413,I159746,);
not I_8836 (I159755,I159746);
not I_8837 (I159773,I159728);
nand I_8838 (I159791,I159773,I159593);
nor I_8839 (I159809,I159026,I159359);
not I_8840 (I159827,I159809);
nor I_8841 (I159845,I159773,I159827);
nor I_8842 (I159863,I159449,I159845);
DFFARX1 I_8843 (I159863,I691,I159413,I159890,);
nor I_8844 (I159899,I159512,I159827);
nor I_8845 (I159917,I159728,I159899);
nor I_8846 (I159935,I159656,I159809);
nor I_8847 (I159953,I159512,I159809);
not I_8848 (I159971,I698);
DFFARX1 I_8849 (I159755,I691,I159971,I159998,);
and I_8850 (I160007,I159998,I159584);
DFFARX1 I_8851 (I160007,I691,I159971,I160034,);
DFFARX1 I_8852 (I159890,I691,I159971,I160052,);
not I_8853 (I160061,I159917);
not I_8854 (I160079,I159953);
nand I_8855 (I160097,I160079,I160061);
nor I_8856 (I160115,I160052,I160097);
DFFARX1 I_8857 (I160097,I691,I159971,I160142,);
not I_8858 (I160151,I160142);
not I_8859 (I160169,I159629);
nand I_8860 (I160187,I160079,I160169);
DFFARX1 I_8861 (I160187,I691,I159971,I160214,);
not I_8862 (I160223,I160214);
not I_8863 (I160241,I159953);
nand I_8864 (I160259,I160241,I159674);
and I_8865 (I160277,I160061,I160259);
nor I_8866 (I160295,I160187,I160277);
DFFARX1 I_8867 (I160295,I691,I159971,I160322,);
DFFARX1 I_8868 (I160277,I691,I159971,I160340,);
nor I_8869 (I160349,I159953,I159935);
nor I_8870 (I160367,I160187,I160349);
or I_8871 (I160385,I159953,I159935);
nor I_8872 (I160403,I159791,I159584);
DFFARX1 I_8873 (I160403,I691,I159971,I160430,);
not I_8874 (I160439,I160430);
nor I_8875 (I160457,I160439,I160223);
nand I_8876 (I160475,I160439,I160052);
not I_8877 (I160493,I159791);
nand I_8878 (I160511,I160493,I160169);
nand I_8879 (I160529,I160439,I160511);
nand I_8880 (I160547,I160529,I160475);
nand I_8881 (I160565,I160511,I160385);
not I_8882 (I160583,I698);
DFFARX1 I_8883 (I160115,I691,I160583,I160610,);
DFFARX1 I_8884 (I160034,I691,I160583,I160628,);
not I_8885 (I160637,I160628);
nor I_8886 (I160655,I160610,I160637);
DFFARX1 I_8887 (I160637,I691,I160583,I160682,);
nor I_8888 (I160691,I160367,I160565);
and I_8889 (I160709,I160691,I160322);
nor I_8890 (I160727,I160709,I160367);
not I_8891 (I160745,I160367);
and I_8892 (I160763,I160745,I160547);
nand I_8893 (I160781,I160763,I160322);
nor I_8894 (I160799,I160745,I160781);
DFFARX1 I_8895 (I160799,I691,I160583,I160826,);
not I_8896 (I160835,I160781);
nand I_8897 (I160853,I160637,I160835);
nand I_8898 (I160871,I160709,I160835);
DFFARX1 I_8899 (I160745,I691,I160583,I160898,);
not I_8900 (I160907,I160151);
nor I_8901 (I160925,I160907,I160547);
nor I_8902 (I160943,I160925,I160727);
DFFARX1 I_8903 (I160943,I691,I160583,I160970,);
not I_8904 (I160979,I160925);
DFFARX1 I_8905 (I160979,I691,I160583,I161006,);
not I_8906 (I161015,I161006);
nor I_8907 (I161033,I161015,I160925);
nor I_8908 (I161051,I160907,I160457);
and I_8909 (I161069,I161051,I160340);
or I_8910 (I161087,I161069,I160115);
DFFARX1 I_8911 (I161087,I691,I160583,I161114,);
not I_8912 (I161123,I161114);
nand I_8913 (I161141,I161123,I160835);
not I_8914 (I161159,I161141);
nand I_8915 (I161177,I161141,I160853);
nand I_8916 (I161195,I161123,I160709);
not I_8917 (I161213,I698);
DFFARX1 I_8918 (I161159,I691,I161213,I161240,);
nand I_8919 (I161249,I161240,I161195);
not I_8920 (I161267,I161249);
DFFARX1 I_8921 (I161267,I691,I161213,I161294,);
DFFARX1 I_8922 (I161177,I691,I161213,I161312,);
not I_8923 (I161321,I161312);
not I_8924 (I161339,I161033);
not I_8925 (I161357,I160871);
nand I_8926 (I161375,I161321,I161357);
nor I_8927 (I161393,I161375,I161033);
DFFARX1 I_8928 (I161393,I691,I161213,I161420,);
nor I_8929 (I161429,I160871,I161033);
nand I_8930 (I161447,I161312,I161429);
nor I_8931 (I161465,I160826,I160826);
nor I_8932 (I161483,I161375,I160826);
not I_8933 (I161501,I160826);
not I_8934 (I161519,I160970);
nand I_8935 (I161537,I161519,I160655);
nand I_8936 (I161555,I161339,I161537);
not I_8937 (I161573,I161555);
nor I_8938 (I161591,I160970,I160826);
nor I_8939 (I161609,I161573,I161591);
nor I_8940 (I161627,I160682,I160970);
and I_8941 (I161645,I161627,I161465);
nor I_8942 (I161663,I161555,I161645);
DFFARX1 I_8943 (I161663,I691,I161213,I161690,);
nor I_8944 (I161699,I161249,I161645);
DFFARX1 I_8945 (I161699,I691,I161213,I161726,);
nor I_8946 (I161735,I160682,I160898);
DFFARX1 I_8947 (I161735,I691,I161213,I161762,);
nor I_8948 (I161771,I161762,I160871);
nand I_8949 (I161789,I161771,I161339);
nand I_8950 (I161807,I161789,I161447);
nand I_8951 (I161825,I161771,I161501);
not I_8952 (I161843,I698);
DFFARX1 I_8953 (I161825,I691,I161843,I161870,);
not I_8954 (I161879,I161870);
nand I_8955 (I161897,I161807,I161294);
and I_8956 (I161915,I161897,I161420);
DFFARX1 I_8957 (I161915,I691,I161843,I161942,);
not I_8958 (I161951,I161420);
DFFARX1 I_8959 (I161483,I691,I161843,I161978,);
not I_8960 (I161987,I161978);
nor I_8961 (I162005,I161987,I161879);
and I_8962 (I162023,I162005,I161420);
nor I_8963 (I162041,I161987,I161951);
nor I_8964 (I162059,I161942,I162041);
DFFARX1 I_8965 (I161726,I691,I161843,I162086,);
nor I_8966 (I162095,I162086,I161942);
not I_8967 (I162113,I162095);
not I_8968 (I162131,I162086);
nor I_8969 (I162149,I162131,I162023);
DFFARX1 I_8970 (I162149,I691,I161843,I162176,);
nand I_8971 (I162185,I161690,I161483);
and I_8972 (I162203,I162185,I161609);
DFFARX1 I_8973 (I162203,I691,I161843,I162230,);
nor I_8974 (I162239,I162230,I162086);
DFFARX1 I_8975 (I162239,I691,I161843,I162266,);
nand I_8976 (I162275,I162230,I162131);
nand I_8977 (I162293,I162113,I162275);
not I_8978 (I162311,I162230);
nor I_8979 (I162329,I162311,I162023);
DFFARX1 I_8980 (I162329,I691,I161843,I162356,);
nor I_8981 (I162365,I161825,I161483);
or I_8982 (I162383,I162086,I162365);
nor I_8983 (I162401,I162230,I162365);
or I_8984 (I162419,I161942,I162365);
DFFARX1 I_8985 (I162365,I691,I161843,I162446,);
not I_8986 (I162455,I698);
DFFARX1 I_8987 (I162401,I691,I162455,I162482,);
DFFARX1 I_8988 (I162482,I691,I162455,I162500,);
not I_8989 (I162509,I162500);
not I_8990 (I162527,I162482);
nand I_8991 (I162545,I162446,I162059);
and I_8992 (I162563,I162545,I162401);
DFFARX1 I_8993 (I162563,I691,I162455,I162590,);
not I_8994 (I162599,I162590);
DFFARX1 I_8995 (I162293,I691,I162455,I162626,);
and I_8996 (I162635,I162626,I162419);
nand I_8997 (I162653,I162626,I162419);
nand I_8998 (I162671,I162599,I162653);
DFFARX1 I_8999 (I162266,I691,I162455,I162698,);
nor I_9000 (I162707,I162698,I162635);
DFFARX1 I_9001 (I162707,I691,I162455,I162734,);
nor I_9002 (I162743,I162698,I162590);
nand I_9003 (I162761,I162266,I162383);
and I_9004 (I162779,I162761,I162356);
DFFARX1 I_9005 (I162779,I691,I162455,I162806,);
nor I_9006 (I162815,I162806,I162698);
not I_9007 (I162833,I162806);
nor I_9008 (I162851,I162833,I162599);
nor I_9009 (I162869,I162527,I162851);
DFFARX1 I_9010 (I162869,I691,I162455,I162896,);
nor I_9011 (I162905,I162833,I162698);
nor I_9012 (I162923,I162176,I162383);
nor I_9013 (I162941,I162923,I162905);
not I_9014 (I162959,I162923);
nand I_9015 (I162977,I162653,I162959);
DFFARX1 I_9016 (I162923,I691,I162455,I163004,);
DFFARX1 I_9017 (I162923,I691,I162455,I163022,);
not I_9018 (I163031,I698);
DFFARX1 I_9019 (I162896,I691,I163031,I163058,);
not I_9020 (I163067,I163058);
nand I_9021 (I163085,I162977,I162815);
and I_9022 (I163103,I163085,I163004);
DFFARX1 I_9023 (I163103,I691,I163031,I163130,);
DFFARX1 I_9024 (I162671,I691,I163031,I163148,);
and I_9025 (I163157,I163148,I162734);
nor I_9026 (I163175,I163130,I163157);
DFFARX1 I_9027 (I163175,I691,I163031,I163202,);
nand I_9028 (I163211,I163148,I162734);
nand I_9029 (I163229,I163067,I163211);
not I_9030 (I163247,I163229);
DFFARX1 I_9031 (I162734,I691,I163031,I163274,);
DFFARX1 I_9032 (I163274,I691,I163031,I163292,);
nand I_9033 (I163301,I162509,I162941);
and I_9034 (I163319,I163301,I162743);
DFFARX1 I_9035 (I163319,I691,I163031,I163346,);
DFFARX1 I_9036 (I163346,I691,I163031,I163364,);
not I_9037 (I163373,I163364);
not I_9038 (I163391,I163346);
nand I_9039 (I163409,I163391,I163211);
nor I_9040 (I163427,I163022,I162941);
not I_9041 (I163445,I163427);
nor I_9042 (I163463,I163391,I163445);
nor I_9043 (I163481,I163067,I163463);
DFFARX1 I_9044 (I163481,I691,I163031,I163508,);
nor I_9045 (I163517,I163130,I163445);
nor I_9046 (I163535,I163346,I163517);
nor I_9047 (I163553,I163274,I163427);
nor I_9048 (I163571,I163130,I163427);
not I_9049 (I163589,I698);
DFFARX1 I_9050 (I163292,I691,I163589,I163616,);
nand I_9051 (I163625,I163616,I163571);
DFFARX1 I_9052 (I163202,I691,I163589,I163652,);
DFFARX1 I_9053 (I163652,I691,I163589,I163670,);
not I_9054 (I163679,I163670);
not I_9055 (I163697,I163508);
nor I_9056 (I163715,I163508,I163247);
not I_9057 (I163733,I163202);
nand I_9058 (I163751,I163697,I163733);
nor I_9059 (I163769,I163202,I163508);
and I_9060 (I163787,I163769,I163625);
not I_9061 (I163805,I163409);
nand I_9062 (I163823,I163805,I163553);
nor I_9063 (I163841,I163409,I163571);
not I_9064 (I163859,I163841);
nand I_9065 (I163877,I163715,I163859);
DFFARX1 I_9066 (I163841,I691,I163589,I163904,);
nor I_9067 (I163913,I163535,I163202);
nor I_9068 (I163931,I163913,I163247);
and I_9069 (I163949,I163931,I163823);
DFFARX1 I_9070 (I163949,I691,I163589,I163976,);
nor I_9071 (I163985,I163913,I163751);
or I_9072 (I164003,I163841,I163913);
nor I_9073 (I164021,I163535,I163373);
DFFARX1 I_9074 (I164021,I691,I163589,I164048,);
not I_9075 (I164057,I164048);
nand I_9076 (I164075,I164057,I163697);
nor I_9077 (I164093,I164075,I163247);
DFFARX1 I_9078 (I164093,I691,I163589,I164120,);
nor I_9079 (I164129,I164057,I163751);
nor I_9080 (I164147,I163913,I164129);
not I_9081 (I164165,I698);
DFFARX1 I_9082 (I164120,I691,I164165,I164192,);
not I_9083 (I164201,I164192);
nand I_9084 (I164219,I163787,I164003);
and I_9085 (I164237,I164219,I163985);
DFFARX1 I_9086 (I164237,I691,I164165,I164264,);
not I_9087 (I164273,I163679);
DFFARX1 I_9088 (I163877,I691,I164165,I164300,);
not I_9089 (I164309,I164300);
nor I_9090 (I164327,I164309,I164201);
and I_9091 (I164345,I164327,I163679);
nor I_9092 (I164363,I164309,I164273);
nor I_9093 (I164381,I164264,I164363);
DFFARX1 I_9094 (I163787,I691,I164165,I164408,);
nor I_9095 (I164417,I164408,I164264);
not I_9096 (I164435,I164417);
not I_9097 (I164453,I164408);
nor I_9098 (I164471,I164453,I164345);
DFFARX1 I_9099 (I164471,I691,I164165,I164498,);
nand I_9100 (I164507,I163904,I164120);
and I_9101 (I164525,I164507,I163976);
DFFARX1 I_9102 (I164525,I691,I164165,I164552,);
nor I_9103 (I164561,I164552,I164408);
DFFARX1 I_9104 (I164561,I691,I164165,I164588,);
nand I_9105 (I164597,I164552,I164453);
nand I_9106 (I164615,I164435,I164597);
not I_9107 (I164633,I164552);
nor I_9108 (I164651,I164633,I164345);
DFFARX1 I_9109 (I164651,I691,I164165,I164678,);
nor I_9110 (I164687,I164147,I164120);
or I_9111 (I164705,I164408,I164687);
nor I_9112 (I164723,I164552,I164687);
or I_9113 (I164741,I164264,I164687);
DFFARX1 I_9114 (I164687,I691,I164165,I164768,);
endmodule


