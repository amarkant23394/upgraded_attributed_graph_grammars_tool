module test_I7269(I1477,I1470,I3377,I7269);
input I1477,I1470,I3377;
output I7269;
wire I5625,I5067,I6907,I5105,I5642;
DFFARX1 I_0(I3377,I1470,I5105,,,I5625,);
DFFARX1 I_1(I5642,I1470,I5105,,,I5067,);
not I_2(I6907,I1477);
DFFARX1 I_3(I5067,I1470,I6907,,,I7269,);
not I_4(I5105,I1477);
not I_5(I5642,I5625);
endmodule


