module test_I3356(I1477,I1470,I1489,I2103,I3538,I3487,I3356);
input I1477,I1470,I1489,I2103,I3538,I3487;
output I3356;
wire I1518,I3388,I1480,I3521,I3504,I3405,I3555,I3589,I1495,I3572;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
DFFARX1 I_2(I1470,I1518,,,I1480,);
nor I_3(I3521,I3504,I1495);
and I_4(I3504,I3487,I1489);
or I_5(I3405,I1480,I1495);
DFFARX1 I_6(I3538,I1470,I3388,,,I3555,);
and I_7(I3589,I3521,I3572);
DFFARX1 I_8(I2103,I1470,I1518,,,I1495,);
DFFARX1 I_9(I3589,I1470,I3388,,,I3356,);
nand I_10(I3572,I3555,I3405);
endmodule


