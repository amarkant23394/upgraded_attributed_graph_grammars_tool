module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_6_1_l_11,IN_1_5_l_11,IN_2_5_l_11,IN_3_5_l_11,IN_6_5_l_11,blif_reset_net_0_r_6,blif_clk_net_0_r_6,ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6);
input IN_1_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_6_1_l_11,IN_1_5_l_11,IN_2_5_l_11,IN_3_5_l_11,IN_6_5_l_11,blif_reset_net_0_r_6,blif_clk_net_0_r_6;
output ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6;
wire G199_1_r_11,G214_1_r_11,ACVQN1_2_r_11,P6_2_r_11,n_429_or_0_3_r_11,G78_3_r_11,n_576_3_r_11,n_102_3_r_11,n_547_3_r_11,n_42_5_r_11,G199_5_r_11,ACVQN2_0_l_11,n_266_and_0_0_l_11,ACVQN1_0_l_11,N1_1_l_11,G199_1_l_11,G214_1_l_11,n3_1_l_11,n_42_5_l_11,N3_5_l_11,G199_5_l_11,n3_5_l_11,N1_1_r_11,n3_1_r_11,P6_internal_2_r_11,n12_3_r_11,n_431_3_r_11,n11_3_r_11,n13_3_r_11,n14_3_r_11,n15_3_r_11,n16_3_r_11,N3_5_r_11,n3_5_r_11,n1_0_r_6,ACVQN1_2_l_6,P6_2_l_6,P6_internal_2_l_6,n_429_or_0_3_l_6,n12_3_l_6,n_431_3_l_6,G78_3_l_6,n_576_3_l_6,n11_3_l_6,n_102_3_l_6,n_547_3_l_6,n13_3_l_6,n14_3_l_6,n15_3_l_6,n16_3_l_6,ACVQN1_0_r_6,P6_internal_2_r_6,n12_3_r_6,n_431_3_r_6,n11_3_r_6,n13_3_r_6,n14_3_r_6,n15_3_r_6,n16_3_r_6,N3_5_r_6,n3_5_r_6;
DFFARX1 I_0(N1_1_r_11,blif_clk_net_0_r_6,n1_0_r_6,G199_1_r_11,);
DFFARX1 I_1(ACVQN2_0_l_11,blif_clk_net_0_r_6,n1_0_r_6,G214_1_r_11,);
DFFARX1 I_2(G214_1_l_11,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_r_11,);
not I_3(P6_2_r_11,P6_internal_2_r_11);
nand I_4(n_429_or_0_3_r_11,ACVQN2_0_l_11,n12_3_r_11);
DFFARX1 I_5(n_431_3_r_11,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_11,);
nand I_6(n_576_3_r_11,G199_1_l_11,n11_3_r_11);
not I_7(n_102_3_r_11,n_42_5_l_11);
nand I_8(n_547_3_r_11,G214_1_l_11,n13_3_r_11);
nor I_9(n_42_5_r_11,G199_1_l_11,G199_5_l_11);
DFFARX1 I_10(N3_5_r_11,blif_clk_net_0_r_6,n1_0_r_6,G199_5_r_11,);
DFFARX1 I_11(IN_1_0_l_11,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_l_11,);
and I_12(n_266_and_0_0_l_11,IN_4_0_l_11,ACVQN1_0_l_11);
DFFARX1 I_13(IN_2_0_l_11,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_l_11,);
and I_14(N1_1_l_11,IN_6_1_l_11,n3_1_l_11);
DFFARX1 I_15(N1_1_l_11,blif_clk_net_0_r_6,n1_0_r_6,G199_1_l_11,);
DFFARX1 I_16(IN_3_1_l_11,blif_clk_net_0_r_6,n1_0_r_6,G214_1_l_11,);
nand I_17(n3_1_l_11,IN_1_1_l_11,IN_2_1_l_11);
nor I_18(n_42_5_l_11,IN_1_5_l_11,IN_3_5_l_11);
and I_19(N3_5_l_11,IN_6_5_l_11,n3_5_l_11);
DFFARX1 I_20(N3_5_l_11,blif_clk_net_0_r_6,n1_0_r_6,G199_5_l_11,);
nand I_21(n3_5_l_11,IN_2_5_l_11,IN_3_5_l_11);
and I_22(N1_1_r_11,G199_5_l_11,n3_1_r_11);
nand I_23(n3_1_r_11,n_266_and_0_0_l_11,G199_1_l_11);
DFFARX1 I_24(n_266_and_0_0_l_11,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_r_11,);
not I_25(n12_3_r_11,G214_1_l_11);
or I_26(n_431_3_r_11,n_266_and_0_0_l_11,n14_3_r_11);
nor I_27(n11_3_r_11,n_42_5_l_11,n12_3_r_11);
nor I_28(n13_3_r_11,n_42_5_l_11,G199_5_l_11);
and I_29(n14_3_r_11,ACVQN2_0_l_11,n15_3_r_11);
nor I_30(n15_3_r_11,n_42_5_l_11,n16_3_r_11);
not I_31(n16_3_r_11,ACVQN2_0_l_11);
and I_32(N3_5_r_11,G199_1_l_11,n3_5_r_11);
nand I_33(n3_5_r_11,ACVQN2_0_l_11,G199_5_l_11);
DFFARX1 I_34(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_r_6,);
and I_35(n_266_and_0_0_r_6,n_429_or_0_3_l_6,ACVQN1_0_r_6);
DFFARX1 I_36(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_r_6,);
not I_37(P6_2_r_6,P6_internal_2_r_6);
nand I_38(n_429_or_0_3_r_6,n_102_3_l_6,n12_3_r_6);
DFFARX1 I_39(n_431_3_r_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_6,);
nand I_40(n_576_3_r_6,P6_2_l_6,n11_3_r_6);
not I_41(n_102_3_r_6,ACVQN1_2_l_6);
nand I_42(n_547_3_r_6,n_576_3_l_6,n13_3_r_6);
nor I_43(n_42_5_r_6,ACVQN1_2_l_6,n_429_or_0_3_l_6);
DFFARX1 I_44(N3_5_r_6,blif_clk_net_0_r_6,n1_0_r_6,G199_5_r_6,);
not I_45(n1_0_r_6,blif_reset_net_0_r_6);
DFFARX1 I_46(n_576_3_r_11,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_l_6,);
not I_47(P6_2_l_6,P6_internal_2_l_6);
DFFARX1 I_48(n_429_or_0_3_r_11,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_l_6,);
nand I_49(n_429_or_0_3_l_6,n12_3_l_6,n_547_3_r_11);
not I_50(n12_3_l_6,P6_2_r_11);
or I_51(n_431_3_l_6,n14_3_l_6,G199_5_r_11);
DFFARX1 I_52(n_431_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_l_6,);
nand I_53(n_576_3_l_6,n11_3_l_6,n_42_5_r_11);
nor I_54(n11_3_l_6,n12_3_l_6,n_102_3_r_11);
not I_55(n_102_3_l_6,n_102_3_r_11);
nand I_56(n_547_3_l_6,n13_3_l_6,G199_1_r_11);
nor I_57(n13_3_l_6,G78_3_r_11,n_102_3_r_11);
and I_58(n14_3_l_6,n15_3_l_6,G214_1_r_11);
nor I_59(n15_3_l_6,n16_3_l_6,ACVQN1_2_r_11);
not I_60(n16_3_l_6,n_547_3_r_11);
DFFARX1 I_61(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_r_6,);
DFFARX1 I_62(n_576_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_r_6,);
not I_63(n12_3_r_6,P6_2_l_6);
or I_64(n_431_3_r_6,n_429_or_0_3_l_6,n14_3_r_6);
nor I_65(n11_3_r_6,ACVQN1_2_l_6,n12_3_r_6);
nor I_66(n13_3_r_6,ACVQN1_2_l_6,n_547_3_l_6);
and I_67(n14_3_r_6,ACVQN1_2_l_6,n15_3_r_6);
nor I_68(n15_3_r_6,P6_2_l_6,n16_3_r_6);
not I_69(n16_3_r_6,n_102_3_l_6);
and I_70(N3_5_r_6,n_102_3_l_6,n3_5_r_6);
nand I_71(n3_5_r_6,n_429_or_0_3_l_6,n_547_3_l_6);
endmodule


