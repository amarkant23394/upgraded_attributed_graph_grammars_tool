module test_I1620(I1423,I1215,I1455,I1620);
input I1423,I1215,I1455;
output I1620;
wire I1603,I1586,I1535;
nand I_0(I1603,I1586,I1423);
not I_1(I1620,I1603);
nor I_2(I1586,I1535,I1215);
not I_3(I1535,I1455);
endmodule


