module test_I17662(I17594,I15730,I1477,I15832,I13746,I1470,I17662);
input I17594,I15730,I1477,I15832,I13746,I1470;
output I17662;
wire I15582,I17413,I15591,I17628,I17645,I15611,I15573,I15928,I17611;
not I_0(I15582,I15928);
not I_1(I17413,I1477);
nor I_2(I15591,I15832);
and I_3(I17628,I17611,I15573);
or I_4(I17645,I17628,I15582);
not I_5(I15611,I1477);
nand I_6(I15573,I15832,I15730);
DFFARX1 I_7(I17645,I1470,I17413,,,I17662,);
DFFARX1 I_8(I13746,I1470,I15611,,,I15928,);
nor I_9(I17611,I17594,I15591);
endmodule


