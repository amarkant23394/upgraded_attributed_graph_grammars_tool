module test_I1504(I1439,I1477,I1215,I1423,I1279,I1470,I1716,I1535,I1383,I1504);
input I1439,I1477,I1215,I1423,I1279,I1470,I1716,I1535,I1383;
output I1504;
wire I1518,I1750,I1733,I1880,I1603,I1586,I1897,I1767;
not I_0(I1518,I1477);
or I_1(I1750,I1733,I1279);
and I_2(I1733,I1716,I1439);
nand I_3(I1504,I1767,I1897);
DFFARX1 I_4(I1383,I1470,I1518,,,I1880,);
nand I_5(I1603,I1586,I1423);
nor I_6(I1586,I1535,I1215);
nor I_7(I1897,I1880,I1603);
DFFARX1 I_8(I1750,I1470,I1518,,,I1767,);
endmodule


