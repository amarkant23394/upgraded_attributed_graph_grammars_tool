module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_5_r_7,n6_7,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_7,n53_7,n52_7);
nor I_37(N1508_0_r_7,n51_7,n52_7);
nand I_38(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_39(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_40(n_576_5_r_7,n31_7,n32_7);
nor I_41(n_102_5_r_7,N1372_1_r_5,n_452_7_r_5);
nand I_42(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_43(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_44(n_572_7_r_7,n54_7,n33_7);
nand I_45(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_46(n_549_7_r_7,n53_7,n36_7);
nand I_47(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_48(n_452_7_r_7,N1508_1_r_5,N1372_1_r_5);
nor I_49(n4_7_l_7,G42_7_r_5,n_569_7_r_5);
not I_50(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_51(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_52(n30_7,n53_7);
and I_53(N3_8_l_7,n50_7,n_573_7_r_5);
DFFARX1 I_54(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_55(n_431_5_r_7,n40_7,n41_7);
nor I_56(n4_7_r_7,n54_7,n49_7);
and I_57(n31_7,n_102_5_r_7,n39_7);
not I_58(n32_7,G42_7_r_5);
nor I_59(n33_7,n34_7,N1508_0_r_5);
and I_60(n34_7,n35_7,N6147_2_r_5);
not I_61(n35_7,N1508_0_r_5);
nor I_62(n36_7,n37_7,G42_7_r_5);
or I_63(n37_7,n54_7,N1372_1_r_5);
or I_64(n38_7,N1371_0_r_5,N1508_6_r_5);
nor I_65(n39_7,n_452_7_r_7,N1371_0_r_5);
nand I_66(n40_7,n46_7,n47_7);
nand I_67(n41_7,n42_7,n43_7);
nor I_68(n42_7,n44_7,n45_7);
nor I_69(n43_7,N1371_0_r_5,N1508_6_r_5);
nor I_70(n44_7,N1508_0_r_5,N1507_6_r_5);
nor I_71(n45_7,n_452_7_r_5,N1508_0_r_5);
nand I_72(n46_7,n35_7,N6147_2_r_5);
not I_73(n47_7,N1508_0_r_5);
or I_74(n48_7,n_452_7_r_7,N1371_0_r_5);
not I_75(n49_7,n_452_7_r_7);
nand I_76(n50_7,N1508_6_r_5,n_572_7_r_5);
and I_77(n51_7,n_452_7_r_7,n45_7);
not I_78(n52_7,n44_7);
endmodule


