module Benchmark_testing100(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I2128,I2138,I2148,I2158,I2168,I2178,I2188,I2198,I2208);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458;
output I2128,I2138,I2148,I2158,I2168,I2178,I2188,I2198,I2208;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I1468,I1478,I1488,I1498,I1508,I1518,I1528,I1538,I1548,I1558,I1568,I1608,I1611,I1614,I1617,I1620,I1623,I1626,I1629,I1632,I1648,I1658,I1668,I1678,I1688,I1698,I1708,I1718,I1728,I1768,I1771,I1774,I1777,I1780,I1783,I1786,I1789,I1792,I1808,I1818,I1828,I1838,I1848,I1858,I1868,I1878,I1888,I1928,I1931,I1934,I1937,I1940,I1943,I1946,I1949,I1952,I1968,I1978,I1988,I1998,I2008,I2018,I2028,I2038,I2048,I2088,I2091,I2094,I2097,I2100,I2103,I2106,I2109,I2112,I2243,I2269,I2277,I2294,I2311,I2337,I2345,I2371,I2379,I2396,I2413,I2430,I2226,I2470,I2478,I2495,I2512,I2529,I2229,I2560,I2577,I2603,I2611,I2211,I2642,I2220,I2673,I2690,I2232,I2721,I2223,I2214,I2217,I2235;
IN_INSTANCE I_0 (I1420,I1468);
IN_INSTANCE I_1 (I1444,I1478);
IN_INSTANCE I_2 (I1388,I1488);
IN_INSTANCE I_3 (I1380,I1498);
IN_INSTANCE I_4 (I1404,I1508);
IN_INSTANCE I_5 (I1412,I1518);
IN_INSTANCE I_6 (I1436,I1528);
IN_INSTANCE I_7 (I1372,I1538);
IN_INSTANCE I_8 (I1428,I1548);
IN_INSTANCE I_9 (I1396,I1558);
IN_INSTANCE I_10 (I1364,I1568);
PAT_9 I_11 (I1468,I1478,I1488,I1498,I1508,I1518,I1528,I1538,I1548,I1558,I1568,I1608,I1611,I1614,I1617,I1620,I1623,I1626,I1629,I1632,I1451,I1458);
OUT_INSTANCE I_12 (I1608,I1648);
OUT_INSTANCE I_13 (I1611,I1658);
OUT_INSTANCE I_14 (I1614,I1668);
OUT_INSTANCE I_15 (I1617,I1678);
OUT_INSTANCE I_16 (I1620,I1688);
OUT_INSTANCE I_17 (I1623,I1698);
OUT_INSTANCE I_18 (I1626,I1708);
OUT_INSTANCE I_19 (I1629,I1718);
OUT_INSTANCE I_20 (I1632,I1728);
PAT_2 I_21 (I1698,I1708,I1678,I1728,I1648,I1658,I1668,I1658,I1718,I1688,I1648,I1768,I1771,I1774,I1777,I1780,I1783,I1786,I1789,I1792,I1451,I1458);
OUT_INSTANCE I_22 (I1768,I1808);
OUT_INSTANCE I_23 (I1771,I1818);
OUT_INSTANCE I_24 (I1774,I1828);
OUT_INSTANCE I_25 (I1777,I1838);
OUT_INSTANCE I_26 (I1780,I1848);
OUT_INSTANCE I_27 (I1783,I1858);
OUT_INSTANCE I_28 (I1786,I1868);
OUT_INSTANCE I_29 (I1789,I1878);
OUT_INSTANCE I_30 (I1792,I1888);
PAT_8 I_31 (I1848,I1818,I1838,I1808,I1828,I1878,I1868,I1808,I1858,I1818,I1888,I1928,I1931,I1934,I1937,I1940,I1943,I1946,I1949,I1952,I1451,I1458);
OUT_INSTANCE I_32 (I1928,I1968);
OUT_INSTANCE I_33 (I1931,I1978);
OUT_INSTANCE I_34 (I1934,I1988);
OUT_INSTANCE I_35 (I1937,I1998);
OUT_INSTANCE I_36 (I1940,I2008);
OUT_INSTANCE I_37 (I1943,I2018);
OUT_INSTANCE I_38 (I1946,I2028);
OUT_INSTANCE I_39 (I1949,I2038);
OUT_INSTANCE I_40 (I1952,I2048);
PAT_4 I_41 (I2028,I1978,I1998,I1968,I1968,I2008,I1978,I2038,I2048,I1988,I2018,I2088,I2091,I2094,I2097,I2100,I2103,I2106,I2109,I2112,I1451,I1458);
OUT_INSTANCE I_42 (I2088,I2128);
OUT_INSTANCE I_43 (I2091,I2138);
OUT_INSTANCE I_44 (I2094,I2148);
OUT_INSTANCE I_45 (I2097,I2158);
OUT_INSTANCE I_46 (I2100,I2168);
OUT_INSTANCE I_47 (I2103,I2178);
OUT_INSTANCE I_48 (I2106,I2188);
OUT_INSTANCE I_49 (I2109,I2198);
OUT_INSTANCE I_50 (I2112,I2208);
not I_51 (I2243,I1458);
DFFARX1 I_52 (I1558,I1451,I2243,I2269,);
not I_53 (I2277,I2269);
nand I_54 (I2294,I1538,I1548);
and I_55 (I2311,I2294,I1568);
DFFARX1 I_56 (I2311,I1451,I2243,I2337,);
not I_57 (I2345,I1528);
DFFARX1 I_58 (I1518,I1451,I2243,I2371,);
not I_59 (I2379,I2371);
nor I_60 (I2396,I2379,I2277);
and I_61 (I2413,I2396,I1528);
nor I_62 (I2430,I2379,I2345);
nor I_63 (I2226,I2337,I2430);
DFFARX1 I_64 (I1508,I1451,I2243,I2470,);
nor I_65 (I2478,I2470,I2337);
not I_66 (I2495,I2478);
not I_67 (I2512,I2470);
nor I_68 (I2529,I2512,I2413);
DFFARX1 I_69 (I2529,I1451,I2243,I2229,);
nand I_70 (I2560,I1478,I1488);
and I_71 (I2577,I2560,I1498);
DFFARX1 I_72 (I2577,I1451,I2243,I2603,);
nor I_73 (I2611,I2603,I2470);
DFFARX1 I_74 (I2611,I1451,I2243,I2211,);
nand I_75 (I2642,I2603,I2512);
nand I_76 (I2220,I2495,I2642);
not I_77 (I2673,I2603);
nor I_78 (I2690,I2673,I2413);
DFFARX1 I_79 (I2690,I1451,I2243,I2232,);
nor I_80 (I2721,I1468,I1488);
or I_81 (I2223,I2470,I2721);
nor I_82 (I2214,I2603,I2721);
or I_83 (I2217,I2337,I2721);
DFFARX1 I_84 (I2721,I1451,I2243,I2235,);
endmodule


