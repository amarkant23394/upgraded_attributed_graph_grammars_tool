module test_I4612(I2173,I1477,I1470,I2311,I4612);
input I2173,I1477,I1470,I2311;
output I4612;
wire I4595,I4544,I4561,I2152,I2345,I4578,I2161;
DFFARX1 I_0(I4578,I1470,I4544,,,I4595,);
not I_1(I4544,I1477);
nand I_2(I4561,I2152,I2173);
DFFARX1 I_3(I1470,,,I2152,);
DFFARX1 I_4(I1470,,,I2345,);
and I_5(I4578,I4561,I2161);
nand I_6(I2161,I2345,I2311);
not I_7(I4612,I4595);
endmodule


