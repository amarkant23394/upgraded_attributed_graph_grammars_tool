module test_final(G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12,n_431_0_l_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_12,blif_clk_net_1_r_17,n6_17,G42_1_r_12,);
nor I_1(n_572_1_r_12,n29_12,n30_12);
nand I_2(n_573_1_r_12,n26_12,n27_12);
nor I_3(n_549_1_r_12,n33_12,n34_12);
and I_4(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_5(N3_2_r_12,blif_clk_net_1_r_17,n6_17,G199_2_r_12,);
DFFARX1 I_6(n3_12,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_12,);
not I_7(P6_5_r_12,P6_5_r_internal_12);
or I_8(n_431_0_l_12,IN_8_0_l_12,n36_12);
DFFARX1 I_9(n_431_0_l_12,blif_clk_net_1_r_17,n6_17,n41_12,);
DFFARX1 I_10(IN_2_5_l_12,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_12,);
not I_11(n22_12,ACVQN1_5_l_12);
DFFARX1 I_12(IN_1_5_l_12,blif_clk_net_1_r_17,n6_17,n42_12,);
nor I_13(n4_1_r_12,n41_12,n31_12);
nor I_14(N3_2_r_12,n22_12,n40_12);
not I_15(n3_12,n39_12);
DFFARX1 I_16(ACVQN1_5_l_12,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_12,);
and I_17(n26_12,IN_5_0_l_12,IN_7_0_l_12);
nor I_18(n27_12,n28_12,n29_12);
not I_19(n28_12,IN_11_0_l_12);
nand I_20(n29_12,n31_12,n32_12);
nand I_21(n30_12,IN_11_0_l_12,n42_12);
not I_22(n31_12,G2_0_l_12);
not I_23(n32_12,IN_10_0_l_12);
nand I_24(n33_12,n31_12,n35_12);
nand I_25(n34_12,IN_5_0_l_12,IN_7_0_l_12);
nand I_26(n35_12,n41_12,n42_12);
and I_27(n36_12,IN_2_0_l_12,n37_12);
nor I_28(n37_12,IN_4_0_l_12,n38_12);
not I_29(n38_12,G1_0_l_12);
nor I_30(n39_12,IN_5_0_l_12,n38_12);
nor I_31(n40_12,G2_0_l_12,n39_12);
DFFARX1 I_32(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_33(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_34(n_573_1_r_17,n20_17,n21_17);
nand I_35(n_549_1_r_17,n23_17,n24_17);
nand I_36(n_569_1_r_17,n21_17,n22_17);
not I_37(n_452_1_r_17,n23_17);
DFFARX1 I_38(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_39(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_40(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_41(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_42(n_431_0_l_17,n26_17,ACVQN1_5_r_12);
not I_43(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_44(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_45(n20_17,n20_internal_17);
DFFARX1 I_46(n_549_1_r_12,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_47(G42_1_r_12,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_48(n19_17,n19_internal_17);
nor I_49(n4_1_r_17,n5_17,n25_17);
not I_50(n2_17,n29_17);
DFFARX1 I_51(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_52(n17_17,n17_internal_17);
nor I_53(N1_4_r_17,n29_17,n31_17);
not I_54(n5_17,G42_1_r_12);
and I_55(n21_17,n32_17,n_572_1_r_12);
not I_56(n22_17,n25_17);
nand I_57(n23_17,n20_17,n22_17);
nand I_58(n24_17,n19_17,n22_17);
nand I_59(n25_17,n30_17,n_573_1_r_12);
and I_60(n26_17,n27_17,n_572_1_r_12);
nor I_61(n27_17,n28_17,n_42_2_r_12);
not I_62(n28_17,n_573_1_r_12);
nor I_63(n29_17,n28_17,G199_2_r_12);
and I_64(n30_17,n5_17,G199_2_r_12);
nor I_65(n31_17,n21_17,G42_1_r_12);
nor I_66(n32_17,P6_5_r_12,G42_1_r_12);
endmodule


