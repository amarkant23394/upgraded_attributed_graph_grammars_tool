module test_I1342_rst(I1301_rst,I1342_rst);
,I1342_rst);
input I1301_rst;
output I1342_rst;
wire ;
not I_0(I1342_rst,I1301_rst);
endmodule


