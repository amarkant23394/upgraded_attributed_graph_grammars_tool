module test_I5433(I3422,I1477,I3521,I1470,I3365,I3685,I3572,I5300,I5433);
input I3422,I1477,I3521,I1470,I3365,I3685,I3572,I5300;
output I5433;
wire I5416,I3388,I5351,I3362,I3350,I5334,I5122,I3589,I5317,I3356,I5105;
nand I_0(I5416,I5122,I3356);
not I_1(I3388,I1477);
DFFARX1 I_2(I5334,I1470,I5105,,,I5351,);
DFFARX1 I_3(I3422,I1470,I3388,,,I3362,);
DFFARX1 I_4(I3685,I1470,I3388,,,I3350,);
or I_5(I5334,I5317,I3362);
nand I_6(I5433,I5416,I5351);
not I_7(I5122,I3350);
and I_8(I3589,I3521,I3572);
and I_9(I5317,I5300,I3365);
DFFARX1 I_10(I3589,I1470,I3388,,,I3356,);
not I_11(I5105,I1477);
endmodule


