module test_I13925(I1477,I12024,I12041,I10026,I12106,I1470,I13925);
input I1477,I12024,I12041,I10026,I12106,I1470;
output I13925;
wire I13908,I13891,I12058,I12380,I13775,I13843,I11965,I11944,I12287,I12349,I12304,I11973,I12075,I11959;
not I_0(I13908,I13891);
DFFARX1 I_1(I11944,I1470,I13775,,,I13891,);
nand I_2(I12058,I12041,I10026);
nor I_3(I12380,I12349,I12024);
not I_4(I13775,I1477);
nor I_5(I13843,I11959,I11965);
DFFARX1 I_6(I12304,I1470,I11973,,,I11965,);
not I_7(I11944,I12075);
nand I_8(I12287,I12024);
DFFARX1 I_9(I1470,I11973,,,I12349,);
and I_10(I12304,I12106,I12287);
not I_11(I11973,I1477);
DFFARX1 I_12(I12058,I1470,I11973,,,I12075,);
nand I_13(I11959,I12058,I12380);
nor I_14(I13925,I13843,I13908);
endmodule


