module Benchmark_testing25000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2683,I2690,I28856,I28868,I28877,I28880,I28865,I28874,I28862,I28871,I28859,I53683,I53659,I53671,I53665,I53680,I53674,I53668,I53662,I53677,I71533,I71509,I71521,I71515,I71530,I71524,I71518,I71512,I71527,I81648,I81624,I81636,I81630,I81645,I81639,I81633,I81627,I81642,I111088,I111112,I111094,I111097,I111085,I111103,I111106,I111091,I111100,I111109,I148138,I148117,I148111,I148126,I148114,I148129,I148120,I148123,I148135,I148132,I198446,I198449,I198431,I198440,I198452,I198443,I198434,I198437,I198455,I206538,I206541,I206523,I206532,I206544,I206535,I206526,I206529,I206547,I250826,I250829,I250820,I250811,I250814,I250823,I250808,I250817,I255042,I255045,I255036,I255027,I255030,I255039,I255024,I255033,I257150,I257153,I257144,I257135,I257138,I257147,I257132,I257141,I323872,I323860,I323881,I323857,I323878,I323869,I323875,I323866,I323863,I327918,I327906,I327927,I327903,I327924,I327915,I327921,I327912,I327909,I354506,I354494,I354515,I354491,I354512,I354503,I354509,I354500,I354497,I361442,I361430,I361451,I361427,I361448,I361439,I361445,I361436,I361433);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2683,I2690;
output I28856,I28868,I28877,I28880,I28865,I28874,I28862,I28871,I28859,I53683,I53659,I53671,I53665,I53680,I53674,I53668,I53662,I53677,I71533,I71509,I71521,I71515,I71530,I71524,I71518,I71512,I71527,I81648,I81624,I81636,I81630,I81645,I81639,I81633,I81627,I81642,I111088,I111112,I111094,I111097,I111085,I111103,I111106,I111091,I111100,I111109,I148138,I148117,I148111,I148126,I148114,I148129,I148120,I148123,I148135,I148132,I198446,I198449,I198431,I198440,I198452,I198443,I198434,I198437,I198455,I206538,I206541,I206523,I206532,I206544,I206535,I206526,I206529,I206547,I250826,I250829,I250820,I250811,I250814,I250823,I250808,I250817,I255042,I255045,I255036,I255027,I255030,I255039,I255024,I255033,I257150,I257153,I257144,I257135,I257138,I257147,I257132,I257141,I323872,I323860,I323881,I323857,I323878,I323869,I323875,I323866,I323863,I327918,I327906,I327927,I327903,I327924,I327915,I327921,I327912,I327909,I354506,I354494,I354515,I354491,I354512,I354503,I354509,I354500,I354497,I361442,I361430,I361451,I361427,I361448,I361439,I361445,I361436,I361433;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2683,I2690,I2722,I42043,I2748,I2756,I42034,I2773,I2714,I42055,I2813,I2821,I2838,I42031,I2855,I2872,I2889,I2693,I2920,I2937,I2954,I42040,I2696,I2985,I3002,I42052,I3019,I42049,I3036,I3053,I3070,I2705,I3101,I42046,I3118,I3135,I2711,I3166,I2708,I3197,I42037,I3223,I3231,I3248,I2702,I2699,I3317,I373045,I3343,I3351,I373033,I3368,I3309,I373021,I3408,I3416,I3433,I3450,I373027,I3467,I3484,I3288,I3515,I3532,I3549,I373024,I373039,I3291,I3580,I3597,I373030,I3614,I373042,I3631,I3648,I3665,I3300,I3696,I373036,I3713,I3730,I3306,I3761,I3303,I3792,I3818,I3826,I3843,I3297,I3294,I3912,I63182,I3938,I3946,I3963,I3904,I63188,I4003,I4011,I4028,I63197,I4045,I63191,I4062,I4079,I3883,I4110,I4127,I4144,I63194,I63200,I3886,I4175,I4192,I63203,I4209,I63179,I4226,I4243,I4260,I3895,I4291,I63185,I4308,I4325,I3901,I4356,I3898,I4387,I4413,I4421,I4438,I3892,I3889,I4507,I190920,I4533,I4541,I190938,I4558,I4499,I190932,I4598,I4606,I4623,I190923,I4640,I4657,I4674,I4478,I4705,I4722,I4739,I190929,I190917,I4481,I4770,I4787,I190935,I4804,I190941,I4821,I4838,I4855,I4490,I4886,I4903,I4920,I4496,I4951,I4493,I4982,I190926,I5008,I5016,I5033,I4487,I4484,I5102,I27814,I5128,I5136,I27805,I5153,I5094,I27826,I5193,I5201,I5218,I27802,I5235,I5252,I5269,I5073,I5300,I5317,I5334,I27811,I5076,I5365,I5382,I27823,I5399,I27820,I5416,I5433,I5450,I5085,I5481,I27817,I5498,I5515,I5091,I5546,I5088,I5577,I27808,I5603,I5611,I5628,I5082,I5079,I5700,I399184,I5726,I5743,I5751,I5768,I399187,I399193,I5785,I399202,I5811,I5692,I5683,I399205,I5856,I5864,I399196,I5881,I5680,I5921,I5929,I5686,I5674,I5974,I399211,I399190,I5991,I399199,I6017,I6025,I5668,I6056,I6073,I399208,I6090,I6107,I6124,I5689,I6155,I5677,I5671,I6227,I163573,I6253,I6270,I6278,I6295,I163579,I163567,I6312,I163564,I6338,I6219,I6210,I163576,I6383,I6391,I163570,I6408,I6207,I163588,I6448,I6456,I6213,I6201,I6501,I163582,I163585,I6518,I6544,I6552,I6195,I6583,I6600,I6617,I6634,I6651,I6216,I6682,I6204,I6198,I6754,I256614,I6780,I6797,I6805,I6822,I256605,I256626,I6839,I256608,I6865,I6746,I6737,I6910,I6918,I256623,I6935,I6734,I256617,I6975,I6983,I6740,I6728,I7028,I256611,I256620,I7045,I7071,I7079,I6722,I7110,I7127,I7144,I7161,I7178,I6743,I7209,I6731,I6725,I7281,I285308,I7307,I7324,I7332,I7349,I285284,I285311,I7366,I285296,I7392,I7273,I7264,I285302,I7437,I7445,I285287,I7462,I7261,I285305,I7502,I7510,I7267,I7255,I7555,I285290,I285293,I7572,I7598,I7606,I7249,I7637,I7654,I285299,I7671,I7688,I7705,I7270,I7736,I7258,I7252,I7808,I370301,I7834,I7851,I7859,I7876,I370319,I370313,I7893,I370322,I7919,I7800,I7791,I370307,I7964,I7972,I370316,I7989,I7788,I370304,I8029,I8037,I7794,I7782,I8082,I370325,I370310,I8099,I8125,I8133,I7776,I8164,I8181,I8198,I8215,I8232,I7797,I8263,I7785,I7779,I8335,I304042,I8361,I8378,I8386,I8403,I304018,I304045,I8420,I304030,I8446,I8327,I8318,I304036,I8491,I8499,I304021,I8516,I8315,I304039,I8556,I8564,I8321,I8309,I8609,I304024,I304027,I8626,I8652,I8660,I8303,I8691,I8708,I304033,I8725,I8742,I8759,I8324,I8790,I8312,I8306,I8862,I104261,I8888,I8905,I8913,I8930,I104258,I104252,I8947,I104246,I8973,I8854,I8845,I104234,I9018,I9026,I104243,I9043,I8842,I104240,I9083,I9091,I8848,I8836,I9136,I104237,I104255,I9153,I9179,I9187,I8830,I9218,I9235,I104249,I9252,I9269,I9286,I8851,I9317,I8839,I8833,I9389,I218667,I9415,I9432,I9440,I9457,I218682,I218685,I9474,I218664,I9500,I9381,I9372,I218670,I9545,I9553,I218676,I9570,I9369,I9610,I9618,I9375,I9363,I9663,I218679,I218661,I9680,I218673,I9706,I9714,I9357,I9745,I9762,I9779,I9796,I9813,I9378,I9844,I9366,I9360,I9916,I151919,I9942,I9959,I9967,I9984,I151922,I10001,I151943,I10027,I9908,I9899,I151931,I10072,I10080,I151934,I10097,I9896,I151940,I10137,I10145,I9902,I9890,I10190,I151937,I151925,I10207,I151928,I10233,I10241,I9884,I10272,I10289,I151946,I10306,I10323,I10340,I9905,I10371,I9893,I9887,I10443,I239223,I10469,I10486,I10494,I10511,I239214,I239235,I10528,I239217,I10554,I10435,I10426,I10599,I10607,I239232,I10624,I10423,I239226,I10664,I10672,I10429,I10417,I10717,I239220,I239229,I10734,I10760,I10768,I10411,I10799,I10816,I10833,I10850,I10867,I10432,I10898,I10420,I10414,I10970,I415844,I10996,I11013,I11021,I11038,I415847,I415853,I11055,I415862,I11081,I10962,I10953,I415865,I11126,I11134,I415856,I11151,I10950,I11191,I11199,I10956,I10944,I11244,I415871,I415850,I11261,I415859,I11287,I11295,I10938,I11326,I11343,I415868,I11360,I11377,I11394,I10959,I11425,I10947,I10941,I11497,I330817,I11523,I11540,I11548,I11565,I330805,I330796,I11582,I330793,I11608,I11489,I11480,I330799,I11653,I11661,I330811,I11678,I11477,I330808,I11718,I11726,I11483,I11471,I11771,I330802,I11788,I330814,I11814,I11822,I11465,I11853,I11870,I11887,I11904,I11921,I11486,I11952,I11474,I11468,I12024,I26224,I12050,I12067,I12075,I12092,I26239,I12109,I26242,I12135,I12016,I12007,I26236,I12180,I12188,I26245,I12205,I12004,I26221,I12245,I12253,I12010,I11998,I12298,I26227,I12315,I26230,I12341,I12349,I11992,I12380,I12397,I26233,I12414,I12431,I12448,I12013,I12479,I12001,I11995,I12551,I362607,I12577,I12594,I12602,I12619,I362595,I362586,I12636,I362583,I12662,I12543,I12534,I362589,I12707,I12715,I362601,I12732,I12531,I362598,I12772,I12780,I12537,I12525,I12825,I362592,I12842,I362604,I12868,I12876,I12519,I12907,I12924,I12941,I12958,I12975,I12540,I13006,I12528,I12522,I13078,I82225,I13104,I13121,I13129,I13146,I82243,I82228,I13163,I82231,I13189,I13070,I13061,I82219,I13234,I13242,I82222,I13259,I13058,I82234,I13299,I13307,I13064,I13052,I13352,I82240,I82237,I13369,I13395,I13403,I13046,I13434,I13451,I13468,I13485,I13502,I13067,I13533,I13055,I13049,I13605,I39926,I13631,I13648,I13656,I13673,I39941,I13690,I39944,I13716,I13597,I13588,I39938,I13761,I13769,I39947,I13786,I13585,I39923,I13826,I13834,I13591,I13579,I13879,I39929,I13896,I39932,I13922,I13930,I13573,I13961,I13978,I39935,I13995,I14012,I14029,I13594,I14060,I13582,I13576,I14132,I269262,I14158,I14175,I14183,I14200,I269253,I269274,I14217,I269256,I14243,I14124,I14115,I14288,I14296,I269271,I14313,I14112,I269265,I14353,I14361,I14118,I14106,I14406,I269259,I269268,I14423,I14449,I14457,I14100,I14488,I14505,I14522,I14539,I14556,I14121,I14587,I14109,I14103,I14659,I240277,I14685,I14702,I14710,I14727,I240268,I240289,I14744,I240271,I14770,I14651,I14642,I14815,I14823,I240286,I14840,I14639,I240280,I14880,I14888,I14645,I14633,I14933,I240274,I240283,I14950,I14976,I14984,I14627,I15015,I15032,I15049,I15066,I15083,I14648,I15114,I14636,I14630,I15186,I266627,I15212,I15229,I15237,I15254,I266618,I266639,I15271,I266621,I15297,I15178,I15169,I15342,I15350,I266636,I15367,I15166,I266630,I15407,I15415,I15172,I15160,I15460,I266624,I266633,I15477,I15503,I15511,I15154,I15542,I15559,I15576,I15593,I15610,I15175,I15641,I15163,I15157,I15713,I90032,I15739,I15756,I15764,I15781,I90029,I90023,I15798,I90017,I15824,I15705,I15696,I90005,I15869,I15877,I90014,I15894,I15693,I90011,I15934,I15942,I15699,I15687,I15987,I90008,I90026,I16004,I16030,I16038,I15681,I16069,I16086,I90020,I16103,I16120,I16137,I15702,I16168,I15690,I15684,I16240,I125868,I16266,I16283,I16291,I16308,I125865,I125859,I16325,I125853,I16351,I16232,I16223,I125841,I16396,I16404,I125850,I16421,I16220,I125847,I16461,I16469,I16226,I16214,I16514,I125844,I125862,I16531,I16557,I16565,I16208,I16596,I16613,I125856,I16630,I16647,I16664,I16229,I16695,I16217,I16211,I16767,I147567,I16793,I16810,I16818,I16835,I147570,I16852,I147591,I16878,I16759,I16750,I147579,I16923,I16931,I147582,I16948,I16747,I147588,I16988,I16996,I16753,I16741,I17041,I147585,I147573,I17058,I147576,I17084,I17092,I16735,I17123,I17140,I147594,I17157,I17174,I17191,I16756,I17222,I16744,I16738,I17294,I285954,I17320,I17337,I17345,I17362,I285930,I285957,I17379,I285942,I17405,I17286,I17277,I285948,I17450,I17458,I285933,I17475,I17274,I285951,I17515,I17523,I17280,I17268,I17568,I285936,I285939,I17585,I17611,I17619,I17262,I17650,I17667,I285945,I17684,I17701,I17718,I17283,I17749,I17271,I17265,I17821,I353359,I17847,I17864,I17872,I17889,I353347,I353338,I17906,I353335,I17932,I17813,I17804,I353341,I17977,I17985,I353353,I18002,I17801,I353350,I18042,I18050,I17807,I17795,I18095,I353344,I18112,I353356,I18138,I18146,I17789,I18177,I18194,I18211,I18228,I18245,I17810,I18276,I17798,I17792,I18348,I246601,I18374,I18391,I18399,I18416,I246592,I246613,I18433,I246595,I18459,I18340,I18331,I18504,I18512,I246610,I18529,I18328,I246604,I18569,I18577,I18334,I18322,I18622,I246598,I246607,I18639,I18665,I18673,I18316,I18704,I18721,I18738,I18755,I18772,I18337,I18803,I18325,I18319,I18875,I410501,I18901,I18909,I18926,I410495,I410516,I18943,I410492,I18969,I410513,I18986,I18994,I410510,I19011,I18843,I19042,I19059,I18855,I410498,I19099,I18864,I19121,I410507,I410504,I19138,I410489,I19164,I19181,I18867,I19203,I18852,I19234,I19251,I19268,I19285,I18861,I19316,I18849,I18858,I18846,I19402,I139425,I19428,I19436,I19453,I139419,I139410,I19470,I139431,I19496,I139413,I19513,I19521,I139407,I19538,I19370,I19569,I19586,I19382,I19626,I19391,I19648,I139434,I139416,I19665,I139422,I19691,I19708,I19394,I19730,I19379,I19761,I139428,I19778,I19795,I19812,I19388,I19843,I19376,I19385,I19373,I19929,I348139,I19955,I19963,I19980,I348154,I348133,I19997,I348136,I20023,I348157,I20040,I20048,I20065,I19897,I20096,I20113,I19909,I20153,I19918,I20175,I348145,I348142,I20192,I348148,I20218,I20235,I19921,I20257,I19906,I20288,I348151,I20305,I20322,I20339,I19915,I20370,I19903,I19912,I19900,I20456,I164162,I20482,I20490,I20507,I164183,I164177,I20524,I164159,I20550,I20567,I20575,I164171,I20592,I20424,I20623,I20640,I20436,I164168,I20680,I20445,I20702,I164174,I164165,I20719,I20745,I20762,I20448,I20784,I20433,I20815,I164180,I20832,I20849,I20866,I20442,I20897,I20430,I20439,I20427,I20983,I80446,I21009,I21017,I21034,I80440,I80434,I21051,I80455,I21077,I80452,I21094,I21102,I80449,I21119,I20951,I21150,I21167,I20963,I21207,I20972,I21229,I80437,I21246,I80458,I21272,I21289,I20975,I21311,I20960,I21342,I80443,I21359,I21376,I21393,I20969,I21424,I20957,I20966,I20954,I21510,I155237,I21536,I21544,I21561,I155258,I155252,I21578,I155234,I21604,I21621,I21629,I155246,I21646,I21478,I21677,I21694,I21490,I155243,I21734,I21499,I21756,I155249,I155240,I21773,I21799,I21816,I21502,I21838,I21487,I21869,I155255,I21886,I21903,I21920,I21496,I21951,I21484,I21493,I21481,I22037,I415261,I22063,I22071,I22088,I415255,I415276,I22105,I415252,I22131,I415273,I22148,I22156,I415270,I22173,I22005,I22204,I22221,I22017,I415258,I22261,I22026,I22283,I415267,I415264,I22300,I415249,I22326,I22343,I22029,I22365,I22014,I22396,I22413,I22430,I22447,I22023,I22478,I22011,I22020,I22008,I22564,I290461,I22590,I22598,I22615,I290479,I290473,I22632,I290452,I22658,I290470,I22675,I22683,I290455,I22700,I22532,I22731,I22748,I22544,I290467,I22788,I22553,I22810,I290476,I290464,I22827,I290458,I22853,I22870,I22556,I22892,I22541,I22923,I22940,I22957,I22974,I22550,I23005,I22538,I22547,I22535,I23091,I318811,I23117,I23125,I23142,I318808,I318814,I23159,I23185,I23202,I23210,I23227,I23059,I23258,I23275,I23071,I318817,I23315,I23080,I23337,I318820,I318829,I23354,I318823,I23380,I23397,I23083,I23419,I23068,I23450,I318826,I23467,I23484,I23501,I23077,I23532,I23065,I23074,I23062,I23618,I158807,I23644,I23652,I23669,I158828,I158822,I23686,I158804,I23712,I23729,I23737,I158816,I23754,I23586,I23785,I23802,I23598,I158813,I23842,I23607,I23864,I158819,I158810,I23881,I23907,I23924,I23610,I23946,I23595,I23977,I158825,I23994,I24011,I24028,I23604,I24059,I23592,I23601,I23589,I24145,I132897,I24171,I24179,I24196,I132891,I132882,I24213,I132903,I24239,I132885,I24256,I24264,I132879,I24281,I24113,I24312,I24329,I24125,I24369,I24134,I24391,I132906,I132888,I24408,I132894,I24434,I24451,I24137,I24473,I24122,I24504,I132900,I24521,I24538,I24555,I24131,I24586,I24119,I24128,I24116,I24672,I326753,I24698,I24706,I24723,I326768,I326747,I24740,I326750,I24766,I326771,I24783,I24791,I24808,I24640,I24839,I24856,I24652,I24896,I24661,I24918,I326759,I326756,I24935,I326762,I24961,I24978,I24664,I25000,I24649,I25031,I326765,I25048,I25065,I25082,I24658,I25113,I24646,I24655,I24643,I25199,I388274,I25225,I25233,I25250,I388277,I388271,I25267,I388268,I25293,I388253,I25310,I25318,I388262,I25335,I25167,I25366,I25383,I25179,I25423,I25188,I25445,I388256,I388259,I25462,I388265,I25488,I25505,I25191,I25527,I25176,I25558,I25575,I25592,I25609,I25185,I25640,I25173,I25182,I25170,I25726,I302089,I25752,I25760,I25777,I302107,I302101,I25794,I302080,I25820,I302098,I25837,I25845,I302083,I25862,I25694,I25893,I25910,I25706,I302095,I25950,I25715,I25972,I302104,I302092,I25989,I302086,I26015,I26032,I25718,I26054,I25703,I26085,I26102,I26119,I26136,I25712,I26167,I25700,I25709,I25697,I26253,I368675,I26279,I26287,I26304,I368669,I368690,I26321,I368681,I26347,I368672,I26364,I26372,I368684,I26389,I26420,I26437,I26477,I26499,I368693,I368678,I26516,I26542,I26559,I26581,I26612,I368687,I26629,I26646,I26663,I26694,I26780,I72711,I26806,I26814,I26831,I72705,I72699,I26848,I72720,I26874,I72717,I26891,I26899,I72714,I26916,I26748,I26947,I26964,I26760,I27004,I26769,I27026,I72702,I27043,I72723,I27069,I27086,I26772,I27108,I26757,I27139,I72708,I27156,I27173,I27190,I26766,I27221,I26754,I26763,I26751,I27307,I234857,I27333,I27341,I27358,I234848,I234866,I27375,I234845,I27401,I27418,I27426,I234851,I27443,I27275,I27474,I27491,I27287,I27531,I27296,I27553,I234863,I234854,I27570,I234869,I27596,I27613,I27299,I27635,I27284,I27666,I234860,I27683,I27700,I27717,I27293,I27748,I27281,I27290,I27278,I27834,I323299,I27860,I27868,I27885,I323296,I323302,I27902,I27928,I27945,I27953,I27970,I28001,I28018,I323305,I28058,I28080,I323308,I323317,I28097,I323311,I28123,I28140,I28162,I28193,I323314,I28210,I28227,I28244,I28275,I28361,I100045,I28387,I28395,I28412,I100027,I100042,I28429,I100018,I28455,I100021,I28472,I28480,I100036,I28497,I28329,I28528,I28545,I28341,I100039,I28585,I28350,I28607,I100030,I28624,I100024,I28650,I28667,I28353,I28689,I28338,I28720,I100033,I28737,I28754,I28771,I28347,I28802,I28335,I28344,I28332,I28888,I246074,I28914,I28922,I28939,I246071,I246086,I28956,I246068,I28982,I246065,I28999,I29007,I29024,I29055,I29072,I29112,I29134,I246080,I29151,I246083,I29177,I29194,I29216,I29247,I246077,I29264,I29281,I29298,I29329,I29415,I168327,I29441,I29449,I29466,I168348,I168342,I29483,I168324,I29509,I29526,I29534,I168336,I29551,I29383,I29582,I29599,I29395,I168333,I29639,I29404,I29661,I168339,I168330,I29678,I29704,I29721,I29407,I29743,I29392,I29774,I168345,I29791,I29808,I29825,I29401,I29856,I29389,I29398,I29386,I29942,I44160,I29968,I29976,I29993,I44157,I44139,I30010,I44145,I30036,I44154,I30053,I30061,I44148,I30078,I29910,I30109,I30126,I29922,I44163,I30166,I29931,I30188,I44151,I44142,I30205,I30231,I30248,I29934,I30270,I29919,I30301,I44166,I30318,I30335,I30352,I29928,I30383,I29916,I29925,I29913,I30469,I84016,I30495,I30503,I30520,I84010,I84004,I30537,I84025,I30563,I84022,I30580,I30588,I84019,I30605,I30437,I30636,I30653,I30449,I30693,I30458,I30715,I84007,I30732,I84028,I30758,I30775,I30461,I30797,I30446,I30828,I84013,I30845,I30862,I30879,I30455,I30910,I30443,I30452,I30440,I30996,I224453,I31022,I31030,I31047,I224444,I224462,I31064,I224441,I31090,I31107,I31115,I224447,I31132,I30964,I31163,I31180,I30976,I31220,I30985,I31242,I224459,I224450,I31259,I224465,I31285,I31302,I30988,I31324,I30973,I31355,I224456,I31372,I31389,I31406,I30982,I31437,I30970,I30979,I30967,I31523,I258722,I31549,I31557,I31574,I258719,I258734,I31591,I258716,I31617,I258713,I31634,I31642,I31659,I31491,I31690,I31707,I31503,I31747,I31512,I31769,I258728,I31786,I258731,I31812,I31829,I31515,I31851,I31500,I31882,I258725,I31899,I31916,I31933,I31509,I31964,I31497,I31506,I31494,I32050,I242912,I32076,I32084,I32101,I242909,I242924,I32118,I242906,I32144,I242903,I32161,I32169,I32186,I32018,I32217,I32234,I32030,I32274,I32039,I32296,I242918,I32313,I242921,I32339,I32356,I32042,I32378,I32027,I32409,I242915,I32426,I32443,I32460,I32036,I32491,I32024,I32033,I32021,I32577,I183990,I32603,I32611,I32628,I184002,I183987,I32645,I183981,I32671,I183996,I32688,I32696,I183984,I32713,I32545,I32744,I32761,I32557,I183993,I32801,I32566,I32823,I183999,I184005,I32840,I32866,I32883,I32569,I32905,I32554,I32936,I32953,I32970,I32987,I32563,I33018,I32551,I32560,I32548,I33104,I196131,I33130,I33138,I33155,I196122,I196140,I33172,I196119,I33198,I33215,I33223,I196125,I33240,I33072,I33271,I33288,I33084,I33328,I33093,I33350,I196137,I196128,I33367,I196143,I33393,I33410,I33096,I33432,I33081,I33463,I196134,I33480,I33497,I33514,I33090,I33545,I33078,I33087,I33075,I33631,I396816,I33657,I33665,I33682,I396810,I396831,I33699,I396807,I33725,I396828,I33742,I33750,I396825,I33767,I33599,I33798,I33815,I33611,I396813,I33855,I33620,I33877,I396822,I396819,I33894,I396804,I33920,I33937,I33623,I33959,I33608,I33990,I34007,I34024,I34041,I33617,I34072,I33605,I33614,I33602,I34158,I291753,I34184,I34192,I34209,I291771,I291765,I34226,I291744,I34252,I291762,I34269,I34277,I291747,I34294,I34126,I34325,I34342,I34138,I291759,I34382,I34147,I34404,I291768,I291756,I34421,I291750,I34447,I34464,I34150,I34486,I34135,I34517,I34534,I34551,I34568,I34144,I34599,I34132,I34141,I34129,I34685,I342937,I34711,I34719,I34736,I342952,I342931,I34753,I342934,I34779,I342955,I34796,I34804,I34821,I34653,I34852,I34869,I34665,I34909,I34674,I34931,I342943,I342940,I34948,I342946,I34974,I34991,I34677,I35013,I34662,I35044,I342949,I35061,I35078,I35095,I34671,I35126,I34659,I34668,I34656,I35212,I244493,I35238,I35246,I35263,I244490,I244505,I35280,I244487,I35306,I244484,I35323,I35331,I35348,I35180,I35379,I35396,I35192,I35436,I35201,I35458,I244499,I35475,I244502,I35501,I35518,I35204,I35540,I35189,I35571,I244496,I35588,I35605,I35622,I35198,I35653,I35186,I35195,I35183,I35739,I269789,I35765,I35773,I35790,I269807,I269801,I35807,I269780,I35833,I269798,I35850,I35858,I269783,I35875,I35707,I35906,I35923,I35719,I269795,I35963,I35728,I35985,I269804,I269792,I36002,I269786,I36028,I36045,I35731,I36067,I35716,I36098,I36115,I36132,I36149,I35725,I36180,I35713,I35722,I35710,I36266,I64381,I36292,I36300,I36317,I64375,I64369,I36334,I64390,I36360,I64387,I36377,I36385,I64384,I36402,I36234,I36433,I36450,I36246,I36490,I36255,I36512,I64372,I36529,I64393,I36555,I36572,I36258,I36594,I36243,I36625,I64378,I36642,I36659,I36676,I36252,I36707,I36240,I36249,I36237,I36793,I174742,I36819,I36827,I36844,I174754,I174739,I36861,I174733,I36887,I174748,I36904,I36912,I174736,I36929,I36761,I36960,I36977,I36773,I174745,I37017,I36782,I37039,I174751,I174757,I37056,I37082,I37099,I36785,I37121,I36770,I37152,I37169,I37186,I37203,I36779,I37234,I36767,I36776,I36764,I37320,I201333,I37346,I37354,I37371,I201324,I201342,I37388,I201321,I37414,I37431,I37439,I201327,I37456,I37288,I37487,I37504,I37300,I37544,I37309,I37566,I201339,I201330,I37583,I201345,I37609,I37626,I37312,I37648,I37297,I37679,I201336,I37696,I37713,I37730,I37306,I37761,I37294,I37303,I37291,I37847,I258195,I37873,I37881,I37898,I258192,I258207,I37915,I258189,I37941,I258186,I37958,I37966,I37983,I37815,I38014,I38031,I37827,I38071,I37836,I38093,I258201,I38110,I258204,I38136,I38153,I37839,I38175,I37824,I38206,I258198,I38223,I38240,I38257,I37833,I38288,I37821,I37830,I37818,I38374,I122179,I38400,I38408,I38425,I122161,I122176,I38442,I122152,I38468,I122155,I38485,I38493,I122170,I38510,I38342,I38541,I38558,I38354,I122173,I38598,I38363,I38620,I122164,I38637,I122158,I38663,I38680,I38366,I38702,I38351,I38733,I122167,I38750,I38767,I38784,I38360,I38815,I38348,I38357,I38345,I38901,I376835,I38927,I38935,I38952,I376829,I376850,I38969,I376841,I38995,I376832,I39012,I39020,I376844,I39037,I38869,I39068,I39085,I38881,I39125,I38890,I39147,I376853,I376838,I39164,I39190,I39207,I38893,I39229,I38878,I39260,I376847,I39277,I39294,I39311,I38887,I39342,I38875,I38884,I38872,I39428,I233701,I39454,I39462,I39479,I233692,I233710,I39496,I233689,I39522,I39539,I39547,I233695,I39564,I39396,I39595,I39612,I39408,I39652,I39417,I39674,I233707,I233698,I39691,I233713,I39717,I39734,I39420,I39756,I39405,I39787,I233704,I39804,I39821,I39838,I39414,I39869,I39402,I39411,I39399,I39955,I263465,I39981,I39989,I40006,I263462,I263477,I40023,I263459,I40049,I263456,I40066,I40074,I40091,I40122,I40139,I40179,I40201,I263471,I40218,I263474,I40244,I40261,I40283,I40314,I263468,I40331,I40348,I40365,I40396,I40482,I209425,I40508,I40516,I40533,I209416,I209434,I40550,I209413,I40576,I40593,I40601,I209419,I40618,I40450,I40649,I40666,I40462,I40706,I40471,I40728,I209431,I209422,I40745,I209437,I40771,I40788,I40474,I40810,I40459,I40841,I209428,I40858,I40875,I40892,I40468,I40923,I40456,I40465,I40453,I41009,I84611,I41035,I41043,I41060,I84605,I84599,I41077,I84620,I41103,I84617,I41120,I41128,I84614,I41145,I40977,I41176,I41193,I40989,I41233,I40998,I41255,I84602,I41272,I84623,I41298,I41315,I41001,I41337,I40986,I41368,I84608,I41385,I41402,I41419,I40995,I41450,I40983,I40992,I40980,I41536,I307903,I41562,I41570,I41587,I307921,I307915,I41604,I307894,I41630,I307912,I41647,I41655,I307897,I41672,I41504,I41703,I41720,I41516,I307909,I41760,I41525,I41782,I307918,I307906,I41799,I307900,I41825,I41842,I41528,I41864,I41513,I41895,I41912,I41929,I41946,I41522,I41977,I41510,I41519,I41507,I42063,I119544,I42089,I42097,I42114,I119526,I119541,I42131,I119517,I42157,I119520,I42174,I42182,I119535,I42199,I42230,I42247,I119538,I42287,I42309,I119529,I42326,I119523,I42352,I42369,I42391,I42422,I119532,I42439,I42456,I42473,I42504,I42590,I243966,I42616,I42624,I42641,I243963,I243978,I42658,I243960,I42684,I243957,I42701,I42709,I42726,I42558,I42757,I42774,I42570,I42814,I42579,I42836,I243972,I42853,I243975,I42879,I42896,I42582,I42918,I42567,I42949,I243969,I42966,I42983,I43000,I42576,I43031,I42564,I42573,I42561,I43117,I114801,I43143,I43151,I43168,I114783,I114798,I43185,I114774,I43211,I114777,I43228,I43236,I114792,I43253,I43085,I43284,I43301,I43097,I114795,I43341,I43106,I43363,I114786,I43380,I114780,I43406,I43423,I43109,I43445,I43094,I43476,I114789,I43493,I43510,I43527,I43103,I43558,I43091,I43100,I43088,I43644,I78066,I43670,I43678,I43695,I78060,I78054,I43712,I78075,I43738,I78072,I43755,I43763,I78069,I43780,I43612,I43811,I43828,I43624,I43868,I43633,I43890,I78057,I43907,I78078,I43933,I43950,I43636,I43972,I43621,I44003,I78063,I44020,I44037,I44054,I43630,I44085,I43618,I43627,I43615,I44174,I61418,I44200,I44208,I61412,I44234,I44242,I61397,I44259,I61406,I44276,I44307,I61394,I44338,I61400,I44355,I44372,I61403,I61415,I44389,I44406,I44423,I44482,I44499,I44516,I61409,I44542,I44573,I44581,I44612,I44629,I44646,I44677,I44694,I44769,I248179,I44795,I44803,I44829,I44837,I248176,I44854,I248188,I44871,I44746,I44902,I248182,I44740,I44933,I248194,I44950,I44967,I248185,I248173,I44984,I45001,I45018,I44755,I44752,I44758,I45077,I45094,I45111,I45137,I44737,I45168,I45176,I248191,I44761,I45207,I45224,I45241,I44743,I45272,I45289,I44734,I44749,I45364,I329062,I45390,I45398,I329059,I45424,I45432,I329068,I45449,I45466,I45341,I45497,I329071,I45335,I45528,I329065,I45545,I45562,I329080,I45579,I45596,I45613,I45350,I45347,I45353,I45672,I45689,I45706,I329083,I329077,I45732,I45332,I45763,I45771,I329074,I45356,I45802,I45819,I45836,I45338,I45867,I45884,I45329,I45344,I45959,I287874,I45985,I45993,I287895,I46019,I46027,I287877,I46044,I287868,I46061,I45936,I46092,I287880,I45930,I46123,I287871,I46140,I46157,I287889,I287892,I46174,I46191,I46208,I45945,I45942,I45948,I46267,I46284,I46301,I287883,I287886,I46327,I45927,I46358,I46366,I45951,I46397,I46414,I46431,I45933,I46462,I46479,I45924,I45939,I46554,I207679,I46580,I46588,I207700,I46614,I46622,I46639,I207691,I46656,I46531,I46687,I207688,I46525,I46718,I207697,I46735,I46752,I207682,I46769,I46786,I46803,I46540,I46537,I46543,I46862,I46879,I46896,I207703,I207685,I46922,I46522,I46953,I46961,I207694,I46546,I46992,I47009,I47026,I46528,I47057,I47074,I46519,I46534,I47149,I352760,I47175,I47183,I352757,I47209,I47217,I352766,I47234,I47251,I47126,I47282,I352769,I47120,I47313,I352763,I47330,I47347,I352778,I47364,I47381,I47398,I47135,I47132,I47138,I47457,I47474,I47491,I352781,I352775,I47517,I47117,I47548,I47556,I352772,I47141,I47587,I47604,I47621,I47123,I47652,I47669,I47114,I47129,I47744,I271078,I47770,I47778,I271099,I47804,I47812,I271081,I47829,I271072,I47846,I47721,I47877,I271084,I47715,I47908,I271075,I47925,I47942,I271093,I271096,I47959,I47976,I47993,I47730,I47727,I47733,I48052,I48069,I48086,I271087,I271090,I48112,I47712,I48143,I48151,I47736,I48182,I48199,I48216,I47718,I48247,I48264,I47709,I47724,I48336,I305325,I48362,I48379,I48328,I48401,I305334,I48427,I48435,I48452,I305322,I48469,I305313,I48486,I48503,I305319,I48520,I305337,I48537,I305310,I48554,I48304,I48585,I48602,I48619,I48636,I48316,I48310,I48681,I305316,I48325,I48319,I48726,I48743,I305328,I48760,I48777,I305331,I48803,I48811,I48313,I48307,I48865,I48873,I48322,I48931,I259773,I48957,I48974,I48923,I48996,I259767,I49022,I49030,I49047,I259785,I49064,I49081,I49098,I49115,I259779,I49132,I259770,I49149,I48899,I49180,I49197,I49214,I49231,I48911,I48905,I49276,I259782,I48920,I48914,I49321,I49338,I259788,I49355,I49372,I259776,I49398,I49406,I48908,I48902,I49460,I49468,I48917,I49526,I223875,I49552,I49569,I49518,I49591,I223872,I49617,I49625,I49642,I223878,I49659,I223863,I49676,I49693,I223866,I49710,I223887,I49727,I223884,I49744,I49494,I49775,I49792,I49809,I49826,I49506,I49500,I49871,I49515,I49509,I49916,I49933,I223869,I49950,I223881,I49967,I49993,I50001,I49503,I49497,I50055,I50063,I49512,I50121,I157031,I50147,I50164,I50113,I50186,I157025,I50212,I50220,I50237,I157040,I50254,I157037,I50271,I50288,I157028,I50305,I157019,I50322,I157022,I50339,I50089,I50370,I50387,I50404,I50421,I50101,I50095,I50466,I157043,I50110,I50104,I50511,I50528,I157034,I50545,I50562,I50588,I50596,I50098,I50092,I50650,I50658,I50107,I50716,I193819,I50742,I50759,I50708,I50781,I193816,I50807,I50815,I50832,I193822,I50849,I193807,I50866,I50883,I193810,I50900,I193831,I50917,I193828,I50934,I50684,I50965,I50982,I50999,I51016,I50696,I50690,I51061,I50705,I50699,I51106,I51123,I193813,I51140,I193825,I51157,I51183,I51191,I50693,I50687,I51245,I51253,I50702,I51311,I130727,I51337,I51354,I51303,I51376,I130715,I51402,I51410,I51427,I130724,I51444,I130721,I51461,I51478,I130712,I51495,I130718,I51512,I130703,I51529,I51279,I51560,I51577,I51594,I51611,I51291,I51285,I51656,I51300,I51294,I51701,I51718,I130709,I51735,I130706,I51752,I130730,I51778,I51786,I51288,I51282,I51840,I51848,I51297,I51906,I359115,I51932,I51949,I51898,I51971,I51997,I52005,I52022,I359118,I52039,I359130,I52056,I52073,I359136,I52090,I359127,I52107,I359133,I52124,I51874,I52155,I52172,I52189,I52206,I51886,I51880,I52251,I359124,I51895,I51889,I52296,I52313,I359121,I52330,I359139,I52347,I52373,I52381,I51883,I51877,I52435,I52443,I51892,I52501,I238693,I52527,I52544,I52493,I52566,I238687,I52592,I52600,I52617,I238705,I52634,I52651,I52668,I52685,I238699,I52702,I238690,I52719,I52469,I52750,I52767,I52784,I52801,I52481,I52475,I52846,I238702,I52490,I52484,I52891,I52908,I238708,I52925,I52942,I238696,I52968,I52976,I52478,I52472,I53030,I53038,I52487,I53096,I94748,I53122,I53139,I53088,I53161,I94763,I53187,I53195,I53212,I94760,I53229,I53246,I53263,I94757,I53280,I94772,I53297,I94769,I53314,I53064,I53345,I53362,I53379,I53396,I53076,I53070,I53441,I94766,I53085,I53079,I53486,I53503,I94754,I53520,I94775,I53537,I94751,I53563,I53571,I53073,I53067,I53625,I53633,I53082,I53691,I252922,I53717,I53734,I53756,I252916,I53782,I53790,I53807,I252934,I53824,I53841,I53858,I53875,I252928,I53892,I252919,I53909,I53940,I53957,I53974,I53991,I54036,I252931,I54081,I54098,I252937,I54115,I54132,I252925,I54158,I54166,I54220,I54228,I54286,I126919,I54312,I54329,I54278,I54351,I126907,I54377,I54385,I54402,I126916,I54419,I126913,I54436,I54453,I126904,I54470,I126910,I54487,I126895,I54504,I54254,I54535,I54552,I54569,I54586,I54266,I54260,I54631,I54275,I54269,I54676,I54693,I126901,I54710,I126898,I54727,I126922,I54753,I54761,I54263,I54257,I54815,I54823,I54272,I54881,I102126,I54907,I54924,I54873,I54946,I102141,I54972,I54980,I54997,I102138,I55014,I55031,I55048,I102135,I55065,I102150,I55082,I102147,I55099,I54849,I55130,I55147,I55164,I55181,I54861,I54855,I55226,I102144,I54870,I54864,I55271,I55288,I102132,I55305,I102153,I55322,I102129,I55348,I55356,I54858,I54852,I55410,I55418,I54867,I55476,I154651,I55502,I55519,I55468,I55541,I154645,I55567,I55575,I55592,I154660,I55609,I154657,I55626,I55643,I154648,I55660,I154639,I55677,I154642,I55694,I55444,I55725,I55742,I55759,I55776,I55456,I55450,I55821,I154663,I55465,I55459,I55866,I55883,I154654,I55900,I55917,I55943,I55951,I55453,I55447,I56005,I56013,I55462,I56071,I364879,I56097,I56114,I56063,I56136,I364864,I56162,I56170,I56187,I364882,I56204,I56221,I56238,I364885,I56255,I364876,I56272,I364873,I56289,I56039,I56320,I56337,I56354,I56371,I56051,I56045,I56416,I364870,I56060,I56054,I56461,I56478,I364861,I56495,I364867,I56512,I56538,I56546,I56048,I56042,I56600,I56608,I56057,I56666,I329637,I56692,I56709,I56658,I56731,I56757,I56765,I56782,I329640,I56799,I329652,I56816,I56833,I329658,I56850,I329649,I56867,I329655,I56884,I56634,I56915,I56932,I56949,I56966,I56646,I56640,I57011,I329646,I56655,I56649,I57056,I57073,I329643,I57090,I329661,I57107,I57133,I57141,I56643,I56637,I57195,I57203,I56652,I57261,I144871,I57287,I57304,I57253,I57326,I144859,I57352,I57360,I57377,I144868,I57394,I144865,I57411,I57428,I144856,I57445,I144862,I57462,I144847,I57479,I57229,I57510,I57527,I57544,I57561,I57241,I57235,I57606,I57250,I57244,I57651,I57668,I144853,I57685,I144850,I57702,I144874,I57728,I57736,I57238,I57232,I57790,I57798,I57247,I57856,I97383,I57882,I57899,I57848,I57921,I97398,I57947,I57955,I57972,I97395,I57989,I58006,I58023,I97392,I58040,I97407,I58057,I97404,I58074,I57824,I58105,I58122,I58139,I58156,I57836,I57830,I58201,I97401,I57845,I57839,I58246,I58263,I97389,I58280,I97410,I58297,I97386,I58323,I58331,I57833,I57827,I58385,I58393,I57842,I58451,I324435,I58477,I58494,I58443,I58516,I58542,I58550,I58567,I324438,I58584,I324450,I58601,I58618,I324456,I58635,I324447,I58652,I324453,I58669,I58419,I58700,I58717,I58734,I58751,I58431,I58425,I58796,I324444,I58440,I58434,I58841,I58858,I324441,I58875,I324459,I58892,I58918,I58926,I58428,I58422,I58980,I58988,I58437,I59046,I156436,I59072,I59089,I59038,I59111,I156430,I59137,I59145,I59162,I156445,I59179,I156442,I59196,I59213,I156433,I59230,I156424,I59247,I156427,I59264,I59014,I59295,I59312,I59329,I59346,I59026,I59020,I59391,I156448,I59035,I59029,I59436,I59453,I156439,I59470,I59487,I59513,I59521,I59023,I59017,I59575,I59583,I59032,I59641,I296927,I59667,I59684,I59633,I59706,I296936,I59732,I59740,I59757,I296924,I59774,I296915,I59791,I59808,I296921,I59825,I296939,I59842,I296912,I59859,I59609,I59890,I59907,I59924,I59941,I59621,I59615,I59986,I296918,I59630,I59624,I60031,I60048,I296930,I60065,I60082,I296933,I60108,I60116,I59618,I59612,I60170,I60178,I59627,I60236,I115828,I60262,I60279,I60228,I60301,I115843,I60327,I60335,I60352,I115840,I60369,I60386,I60403,I115837,I60420,I115852,I60437,I115849,I60454,I60204,I60485,I60502,I60519,I60536,I60216,I60210,I60581,I115846,I60225,I60219,I60626,I60643,I115834,I60660,I115855,I60677,I115831,I60703,I60711,I60213,I60207,I60765,I60773,I60222,I60831,I136167,I60857,I60874,I60823,I60896,I136155,I60922,I60930,I60947,I136164,I60964,I136161,I60981,I60998,I136152,I61015,I136158,I61032,I136143,I61049,I60799,I61080,I61097,I61114,I61131,I60811,I60805,I61176,I60820,I60814,I61221,I61238,I136149,I61255,I136146,I61272,I136170,I61298,I61306,I60808,I60802,I61360,I61368,I60817,I61426,I61452,I61469,I61491,I61517,I61525,I61542,I61559,I61576,I61593,I61610,I61627,I61644,I61675,I61692,I61709,I61726,I61771,I61816,I61833,I61850,I61867,I61893,I61901,I61955,I61963,I62021,I62047,I62064,I62013,I62086,I62112,I62120,I62137,I62154,I62171,I62188,I62205,I62222,I62239,I61989,I62270,I62287,I62304,I62321,I62001,I61995,I62366,I62010,I62004,I62411,I62428,I62445,I62462,I62488,I62496,I61998,I61992,I62550,I62558,I62007,I62616,I236013,I62642,I62659,I62608,I62681,I236010,I62707,I62715,I62732,I236016,I62749,I236001,I62766,I62783,I236004,I62800,I236025,I62817,I236022,I62834,I62584,I62865,I62882,I62899,I62916,I62596,I62590,I62961,I62605,I62599,I63006,I63023,I236007,I63040,I236019,I63057,I63083,I63091,I62593,I62587,I63145,I63153,I62602,I63211,I63237,I63254,I63276,I63302,I63310,I63327,I63344,I63361,I63378,I63395,I63412,I63429,I63460,I63477,I63494,I63511,I63556,I63601,I63618,I63635,I63652,I63678,I63686,I63740,I63748,I63806,I197865,I63832,I63849,I63798,I63871,I197862,I63897,I63905,I63922,I197868,I63939,I197853,I63956,I63973,I197856,I63990,I197877,I64007,I197874,I64024,I63774,I64055,I64072,I64089,I64106,I63786,I63780,I64151,I63795,I63789,I64196,I64213,I197859,I64230,I197871,I64247,I64273,I64281,I63783,I63777,I64335,I64343,I63792,I64401,I372495,I64427,I64444,I64466,I372480,I64492,I64500,I64517,I372498,I64534,I64551,I64568,I372501,I64585,I372492,I64602,I372489,I64619,I64650,I64667,I64684,I64701,I64746,I372486,I64791,I64808,I372477,I64825,I372483,I64842,I64868,I64876,I64930,I64938,I64996,I222141,I65022,I65039,I64988,I65061,I222138,I65087,I65095,I65112,I222144,I65129,I222129,I65146,I65163,I222132,I65180,I222153,I65197,I222150,I65214,I64964,I65245,I65262,I65279,I65296,I64976,I64970,I65341,I64985,I64979,I65386,I65403,I222135,I65420,I222147,I65437,I65463,I65471,I64973,I64967,I65525,I65533,I64982,I65591,I215205,I65617,I65634,I65583,I65656,I215202,I65682,I65690,I65707,I215208,I65724,I215193,I65741,I65758,I215196,I65775,I215217,I65792,I215214,I65809,I65559,I65840,I65857,I65874,I65891,I65571,I65565,I65936,I65580,I65574,I65981,I65998,I215199,I66015,I215211,I66032,I66058,I66066,I65568,I65562,I66120,I66128,I65577,I66186,I153575,I66212,I66229,I66178,I66251,I153563,I66277,I66285,I66302,I153572,I66319,I153569,I66336,I66353,I153560,I66370,I153566,I66387,I153551,I66404,I66154,I66435,I66452,I66469,I66486,I66166,I66160,I66531,I66175,I66169,I66576,I66593,I153557,I66610,I153554,I66627,I153578,I66653,I66661,I66163,I66157,I66715,I66723,I66172,I66781,I177060,I66807,I66824,I66773,I66846,I177051,I66872,I66880,I66897,I177069,I66914,I177066,I66931,I66948,I177045,I66965,I177048,I66982,I177057,I66999,I66749,I67030,I67047,I67064,I67081,I66761,I66755,I67126,I177063,I66770,I66764,I67171,I67188,I67205,I177054,I67222,I67248,I67256,I66758,I66752,I67310,I67318,I66767,I67376,I279485,I67402,I67419,I67368,I67441,I279494,I67467,I67475,I67492,I279482,I67509,I279473,I67526,I67543,I279479,I67560,I279497,I67577,I279470,I67594,I67344,I67625,I67642,I67659,I67676,I67356,I67350,I67721,I279476,I67365,I67359,I67766,I67783,I279488,I67800,I67817,I279491,I67843,I67851,I67353,I67347,I67905,I67913,I67362,I67971,I333683,I67997,I68014,I67963,I68036,I68062,I68070,I68087,I333686,I68104,I333698,I68121,I68138,I333704,I68155,I333695,I68172,I333701,I68189,I67939,I68220,I68237,I68254,I68271,I67951,I67945,I68316,I333692,I67960,I67954,I68361,I68378,I333689,I68395,I333707,I68412,I68438,I68446,I67948,I67942,I68500,I68508,I67957,I68566,I146503,I68592,I68609,I68558,I68631,I146491,I68657,I68665,I68682,I146500,I68699,I146497,I68716,I68733,I146488,I68750,I146494,I68767,I146479,I68784,I68534,I68815,I68832,I68849,I68866,I68546,I68540,I68911,I68555,I68549,I68956,I68973,I146485,I68990,I146482,I69007,I146506,I69033,I69041,I68543,I68537,I69095,I69103,I68552,I69161,I315445,I69187,I69204,I69153,I69226,I315454,I69252,I69260,I69277,I315448,I69294,I315442,I69311,I69328,I315457,I69345,I69362,I315451,I69379,I69129,I69410,I69427,I69444,I69461,I69141,I69135,I69506,I69150,I69144,I69551,I69568,I315463,I69585,I315460,I69602,I69628,I69636,I69138,I69132,I69690,I69698,I69147,I69756,I220985,I69782,I69799,I69748,I69821,I220982,I69847,I69855,I69872,I220988,I69889,I220973,I69906,I69923,I220976,I69940,I220997,I69957,I220994,I69974,I69724,I70005,I70022,I70039,I70056,I69736,I69730,I70101,I69745,I69739,I70146,I70163,I220979,I70180,I220991,I70197,I70223,I70231,I69733,I69727,I70285,I70293,I69742,I70351,I229655,I70377,I70394,I70343,I70416,I229652,I70442,I70450,I70467,I229658,I70484,I229643,I70501,I70518,I229646,I70535,I229667,I70552,I229664,I70569,I70319,I70600,I70617,I70634,I70651,I70331,I70325,I70696,I70340,I70334,I70741,I70758,I229649,I70775,I229661,I70792,I70818,I70826,I70328,I70322,I70880,I70888,I70337,I70946,I157626,I70972,I70989,I70938,I71011,I157620,I71037,I71045,I71062,I157635,I71079,I157632,I71096,I71113,I157623,I71130,I157614,I71147,I157617,I71164,I70914,I71195,I71212,I71229,I71246,I70926,I70920,I71291,I157638,I70935,I70929,I71336,I71353,I157629,I71370,I71387,I71413,I71421,I70923,I70917,I71475,I71483,I70932,I71541,I360849,I71567,I71584,I71606,I71632,I71640,I71657,I360852,I71674,I360864,I71691,I71708,I360870,I71725,I360861,I71742,I360867,I71759,I71790,I71807,I71824,I71841,I71886,I360858,I71931,I71948,I360855,I71965,I360873,I71982,I72008,I72016,I72070,I72078,I72136,I181106,I72162,I72179,I72128,I72201,I181097,I72227,I72235,I72252,I181115,I72269,I181112,I72286,I72303,I181091,I72320,I181094,I72337,I181103,I72354,I72104,I72385,I72402,I72419,I72436,I72116,I72110,I72481,I181109,I72125,I72119,I72526,I72543,I72560,I181100,I72577,I72603,I72611,I72113,I72107,I72665,I72673,I72122,I72731,I121098,I72757,I72774,I72796,I121113,I72822,I72830,I72847,I121110,I72864,I72881,I72898,I121107,I72915,I121122,I72932,I121119,I72949,I72980,I72997,I73014,I73031,I73076,I121116,I73121,I73138,I121104,I73155,I121125,I73172,I121101,I73198,I73206,I73260,I73268,I73326,I282715,I73352,I73369,I73318,I73391,I282724,I73417,I73425,I73442,I282712,I73459,I282703,I73476,I73493,I282709,I73510,I282727,I73527,I282700,I73544,I73294,I73575,I73592,I73609,I73626,I73306,I73300,I73671,I282706,I73315,I73309,I73716,I73733,I282718,I73750,I73767,I282721,I73793,I73801,I73303,I73297,I73855,I73863,I73312,I73921,I367599,I73947,I73964,I73913,I73986,I367584,I74012,I74020,I74037,I367602,I74054,I74071,I74088,I367605,I74105,I367596,I74122,I367593,I74139,I73889,I74170,I74187,I74204,I74221,I73901,I73895,I74266,I367590,I73910,I73904,I74311,I74328,I367581,I74345,I367587,I74362,I74388,I74396,I73898,I73892,I74450,I74458,I73907,I74516,I216939,I74542,I74559,I74508,I74581,I216936,I74607,I74615,I74632,I216942,I74649,I216927,I74666,I74683,I216930,I74700,I216951,I74717,I216948,I74734,I74484,I74765,I74782,I74799,I74816,I74496,I74490,I74861,I74505,I74499,I74906,I74923,I216933,I74940,I216945,I74957,I74983,I74991,I74493,I74487,I75045,I75053,I74502,I75111,I309201,I75137,I75154,I75103,I75176,I309210,I75202,I75210,I75227,I309198,I75244,I309189,I75261,I75278,I309195,I75295,I309213,I75312,I309186,I75329,I75079,I75360,I75377,I75394,I75411,I75091,I75085,I75456,I309192,I75100,I75094,I75501,I75518,I309204,I75535,I75552,I309207,I75578,I75586,I75088,I75082,I75640,I75648,I75097,I75706,I112139,I75732,I75749,I75698,I75771,I112154,I75797,I75805,I75822,I112151,I75839,I75856,I75873,I112148,I75890,I112163,I75907,I112160,I75924,I75674,I75955,I75972,I75989,I76006,I75686,I75680,I76051,I112157,I75695,I75689,I76096,I76113,I112145,I76130,I112166,I76147,I112142,I76173,I76181,I75683,I75677,I76235,I76243,I75692,I76301,I253976,I76327,I76344,I76293,I76366,I253970,I76392,I76400,I76417,I253988,I76434,I76451,I76468,I76485,I253982,I76502,I253973,I76519,I76269,I76550,I76567,I76584,I76601,I76281,I76275,I76646,I253985,I76290,I76284,I76691,I76708,I253991,I76725,I76742,I253979,I76768,I76776,I76278,I76272,I76830,I76838,I76287,I76896,I173014,I76922,I76939,I76888,I76961,I173005,I76987,I76995,I77012,I173023,I77029,I173020,I77046,I77063,I172999,I77080,I173002,I77097,I173011,I77114,I76864,I77145,I77162,I77179,I77196,I76876,I76870,I77241,I173017,I76885,I76879,I77286,I77303,I77320,I173008,I77337,I77363,I77371,I76873,I76867,I77425,I77433,I76882,I77491,I115301,I77517,I77534,I77483,I77556,I115316,I77582,I77590,I77607,I115313,I77624,I77641,I77658,I115310,I77675,I115325,I77692,I115322,I77709,I77459,I77740,I77757,I77774,I77791,I77471,I77465,I77836,I115319,I77480,I77474,I77881,I77898,I115307,I77915,I115328,I77932,I115304,I77958,I77966,I77468,I77462,I78020,I78028,I77477,I78086,I298219,I78112,I78129,I78151,I298228,I78177,I78185,I78202,I298216,I78219,I298207,I78236,I78253,I298213,I78270,I298231,I78287,I298204,I78304,I78335,I78352,I78369,I78386,I78431,I298210,I78476,I78493,I298222,I78510,I78527,I298225,I78553,I78561,I78615,I78623,I78681,I292405,I78707,I78724,I78673,I78746,I292414,I78772,I78780,I78797,I292402,I78814,I292393,I78831,I78848,I292399,I78865,I292417,I78882,I292390,I78899,I78649,I78930,I78947,I78964,I78981,I78661,I78655,I79026,I292396,I78670,I78664,I79071,I79088,I292408,I79105,I79122,I292411,I79148,I79156,I78658,I78652,I79210,I79218,I78667,I79276,I261881,I79302,I79319,I79268,I79341,I261875,I79367,I79375,I79392,I261893,I79409,I79426,I79443,I79460,I261887,I79477,I261878,I79494,I79244,I79525,I79542,I79559,I79576,I79256,I79250,I79621,I261890,I79265,I79259,I79666,I79683,I261896,I79700,I79717,I261884,I79743,I79751,I79253,I79247,I79805,I79813,I79262,I79871,I79897,I79914,I79863,I79936,I79962,I79970,I79987,I80004,I80021,I80038,I80055,I80072,I80089,I79839,I80120,I80137,I80154,I80171,I79851,I79845,I80216,I79860,I79854,I80261,I80278,I80295,I80312,I80338,I80346,I79848,I79842,I80400,I80408,I79857,I80466,I400990,I80492,I80509,I80531,I400981,I80557,I80565,I80582,I400975,I80599,I400969,I80616,I80633,I400996,I80650,I80667,I400993,I80684,I80715,I80732,I80749,I80766,I80811,I400978,I80856,I80873,I400984,I80890,I400987,I80907,I400972,I80933,I80941,I80995,I81003,I81061,I81087,I81104,I81053,I81126,I81152,I81160,I81177,I81194,I81211,I81228,I81245,I81262,I81279,I81029,I81310,I81327,I81344,I81361,I81041,I81035,I81406,I81050,I81044,I81451,I81468,I81485,I81502,I81528,I81536,I81038,I81032,I81590,I81598,I81047,I81656,I164766,I81682,I81699,I81721,I164760,I81747,I81755,I81772,I164775,I81789,I164772,I81806,I81823,I164763,I81840,I164754,I81857,I164757,I81874,I81905,I81922,I81939,I81956,I82001,I164778,I82046,I82063,I164769,I82080,I82097,I82123,I82131,I82185,I82193,I82251,I182262,I82277,I82294,I82316,I182253,I82342,I82350,I82367,I182271,I82384,I182268,I82401,I82418,I182247,I82435,I182250,I82452,I182259,I82469,I82500,I82517,I82534,I82551,I82596,I182265,I82641,I82658,I82675,I182256,I82692,I82718,I82726,I82780,I82788,I82846,I91586,I82872,I82889,I82838,I82911,I91601,I82937,I82945,I82962,I91598,I82979,I82996,I83013,I91595,I83030,I91610,I83047,I91607,I83064,I82814,I83095,I83112,I83129,I83146,I82826,I82820,I83191,I91604,I82835,I82829,I83236,I83253,I91592,I83270,I91613,I83287,I91589,I83313,I83321,I82823,I82817,I83375,I83383,I82832,I83441,I300157,I83467,I83484,I83433,I83506,I300166,I83532,I83540,I83557,I300154,I83574,I300145,I83591,I83608,I300151,I83625,I300169,I83642,I300142,I83659,I83409,I83690,I83707,I83724,I83741,I83421,I83415,I83786,I300148,I83430,I83424,I83831,I83848,I300160,I83865,I83882,I300163,I83908,I83916,I83418,I83412,I83970,I83978,I83427,I84036,I409915,I84062,I84079,I84101,I409906,I84127,I84135,I84152,I409900,I84169,I409894,I84186,I84203,I409921,I84220,I84237,I409918,I84254,I84285,I84302,I84319,I84336,I84381,I409903,I84426,I84443,I409909,I84460,I409912,I84477,I409897,I84503,I84511,I84565,I84573,I84631,I406940,I84657,I84674,I84696,I406931,I84722,I84730,I84747,I406925,I84764,I406919,I84781,I84798,I406946,I84815,I84832,I406943,I84849,I84880,I84897,I84914,I84931,I84976,I406928,I85021,I85038,I406934,I85055,I406937,I85072,I406922,I85098,I85106,I85160,I85168,I85226,I85252,I85269,I85218,I85291,I85317,I85325,I85342,I85359,I85376,I85393,I85410,I85427,I85444,I85194,I85475,I85492,I85509,I85526,I85206,I85200,I85571,I85215,I85209,I85616,I85633,I85650,I85667,I85693,I85701,I85203,I85197,I85755,I85763,I85212,I85824,I237109,I85850,I85858,I237112,I237106,I85875,I237118,I85901,I85792,I85923,I237121,I85949,I85957,I85974,I86000,I85816,I86022,I85798,I237124,I86062,I86079,I86087,I86104,I85801,I86135,I237115,I86152,I86178,I86186,I85789,I85807,I86231,I237127,I86248,I85810,I85795,I85804,I85813,I86351,I390002,I86377,I86385,I389999,I389990,I86402,I389987,I86428,I86319,I86450,I389996,I86476,I86484,I390005,I86501,I86527,I86343,I86549,I86325,I390008,I86589,I86606,I86614,I86631,I86328,I86662,I389993,I86679,I390011,I86705,I86713,I86316,I86334,I86758,I86775,I86337,I86322,I86331,I86340,I86878,I385378,I86904,I86912,I385375,I385366,I86929,I385363,I86955,I86846,I86977,I385372,I87003,I87011,I385381,I87028,I87054,I86870,I87076,I86852,I385384,I87116,I87133,I87141,I87158,I86855,I87189,I385369,I87206,I385387,I87232,I87240,I86843,I86861,I87285,I87302,I86864,I86849,I86858,I86867,I87405,I207113,I87431,I87439,I207104,I207119,I87456,I207125,I87482,I87373,I87504,I207110,I87530,I87538,I87555,I87581,I87397,I87603,I87379,I207107,I87643,I87660,I87668,I87685,I87382,I87716,I207101,I207116,I87733,I87759,I87767,I87370,I87388,I87812,I207122,I87829,I87391,I87376,I87385,I87394,I87932,I384222,I87958,I87966,I384219,I384210,I87983,I384207,I88009,I87900,I88031,I384216,I88057,I88065,I384225,I88082,I88108,I87924,I88130,I87906,I384228,I88170,I88187,I88195,I88212,I87909,I88243,I384213,I88260,I384231,I88286,I88294,I87897,I87915,I88339,I88356,I87918,I87903,I87912,I87921,I88459,I399800,I88485,I88493,I399779,I88510,I399806,I88536,I88427,I88558,I399794,I88584,I88592,I399797,I88609,I88635,I88451,I88657,I88433,I399788,I88697,I88714,I88722,I88739,I88436,I88770,I399785,I399782,I88787,I399803,I88813,I88821,I88424,I88442,I88866,I399791,I88883,I88445,I88430,I88439,I88448,I88986,I407535,I89012,I89020,I407514,I89037,I407541,I89063,I88954,I89085,I407529,I89111,I89119,I407532,I89136,I89162,I88978,I89184,I88960,I407523,I89224,I89241,I89249,I89266,I88963,I89297,I407520,I407517,I89314,I407538,I89340,I89348,I88951,I88969,I89393,I407526,I89410,I88972,I88957,I88966,I88975,I89513,I141595,I89539,I89547,I141607,I141586,I89564,I141610,I89590,I89481,I89612,I141601,I89638,I89646,I141583,I89663,I89689,I89505,I89711,I89487,I141598,I89751,I89768,I89776,I89793,I89490,I89824,I141589,I89841,I141592,I89867,I89875,I89478,I89496,I89920,I141604,I89937,I89499,I89484,I89493,I89502,I90040,I408130,I90066,I90074,I408109,I90091,I408136,I90117,I90139,I408124,I90165,I90173,I408127,I90190,I90216,I90238,I408118,I90278,I90295,I90303,I90320,I90351,I408115,I408112,I90368,I408133,I90394,I90402,I90447,I408121,I90464,I90567,I392314,I90593,I90601,I392311,I392302,I90618,I392299,I90644,I90535,I90666,I392308,I90692,I90700,I392317,I90717,I90743,I90559,I90765,I90541,I392320,I90805,I90822,I90830,I90847,I90544,I90878,I392305,I90895,I392323,I90921,I90929,I90532,I90550,I90974,I90991,I90553,I90538,I90547,I90556,I91094,I91120,I91128,I91145,I91171,I91062,I91193,I91219,I91227,I91244,I91270,I91086,I91292,I91068,I91332,I91349,I91357,I91374,I91071,I91405,I91422,I91448,I91456,I91059,I91077,I91501,I91518,I91080,I91065,I91074,I91083,I91621,I260297,I91647,I91655,I260300,I260294,I91672,I260306,I91698,I91720,I260309,I91746,I91754,I91771,I91797,I91819,I260312,I91859,I91876,I91884,I91901,I91932,I260303,I91949,I91975,I91983,I92028,I260315,I92045,I92148,I418245,I92174,I92182,I418224,I92199,I418251,I92225,I92116,I92247,I418239,I92273,I92281,I418242,I92298,I92324,I92140,I92346,I92122,I418233,I92386,I92403,I92411,I92428,I92125,I92459,I418230,I418227,I92476,I418248,I92502,I92510,I92113,I92131,I92555,I418236,I92572,I92134,I92119,I92128,I92137,I92675,I337151,I92701,I92709,I337166,I92726,I337169,I92752,I92643,I92774,I337175,I92800,I92808,I337157,I92825,I92851,I92667,I92873,I92649,I337154,I92913,I92930,I92938,I92955,I92652,I92986,I337160,I93003,I337172,I93029,I93037,I92640,I92658,I93082,I337163,I93099,I92661,I92646,I92655,I92664,I93202,I299499,I93228,I93236,I299496,I299514,I93253,I299505,I93279,I93170,I93301,I299520,I93327,I93335,I299502,I93352,I93378,I93194,I93400,I93176,I299508,I93440,I93457,I93465,I93482,I93179,I93513,I299523,I93530,I299511,I93556,I93564,I93167,I93185,I93609,I299517,I93626,I93188,I93173,I93182,I93191,I93729,I93755,I93763,I93780,I93806,I93697,I93828,I93854,I93862,I93879,I93905,I93721,I93927,I93703,I93967,I93984,I93992,I94009,I93706,I94040,I94057,I94083,I94091,I93694,I93712,I94136,I94153,I93715,I93700,I93709,I93718,I94256,I388846,I94282,I94290,I388843,I388834,I94307,I388831,I94333,I94224,I94355,I388840,I94381,I94389,I388849,I94406,I94432,I94248,I94454,I94230,I388852,I94494,I94511,I94519,I94536,I94233,I94567,I388837,I94584,I388855,I94610,I94618,I94221,I94239,I94663,I94680,I94242,I94227,I94236,I94245,I94783,I94809,I94817,I94834,I94860,I94882,I94908,I94916,I94933,I94959,I94981,I95021,I95038,I95046,I95063,I95094,I95111,I95137,I95145,I95190,I95207,I95310,I330215,I95336,I95344,I330230,I95361,I330233,I95387,I95278,I95409,I330239,I95435,I95443,I330221,I95460,I95486,I95302,I95508,I95284,I330218,I95548,I95565,I95573,I95590,I95287,I95621,I330224,I95638,I330236,I95664,I95672,I95275,I95293,I95717,I330227,I95734,I95296,I95281,I95290,I95299,I95837,I169517,I95863,I95871,I169529,I95888,I169514,I95914,I95805,I95936,I169538,I95962,I95970,I169535,I95987,I96013,I95829,I96035,I95811,I169526,I96075,I96092,I96100,I96117,I95814,I96148,I169523,I96165,I169532,I96191,I96199,I95802,I95820,I96244,I169520,I96261,I95823,I95808,I95817,I95826,I96364,I96390,I96398,I96415,I96441,I96332,I96463,I96489,I96497,I96514,I96540,I96356,I96562,I96338,I96602,I96619,I96627,I96644,I96341,I96675,I96692,I96718,I96726,I96329,I96347,I96771,I96788,I96350,I96335,I96344,I96353,I96891,I294977,I96917,I96925,I294974,I294992,I96942,I294983,I96968,I96859,I96990,I294998,I97016,I97024,I294980,I97041,I97067,I96883,I97089,I96865,I294986,I97129,I97146,I97154,I97171,I96868,I97202,I295001,I97219,I294989,I97245,I97253,I96856,I96874,I97298,I294995,I97315,I96877,I96862,I96871,I96880,I97418,I387690,I97444,I97452,I387687,I387678,I97469,I387675,I97495,I97517,I387684,I97543,I97551,I387693,I97568,I97594,I97616,I387696,I97656,I97673,I97681,I97698,I97729,I387681,I97746,I387699,I97772,I97780,I97825,I97842,I97945,I97971,I97979,I97996,I98022,I97913,I98044,I98070,I98078,I98095,I98121,I97937,I98143,I97919,I98183,I98200,I98208,I98225,I97922,I98256,I98273,I98299,I98307,I97910,I97928,I98352,I98369,I97931,I97916,I97925,I97934,I98472,I307251,I98498,I98506,I307248,I307266,I98523,I307257,I98549,I98440,I98571,I307272,I98597,I98605,I307254,I98622,I98648,I98464,I98670,I98446,I307260,I98710,I98727,I98735,I98752,I98449,I98783,I307275,I98800,I307263,I98826,I98834,I98437,I98455,I98879,I307269,I98896,I98458,I98443,I98452,I98461,I98999,I405155,I99025,I99033,I405134,I99050,I405161,I99076,I98967,I99098,I405149,I99124,I99132,I405152,I99149,I99175,I98991,I99197,I98973,I405143,I99237,I99254,I99262,I99279,I98976,I99310,I405140,I405137,I99327,I405158,I99353,I99361,I98964,I98982,I99406,I405146,I99423,I98985,I98970,I98979,I98988,I99526,I130171,I99552,I99560,I130183,I130162,I99577,I130186,I99603,I99494,I99625,I130177,I99651,I99659,I130159,I99676,I99702,I99518,I99724,I99500,I130174,I99764,I99781,I99789,I99806,I99503,I99837,I130165,I99854,I130168,I99880,I99888,I99491,I99509,I99933,I130180,I99950,I99512,I99497,I99506,I99515,I100053,I204223,I100079,I100087,I204214,I204229,I100104,I204235,I100130,I100152,I204220,I100178,I100186,I100203,I100229,I100251,I204217,I100291,I100308,I100316,I100333,I100364,I204211,I204226,I100381,I100407,I100415,I100460,I204232,I100477,I100580,I310396,I100606,I100614,I310393,I100631,I310405,I100657,I100548,I100679,I100705,I100713,I310411,I100730,I100756,I100572,I100778,I100554,I310399,I100818,I100835,I100843,I100860,I100557,I100891,I310408,I310414,I100908,I100934,I100942,I100545,I100563,I100987,I310402,I101004,I100566,I100551,I100560,I100569,I101107,I316006,I101133,I101141,I316003,I101158,I316015,I101184,I101075,I101206,I101232,I101240,I316021,I101257,I101283,I101099,I101305,I101081,I316009,I101345,I101362,I101370,I101387,I101084,I101418,I316018,I316024,I101435,I101461,I101469,I101072,I101090,I101514,I316012,I101531,I101093,I101078,I101087,I101096,I101634,I314884,I101660,I101668,I314881,I101685,I314893,I101711,I101602,I101733,I101759,I101767,I314899,I101784,I101810,I101626,I101832,I101608,I314887,I101872,I101889,I101897,I101914,I101611,I101945,I314896,I314902,I101962,I101988,I101996,I101599,I101617,I102041,I314890,I102058,I101620,I101605,I101614,I101623,I102161,I102187,I102195,I102212,I102238,I102260,I102286,I102294,I102311,I102337,I102359,I102399,I102416,I102424,I102441,I102472,I102489,I102515,I102523,I102568,I102585,I102688,I102714,I102722,I102739,I102765,I102656,I102787,I102813,I102821,I102838,I102864,I102680,I102886,I102662,I102926,I102943,I102951,I102968,I102665,I102999,I103016,I103042,I103050,I102653,I102671,I103095,I103112,I102674,I102659,I102668,I102677,I103215,I371951,I103241,I103249,I371933,I371957,I103266,I371948,I103292,I103183,I103314,I371954,I103340,I103348,I371942,I103365,I103391,I103207,I103413,I103189,I103453,I103470,I103478,I103495,I103192,I103526,I371939,I371936,I103543,I371945,I103569,I103577,I103180,I103198,I103622,I103639,I103201,I103186,I103195,I103204,I103742,I364335,I103768,I103776,I364317,I364341,I103793,I364332,I103819,I103710,I103841,I364338,I103867,I103875,I364326,I103892,I103918,I103734,I103940,I103716,I103980,I103997,I104005,I104022,I103719,I104053,I364323,I364320,I104070,I364329,I104096,I104104,I103707,I103725,I104149,I104166,I103728,I103713,I103722,I103731,I104269,I171280,I104295,I104303,I171265,I171268,I104320,I171283,I104346,I104368,I171277,I104394,I104402,I104419,I104445,I104467,I171274,I104507,I104524,I104532,I104549,I104580,I171289,I104597,I171286,I104623,I104631,I104676,I171271,I104693,I104796,I104822,I104830,I104847,I104873,I104764,I104895,I104921,I104929,I104946,I104972,I104788,I104994,I104770,I105034,I105051,I105059,I105076,I104773,I105107,I105124,I105150,I105158,I104761,I104779,I105203,I105220,I104782,I104767,I104776,I104785,I105323,I105349,I105357,I105374,I105400,I105291,I105422,I105448,I105456,I105473,I105499,I105315,I105521,I105297,I105561,I105578,I105586,I105603,I105300,I105634,I105651,I105677,I105685,I105288,I105306,I105730,I105747,I105309,I105294,I105303,I105312,I105850,I241325,I105876,I105884,I241328,I241322,I105901,I241334,I105927,I105818,I105949,I241337,I105975,I105983,I106000,I106026,I105842,I106048,I105824,I241340,I106088,I106105,I106113,I106130,I105827,I106161,I241331,I106178,I106204,I106212,I105815,I105833,I106257,I241343,I106274,I105836,I105821,I105830,I105839,I106377,I303375,I106403,I106411,I303372,I303390,I106428,I303381,I106454,I106345,I106476,I303396,I106502,I106510,I303378,I106527,I106553,I106369,I106575,I106351,I303384,I106615,I106632,I106640,I106657,I106354,I106688,I303399,I106705,I303387,I106731,I106739,I106342,I106360,I106784,I303393,I106801,I106363,I106348,I106357,I106366,I106904,I352179,I106930,I106938,I352194,I106955,I352197,I106981,I106872,I107003,I352203,I107029,I107037,I352185,I107054,I107080,I106896,I107102,I106878,I352182,I107142,I107159,I107167,I107184,I106881,I107215,I352188,I107232,I352200,I107258,I107266,I106869,I106887,I107311,I352191,I107328,I106890,I106875,I106884,I106893,I107431,I145947,I107457,I107465,I145959,I145938,I107482,I145962,I107508,I107399,I107530,I145953,I107556,I107564,I145935,I107581,I107607,I107423,I107629,I107405,I145950,I107669,I107686,I107694,I107711,I107408,I107742,I145941,I107759,I145944,I107785,I107793,I107396,I107414,I107838,I145956,I107855,I107417,I107402,I107411,I107420,I107958,I142139,I107984,I107992,I142151,I142130,I108009,I142154,I108035,I107926,I108057,I142145,I108083,I108091,I142127,I108108,I108134,I107950,I108156,I107932,I142142,I108196,I108213,I108221,I108238,I107935,I108269,I142133,I108286,I142136,I108312,I108320,I107923,I107941,I108365,I142148,I108382,I107944,I107929,I107938,I107947,I108485,I237636,I108511,I108519,I237639,I237633,I108536,I237645,I108562,I108453,I108584,I237648,I108610,I108618,I108635,I108661,I108477,I108683,I108459,I237651,I108723,I108740,I108748,I108765,I108462,I108796,I237642,I108813,I108839,I108847,I108450,I108468,I108892,I237654,I108909,I108471,I108456,I108465,I108474,I109012,I194975,I109038,I109046,I194966,I194981,I109063,I194987,I109089,I108980,I109111,I194972,I109137,I109145,I109162,I109188,I109004,I109210,I108986,I194969,I109250,I109267,I109275,I109292,I108989,I109323,I194963,I194978,I109340,I109366,I109374,I108977,I108995,I109419,I194984,I109436,I108998,I108983,I108992,I109001,I109539,I109565,I109573,I109590,I109616,I109507,I109638,I109664,I109672,I109689,I109715,I109531,I109737,I109513,I109777,I109794,I109802,I109819,I109516,I109850,I109867,I109893,I109901,I109504,I109522,I109946,I109963,I109525,I109510,I109519,I109528,I110066,I165947,I110092,I110100,I165959,I110117,I165944,I110143,I110034,I110165,I165968,I110191,I110199,I165965,I110216,I110242,I110058,I110264,I110040,I165956,I110304,I110321,I110329,I110346,I110043,I110377,I165953,I110394,I165962,I110420,I110428,I110031,I110049,I110473,I165950,I110490,I110052,I110037,I110046,I110055,I110593,I374127,I110619,I110627,I374109,I374133,I110644,I374124,I110670,I110561,I110692,I374130,I110718,I110726,I374118,I110743,I110769,I110585,I110791,I110567,I110831,I110848,I110856,I110873,I110570,I110904,I374115,I374112,I110921,I374121,I110947,I110955,I110558,I110576,I111000,I111017,I110579,I110564,I110573,I110582,I111120,I208269,I111146,I111154,I208260,I208275,I111171,I208281,I111197,I111219,I208266,I111245,I111253,I111270,I111296,I111318,I208263,I111358,I111375,I111383,I111400,I111431,I208257,I208272,I111448,I111474,I111482,I111527,I208278,I111544,I111647,I226187,I111673,I111681,I226178,I226193,I111698,I226199,I111724,I111615,I111746,I226184,I111772,I111780,I111797,I111823,I111639,I111845,I111621,I226181,I111885,I111902,I111910,I111927,I111624,I111958,I226175,I226190,I111975,I112001,I112009,I111612,I111630,I112054,I226196,I112071,I111633,I111618,I111627,I111636,I112174,I316567,I112200,I112208,I316564,I112225,I316576,I112251,I112273,I112299,I112307,I316582,I112324,I112350,I112372,I316570,I112412,I112429,I112437,I112454,I112485,I316579,I316585,I112502,I112528,I112536,I112581,I316573,I112598,I112701,I167732,I112727,I112735,I167744,I112752,I167729,I112778,I112669,I112800,I167753,I112826,I112834,I167750,I112851,I112877,I112693,I112899,I112675,I167741,I112939,I112956,I112964,I112981,I112678,I113012,I167738,I113029,I167747,I113055,I113063,I112666,I112684,I113108,I167735,I113125,I112687,I112672,I112681,I112690,I113228,I113254,I113262,I113279,I113305,I113196,I113327,I113353,I113361,I113378,I113404,I113220,I113426,I113202,I113466,I113483,I113491,I113508,I113205,I113539,I113556,I113582,I113590,I113193,I113211,I113635,I113652,I113214,I113199,I113208,I113217,I113755,I231389,I113781,I113789,I231380,I231395,I113806,I231401,I113832,I113723,I113854,I231386,I113880,I113888,I113905,I113931,I113747,I113953,I113729,I231383,I113993,I114010,I114018,I114035,I113732,I114066,I231377,I231392,I114083,I114109,I114117,I113720,I113738,I114162,I231398,I114179,I113741,I113726,I113735,I113744,I114282,I200755,I114308,I114316,I200746,I200761,I114333,I200767,I114359,I114250,I114381,I200752,I114407,I114415,I114432,I114458,I114274,I114480,I114256,I200749,I114520,I114537,I114545,I114562,I114259,I114593,I200743,I200758,I114610,I114636,I114644,I114247,I114265,I114689,I200764,I114706,I114268,I114253,I114262,I114271,I114809,I362005,I114835,I114843,I362020,I114860,I362023,I114886,I114908,I362029,I114934,I114942,I362011,I114959,I114985,I115007,I362008,I115047,I115064,I115072,I115089,I115120,I362014,I115137,I362026,I115163,I115171,I115216,I362017,I115233,I115336,I281411,I115362,I115370,I281408,I281426,I115387,I281417,I115413,I115435,I281432,I115461,I115469,I281414,I115486,I115512,I115534,I281420,I115574,I115591,I115599,I115616,I115647,I281435,I115664,I281423,I115690,I115698,I115743,I281429,I115760,I115863,I385956,I115889,I115897,I385953,I385944,I115914,I385941,I115940,I115962,I385950,I115988,I115996,I385959,I116013,I116039,I116061,I385962,I116101,I116118,I116126,I116143,I116174,I385947,I116191,I385965,I116217,I116225,I116270,I116287,I116390,I376303,I116416,I116424,I376285,I376309,I116441,I376300,I116467,I116358,I116489,I376306,I116515,I116523,I376294,I116540,I116566,I116382,I116588,I116364,I116628,I116645,I116653,I116670,I116367,I116701,I376291,I376288,I116718,I376297,I116744,I116752,I116355,I116373,I116797,I116814,I116376,I116361,I116370,I116379,I116917,I149755,I116943,I116951,I149767,I149746,I116968,I149770,I116994,I116885,I117016,I149761,I117042,I117050,I149743,I117067,I117093,I116909,I117115,I116891,I149758,I117155,I117172,I117180,I117197,I116894,I117228,I149749,I117245,I149752,I117271,I117279,I116882,I116900,I117324,I149764,I117341,I116903,I116888,I116897,I116906,I117444,I203067,I117470,I117478,I203058,I203073,I117495,I203079,I117521,I117412,I117543,I203064,I117569,I117577,I117594,I117620,I117436,I117642,I117418,I203061,I117682,I117699,I117707,I117724,I117421,I117755,I203055,I203070,I117772,I117798,I117806,I117409,I117427,I117851,I203076,I117868,I117430,I117415,I117424,I117433,I117971,I117997,I118005,I118022,I118048,I117939,I118070,I118096,I118104,I118121,I118147,I117963,I118169,I117945,I118209,I118226,I118234,I118251,I117948,I118282,I118299,I118325,I118333,I117936,I117954,I118378,I118395,I117957,I117942,I117951,I117960,I118498,I131259,I118524,I118532,I131271,I131250,I118549,I131274,I118575,I118466,I118597,I131265,I118623,I118631,I131247,I118648,I118674,I118490,I118696,I118472,I131262,I118736,I118753,I118761,I118778,I118475,I118809,I131253,I118826,I131256,I118852,I118860,I118463,I118481,I118905,I131268,I118922,I118484,I118469,I118478,I118487,I119025,I119051,I119059,I119076,I119102,I118993,I119124,I119150,I119158,I119175,I119201,I119017,I119223,I118999,I119263,I119280,I119288,I119305,I119002,I119336,I119353,I119379,I119387,I118990,I119008,I119432,I119449,I119011,I118996,I119005,I119014,I119552,I321055,I119578,I119586,I321052,I119603,I321064,I119629,I119651,I119677,I119685,I321070,I119702,I119728,I119750,I321058,I119790,I119807,I119815,I119832,I119863,I321067,I321073,I119880,I119906,I119914,I119959,I321061,I119976,I120079,I322738,I120105,I120113,I322735,I120130,I322747,I120156,I120047,I120178,I120204,I120212,I322753,I120229,I120255,I120071,I120277,I120053,I322741,I120317,I120334,I120342,I120359,I120056,I120390,I322750,I322756,I120407,I120433,I120441,I120044,I120062,I120486,I322744,I120503,I120065,I120050,I120059,I120068,I120606,I120632,I120640,I120657,I120683,I120574,I120705,I120731,I120739,I120756,I120782,I120598,I120804,I120580,I120844,I120861,I120869,I120886,I120583,I120917,I120934,I120960,I120968,I120571,I120589,I121013,I121030,I120592,I120577,I120586,I120595,I121133,I188042,I121159,I121167,I188027,I188030,I121184,I188045,I121210,I121232,I188039,I121258,I121266,I121283,I121309,I121331,I188036,I121371,I121388,I121396,I121413,I121444,I188051,I121461,I188048,I121487,I121495,I121540,I188033,I121557,I121660,I351023,I121686,I121694,I351038,I121711,I351041,I121737,I121628,I121759,I351047,I121785,I121793,I351029,I121810,I121836,I121652,I121858,I121634,I351026,I121898,I121915,I121923,I121940,I121637,I121971,I351032,I121988,I351044,I122014,I122022,I121625,I121643,I122067,I351035,I122084,I121646,I121631,I121640,I121649,I122187,I184574,I122213,I122221,I184559,I184562,I122238,I184577,I122264,I122286,I184571,I122312,I122320,I122337,I122363,I122385,I184568,I122425,I122442,I122450,I122467,I122498,I184583,I122515,I184580,I122541,I122549,I122594,I184565,I122611,I122714,I171858,I122740,I122748,I171843,I171846,I122765,I171861,I122791,I122682,I122813,I171855,I122839,I122847,I122864,I122890,I122706,I122912,I122688,I171852,I122952,I122969,I122977,I122994,I122691,I123025,I171867,I123042,I171864,I123068,I123076,I122679,I122697,I123121,I171849,I123138,I122700,I122685,I122694,I122703,I123241,I137243,I123267,I123275,I137255,I137234,I123292,I137258,I123318,I123209,I123340,I137249,I123366,I123374,I137231,I123391,I123417,I123233,I123439,I123215,I137246,I123479,I123496,I123504,I123521,I123218,I123552,I137237,I123569,I137240,I123595,I123603,I123206,I123224,I123648,I137252,I123665,I123227,I123212,I123221,I123230,I123768,I355069,I123794,I123802,I355084,I123819,I355087,I123845,I123736,I123867,I355093,I123893,I123901,I355075,I123918,I123944,I123760,I123966,I123742,I355072,I124006,I124023,I124031,I124048,I123745,I124079,I355078,I124096,I355090,I124122,I124130,I123733,I123751,I124175,I355081,I124192,I123754,I123739,I123748,I123757,I124295,I203645,I124321,I124329,I203636,I203651,I124346,I203657,I124372,I124263,I124394,I203642,I124420,I124428,I124445,I124471,I124287,I124493,I124269,I203639,I124533,I124550,I124558,I124575,I124272,I124606,I203633,I203648,I124623,I124649,I124657,I124260,I124278,I124702,I203654,I124719,I124281,I124266,I124275,I124284,I124822,I205379,I124848,I124856,I205370,I205385,I124873,I205391,I124899,I124790,I124921,I205376,I124947,I124955,I124972,I124998,I124814,I125020,I124796,I205373,I125060,I125077,I125085,I125102,I124799,I125133,I205367,I205382,I125150,I125176,I125184,I124787,I124805,I125229,I205388,I125246,I124808,I124793,I124802,I124811,I125349,I177638,I125375,I125383,I177623,I177626,I125400,I177641,I125426,I125317,I125448,I177635,I125474,I125482,I125499,I125525,I125341,I125547,I125323,I177632,I125587,I125604,I125612,I125629,I125326,I125660,I177647,I125677,I177644,I125703,I125711,I125314,I125332,I125756,I177629,I125773,I125335,I125320,I125329,I125338,I125876,I125902,I125910,I125927,I125953,I125975,I126001,I126009,I126026,I126052,I126074,I126114,I126131,I126139,I126156,I126187,I126204,I126230,I126238,I126283,I126300,I126403,I126429,I126437,I126454,I126480,I126371,I126502,I126528,I126536,I126553,I126579,I126395,I126601,I126377,I126641,I126658,I126666,I126683,I126380,I126714,I126731,I126757,I126765,I126368,I126386,I126810,I126827,I126389,I126374,I126383,I126392,I126930,I170690,I126956,I126973,I126995,I127012,I170687,I170708,I127029,I170711,I127055,I127063,I170696,I127089,I127097,I170699,I127114,I170702,I127154,I127162,I127207,I170693,I127224,I170705,I127250,I127272,I127289,I127306,I127337,I127354,I127385,I127474,I127500,I127517,I127466,I127539,I127556,I127573,I127599,I127607,I127633,I127641,I127658,I127445,I127698,I127706,I127439,I127454,I127751,I127768,I127794,I127442,I127816,I127833,I127850,I127457,I127881,I127898,I127448,I127929,I127451,I127463,I127460,I128018,I128044,I128061,I128010,I128083,I128100,I128117,I128143,I128151,I128177,I128185,I128202,I127989,I128242,I128250,I127983,I127998,I128295,I128312,I128338,I127986,I128360,I128377,I128394,I128001,I128425,I128442,I127992,I128473,I127995,I128007,I128004,I128562,I263995,I128588,I128605,I128554,I128627,I128644,I263989,I263986,I128661,I264001,I128687,I128695,I128721,I128729,I263983,I128746,I128533,I128786,I128794,I128527,I128542,I128839,I263998,I263992,I128856,I128882,I128530,I128904,I128921,I128938,I128545,I128969,I128986,I264004,I128536,I129017,I128539,I128551,I128548,I129106,I402186,I129132,I129149,I129098,I129171,I129188,I402162,I402183,I129205,I402180,I129231,I129239,I402159,I129265,I129273,I402171,I129290,I129077,I402174,I129330,I129338,I129071,I129086,I129383,I402177,I402165,I129400,I402168,I129426,I129074,I129448,I129465,I129482,I129089,I129513,I129530,I129080,I129561,I129083,I129095,I129092,I129650,I129676,I129693,I129642,I129715,I129732,I129749,I129775,I129783,I129809,I129817,I129834,I129621,I129874,I129882,I129615,I129630,I129927,I129944,I129970,I129618,I129992,I130009,I130026,I129633,I130057,I130074,I129624,I130105,I129627,I129639,I129636,I130194,I130220,I130237,I130259,I130276,I130293,I130319,I130327,I130353,I130361,I130378,I130418,I130426,I130471,I130488,I130514,I130536,I130553,I130570,I130601,I130618,I130649,I130738,I199012,I130764,I130781,I130803,I130820,I199033,I199024,I130837,I130863,I130871,I199018,I130897,I130905,I199015,I130922,I199009,I130962,I130970,I131015,I199021,I131032,I199030,I131058,I131080,I131097,I131114,I131145,I131162,I199027,I131193,I131282,I131308,I131325,I131347,I131364,I131381,I131407,I131415,I131441,I131449,I131466,I131506,I131514,I131559,I131576,I131602,I131624,I131641,I131658,I131689,I131706,I131737,I131826,I332530,I131852,I131869,I131818,I131891,I131908,I332542,I131925,I332533,I131951,I131959,I332551,I131985,I131993,I332527,I132010,I131797,I332545,I132050,I132058,I131791,I131806,I132103,I332539,I332536,I132120,I332548,I132146,I131794,I132168,I132185,I132202,I131809,I132233,I132250,I131800,I132281,I131803,I131815,I131812,I132370,I161187,I132396,I132413,I132362,I132435,I132452,I161190,I161208,I132469,I161196,I132495,I132503,I132529,I132537,I161205,I132554,I132341,I161199,I132594,I132602,I132335,I132350,I132647,I161202,I161184,I132664,I161193,I132690,I132338,I132712,I132729,I132746,I132353,I132777,I132794,I132344,I132825,I132347,I132359,I132356,I132914,I248712,I132940,I132957,I132979,I132996,I248706,I248703,I133013,I248718,I133039,I133047,I133073,I133081,I248700,I133098,I133138,I133146,I133191,I248715,I248709,I133208,I133234,I133256,I133273,I133290,I133321,I133338,I248721,I133369,I133458,I325016,I133484,I133501,I133450,I133523,I133540,I325028,I133557,I325019,I133583,I133591,I325037,I133617,I133625,I325013,I133642,I133429,I325031,I133682,I133690,I133423,I133438,I133735,I325025,I325022,I133752,I325034,I133778,I133426,I133800,I133817,I133834,I133441,I133865,I133882,I133432,I133913,I133435,I133447,I133444,I134002,I134028,I134045,I133994,I134067,I134084,I134101,I134127,I134135,I134161,I134169,I134186,I133973,I134226,I134234,I133967,I133982,I134279,I134296,I134322,I133970,I134344,I134361,I134378,I133985,I134409,I134426,I133976,I134457,I133979,I133991,I133988,I134546,I321613,I134572,I134589,I134538,I134611,I134628,I321631,I134645,I321625,I134671,I134679,I321619,I134705,I134713,I321628,I134730,I134517,I321616,I134770,I134778,I134511,I134526,I134823,I321634,I134840,I134866,I134514,I134888,I134905,I134922,I134529,I134953,I134970,I321622,I134520,I135001,I134523,I134535,I134532,I135090,I211728,I135116,I135133,I135082,I135155,I135172,I211749,I211740,I135189,I135215,I135223,I211734,I135249,I135257,I211731,I135274,I135061,I211725,I135314,I135322,I135055,I135070,I135367,I211737,I135384,I211746,I135410,I135058,I135432,I135449,I135466,I135073,I135497,I135514,I211743,I135064,I135545,I135067,I135079,I135076,I135634,I265576,I135660,I135677,I135626,I135699,I135716,I265570,I265567,I135733,I265582,I135759,I135767,I135793,I135801,I265564,I135818,I135605,I135858,I135866,I135599,I135614,I135911,I265579,I265573,I135928,I135954,I135602,I135976,I135993,I136010,I135617,I136041,I136058,I265585,I135608,I136089,I135611,I135623,I135620,I136178,I196700,I136204,I136221,I136243,I136260,I196721,I196712,I136277,I136303,I136311,I196706,I136337,I136345,I196703,I136362,I196697,I136402,I136410,I136455,I196709,I136472,I196718,I136498,I136520,I136537,I136554,I136585,I136602,I196715,I136633,I136722,I347558,I136748,I136765,I136714,I136787,I136804,I347570,I136821,I347561,I136847,I136855,I347579,I136881,I136889,I347555,I136906,I136693,I347573,I136946,I136954,I136687,I136702,I136999,I347567,I347564,I137016,I347576,I137042,I136690,I137064,I137081,I137098,I136705,I137129,I137146,I136696,I137177,I136699,I136711,I136708,I137266,I137292,I137309,I137331,I137348,I137365,I137391,I137399,I137425,I137433,I137450,I137490,I137498,I137543,I137560,I137586,I137608,I137625,I137642,I137673,I137690,I137721,I137810,I174158,I137836,I137853,I137802,I137875,I137892,I174155,I174176,I137909,I174179,I137935,I137943,I174164,I137969,I137977,I174167,I137994,I137781,I174170,I138034,I138042,I137775,I137790,I138087,I174161,I138104,I174173,I138130,I137778,I138152,I138169,I138186,I137793,I138217,I138234,I137784,I138265,I137787,I137799,I137796,I138354,I200168,I138380,I138397,I138346,I138419,I138436,I200189,I200180,I138453,I138479,I138487,I200174,I138513,I138521,I200171,I138538,I138325,I200165,I138578,I138586,I138319,I138334,I138631,I200177,I138648,I200186,I138674,I138322,I138696,I138713,I138730,I138337,I138761,I138778,I200183,I138328,I138809,I138331,I138343,I138340,I138898,I208838,I138924,I138941,I138890,I138963,I138980,I208859,I208850,I138997,I139023,I139031,I208844,I139057,I139065,I208841,I139082,I138869,I208835,I139122,I139130,I138863,I138878,I139175,I208847,I139192,I208856,I139218,I138866,I139240,I139257,I139274,I138881,I139305,I139322,I208853,I138872,I139353,I138875,I138887,I138884,I139442,I139468,I139485,I139507,I139524,I139541,I139567,I139575,I139601,I139609,I139626,I139666,I139674,I139719,I139736,I139762,I139784,I139801,I139818,I139849,I139866,I139897,I139986,I266103,I140012,I140029,I139978,I140051,I140068,I266097,I266094,I140085,I266109,I140111,I140119,I140145,I140153,I266091,I140170,I139957,I140210,I140218,I139951,I139966,I140263,I266106,I266100,I140280,I140306,I139954,I140328,I140345,I140362,I139969,I140393,I140410,I266112,I139960,I140441,I139963,I139975,I139972,I140530,I312637,I140556,I140573,I140522,I140595,I140612,I312655,I140629,I312649,I140655,I140663,I312643,I140689,I140697,I312652,I140714,I140501,I312640,I140754,I140762,I140495,I140510,I140807,I312658,I140824,I140850,I140498,I140872,I140889,I140906,I140513,I140937,I140954,I312646,I140504,I140985,I140507,I140519,I140516,I141074,I272370,I141100,I141117,I141066,I141139,I141156,I272385,I272373,I141173,I272364,I141199,I141207,I272376,I141233,I141241,I272367,I141258,I141045,I272382,I141298,I141306,I141039,I141054,I141351,I272391,I272379,I141368,I272388,I141394,I141042,I141416,I141433,I141450,I141057,I141481,I141498,I141048,I141529,I141051,I141063,I141060,I141618,I386537,I141644,I141661,I141683,I141700,I386534,I386531,I141717,I386519,I141743,I141751,I386543,I141777,I141785,I386528,I141802,I386522,I141842,I141850,I141895,I386525,I141912,I386540,I141938,I141960,I141977,I141994,I142025,I142042,I142073,I142162,I142188,I142205,I142227,I142244,I142261,I142287,I142295,I142321,I142329,I142346,I142386,I142394,I142439,I142456,I142482,I142504,I142521,I142538,I142569,I142586,I142617,I142706,I176470,I142732,I142749,I142698,I142771,I142788,I176467,I176488,I142805,I176491,I142831,I142839,I176476,I142865,I142873,I176479,I142890,I142677,I176482,I142930,I142938,I142671,I142686,I142983,I176473,I143000,I176485,I143026,I142674,I143048,I143065,I143082,I142689,I143113,I143130,I142680,I143161,I142683,I142695,I142692,I143250,I143276,I143293,I143242,I143315,I143332,I143349,I143375,I143383,I143409,I143417,I143434,I143221,I143474,I143482,I143215,I143230,I143527,I143544,I143570,I143218,I143592,I143609,I143626,I143233,I143657,I143674,I143224,I143705,I143227,I143239,I143236,I143794,I212306,I143820,I143837,I143786,I143859,I143876,I212327,I212318,I143893,I143919,I143927,I212312,I143953,I143961,I212309,I143978,I143765,I212303,I144018,I144026,I143759,I143774,I144071,I212315,I144088,I212324,I144114,I143762,I144136,I144153,I144170,I143777,I144201,I144218,I212321,I143768,I144249,I143771,I143783,I143780,I144338,I419441,I144364,I144381,I144330,I144403,I144420,I419417,I419438,I144437,I419435,I144463,I144471,I419414,I144497,I144505,I419426,I144522,I144309,I419429,I144562,I144570,I144303,I144318,I144615,I419432,I419420,I144632,I419423,I144658,I144306,I144680,I144697,I144714,I144321,I144745,I144762,I144312,I144793,I144315,I144327,I144324,I144882,I300794,I144908,I144925,I144947,I144964,I300809,I300797,I144981,I300788,I145007,I145015,I300800,I145041,I145049,I300791,I145066,I300806,I145106,I145114,I145159,I300815,I300803,I145176,I300812,I145202,I145224,I145241,I145258,I145289,I145306,I145337,I145426,I145452,I145469,I145418,I145491,I145508,I145525,I145551,I145559,I145585,I145593,I145610,I145397,I145650,I145658,I145391,I145406,I145703,I145720,I145746,I145394,I145768,I145785,I145802,I145409,I145833,I145850,I145400,I145881,I145403,I145415,I145412,I145970,I145996,I146013,I146035,I146052,I146069,I146095,I146103,I146129,I146137,I146154,I146194,I146202,I146247,I146264,I146290,I146312,I146329,I146346,I146377,I146394,I146425,I146514,I345824,I146540,I146557,I146579,I146596,I345836,I146613,I345827,I146639,I146647,I345845,I146673,I146681,I345821,I146698,I345839,I146738,I146746,I146791,I345833,I345830,I146808,I345842,I146834,I146856,I146873,I146890,I146921,I146938,I146969,I147058,I287228,I147084,I147101,I147050,I147123,I147140,I287243,I287231,I147157,I287222,I147183,I147191,I287234,I147217,I147225,I287225,I147242,I147029,I287240,I147282,I147290,I147023,I147038,I147335,I287249,I287237,I147352,I287246,I147378,I147026,I147400,I147417,I147434,I147041,I147465,I147482,I147032,I147513,I147035,I147047,I147044,I147602,I414681,I147628,I147645,I147667,I147684,I414657,I414678,I147701,I414675,I147727,I147735,I414654,I147761,I147769,I414666,I147786,I414669,I147826,I147834,I147879,I414672,I414660,I147896,I414663,I147922,I147944,I147961,I147978,I148009,I148026,I148057,I148146,I344668,I148172,I148189,I148211,I148228,I344680,I148245,I344671,I148271,I148279,I344689,I148305,I148313,I344665,I148330,I344683,I148370,I148378,I148423,I344677,I344674,I148440,I344686,I148466,I148488,I148505,I148522,I148553,I148570,I148601,I148690,I304670,I148716,I148733,I148682,I148755,I148772,I304685,I304673,I148789,I304664,I148815,I148823,I304676,I148849,I148857,I304667,I148874,I148661,I304682,I148914,I148922,I148655,I148670,I148967,I304691,I304679,I148984,I304688,I149010,I148658,I149032,I149049,I149066,I148673,I149097,I149114,I148664,I149145,I148667,I148679,I148676,I149234,I267157,I149260,I149277,I149226,I149299,I149316,I267151,I267148,I149333,I267163,I149359,I149367,I149393,I149401,I267145,I149418,I149205,I149458,I149466,I149199,I149214,I149511,I267160,I267154,I149528,I149554,I149202,I149576,I149593,I149610,I149217,I149641,I149658,I267166,I149208,I149689,I149211,I149223,I149220,I149778,I268738,I149804,I149821,I149843,I149860,I268732,I268729,I149877,I268744,I149903,I149911,I149937,I149945,I268726,I149962,I150002,I150010,I150055,I268741,I268735,I150072,I150098,I150120,I150137,I150154,I150185,I150202,I268747,I150233,I150322,I260833,I150348,I150365,I150314,I150387,I150404,I260827,I260824,I150421,I260839,I150447,I150455,I150481,I150489,I260821,I150506,I150293,I150546,I150554,I150287,I150302,I150599,I260836,I260830,I150616,I150642,I150290,I150664,I150681,I150698,I150305,I150729,I150746,I260842,I150296,I150777,I150299,I150311,I150308,I150866,I278830,I150892,I150909,I150858,I150931,I150948,I278845,I278833,I150965,I278824,I150991,I150999,I278836,I151025,I151033,I278827,I151050,I150837,I278842,I151090,I151098,I150831,I150846,I151143,I278851,I278839,I151160,I278848,I151186,I150834,I151208,I151225,I151242,I150849,I151273,I151290,I150840,I151321,I150843,I150855,I150852,I151410,I411111,I151436,I151453,I151402,I151475,I151492,I411087,I411108,I151509,I411105,I151535,I151543,I411084,I151569,I151577,I411096,I151594,I151381,I411099,I151634,I151642,I151375,I151390,I151687,I411102,I411090,I151704,I411093,I151730,I151378,I151752,I151769,I151786,I151393,I151817,I151834,I151384,I151865,I151387,I151399,I151396,I151954,I151980,I151997,I152019,I152036,I152053,I152079,I152087,I152113,I152121,I152138,I152178,I152186,I152231,I152248,I152274,I152296,I152313,I152330,I152361,I152378,I152409,I152498,I181672,I152524,I152541,I152490,I152563,I152580,I181669,I181690,I152597,I181693,I152623,I152631,I181678,I152657,I152665,I181681,I152682,I152469,I181684,I152722,I152730,I152463,I152478,I152775,I181675,I152792,I181687,I152818,I152466,I152840,I152857,I152874,I152481,I152905,I152922,I152472,I152953,I152475,I152487,I152484,I153042,I153068,I153085,I153034,I153107,I153124,I153141,I153167,I153175,I153201,I153209,I153226,I153013,I153266,I153274,I153007,I153022,I153319,I153336,I153362,I153010,I153384,I153401,I153418,I153025,I153449,I153466,I153016,I153497,I153019,I153031,I153028,I153586,I153612,I153629,I153651,I153668,I153685,I153711,I153719,I153745,I153753,I153770,I153810,I153818,I153863,I153880,I153906,I153928,I153945,I153962,I153993,I154010,I154041,I154130,I356228,I154156,I154173,I154122,I154195,I154212,I356240,I154229,I356231,I154255,I154263,I356249,I154289,I154297,I356225,I154314,I154101,I356243,I154354,I154362,I154095,I154110,I154407,I356237,I356234,I154424,I356246,I154450,I154098,I154472,I154489,I154506,I154113,I154537,I154554,I154104,I154585,I154107,I154119,I154116,I154671,I358555,I154697,I154714,I358537,I154745,I154753,I358543,I154770,I154787,I358558,I154804,I358549,I154821,I154838,I154855,I154886,I358561,I154903,I358540,I154920,I154965,I154982,I155013,I358546,I155030,I155061,I358552,I155078,I155095,I155121,I155129,I155160,I155177,I155208,I155266,I403349,I155292,I155309,I403355,I155340,I155348,I403370,I155365,I155382,I403361,I155399,I403358,I155416,I155433,I155450,I155481,I155498,I403373,I155515,I155560,I155577,I155608,I403367,I155625,I155656,I403352,I155673,I403364,I155690,I403376,I155716,I155724,I155755,I155772,I155803,I155861,I155887,I155904,I155853,I155935,I155943,I155960,I155977,I155994,I156011,I156028,I156045,I155850,I156076,I156093,I156110,I155835,I155847,I156155,I156172,I155841,I156203,I156220,I155829,I156251,I156268,I156285,I156311,I156319,I155838,I156350,I156367,I155844,I156398,I155832,I156456,I156482,I156499,I156530,I156538,I156555,I156572,I156589,I156606,I156623,I156640,I156671,I156688,I156705,I156750,I156767,I156798,I156815,I156846,I156863,I156880,I156906,I156914,I156945,I156962,I156993,I157051,I293051,I157077,I157094,I293039,I157125,I157133,I293036,I157150,I157167,I293048,I157184,I293045,I157201,I157218,I157235,I157266,I293054,I157283,I293057,I157300,I157345,I157362,I157393,I293060,I157410,I157441,I293063,I157458,I293042,I157475,I157501,I157509,I157540,I157557,I157588,I157646,I371389,I157672,I157689,I371404,I157720,I157728,I371413,I157745,I157762,I371392,I157779,I371398,I157796,I157813,I157830,I157861,I371410,I157878,I371407,I157895,I157940,I157957,I157988,I158005,I158036,I371401,I158053,I371395,I158070,I158096,I158104,I158135,I158152,I158183,I158241,I158267,I158284,I158233,I158315,I158323,I158340,I158357,I158374,I158391,I158408,I158425,I158230,I158456,I158473,I158490,I158215,I158227,I158535,I158552,I158221,I158583,I158600,I158209,I158631,I158648,I158665,I158691,I158699,I158218,I158730,I158747,I158224,I158778,I158212,I158836,I212890,I158862,I158879,I212884,I158910,I158918,I212881,I158935,I158952,I212893,I158969,I212896,I158986,I159003,I159020,I159051,I212905,I159068,I212899,I159085,I159130,I159147,I159178,I212887,I159195,I159226,I212902,I159243,I159260,I159286,I159294,I159325,I159342,I159373,I159431,I313759,I159457,I159474,I159423,I313762,I159505,I159513,I313765,I159530,I159547,I313777,I159564,I313768,I159581,I159598,I159615,I159420,I159646,I313774,I159663,I159680,I159405,I159417,I159725,I159742,I159411,I159773,I159790,I159399,I159821,I313771,I159838,I159855,I313780,I159881,I159889,I159408,I159920,I159937,I159414,I159968,I159402,I160026,I160052,I160069,I160018,I160100,I160108,I160125,I160142,I160159,I160176,I160193,I160210,I160015,I160241,I160258,I160275,I160000,I160012,I160320,I160337,I160006,I160368,I160385,I159994,I160416,I160433,I160450,I160476,I160484,I160003,I160515,I160532,I160009,I160563,I159997,I160621,I382482,I160647,I160664,I160613,I382488,I160695,I160703,I382476,I160720,I160737,I382479,I160754,I382485,I160771,I160788,I160805,I160610,I160836,I160853,I382494,I160870,I160595,I160607,I160915,I160932,I160601,I160963,I382473,I160980,I160589,I161011,I382497,I161028,I161045,I382491,I161071,I161079,I160598,I161110,I161127,I160604,I161158,I160592,I161216,I161242,I161259,I161290,I161298,I161315,I161332,I161349,I161366,I161383,I161400,I161431,I161448,I161465,I161510,I161527,I161558,I161575,I161606,I161623,I161640,I161666,I161674,I161705,I161722,I161753,I161811,I161837,I161854,I161803,I161885,I161893,I161910,I161927,I161944,I161961,I161978,I161995,I161800,I162026,I162043,I162060,I161785,I161797,I162105,I162122,I161791,I162153,I162170,I161779,I162201,I162218,I162235,I162261,I162269,I161788,I162300,I162317,I161794,I162348,I161782,I162406,I249763,I162432,I162449,I162398,I249760,I162480,I162488,I162505,I162522,I249757,I162539,I249772,I162556,I162573,I162590,I162395,I162621,I249766,I162638,I249754,I162655,I162380,I162392,I162700,I162717,I162386,I162748,I249775,I162765,I162374,I162796,I162813,I249769,I162830,I162856,I162864,I162383,I162895,I162912,I162389,I162943,I162377,I163001,I163027,I163044,I162993,I163075,I163083,I163100,I163117,I163134,I163151,I163168,I163185,I162990,I163216,I163233,I163250,I162975,I162987,I163295,I163312,I162981,I163343,I163360,I162969,I163391,I163408,I163425,I163451,I163459,I162978,I163490,I163507,I162984,I163538,I162972,I163596,I163622,I163639,I163670,I163678,I163695,I163712,I163729,I163746,I163763,I163780,I163811,I163828,I163845,I163890,I163907,I163938,I163955,I163986,I164003,I164020,I164046,I164054,I164085,I164102,I164133,I164191,I314320,I164217,I164234,I314323,I164265,I164273,I314326,I164290,I164307,I314338,I164324,I314329,I164341,I164358,I164375,I164406,I314335,I164423,I164440,I164485,I164502,I164533,I164550,I164581,I314332,I164598,I164615,I314341,I164641,I164649,I164680,I164697,I164728,I164786,I164812,I164829,I164860,I164868,I164885,I164902,I164919,I164936,I164953,I164970,I165001,I165018,I165035,I165080,I165097,I165128,I165145,I165176,I165193,I165210,I165236,I165244,I165275,I165292,I165323,I165381,I165407,I165424,I165373,I165455,I165463,I165480,I165497,I165514,I165531,I165548,I165565,I165370,I165596,I165613,I165630,I165355,I165367,I165675,I165692,I165361,I165723,I165740,I165349,I165771,I165788,I165805,I165831,I165839,I165358,I165870,I165887,I165364,I165918,I165352,I165976,I333123,I166002,I166019,I333105,I166050,I166058,I333111,I166075,I166092,I333126,I166109,I333117,I166126,I166143,I166160,I166191,I333129,I166208,I333108,I166225,I166270,I166287,I166318,I333114,I166335,I166366,I333120,I166383,I166400,I166426,I166434,I166465,I166482,I166513,I166571,I274963,I166597,I166614,I166563,I274951,I166645,I166653,I274948,I166670,I166687,I274960,I166704,I274957,I166721,I166738,I166755,I166560,I166786,I274966,I166803,I274969,I166820,I166545,I166557,I166865,I166882,I166551,I166913,I274972,I166930,I166539,I166961,I274975,I166978,I274954,I166995,I167021,I167029,I166548,I167060,I167077,I166554,I167108,I166542,I167166,I167192,I167209,I167158,I167240,I167248,I167265,I167282,I167299,I167316,I167333,I167350,I167155,I167381,I167398,I167415,I167140,I167152,I167460,I167477,I167146,I167508,I167525,I167134,I167556,I167573,I167590,I167616,I167624,I167143,I167655,I167672,I167149,I167703,I167137,I167761,I267681,I167787,I167804,I267678,I167835,I167843,I167860,I167877,I267675,I167894,I267690,I167911,I167928,I167945,I167976,I267684,I167993,I267672,I168010,I168055,I168072,I168103,I267693,I168120,I168151,I168168,I267687,I168185,I168211,I168219,I168250,I168267,I168298,I168356,I168382,I168399,I168430,I168438,I168455,I168472,I168489,I168506,I168523,I168540,I168571,I168588,I168605,I168650,I168667,I168698,I168715,I168746,I168763,I168780,I168806,I168814,I168845,I168862,I168893,I168951,I195550,I168977,I168994,I168943,I195544,I169025,I169033,I195541,I169050,I169067,I195553,I169084,I195556,I169101,I169118,I169135,I168940,I169166,I195565,I169183,I195559,I169200,I168925,I168937,I169245,I169262,I168931,I169293,I195547,I169310,I168919,I169341,I195562,I169358,I169375,I169401,I169409,I168928,I169440,I169457,I168934,I169488,I168922,I169546,I169572,I169589,I169620,I169628,I169645,I169662,I169679,I169696,I169713,I169730,I169761,I169778,I169795,I169840,I169857,I169888,I169905,I169936,I169953,I169970,I169996,I170004,I170035,I170052,I170083,I170141,I265043,I170167,I170175,I170201,I170209,I265040,I170226,I265055,I170243,I170260,I265049,I170277,I170127,I170308,I170325,I170342,I265046,I170359,I265037,I170124,I170115,I170404,I170118,I170112,I170449,I265058,I170466,I170483,I170121,I170514,I170531,I170548,I265052,I170574,I170582,I170109,I170133,I170627,I170644,I170661,I170130,I170719,I337729,I170745,I170753,I337735,I170779,I170787,I170804,I337732,I170821,I170838,I337750,I170855,I170886,I170903,I170920,I337753,I170937,I170982,I171027,I337738,I171044,I171061,I171092,I337744,I171109,I337741,I171126,I337747,I171152,I171160,I171205,I171222,I171239,I171297,I171323,I171331,I171357,I171365,I171382,I171399,I171416,I171433,I171464,I171481,I171498,I171515,I171560,I171605,I171622,I171639,I171670,I171687,I171704,I171730,I171738,I171783,I171800,I171817,I171875,I171901,I171909,I171935,I171943,I171960,I171977,I171994,I172011,I172042,I172059,I172076,I172093,I172138,I172183,I172200,I172217,I172248,I172265,I172282,I172308,I172316,I172361,I172378,I172395,I172453,I213459,I172479,I172487,I213471,I172513,I172521,I213462,I172538,I213465,I172555,I172572,I213468,I172589,I172439,I172620,I172637,I172654,I172671,I213474,I172436,I172427,I172716,I172430,I172424,I172761,I213480,I172778,I172795,I172433,I172826,I172843,I213477,I172860,I213483,I172886,I172894,I172421,I172445,I172939,I172956,I172973,I172442,I173031,I173057,I173065,I173091,I173099,I173116,I173133,I173150,I173167,I173198,I173215,I173232,I173249,I173294,I173339,I173356,I173373,I173404,I173421,I173438,I173464,I173472,I173517,I173534,I173551,I173609,I173635,I173643,I173669,I173677,I173694,I173711,I173728,I173745,I173595,I173776,I173793,I173810,I173827,I173592,I173583,I173872,I173586,I173580,I173917,I173934,I173951,I173589,I173982,I173999,I174016,I174042,I174050,I173577,I173601,I174095,I174112,I174129,I173598,I174187,I174213,I174221,I174247,I174255,I174272,I174289,I174306,I174323,I174354,I174371,I174388,I174405,I174450,I174495,I174512,I174529,I174560,I174577,I174594,I174620,I174628,I174673,I174690,I174707,I174765,I412274,I174791,I174799,I174825,I174833,I412298,I174850,I412280,I174867,I174884,I412295,I174901,I174932,I174949,I174966,I412277,I174983,I412286,I175028,I175073,I412283,I175090,I175107,I175138,I412292,I175155,I412301,I175172,I412289,I175198,I175206,I175251,I175268,I175285,I175343,I357381,I175369,I175377,I357387,I175403,I175411,I175428,I357384,I175445,I175462,I357402,I175479,I175329,I175510,I175527,I175544,I357405,I175561,I175326,I175317,I175606,I175320,I175314,I175651,I357390,I175668,I175685,I175323,I175716,I357396,I175733,I357393,I175750,I357399,I175776,I175784,I175311,I175335,I175829,I175846,I175863,I175332,I175921,I175947,I175955,I175981,I175989,I176006,I176023,I176040,I176057,I175907,I176088,I176105,I176122,I176139,I175904,I175895,I176184,I175898,I175892,I176229,I176246,I176263,I175901,I176294,I176311,I176328,I176354,I176362,I175889,I175913,I176407,I176424,I176441,I175910,I176499,I176525,I176533,I176559,I176567,I176584,I176601,I176618,I176635,I176666,I176683,I176700,I176717,I176762,I176807,I176824,I176841,I176872,I176889,I176906,I176932,I176940,I176985,I177002,I177019,I177077,I369775,I177103,I177111,I369769,I177137,I177145,I369778,I177162,I369757,I177179,I177196,I369766,I177213,I177244,I177261,I177278,I369781,I177295,I369760,I177340,I177385,I369763,I177402,I177419,I177450,I369772,I177467,I177484,I177510,I177518,I177563,I177580,I177597,I177655,I375215,I177681,I177689,I375209,I177715,I177723,I375218,I177740,I375197,I177757,I177774,I375206,I177791,I177822,I177839,I177856,I375221,I177873,I375200,I177918,I177963,I375203,I177980,I177997,I178028,I375212,I178045,I178062,I178088,I178096,I178141,I178158,I178175,I178233,I243436,I178259,I178267,I178293,I178301,I243433,I178318,I243448,I178335,I178352,I243442,I178369,I178219,I178400,I178417,I178434,I243439,I178451,I243430,I178216,I178207,I178496,I178210,I178204,I178541,I243451,I178558,I178575,I178213,I178606,I178623,I178640,I243445,I178666,I178674,I178201,I178225,I178719,I178736,I178753,I178222,I178811,I178837,I178845,I178871,I178879,I178896,I178913,I178930,I178947,I178797,I178978,I178995,I179012,I179029,I178794,I178785,I179074,I178788,I178782,I179119,I179136,I179153,I178791,I179184,I179201,I179218,I179244,I179252,I178779,I178803,I179297,I179314,I179331,I178800,I179389,I179415,I179423,I179449,I179457,I179474,I179491,I179508,I179525,I179375,I179556,I179573,I179590,I179607,I179372,I179363,I179652,I179366,I179360,I179697,I179714,I179731,I179369,I179762,I179779,I179796,I179822,I179830,I179357,I179381,I179875,I179892,I179909,I179378,I179967,I179993,I180001,I180027,I180035,I180052,I180069,I180086,I180103,I179953,I180134,I180151,I180168,I180185,I179950,I179941,I180230,I179944,I179938,I180275,I180292,I180309,I179947,I180340,I180357,I180374,I180400,I180408,I179935,I179959,I180453,I180470,I180487,I179956,I180545,I180571,I180579,I180605,I180613,I180630,I180647,I180664,I180681,I180531,I180712,I180729,I180746,I180763,I180528,I180519,I180808,I180522,I180516,I180853,I180870,I180887,I180525,I180918,I180935,I180952,I180978,I180986,I180513,I180537,I181031,I181048,I181065,I180534,I181123,I405729,I181149,I181157,I181183,I181191,I405753,I181208,I405735,I181225,I181242,I405750,I181259,I181290,I181307,I181324,I405732,I181341,I405741,I181386,I181431,I405738,I181448,I181465,I181496,I405747,I181513,I405756,I181530,I405744,I181556,I181564,I181609,I181626,I181643,I181701,I214615,I181727,I181735,I214627,I181761,I181769,I214618,I181786,I214621,I181803,I181820,I214624,I181837,I181868,I181885,I181902,I181919,I214630,I181964,I182009,I214636,I182026,I182043,I182074,I182091,I214633,I182108,I214639,I182134,I182142,I182187,I182204,I182221,I182279,I182305,I182313,I182339,I182347,I182364,I182381,I182398,I182415,I182446,I182463,I182480,I182497,I182542,I182587,I182604,I182621,I182652,I182669,I182686,I182712,I182720,I182765,I182782,I182799,I182857,I182883,I182891,I182917,I182925,I182942,I182959,I182976,I182993,I182843,I183024,I183041,I183058,I183075,I182840,I182831,I183120,I182834,I182828,I183165,I183182,I183199,I182837,I183230,I183247,I183264,I183290,I183298,I182825,I182849,I183343,I183360,I183377,I182846,I183435,I183461,I183469,I183495,I183503,I183520,I183537,I183554,I183571,I183421,I183602,I183619,I183636,I183653,I183418,I183409,I183698,I183412,I183406,I183743,I183760,I183777,I183415,I183808,I183825,I183842,I183868,I183876,I183403,I183427,I183921,I183938,I183955,I183424,I184013,I184039,I184047,I184073,I184081,I184098,I184115,I184132,I184149,I184180,I184197,I184214,I184231,I184276,I184321,I184338,I184355,I184386,I184403,I184420,I184446,I184454,I184499,I184516,I184533,I184591,I184617,I184625,I184651,I184659,I184676,I184693,I184710,I184727,I184758,I184775,I184792,I184809,I184854,I184899,I184916,I184933,I184964,I184981,I184998,I185024,I185032,I185077,I185094,I185111,I185169,I251341,I185195,I185203,I185229,I185237,I251338,I185254,I251353,I185271,I185288,I251347,I185305,I185155,I185336,I185353,I185370,I251344,I185387,I251335,I185152,I185143,I185432,I185146,I185140,I185477,I251356,I185494,I185511,I185149,I185542,I185559,I185576,I251350,I185602,I185610,I185137,I185161,I185655,I185672,I185689,I185158,I185747,I185773,I185781,I185807,I185815,I185832,I185849,I185866,I185883,I185733,I185914,I185931,I185948,I185965,I185730,I185721,I186010,I185724,I185718,I186055,I186072,I186089,I185727,I186120,I186137,I186154,I186180,I186188,I185715,I185739,I186233,I186250,I186267,I185736,I186325,I186351,I186359,I186385,I186393,I186410,I186427,I186444,I186461,I186311,I186492,I186509,I186526,I186543,I186308,I186299,I186588,I186302,I186296,I186633,I186650,I186667,I186305,I186698,I186715,I186732,I186758,I186766,I186293,I186317,I186811,I186828,I186845,I186314,I186903,I232533,I186929,I186937,I232545,I186963,I186971,I232536,I186988,I232539,I187005,I187022,I232542,I187039,I186889,I187070,I187087,I187104,I187121,I232548,I186886,I186877,I187166,I186880,I186874,I187211,I232554,I187228,I187245,I186883,I187276,I187293,I232551,I187310,I232557,I187336,I187344,I186871,I186895,I187389,I187406,I187423,I186892,I187481,I187507,I187515,I187541,I187549,I187566,I187583,I187600,I187617,I187467,I187648,I187665,I187682,I187699,I187464,I187455,I187744,I187458,I187452,I187789,I187806,I187823,I187461,I187854,I187871,I187888,I187914,I187922,I187449,I187473,I187967,I187984,I188001,I187470,I188059,I346977,I188085,I188093,I346983,I188119,I188127,I188144,I346980,I188161,I188178,I346998,I188195,I188226,I188243,I188260,I347001,I188277,I188322,I188367,I346986,I188384,I188401,I188432,I346992,I188449,I346989,I188466,I346995,I188492,I188500,I188545,I188562,I188579,I188637,I188663,I188671,I188697,I188705,I188722,I188739,I188756,I188773,I188623,I188804,I188821,I188838,I188855,I188620,I188611,I188900,I188614,I188608,I188945,I188962,I188979,I188617,I189010,I189027,I189044,I189070,I189078,I188605,I188629,I189123,I189140,I189157,I188626,I189215,I282060,I189241,I189249,I282057,I189275,I189283,I282054,I189300,I282081,I189317,I189334,I282069,I189351,I189201,I189382,I189399,I189416,I282075,I189433,I282066,I189198,I189189,I189478,I189192,I189186,I189523,I282063,I189540,I189557,I189195,I189588,I282078,I189605,I282072,I189622,I189648,I189656,I189183,I189207,I189701,I189718,I189735,I189204,I189793,I189819,I189827,I189853,I189861,I189878,I189895,I189912,I189929,I189779,I189960,I189977,I189994,I190011,I189776,I189767,I190056,I189770,I189764,I190101,I190118,I190135,I189773,I190166,I190183,I190200,I190226,I190234,I189761,I189785,I190279,I190296,I190313,I189782,I190371,I339463,I190397,I190405,I339469,I190431,I190439,I190456,I339466,I190473,I190490,I339484,I190507,I190357,I190538,I190555,I190572,I339487,I190589,I190354,I190345,I190634,I190348,I190342,I190679,I339472,I190696,I190713,I190351,I190744,I339478,I190761,I339475,I190778,I339481,I190804,I190812,I190339,I190363,I190857,I190874,I190891,I190360,I190949,I313219,I190975,I190983,I313210,I191009,I191017,I313204,I191034,I313216,I191051,I191068,I313207,I191085,I191116,I191133,I191150,I313213,I191167,I313198,I191212,I191257,I191274,I191291,I191322,I313201,I191339,I191356,I191382,I191390,I191435,I191452,I191469,I191527,I191553,I191561,I191587,I191595,I191612,I191629,I191646,I191663,I191513,I191694,I191711,I191728,I191745,I191510,I191501,I191790,I191504,I191498,I191835,I191852,I191869,I191507,I191900,I191917,I191934,I191960,I191968,I191495,I191519,I192013,I192030,I192047,I191516,I192105,I335417,I192131,I192139,I335423,I192165,I192173,I192190,I335420,I192207,I192224,I335438,I192241,I192091,I192272,I192289,I192306,I335441,I192323,I192088,I192079,I192368,I192082,I192076,I192413,I335426,I192430,I192447,I192085,I192478,I335432,I192495,I335429,I192512,I335435,I192538,I192546,I192073,I192097,I192591,I192608,I192625,I192094,I192683,I325591,I192709,I192717,I325597,I192743,I192751,I192768,I325594,I192785,I192802,I325612,I192819,I192669,I192850,I192867,I192884,I325615,I192901,I192666,I192657,I192946,I192660,I192654,I192991,I325600,I193008,I193025,I192663,I193056,I325606,I193073,I325603,I193090,I325609,I193116,I193124,I192651,I192675,I193169,I193186,I193203,I192672,I193261,I193287,I193295,I193321,I193329,I193346,I193363,I193380,I193397,I193247,I193428,I193445,I193462,I193479,I193244,I193235,I193524,I193238,I193232,I193569,I193586,I193603,I193241,I193634,I193651,I193668,I193694,I193702,I193229,I193253,I193747,I193764,I193781,I193250,I193839,I363757,I193865,I193873,I193890,I363739,I363751,I193907,I363754,I193933,I193941,I363748,I363745,I193967,I193975,I193992,I194009,I194026,I363763,I194066,I194074,I194091,I194108,I194125,I194156,I363742,I194173,I194199,I194207,I194238,I194269,I194286,I194317,I363760,I194417,I194443,I194451,I194468,I194485,I194511,I194519,I194545,I194553,I194570,I194587,I194604,I194400,I194644,I194652,I194669,I194686,I194703,I194403,I194734,I194751,I194777,I194785,I194385,I194816,I194394,I194847,I194864,I194406,I194895,I194397,I194388,I194391,I194409,I194995,I195021,I195029,I195046,I195063,I195089,I195097,I195123,I195131,I195148,I195165,I195182,I195222,I195230,I195247,I195264,I195281,I195312,I195329,I195355,I195363,I195394,I195425,I195442,I195473,I195573,I195599,I195607,I195624,I195641,I195667,I195675,I195701,I195709,I195726,I195743,I195760,I195800,I195808,I195825,I195842,I195859,I195890,I195907,I195933,I195941,I195972,I196003,I196020,I196051,I196151,I196177,I196185,I196202,I196219,I196245,I196253,I196279,I196287,I196304,I196321,I196338,I196378,I196386,I196403,I196420,I196437,I196468,I196485,I196511,I196519,I196550,I196581,I196598,I196629,I196729,I273034,I196755,I196763,I196780,I273010,I273025,I196797,I273037,I196823,I196831,I273022,I273013,I196857,I196865,I196882,I196899,I196916,I196956,I196964,I196981,I196998,I197015,I197046,I273028,I273019,I197063,I273031,I197089,I197097,I197128,I197159,I197176,I197207,I273016,I197307,I197333,I197341,I197358,I197375,I197401,I197409,I197435,I197443,I197460,I197477,I197494,I197290,I197534,I197542,I197559,I197576,I197593,I197293,I197624,I197641,I197667,I197675,I197275,I197706,I197284,I197737,I197754,I197296,I197785,I197287,I197278,I197281,I197299,I197885,I197911,I197919,I197936,I197953,I197979,I197987,I198013,I198021,I198038,I198055,I198072,I198112,I198120,I198137,I198154,I198171,I198202,I198219,I198245,I198253,I198284,I198315,I198332,I198363,I198463,I360289,I198489,I198497,I198514,I360271,I360283,I198531,I360286,I198557,I198565,I360280,I360277,I198591,I198599,I198616,I198633,I198650,I360295,I198690,I198698,I198715,I198732,I198749,I198780,I360274,I198797,I198823,I198831,I198862,I198893,I198910,I198941,I360292,I199041,I199067,I199075,I199092,I199109,I199135,I199143,I199169,I199177,I199194,I199211,I199228,I199268,I199276,I199293,I199310,I199327,I199358,I199375,I199401,I199409,I199440,I199471,I199488,I199519,I199619,I370845,I199645,I199653,I199670,I370848,I370857,I199687,I370860,I199713,I199721,I370869,I370851,I199747,I199755,I199772,I199789,I199806,I199602,I199846,I199854,I199871,I199888,I199905,I199605,I199936,I370866,I199953,I370863,I199979,I199987,I199587,I200018,I199596,I200049,I200066,I199608,I200097,I370854,I199599,I199590,I199593,I199611,I200197,I200223,I200231,I200248,I200265,I200291,I200299,I200325,I200333,I200350,I200367,I200384,I200424,I200432,I200449,I200466,I200483,I200514,I200531,I200557,I200565,I200596,I200627,I200644,I200675,I200775,I308564,I200801,I200809,I200826,I308540,I308555,I200843,I308567,I200869,I200877,I308552,I308543,I200903,I200911,I200928,I200945,I200962,I201002,I201010,I201027,I201044,I201061,I201092,I308558,I308549,I201109,I308561,I201135,I201143,I201174,I201205,I201222,I201253,I308546,I201353,I201379,I201387,I201404,I201421,I201447,I201455,I201481,I201489,I201506,I201523,I201540,I201580,I201588,I201605,I201622,I201639,I201670,I201687,I201713,I201721,I201752,I201783,I201800,I201831,I201931,I201957,I201965,I201982,I201999,I202025,I202033,I202059,I202067,I202084,I202101,I202118,I201914,I202158,I202166,I202183,I202200,I202217,I201917,I202248,I202265,I202291,I202299,I201899,I202330,I201908,I202361,I202378,I201920,I202409,I201911,I201902,I201905,I201923,I202509,I381895,I202535,I202543,I202560,I381919,I381901,I202577,I381907,I202603,I202611,I381913,I381898,I202637,I202645,I202662,I202679,I202696,I202492,I381910,I202736,I202744,I202761,I202778,I202795,I202495,I202826,I381916,I381904,I202843,I202869,I202877,I202477,I202908,I202486,I202939,I202956,I202498,I202987,I202489,I202480,I202483,I202501,I203087,I409326,I203113,I203121,I203138,I409311,I409299,I203155,I409314,I203181,I203189,I409317,I203215,I203223,I203240,I203257,I203274,I409305,I203314,I203322,I203339,I203356,I203373,I203404,I409302,I409308,I203421,I409323,I203447,I203455,I203486,I203517,I203534,I203565,I409320,I203665,I203691,I203699,I203716,I203733,I203759,I203767,I203793,I203801,I203818,I203835,I203852,I203892,I203900,I203917,I203934,I203951,I203982,I203999,I204025,I204033,I204064,I204095,I204112,I204143,I204243,I204269,I204277,I204294,I204311,I204337,I204345,I204371,I204379,I204396,I204413,I204430,I204470,I204478,I204495,I204512,I204529,I204560,I204577,I204603,I204611,I204642,I204673,I204690,I204721,I204821,I349307,I204847,I204855,I204872,I349289,I349301,I204889,I349304,I204915,I204923,I349298,I349295,I204949,I204957,I204974,I204991,I205008,I204804,I349313,I205048,I205056,I205073,I205090,I205107,I204807,I205138,I349292,I205155,I205181,I205189,I204789,I205220,I204798,I205251,I205268,I204810,I205299,I349310,I204801,I204792,I204795,I204813,I205399,I205425,I205433,I205450,I205467,I205493,I205501,I205527,I205535,I205552,I205569,I205586,I205626,I205634,I205651,I205668,I205685,I205716,I205733,I205759,I205767,I205798,I205829,I205846,I205877,I205977,I383051,I206003,I206011,I206028,I383075,I383057,I206045,I383063,I206071,I206079,I383069,I383054,I206105,I206113,I206130,I206147,I206164,I205960,I383066,I206204,I206212,I206229,I206246,I206263,I205963,I206294,I383072,I383060,I206311,I206337,I206345,I205945,I206376,I205954,I206407,I206424,I205966,I206455,I205957,I205948,I205951,I205969,I206555,I206581,I206589,I206606,I206623,I206649,I206657,I206683,I206691,I206708,I206725,I206742,I206782,I206790,I206807,I206824,I206841,I206872,I206889,I206915,I206923,I206954,I206985,I207002,I207033,I207133,I207159,I207167,I207184,I207201,I207227,I207235,I207261,I207269,I207286,I207303,I207320,I207360,I207368,I207385,I207402,I207419,I207450,I207467,I207493,I207501,I207532,I207563,I207580,I207611,I207711,I207737,I207745,I207762,I207779,I207805,I207813,I207839,I207847,I207864,I207881,I207898,I207938,I207946,I207963,I207980,I207997,I208028,I208045,I208071,I208079,I208110,I208141,I208158,I208189,I208289,I208315,I208323,I208340,I208357,I208383,I208391,I208417,I208425,I208442,I208459,I208476,I208516,I208524,I208541,I208558,I208575,I208606,I208623,I208649,I208657,I208688,I208719,I208736,I208767,I208867,I359711,I208893,I208901,I208918,I359693,I359705,I208935,I359708,I208961,I208969,I359702,I359699,I208995,I209003,I209020,I209037,I209054,I359717,I209094,I209102,I209119,I209136,I209153,I209184,I359696,I209201,I209227,I209235,I209266,I209297,I209314,I209345,I359714,I209445,I209471,I209479,I209496,I209513,I209539,I209547,I209573,I209581,I209598,I209615,I209632,I209672,I209680,I209697,I209714,I209731,I209762,I209779,I209805,I209813,I209844,I209875,I209892,I209923,I210023,I391721,I210049,I210057,I210074,I391745,I391727,I210091,I391733,I210117,I210125,I391739,I391724,I210151,I210159,I210176,I210193,I210210,I210006,I391736,I210250,I210258,I210275,I210292,I210309,I210009,I210340,I391742,I391730,I210357,I210383,I210391,I209991,I210422,I210000,I210453,I210470,I210012,I210501,I210003,I209994,I209997,I210015,I210601,I210627,I210635,I210652,I210669,I210695,I210703,I210729,I210737,I210754,I210771,I210788,I210584,I210828,I210836,I210853,I210870,I210887,I210587,I210918,I210935,I210961,I210969,I210569,I211000,I210578,I211031,I211048,I210590,I211079,I210581,I210572,I210575,I210593,I211179,I211205,I211213,I211230,I211247,I211273,I211281,I211307,I211315,I211332,I211349,I211366,I211162,I211406,I211414,I211431,I211448,I211465,I211165,I211496,I211513,I211539,I211547,I211147,I211578,I211156,I211609,I211626,I211168,I211657,I211159,I211150,I211153,I211171,I211757,I250296,I211783,I211791,I211808,I250284,I250302,I211825,I250299,I211851,I211859,I250290,I250287,I211885,I211893,I211910,I211927,I211944,I250281,I211984,I211992,I212009,I212026,I212043,I212074,I212091,I212117,I212125,I212156,I212187,I212204,I212235,I250293,I212335,I268214,I212361,I212369,I212386,I268202,I268220,I212403,I268217,I212429,I212437,I268208,I268205,I212463,I212471,I212488,I212505,I212522,I268199,I212562,I212570,I212587,I212604,I212621,I212652,I212669,I212695,I212703,I212734,I212765,I212782,I212813,I268211,I212913,I414086,I212939,I212947,I212964,I414071,I414059,I212981,I414074,I213007,I213015,I414077,I213041,I213049,I213066,I213083,I213100,I414065,I213140,I213148,I213165,I213182,I213199,I213230,I414062,I414068,I213247,I414083,I213273,I213281,I213312,I213343,I213360,I213391,I414080,I213491,I213517,I213525,I213542,I213559,I213585,I213593,I213619,I213627,I213644,I213661,I213678,I213718,I213726,I213743,I213760,I213777,I213808,I213825,I213851,I213859,I213890,I213921,I213938,I213969,I214069,I214095,I214103,I214120,I214137,I214163,I214171,I214197,I214205,I214222,I214239,I214256,I214052,I214296,I214304,I214321,I214338,I214355,I214055,I214386,I214403,I214429,I214437,I214037,I214468,I214046,I214499,I214516,I214058,I214547,I214049,I214040,I214043,I214061,I214647,I214673,I214681,I214698,I214715,I214741,I214749,I214775,I214783,I214800,I214817,I214834,I214874,I214882,I214899,I214916,I214933,I214964,I214981,I215007,I215015,I215046,I215077,I215094,I215125,I215225,I215251,I215259,I215276,I215293,I215319,I215327,I215353,I215361,I215378,I215395,I215412,I215452,I215460,I215477,I215494,I215511,I215542,I215559,I215585,I215593,I215624,I215655,I215672,I215703,I215803,I215829,I215837,I215854,I215871,I215897,I215905,I215931,I215939,I215956,I215973,I215990,I215786,I216030,I216038,I216055,I216072,I216089,I215789,I216120,I216137,I216163,I216171,I215771,I216202,I215780,I216233,I216250,I215792,I216281,I215783,I215774,I215777,I215795,I216381,I398616,I216407,I216415,I216432,I398601,I398589,I216449,I398604,I216475,I216483,I398607,I216509,I216517,I216534,I216551,I216568,I216364,I398595,I216608,I216616,I216633,I216650,I216667,I216367,I216698,I398592,I398598,I216715,I398613,I216741,I216749,I216349,I216780,I216358,I216811,I216828,I216370,I216859,I398610,I216361,I216352,I216355,I216373,I216959,I216985,I216993,I217010,I217027,I217053,I217061,I217087,I217095,I217112,I217129,I217146,I217186,I217194,I217211,I217228,I217245,I217276,I217293,I217319,I217327,I217358,I217389,I217406,I217437,I217537,I355665,I217563,I217571,I217588,I355647,I355659,I217605,I355662,I217631,I217639,I355656,I355653,I217665,I217673,I217690,I217707,I217724,I217520,I355671,I217764,I217772,I217789,I217806,I217823,I217523,I217854,I355650,I217871,I217897,I217905,I217505,I217936,I217514,I217967,I217984,I217526,I218015,I355668,I217517,I217508,I217511,I217529,I218115,I218141,I218149,I218166,I218183,I218209,I218217,I218243,I218251,I218268,I218285,I218302,I218098,I218342,I218350,I218367,I218384,I218401,I218101,I218432,I218449,I218475,I218483,I218083,I218514,I218092,I218545,I218562,I218104,I218593,I218095,I218086,I218089,I218107,I218693,I218719,I218727,I218744,I218761,I218787,I218795,I218821,I218829,I218846,I218863,I218880,I218920,I218928,I218945,I218962,I218979,I219010,I219027,I219053,I219061,I219092,I219123,I219140,I219171,I219271,I219297,I219305,I219322,I219339,I219365,I219373,I219399,I219407,I219424,I219441,I219458,I219254,I219498,I219506,I219523,I219540,I219557,I219257,I219588,I219605,I219631,I219639,I219239,I219670,I219248,I219701,I219718,I219260,I219749,I219251,I219242,I219245,I219263,I219849,I249242,I219875,I219883,I219900,I249230,I249248,I219917,I249245,I219943,I219951,I249236,I249233,I219977,I219985,I220002,I220019,I220036,I219832,I249227,I220076,I220084,I220101,I220118,I220135,I219835,I220166,I220183,I220209,I220217,I219817,I220248,I219826,I220279,I220296,I219838,I220327,I249239,I219829,I219820,I219823,I219841,I220427,I284662,I220453,I220461,I220478,I284638,I284653,I220495,I284665,I220521,I220529,I284650,I284641,I220555,I220563,I220580,I220597,I220614,I220410,I220654,I220662,I220679,I220696,I220713,I220413,I220744,I284656,I284647,I220761,I284659,I220787,I220795,I220395,I220826,I220404,I220857,I220874,I220416,I220905,I284644,I220407,I220398,I220401,I220419,I221005,I363179,I221031,I221039,I221056,I363161,I363173,I221073,I363176,I221099,I221107,I363170,I363167,I221133,I221141,I221158,I221175,I221192,I363185,I221232,I221240,I221257,I221274,I221291,I221322,I363164,I221339,I221365,I221373,I221404,I221435,I221452,I221483,I363182,I221583,I221609,I221617,I221634,I221651,I221677,I221685,I221711,I221719,I221736,I221753,I221770,I221566,I221810,I221818,I221835,I221852,I221869,I221569,I221900,I221917,I221943,I221951,I221551,I221982,I221560,I222013,I222030,I221572,I222061,I221563,I221554,I221557,I221575,I222161,I251877,I222187,I222195,I222212,I251865,I251883,I222229,I251880,I222255,I222263,I251871,I251868,I222289,I222297,I222314,I222331,I222348,I251862,I222388,I222396,I222413,I222430,I222447,I222478,I222495,I222521,I222529,I222560,I222591,I222608,I222639,I251874,I222739,I222765,I222773,I222790,I222807,I222833,I222841,I222867,I222875,I222892,I222909,I222926,I222722,I222966,I222974,I222991,I223008,I223025,I222725,I223056,I223073,I223099,I223107,I222707,I223138,I222716,I223169,I223186,I222728,I223217,I222719,I222710,I222713,I222731,I223317,I223343,I223351,I223368,I223385,I223411,I223419,I223445,I223453,I223470,I223487,I223504,I223300,I223544,I223552,I223569,I223586,I223603,I223303,I223634,I223651,I223677,I223685,I223285,I223716,I223294,I223747,I223764,I223306,I223795,I223297,I223288,I223291,I223309,I223895,I288538,I223921,I223929,I223946,I288514,I288529,I223963,I288541,I223989,I223997,I288526,I288517,I224023,I224031,I224048,I224065,I224082,I224122,I224130,I224147,I224164,I224181,I224212,I288532,I288523,I224229,I288535,I224255,I224263,I224294,I224325,I224342,I224373,I288520,I224473,I224499,I224507,I224524,I224541,I224567,I224575,I224601,I224609,I224626,I224643,I224660,I224700,I224708,I224725,I224742,I224759,I224790,I224807,I224833,I224841,I224872,I224903,I224920,I224951,I225051,I225077,I225085,I225102,I225119,I225145,I225153,I225179,I225187,I225204,I225221,I225238,I225034,I225278,I225286,I225303,I225320,I225337,I225037,I225368,I225385,I225411,I225419,I225019,I225450,I225028,I225481,I225498,I225040,I225529,I225031,I225022,I225025,I225043,I225629,I276264,I225655,I225663,I225680,I276240,I276255,I225697,I276267,I225723,I225731,I276252,I276243,I225757,I225765,I225782,I225799,I225816,I225612,I225856,I225864,I225881,I225898,I225915,I225615,I225946,I276258,I276249,I225963,I276261,I225989,I225997,I225597,I226028,I225606,I226059,I226076,I225618,I226107,I276246,I225609,I225600,I225603,I225621,I226207,I226233,I226241,I226258,I226275,I226301,I226309,I226335,I226343,I226360,I226377,I226394,I226434,I226442,I226459,I226476,I226493,I226524,I226541,I226567,I226575,I226606,I226637,I226654,I226685,I226785,I239756,I226811,I226819,I226836,I239744,I239762,I226853,I239759,I226879,I226887,I239750,I239747,I226913,I226921,I226938,I226955,I226972,I226768,I239741,I227012,I227020,I227037,I227054,I227071,I226771,I227102,I227119,I227145,I227153,I226753,I227184,I226762,I227215,I227232,I226774,I227263,I239753,I226765,I226756,I226759,I226777,I227363,I280140,I227389,I227397,I227414,I280116,I280131,I227431,I280143,I227457,I227465,I280128,I280119,I227491,I227499,I227516,I227533,I227550,I227346,I227590,I227598,I227615,I227632,I227649,I227349,I227680,I280134,I280125,I227697,I280137,I227723,I227731,I227331,I227762,I227340,I227793,I227810,I227352,I227841,I280122,I227343,I227334,I227337,I227355,I227941,I256093,I227967,I227975,I227992,I256081,I256099,I228009,I256096,I228035,I228043,I256087,I256084,I228069,I228077,I228094,I228111,I228128,I227924,I256078,I228168,I228176,I228193,I228210,I228227,I227927,I228258,I228275,I228301,I228309,I227909,I228340,I227918,I228371,I228388,I227930,I228419,I256090,I227921,I227912,I227915,I227933,I228519,I236594,I228545,I228553,I228570,I236582,I236600,I228587,I236597,I228613,I228621,I236588,I236585,I228647,I228655,I228672,I228689,I228706,I228502,I236579,I228746,I228754,I228771,I228788,I228805,I228505,I228836,I228853,I228879,I228887,I228487,I228918,I228496,I228949,I228966,I228508,I228997,I236591,I228499,I228490,I228493,I228511,I229097,I229123,I229131,I229148,I229165,I229191,I229199,I229225,I229233,I229250,I229267,I229284,I229080,I229324,I229332,I229349,I229366,I229383,I229083,I229414,I229431,I229457,I229465,I229065,I229496,I229074,I229527,I229544,I229086,I229575,I229077,I229068,I229071,I229089,I229675,I416466,I229701,I229709,I229726,I416451,I416439,I229743,I416454,I229769,I229777,I416457,I229803,I229811,I229828,I229845,I229862,I416445,I229902,I229910,I229927,I229944,I229961,I229992,I416442,I416448,I230009,I416463,I230035,I230043,I230074,I230105,I230122,I230153,I416460,I230253,I230279,I230287,I230304,I230321,I230347,I230355,I230381,I230389,I230406,I230423,I230440,I230236,I230480,I230488,I230505,I230522,I230539,I230239,I230570,I230587,I230613,I230621,I230221,I230652,I230230,I230683,I230700,I230242,I230731,I230233,I230224,I230227,I230245,I230831,I274326,I230857,I230865,I230882,I274302,I274317,I230899,I274329,I230925,I230933,I274314,I274305,I230959,I230967,I230984,I231001,I231018,I230814,I231058,I231066,I231083,I231100,I231117,I230817,I231148,I274320,I274311,I231165,I274323,I231191,I231199,I230799,I231230,I230808,I231261,I231278,I230820,I231309,I274308,I230811,I230802,I230805,I230823,I231409,I231435,I231443,I231460,I231477,I231503,I231511,I231537,I231545,I231562,I231579,I231596,I231636,I231644,I231661,I231678,I231695,I231726,I231743,I231769,I231777,I231808,I231839,I231856,I231887,I231987,I394014,I232013,I232021,I232038,I394002,I394020,I232055,I394011,I232081,I232089,I394026,I394023,I232115,I232123,I232140,I232157,I232174,I231970,I394005,I232214,I232222,I232239,I232256,I232273,I231973,I232304,I393999,I232321,I394008,I232347,I232355,I231955,I232386,I231964,I232417,I232434,I231976,I232465,I394017,I231967,I231958,I231961,I231979,I232565,I232591,I232599,I232616,I232633,I232659,I232667,I232693,I232701,I232718,I232735,I232752,I232792,I232800,I232817,I232834,I232851,I232882,I232899,I232925,I232933,I232964,I232995,I233012,I233043,I233143,I233169,I233177,I233194,I233211,I233237,I233245,I233271,I233279,I233296,I233313,I233330,I233126,I233370,I233378,I233395,I233412,I233429,I233129,I233460,I233477,I233503,I233511,I233111,I233542,I233120,I233573,I233590,I233132,I233621,I233123,I233114,I233117,I233135,I233721,I233747,I233755,I233772,I233789,I233815,I233823,I233849,I233857,I233874,I233891,I233908,I233948,I233956,I233973,I233990,I234007,I234038,I234055,I234081,I234089,I234120,I234151,I234168,I234199,I234299,I234325,I234333,I234350,I234367,I234393,I234401,I234427,I234435,I234452,I234469,I234486,I234282,I234526,I234534,I234551,I234568,I234585,I234285,I234616,I234633,I234659,I234667,I234267,I234698,I234276,I234729,I234746,I234288,I234777,I234279,I234270,I234273,I234291,I234877,I234903,I234911,I234928,I234945,I234971,I234979,I235005,I235013,I235030,I235047,I235064,I235104,I235112,I235129,I235146,I235163,I235194,I235211,I235237,I235245,I235276,I235307,I235324,I235355,I235455,I235481,I235489,I235506,I235523,I235549,I235557,I235583,I235591,I235608,I235625,I235642,I235438,I235682,I235690,I235707,I235724,I235741,I235441,I235772,I235789,I235815,I235823,I235423,I235854,I235432,I235885,I235902,I235444,I235933,I235435,I235426,I235429,I235447,I236033,I236059,I236067,I236084,I236101,I236127,I236135,I236161,I236169,I236186,I236203,I236220,I236260,I236268,I236285,I236302,I236319,I236350,I236367,I236393,I236401,I236432,I236463,I236480,I236511,I236608,I286579,I236634,I236642,I236659,I286594,I286576,I236676,I236702,I286585,I236733,I236741,I286603,I236758,I236784,I236792,I286600,I236832,I236868,I286597,I286588,I236885,I286582,I236911,I236919,I236936,I236967,I286591,I236984,I237001,I237032,I237063,I237080,I237135,I237161,I237169,I237186,I237203,I237229,I237260,I237268,I237285,I237311,I237319,I237359,I237395,I237412,I237438,I237446,I237463,I237494,I237511,I237528,I237559,I237590,I237607,I237662,I237688,I237696,I237713,I237730,I237756,I237787,I237795,I237812,I237838,I237846,I237886,I237922,I237939,I237965,I237973,I237990,I238021,I238038,I238055,I238086,I238117,I238134,I238189,I238215,I238223,I238240,I238257,I238283,I238178,I238314,I238322,I238339,I238365,I238373,I238181,I238413,I238172,I238163,I238449,I238466,I238492,I238500,I238517,I238166,I238548,I238565,I238582,I238175,I238613,I238160,I238644,I238661,I238169,I238716,I311524,I238742,I238750,I238767,I311533,I311521,I238784,I311518,I238810,I238841,I238849,I311515,I238866,I238892,I238900,I238940,I238976,I311536,I311527,I238993,I311530,I239019,I239027,I239044,I239075,I239092,I239109,I239140,I239171,I239188,I239243,I239269,I239277,I239294,I239311,I239337,I239368,I239376,I239393,I239419,I239427,I239467,I239503,I239520,I239546,I239554,I239571,I239602,I239619,I239636,I239667,I239698,I239715,I239770,I283349,I239796,I239804,I239821,I283364,I283346,I239838,I239864,I283355,I239895,I239903,I283373,I239920,I239946,I239954,I283370,I239994,I240030,I283367,I283358,I240047,I283352,I240073,I240081,I240098,I240129,I283361,I240146,I240163,I240194,I240225,I240242,I240297,I240323,I240331,I240348,I240365,I240391,I240422,I240430,I240447,I240473,I240481,I240521,I240557,I240574,I240600,I240608,I240625,I240656,I240673,I240690,I240721,I240752,I240769,I240824,I240850,I240858,I240875,I240892,I240918,I240813,I240949,I240957,I240974,I241000,I241008,I240816,I241048,I240807,I240798,I241084,I241101,I241127,I241135,I241152,I240801,I241183,I241200,I241217,I240810,I241248,I240795,I241279,I241296,I240804,I241351,I380757,I241377,I241385,I241402,I380739,I380742,I241419,I380754,I241445,I380763,I241476,I241484,I380748,I241501,I241527,I241535,I380760,I241575,I241611,I380751,I380745,I241628,I241654,I241662,I241679,I241710,I241727,I241744,I241775,I241806,I241823,I241878,I402769,I241904,I241912,I241929,I402766,I402775,I241946,I402754,I241972,I241867,I402757,I242003,I242011,I402772,I242028,I242054,I242062,I241870,I402778,I242102,I241861,I241852,I242138,I402760,I402781,I242155,I402763,I242181,I242189,I242206,I241855,I242237,I242254,I242271,I241864,I242302,I241849,I242333,I242350,I241858,I242405,I242431,I242439,I242456,I242473,I242499,I242394,I242530,I242538,I242555,I242581,I242589,I242397,I242629,I242388,I242379,I242665,I242682,I242708,I242716,I242733,I242382,I242764,I242781,I242798,I242391,I242829,I242376,I242860,I242877,I242385,I242932,I357977,I242958,I242966,I242983,I357959,I243000,I357965,I243026,I357962,I243057,I243065,I357971,I243082,I243108,I243116,I357983,I243156,I243192,I357974,I357968,I243209,I243235,I243243,I243260,I243291,I357980,I243308,I243325,I243356,I243387,I243404,I243459,I294331,I243485,I243493,I243510,I294346,I294328,I243527,I243553,I294337,I243584,I243592,I294355,I243609,I243635,I243643,I294352,I243683,I243719,I294349,I294340,I243736,I294334,I243762,I243770,I243787,I243818,I294343,I243835,I243852,I243883,I243914,I243931,I243986,I244012,I244020,I244037,I244054,I244080,I244111,I244119,I244136,I244162,I244170,I244210,I244246,I244263,I244289,I244297,I244314,I244345,I244362,I244379,I244410,I244441,I244458,I244513,I244539,I244547,I244564,I244581,I244607,I244638,I244646,I244663,I244689,I244697,I244737,I244773,I244790,I244816,I244824,I244841,I244872,I244889,I244906,I244937,I244968,I244985,I245040,I379601,I245066,I245074,I245091,I379583,I379586,I245108,I379598,I245134,I245029,I379607,I245165,I245173,I379592,I245190,I245216,I245224,I245032,I379604,I245264,I245023,I245014,I245300,I379595,I379589,I245317,I245343,I245351,I245368,I245017,I245399,I245416,I245433,I245026,I245464,I245011,I245495,I245512,I245020,I245567,I245593,I245601,I245618,I245635,I245661,I245556,I245692,I245700,I245717,I245743,I245751,I245559,I245791,I245550,I245541,I245827,I245844,I245870,I245878,I245895,I245544,I245926,I245943,I245960,I245553,I245991,I245538,I246022,I246039,I245547,I246094,I246120,I246128,I246145,I246162,I246188,I246219,I246227,I246244,I246270,I246278,I246318,I246354,I246371,I246397,I246405,I246422,I246453,I246470,I246487,I246518,I246549,I246566,I246621,I246647,I246655,I246672,I246689,I246715,I246746,I246754,I246771,I246797,I246805,I246845,I246881,I246898,I246924,I246932,I246949,I246980,I246997,I247014,I247045,I247076,I247093,I247148,I392883,I247174,I247182,I247199,I392877,I392895,I247216,I392880,I247242,I247137,I392901,I247273,I247281,I392886,I247298,I247324,I247332,I247140,I392898,I247372,I247131,I247122,I247408,I392889,I392904,I247425,I392892,I247451,I247459,I247476,I247125,I247507,I247524,I247541,I247134,I247572,I247119,I247603,I247620,I247128,I247675,I247701,I247709,I247726,I247743,I247769,I247664,I247800,I247808,I247825,I247851,I247859,I247667,I247899,I247658,I247649,I247935,I247952,I247978,I247986,I248003,I247652,I248034,I248051,I248068,I247661,I248099,I247646,I248130,I248147,I247655,I248202,I353931,I248228,I248236,I248253,I353913,I248270,I353919,I248296,I353916,I248327,I248335,I353925,I248352,I248378,I248386,I353937,I248426,I248462,I353928,I353922,I248479,I248505,I248513,I248530,I248561,I353934,I248578,I248595,I248626,I248657,I248674,I248729,I379023,I248755,I248763,I248780,I379005,I379008,I248797,I379020,I248823,I379029,I248854,I248862,I379014,I248879,I248905,I248913,I379026,I248953,I248989,I379017,I379011,I249006,I249032,I249040,I249057,I249088,I249105,I249122,I249153,I249184,I249201,I249256,I249282,I249290,I249307,I249324,I249350,I249381,I249389,I249406,I249432,I249440,I249480,I249516,I249533,I249559,I249567,I249584,I249615,I249632,I249649,I249680,I249711,I249728,I249783,I249809,I249817,I249834,I249851,I249877,I249908,I249916,I249933,I249959,I249967,I250007,I250043,I250060,I250086,I250094,I250111,I250142,I250159,I250176,I250207,I250238,I250255,I250310,I250336,I250344,I250361,I250378,I250404,I250435,I250443,I250460,I250486,I250494,I250534,I250570,I250587,I250613,I250621,I250638,I250669,I250686,I250703,I250734,I250765,I250782,I250837,I250863,I250871,I250888,I250905,I250931,I250962,I250970,I250987,I251013,I251021,I251061,I251097,I251114,I251140,I251148,I251165,I251196,I251213,I251230,I251261,I251292,I251309,I251364,I251390,I251398,I251415,I251432,I251458,I251489,I251497,I251514,I251540,I251548,I251588,I251624,I251641,I251667,I251675,I251692,I251723,I251740,I251757,I251788,I251819,I251836,I251891,I406339,I251917,I251925,I251942,I406336,I406345,I251959,I406324,I251985,I406327,I252016,I252024,I406342,I252041,I252067,I252075,I406348,I252115,I252151,I406330,I406351,I252168,I406333,I252194,I252202,I252219,I252250,I252267,I252284,I252315,I252346,I252363,I252418,I252444,I252452,I252469,I252486,I252512,I252407,I252543,I252551,I252568,I252594,I252602,I252410,I252642,I252401,I252392,I252678,I252695,I252721,I252729,I252746,I252395,I252777,I252794,I252811,I252404,I252842,I252389,I252873,I252890,I252398,I252945,I384803,I252971,I252979,I252996,I384785,I384788,I253013,I384800,I253039,I384809,I253070,I253078,I384794,I253095,I253121,I253129,I384806,I253169,I253205,I384797,I384791,I253222,I253248,I253256,I253273,I253304,I253321,I253338,I253369,I253400,I253417,I253472,I253498,I253506,I253523,I253540,I253566,I253461,I253597,I253605,I253622,I253648,I253656,I253464,I253696,I253455,I253446,I253732,I253749,I253775,I253783,I253800,I253449,I253831,I253848,I253865,I253458,I253896,I253443,I253927,I253944,I253452,I253999,I254025,I254033,I254050,I254067,I254093,I254124,I254132,I254149,I254175,I254183,I254223,I254259,I254276,I254302,I254310,I254327,I254358,I254375,I254392,I254423,I254454,I254471,I254526,I254552,I254560,I254577,I254594,I254620,I254515,I254651,I254659,I254676,I254702,I254710,I254518,I254750,I254509,I254500,I254786,I254803,I254829,I254837,I254854,I254503,I254885,I254902,I254919,I254512,I254950,I254497,I254981,I254998,I254506,I255053,I366505,I255079,I255087,I255104,I366511,I366493,I255121,I366502,I255147,I366508,I255178,I255186,I366496,I255203,I255229,I255237,I366514,I255277,I255313,I366499,I255330,I366517,I255356,I255364,I255381,I255412,I255429,I255446,I255477,I255508,I255525,I255580,I331389,I255606,I255614,I255631,I331371,I255648,I331377,I255674,I255569,I331374,I255705,I255713,I331383,I255730,I255756,I255764,I255572,I331395,I255804,I255563,I255554,I255840,I331386,I331380,I255857,I255883,I255891,I255908,I255557,I255939,I331392,I255956,I255973,I255566,I256004,I255551,I256035,I256052,I255560,I256107,I256133,I256141,I256158,I256175,I256201,I256232,I256240,I256257,I256283,I256291,I256331,I256367,I256384,I256410,I256418,I256435,I256466,I256483,I256500,I256531,I256562,I256579,I256634,I338903,I256660,I256668,I256685,I338885,I256702,I338891,I256728,I338888,I256759,I256767,I338897,I256784,I256810,I256818,I338909,I256858,I256894,I338900,I338894,I256911,I256937,I256945,I256962,I256993,I338906,I257010,I257027,I257058,I257089,I257106,I257161,I257187,I257195,I257212,I257229,I257255,I257286,I257294,I257311,I257337,I257345,I257385,I257421,I257438,I257464,I257472,I257489,I257520,I257537,I257554,I257585,I257616,I257633,I257688,I296269,I257714,I257722,I257739,I296284,I296266,I257756,I257782,I257677,I296275,I257813,I257821,I296293,I257838,I257864,I257872,I257680,I296290,I257912,I257671,I257662,I257948,I296287,I296278,I257965,I296272,I257991,I257999,I258016,I257665,I258047,I296281,I258064,I258081,I257674,I258112,I257659,I258143,I258160,I257668,I258215,I258241,I258249,I258266,I258283,I258309,I258340,I258348,I258365,I258391,I258399,I258439,I258475,I258492,I258518,I258526,I258543,I258574,I258591,I258608,I258639,I258670,I258687,I258742,I258768,I258776,I258793,I258810,I258836,I258867,I258875,I258892,I258918,I258926,I258966,I259002,I259019,I259045,I259053,I259070,I259101,I259118,I259135,I259166,I259197,I259214,I259269,I259295,I259303,I259320,I259337,I259363,I259258,I259394,I259402,I259419,I259445,I259453,I259261,I259493,I259252,I259243,I259529,I259546,I259572,I259580,I259597,I259246,I259628,I259645,I259662,I259255,I259693,I259240,I259724,I259741,I259249,I259796,I343527,I259822,I259830,I259847,I343509,I259864,I343515,I259890,I343512,I259921,I259929,I343521,I259946,I259972,I259980,I343533,I260020,I260056,I343524,I343518,I260073,I260099,I260107,I260124,I260155,I343530,I260172,I260189,I260220,I260251,I260268,I260323,I260349,I260357,I260374,I260391,I260417,I260448,I260456,I260473,I260499,I260507,I260547,I260583,I260600,I260626,I260634,I260651,I260682,I260699,I260716,I260747,I260778,I260795,I260850,I260876,I260884,I260901,I260918,I260944,I260975,I260983,I261000,I261026,I261034,I261074,I261110,I261127,I261153,I261161,I261178,I261209,I261226,I261243,I261274,I261305,I261322,I261377,I261403,I261411,I261428,I261445,I261471,I261366,I261502,I261510,I261527,I261553,I261561,I261369,I261601,I261360,I261351,I261637,I261654,I261680,I261688,I261705,I261354,I261736,I261753,I261770,I261363,I261801,I261348,I261832,I261849,I261357,I261904,I261930,I261938,I261955,I261972,I261998,I262029,I262037,I262054,I262080,I262088,I262128,I262164,I262181,I262207,I262215,I262232,I262263,I262280,I262297,I262328,I262359,I262376,I262431,I262457,I262465,I262482,I262499,I262525,I262420,I262556,I262564,I262581,I262607,I262615,I262423,I262655,I262414,I262405,I262691,I262708,I262734,I262742,I262759,I262408,I262790,I262807,I262824,I262417,I262855,I262402,I262886,I262903,I262411,I262958,I381335,I262984,I262992,I263009,I381317,I381320,I263026,I381332,I263052,I262947,I381341,I263083,I263091,I381326,I263108,I263134,I263142,I262950,I381338,I263182,I262941,I262932,I263218,I381329,I381323,I263235,I263261,I263269,I263286,I262935,I263317,I263334,I263351,I262944,I263382,I262929,I263413,I263430,I262938,I263485,I263511,I263519,I263536,I263553,I263579,I263610,I263618,I263635,I263661,I263669,I263709,I263745,I263762,I263788,I263796,I263813,I263844,I263861,I263878,I263909,I263940,I263957,I264012,I264038,I264046,I264063,I264080,I264106,I264137,I264145,I264162,I264188,I264196,I264236,I264272,I264289,I264315,I264323,I264340,I264371,I264388,I264405,I264436,I264467,I264484,I264539,I264565,I264573,I264590,I264607,I264633,I264528,I264664,I264672,I264689,I264715,I264723,I264531,I264763,I264522,I264513,I264799,I264816,I264842,I264850,I264867,I264516,I264898,I264915,I264932,I264525,I264963,I264510,I264994,I265011,I264519,I265066,I265092,I265100,I265117,I265134,I265160,I265191,I265199,I265216,I265242,I265250,I265290,I265326,I265343,I265369,I265377,I265394,I265425,I265442,I265459,I265490,I265521,I265538,I265593,I265619,I265627,I265644,I265661,I265687,I265718,I265726,I265743,I265769,I265777,I265817,I265853,I265870,I265896,I265904,I265921,I265952,I265969,I265986,I266017,I266048,I266065,I266120,I336013,I266146,I266154,I266171,I335995,I266188,I336001,I266214,I335998,I266245,I266253,I336007,I266270,I266296,I266304,I336019,I266344,I266380,I336010,I336004,I266397,I266423,I266431,I266448,I266479,I336016,I266496,I266513,I266544,I266575,I266592,I266647,I266673,I266681,I266698,I266715,I266741,I266772,I266780,I266797,I266823,I266831,I266871,I266907,I266924,I266950,I266958,I266975,I267006,I267023,I267040,I267071,I267102,I267119,I267174,I267200,I267208,I267225,I267242,I267268,I267299,I267307,I267324,I267350,I267358,I267398,I267434,I267451,I267477,I267485,I267502,I267533,I267550,I267567,I267598,I267629,I267646,I267701,I267727,I267735,I267752,I267769,I267795,I267826,I267834,I267851,I267877,I267885,I267925,I267961,I267978,I268004,I268012,I268029,I268060,I268077,I268094,I268125,I268156,I268173,I268228,I268254,I268262,I268279,I268296,I268322,I268353,I268361,I268378,I268404,I268412,I268452,I268488,I268505,I268531,I268539,I268556,I268587,I268604,I268621,I268652,I268683,I268700,I268755,I268781,I268789,I268806,I268823,I268849,I268880,I268888,I268905,I268931,I268939,I268979,I269015,I269032,I269058,I269066,I269083,I269114,I269131,I269148,I269179,I269210,I269227,I269282,I269308,I269316,I269333,I269350,I269376,I269407,I269415,I269432,I269458,I269466,I269506,I269542,I269559,I269585,I269593,I269610,I269641,I269658,I269675,I269706,I269737,I269754,I269815,I269841,I269858,I269866,I269883,I269900,I269917,I269934,I269951,I269982,I269999,I270030,I270047,I270064,I270095,I270135,I270143,I270160,I270177,I270194,I270225,I270242,I270259,I270285,I270307,I270324,I270355,I270400,I270461,I270487,I270504,I270512,I270529,I270546,I270563,I270580,I270597,I270447,I270628,I270645,I270450,I270676,I270693,I270710,I270426,I270741,I270438,I270781,I270789,I270806,I270823,I270840,I270453,I270871,I270888,I270905,I270931,I270441,I270953,I270970,I270435,I271001,I270429,I270432,I271046,I270444,I271107,I271133,I271150,I271158,I271175,I271192,I271209,I271226,I271243,I271274,I271291,I271322,I271339,I271356,I271387,I271427,I271435,I271452,I271469,I271486,I271517,I271534,I271551,I271577,I271599,I271616,I271647,I271692,I271753,I271779,I271796,I271804,I271821,I271838,I271855,I271872,I271889,I271739,I271920,I271937,I271742,I271968,I271985,I272002,I271718,I272033,I271730,I272073,I272081,I272098,I272115,I272132,I271745,I272163,I272180,I272197,I272223,I271733,I272245,I272262,I271727,I272293,I271721,I271724,I272338,I271736,I272399,I272425,I272442,I272450,I272467,I272484,I272501,I272518,I272535,I272566,I272583,I272614,I272631,I272648,I272679,I272719,I272727,I272744,I272761,I272778,I272809,I272826,I272843,I272869,I272891,I272908,I272939,I272984,I273045,I334279,I273071,I334261,I273088,I273096,I273113,I334270,I273130,I334282,I273147,I334264,I273164,I334273,I273181,I273212,I273229,I273260,I273277,I334285,I273294,I273325,I273365,I273373,I273390,I273407,I273424,I273455,I334267,I273472,I334276,I273489,I273515,I273537,I273554,I273585,I273630,I273691,I273717,I273734,I273742,I273759,I273776,I273793,I273810,I273827,I273677,I273858,I273875,I273680,I273906,I273923,I273940,I273656,I273971,I273668,I274011,I274019,I274036,I274053,I274070,I273683,I274101,I274118,I274135,I274161,I273671,I274183,I274200,I273665,I274231,I273659,I273662,I274276,I273674,I274337,I274363,I274380,I274388,I274405,I274422,I274439,I274456,I274473,I274504,I274521,I274552,I274569,I274586,I274617,I274657,I274665,I274682,I274699,I274716,I274747,I274764,I274781,I274807,I274829,I274846,I274877,I274922,I274983,I275009,I275026,I275034,I275051,I275068,I275085,I275102,I275119,I275150,I275167,I275198,I275215,I275232,I275263,I275303,I275311,I275328,I275345,I275362,I275393,I275410,I275427,I275453,I275475,I275492,I275523,I275568,I275629,I403944,I275655,I403968,I275672,I275680,I275697,I403950,I275714,I403959,I275731,I275748,I403965,I275765,I275615,I275796,I275813,I275618,I275844,I275861,I403962,I275878,I275594,I275909,I275606,I275949,I275957,I275974,I275991,I403956,I276008,I275621,I276039,I403947,I276056,I403971,I276073,I403953,I276099,I275609,I276121,I276138,I275603,I276169,I275597,I275600,I276214,I275612,I276275,I276301,I276318,I276326,I276343,I276360,I276377,I276394,I276411,I276442,I276459,I276490,I276507,I276524,I276555,I276595,I276603,I276620,I276637,I276654,I276685,I276702,I276719,I276745,I276767,I276784,I276815,I276860,I276921,I276947,I276964,I276972,I276989,I277006,I277023,I277040,I277057,I276907,I277088,I277105,I276910,I277136,I277153,I277170,I276886,I277201,I276898,I277241,I277249,I277266,I277283,I277300,I276913,I277331,I277348,I277365,I277391,I276901,I277413,I277430,I276895,I277461,I276889,I276892,I277506,I276904,I277567,I277593,I277610,I277618,I277635,I277652,I277669,I277686,I277703,I277553,I277734,I277751,I277556,I277782,I277799,I277816,I277532,I277847,I277544,I277887,I277895,I277912,I277929,I277946,I277559,I277977,I277994,I278011,I278037,I277547,I278059,I278076,I277541,I278107,I277535,I277538,I278152,I277550,I278213,I278239,I278256,I278264,I278281,I278298,I278315,I278332,I278349,I278199,I278380,I278397,I278202,I278428,I278445,I278462,I278178,I278493,I278190,I278533,I278541,I278558,I278575,I278592,I278205,I278623,I278640,I278657,I278683,I278193,I278705,I278722,I278187,I278753,I278181,I278184,I278798,I278196,I278859,I278885,I278902,I278910,I278927,I278944,I278961,I278978,I278995,I279026,I279043,I279074,I279091,I279108,I279139,I279179,I279187,I279204,I279221,I279238,I279269,I279286,I279303,I279329,I279351,I279368,I279399,I279444,I279505,I279531,I279548,I279556,I279573,I279590,I279607,I279624,I279641,I279672,I279689,I279720,I279737,I279754,I279785,I279825,I279833,I279850,I279867,I279884,I279915,I279932,I279949,I279975,I279997,I280014,I280045,I280090,I280151,I280177,I280194,I280202,I280219,I280236,I280253,I280270,I280287,I280318,I280335,I280366,I280383,I280400,I280431,I280471,I280479,I280496,I280513,I280530,I280561,I280578,I280595,I280621,I280643,I280660,I280691,I280736,I280797,I378479,I280823,I378485,I280840,I280848,I280865,I378482,I280882,I378461,I280899,I378464,I280916,I378470,I280933,I280783,I280964,I280981,I280786,I281012,I281029,I281046,I280762,I281077,I280774,I281117,I281125,I281142,I281159,I378473,I281176,I280789,I281207,I281224,I378467,I281241,I378476,I281267,I280777,I281289,I281306,I280771,I281337,I280765,I280768,I281382,I280780,I281443,I281469,I281486,I281494,I281511,I281528,I281545,I281562,I281579,I281610,I281627,I281658,I281675,I281692,I281723,I281763,I281771,I281788,I281805,I281822,I281853,I281870,I281887,I281913,I281935,I281952,I281983,I282028,I282089,I282115,I282132,I282140,I282157,I282174,I282191,I282208,I282225,I282256,I282273,I282304,I282321,I282338,I282369,I282409,I282417,I282434,I282451,I282468,I282499,I282516,I282533,I282559,I282581,I282598,I282629,I282674,I282735,I282761,I282778,I282786,I282803,I282820,I282837,I282854,I282871,I282902,I282919,I282950,I282967,I282984,I283015,I283055,I283063,I283080,I283097,I283114,I283145,I283162,I283179,I283205,I283227,I283244,I283275,I283320,I283381,I283407,I283424,I283432,I283449,I283466,I283483,I283500,I283517,I283548,I283565,I283596,I283613,I283630,I283661,I283701,I283709,I283726,I283743,I283760,I283791,I283808,I283825,I283851,I283873,I283890,I283921,I283966,I284027,I368143,I284053,I368149,I284070,I284078,I284095,I368146,I284112,I368125,I284129,I368128,I284146,I368134,I284163,I284013,I284194,I284211,I284016,I284242,I284259,I284276,I283992,I284307,I284004,I284347,I284355,I284372,I284389,I368137,I284406,I284019,I284437,I284454,I368131,I284471,I368140,I284497,I284007,I284519,I284536,I284001,I284567,I283995,I283998,I284612,I284010,I284673,I284699,I284716,I284724,I284741,I284758,I284775,I284792,I284809,I284840,I284857,I284888,I284905,I284922,I284953,I284993,I285001,I285018,I285035,I285052,I285083,I285100,I285117,I285143,I285165,I285182,I285213,I285258,I285319,I285345,I285362,I285370,I285387,I285404,I285421,I285438,I285455,I285486,I285503,I285534,I285551,I285568,I285599,I285639,I285647,I285664,I285681,I285698,I285729,I285746,I285763,I285789,I285811,I285828,I285859,I285904,I285965,I317686,I285991,I317689,I286008,I286016,I286033,I286050,I317698,I286067,I317707,I286084,I317695,I286101,I286132,I286149,I286180,I286197,I317701,I286214,I286245,I286285,I286293,I286310,I286327,I317692,I286344,I286375,I317704,I286392,I286409,I286435,I286457,I286474,I286505,I286550,I286611,I286637,I286654,I286662,I286679,I286696,I286713,I286730,I286747,I286778,I286795,I286826,I286843,I286860,I286891,I286931,I286939,I286956,I286973,I286990,I287021,I287038,I287055,I287081,I287103,I287120,I287151,I287196,I287257,I287283,I287300,I287308,I287325,I287342,I287359,I287376,I287393,I287424,I287441,I287472,I287489,I287506,I287537,I287577,I287585,I287602,I287619,I287636,I287667,I287684,I287701,I287727,I287749,I287766,I287797,I287842,I287903,I346417,I287929,I346399,I287946,I287954,I287971,I346408,I287988,I346420,I288005,I346402,I288022,I346411,I288039,I288070,I288087,I288118,I288135,I346423,I288152,I288183,I288223,I288231,I288248,I288265,I288282,I288313,I346405,I288330,I346414,I288347,I288373,I288395,I288412,I288443,I288488,I288549,I288575,I288592,I288600,I288617,I288634,I288651,I288668,I288685,I288716,I288733,I288764,I288781,I288798,I288829,I288869,I288877,I288894,I288911,I288928,I288959,I288976,I288993,I289019,I289041,I289058,I289089,I289134,I289195,I289221,I289238,I289246,I289263,I289280,I289297,I289314,I289331,I289181,I289362,I289379,I289184,I289410,I289427,I289444,I289160,I289475,I289172,I289515,I289523,I289540,I289557,I289574,I289187,I289605,I289622,I289639,I289665,I289175,I289687,I289704,I289169,I289735,I289163,I289166,I289780,I289178,I289841,I289867,I289884,I289892,I289909,I289926,I289943,I289960,I289977,I289827,I290008,I290025,I289830,I290056,I290073,I290090,I289806,I290121,I289818,I290161,I290169,I290186,I290203,I290220,I289833,I290251,I290268,I290285,I290311,I289821,I290333,I290350,I289815,I290381,I289809,I289812,I290426,I289824,I290487,I395697,I290513,I395694,I290530,I290538,I290555,I395691,I290572,I395682,I290589,I395703,I290606,I290623,I290654,I290671,I290702,I290719,I395706,I290736,I290767,I290807,I290815,I290832,I290849,I395685,I290866,I290897,I395688,I290914,I395709,I290931,I395700,I290957,I290979,I290996,I291027,I291072,I291133,I291159,I291176,I291184,I291201,I291218,I291235,I291252,I291269,I291119,I291300,I291317,I291122,I291348,I291365,I291382,I291098,I291413,I291110,I291453,I291461,I291478,I291495,I291512,I291125,I291543,I291560,I291577,I291603,I291113,I291625,I291642,I291107,I291673,I291101,I291104,I291718,I291116,I291779,I291805,I291822,I291830,I291847,I291864,I291881,I291898,I291915,I291946,I291963,I291994,I292011,I292028,I292059,I292099,I292107,I292124,I292141,I292158,I292189,I292206,I292223,I292249,I292271,I292288,I292319,I292364,I292425,I292451,I292468,I292476,I292493,I292510,I292527,I292544,I292561,I292592,I292609,I292640,I292657,I292674,I292705,I292745,I292753,I292770,I292787,I292804,I292835,I292852,I292869,I292895,I292917,I292934,I292965,I293010,I293071,I293097,I293114,I293122,I293139,I293156,I293173,I293190,I293207,I293238,I293255,I293286,I293303,I293320,I293351,I293391,I293399,I293416,I293433,I293450,I293481,I293498,I293515,I293541,I293563,I293580,I293611,I293656,I293717,I293743,I293760,I293768,I293785,I293802,I293819,I293836,I293853,I293703,I293884,I293901,I293706,I293932,I293949,I293966,I293682,I293997,I293694,I294037,I294045,I294062,I294079,I294096,I293709,I294127,I294144,I294161,I294187,I293697,I294209,I294226,I293691,I294257,I293685,I293688,I294302,I293700,I294363,I341793,I294389,I341775,I294406,I294414,I294431,I341784,I294448,I341796,I294465,I341778,I294482,I341787,I294499,I294530,I294547,I294578,I294595,I341799,I294612,I294643,I294683,I294691,I294708,I294725,I294742,I294773,I341781,I294790,I341790,I294807,I294833,I294855,I294872,I294903,I294948,I295009,I319930,I295035,I319933,I295052,I295060,I295077,I295094,I319942,I295111,I319951,I295128,I319939,I295145,I295176,I295193,I295224,I295241,I319945,I295258,I295289,I295329,I295337,I295354,I295371,I319936,I295388,I295419,I319948,I295436,I295453,I295479,I295501,I295518,I295549,I295594,I295655,I295681,I295698,I295706,I295723,I295740,I295757,I295774,I295791,I295641,I295822,I295839,I295644,I295870,I295887,I295904,I295620,I295935,I295632,I295975,I295983,I296000,I296017,I296034,I295647,I296065,I296082,I296099,I296125,I295635,I296147,I296164,I295629,I296195,I295623,I295626,I296240,I295638,I296301,I296327,I296344,I296352,I296369,I296386,I296403,I296420,I296437,I296468,I296485,I296516,I296533,I296550,I296581,I296621,I296629,I296646,I296663,I296680,I296711,I296728,I296745,I296771,I296793,I296810,I296841,I296886,I296947,I296973,I296990,I296998,I297015,I297032,I297049,I297066,I297083,I297114,I297131,I297162,I297179,I297196,I297227,I297267,I297275,I297292,I297309,I297326,I297357,I297374,I297391,I297417,I297439,I297456,I297487,I297532,I297593,I334857,I297619,I334839,I297636,I297644,I297661,I334848,I297678,I334860,I297695,I334842,I297712,I334851,I297729,I297579,I297760,I297777,I297582,I297808,I297825,I334863,I297842,I297558,I297873,I297570,I297913,I297921,I297938,I297955,I297972,I297585,I298003,I334845,I298020,I334854,I298037,I298063,I297573,I298085,I298102,I297567,I298133,I297561,I297564,I298178,I297576,I298239,I320491,I298265,I320494,I298282,I298290,I298307,I298324,I320503,I298341,I320512,I298358,I320500,I298375,I298406,I298423,I298454,I298471,I320506,I298488,I298519,I298559,I298567,I298584,I298601,I320497,I298618,I298649,I320509,I298666,I298683,I298709,I298731,I298748,I298779,I298824,I298885,I400374,I298911,I400398,I298928,I298936,I298953,I400380,I298970,I400389,I298987,I299004,I400395,I299021,I298871,I299052,I299069,I298874,I299100,I299117,I400392,I299134,I298850,I299165,I298862,I299205,I299213,I299230,I299247,I400386,I299264,I298877,I299295,I400377,I299312,I400401,I299329,I400383,I299355,I298865,I299377,I299394,I298859,I299425,I298853,I298856,I299470,I298868,I299531,I299557,I299574,I299582,I299599,I299616,I299633,I299650,I299667,I299698,I299715,I299746,I299763,I299780,I299811,I299851,I299859,I299876,I299893,I299910,I299941,I299958,I299975,I300001,I300023,I300040,I300071,I300116,I300177,I300203,I300220,I300228,I300245,I300262,I300279,I300296,I300313,I300344,I300361,I300392,I300409,I300426,I300457,I300497,I300505,I300522,I300539,I300556,I300587,I300604,I300621,I300647,I300669,I300686,I300717,I300762,I300823,I300849,I300866,I300874,I300891,I300908,I300925,I300942,I300959,I300990,I301007,I301038,I301055,I301072,I301103,I301143,I301151,I301168,I301185,I301202,I301233,I301250,I301267,I301293,I301315,I301332,I301363,I301408,I301469,I391152,I301495,I391146,I301512,I301520,I301537,I391155,I301554,I391167,I301571,I391149,I301588,I301605,I301455,I301636,I301653,I301458,I301684,I301701,I391143,I301718,I301434,I301749,I301446,I301789,I301797,I301814,I301831,I391164,I301848,I301461,I301879,I391158,I301896,I301913,I391161,I301939,I301449,I301961,I301978,I301443,I302009,I301437,I301440,I302054,I301452,I302115,I310954,I302141,I310957,I302158,I302166,I302183,I302200,I310966,I302217,I310975,I302234,I310963,I302251,I302282,I302299,I302330,I302347,I310969,I302364,I302395,I302435,I302443,I302460,I302477,I310960,I302494,I302525,I310972,I302542,I302559,I302585,I302607,I302624,I302655,I302700,I302761,I302787,I302804,I302812,I302829,I302846,I302863,I302880,I302897,I302747,I302928,I302945,I302750,I302976,I302993,I303010,I302726,I303041,I302738,I303081,I303089,I303106,I303123,I303140,I302753,I303171,I303188,I303205,I303231,I302741,I303253,I303270,I302735,I303301,I302729,I302732,I303346,I302744,I303407,I369231,I303433,I369237,I303450,I303458,I303475,I369234,I303492,I369213,I303509,I369216,I303526,I369222,I303543,I303574,I303591,I303622,I303639,I303656,I303687,I303727,I303735,I303752,I303769,I369225,I303786,I303817,I303834,I369219,I303851,I369228,I303877,I303899,I303916,I303947,I303992,I304053,I304079,I304096,I304104,I304121,I304138,I304155,I304172,I304189,I304220,I304237,I304268,I304285,I304302,I304333,I304373,I304381,I304398,I304415,I304432,I304463,I304480,I304497,I304523,I304545,I304562,I304593,I304638,I304699,I304725,I304742,I304750,I304767,I304784,I304801,I304818,I304835,I304866,I304883,I304914,I304931,I304948,I304979,I305019,I305027,I305044,I305061,I305078,I305109,I305126,I305143,I305169,I305191,I305208,I305239,I305284,I305345,I365423,I305371,I365429,I305388,I305396,I305413,I365426,I305430,I365405,I305447,I365408,I305464,I365414,I305481,I305512,I305529,I305560,I305577,I305594,I305625,I305665,I305673,I305690,I305707,I365417,I305724,I305755,I305772,I365411,I305789,I365420,I305815,I305837,I305854,I305885,I305930,I305991,I306017,I306034,I306042,I306059,I306076,I306093,I306110,I306127,I305977,I306158,I306175,I305980,I306206,I306223,I306240,I305956,I306271,I305968,I306311,I306319,I306336,I306353,I306370,I305983,I306401,I306418,I306435,I306461,I305971,I306483,I306500,I305965,I306531,I305959,I305962,I306576,I305974,I306637,I350463,I306663,I350445,I306680,I306688,I306705,I350454,I306722,I350466,I306739,I350448,I306756,I350457,I306773,I306623,I306804,I306821,I306626,I306852,I306869,I350469,I306886,I306602,I306917,I306614,I306957,I306965,I306982,I306999,I307016,I306629,I307047,I350451,I307064,I350460,I307081,I307107,I306617,I307129,I307146,I306611,I307177,I306605,I306608,I307222,I306620,I307283,I377391,I307309,I377397,I307326,I307334,I307351,I377394,I307368,I377373,I307385,I377376,I307402,I377382,I307419,I307450,I307467,I307498,I307515,I307532,I307563,I307603,I307611,I307628,I307645,I377385,I307662,I307693,I307710,I377379,I307727,I377388,I307753,I307775,I307792,I307823,I307868,I307929,I307955,I307972,I307980,I307997,I308014,I308031,I308048,I308065,I308096,I308113,I308144,I308161,I308178,I308209,I308249,I308257,I308274,I308291,I308308,I308339,I308356,I308373,I308399,I308421,I308438,I308469,I308514,I308575,I308601,I308618,I308626,I308643,I308660,I308677,I308694,I308711,I308742,I308759,I308790,I308807,I308824,I308855,I308895,I308903,I308920,I308937,I308954,I308985,I309002,I309019,I309045,I309067,I309084,I309115,I309160,I309221,I309247,I309264,I309272,I309289,I309306,I309323,I309340,I309357,I309388,I309405,I309436,I309453,I309470,I309501,I309541,I309549,I309566,I309583,I309600,I309631,I309648,I309665,I309691,I309713,I309730,I309761,I309806,I309861,I309887,I309904,I309853,I309926,I309952,I309960,I309977,I309994,I310011,I310028,I310045,I310062,I309835,I310093,I309838,I310124,I310141,I310158,I310175,I309847,I310206,I309850,I309844,I310251,I310268,I310285,I310311,I310319,I309832,I310350,I310367,I309841,I310422,I417644,I310448,I310465,I310487,I417638,I310513,I310521,I417629,I310538,I310555,I417656,I310572,I417641,I417650,I310589,I310606,I417635,I310623,I310654,I310685,I417653,I310702,I310719,I310736,I310767,I310812,I417647,I310829,I310846,I417632,I310872,I310880,I310911,I310928,I310983,I311009,I311026,I311048,I311074,I311082,I311099,I311116,I311133,I311150,I311167,I311184,I311215,I311246,I311263,I311280,I311297,I311328,I311373,I311390,I311407,I311433,I311441,I311472,I311489,I311544,I311570,I311587,I311609,I311635,I311643,I311660,I311677,I311694,I311711,I311728,I311745,I311776,I311807,I311824,I311841,I311858,I311889,I311934,I311951,I311968,I311994,I312002,I312033,I312050,I312105,I312131,I312148,I312097,I312170,I312196,I312204,I312221,I312238,I312255,I312272,I312289,I312306,I312079,I312337,I312082,I312368,I312385,I312402,I312419,I312091,I312450,I312094,I312088,I312495,I312512,I312529,I312555,I312563,I312076,I312594,I312611,I312085,I312666,I312692,I312709,I312731,I312757,I312765,I312782,I312799,I312816,I312833,I312850,I312867,I312898,I312929,I312946,I312963,I312980,I313011,I313056,I313073,I313090,I313116,I313124,I313155,I313172,I313227,I365955,I313253,I313270,I313292,I365961,I313318,I313326,I365970,I313343,I313360,I365949,I313377,I365952,I313394,I313411,I365964,I313428,I313459,I313490,I365958,I313507,I313524,I313541,I313572,I313617,I365973,I313634,I313651,I365967,I313677,I313685,I313716,I313733,I313788,I313814,I313831,I313853,I313879,I313887,I313904,I313921,I313938,I313955,I313972,I313989,I314020,I314051,I314068,I314085,I314102,I314133,I314178,I314195,I314212,I314238,I314246,I314277,I314294,I314349,I314375,I314392,I314414,I314440,I314448,I314465,I314482,I314499,I314516,I314533,I314550,I314581,I314612,I314629,I314646,I314663,I314694,I314739,I314756,I314773,I314799,I314807,I314838,I314855,I314910,I314936,I314953,I314975,I315001,I315009,I315026,I315043,I315060,I315077,I315094,I315111,I315142,I315173,I315190,I315207,I315224,I315255,I315300,I315317,I315334,I315360,I315368,I315399,I315416,I315471,I315497,I315514,I315536,I315562,I315570,I315587,I315604,I315621,I315638,I315655,I315672,I315703,I315734,I315751,I315768,I315785,I315816,I315861,I315878,I315895,I315921,I315929,I315960,I315977,I316032,I316058,I316075,I316097,I316123,I316131,I316148,I316165,I316182,I316199,I316216,I316233,I316264,I316295,I316312,I316329,I316346,I316377,I316422,I316439,I316456,I316482,I316490,I316521,I316538,I316593,I413479,I316619,I316636,I316658,I413473,I316684,I316692,I413464,I316709,I316726,I413491,I316743,I413476,I413485,I316760,I316777,I413470,I316794,I316825,I316856,I413488,I316873,I316890,I316907,I316938,I316983,I413482,I317000,I317017,I413467,I317043,I317051,I317082,I317099,I317154,I317180,I317197,I317146,I317219,I317245,I317253,I317270,I317287,I317304,I317321,I317338,I317355,I317128,I317386,I317131,I317417,I317434,I317451,I317468,I317140,I317499,I317143,I317137,I317544,I317561,I317578,I317604,I317612,I317125,I317643,I317660,I317134,I317715,I317741,I317758,I317780,I317806,I317814,I317831,I317848,I317865,I317882,I317899,I317916,I317947,I317978,I317995,I318012,I318029,I318060,I318105,I318122,I318139,I318165,I318173,I318204,I318221,I318276,I327340,I318302,I318319,I318268,I318341,I327331,I318367,I318375,I327328,I318392,I318409,I327337,I318426,I327346,I318443,I318460,I327325,I318477,I318250,I318508,I318253,I318539,I327334,I318556,I318573,I318590,I318262,I318621,I318265,I318259,I318666,I327349,I318683,I318700,I327343,I318726,I318734,I318247,I318765,I318782,I318256,I318837,I341212,I318863,I318880,I318902,I341203,I318928,I318936,I341200,I318953,I318970,I341209,I318987,I341218,I319004,I319021,I341197,I319038,I319069,I319100,I341206,I319117,I319134,I319151,I319182,I319227,I341221,I319244,I319261,I341215,I319287,I319295,I319326,I319343,I319398,I319424,I319441,I319390,I319463,I319489,I319497,I319514,I319531,I319548,I319565,I319582,I319599,I319372,I319630,I319375,I319661,I319678,I319695,I319712,I319384,I319743,I319387,I319381,I319788,I319805,I319822,I319848,I319856,I319369,I319887,I319904,I319378,I319959,I319985,I320002,I320024,I320050,I320058,I320075,I320092,I320109,I320126,I320143,I320160,I320191,I320222,I320239,I320256,I320273,I320304,I320349,I320366,I320383,I320409,I320417,I320448,I320465,I320520,I351616,I320546,I320563,I320585,I351607,I320611,I320619,I351604,I320636,I320653,I351613,I320670,I351622,I320687,I320704,I351601,I320721,I320752,I320783,I351610,I320800,I320817,I320834,I320865,I320910,I351625,I320927,I320944,I351619,I320970,I320978,I321009,I321026,I321081,I321107,I321124,I321146,I321172,I321180,I321197,I321214,I321231,I321248,I321265,I321282,I321313,I321344,I321361,I321378,I321395,I321426,I321471,I321488,I321505,I321531,I321539,I321570,I321587,I321642,I321668,I321685,I321707,I321733,I321741,I321758,I321775,I321792,I321809,I321826,I321843,I321874,I321905,I321922,I321939,I321956,I321987,I322032,I322049,I322066,I322092,I322100,I322131,I322148,I322203,I322229,I322246,I322195,I322268,I322294,I322302,I322319,I322336,I322353,I322370,I322387,I322404,I322177,I322435,I322180,I322466,I322483,I322500,I322517,I322189,I322548,I322192,I322186,I322593,I322610,I322627,I322653,I322661,I322174,I322692,I322709,I322183,I322764,I322790,I322807,I322829,I322855,I322863,I322880,I322897,I322914,I322931,I322948,I322965,I322996,I323027,I323044,I323061,I323078,I323109,I323154,I323171,I323188,I323214,I323222,I323253,I323270,I323325,I340056,I323351,I323368,I323390,I340047,I323416,I323424,I340044,I323441,I323458,I340053,I323475,I340062,I323492,I323509,I340041,I323526,I323557,I323588,I340050,I323605,I323622,I323639,I323670,I323715,I340065,I323732,I323749,I340059,I323775,I323783,I323814,I323831,I323889,I323915,I323923,I323963,I323971,I323988,I324005,I324045,I324067,I324084,I324110,I324118,I324135,I324152,I324169,I324186,I324231,I324262,I324279,I324305,I324313,I324344,I324361,I324378,I324395,I324467,I324493,I324501,I324541,I324549,I324566,I324583,I324623,I324645,I324662,I324688,I324696,I324713,I324730,I324747,I324764,I324809,I324840,I324857,I324883,I324891,I324922,I324939,I324956,I324973,I325045,I325071,I325079,I325119,I325127,I325144,I325161,I325201,I325223,I325240,I325266,I325274,I325291,I325308,I325325,I325342,I325387,I325418,I325435,I325461,I325469,I325500,I325517,I325534,I325551,I325623,I393438,I325649,I325657,I393465,I393447,I325697,I325705,I393456,I325722,I393459,I325739,I325779,I325801,I393453,I325818,I325844,I325852,I325869,I393441,I325886,I393444,I325903,I325920,I325965,I393462,I325996,I326013,I393450,I326039,I326047,I326078,I326095,I326112,I326129,I326201,I326227,I326235,I326184,I326275,I326283,I326300,I326317,I326172,I326357,I326193,I326379,I326396,I326422,I326430,I326447,I326464,I326481,I326498,I326169,I326190,I326543,I326181,I326574,I326591,I326617,I326625,I326187,I326656,I326673,I326690,I326707,I326178,I326175,I326779,I326805,I326813,I326853,I326861,I326878,I326895,I326935,I326957,I326974,I327000,I327008,I327025,I327042,I327059,I327076,I327121,I327152,I327169,I327195,I327203,I327234,I327251,I327268,I327285,I327357,I327383,I327391,I327431,I327439,I327456,I327473,I327513,I327535,I327552,I327578,I327586,I327603,I327620,I327637,I327654,I327699,I327730,I327747,I327773,I327781,I327812,I327829,I327846,I327863,I327935,I327961,I327969,I328009,I328017,I328034,I328051,I328091,I328113,I328130,I328156,I328164,I328181,I328198,I328215,I328232,I328277,I328308,I328325,I328351,I328359,I328390,I328407,I328424,I328441,I328513,I328539,I328547,I328496,I328587,I328595,I328612,I328629,I328484,I328669,I328505,I328691,I328708,I328734,I328742,I328759,I328776,I328793,I328810,I328481,I328502,I328855,I328493,I328886,I328903,I328929,I328937,I328499,I328968,I328985,I329002,I329019,I328490,I328487,I329091,I329117,I329125,I329165,I329173,I329190,I329207,I329247,I329269,I329286,I329312,I329320,I329337,I329354,I329371,I329388,I329433,I329464,I329481,I329507,I329515,I329546,I329563,I329580,I329597,I329669,I390589,I329695,I329703,I390571,I390580,I329743,I329751,I390565,I329768,I390577,I329785,I329825,I329847,I390568,I329864,I329890,I329898,I329915,I329932,I329949,I329966,I330011,I390586,I330042,I330059,I390574,I390583,I330085,I330093,I330124,I330141,I330158,I330175,I330247,I330273,I330281,I330321,I330329,I330346,I330363,I330403,I330425,I330442,I330468,I330476,I330493,I330510,I330527,I330544,I330589,I330620,I330637,I330663,I330671,I330702,I330719,I330736,I330753,I330825,I330851,I330859,I330899,I330907,I330924,I330941,I330981,I331003,I331020,I331046,I331054,I331071,I331088,I331105,I331122,I331167,I331198,I331215,I331241,I331249,I331280,I331297,I331314,I331331,I331403,I331429,I331437,I331477,I331485,I331502,I331519,I331559,I331581,I331598,I331624,I331632,I331649,I331666,I331683,I331700,I331745,I331776,I331793,I331819,I331827,I331858,I331875,I331892,I331909,I331981,I332007,I332015,I331964,I332055,I332063,I332080,I332097,I331952,I332137,I331973,I332159,I332176,I332202,I332210,I332227,I332244,I332261,I332278,I331949,I331970,I332323,I331961,I332354,I332371,I332397,I332405,I331967,I332436,I332453,I332470,I332487,I331958,I331955,I332559,I332585,I332593,I332633,I332641,I332658,I332675,I332715,I332737,I332754,I332780,I332788,I332805,I332822,I332839,I332856,I332901,I332932,I332949,I332975,I332983,I333014,I333031,I333048,I333065,I333137,I333163,I333171,I333211,I333219,I333236,I333253,I333293,I333315,I333332,I333358,I333366,I333383,I333400,I333417,I333434,I333479,I333510,I333527,I333553,I333561,I333592,I333609,I333626,I333643,I333715,I333741,I333749,I333789,I333797,I333814,I333831,I333871,I333893,I333910,I333936,I333944,I333961,I333978,I333995,I334012,I334057,I334088,I334105,I334131,I334139,I334170,I334187,I334204,I334221,I334293,I334319,I334327,I334367,I334375,I334392,I334409,I334449,I334471,I334488,I334514,I334522,I334539,I334556,I334573,I334590,I334635,I334666,I334683,I334709,I334717,I334748,I334765,I334782,I334799,I334871,I334897,I334905,I334945,I334953,I334970,I334987,I335027,I335049,I335066,I335092,I335100,I335117,I335134,I335151,I335168,I335213,I335244,I335261,I335287,I335295,I335326,I335343,I335360,I335377,I335449,I335475,I335483,I335523,I335531,I335548,I335565,I335605,I335627,I335644,I335670,I335678,I335695,I335712,I335729,I335746,I335791,I335822,I335839,I335865,I335873,I335904,I335921,I335938,I335955,I336027,I394560,I336053,I336061,I394587,I394569,I336101,I336109,I394578,I336126,I394581,I336143,I336183,I336205,I394575,I336222,I336248,I336256,I336273,I394563,I336290,I394566,I336307,I336324,I336369,I394584,I336400,I336417,I394572,I336443,I336451,I336482,I336499,I336516,I336533,I336605,I336631,I336639,I336588,I336679,I336687,I336704,I336721,I336576,I336761,I336597,I336783,I336800,I336826,I336834,I336851,I336868,I336885,I336902,I336573,I336594,I336947,I336585,I336978,I336995,I337021,I337029,I336591,I337060,I337077,I337094,I337111,I336582,I336579,I337183,I337209,I337217,I337257,I337265,I337282,I337299,I337339,I337361,I337378,I337404,I337412,I337429,I337446,I337463,I337480,I337525,I337556,I337573,I337599,I337607,I337638,I337655,I337672,I337689,I337761,I387121,I337787,I337795,I387103,I387112,I337835,I337843,I387097,I337860,I387109,I337877,I337917,I337939,I387100,I337956,I337982,I337990,I338007,I338024,I338041,I338058,I338103,I387118,I338134,I338151,I387106,I387115,I338177,I338185,I338216,I338233,I338250,I338267,I338339,I338365,I338373,I338322,I338413,I338421,I338438,I338455,I338310,I338495,I338331,I338517,I338534,I338560,I338568,I338585,I338602,I338619,I338636,I338307,I338328,I338681,I338319,I338712,I338729,I338755,I338763,I338325,I338794,I338811,I338828,I338845,I338316,I338313,I338917,I338943,I338951,I338991,I338999,I339016,I339033,I339073,I339095,I339112,I339138,I339146,I339163,I339180,I339197,I339214,I339259,I339290,I339307,I339333,I339341,I339372,I339389,I339406,I339423,I339495,I339521,I339529,I339569,I339577,I339594,I339611,I339651,I339673,I339690,I339716,I339724,I339741,I339758,I339775,I339792,I339837,I339868,I339885,I339911,I339919,I339950,I339967,I339984,I340001,I340073,I375762,I340099,I340107,I375756,I375741,I340147,I340155,I375747,I340172,I375759,I340189,I340229,I340251,I340268,I340294,I340302,I340319,I375765,I340336,I375753,I340353,I340370,I340415,I375744,I340446,I340463,I375750,I340489,I340497,I340528,I340545,I340562,I340579,I340651,I340677,I340685,I340634,I340725,I340733,I340750,I340767,I340622,I340807,I340643,I340829,I340846,I340872,I340880,I340897,I340914,I340931,I340948,I340619,I340640,I340993,I340631,I341024,I341041,I341067,I341075,I340637,I341106,I341123,I341140,I341157,I340628,I340625,I341229,I341255,I341263,I341303,I341311,I341328,I341345,I341385,I341407,I341424,I341450,I341458,I341475,I341492,I341509,I341526,I341571,I341602,I341619,I341645,I341653,I341684,I341701,I341718,I341735,I341807,I341833,I341841,I341881,I341889,I341906,I341923,I341963,I341985,I342002,I342028,I342036,I342053,I342070,I342087,I342104,I342149,I342180,I342197,I342223,I342231,I342262,I342279,I342296,I342313,I342385,I396243,I342411,I342419,I396270,I342368,I396252,I342459,I342467,I396261,I342484,I396264,I342501,I342356,I342541,I342377,I342563,I396258,I342580,I342606,I342614,I342631,I396246,I342648,I396249,I342665,I342682,I342353,I342374,I342727,I396267,I342365,I342758,I342775,I396255,I342801,I342809,I342371,I342840,I342857,I342874,I342891,I342362,I342359,I342963,I418846,I342989,I342997,I418828,I418819,I343037,I343045,I418834,I343062,I418822,I343079,I343119,I343141,I418831,I343158,I343184,I343192,I343209,I418840,I343226,I343243,I343260,I343305,I418843,I343336,I343353,I418837,I418825,I343379,I343387,I343418,I343435,I343452,I343469,I343541,I417061,I343567,I343575,I417043,I417034,I343615,I343623,I417049,I343640,I417037,I343657,I343697,I343719,I417046,I343736,I343762,I343770,I343787,I417055,I343804,I343821,I343838,I343883,I417058,I343914,I343931,I417052,I417040,I343957,I343965,I343996,I344013,I344030,I344047,I344119,I344145,I344153,I344102,I344193,I344201,I344218,I344235,I344090,I344275,I344111,I344297,I344314,I344340,I344348,I344365,I344382,I344399,I344416,I344087,I344108,I344461,I344099,I344492,I344509,I344535,I344543,I344105,I344574,I344591,I344608,I344625,I344096,I344093,I344697,I389433,I344723,I344731,I389415,I389424,I344771,I344779,I389409,I344796,I389421,I344813,I344853,I344875,I389412,I344892,I344918,I344926,I344943,I344960,I344977,I344994,I345039,I389430,I345070,I345087,I389418,I389427,I345113,I345121,I345152,I345169,I345186,I345203,I345275,I345301,I345309,I345258,I345349,I345357,I345374,I345391,I345246,I345431,I345267,I345453,I345470,I345496,I345504,I345521,I345538,I345555,I345572,I345243,I345264,I345617,I345255,I345648,I345665,I345691,I345699,I345261,I345730,I345747,I345764,I345781,I345252,I345249,I345853,I345879,I345887,I345927,I345935,I345952,I345969,I346009,I346031,I346048,I346074,I346082,I346099,I346116,I346133,I346150,I346195,I346226,I346243,I346269,I346277,I346308,I346325,I346342,I346359,I346431,I346457,I346465,I346505,I346513,I346530,I346547,I346587,I346609,I346626,I346652,I346660,I346677,I346694,I346711,I346728,I346773,I346804,I346821,I346847,I346855,I346886,I346903,I346920,I346937,I347009,I412896,I347035,I347043,I412878,I412869,I347083,I347091,I412884,I347108,I412872,I347125,I347165,I347187,I412881,I347204,I347230,I347238,I347255,I412890,I347272,I347289,I347306,I347351,I412893,I347382,I347399,I412887,I412875,I347425,I347433,I347464,I347481,I347498,I347515,I347587,I398021,I347613,I347621,I398003,I397994,I347661,I347669,I398009,I347686,I397997,I347703,I347743,I347765,I398006,I347782,I347808,I347816,I347833,I398015,I347850,I347867,I347884,I347929,I398018,I347960,I347977,I398012,I398000,I348003,I348011,I348042,I348059,I348076,I348093,I348165,I348191,I348199,I348239,I348247,I348264,I348281,I348321,I348343,I348360,I348386,I348394,I348411,I348428,I348445,I348462,I348507,I348538,I348555,I348581,I348589,I348620,I348637,I348654,I348671,I348743,I348769,I348777,I348726,I348817,I348825,I348842,I348859,I348714,I348899,I348735,I348921,I348938,I348964,I348972,I348989,I349006,I349023,I349040,I348711,I348732,I349085,I348723,I349116,I349133,I349159,I349167,I348729,I349198,I349215,I349232,I349249,I348720,I348717,I349321,I349347,I349355,I349395,I349403,I349420,I349437,I349477,I349499,I349516,I349542,I349550,I349567,I349584,I349601,I349618,I349663,I349694,I349711,I349737,I349745,I349776,I349793,I349810,I349827,I349899,I349925,I349933,I349882,I349973,I349981,I349998,I350015,I349870,I350055,I349891,I350077,I350094,I350120,I350128,I350145,I350162,I350179,I350196,I349867,I349888,I350241,I349879,I350272,I350289,I350315,I350323,I349885,I350354,I350371,I350388,I350405,I349876,I349873,I350477,I350503,I350511,I350551,I350559,I350576,I350593,I350633,I350655,I350672,I350698,I350706,I350723,I350740,I350757,I350774,I350819,I350850,I350867,I350893,I350901,I350932,I350949,I350966,I350983,I351055,I351081,I351089,I351129,I351137,I351154,I351171,I351211,I351233,I351250,I351276,I351284,I351301,I351318,I351335,I351352,I351397,I351428,I351445,I351471,I351479,I351510,I351527,I351544,I351561,I351633,I351659,I351667,I351707,I351715,I351732,I351749,I351789,I351811,I351828,I351854,I351862,I351879,I351896,I351913,I351930,I351975,I352006,I352023,I352049,I352057,I352088,I352105,I352122,I352139,I352211,I352237,I352245,I352285,I352293,I352310,I352327,I352367,I352389,I352406,I352432,I352440,I352457,I352474,I352491,I352508,I352553,I352584,I352601,I352627,I352635,I352666,I352683,I352700,I352717,I352789,I380185,I352815,I352823,I380167,I380176,I352863,I352871,I380161,I352888,I380173,I352905,I352945,I352967,I380164,I352984,I353010,I353018,I353035,I353052,I353069,I353086,I353131,I380182,I353162,I353179,I380170,I380179,I353205,I353213,I353244,I353261,I353278,I353295,I353367,I353393,I353401,I353441,I353449,I353466,I353483,I353523,I353545,I353562,I353588,I353596,I353613,I353630,I353647,I353664,I353709,I353740,I353757,I353783,I353791,I353822,I353839,I353856,I353873,I353945,I353971,I353979,I354019,I354027,I354044,I354061,I354101,I354123,I354140,I354166,I354174,I354191,I354208,I354225,I354242,I354287,I354318,I354335,I354361,I354369,I354400,I354417,I354434,I354451,I354523,I354549,I354557,I354597,I354605,I354622,I354639,I354679,I354701,I354718,I354744,I354752,I354769,I354786,I354803,I354820,I354865,I354896,I354913,I354939,I354947,I354978,I354995,I355012,I355029,I355101,I355127,I355135,I355175,I355183,I355200,I355217,I355257,I355279,I355296,I355322,I355330,I355347,I355364,I355381,I355398,I355443,I355474,I355491,I355517,I355525,I355556,I355573,I355590,I355607,I355679,I355705,I355713,I355753,I355761,I355778,I355795,I355835,I355857,I355874,I355900,I355908,I355925,I355942,I355959,I355976,I356021,I356052,I356069,I356095,I356103,I356134,I356151,I356168,I356185,I356257,I397426,I356283,I356291,I397408,I397399,I356331,I356339,I397414,I356356,I397402,I356373,I356413,I356435,I397411,I356452,I356478,I356486,I356503,I397420,I356520,I356537,I356554,I356599,I397423,I356630,I356647,I397417,I397405,I356673,I356681,I356712,I356729,I356746,I356763,I356835,I408731,I356861,I356869,I408713,I356818,I408704,I356909,I356917,I408719,I356934,I408707,I356951,I356806,I356991,I356827,I357013,I408716,I357030,I357056,I357064,I357081,I408725,I357098,I357115,I357132,I356803,I356824,I357177,I408728,I356815,I357208,I357225,I408722,I408710,I357251,I357259,I356821,I357290,I357307,I357324,I357341,I356812,I356809,I357413,I404566,I357439,I357447,I404548,I404539,I357487,I357495,I404554,I357512,I404542,I357529,I357569,I357591,I404551,I357608,I357634,I357642,I357659,I404560,I357676,I357693,I357710,I357755,I404563,I357786,I357803,I404557,I404545,I357829,I357837,I357868,I357885,I357902,I357919,I357991,I358017,I358025,I358065,I358073,I358090,I358107,I358147,I358169,I358186,I358212,I358220,I358237,I358254,I358271,I358288,I358333,I358364,I358381,I358407,I358415,I358446,I358463,I358480,I358497,I358569,I358595,I358603,I358643,I358651,I358668,I358685,I358725,I358747,I358764,I358790,I358798,I358815,I358832,I358849,I358866,I358911,I358942,I358959,I358985,I358993,I359024,I359041,I359058,I359075,I359147,I359173,I359181,I359221,I359229,I359246,I359263,I359303,I359325,I359342,I359368,I359376,I359393,I359410,I359427,I359444,I359489,I359520,I359537,I359563,I359571,I359602,I359619,I359636,I359653,I359725,I383653,I359751,I359759,I383635,I383644,I359799,I359807,I383629,I359824,I383641,I359841,I359881,I359903,I383632,I359920,I359946,I359954,I359971,I359988,I360005,I360022,I360067,I383650,I360098,I360115,I383638,I383647,I360141,I360149,I360180,I360197,I360214,I360231,I360303,I360329,I360337,I360377,I360385,I360402,I360419,I360459,I360481,I360498,I360524,I360532,I360549,I360566,I360583,I360600,I360645,I360676,I360693,I360719,I360727,I360758,I360775,I360792,I360809,I360881,I360907,I360915,I360955,I360963,I360980,I360997,I361037,I361059,I361076,I361102,I361110,I361127,I361144,I361161,I361178,I361223,I361254,I361271,I361297,I361305,I361336,I361353,I361370,I361387,I361459,I361485,I361493,I361533,I361541,I361558,I361575,I361615,I361637,I361654,I361680,I361688,I361705,I361722,I361739,I361756,I361801,I361832,I361849,I361875,I361883,I361914,I361931,I361948,I361965,I362037,I362063,I362071,I362111,I362119,I362136,I362153,I362193,I362215,I362232,I362258,I362266,I362283,I362300,I362317,I362334,I362379,I362410,I362427,I362453,I362461,I362492,I362509,I362526,I362543,I362615,I377938,I362641,I362649,I377932,I377917,I362689,I362697,I377923,I362714,I377935,I362731,I362771,I362793,I362810,I362836,I362844,I362861,I377941,I362878,I377929,I362895,I362912,I362957,I377920,I362988,I363005,I377926,I363031,I363039,I363070,I363087,I363104,I363121,I363193,I401591,I363219,I363227,I401573,I401564,I363267,I363275,I401579,I363292,I401567,I363309,I363349,I363371,I401576,I363388,I363414,I363422,I363439,I401585,I363456,I363473,I363490,I363535,I401588,I363566,I363583,I401582,I401570,I363609,I363617,I363648,I363665,I363682,I363699,I363771,I363797,I363805,I363845,I363853,I363870,I363887,I363927,I363949,I363966,I363992,I364000,I364017,I364034,I364051,I364068,I364113,I364144,I364161,I364187,I364195,I364226,I364243,I364260,I364277,I364349,I364375,I364383,I364409,I364426,I364448,I364465,I364482,I364499,I364516,I364547,I364564,I364581,I364598,I364643,I364660,I364677,I364736,I364762,I364770,I364787,I364804,I364835,I364893,I364919,I364927,I364953,I364970,I364992,I365009,I365026,I365043,I365060,I365091,I365108,I365125,I365142,I365187,I365204,I365221,I365280,I365306,I365314,I365331,I365348,I365379,I365437,I365463,I365471,I365497,I365514,I365536,I365553,I365570,I365587,I365604,I365635,I365652,I365669,I365686,I365731,I365748,I365765,I365824,I365850,I365858,I365875,I365892,I365923,I365981,I366007,I366015,I366041,I366058,I366080,I366097,I366114,I366131,I366148,I366179,I366196,I366213,I366230,I366275,I366292,I366309,I366368,I366394,I366402,I366419,I366436,I366467,I366525,I366551,I366559,I366585,I366602,I366624,I366641,I366658,I366675,I366692,I366723,I366740,I366757,I366774,I366819,I366836,I366853,I366912,I366938,I366946,I366963,I366980,I367011,I367069,I367095,I367103,I367129,I367146,I367061,I367168,I367185,I367202,I367219,I367236,I367040,I367267,I367284,I367301,I367318,I367043,I367058,I367363,I367380,I367397,I367055,I367052,I367049,I367456,I367482,I367490,I367507,I367524,I367037,I367555,I367046,I367613,I367639,I367647,I367673,I367690,I367712,I367729,I367746,I367763,I367780,I367811,I367828,I367845,I367862,I367907,I367924,I367941,I368000,I368026,I368034,I368051,I368068,I368099,I368157,I368183,I368191,I368217,I368234,I368256,I368273,I368290,I368307,I368324,I368355,I368372,I368389,I368406,I368451,I368468,I368485,I368544,I368570,I368578,I368595,I368612,I368643,I368701,I368727,I368735,I368761,I368778,I368800,I368817,I368834,I368851,I368868,I368899,I368916,I368933,I368950,I368995,I369012,I369029,I369088,I369114,I369122,I369139,I369156,I369187,I369245,I369271,I369279,I369305,I369322,I369344,I369361,I369378,I369395,I369412,I369443,I369460,I369477,I369494,I369539,I369556,I369573,I369632,I369658,I369666,I369683,I369700,I369731,I369789,I369815,I369823,I369849,I369866,I369888,I369905,I369922,I369939,I369956,I369987,I370004,I370021,I370038,I370083,I370100,I370117,I370176,I370202,I370210,I370227,I370244,I370275,I370333,I370359,I370367,I370393,I370410,I370432,I370449,I370466,I370483,I370500,I370531,I370548,I370565,I370582,I370627,I370644,I370661,I370720,I370746,I370754,I370771,I370788,I370819,I370877,I370903,I370911,I370937,I370954,I370976,I370993,I371010,I371027,I371044,I371075,I371092,I371109,I371126,I371171,I371188,I371205,I371264,I371290,I371298,I371315,I371332,I371363,I371421,I371447,I371455,I371481,I371498,I371520,I371537,I371554,I371571,I371588,I371619,I371636,I371653,I371670,I371715,I371732,I371749,I371808,I371834,I371842,I371859,I371876,I371907,I371965,I371991,I371999,I372025,I372042,I372064,I372081,I372098,I372115,I372132,I372163,I372180,I372197,I372214,I372259,I372276,I372293,I372352,I372378,I372386,I372403,I372420,I372451,I372509,I372535,I372543,I372569,I372586,I372608,I372625,I372642,I372659,I372676,I372707,I372724,I372741,I372758,I372803,I372820,I372837,I372896,I372922,I372930,I372947,I372964,I372995,I373053,I373079,I373087,I373113,I373130,I373152,I373169,I373186,I373203,I373220,I373251,I373268,I373285,I373302,I373347,I373364,I373381,I373440,I373466,I373474,I373491,I373508,I373539,I373597,I373623,I373631,I373657,I373674,I373589,I373696,I373713,I373730,I373747,I373764,I373568,I373795,I373812,I373829,I373846,I373571,I373586,I373891,I373908,I373925,I373583,I373580,I373577,I373984,I374010,I374018,I374035,I374052,I373565,I374083,I373574,I374141,I374167,I374175,I374201,I374218,I374240,I374257,I374274,I374291,I374308,I374339,I374356,I374373,I374390,I374435,I374452,I374469,I374528,I374554,I374562,I374579,I374596,I374627,I374685,I374711,I374719,I374745,I374762,I374677,I374784,I374801,I374818,I374835,I374852,I374656,I374883,I374900,I374917,I374934,I374659,I374674,I374979,I374996,I375013,I374671,I374668,I374665,I375072,I375098,I375106,I375123,I375140,I374653,I375171,I374662,I375229,I375255,I375263,I375289,I375306,I375328,I375345,I375362,I375379,I375396,I375427,I375444,I375461,I375478,I375523,I375540,I375557,I375616,I375642,I375650,I375667,I375684,I375715,I375773,I375799,I375807,I375833,I375850,I375872,I375889,I375906,I375923,I375940,I375971,I375988,I376005,I376022,I376067,I376084,I376101,I376160,I376186,I376194,I376211,I376228,I376259,I376317,I376343,I376351,I376377,I376394,I376416,I376433,I376450,I376467,I376484,I376515,I376532,I376549,I376566,I376611,I376628,I376645,I376704,I376730,I376738,I376755,I376772,I376803,I376861,I376887,I376895,I376921,I376938,I376960,I376977,I376994,I377011,I377028,I377059,I377076,I377093,I377110,I377155,I377172,I377189,I377248,I377274,I377282,I377299,I377316,I377347,I377405,I377431,I377439,I377465,I377482,I377504,I377521,I377538,I377555,I377572,I377603,I377620,I377637,I377654,I377699,I377716,I377733,I377792,I377818,I377826,I377843,I377860,I377891,I377949,I377975,I377983,I378009,I378026,I378048,I378065,I378082,I378099,I378116,I378147,I378164,I378181,I378198,I378243,I378260,I378277,I378336,I378362,I378370,I378387,I378404,I378435,I378493,I378519,I378527,I378553,I378570,I378592,I378609,I378626,I378643,I378660,I378691,I378708,I378725,I378742,I378787,I378804,I378821,I378880,I378906,I378914,I378931,I378948,I378979,I379037,I379063,I379071,I379088,I379114,I379122,I379139,I379156,I379173,I379190,I379221,I379238,I379255,I379286,I379303,I379343,I379351,I379382,I379399,I379416,I379433,I379464,I379495,I379521,I379543,I379615,I379641,I379649,I379666,I379692,I379700,I379717,I379734,I379751,I379768,I379799,I379816,I379833,I379864,I379881,I379921,I379929,I379960,I379977,I379994,I380011,I380042,I380073,I380099,I380121,I380193,I395139,I380219,I380227,I395133,I380244,I395148,I380270,I380278,I380295,I395124,I380312,I395121,I380329,I380346,I395127,I380377,I380394,I395136,I380411,I380442,I395130,I380459,I380499,I380507,I380538,I395145,I380555,I380572,I380589,I380620,I380651,I395142,I380677,I380699,I380771,I380797,I380805,I380822,I380848,I380856,I380873,I380890,I380907,I380924,I380955,I380972,I380989,I381020,I381037,I381077,I381085,I381116,I381133,I381150,I381167,I381198,I381229,I381255,I381277,I381349,I381375,I381383,I381400,I381426,I381434,I381451,I381468,I381485,I381502,I381533,I381550,I381567,I381598,I381615,I381655,I381663,I381694,I381711,I381728,I381745,I381776,I381807,I381833,I381855,I381927,I381953,I381961,I381978,I382004,I382012,I382029,I382046,I382063,I382080,I382111,I382128,I382145,I382176,I382193,I382233,I382241,I382272,I382289,I382306,I382323,I382354,I382385,I382411,I382433,I382505,I382531,I382539,I382556,I382582,I382590,I382607,I382624,I382641,I382658,I382689,I382706,I382723,I382754,I382771,I382811,I382819,I382850,I382867,I382884,I382901,I382932,I382963,I382989,I383011,I383083,I383109,I383117,I383134,I383160,I383168,I383185,I383202,I383219,I383236,I383267,I383284,I383301,I383332,I383349,I383389,I383397,I383428,I383445,I383462,I383479,I383510,I383541,I383567,I383589,I383661,I383687,I383695,I383712,I383738,I383746,I383763,I383780,I383797,I383814,I383845,I383862,I383879,I383910,I383927,I383967,I383975,I384006,I384023,I384040,I384057,I384088,I384119,I384145,I384167,I384239,I384265,I384273,I384290,I384316,I384324,I384341,I384358,I384375,I384392,I384423,I384440,I384457,I384488,I384505,I384545,I384553,I384584,I384601,I384618,I384635,I384666,I384697,I384723,I384745,I384817,I384843,I384851,I384868,I384894,I384902,I384919,I384936,I384953,I384970,I385001,I385018,I385035,I385066,I385083,I385123,I385131,I385162,I385179,I385196,I385213,I385244,I385275,I385301,I385323,I385395,I385421,I385429,I385446,I385472,I385480,I385497,I385514,I385531,I385548,I385579,I385596,I385613,I385644,I385661,I385701,I385709,I385740,I385757,I385774,I385791,I385822,I385853,I385879,I385901,I385973,I411703,I385999,I386007,I411694,I386024,I411679,I386050,I386058,I386075,I411682,I386092,I411691,I386109,I386126,I411688,I386157,I411700,I386174,I386191,I386222,I411685,I386239,I386279,I386287,I386318,I411706,I386335,I386352,I386369,I386400,I386431,I411697,I386457,I386479,I386551,I386577,I386585,I386602,I386628,I386636,I386653,I386670,I386687,I386704,I386735,I386752,I386769,I386800,I386817,I386857,I386865,I386896,I386913,I386930,I386947,I386978,I387009,I387035,I387057,I387129,I387155,I387163,I387180,I387206,I387214,I387231,I387248,I387265,I387282,I387313,I387330,I387347,I387378,I387395,I387435,I387443,I387474,I387491,I387508,I387525,I387556,I387587,I387613,I387635,I387707,I387733,I387741,I387758,I387784,I387792,I387809,I387826,I387843,I387860,I387891,I387908,I387925,I387956,I387973,I388013,I388021,I388052,I388069,I388086,I388103,I388134,I388165,I388191,I388213,I388285,I388311,I388319,I388336,I388362,I388370,I388387,I388404,I388421,I388438,I388469,I388486,I388503,I388534,I388551,I388591,I388599,I388630,I388647,I388664,I388681,I388712,I388743,I388769,I388791,I388863,I388889,I388897,I388914,I388940,I388948,I388965,I388982,I388999,I389016,I389047,I389064,I389081,I389112,I389129,I389169,I389177,I389208,I389225,I389242,I389259,I389290,I389321,I389347,I389369,I389441,I389467,I389475,I389492,I389518,I389526,I389543,I389560,I389577,I389594,I389625,I389642,I389659,I389690,I389707,I389747,I389755,I389786,I389803,I389820,I389837,I389868,I389899,I389925,I389947,I390019,I390045,I390053,I390070,I390096,I390104,I390121,I390138,I390155,I390172,I390203,I390220,I390237,I390268,I390285,I390325,I390333,I390364,I390381,I390398,I390415,I390446,I390477,I390503,I390525,I390597,I390623,I390631,I390648,I390674,I390682,I390699,I390716,I390733,I390750,I390781,I390798,I390815,I390846,I390863,I390903,I390911,I390942,I390959,I390976,I390993,I391024,I391055,I391081,I391103,I391175,I391201,I391209,I391226,I391252,I391260,I391277,I391294,I391311,I391328,I391359,I391376,I391393,I391424,I391441,I391481,I391489,I391520,I391537,I391554,I391571,I391602,I391633,I391659,I391681,I391753,I391779,I391787,I391804,I391830,I391838,I391855,I391872,I391889,I391906,I391937,I391954,I391971,I392002,I392019,I392059,I392067,I392098,I392115,I392132,I392149,I392180,I392211,I392237,I392259,I392331,I392357,I392365,I392382,I392408,I392416,I392433,I392450,I392467,I392484,I392515,I392532,I392549,I392580,I392597,I392637,I392645,I392676,I392693,I392710,I392727,I392758,I392789,I392815,I392837,I392912,I392938,I392946,I392963,I392989,I392997,I393014,I393031,I393062,I393093,I393110,I393127,I393144,I393161,I393192,I393251,I393268,I393294,I393316,I393342,I393350,I393367,I393398,I393473,I393499,I393507,I393524,I393550,I393558,I393575,I393592,I393623,I393654,I393671,I393688,I393705,I393722,I393753,I393812,I393829,I393855,I393877,I393903,I393911,I393928,I393959,I394034,I394060,I394068,I394085,I394111,I394119,I394136,I394153,I394184,I394215,I394232,I394249,I394266,I394283,I394314,I394373,I394390,I394416,I394438,I394464,I394472,I394489,I394520,I394595,I394621,I394629,I394646,I394672,I394680,I394697,I394714,I394745,I394776,I394793,I394810,I394827,I394844,I394875,I394934,I394951,I394977,I394999,I395025,I395033,I395050,I395081,I395156,I395182,I395190,I395207,I395233,I395241,I395258,I395275,I395306,I395337,I395354,I395371,I395388,I395405,I395436,I395495,I395512,I395538,I395560,I395586,I395594,I395611,I395642,I395717,I395743,I395751,I395768,I395794,I395802,I395819,I395836,I395867,I395898,I395915,I395932,I395949,I395966,I395997,I396056,I396073,I396099,I396121,I396147,I396155,I396172,I396203,I396278,I396304,I396312,I396329,I396355,I396363,I396380,I396397,I396428,I396459,I396476,I396493,I396510,I396527,I396558,I396617,I396634,I396660,I396682,I396708,I396716,I396733,I396764,I396839,I396865,I396882,I396890,I396935,I396952,I396969,I396986,I397003,I397020,I397037,I397068,I397085,I397130,I397147,I397164,I397195,I397221,I397229,I397260,I397277,I397294,I397320,I397328,I397345,I397434,I397460,I397477,I397485,I397530,I397547,I397564,I397581,I397598,I397615,I397632,I397663,I397680,I397725,I397742,I397759,I397790,I397816,I397824,I397855,I397872,I397889,I397915,I397923,I397940,I398029,I398055,I398072,I398080,I398125,I398142,I398159,I398176,I398193,I398210,I398227,I398258,I398275,I398320,I398337,I398354,I398385,I398411,I398419,I398450,I398467,I398484,I398510,I398518,I398535,I398624,I398650,I398667,I398675,I398720,I398737,I398754,I398771,I398788,I398805,I398822,I398853,I398870,I398915,I398932,I398949,I398980,I399006,I399014,I399045,I399062,I399079,I399105,I399113,I399130,I399219,I399245,I399262,I399270,I399315,I399332,I399349,I399366,I399383,I399400,I399417,I399448,I399465,I399510,I399527,I399544,I399575,I399601,I399609,I399640,I399657,I399674,I399700,I399708,I399725,I399814,I399840,I399857,I399865,I399910,I399927,I399944,I399961,I399978,I399995,I400012,I400043,I400060,I400105,I400122,I400139,I400170,I400196,I400204,I400235,I400252,I400269,I400295,I400303,I400320,I400409,I400435,I400452,I400460,I400505,I400522,I400539,I400556,I400573,I400590,I400607,I400638,I400655,I400700,I400717,I400734,I400765,I400791,I400799,I400830,I400847,I400864,I400890,I400898,I400915,I401004,I401030,I401047,I401055,I401100,I401117,I401134,I401151,I401168,I401185,I401202,I401233,I401250,I401295,I401312,I401329,I401360,I401386,I401394,I401425,I401442,I401459,I401485,I401493,I401510,I401599,I401625,I401642,I401650,I401695,I401712,I401729,I401746,I401763,I401780,I401797,I401828,I401845,I401890,I401907,I401924,I401955,I401981,I401989,I402020,I402037,I402054,I402080,I402088,I402105,I402194,I402220,I402237,I402245,I402290,I402307,I402324,I402341,I402358,I402375,I402392,I402423,I402440,I402485,I402502,I402519,I402550,I402576,I402584,I402615,I402632,I402649,I402675,I402683,I402700,I402789,I402815,I402832,I402840,I402885,I402902,I402919,I402936,I402953,I402970,I402987,I403018,I403035,I403080,I403097,I403114,I403145,I403171,I403179,I403210,I403227,I403244,I403270,I403278,I403295,I403384,I403410,I403427,I403435,I403480,I403497,I403514,I403531,I403548,I403565,I403582,I403613,I403630,I403675,I403692,I403709,I403740,I403766,I403774,I403805,I403822,I403839,I403865,I403873,I403890,I403979,I404005,I404022,I404030,I404075,I404092,I404109,I404126,I404143,I404160,I404177,I404208,I404225,I404270,I404287,I404304,I404335,I404361,I404369,I404400,I404417,I404434,I404460,I404468,I404485,I404574,I404600,I404617,I404625,I404670,I404687,I404704,I404721,I404738,I404755,I404772,I404803,I404820,I404865,I404882,I404899,I404930,I404956,I404964,I404995,I405012,I405029,I405055,I405063,I405080,I405169,I405195,I405212,I405220,I405265,I405282,I405299,I405316,I405333,I405350,I405367,I405398,I405415,I405460,I405477,I405494,I405525,I405551,I405559,I405590,I405607,I405624,I405650,I405658,I405675,I405764,I405790,I405807,I405815,I405860,I405877,I405894,I405911,I405928,I405945,I405962,I405993,I406010,I406055,I406072,I406089,I406120,I406146,I406154,I406185,I406202,I406219,I406245,I406253,I406270,I406359,I406385,I406402,I406410,I406455,I406472,I406489,I406506,I406523,I406540,I406557,I406588,I406605,I406650,I406667,I406684,I406715,I406741,I406749,I406780,I406797,I406814,I406840,I406848,I406865,I406954,I406980,I406997,I407005,I407050,I407067,I407084,I407101,I407118,I407135,I407152,I407183,I407200,I407245,I407262,I407279,I407310,I407336,I407344,I407375,I407392,I407409,I407435,I407443,I407460,I407549,I407575,I407592,I407600,I407645,I407662,I407679,I407696,I407713,I407730,I407747,I407778,I407795,I407840,I407857,I407874,I407905,I407931,I407939,I407970,I407987,I408004,I408030,I408038,I408055,I408144,I408170,I408187,I408195,I408240,I408257,I408274,I408291,I408308,I408325,I408342,I408373,I408390,I408435,I408452,I408469,I408500,I408526,I408534,I408565,I408582,I408599,I408625,I408633,I408650,I408739,I408765,I408782,I408790,I408835,I408852,I408869,I408886,I408903,I408920,I408937,I408968,I408985,I409030,I409047,I409064,I409095,I409121,I409129,I409160,I409177,I409194,I409220,I409228,I409245,I409334,I409360,I409377,I409385,I409430,I409447,I409464,I409481,I409498,I409515,I409532,I409563,I409580,I409625,I409642,I409659,I409690,I409716,I409724,I409755,I409772,I409789,I409815,I409823,I409840,I409929,I409955,I409972,I409980,I410025,I410042,I410059,I410076,I410093,I410110,I410127,I410158,I410175,I410220,I410237,I410254,I410285,I410311,I410319,I410350,I410367,I410384,I410410,I410418,I410435,I410524,I410550,I410567,I410575,I410620,I410637,I410654,I410671,I410688,I410705,I410722,I410753,I410770,I410815,I410832,I410849,I410880,I410906,I410914,I410945,I410962,I410979,I411005,I411013,I411030,I411119,I411145,I411162,I411170,I411215,I411232,I411249,I411266,I411283,I411300,I411317,I411348,I411365,I411410,I411427,I411444,I411475,I411501,I411509,I411540,I411557,I411574,I411600,I411608,I411625,I411714,I411740,I411757,I411765,I411810,I411827,I411844,I411861,I411878,I411895,I411912,I411943,I411960,I412005,I412022,I412039,I412070,I412096,I412104,I412135,I412152,I412169,I412195,I412203,I412220,I412309,I412335,I412352,I412360,I412405,I412422,I412439,I412456,I412473,I412490,I412507,I412538,I412555,I412600,I412617,I412634,I412665,I412691,I412699,I412730,I412747,I412764,I412790,I412798,I412815,I412904,I412930,I412947,I412955,I413000,I413017,I413034,I413051,I413068,I413085,I413102,I413133,I413150,I413195,I413212,I413229,I413260,I413286,I413294,I413325,I413342,I413359,I413385,I413393,I413410,I413499,I413525,I413542,I413550,I413595,I413612,I413629,I413646,I413663,I413680,I413697,I413728,I413745,I413790,I413807,I413824,I413855,I413881,I413889,I413920,I413937,I413954,I413980,I413988,I414005,I414094,I414120,I414137,I414145,I414190,I414207,I414224,I414241,I414258,I414275,I414292,I414323,I414340,I414385,I414402,I414419,I414450,I414476,I414484,I414515,I414532,I414549,I414575,I414583,I414600,I414689,I414715,I414732,I414740,I414785,I414802,I414819,I414836,I414853,I414870,I414887,I414918,I414935,I414980,I414997,I415014,I415045,I415071,I415079,I415110,I415127,I415144,I415170,I415178,I415195,I415284,I415310,I415327,I415335,I415380,I415397,I415414,I415431,I415448,I415465,I415482,I415513,I415530,I415575,I415592,I415609,I415640,I415666,I415674,I415705,I415722,I415739,I415765,I415773,I415790,I415879,I415905,I415922,I415930,I415975,I415992,I416009,I416026,I416043,I416060,I416077,I416108,I416125,I416170,I416187,I416204,I416235,I416261,I416269,I416300,I416317,I416334,I416360,I416368,I416385,I416474,I416500,I416517,I416525,I416570,I416587,I416604,I416621,I416638,I416655,I416672,I416703,I416720,I416765,I416782,I416799,I416830,I416856,I416864,I416895,I416912,I416929,I416955,I416963,I416980,I417069,I417095,I417112,I417120,I417165,I417182,I417199,I417216,I417233,I417250,I417267,I417298,I417315,I417360,I417377,I417394,I417425,I417451,I417459,I417490,I417507,I417524,I417550,I417558,I417575,I417664,I417690,I417707,I417715,I417760,I417777,I417794,I417811,I417828,I417845,I417862,I417893,I417910,I417955,I417972,I417989,I418020,I418046,I418054,I418085,I418102,I418119,I418145,I418153,I418170,I418259,I418285,I418302,I418310,I418355,I418372,I418389,I418406,I418423,I418440,I418457,I418488,I418505,I418550,I418567,I418584,I418615,I418641,I418649,I418680,I418697,I418714,I418740,I418748,I418765,I418854,I418880,I418897,I418905,I418950,I418967,I418984,I419001,I419018,I419035,I419052,I419083,I419100,I419145,I419162,I419179,I419210,I419236,I419244,I419275,I419292,I419309,I419335,I419343,I419360,I419449,I419475,I419492,I419500,I419545,I419562,I419579,I419596,I419613,I419630,I419647,I419678,I419695,I419740,I419757,I419774,I419805,I419831,I419839,I419870,I419887,I419904,I419930,I419938,I419955;
not I_0 (I2722,I2690);
DFFARX1 I_1 (I42043,I2683,I2722,I2748,);
nand I_2 (I2756,I2748,I42034);
not I_3 (I2773,I2756);
DFFARX1 I_4 (I2773,I2683,I2722,I2714,);
DFFARX1 I_5 (I42055,I2683,I2722,I2813,);
not I_6 (I2821,I2813);
not I_7 (I2838,I42031);
not I_8 (I2855,I42031);
nand I_9 (I2872,I2821,I2855);
nor I_10 (I2889,I2872,I42031);
DFFARX1 I_11 (I2889,I2683,I2722,I2693,);
nor I_12 (I2920,I42031,I42031);
nand I_13 (I2937,I2813,I2920);
nor I_14 (I2954,I42040,I42034);
nor I_15 (I2696,I2872,I42040);
not I_16 (I2985,I42040);
not I_17 (I3002,I42052);
nand I_18 (I3019,I3002,I42049);
nand I_19 (I3036,I2838,I3019);
not I_20 (I3053,I3036);
nor I_21 (I3070,I42052,I42034);
nor I_22 (I2705,I3053,I3070);
nor I_23 (I3101,I42046,I42052);
and I_24 (I3118,I3101,I2954);
nor I_25 (I3135,I3036,I3118);
DFFARX1 I_26 (I3135,I2683,I2722,I2711,);
nor I_27 (I3166,I2756,I3118);
DFFARX1 I_28 (I3166,I2683,I2722,I2708,);
nor I_29 (I3197,I42046,I42037);
DFFARX1 I_30 (I3197,I2683,I2722,I3223,);
nor I_31 (I3231,I3223,I42031);
nand I_32 (I3248,I3231,I2838);
nand I_33 (I2702,I3248,I2937);
nand I_34 (I2699,I3231,I2985);
not I_35 (I3317,I2690);
DFFARX1 I_36 (I373045,I2683,I3317,I3343,);
nand I_37 (I3351,I3343,I373033);
not I_38 (I3368,I3351);
DFFARX1 I_39 (I3368,I2683,I3317,I3309,);
DFFARX1 I_40 (I373021,I2683,I3317,I3408,);
not I_41 (I3416,I3408);
not I_42 (I3433,I373021);
not I_43 (I3450,I373027);
nand I_44 (I3467,I3416,I3450);
nor I_45 (I3484,I3467,I373021);
DFFARX1 I_46 (I3484,I2683,I3317,I3288,);
nor I_47 (I3515,I373027,I373021);
nand I_48 (I3532,I3408,I3515);
nor I_49 (I3549,I373024,I373039);
nor I_50 (I3291,I3467,I373024);
not I_51 (I3580,I373024);
not I_52 (I3597,I373030);
nand I_53 (I3614,I3597,I373042);
nand I_54 (I3631,I3433,I3614);
not I_55 (I3648,I3631);
nor I_56 (I3665,I373030,I373039);
nor I_57 (I3300,I3648,I3665);
nor I_58 (I3696,I373036,I373030);
and I_59 (I3713,I3696,I3549);
nor I_60 (I3730,I3631,I3713);
DFFARX1 I_61 (I3730,I2683,I3317,I3306,);
nor I_62 (I3761,I3351,I3713);
DFFARX1 I_63 (I3761,I2683,I3317,I3303,);
nor I_64 (I3792,I373036,I373024);
DFFARX1 I_65 (I3792,I2683,I3317,I3818,);
nor I_66 (I3826,I3818,I373027);
nand I_67 (I3843,I3826,I3433);
nand I_68 (I3297,I3843,I3532);
nand I_69 (I3294,I3826,I3580);
not I_70 (I3912,I2690);
DFFARX1 I_71 (I63182,I2683,I3912,I3938,);
nand I_72 (I3946,I3938,I63182);
not I_73 (I3963,I3946);
DFFARX1 I_74 (I3963,I2683,I3912,I3904,);
DFFARX1 I_75 (I63188,I2683,I3912,I4003,);
not I_76 (I4011,I4003);
not I_77 (I4028,I63197);
not I_78 (I4045,I63191);
nand I_79 (I4062,I4011,I4045);
nor I_80 (I4079,I4062,I63197);
DFFARX1 I_81 (I4079,I2683,I3912,I3883,);
nor I_82 (I4110,I63191,I63197);
nand I_83 (I4127,I4003,I4110);
nor I_84 (I4144,I63194,I63200);
nor I_85 (I3886,I4062,I63194);
not I_86 (I4175,I63194);
not I_87 (I4192,I63203);
nand I_88 (I4209,I4192,I63179);
nand I_89 (I4226,I4028,I4209);
not I_90 (I4243,I4226);
nor I_91 (I4260,I63203,I63200);
nor I_92 (I3895,I4243,I4260);
nor I_93 (I4291,I63185,I63203);
and I_94 (I4308,I4291,I4144);
nor I_95 (I4325,I4226,I4308);
DFFARX1 I_96 (I4325,I2683,I3912,I3901,);
nor I_97 (I4356,I3946,I4308);
DFFARX1 I_98 (I4356,I2683,I3912,I3898,);
nor I_99 (I4387,I63185,I63179);
DFFARX1 I_100 (I4387,I2683,I3912,I4413,);
nor I_101 (I4421,I4413,I63191);
nand I_102 (I4438,I4421,I4028);
nand I_103 (I3892,I4438,I4127);
nand I_104 (I3889,I4421,I4175);
not I_105 (I4507,I2690);
DFFARX1 I_106 (I190920,I2683,I4507,I4533,);
nand I_107 (I4541,I4533,I190938);
not I_108 (I4558,I4541);
DFFARX1 I_109 (I4558,I2683,I4507,I4499,);
DFFARX1 I_110 (I190932,I2683,I4507,I4598,);
not I_111 (I4606,I4598);
not I_112 (I4623,I190923);
not I_113 (I4640,I190920);
nand I_114 (I4657,I4606,I4640);
nor I_115 (I4674,I4657,I190923);
DFFARX1 I_116 (I4674,I2683,I4507,I4478,);
nor I_117 (I4705,I190920,I190923);
nand I_118 (I4722,I4598,I4705);
nor I_119 (I4739,I190929,I190917);
nor I_120 (I4481,I4657,I190929);
not I_121 (I4770,I190929);
not I_122 (I4787,I190935);
nand I_123 (I4804,I4787,I190941);
nand I_124 (I4821,I4623,I4804);
not I_125 (I4838,I4821);
nor I_126 (I4855,I190935,I190917);
nor I_127 (I4490,I4838,I4855);
nor I_128 (I4886,I190917,I190935);
and I_129 (I4903,I4886,I4739);
nor I_130 (I4920,I4821,I4903);
DFFARX1 I_131 (I4920,I2683,I4507,I4496,);
nor I_132 (I4951,I4541,I4903);
DFFARX1 I_133 (I4951,I2683,I4507,I4493,);
nor I_134 (I4982,I190917,I190926);
DFFARX1 I_135 (I4982,I2683,I4507,I5008,);
nor I_136 (I5016,I5008,I190920);
nand I_137 (I5033,I5016,I4623);
nand I_138 (I4487,I5033,I4722);
nand I_139 (I4484,I5016,I4770);
not I_140 (I5102,I2690);
DFFARX1 I_141 (I27814,I2683,I5102,I5128,);
nand I_142 (I5136,I5128,I27805);
not I_143 (I5153,I5136);
DFFARX1 I_144 (I5153,I2683,I5102,I5094,);
DFFARX1 I_145 (I27826,I2683,I5102,I5193,);
not I_146 (I5201,I5193);
not I_147 (I5218,I27802);
not I_148 (I5235,I27802);
nand I_149 (I5252,I5201,I5235);
nor I_150 (I5269,I5252,I27802);
DFFARX1 I_151 (I5269,I2683,I5102,I5073,);
nor I_152 (I5300,I27802,I27802);
nand I_153 (I5317,I5193,I5300);
nor I_154 (I5334,I27811,I27805);
nor I_155 (I5076,I5252,I27811);
not I_156 (I5365,I27811);
not I_157 (I5382,I27823);
nand I_158 (I5399,I5382,I27820);
nand I_159 (I5416,I5218,I5399);
not I_160 (I5433,I5416);
nor I_161 (I5450,I27823,I27805);
nor I_162 (I5085,I5433,I5450);
nor I_163 (I5481,I27817,I27823);
and I_164 (I5498,I5481,I5334);
nor I_165 (I5515,I5416,I5498);
DFFARX1 I_166 (I5515,I2683,I5102,I5091,);
nor I_167 (I5546,I5136,I5498);
DFFARX1 I_168 (I5546,I2683,I5102,I5088,);
nor I_169 (I5577,I27817,I27808);
DFFARX1 I_170 (I5577,I2683,I5102,I5603,);
nor I_171 (I5611,I5603,I27802);
nand I_172 (I5628,I5611,I5218);
nand I_173 (I5082,I5628,I5317);
nand I_174 (I5079,I5611,I5365);
not I_175 (I5700,I2690);
DFFARX1 I_176 (I399184,I2683,I5700,I5726,);
DFFARX1 I_177 (I5726,I2683,I5700,I5743,);
not I_178 (I5751,I5743);
nand I_179 (I5768,I399187,I399193);
and I_180 (I5785,I5768,I399202);
DFFARX1 I_181 (I5785,I2683,I5700,I5811,);
DFFARX1 I_182 (I5811,I2683,I5700,I5692,);
DFFARX1 I_183 (I5811,I2683,I5700,I5683,);
DFFARX1 I_184 (I399205,I2683,I5700,I5856,);
nand I_185 (I5864,I5856,I399196);
not I_186 (I5881,I5864);
nor I_187 (I5680,I5726,I5881);
DFFARX1 I_188 (I399184,I2683,I5700,I5921,);
not I_189 (I5929,I5921);
nor I_190 (I5686,I5929,I5751);
nand I_191 (I5674,I5929,I5864);
nand I_192 (I5974,I399211,I399190);
and I_193 (I5991,I5974,I399199);
DFFARX1 I_194 (I5991,I2683,I5700,I6017,);
nor I_195 (I6025,I6017,I5726);
DFFARX1 I_196 (I6025,I2683,I5700,I5668,);
not I_197 (I6056,I6017);
nor I_198 (I6073,I399208,I399190);
not I_199 (I6090,I6073);
nor I_200 (I6107,I5864,I6090);
nor I_201 (I6124,I6056,I6107);
DFFARX1 I_202 (I6124,I2683,I5700,I5689,);
nor I_203 (I6155,I6017,I6090);
nor I_204 (I5677,I5881,I6155);
nor I_205 (I5671,I6017,I6073);
not I_206 (I6227,I2690);
DFFARX1 I_207 (I163573,I2683,I6227,I6253,);
DFFARX1 I_208 (I6253,I2683,I6227,I6270,);
not I_209 (I6278,I6270);
nand I_210 (I6295,I163579,I163567);
and I_211 (I6312,I6295,I163564);
DFFARX1 I_212 (I6312,I2683,I6227,I6338,);
DFFARX1 I_213 (I6338,I2683,I6227,I6219,);
DFFARX1 I_214 (I6338,I2683,I6227,I6210,);
DFFARX1 I_215 (I163576,I2683,I6227,I6383,);
nand I_216 (I6391,I6383,I163570);
not I_217 (I6408,I6391);
nor I_218 (I6207,I6253,I6408);
DFFARX1 I_219 (I163588,I2683,I6227,I6448,);
not I_220 (I6456,I6448);
nor I_221 (I6213,I6456,I6278);
nand I_222 (I6201,I6456,I6391);
nand I_223 (I6501,I163582,I163585);
and I_224 (I6518,I6501,I163567);
DFFARX1 I_225 (I6518,I2683,I6227,I6544,);
nor I_226 (I6552,I6544,I6253);
DFFARX1 I_227 (I6552,I2683,I6227,I6195,);
not I_228 (I6583,I6544);
nor I_229 (I6600,I163564,I163585);
not I_230 (I6617,I6600);
nor I_231 (I6634,I6391,I6617);
nor I_232 (I6651,I6583,I6634);
DFFARX1 I_233 (I6651,I2683,I6227,I6216,);
nor I_234 (I6682,I6544,I6617);
nor I_235 (I6204,I6408,I6682);
nor I_236 (I6198,I6544,I6600);
not I_237 (I6754,I2690);
DFFARX1 I_238 (I256614,I2683,I6754,I6780,);
DFFARX1 I_239 (I6780,I2683,I6754,I6797,);
not I_240 (I6805,I6797);
nand I_241 (I6822,I256605,I256626);
and I_242 (I6839,I6822,I256608);
DFFARX1 I_243 (I6839,I2683,I6754,I6865,);
DFFARX1 I_244 (I6865,I2683,I6754,I6746,);
DFFARX1 I_245 (I6865,I2683,I6754,I6737,);
DFFARX1 I_246 (I256608,I2683,I6754,I6910,);
nand I_247 (I6918,I6910,I256623);
not I_248 (I6935,I6918);
nor I_249 (I6734,I6780,I6935);
DFFARX1 I_250 (I256617,I2683,I6754,I6975,);
not I_251 (I6983,I6975);
nor I_252 (I6740,I6983,I6805);
nand I_253 (I6728,I6983,I6918);
nand I_254 (I7028,I256611,I256620);
and I_255 (I7045,I7028,I256605);
DFFARX1 I_256 (I7045,I2683,I6754,I7071,);
nor I_257 (I7079,I7071,I6780);
DFFARX1 I_258 (I7079,I2683,I6754,I6722,);
not I_259 (I7110,I7071);
nor I_260 (I7127,I256611,I256620);
not I_261 (I7144,I7127);
nor I_262 (I7161,I6918,I7144);
nor I_263 (I7178,I7110,I7161);
DFFARX1 I_264 (I7178,I2683,I6754,I6743,);
nor I_265 (I7209,I7071,I7144);
nor I_266 (I6731,I6935,I7209);
nor I_267 (I6725,I7071,I7127);
not I_268 (I7281,I2690);
DFFARX1 I_269 (I285308,I2683,I7281,I7307,);
DFFARX1 I_270 (I7307,I2683,I7281,I7324,);
not I_271 (I7332,I7324);
nand I_272 (I7349,I285284,I285311);
and I_273 (I7366,I7349,I285296);
DFFARX1 I_274 (I7366,I2683,I7281,I7392,);
DFFARX1 I_275 (I7392,I2683,I7281,I7273,);
DFFARX1 I_276 (I7392,I2683,I7281,I7264,);
DFFARX1 I_277 (I285302,I2683,I7281,I7437,);
nand I_278 (I7445,I7437,I285287);
not I_279 (I7462,I7445);
nor I_280 (I7261,I7307,I7462);
DFFARX1 I_281 (I285305,I2683,I7281,I7502,);
not I_282 (I7510,I7502);
nor I_283 (I7267,I7510,I7332);
nand I_284 (I7255,I7510,I7445);
nand I_285 (I7555,I285290,I285293);
and I_286 (I7572,I7555,I285284);
DFFARX1 I_287 (I7572,I2683,I7281,I7598,);
nor I_288 (I7606,I7598,I7307);
DFFARX1 I_289 (I7606,I2683,I7281,I7249,);
not I_290 (I7637,I7598);
nor I_291 (I7654,I285299,I285293);
not I_292 (I7671,I7654);
nor I_293 (I7688,I7445,I7671);
nor I_294 (I7705,I7637,I7688);
DFFARX1 I_295 (I7705,I2683,I7281,I7270,);
nor I_296 (I7736,I7598,I7671);
nor I_297 (I7258,I7462,I7736);
nor I_298 (I7252,I7598,I7654);
not I_299 (I7808,I2690);
DFFARX1 I_300 (I370301,I2683,I7808,I7834,);
DFFARX1 I_301 (I7834,I2683,I7808,I7851,);
not I_302 (I7859,I7851);
nand I_303 (I7876,I370319,I370313);
and I_304 (I7893,I7876,I370322);
DFFARX1 I_305 (I7893,I2683,I7808,I7919,);
DFFARX1 I_306 (I7919,I2683,I7808,I7800,);
DFFARX1 I_307 (I7919,I2683,I7808,I7791,);
DFFARX1 I_308 (I370307,I2683,I7808,I7964,);
nand I_309 (I7972,I7964,I370316);
not I_310 (I7989,I7972);
nor I_311 (I7788,I7834,I7989);
DFFARX1 I_312 (I370304,I2683,I7808,I8029,);
not I_313 (I8037,I8029);
nor I_314 (I7794,I8037,I7859);
nand I_315 (I7782,I8037,I7972);
nand I_316 (I8082,I370325,I370310);
and I_317 (I8099,I8082,I370304);
DFFARX1 I_318 (I8099,I2683,I7808,I8125,);
nor I_319 (I8133,I8125,I7834);
DFFARX1 I_320 (I8133,I2683,I7808,I7776,);
not I_321 (I8164,I8125);
nor I_322 (I8181,I370301,I370310);
not I_323 (I8198,I8181);
nor I_324 (I8215,I7972,I8198);
nor I_325 (I8232,I8164,I8215);
DFFARX1 I_326 (I8232,I2683,I7808,I7797,);
nor I_327 (I8263,I8125,I8198);
nor I_328 (I7785,I7989,I8263);
nor I_329 (I7779,I8125,I8181);
not I_330 (I8335,I2690);
DFFARX1 I_331 (I304042,I2683,I8335,I8361,);
DFFARX1 I_332 (I8361,I2683,I8335,I8378,);
not I_333 (I8386,I8378);
nand I_334 (I8403,I304018,I304045);
and I_335 (I8420,I8403,I304030);
DFFARX1 I_336 (I8420,I2683,I8335,I8446,);
DFFARX1 I_337 (I8446,I2683,I8335,I8327,);
DFFARX1 I_338 (I8446,I2683,I8335,I8318,);
DFFARX1 I_339 (I304036,I2683,I8335,I8491,);
nand I_340 (I8499,I8491,I304021);
not I_341 (I8516,I8499);
nor I_342 (I8315,I8361,I8516);
DFFARX1 I_343 (I304039,I2683,I8335,I8556,);
not I_344 (I8564,I8556);
nor I_345 (I8321,I8564,I8386);
nand I_346 (I8309,I8564,I8499);
nand I_347 (I8609,I304024,I304027);
and I_348 (I8626,I8609,I304018);
DFFARX1 I_349 (I8626,I2683,I8335,I8652,);
nor I_350 (I8660,I8652,I8361);
DFFARX1 I_351 (I8660,I2683,I8335,I8303,);
not I_352 (I8691,I8652);
nor I_353 (I8708,I304033,I304027);
not I_354 (I8725,I8708);
nor I_355 (I8742,I8499,I8725);
nor I_356 (I8759,I8691,I8742);
DFFARX1 I_357 (I8759,I2683,I8335,I8324,);
nor I_358 (I8790,I8652,I8725);
nor I_359 (I8312,I8516,I8790);
nor I_360 (I8306,I8652,I8708);
not I_361 (I8862,I2690);
DFFARX1 I_362 (I104261,I2683,I8862,I8888,);
DFFARX1 I_363 (I8888,I2683,I8862,I8905,);
not I_364 (I8913,I8905);
nand I_365 (I8930,I104258,I104252);
and I_366 (I8947,I8930,I104246);
DFFARX1 I_367 (I8947,I2683,I8862,I8973,);
DFFARX1 I_368 (I8973,I2683,I8862,I8854,);
DFFARX1 I_369 (I8973,I2683,I8862,I8845,);
DFFARX1 I_370 (I104234,I2683,I8862,I9018,);
nand I_371 (I9026,I9018,I104243);
not I_372 (I9043,I9026);
nor I_373 (I8842,I8888,I9043);
DFFARX1 I_374 (I104240,I2683,I8862,I9083,);
not I_375 (I9091,I9083);
nor I_376 (I8848,I9091,I8913);
nand I_377 (I8836,I9091,I9026);
nand I_378 (I9136,I104237,I104255);
and I_379 (I9153,I9136,I104234);
DFFARX1 I_380 (I9153,I2683,I8862,I9179,);
nor I_381 (I9187,I9179,I8888);
DFFARX1 I_382 (I9187,I2683,I8862,I8830,);
not I_383 (I9218,I9179);
nor I_384 (I9235,I104249,I104255);
not I_385 (I9252,I9235);
nor I_386 (I9269,I9026,I9252);
nor I_387 (I9286,I9218,I9269);
DFFARX1 I_388 (I9286,I2683,I8862,I8851,);
nor I_389 (I9317,I9179,I9252);
nor I_390 (I8839,I9043,I9317);
nor I_391 (I8833,I9179,I9235);
not I_392 (I9389,I2690);
DFFARX1 I_393 (I218667,I2683,I9389,I9415,);
DFFARX1 I_394 (I9415,I2683,I9389,I9432,);
not I_395 (I9440,I9432);
nand I_396 (I9457,I218682,I218685);
and I_397 (I9474,I9457,I218664);
DFFARX1 I_398 (I9474,I2683,I9389,I9500,);
DFFARX1 I_399 (I9500,I2683,I9389,I9381,);
DFFARX1 I_400 (I9500,I2683,I9389,I9372,);
DFFARX1 I_401 (I218670,I2683,I9389,I9545,);
nand I_402 (I9553,I9545,I218676);
not I_403 (I9570,I9553);
nor I_404 (I9369,I9415,I9570);
DFFARX1 I_405 (I218664,I2683,I9389,I9610,);
not I_406 (I9618,I9610);
nor I_407 (I9375,I9618,I9440);
nand I_408 (I9363,I9618,I9553);
nand I_409 (I9663,I218679,I218661);
and I_410 (I9680,I9663,I218673);
DFFARX1 I_411 (I9680,I2683,I9389,I9706,);
nor I_412 (I9714,I9706,I9415);
DFFARX1 I_413 (I9714,I2683,I9389,I9357,);
not I_414 (I9745,I9706);
nor I_415 (I9762,I218661,I218661);
not I_416 (I9779,I9762);
nor I_417 (I9796,I9553,I9779);
nor I_418 (I9813,I9745,I9796);
DFFARX1 I_419 (I9813,I2683,I9389,I9378,);
nor I_420 (I9844,I9706,I9779);
nor I_421 (I9366,I9570,I9844);
nor I_422 (I9360,I9706,I9762);
not I_423 (I9916,I2690);
DFFARX1 I_424 (I151919,I2683,I9916,I9942,);
DFFARX1 I_425 (I9942,I2683,I9916,I9959,);
not I_426 (I9967,I9959);
nand I_427 (I9984,I151919,I151922);
and I_428 (I10001,I9984,I151943);
DFFARX1 I_429 (I10001,I2683,I9916,I10027,);
DFFARX1 I_430 (I10027,I2683,I9916,I9908,);
DFFARX1 I_431 (I10027,I2683,I9916,I9899,);
DFFARX1 I_432 (I151931,I2683,I9916,I10072,);
nand I_433 (I10080,I10072,I151934);
not I_434 (I10097,I10080);
nor I_435 (I9896,I9942,I10097);
DFFARX1 I_436 (I151940,I2683,I9916,I10137,);
not I_437 (I10145,I10137);
nor I_438 (I9902,I10145,I9967);
nand I_439 (I9890,I10145,I10080);
nand I_440 (I10190,I151937,I151925);
and I_441 (I10207,I10190,I151928);
DFFARX1 I_442 (I10207,I2683,I9916,I10233,);
nor I_443 (I10241,I10233,I9942);
DFFARX1 I_444 (I10241,I2683,I9916,I9884,);
not I_445 (I10272,I10233);
nor I_446 (I10289,I151946,I151925);
not I_447 (I10306,I10289);
nor I_448 (I10323,I10080,I10306);
nor I_449 (I10340,I10272,I10323);
DFFARX1 I_450 (I10340,I2683,I9916,I9905,);
nor I_451 (I10371,I10233,I10306);
nor I_452 (I9893,I10097,I10371);
nor I_453 (I9887,I10233,I10289);
not I_454 (I10443,I2690);
DFFARX1 I_455 (I239223,I2683,I10443,I10469,);
DFFARX1 I_456 (I10469,I2683,I10443,I10486,);
not I_457 (I10494,I10486);
nand I_458 (I10511,I239214,I239235);
and I_459 (I10528,I10511,I239217);
DFFARX1 I_460 (I10528,I2683,I10443,I10554,);
DFFARX1 I_461 (I10554,I2683,I10443,I10435,);
DFFARX1 I_462 (I10554,I2683,I10443,I10426,);
DFFARX1 I_463 (I239217,I2683,I10443,I10599,);
nand I_464 (I10607,I10599,I239232);
not I_465 (I10624,I10607);
nor I_466 (I10423,I10469,I10624);
DFFARX1 I_467 (I239226,I2683,I10443,I10664,);
not I_468 (I10672,I10664);
nor I_469 (I10429,I10672,I10494);
nand I_470 (I10417,I10672,I10607);
nand I_471 (I10717,I239220,I239229);
and I_472 (I10734,I10717,I239214);
DFFARX1 I_473 (I10734,I2683,I10443,I10760,);
nor I_474 (I10768,I10760,I10469);
DFFARX1 I_475 (I10768,I2683,I10443,I10411,);
not I_476 (I10799,I10760);
nor I_477 (I10816,I239220,I239229);
not I_478 (I10833,I10816);
nor I_479 (I10850,I10607,I10833);
nor I_480 (I10867,I10799,I10850);
DFFARX1 I_481 (I10867,I2683,I10443,I10432,);
nor I_482 (I10898,I10760,I10833);
nor I_483 (I10420,I10624,I10898);
nor I_484 (I10414,I10760,I10816);
not I_485 (I10970,I2690);
DFFARX1 I_486 (I415844,I2683,I10970,I10996,);
DFFARX1 I_487 (I10996,I2683,I10970,I11013,);
not I_488 (I11021,I11013);
nand I_489 (I11038,I415847,I415853);
and I_490 (I11055,I11038,I415862);
DFFARX1 I_491 (I11055,I2683,I10970,I11081,);
DFFARX1 I_492 (I11081,I2683,I10970,I10962,);
DFFARX1 I_493 (I11081,I2683,I10970,I10953,);
DFFARX1 I_494 (I415865,I2683,I10970,I11126,);
nand I_495 (I11134,I11126,I415856);
not I_496 (I11151,I11134);
nor I_497 (I10950,I10996,I11151);
DFFARX1 I_498 (I415844,I2683,I10970,I11191,);
not I_499 (I11199,I11191);
nor I_500 (I10956,I11199,I11021);
nand I_501 (I10944,I11199,I11134);
nand I_502 (I11244,I415871,I415850);
and I_503 (I11261,I11244,I415859);
DFFARX1 I_504 (I11261,I2683,I10970,I11287,);
nor I_505 (I11295,I11287,I10996);
DFFARX1 I_506 (I11295,I2683,I10970,I10938,);
not I_507 (I11326,I11287);
nor I_508 (I11343,I415868,I415850);
not I_509 (I11360,I11343);
nor I_510 (I11377,I11134,I11360);
nor I_511 (I11394,I11326,I11377);
DFFARX1 I_512 (I11394,I2683,I10970,I10959,);
nor I_513 (I11425,I11287,I11360);
nor I_514 (I10947,I11151,I11425);
nor I_515 (I10941,I11287,I11343);
not I_516 (I11497,I2690);
DFFARX1 I_517 (I330817,I2683,I11497,I11523,);
DFFARX1 I_518 (I11523,I2683,I11497,I11540,);
not I_519 (I11548,I11540);
nand I_520 (I11565,I330805,I330796);
and I_521 (I11582,I11565,I330793);
DFFARX1 I_522 (I11582,I2683,I11497,I11608,);
DFFARX1 I_523 (I11608,I2683,I11497,I11489,);
DFFARX1 I_524 (I11608,I2683,I11497,I11480,);
DFFARX1 I_525 (I330799,I2683,I11497,I11653,);
nand I_526 (I11661,I11653,I330811);
not I_527 (I11678,I11661);
nor I_528 (I11477,I11523,I11678);
DFFARX1 I_529 (I330808,I2683,I11497,I11718,);
not I_530 (I11726,I11718);
nor I_531 (I11483,I11726,I11548);
nand I_532 (I11471,I11726,I11661);
nand I_533 (I11771,I330802,I330796);
and I_534 (I11788,I11771,I330814);
DFFARX1 I_535 (I11788,I2683,I11497,I11814,);
nor I_536 (I11822,I11814,I11523);
DFFARX1 I_537 (I11822,I2683,I11497,I11465,);
not I_538 (I11853,I11814);
nor I_539 (I11870,I330793,I330796);
not I_540 (I11887,I11870);
nor I_541 (I11904,I11661,I11887);
nor I_542 (I11921,I11853,I11904);
DFFARX1 I_543 (I11921,I2683,I11497,I11486,);
nor I_544 (I11952,I11814,I11887);
nor I_545 (I11474,I11678,I11952);
nor I_546 (I11468,I11814,I11870);
not I_547 (I12024,I2690);
DFFARX1 I_548 (I26224,I2683,I12024,I12050,);
DFFARX1 I_549 (I12050,I2683,I12024,I12067,);
not I_550 (I12075,I12067);
nand I_551 (I12092,I26224,I26239);
and I_552 (I12109,I12092,I26242);
DFFARX1 I_553 (I12109,I2683,I12024,I12135,);
DFFARX1 I_554 (I12135,I2683,I12024,I12016,);
DFFARX1 I_555 (I12135,I2683,I12024,I12007,);
DFFARX1 I_556 (I26236,I2683,I12024,I12180,);
nand I_557 (I12188,I12180,I26245);
not I_558 (I12205,I12188);
nor I_559 (I12004,I12050,I12205);
DFFARX1 I_560 (I26221,I2683,I12024,I12245,);
not I_561 (I12253,I12245);
nor I_562 (I12010,I12253,I12075);
nand I_563 (I11998,I12253,I12188);
nand I_564 (I12298,I26221,I26227);
and I_565 (I12315,I12298,I26230);
DFFARX1 I_566 (I12315,I2683,I12024,I12341,);
nor I_567 (I12349,I12341,I12050);
DFFARX1 I_568 (I12349,I2683,I12024,I11992,);
not I_569 (I12380,I12341);
nor I_570 (I12397,I26233,I26227);
not I_571 (I12414,I12397);
nor I_572 (I12431,I12188,I12414);
nor I_573 (I12448,I12380,I12431);
DFFARX1 I_574 (I12448,I2683,I12024,I12013,);
nor I_575 (I12479,I12341,I12414);
nor I_576 (I12001,I12205,I12479);
nor I_577 (I11995,I12341,I12397);
not I_578 (I12551,I2690);
DFFARX1 I_579 (I362607,I2683,I12551,I12577,);
DFFARX1 I_580 (I12577,I2683,I12551,I12594,);
not I_581 (I12602,I12594);
nand I_582 (I12619,I362595,I362586);
and I_583 (I12636,I12619,I362583);
DFFARX1 I_584 (I12636,I2683,I12551,I12662,);
DFFARX1 I_585 (I12662,I2683,I12551,I12543,);
DFFARX1 I_586 (I12662,I2683,I12551,I12534,);
DFFARX1 I_587 (I362589,I2683,I12551,I12707,);
nand I_588 (I12715,I12707,I362601);
not I_589 (I12732,I12715);
nor I_590 (I12531,I12577,I12732);
DFFARX1 I_591 (I362598,I2683,I12551,I12772,);
not I_592 (I12780,I12772);
nor I_593 (I12537,I12780,I12602);
nand I_594 (I12525,I12780,I12715);
nand I_595 (I12825,I362592,I362586);
and I_596 (I12842,I12825,I362604);
DFFARX1 I_597 (I12842,I2683,I12551,I12868,);
nor I_598 (I12876,I12868,I12577);
DFFARX1 I_599 (I12876,I2683,I12551,I12519,);
not I_600 (I12907,I12868);
nor I_601 (I12924,I362583,I362586);
not I_602 (I12941,I12924);
nor I_603 (I12958,I12715,I12941);
nor I_604 (I12975,I12907,I12958);
DFFARX1 I_605 (I12975,I2683,I12551,I12540,);
nor I_606 (I13006,I12868,I12941);
nor I_607 (I12528,I12732,I13006);
nor I_608 (I12522,I12868,I12924);
not I_609 (I13078,I2690);
DFFARX1 I_610 (I82225,I2683,I13078,I13104,);
DFFARX1 I_611 (I13104,I2683,I13078,I13121,);
not I_612 (I13129,I13121);
nand I_613 (I13146,I82243,I82228);
and I_614 (I13163,I13146,I82231);
DFFARX1 I_615 (I13163,I2683,I13078,I13189,);
DFFARX1 I_616 (I13189,I2683,I13078,I13070,);
DFFARX1 I_617 (I13189,I2683,I13078,I13061,);
DFFARX1 I_618 (I82219,I2683,I13078,I13234,);
nand I_619 (I13242,I13234,I82222);
not I_620 (I13259,I13242);
nor I_621 (I13058,I13104,I13259);
DFFARX1 I_622 (I82234,I2683,I13078,I13299,);
not I_623 (I13307,I13299);
nor I_624 (I13064,I13307,I13129);
nand I_625 (I13052,I13307,I13242);
nand I_626 (I13352,I82240,I82237);
and I_627 (I13369,I13352,I82222);
DFFARX1 I_628 (I13369,I2683,I13078,I13395,);
nor I_629 (I13403,I13395,I13104);
DFFARX1 I_630 (I13403,I2683,I13078,I13046,);
not I_631 (I13434,I13395);
nor I_632 (I13451,I82219,I82237);
not I_633 (I13468,I13451);
nor I_634 (I13485,I13242,I13468);
nor I_635 (I13502,I13434,I13485);
DFFARX1 I_636 (I13502,I2683,I13078,I13067,);
nor I_637 (I13533,I13395,I13468);
nor I_638 (I13055,I13259,I13533);
nor I_639 (I13049,I13395,I13451);
not I_640 (I13605,I2690);
DFFARX1 I_641 (I39926,I2683,I13605,I13631,);
DFFARX1 I_642 (I13631,I2683,I13605,I13648,);
not I_643 (I13656,I13648);
nand I_644 (I13673,I39926,I39941);
and I_645 (I13690,I13673,I39944);
DFFARX1 I_646 (I13690,I2683,I13605,I13716,);
DFFARX1 I_647 (I13716,I2683,I13605,I13597,);
DFFARX1 I_648 (I13716,I2683,I13605,I13588,);
DFFARX1 I_649 (I39938,I2683,I13605,I13761,);
nand I_650 (I13769,I13761,I39947);
not I_651 (I13786,I13769);
nor I_652 (I13585,I13631,I13786);
DFFARX1 I_653 (I39923,I2683,I13605,I13826,);
not I_654 (I13834,I13826);
nor I_655 (I13591,I13834,I13656);
nand I_656 (I13579,I13834,I13769);
nand I_657 (I13879,I39923,I39929);
and I_658 (I13896,I13879,I39932);
DFFARX1 I_659 (I13896,I2683,I13605,I13922,);
nor I_660 (I13930,I13922,I13631);
DFFARX1 I_661 (I13930,I2683,I13605,I13573,);
not I_662 (I13961,I13922);
nor I_663 (I13978,I39935,I39929);
not I_664 (I13995,I13978);
nor I_665 (I14012,I13769,I13995);
nor I_666 (I14029,I13961,I14012);
DFFARX1 I_667 (I14029,I2683,I13605,I13594,);
nor I_668 (I14060,I13922,I13995);
nor I_669 (I13582,I13786,I14060);
nor I_670 (I13576,I13922,I13978);
not I_671 (I14132,I2690);
DFFARX1 I_672 (I269262,I2683,I14132,I14158,);
DFFARX1 I_673 (I14158,I2683,I14132,I14175,);
not I_674 (I14183,I14175);
nand I_675 (I14200,I269253,I269274);
and I_676 (I14217,I14200,I269256);
DFFARX1 I_677 (I14217,I2683,I14132,I14243,);
DFFARX1 I_678 (I14243,I2683,I14132,I14124,);
DFFARX1 I_679 (I14243,I2683,I14132,I14115,);
DFFARX1 I_680 (I269256,I2683,I14132,I14288,);
nand I_681 (I14296,I14288,I269271);
not I_682 (I14313,I14296);
nor I_683 (I14112,I14158,I14313);
DFFARX1 I_684 (I269265,I2683,I14132,I14353,);
not I_685 (I14361,I14353);
nor I_686 (I14118,I14361,I14183);
nand I_687 (I14106,I14361,I14296);
nand I_688 (I14406,I269259,I269268);
and I_689 (I14423,I14406,I269253);
DFFARX1 I_690 (I14423,I2683,I14132,I14449,);
nor I_691 (I14457,I14449,I14158);
DFFARX1 I_692 (I14457,I2683,I14132,I14100,);
not I_693 (I14488,I14449);
nor I_694 (I14505,I269259,I269268);
not I_695 (I14522,I14505);
nor I_696 (I14539,I14296,I14522);
nor I_697 (I14556,I14488,I14539);
DFFARX1 I_698 (I14556,I2683,I14132,I14121,);
nor I_699 (I14587,I14449,I14522);
nor I_700 (I14109,I14313,I14587);
nor I_701 (I14103,I14449,I14505);
not I_702 (I14659,I2690);
DFFARX1 I_703 (I240277,I2683,I14659,I14685,);
DFFARX1 I_704 (I14685,I2683,I14659,I14702,);
not I_705 (I14710,I14702);
nand I_706 (I14727,I240268,I240289);
and I_707 (I14744,I14727,I240271);
DFFARX1 I_708 (I14744,I2683,I14659,I14770,);
DFFARX1 I_709 (I14770,I2683,I14659,I14651,);
DFFARX1 I_710 (I14770,I2683,I14659,I14642,);
DFFARX1 I_711 (I240271,I2683,I14659,I14815,);
nand I_712 (I14823,I14815,I240286);
not I_713 (I14840,I14823);
nor I_714 (I14639,I14685,I14840);
DFFARX1 I_715 (I240280,I2683,I14659,I14880,);
not I_716 (I14888,I14880);
nor I_717 (I14645,I14888,I14710);
nand I_718 (I14633,I14888,I14823);
nand I_719 (I14933,I240274,I240283);
and I_720 (I14950,I14933,I240268);
DFFARX1 I_721 (I14950,I2683,I14659,I14976,);
nor I_722 (I14984,I14976,I14685);
DFFARX1 I_723 (I14984,I2683,I14659,I14627,);
not I_724 (I15015,I14976);
nor I_725 (I15032,I240274,I240283);
not I_726 (I15049,I15032);
nor I_727 (I15066,I14823,I15049);
nor I_728 (I15083,I15015,I15066);
DFFARX1 I_729 (I15083,I2683,I14659,I14648,);
nor I_730 (I15114,I14976,I15049);
nor I_731 (I14636,I14840,I15114);
nor I_732 (I14630,I14976,I15032);
not I_733 (I15186,I2690);
DFFARX1 I_734 (I266627,I2683,I15186,I15212,);
DFFARX1 I_735 (I15212,I2683,I15186,I15229,);
not I_736 (I15237,I15229);
nand I_737 (I15254,I266618,I266639);
and I_738 (I15271,I15254,I266621);
DFFARX1 I_739 (I15271,I2683,I15186,I15297,);
DFFARX1 I_740 (I15297,I2683,I15186,I15178,);
DFFARX1 I_741 (I15297,I2683,I15186,I15169,);
DFFARX1 I_742 (I266621,I2683,I15186,I15342,);
nand I_743 (I15350,I15342,I266636);
not I_744 (I15367,I15350);
nor I_745 (I15166,I15212,I15367);
DFFARX1 I_746 (I266630,I2683,I15186,I15407,);
not I_747 (I15415,I15407);
nor I_748 (I15172,I15415,I15237);
nand I_749 (I15160,I15415,I15350);
nand I_750 (I15460,I266624,I266633);
and I_751 (I15477,I15460,I266618);
DFFARX1 I_752 (I15477,I2683,I15186,I15503,);
nor I_753 (I15511,I15503,I15212);
DFFARX1 I_754 (I15511,I2683,I15186,I15154,);
not I_755 (I15542,I15503);
nor I_756 (I15559,I266624,I266633);
not I_757 (I15576,I15559);
nor I_758 (I15593,I15350,I15576);
nor I_759 (I15610,I15542,I15593);
DFFARX1 I_760 (I15610,I2683,I15186,I15175,);
nor I_761 (I15641,I15503,I15576);
nor I_762 (I15163,I15367,I15641);
nor I_763 (I15157,I15503,I15559);
not I_764 (I15713,I2690);
DFFARX1 I_765 (I90032,I2683,I15713,I15739,);
DFFARX1 I_766 (I15739,I2683,I15713,I15756,);
not I_767 (I15764,I15756);
nand I_768 (I15781,I90029,I90023);
and I_769 (I15798,I15781,I90017);
DFFARX1 I_770 (I15798,I2683,I15713,I15824,);
DFFARX1 I_771 (I15824,I2683,I15713,I15705,);
DFFARX1 I_772 (I15824,I2683,I15713,I15696,);
DFFARX1 I_773 (I90005,I2683,I15713,I15869,);
nand I_774 (I15877,I15869,I90014);
not I_775 (I15894,I15877);
nor I_776 (I15693,I15739,I15894);
DFFARX1 I_777 (I90011,I2683,I15713,I15934,);
not I_778 (I15942,I15934);
nor I_779 (I15699,I15942,I15764);
nand I_780 (I15687,I15942,I15877);
nand I_781 (I15987,I90008,I90026);
and I_782 (I16004,I15987,I90005);
DFFARX1 I_783 (I16004,I2683,I15713,I16030,);
nor I_784 (I16038,I16030,I15739);
DFFARX1 I_785 (I16038,I2683,I15713,I15681,);
not I_786 (I16069,I16030);
nor I_787 (I16086,I90020,I90026);
not I_788 (I16103,I16086);
nor I_789 (I16120,I15877,I16103);
nor I_790 (I16137,I16069,I16120);
DFFARX1 I_791 (I16137,I2683,I15713,I15702,);
nor I_792 (I16168,I16030,I16103);
nor I_793 (I15690,I15894,I16168);
nor I_794 (I15684,I16030,I16086);
not I_795 (I16240,I2690);
DFFARX1 I_796 (I125868,I2683,I16240,I16266,);
DFFARX1 I_797 (I16266,I2683,I16240,I16283,);
not I_798 (I16291,I16283);
nand I_799 (I16308,I125865,I125859);
and I_800 (I16325,I16308,I125853);
DFFARX1 I_801 (I16325,I2683,I16240,I16351,);
DFFARX1 I_802 (I16351,I2683,I16240,I16232,);
DFFARX1 I_803 (I16351,I2683,I16240,I16223,);
DFFARX1 I_804 (I125841,I2683,I16240,I16396,);
nand I_805 (I16404,I16396,I125850);
not I_806 (I16421,I16404);
nor I_807 (I16220,I16266,I16421);
DFFARX1 I_808 (I125847,I2683,I16240,I16461,);
not I_809 (I16469,I16461);
nor I_810 (I16226,I16469,I16291);
nand I_811 (I16214,I16469,I16404);
nand I_812 (I16514,I125844,I125862);
and I_813 (I16531,I16514,I125841);
DFFARX1 I_814 (I16531,I2683,I16240,I16557,);
nor I_815 (I16565,I16557,I16266);
DFFARX1 I_816 (I16565,I2683,I16240,I16208,);
not I_817 (I16596,I16557);
nor I_818 (I16613,I125856,I125862);
not I_819 (I16630,I16613);
nor I_820 (I16647,I16404,I16630);
nor I_821 (I16664,I16596,I16647);
DFFARX1 I_822 (I16664,I2683,I16240,I16229,);
nor I_823 (I16695,I16557,I16630);
nor I_824 (I16217,I16421,I16695);
nor I_825 (I16211,I16557,I16613);
not I_826 (I16767,I2690);
DFFARX1 I_827 (I147567,I2683,I16767,I16793,);
DFFARX1 I_828 (I16793,I2683,I16767,I16810,);
not I_829 (I16818,I16810);
nand I_830 (I16835,I147567,I147570);
and I_831 (I16852,I16835,I147591);
DFFARX1 I_832 (I16852,I2683,I16767,I16878,);
DFFARX1 I_833 (I16878,I2683,I16767,I16759,);
DFFARX1 I_834 (I16878,I2683,I16767,I16750,);
DFFARX1 I_835 (I147579,I2683,I16767,I16923,);
nand I_836 (I16931,I16923,I147582);
not I_837 (I16948,I16931);
nor I_838 (I16747,I16793,I16948);
DFFARX1 I_839 (I147588,I2683,I16767,I16988,);
not I_840 (I16996,I16988);
nor I_841 (I16753,I16996,I16818);
nand I_842 (I16741,I16996,I16931);
nand I_843 (I17041,I147585,I147573);
and I_844 (I17058,I17041,I147576);
DFFARX1 I_845 (I17058,I2683,I16767,I17084,);
nor I_846 (I17092,I17084,I16793);
DFFARX1 I_847 (I17092,I2683,I16767,I16735,);
not I_848 (I17123,I17084);
nor I_849 (I17140,I147594,I147573);
not I_850 (I17157,I17140);
nor I_851 (I17174,I16931,I17157);
nor I_852 (I17191,I17123,I17174);
DFFARX1 I_853 (I17191,I2683,I16767,I16756,);
nor I_854 (I17222,I17084,I17157);
nor I_855 (I16744,I16948,I17222);
nor I_856 (I16738,I17084,I17140);
not I_857 (I17294,I2690);
DFFARX1 I_858 (I285954,I2683,I17294,I17320,);
DFFARX1 I_859 (I17320,I2683,I17294,I17337,);
not I_860 (I17345,I17337);
nand I_861 (I17362,I285930,I285957);
and I_862 (I17379,I17362,I285942);
DFFARX1 I_863 (I17379,I2683,I17294,I17405,);
DFFARX1 I_864 (I17405,I2683,I17294,I17286,);
DFFARX1 I_865 (I17405,I2683,I17294,I17277,);
DFFARX1 I_866 (I285948,I2683,I17294,I17450,);
nand I_867 (I17458,I17450,I285933);
not I_868 (I17475,I17458);
nor I_869 (I17274,I17320,I17475);
DFFARX1 I_870 (I285951,I2683,I17294,I17515,);
not I_871 (I17523,I17515);
nor I_872 (I17280,I17523,I17345);
nand I_873 (I17268,I17523,I17458);
nand I_874 (I17568,I285936,I285939);
and I_875 (I17585,I17568,I285930);
DFFARX1 I_876 (I17585,I2683,I17294,I17611,);
nor I_877 (I17619,I17611,I17320);
DFFARX1 I_878 (I17619,I2683,I17294,I17262,);
not I_879 (I17650,I17611);
nor I_880 (I17667,I285945,I285939);
not I_881 (I17684,I17667);
nor I_882 (I17701,I17458,I17684);
nor I_883 (I17718,I17650,I17701);
DFFARX1 I_884 (I17718,I2683,I17294,I17283,);
nor I_885 (I17749,I17611,I17684);
nor I_886 (I17271,I17475,I17749);
nor I_887 (I17265,I17611,I17667);
not I_888 (I17821,I2690);
DFFARX1 I_889 (I353359,I2683,I17821,I17847,);
DFFARX1 I_890 (I17847,I2683,I17821,I17864,);
not I_891 (I17872,I17864);
nand I_892 (I17889,I353347,I353338);
and I_893 (I17906,I17889,I353335);
DFFARX1 I_894 (I17906,I2683,I17821,I17932,);
DFFARX1 I_895 (I17932,I2683,I17821,I17813,);
DFFARX1 I_896 (I17932,I2683,I17821,I17804,);
DFFARX1 I_897 (I353341,I2683,I17821,I17977,);
nand I_898 (I17985,I17977,I353353);
not I_899 (I18002,I17985);
nor I_900 (I17801,I17847,I18002);
DFFARX1 I_901 (I353350,I2683,I17821,I18042,);
not I_902 (I18050,I18042);
nor I_903 (I17807,I18050,I17872);
nand I_904 (I17795,I18050,I17985);
nand I_905 (I18095,I353344,I353338);
and I_906 (I18112,I18095,I353356);
DFFARX1 I_907 (I18112,I2683,I17821,I18138,);
nor I_908 (I18146,I18138,I17847);
DFFARX1 I_909 (I18146,I2683,I17821,I17789,);
not I_910 (I18177,I18138);
nor I_911 (I18194,I353335,I353338);
not I_912 (I18211,I18194);
nor I_913 (I18228,I17985,I18211);
nor I_914 (I18245,I18177,I18228);
DFFARX1 I_915 (I18245,I2683,I17821,I17810,);
nor I_916 (I18276,I18138,I18211);
nor I_917 (I17798,I18002,I18276);
nor I_918 (I17792,I18138,I18194);
not I_919 (I18348,I2690);
DFFARX1 I_920 (I246601,I2683,I18348,I18374,);
DFFARX1 I_921 (I18374,I2683,I18348,I18391,);
not I_922 (I18399,I18391);
nand I_923 (I18416,I246592,I246613);
and I_924 (I18433,I18416,I246595);
DFFARX1 I_925 (I18433,I2683,I18348,I18459,);
DFFARX1 I_926 (I18459,I2683,I18348,I18340,);
DFFARX1 I_927 (I18459,I2683,I18348,I18331,);
DFFARX1 I_928 (I246595,I2683,I18348,I18504,);
nand I_929 (I18512,I18504,I246610);
not I_930 (I18529,I18512);
nor I_931 (I18328,I18374,I18529);
DFFARX1 I_932 (I246604,I2683,I18348,I18569,);
not I_933 (I18577,I18569);
nor I_934 (I18334,I18577,I18399);
nand I_935 (I18322,I18577,I18512);
nand I_936 (I18622,I246598,I246607);
and I_937 (I18639,I18622,I246592);
DFFARX1 I_938 (I18639,I2683,I18348,I18665,);
nor I_939 (I18673,I18665,I18374);
DFFARX1 I_940 (I18673,I2683,I18348,I18316,);
not I_941 (I18704,I18665);
nor I_942 (I18721,I246598,I246607);
not I_943 (I18738,I18721);
nor I_944 (I18755,I18512,I18738);
nor I_945 (I18772,I18704,I18755);
DFFARX1 I_946 (I18772,I2683,I18348,I18337,);
nor I_947 (I18803,I18665,I18738);
nor I_948 (I18325,I18529,I18803);
nor I_949 (I18319,I18665,I18721);
not I_950 (I18875,I2690);
DFFARX1 I_951 (I410501,I2683,I18875,I18901,);
not I_952 (I18909,I18901);
nand I_953 (I18926,I410495,I410516);
and I_954 (I18943,I18926,I410492);
DFFARX1 I_955 (I18943,I2683,I18875,I18969,);
DFFARX1 I_956 (I410513,I2683,I18875,I18986,);
and I_957 (I18994,I18986,I410510);
nor I_958 (I19011,I18969,I18994);
DFFARX1 I_959 (I19011,I2683,I18875,I18843,);
nand I_960 (I19042,I18986,I410510);
nand I_961 (I19059,I18909,I19042);
not I_962 (I18855,I19059);
DFFARX1 I_963 (I410498,I2683,I18875,I19099,);
DFFARX1 I_964 (I19099,I2683,I18875,I18864,);
nand I_965 (I19121,I410507,I410504);
and I_966 (I19138,I19121,I410489);
DFFARX1 I_967 (I19138,I2683,I18875,I19164,);
DFFARX1 I_968 (I19164,I2683,I18875,I19181,);
not I_969 (I18867,I19181);
not I_970 (I19203,I19164);
nand I_971 (I18852,I19203,I19042);
nor I_972 (I19234,I410489,I410504);
not I_973 (I19251,I19234);
nor I_974 (I19268,I19203,I19251);
nor I_975 (I19285,I18909,I19268);
DFFARX1 I_976 (I19285,I2683,I18875,I18861,);
nor I_977 (I19316,I18969,I19251);
nor I_978 (I18849,I19164,I19316);
nor I_979 (I18858,I19099,I19234);
nor I_980 (I18846,I18969,I19234);
not I_981 (I19402,I2690);
DFFARX1 I_982 (I139425,I2683,I19402,I19428,);
not I_983 (I19436,I19428);
nand I_984 (I19453,I139419,I139410);
and I_985 (I19470,I19453,I139431);
DFFARX1 I_986 (I19470,I2683,I19402,I19496,);
DFFARX1 I_987 (I139413,I2683,I19402,I19513,);
and I_988 (I19521,I19513,I139407);
nor I_989 (I19538,I19496,I19521);
DFFARX1 I_990 (I19538,I2683,I19402,I19370,);
nand I_991 (I19569,I19513,I139407);
nand I_992 (I19586,I19436,I19569);
not I_993 (I19382,I19586);
DFFARX1 I_994 (I139407,I2683,I19402,I19626,);
DFFARX1 I_995 (I19626,I2683,I19402,I19391,);
nand I_996 (I19648,I139434,I139416);
and I_997 (I19665,I19648,I139422);
DFFARX1 I_998 (I19665,I2683,I19402,I19691,);
DFFARX1 I_999 (I19691,I2683,I19402,I19708,);
not I_1000 (I19394,I19708);
not I_1001 (I19730,I19691);
nand I_1002 (I19379,I19730,I19569);
nor I_1003 (I19761,I139428,I139416);
not I_1004 (I19778,I19761);
nor I_1005 (I19795,I19730,I19778);
nor I_1006 (I19812,I19436,I19795);
DFFARX1 I_1007 (I19812,I2683,I19402,I19388,);
nor I_1008 (I19843,I19496,I19778);
nor I_1009 (I19376,I19691,I19843);
nor I_1010 (I19385,I19626,I19761);
nor I_1011 (I19373,I19496,I19761);
not I_1012 (I19929,I2690);
DFFARX1 I_1013 (I348139,I2683,I19929,I19955,);
not I_1014 (I19963,I19955);
nand I_1015 (I19980,I348154,I348133);
and I_1016 (I19997,I19980,I348136);
DFFARX1 I_1017 (I19997,I2683,I19929,I20023,);
DFFARX1 I_1018 (I348157,I2683,I19929,I20040,);
and I_1019 (I20048,I20040,I348136);
nor I_1020 (I20065,I20023,I20048);
DFFARX1 I_1021 (I20065,I2683,I19929,I19897,);
nand I_1022 (I20096,I20040,I348136);
nand I_1023 (I20113,I19963,I20096);
not I_1024 (I19909,I20113);
DFFARX1 I_1025 (I348133,I2683,I19929,I20153,);
DFFARX1 I_1026 (I20153,I2683,I19929,I19918,);
nand I_1027 (I20175,I348145,I348142);
and I_1028 (I20192,I20175,I348148);
DFFARX1 I_1029 (I20192,I2683,I19929,I20218,);
DFFARX1 I_1030 (I20218,I2683,I19929,I20235,);
not I_1031 (I19921,I20235);
not I_1032 (I20257,I20218);
nand I_1033 (I19906,I20257,I20096);
nor I_1034 (I20288,I348151,I348142);
not I_1035 (I20305,I20288);
nor I_1036 (I20322,I20257,I20305);
nor I_1037 (I20339,I19963,I20322);
DFFARX1 I_1038 (I20339,I2683,I19929,I19915,);
nor I_1039 (I20370,I20023,I20305);
nor I_1040 (I19903,I20218,I20370);
nor I_1041 (I19912,I20153,I20288);
nor I_1042 (I19900,I20023,I20288);
not I_1043 (I20456,I2690);
DFFARX1 I_1044 (I164162,I2683,I20456,I20482,);
not I_1045 (I20490,I20482);
nand I_1046 (I20507,I164183,I164177);
and I_1047 (I20524,I20507,I164159);
DFFARX1 I_1048 (I20524,I2683,I20456,I20550,);
DFFARX1 I_1049 (I164162,I2683,I20456,I20567,);
and I_1050 (I20575,I20567,I164171);
nor I_1051 (I20592,I20550,I20575);
DFFARX1 I_1052 (I20592,I2683,I20456,I20424,);
nand I_1053 (I20623,I20567,I164171);
nand I_1054 (I20640,I20490,I20623);
not I_1055 (I20436,I20640);
DFFARX1 I_1056 (I164168,I2683,I20456,I20680,);
DFFARX1 I_1057 (I20680,I2683,I20456,I20445,);
nand I_1058 (I20702,I164174,I164165);
and I_1059 (I20719,I20702,I164159);
DFFARX1 I_1060 (I20719,I2683,I20456,I20745,);
DFFARX1 I_1061 (I20745,I2683,I20456,I20762,);
not I_1062 (I20448,I20762);
not I_1063 (I20784,I20745);
nand I_1064 (I20433,I20784,I20623);
nor I_1065 (I20815,I164180,I164165);
not I_1066 (I20832,I20815);
nor I_1067 (I20849,I20784,I20832);
nor I_1068 (I20866,I20490,I20849);
DFFARX1 I_1069 (I20866,I2683,I20456,I20442,);
nor I_1070 (I20897,I20550,I20832);
nor I_1071 (I20430,I20745,I20897);
nor I_1072 (I20439,I20680,I20815);
nor I_1073 (I20427,I20550,I20815);
not I_1074 (I20983,I2690);
DFFARX1 I_1075 (I80446,I2683,I20983,I21009,);
not I_1076 (I21017,I21009);
nand I_1077 (I21034,I80440,I80434);
and I_1078 (I21051,I21034,I80455);
DFFARX1 I_1079 (I21051,I2683,I20983,I21077,);
DFFARX1 I_1080 (I80452,I2683,I20983,I21094,);
and I_1081 (I21102,I21094,I80449);
nor I_1082 (I21119,I21077,I21102);
DFFARX1 I_1083 (I21119,I2683,I20983,I20951,);
nand I_1084 (I21150,I21094,I80449);
nand I_1085 (I21167,I21017,I21150);
not I_1086 (I20963,I21167);
DFFARX1 I_1087 (I80434,I2683,I20983,I21207,);
DFFARX1 I_1088 (I21207,I2683,I20983,I20972,);
nand I_1089 (I21229,I80437,I80437);
and I_1090 (I21246,I21229,I80458);
DFFARX1 I_1091 (I21246,I2683,I20983,I21272,);
DFFARX1 I_1092 (I21272,I2683,I20983,I21289,);
not I_1093 (I20975,I21289);
not I_1094 (I21311,I21272);
nand I_1095 (I20960,I21311,I21150);
nor I_1096 (I21342,I80443,I80437);
not I_1097 (I21359,I21342);
nor I_1098 (I21376,I21311,I21359);
nor I_1099 (I21393,I21017,I21376);
DFFARX1 I_1100 (I21393,I2683,I20983,I20969,);
nor I_1101 (I21424,I21077,I21359);
nor I_1102 (I20957,I21272,I21424);
nor I_1103 (I20966,I21207,I21342);
nor I_1104 (I20954,I21077,I21342);
not I_1105 (I21510,I2690);
DFFARX1 I_1106 (I155237,I2683,I21510,I21536,);
not I_1107 (I21544,I21536);
nand I_1108 (I21561,I155258,I155252);
and I_1109 (I21578,I21561,I155234);
DFFARX1 I_1110 (I21578,I2683,I21510,I21604,);
DFFARX1 I_1111 (I155237,I2683,I21510,I21621,);
and I_1112 (I21629,I21621,I155246);
nor I_1113 (I21646,I21604,I21629);
DFFARX1 I_1114 (I21646,I2683,I21510,I21478,);
nand I_1115 (I21677,I21621,I155246);
nand I_1116 (I21694,I21544,I21677);
not I_1117 (I21490,I21694);
DFFARX1 I_1118 (I155243,I2683,I21510,I21734,);
DFFARX1 I_1119 (I21734,I2683,I21510,I21499,);
nand I_1120 (I21756,I155249,I155240);
and I_1121 (I21773,I21756,I155234);
DFFARX1 I_1122 (I21773,I2683,I21510,I21799,);
DFFARX1 I_1123 (I21799,I2683,I21510,I21816,);
not I_1124 (I21502,I21816);
not I_1125 (I21838,I21799);
nand I_1126 (I21487,I21838,I21677);
nor I_1127 (I21869,I155255,I155240);
not I_1128 (I21886,I21869);
nor I_1129 (I21903,I21838,I21886);
nor I_1130 (I21920,I21544,I21903);
DFFARX1 I_1131 (I21920,I2683,I21510,I21496,);
nor I_1132 (I21951,I21604,I21886);
nor I_1133 (I21484,I21799,I21951);
nor I_1134 (I21493,I21734,I21869);
nor I_1135 (I21481,I21604,I21869);
not I_1136 (I22037,I2690);
DFFARX1 I_1137 (I415261,I2683,I22037,I22063,);
not I_1138 (I22071,I22063);
nand I_1139 (I22088,I415255,I415276);
and I_1140 (I22105,I22088,I415252);
DFFARX1 I_1141 (I22105,I2683,I22037,I22131,);
DFFARX1 I_1142 (I415273,I2683,I22037,I22148,);
and I_1143 (I22156,I22148,I415270);
nor I_1144 (I22173,I22131,I22156);
DFFARX1 I_1145 (I22173,I2683,I22037,I22005,);
nand I_1146 (I22204,I22148,I415270);
nand I_1147 (I22221,I22071,I22204);
not I_1148 (I22017,I22221);
DFFARX1 I_1149 (I415258,I2683,I22037,I22261,);
DFFARX1 I_1150 (I22261,I2683,I22037,I22026,);
nand I_1151 (I22283,I415267,I415264);
and I_1152 (I22300,I22283,I415249);
DFFARX1 I_1153 (I22300,I2683,I22037,I22326,);
DFFARX1 I_1154 (I22326,I2683,I22037,I22343,);
not I_1155 (I22029,I22343);
not I_1156 (I22365,I22326);
nand I_1157 (I22014,I22365,I22204);
nor I_1158 (I22396,I415249,I415264);
not I_1159 (I22413,I22396);
nor I_1160 (I22430,I22365,I22413);
nor I_1161 (I22447,I22071,I22430);
DFFARX1 I_1162 (I22447,I2683,I22037,I22023,);
nor I_1163 (I22478,I22131,I22413);
nor I_1164 (I22011,I22326,I22478);
nor I_1165 (I22020,I22261,I22396);
nor I_1166 (I22008,I22131,I22396);
not I_1167 (I22564,I2690);
DFFARX1 I_1168 (I290461,I2683,I22564,I22590,);
not I_1169 (I22598,I22590);
nand I_1170 (I22615,I290479,I290473);
and I_1171 (I22632,I22615,I290452);
DFFARX1 I_1172 (I22632,I2683,I22564,I22658,);
DFFARX1 I_1173 (I290470,I2683,I22564,I22675,);
and I_1174 (I22683,I22675,I290455);
nor I_1175 (I22700,I22658,I22683);
DFFARX1 I_1176 (I22700,I2683,I22564,I22532,);
nand I_1177 (I22731,I22675,I290455);
nand I_1178 (I22748,I22598,I22731);
not I_1179 (I22544,I22748);
DFFARX1 I_1180 (I290467,I2683,I22564,I22788,);
DFFARX1 I_1181 (I22788,I2683,I22564,I22553,);
nand I_1182 (I22810,I290476,I290464);
and I_1183 (I22827,I22810,I290458);
DFFARX1 I_1184 (I22827,I2683,I22564,I22853,);
DFFARX1 I_1185 (I22853,I2683,I22564,I22870,);
not I_1186 (I22556,I22870);
not I_1187 (I22892,I22853);
nand I_1188 (I22541,I22892,I22731);
nor I_1189 (I22923,I290452,I290464);
not I_1190 (I22940,I22923);
nor I_1191 (I22957,I22892,I22940);
nor I_1192 (I22974,I22598,I22957);
DFFARX1 I_1193 (I22974,I2683,I22564,I22550,);
nor I_1194 (I23005,I22658,I22940);
nor I_1195 (I22538,I22853,I23005);
nor I_1196 (I22547,I22788,I22923);
nor I_1197 (I22535,I22658,I22923);
not I_1198 (I23091,I2690);
DFFARX1 I_1199 (I318811,I2683,I23091,I23117,);
not I_1200 (I23125,I23117);
nand I_1201 (I23142,I318808,I318814);
and I_1202 (I23159,I23142,I318811);
DFFARX1 I_1203 (I23159,I2683,I23091,I23185,);
DFFARX1 I_1204 (I318814,I2683,I23091,I23202,);
and I_1205 (I23210,I23202,I318808);
nor I_1206 (I23227,I23185,I23210);
DFFARX1 I_1207 (I23227,I2683,I23091,I23059,);
nand I_1208 (I23258,I23202,I318808);
nand I_1209 (I23275,I23125,I23258);
not I_1210 (I23071,I23275);
DFFARX1 I_1211 (I318817,I2683,I23091,I23315,);
DFFARX1 I_1212 (I23315,I2683,I23091,I23080,);
nand I_1213 (I23337,I318820,I318829);
and I_1214 (I23354,I23337,I318823);
DFFARX1 I_1215 (I23354,I2683,I23091,I23380,);
DFFARX1 I_1216 (I23380,I2683,I23091,I23397,);
not I_1217 (I23083,I23397);
not I_1218 (I23419,I23380);
nand I_1219 (I23068,I23419,I23258);
nor I_1220 (I23450,I318826,I318829);
not I_1221 (I23467,I23450);
nor I_1222 (I23484,I23419,I23467);
nor I_1223 (I23501,I23125,I23484);
DFFARX1 I_1224 (I23501,I2683,I23091,I23077,);
nor I_1225 (I23532,I23185,I23467);
nor I_1226 (I23065,I23380,I23532);
nor I_1227 (I23074,I23315,I23450);
nor I_1228 (I23062,I23185,I23450);
not I_1229 (I23618,I2690);
DFFARX1 I_1230 (I158807,I2683,I23618,I23644,);
not I_1231 (I23652,I23644);
nand I_1232 (I23669,I158828,I158822);
and I_1233 (I23686,I23669,I158804);
DFFARX1 I_1234 (I23686,I2683,I23618,I23712,);
DFFARX1 I_1235 (I158807,I2683,I23618,I23729,);
and I_1236 (I23737,I23729,I158816);
nor I_1237 (I23754,I23712,I23737);
DFFARX1 I_1238 (I23754,I2683,I23618,I23586,);
nand I_1239 (I23785,I23729,I158816);
nand I_1240 (I23802,I23652,I23785);
not I_1241 (I23598,I23802);
DFFARX1 I_1242 (I158813,I2683,I23618,I23842,);
DFFARX1 I_1243 (I23842,I2683,I23618,I23607,);
nand I_1244 (I23864,I158819,I158810);
and I_1245 (I23881,I23864,I158804);
DFFARX1 I_1246 (I23881,I2683,I23618,I23907,);
DFFARX1 I_1247 (I23907,I2683,I23618,I23924,);
not I_1248 (I23610,I23924);
not I_1249 (I23946,I23907);
nand I_1250 (I23595,I23946,I23785);
nor I_1251 (I23977,I158825,I158810);
not I_1252 (I23994,I23977);
nor I_1253 (I24011,I23946,I23994);
nor I_1254 (I24028,I23652,I24011);
DFFARX1 I_1255 (I24028,I2683,I23618,I23604,);
nor I_1256 (I24059,I23712,I23994);
nor I_1257 (I23592,I23907,I24059);
nor I_1258 (I23601,I23842,I23977);
nor I_1259 (I23589,I23712,I23977);
not I_1260 (I24145,I2690);
DFFARX1 I_1261 (I132897,I2683,I24145,I24171,);
not I_1262 (I24179,I24171);
nand I_1263 (I24196,I132891,I132882);
and I_1264 (I24213,I24196,I132903);
DFFARX1 I_1265 (I24213,I2683,I24145,I24239,);
DFFARX1 I_1266 (I132885,I2683,I24145,I24256,);
and I_1267 (I24264,I24256,I132879);
nor I_1268 (I24281,I24239,I24264);
DFFARX1 I_1269 (I24281,I2683,I24145,I24113,);
nand I_1270 (I24312,I24256,I132879);
nand I_1271 (I24329,I24179,I24312);
not I_1272 (I24125,I24329);
DFFARX1 I_1273 (I132879,I2683,I24145,I24369,);
DFFARX1 I_1274 (I24369,I2683,I24145,I24134,);
nand I_1275 (I24391,I132906,I132888);
and I_1276 (I24408,I24391,I132894);
DFFARX1 I_1277 (I24408,I2683,I24145,I24434,);
DFFARX1 I_1278 (I24434,I2683,I24145,I24451,);
not I_1279 (I24137,I24451);
not I_1280 (I24473,I24434);
nand I_1281 (I24122,I24473,I24312);
nor I_1282 (I24504,I132900,I132888);
not I_1283 (I24521,I24504);
nor I_1284 (I24538,I24473,I24521);
nor I_1285 (I24555,I24179,I24538);
DFFARX1 I_1286 (I24555,I2683,I24145,I24131,);
nor I_1287 (I24586,I24239,I24521);
nor I_1288 (I24119,I24434,I24586);
nor I_1289 (I24128,I24369,I24504);
nor I_1290 (I24116,I24239,I24504);
not I_1291 (I24672,I2690);
DFFARX1 I_1292 (I326753,I2683,I24672,I24698,);
not I_1293 (I24706,I24698);
nand I_1294 (I24723,I326768,I326747);
and I_1295 (I24740,I24723,I326750);
DFFARX1 I_1296 (I24740,I2683,I24672,I24766,);
DFFARX1 I_1297 (I326771,I2683,I24672,I24783,);
and I_1298 (I24791,I24783,I326750);
nor I_1299 (I24808,I24766,I24791);
DFFARX1 I_1300 (I24808,I2683,I24672,I24640,);
nand I_1301 (I24839,I24783,I326750);
nand I_1302 (I24856,I24706,I24839);
not I_1303 (I24652,I24856);
DFFARX1 I_1304 (I326747,I2683,I24672,I24896,);
DFFARX1 I_1305 (I24896,I2683,I24672,I24661,);
nand I_1306 (I24918,I326759,I326756);
and I_1307 (I24935,I24918,I326762);
DFFARX1 I_1308 (I24935,I2683,I24672,I24961,);
DFFARX1 I_1309 (I24961,I2683,I24672,I24978,);
not I_1310 (I24664,I24978);
not I_1311 (I25000,I24961);
nand I_1312 (I24649,I25000,I24839);
nor I_1313 (I25031,I326765,I326756);
not I_1314 (I25048,I25031);
nor I_1315 (I25065,I25000,I25048);
nor I_1316 (I25082,I24706,I25065);
DFFARX1 I_1317 (I25082,I2683,I24672,I24658,);
nor I_1318 (I25113,I24766,I25048);
nor I_1319 (I24646,I24961,I25113);
nor I_1320 (I24655,I24896,I25031);
nor I_1321 (I24643,I24766,I25031);
not I_1322 (I25199,I2690);
DFFARX1 I_1323 (I388274,I2683,I25199,I25225,);
not I_1324 (I25233,I25225);
nand I_1325 (I25250,I388277,I388271);
and I_1326 (I25267,I25250,I388268);
DFFARX1 I_1327 (I25267,I2683,I25199,I25293,);
DFFARX1 I_1328 (I388253,I2683,I25199,I25310,);
and I_1329 (I25318,I25310,I388262);
nor I_1330 (I25335,I25293,I25318);
DFFARX1 I_1331 (I25335,I2683,I25199,I25167,);
nand I_1332 (I25366,I25310,I388262);
nand I_1333 (I25383,I25233,I25366);
not I_1334 (I25179,I25383);
DFFARX1 I_1335 (I388253,I2683,I25199,I25423,);
DFFARX1 I_1336 (I25423,I2683,I25199,I25188,);
nand I_1337 (I25445,I388256,I388259);
and I_1338 (I25462,I25445,I388265);
DFFARX1 I_1339 (I25462,I2683,I25199,I25488,);
DFFARX1 I_1340 (I25488,I2683,I25199,I25505,);
not I_1341 (I25191,I25505);
not I_1342 (I25527,I25488);
nand I_1343 (I25176,I25527,I25366);
nor I_1344 (I25558,I388256,I388259);
not I_1345 (I25575,I25558);
nor I_1346 (I25592,I25527,I25575);
nor I_1347 (I25609,I25233,I25592);
DFFARX1 I_1348 (I25609,I2683,I25199,I25185,);
nor I_1349 (I25640,I25293,I25575);
nor I_1350 (I25173,I25488,I25640);
nor I_1351 (I25182,I25423,I25558);
nor I_1352 (I25170,I25293,I25558);
not I_1353 (I25726,I2690);
DFFARX1 I_1354 (I302089,I2683,I25726,I25752,);
not I_1355 (I25760,I25752);
nand I_1356 (I25777,I302107,I302101);
and I_1357 (I25794,I25777,I302080);
DFFARX1 I_1358 (I25794,I2683,I25726,I25820,);
DFFARX1 I_1359 (I302098,I2683,I25726,I25837,);
and I_1360 (I25845,I25837,I302083);
nor I_1361 (I25862,I25820,I25845);
DFFARX1 I_1362 (I25862,I2683,I25726,I25694,);
nand I_1363 (I25893,I25837,I302083);
nand I_1364 (I25910,I25760,I25893);
not I_1365 (I25706,I25910);
DFFARX1 I_1366 (I302095,I2683,I25726,I25950,);
DFFARX1 I_1367 (I25950,I2683,I25726,I25715,);
nand I_1368 (I25972,I302104,I302092);
and I_1369 (I25989,I25972,I302086);
DFFARX1 I_1370 (I25989,I2683,I25726,I26015,);
DFFARX1 I_1371 (I26015,I2683,I25726,I26032,);
not I_1372 (I25718,I26032);
not I_1373 (I26054,I26015);
nand I_1374 (I25703,I26054,I25893);
nor I_1375 (I26085,I302080,I302092);
not I_1376 (I26102,I26085);
nor I_1377 (I26119,I26054,I26102);
nor I_1378 (I26136,I25760,I26119);
DFFARX1 I_1379 (I26136,I2683,I25726,I25712,);
nor I_1380 (I26167,I25820,I26102);
nor I_1381 (I25700,I26015,I26167);
nor I_1382 (I25709,I25950,I26085);
nor I_1383 (I25697,I25820,I26085);
not I_1384 (I26253,I2690);
DFFARX1 I_1385 (I368675,I2683,I26253,I26279,);
not I_1386 (I26287,I26279);
nand I_1387 (I26304,I368669,I368690);
and I_1388 (I26321,I26304,I368681);
DFFARX1 I_1389 (I26321,I2683,I26253,I26347,);
DFFARX1 I_1390 (I368672,I2683,I26253,I26364,);
and I_1391 (I26372,I26364,I368684);
nor I_1392 (I26389,I26347,I26372);
DFFARX1 I_1393 (I26389,I2683,I26253,I26221,);
nand I_1394 (I26420,I26364,I368684);
nand I_1395 (I26437,I26287,I26420);
not I_1396 (I26233,I26437);
DFFARX1 I_1397 (I368672,I2683,I26253,I26477,);
DFFARX1 I_1398 (I26477,I2683,I26253,I26242,);
nand I_1399 (I26499,I368693,I368678);
and I_1400 (I26516,I26499,I368669);
DFFARX1 I_1401 (I26516,I2683,I26253,I26542,);
DFFARX1 I_1402 (I26542,I2683,I26253,I26559,);
not I_1403 (I26245,I26559);
not I_1404 (I26581,I26542);
nand I_1405 (I26230,I26581,I26420);
nor I_1406 (I26612,I368687,I368678);
not I_1407 (I26629,I26612);
nor I_1408 (I26646,I26581,I26629);
nor I_1409 (I26663,I26287,I26646);
DFFARX1 I_1410 (I26663,I2683,I26253,I26239,);
nor I_1411 (I26694,I26347,I26629);
nor I_1412 (I26227,I26542,I26694);
nor I_1413 (I26236,I26477,I26612);
nor I_1414 (I26224,I26347,I26612);
not I_1415 (I26780,I2690);
DFFARX1 I_1416 (I72711,I2683,I26780,I26806,);
not I_1417 (I26814,I26806);
nand I_1418 (I26831,I72705,I72699);
and I_1419 (I26848,I26831,I72720);
DFFARX1 I_1420 (I26848,I2683,I26780,I26874,);
DFFARX1 I_1421 (I72717,I2683,I26780,I26891,);
and I_1422 (I26899,I26891,I72714);
nor I_1423 (I26916,I26874,I26899);
DFFARX1 I_1424 (I26916,I2683,I26780,I26748,);
nand I_1425 (I26947,I26891,I72714);
nand I_1426 (I26964,I26814,I26947);
not I_1427 (I26760,I26964);
DFFARX1 I_1428 (I72699,I2683,I26780,I27004,);
DFFARX1 I_1429 (I27004,I2683,I26780,I26769,);
nand I_1430 (I27026,I72702,I72702);
and I_1431 (I27043,I27026,I72723);
DFFARX1 I_1432 (I27043,I2683,I26780,I27069,);
DFFARX1 I_1433 (I27069,I2683,I26780,I27086,);
not I_1434 (I26772,I27086);
not I_1435 (I27108,I27069);
nand I_1436 (I26757,I27108,I26947);
nor I_1437 (I27139,I72708,I72702);
not I_1438 (I27156,I27139);
nor I_1439 (I27173,I27108,I27156);
nor I_1440 (I27190,I26814,I27173);
DFFARX1 I_1441 (I27190,I2683,I26780,I26766,);
nor I_1442 (I27221,I26874,I27156);
nor I_1443 (I26754,I27069,I27221);
nor I_1444 (I26763,I27004,I27139);
nor I_1445 (I26751,I26874,I27139);
not I_1446 (I27307,I2690);
DFFARX1 I_1447 (I234857,I2683,I27307,I27333,);
not I_1448 (I27341,I27333);
nand I_1449 (I27358,I234848,I234866);
and I_1450 (I27375,I27358,I234845);
DFFARX1 I_1451 (I27375,I2683,I27307,I27401,);
DFFARX1 I_1452 (I234848,I2683,I27307,I27418,);
and I_1453 (I27426,I27418,I234851);
nor I_1454 (I27443,I27401,I27426);
DFFARX1 I_1455 (I27443,I2683,I27307,I27275,);
nand I_1456 (I27474,I27418,I234851);
nand I_1457 (I27491,I27341,I27474);
not I_1458 (I27287,I27491);
DFFARX1 I_1459 (I234845,I2683,I27307,I27531,);
DFFARX1 I_1460 (I27531,I2683,I27307,I27296,);
nand I_1461 (I27553,I234863,I234854);
and I_1462 (I27570,I27553,I234869);
DFFARX1 I_1463 (I27570,I2683,I27307,I27596,);
DFFARX1 I_1464 (I27596,I2683,I27307,I27613,);
not I_1465 (I27299,I27613);
not I_1466 (I27635,I27596);
nand I_1467 (I27284,I27635,I27474);
nor I_1468 (I27666,I234860,I234854);
not I_1469 (I27683,I27666);
nor I_1470 (I27700,I27635,I27683);
nor I_1471 (I27717,I27341,I27700);
DFFARX1 I_1472 (I27717,I2683,I27307,I27293,);
nor I_1473 (I27748,I27401,I27683);
nor I_1474 (I27281,I27596,I27748);
nor I_1475 (I27290,I27531,I27666);
nor I_1476 (I27278,I27401,I27666);
not I_1477 (I27834,I2690);
DFFARX1 I_1478 (I323299,I2683,I27834,I27860,);
not I_1479 (I27868,I27860);
nand I_1480 (I27885,I323296,I323302);
and I_1481 (I27902,I27885,I323299);
DFFARX1 I_1482 (I27902,I2683,I27834,I27928,);
DFFARX1 I_1483 (I323302,I2683,I27834,I27945,);
and I_1484 (I27953,I27945,I323296);
nor I_1485 (I27970,I27928,I27953);
DFFARX1 I_1486 (I27970,I2683,I27834,I27802,);
nand I_1487 (I28001,I27945,I323296);
nand I_1488 (I28018,I27868,I28001);
not I_1489 (I27814,I28018);
DFFARX1 I_1490 (I323305,I2683,I27834,I28058,);
DFFARX1 I_1491 (I28058,I2683,I27834,I27823,);
nand I_1492 (I28080,I323308,I323317);
and I_1493 (I28097,I28080,I323311);
DFFARX1 I_1494 (I28097,I2683,I27834,I28123,);
DFFARX1 I_1495 (I28123,I2683,I27834,I28140,);
not I_1496 (I27826,I28140);
not I_1497 (I28162,I28123);
nand I_1498 (I27811,I28162,I28001);
nor I_1499 (I28193,I323314,I323317);
not I_1500 (I28210,I28193);
nor I_1501 (I28227,I28162,I28210);
nor I_1502 (I28244,I27868,I28227);
DFFARX1 I_1503 (I28244,I2683,I27834,I27820,);
nor I_1504 (I28275,I27928,I28210);
nor I_1505 (I27808,I28123,I28275);
nor I_1506 (I27817,I28058,I28193);
nor I_1507 (I27805,I27928,I28193);
not I_1508 (I28361,I2690);
DFFARX1 I_1509 (I100045,I2683,I28361,I28387,);
not I_1510 (I28395,I28387);
nand I_1511 (I28412,I100027,I100042);
and I_1512 (I28429,I28412,I100018);
DFFARX1 I_1513 (I28429,I2683,I28361,I28455,);
DFFARX1 I_1514 (I100021,I2683,I28361,I28472,);
and I_1515 (I28480,I28472,I100036);
nor I_1516 (I28497,I28455,I28480);
DFFARX1 I_1517 (I28497,I2683,I28361,I28329,);
nand I_1518 (I28528,I28472,I100036);
nand I_1519 (I28545,I28395,I28528);
not I_1520 (I28341,I28545);
DFFARX1 I_1521 (I100039,I2683,I28361,I28585,);
DFFARX1 I_1522 (I28585,I2683,I28361,I28350,);
nand I_1523 (I28607,I100018,I100030);
and I_1524 (I28624,I28607,I100024);
DFFARX1 I_1525 (I28624,I2683,I28361,I28650,);
DFFARX1 I_1526 (I28650,I2683,I28361,I28667,);
not I_1527 (I28353,I28667);
not I_1528 (I28689,I28650);
nand I_1529 (I28338,I28689,I28528);
nor I_1530 (I28720,I100033,I100030);
not I_1531 (I28737,I28720);
nor I_1532 (I28754,I28689,I28737);
nor I_1533 (I28771,I28395,I28754);
DFFARX1 I_1534 (I28771,I2683,I28361,I28347,);
nor I_1535 (I28802,I28455,I28737);
nor I_1536 (I28335,I28650,I28802);
nor I_1537 (I28344,I28585,I28720);
nor I_1538 (I28332,I28455,I28720);
not I_1539 (I28888,I2690);
DFFARX1 I_1540 (I246074,I2683,I28888,I28914,);
not I_1541 (I28922,I28914);
nand I_1542 (I28939,I246071,I246086);
and I_1543 (I28956,I28939,I246068);
DFFARX1 I_1544 (I28956,I2683,I28888,I28982,);
DFFARX1 I_1545 (I246065,I2683,I28888,I28999,);
and I_1546 (I29007,I28999,I246065);
nor I_1547 (I29024,I28982,I29007);
DFFARX1 I_1548 (I29024,I2683,I28888,I28856,);
nand I_1549 (I29055,I28999,I246065);
nand I_1550 (I29072,I28922,I29055);
not I_1551 (I28868,I29072);
DFFARX1 I_1552 (I246068,I2683,I28888,I29112,);
DFFARX1 I_1553 (I29112,I2683,I28888,I28877,);
nand I_1554 (I29134,I246080,I246071);
and I_1555 (I29151,I29134,I246083);
DFFARX1 I_1556 (I29151,I2683,I28888,I29177,);
DFFARX1 I_1557 (I29177,I2683,I28888,I29194,);
not I_1558 (I28880,I29194);
not I_1559 (I29216,I29177);
nand I_1560 (I28865,I29216,I29055);
nor I_1561 (I29247,I246077,I246071);
not I_1562 (I29264,I29247);
nor I_1563 (I29281,I29216,I29264);
nor I_1564 (I29298,I28922,I29281);
DFFARX1 I_1565 (I29298,I2683,I28888,I28874,);
nor I_1566 (I29329,I28982,I29264);
nor I_1567 (I28862,I29177,I29329);
nor I_1568 (I28871,I29112,I29247);
nor I_1569 (I28859,I28982,I29247);
not I_1570 (I29415,I2690);
DFFARX1 I_1571 (I168327,I2683,I29415,I29441,);
not I_1572 (I29449,I29441);
nand I_1573 (I29466,I168348,I168342);
and I_1574 (I29483,I29466,I168324);
DFFARX1 I_1575 (I29483,I2683,I29415,I29509,);
DFFARX1 I_1576 (I168327,I2683,I29415,I29526,);
and I_1577 (I29534,I29526,I168336);
nor I_1578 (I29551,I29509,I29534);
DFFARX1 I_1579 (I29551,I2683,I29415,I29383,);
nand I_1580 (I29582,I29526,I168336);
nand I_1581 (I29599,I29449,I29582);
not I_1582 (I29395,I29599);
DFFARX1 I_1583 (I168333,I2683,I29415,I29639,);
DFFARX1 I_1584 (I29639,I2683,I29415,I29404,);
nand I_1585 (I29661,I168339,I168330);
and I_1586 (I29678,I29661,I168324);
DFFARX1 I_1587 (I29678,I2683,I29415,I29704,);
DFFARX1 I_1588 (I29704,I2683,I29415,I29721,);
not I_1589 (I29407,I29721);
not I_1590 (I29743,I29704);
nand I_1591 (I29392,I29743,I29582);
nor I_1592 (I29774,I168345,I168330);
not I_1593 (I29791,I29774);
nor I_1594 (I29808,I29743,I29791);
nor I_1595 (I29825,I29449,I29808);
DFFARX1 I_1596 (I29825,I2683,I29415,I29401,);
nor I_1597 (I29856,I29509,I29791);
nor I_1598 (I29389,I29704,I29856);
nor I_1599 (I29398,I29639,I29774);
nor I_1600 (I29386,I29509,I29774);
not I_1601 (I29942,I2690);
DFFARX1 I_1602 (I44160,I2683,I29942,I29968,);
not I_1603 (I29976,I29968);
nand I_1604 (I29993,I44157,I44139);
and I_1605 (I30010,I29993,I44145);
DFFARX1 I_1606 (I30010,I2683,I29942,I30036,);
DFFARX1 I_1607 (I44154,I2683,I29942,I30053,);
and I_1608 (I30061,I30053,I44148);
nor I_1609 (I30078,I30036,I30061);
DFFARX1 I_1610 (I30078,I2683,I29942,I29910,);
nand I_1611 (I30109,I30053,I44148);
nand I_1612 (I30126,I29976,I30109);
not I_1613 (I29922,I30126);
DFFARX1 I_1614 (I44163,I2683,I29942,I30166,);
DFFARX1 I_1615 (I30166,I2683,I29942,I29931,);
nand I_1616 (I30188,I44151,I44142);
and I_1617 (I30205,I30188,I44139);
DFFARX1 I_1618 (I30205,I2683,I29942,I30231,);
DFFARX1 I_1619 (I30231,I2683,I29942,I30248,);
not I_1620 (I29934,I30248);
not I_1621 (I30270,I30231);
nand I_1622 (I29919,I30270,I30109);
nor I_1623 (I30301,I44166,I44142);
not I_1624 (I30318,I30301);
nor I_1625 (I30335,I30270,I30318);
nor I_1626 (I30352,I29976,I30335);
DFFARX1 I_1627 (I30352,I2683,I29942,I29928,);
nor I_1628 (I30383,I30036,I30318);
nor I_1629 (I29916,I30231,I30383);
nor I_1630 (I29925,I30166,I30301);
nor I_1631 (I29913,I30036,I30301);
not I_1632 (I30469,I2690);
DFFARX1 I_1633 (I84016,I2683,I30469,I30495,);
not I_1634 (I30503,I30495);
nand I_1635 (I30520,I84010,I84004);
and I_1636 (I30537,I30520,I84025);
DFFARX1 I_1637 (I30537,I2683,I30469,I30563,);
DFFARX1 I_1638 (I84022,I2683,I30469,I30580,);
and I_1639 (I30588,I30580,I84019);
nor I_1640 (I30605,I30563,I30588);
DFFARX1 I_1641 (I30605,I2683,I30469,I30437,);
nand I_1642 (I30636,I30580,I84019);
nand I_1643 (I30653,I30503,I30636);
not I_1644 (I30449,I30653);
DFFARX1 I_1645 (I84004,I2683,I30469,I30693,);
DFFARX1 I_1646 (I30693,I2683,I30469,I30458,);
nand I_1647 (I30715,I84007,I84007);
and I_1648 (I30732,I30715,I84028);
DFFARX1 I_1649 (I30732,I2683,I30469,I30758,);
DFFARX1 I_1650 (I30758,I2683,I30469,I30775,);
not I_1651 (I30461,I30775);
not I_1652 (I30797,I30758);
nand I_1653 (I30446,I30797,I30636);
nor I_1654 (I30828,I84013,I84007);
not I_1655 (I30845,I30828);
nor I_1656 (I30862,I30797,I30845);
nor I_1657 (I30879,I30503,I30862);
DFFARX1 I_1658 (I30879,I2683,I30469,I30455,);
nor I_1659 (I30910,I30563,I30845);
nor I_1660 (I30443,I30758,I30910);
nor I_1661 (I30452,I30693,I30828);
nor I_1662 (I30440,I30563,I30828);
not I_1663 (I30996,I2690);
DFFARX1 I_1664 (I224453,I2683,I30996,I31022,);
not I_1665 (I31030,I31022);
nand I_1666 (I31047,I224444,I224462);
and I_1667 (I31064,I31047,I224441);
DFFARX1 I_1668 (I31064,I2683,I30996,I31090,);
DFFARX1 I_1669 (I224444,I2683,I30996,I31107,);
and I_1670 (I31115,I31107,I224447);
nor I_1671 (I31132,I31090,I31115);
DFFARX1 I_1672 (I31132,I2683,I30996,I30964,);
nand I_1673 (I31163,I31107,I224447);
nand I_1674 (I31180,I31030,I31163);
not I_1675 (I30976,I31180);
DFFARX1 I_1676 (I224441,I2683,I30996,I31220,);
DFFARX1 I_1677 (I31220,I2683,I30996,I30985,);
nand I_1678 (I31242,I224459,I224450);
and I_1679 (I31259,I31242,I224465);
DFFARX1 I_1680 (I31259,I2683,I30996,I31285,);
DFFARX1 I_1681 (I31285,I2683,I30996,I31302,);
not I_1682 (I30988,I31302);
not I_1683 (I31324,I31285);
nand I_1684 (I30973,I31324,I31163);
nor I_1685 (I31355,I224456,I224450);
not I_1686 (I31372,I31355);
nor I_1687 (I31389,I31324,I31372);
nor I_1688 (I31406,I31030,I31389);
DFFARX1 I_1689 (I31406,I2683,I30996,I30982,);
nor I_1690 (I31437,I31090,I31372);
nor I_1691 (I30970,I31285,I31437);
nor I_1692 (I30979,I31220,I31355);
nor I_1693 (I30967,I31090,I31355);
not I_1694 (I31523,I2690);
DFFARX1 I_1695 (I258722,I2683,I31523,I31549,);
not I_1696 (I31557,I31549);
nand I_1697 (I31574,I258719,I258734);
and I_1698 (I31591,I31574,I258716);
DFFARX1 I_1699 (I31591,I2683,I31523,I31617,);
DFFARX1 I_1700 (I258713,I2683,I31523,I31634,);
and I_1701 (I31642,I31634,I258713);
nor I_1702 (I31659,I31617,I31642);
DFFARX1 I_1703 (I31659,I2683,I31523,I31491,);
nand I_1704 (I31690,I31634,I258713);
nand I_1705 (I31707,I31557,I31690);
not I_1706 (I31503,I31707);
DFFARX1 I_1707 (I258716,I2683,I31523,I31747,);
DFFARX1 I_1708 (I31747,I2683,I31523,I31512,);
nand I_1709 (I31769,I258728,I258719);
and I_1710 (I31786,I31769,I258731);
DFFARX1 I_1711 (I31786,I2683,I31523,I31812,);
DFFARX1 I_1712 (I31812,I2683,I31523,I31829,);
not I_1713 (I31515,I31829);
not I_1714 (I31851,I31812);
nand I_1715 (I31500,I31851,I31690);
nor I_1716 (I31882,I258725,I258719);
not I_1717 (I31899,I31882);
nor I_1718 (I31916,I31851,I31899);
nor I_1719 (I31933,I31557,I31916);
DFFARX1 I_1720 (I31933,I2683,I31523,I31509,);
nor I_1721 (I31964,I31617,I31899);
nor I_1722 (I31497,I31812,I31964);
nor I_1723 (I31506,I31747,I31882);
nor I_1724 (I31494,I31617,I31882);
not I_1725 (I32050,I2690);
DFFARX1 I_1726 (I242912,I2683,I32050,I32076,);
not I_1727 (I32084,I32076);
nand I_1728 (I32101,I242909,I242924);
and I_1729 (I32118,I32101,I242906);
DFFARX1 I_1730 (I32118,I2683,I32050,I32144,);
DFFARX1 I_1731 (I242903,I2683,I32050,I32161,);
and I_1732 (I32169,I32161,I242903);
nor I_1733 (I32186,I32144,I32169);
DFFARX1 I_1734 (I32186,I2683,I32050,I32018,);
nand I_1735 (I32217,I32161,I242903);
nand I_1736 (I32234,I32084,I32217);
not I_1737 (I32030,I32234);
DFFARX1 I_1738 (I242906,I2683,I32050,I32274,);
DFFARX1 I_1739 (I32274,I2683,I32050,I32039,);
nand I_1740 (I32296,I242918,I242909);
and I_1741 (I32313,I32296,I242921);
DFFARX1 I_1742 (I32313,I2683,I32050,I32339,);
DFFARX1 I_1743 (I32339,I2683,I32050,I32356,);
not I_1744 (I32042,I32356);
not I_1745 (I32378,I32339);
nand I_1746 (I32027,I32378,I32217);
nor I_1747 (I32409,I242915,I242909);
not I_1748 (I32426,I32409);
nor I_1749 (I32443,I32378,I32426);
nor I_1750 (I32460,I32084,I32443);
DFFARX1 I_1751 (I32460,I2683,I32050,I32036,);
nor I_1752 (I32491,I32144,I32426);
nor I_1753 (I32024,I32339,I32491);
nor I_1754 (I32033,I32274,I32409);
nor I_1755 (I32021,I32144,I32409);
not I_1756 (I32577,I2690);
DFFARX1 I_1757 (I183990,I2683,I32577,I32603,);
not I_1758 (I32611,I32603);
nand I_1759 (I32628,I184002,I183987);
and I_1760 (I32645,I32628,I183981);
DFFARX1 I_1761 (I32645,I2683,I32577,I32671,);
DFFARX1 I_1762 (I183996,I2683,I32577,I32688,);
and I_1763 (I32696,I32688,I183984);
nor I_1764 (I32713,I32671,I32696);
DFFARX1 I_1765 (I32713,I2683,I32577,I32545,);
nand I_1766 (I32744,I32688,I183984);
nand I_1767 (I32761,I32611,I32744);
not I_1768 (I32557,I32761);
DFFARX1 I_1769 (I183993,I2683,I32577,I32801,);
DFFARX1 I_1770 (I32801,I2683,I32577,I32566,);
nand I_1771 (I32823,I183999,I184005);
and I_1772 (I32840,I32823,I183981);
DFFARX1 I_1773 (I32840,I2683,I32577,I32866,);
DFFARX1 I_1774 (I32866,I2683,I32577,I32883,);
not I_1775 (I32569,I32883);
not I_1776 (I32905,I32866);
nand I_1777 (I32554,I32905,I32744);
nor I_1778 (I32936,I183984,I184005);
not I_1779 (I32953,I32936);
nor I_1780 (I32970,I32905,I32953);
nor I_1781 (I32987,I32611,I32970);
DFFARX1 I_1782 (I32987,I2683,I32577,I32563,);
nor I_1783 (I33018,I32671,I32953);
nor I_1784 (I32551,I32866,I33018);
nor I_1785 (I32560,I32801,I32936);
nor I_1786 (I32548,I32671,I32936);
not I_1787 (I33104,I2690);
DFFARX1 I_1788 (I196131,I2683,I33104,I33130,);
not I_1789 (I33138,I33130);
nand I_1790 (I33155,I196122,I196140);
and I_1791 (I33172,I33155,I196119);
DFFARX1 I_1792 (I33172,I2683,I33104,I33198,);
DFFARX1 I_1793 (I196122,I2683,I33104,I33215,);
and I_1794 (I33223,I33215,I196125);
nor I_1795 (I33240,I33198,I33223);
DFFARX1 I_1796 (I33240,I2683,I33104,I33072,);
nand I_1797 (I33271,I33215,I196125);
nand I_1798 (I33288,I33138,I33271);
not I_1799 (I33084,I33288);
DFFARX1 I_1800 (I196119,I2683,I33104,I33328,);
DFFARX1 I_1801 (I33328,I2683,I33104,I33093,);
nand I_1802 (I33350,I196137,I196128);
and I_1803 (I33367,I33350,I196143);
DFFARX1 I_1804 (I33367,I2683,I33104,I33393,);
DFFARX1 I_1805 (I33393,I2683,I33104,I33410,);
not I_1806 (I33096,I33410);
not I_1807 (I33432,I33393);
nand I_1808 (I33081,I33432,I33271);
nor I_1809 (I33463,I196134,I196128);
not I_1810 (I33480,I33463);
nor I_1811 (I33497,I33432,I33480);
nor I_1812 (I33514,I33138,I33497);
DFFARX1 I_1813 (I33514,I2683,I33104,I33090,);
nor I_1814 (I33545,I33198,I33480);
nor I_1815 (I33078,I33393,I33545);
nor I_1816 (I33087,I33328,I33463);
nor I_1817 (I33075,I33198,I33463);
not I_1818 (I33631,I2690);
DFFARX1 I_1819 (I396816,I2683,I33631,I33657,);
not I_1820 (I33665,I33657);
nand I_1821 (I33682,I396810,I396831);
and I_1822 (I33699,I33682,I396807);
DFFARX1 I_1823 (I33699,I2683,I33631,I33725,);
DFFARX1 I_1824 (I396828,I2683,I33631,I33742,);
and I_1825 (I33750,I33742,I396825);
nor I_1826 (I33767,I33725,I33750);
DFFARX1 I_1827 (I33767,I2683,I33631,I33599,);
nand I_1828 (I33798,I33742,I396825);
nand I_1829 (I33815,I33665,I33798);
not I_1830 (I33611,I33815);
DFFARX1 I_1831 (I396813,I2683,I33631,I33855,);
DFFARX1 I_1832 (I33855,I2683,I33631,I33620,);
nand I_1833 (I33877,I396822,I396819);
and I_1834 (I33894,I33877,I396804);
DFFARX1 I_1835 (I33894,I2683,I33631,I33920,);
DFFARX1 I_1836 (I33920,I2683,I33631,I33937,);
not I_1837 (I33623,I33937);
not I_1838 (I33959,I33920);
nand I_1839 (I33608,I33959,I33798);
nor I_1840 (I33990,I396804,I396819);
not I_1841 (I34007,I33990);
nor I_1842 (I34024,I33959,I34007);
nor I_1843 (I34041,I33665,I34024);
DFFARX1 I_1844 (I34041,I2683,I33631,I33617,);
nor I_1845 (I34072,I33725,I34007);
nor I_1846 (I33605,I33920,I34072);
nor I_1847 (I33614,I33855,I33990);
nor I_1848 (I33602,I33725,I33990);
not I_1849 (I34158,I2690);
DFFARX1 I_1850 (I291753,I2683,I34158,I34184,);
not I_1851 (I34192,I34184);
nand I_1852 (I34209,I291771,I291765);
and I_1853 (I34226,I34209,I291744);
DFFARX1 I_1854 (I34226,I2683,I34158,I34252,);
DFFARX1 I_1855 (I291762,I2683,I34158,I34269,);
and I_1856 (I34277,I34269,I291747);
nor I_1857 (I34294,I34252,I34277);
DFFARX1 I_1858 (I34294,I2683,I34158,I34126,);
nand I_1859 (I34325,I34269,I291747);
nand I_1860 (I34342,I34192,I34325);
not I_1861 (I34138,I34342);
DFFARX1 I_1862 (I291759,I2683,I34158,I34382,);
DFFARX1 I_1863 (I34382,I2683,I34158,I34147,);
nand I_1864 (I34404,I291768,I291756);
and I_1865 (I34421,I34404,I291750);
DFFARX1 I_1866 (I34421,I2683,I34158,I34447,);
DFFARX1 I_1867 (I34447,I2683,I34158,I34464,);
not I_1868 (I34150,I34464);
not I_1869 (I34486,I34447);
nand I_1870 (I34135,I34486,I34325);
nor I_1871 (I34517,I291744,I291756);
not I_1872 (I34534,I34517);
nor I_1873 (I34551,I34486,I34534);
nor I_1874 (I34568,I34192,I34551);
DFFARX1 I_1875 (I34568,I2683,I34158,I34144,);
nor I_1876 (I34599,I34252,I34534);
nor I_1877 (I34132,I34447,I34599);
nor I_1878 (I34141,I34382,I34517);
nor I_1879 (I34129,I34252,I34517);
not I_1880 (I34685,I2690);
DFFARX1 I_1881 (I342937,I2683,I34685,I34711,);
not I_1882 (I34719,I34711);
nand I_1883 (I34736,I342952,I342931);
and I_1884 (I34753,I34736,I342934);
DFFARX1 I_1885 (I34753,I2683,I34685,I34779,);
DFFARX1 I_1886 (I342955,I2683,I34685,I34796,);
and I_1887 (I34804,I34796,I342934);
nor I_1888 (I34821,I34779,I34804);
DFFARX1 I_1889 (I34821,I2683,I34685,I34653,);
nand I_1890 (I34852,I34796,I342934);
nand I_1891 (I34869,I34719,I34852);
not I_1892 (I34665,I34869);
DFFARX1 I_1893 (I342931,I2683,I34685,I34909,);
DFFARX1 I_1894 (I34909,I2683,I34685,I34674,);
nand I_1895 (I34931,I342943,I342940);
and I_1896 (I34948,I34931,I342946);
DFFARX1 I_1897 (I34948,I2683,I34685,I34974,);
DFFARX1 I_1898 (I34974,I2683,I34685,I34991,);
not I_1899 (I34677,I34991);
not I_1900 (I35013,I34974);
nand I_1901 (I34662,I35013,I34852);
nor I_1902 (I35044,I342949,I342940);
not I_1903 (I35061,I35044);
nor I_1904 (I35078,I35013,I35061);
nor I_1905 (I35095,I34719,I35078);
DFFARX1 I_1906 (I35095,I2683,I34685,I34671,);
nor I_1907 (I35126,I34779,I35061);
nor I_1908 (I34659,I34974,I35126);
nor I_1909 (I34668,I34909,I35044);
nor I_1910 (I34656,I34779,I35044);
not I_1911 (I35212,I2690);
DFFARX1 I_1912 (I244493,I2683,I35212,I35238,);
not I_1913 (I35246,I35238);
nand I_1914 (I35263,I244490,I244505);
and I_1915 (I35280,I35263,I244487);
DFFARX1 I_1916 (I35280,I2683,I35212,I35306,);
DFFARX1 I_1917 (I244484,I2683,I35212,I35323,);
and I_1918 (I35331,I35323,I244484);
nor I_1919 (I35348,I35306,I35331);
DFFARX1 I_1920 (I35348,I2683,I35212,I35180,);
nand I_1921 (I35379,I35323,I244484);
nand I_1922 (I35396,I35246,I35379);
not I_1923 (I35192,I35396);
DFFARX1 I_1924 (I244487,I2683,I35212,I35436,);
DFFARX1 I_1925 (I35436,I2683,I35212,I35201,);
nand I_1926 (I35458,I244499,I244490);
and I_1927 (I35475,I35458,I244502);
DFFARX1 I_1928 (I35475,I2683,I35212,I35501,);
DFFARX1 I_1929 (I35501,I2683,I35212,I35518,);
not I_1930 (I35204,I35518);
not I_1931 (I35540,I35501);
nand I_1932 (I35189,I35540,I35379);
nor I_1933 (I35571,I244496,I244490);
not I_1934 (I35588,I35571);
nor I_1935 (I35605,I35540,I35588);
nor I_1936 (I35622,I35246,I35605);
DFFARX1 I_1937 (I35622,I2683,I35212,I35198,);
nor I_1938 (I35653,I35306,I35588);
nor I_1939 (I35186,I35501,I35653);
nor I_1940 (I35195,I35436,I35571);
nor I_1941 (I35183,I35306,I35571);
not I_1942 (I35739,I2690);
DFFARX1 I_1943 (I269789,I2683,I35739,I35765,);
not I_1944 (I35773,I35765);
nand I_1945 (I35790,I269807,I269801);
and I_1946 (I35807,I35790,I269780);
DFFARX1 I_1947 (I35807,I2683,I35739,I35833,);
DFFARX1 I_1948 (I269798,I2683,I35739,I35850,);
and I_1949 (I35858,I35850,I269783);
nor I_1950 (I35875,I35833,I35858);
DFFARX1 I_1951 (I35875,I2683,I35739,I35707,);
nand I_1952 (I35906,I35850,I269783);
nand I_1953 (I35923,I35773,I35906);
not I_1954 (I35719,I35923);
DFFARX1 I_1955 (I269795,I2683,I35739,I35963,);
DFFARX1 I_1956 (I35963,I2683,I35739,I35728,);
nand I_1957 (I35985,I269804,I269792);
and I_1958 (I36002,I35985,I269786);
DFFARX1 I_1959 (I36002,I2683,I35739,I36028,);
DFFARX1 I_1960 (I36028,I2683,I35739,I36045,);
not I_1961 (I35731,I36045);
not I_1962 (I36067,I36028);
nand I_1963 (I35716,I36067,I35906);
nor I_1964 (I36098,I269780,I269792);
not I_1965 (I36115,I36098);
nor I_1966 (I36132,I36067,I36115);
nor I_1967 (I36149,I35773,I36132);
DFFARX1 I_1968 (I36149,I2683,I35739,I35725,);
nor I_1969 (I36180,I35833,I36115);
nor I_1970 (I35713,I36028,I36180);
nor I_1971 (I35722,I35963,I36098);
nor I_1972 (I35710,I35833,I36098);
not I_1973 (I36266,I2690);
DFFARX1 I_1974 (I64381,I2683,I36266,I36292,);
not I_1975 (I36300,I36292);
nand I_1976 (I36317,I64375,I64369);
and I_1977 (I36334,I36317,I64390);
DFFARX1 I_1978 (I36334,I2683,I36266,I36360,);
DFFARX1 I_1979 (I64387,I2683,I36266,I36377,);
and I_1980 (I36385,I36377,I64384);
nor I_1981 (I36402,I36360,I36385);
DFFARX1 I_1982 (I36402,I2683,I36266,I36234,);
nand I_1983 (I36433,I36377,I64384);
nand I_1984 (I36450,I36300,I36433);
not I_1985 (I36246,I36450);
DFFARX1 I_1986 (I64369,I2683,I36266,I36490,);
DFFARX1 I_1987 (I36490,I2683,I36266,I36255,);
nand I_1988 (I36512,I64372,I64372);
and I_1989 (I36529,I36512,I64393);
DFFARX1 I_1990 (I36529,I2683,I36266,I36555,);
DFFARX1 I_1991 (I36555,I2683,I36266,I36572,);
not I_1992 (I36258,I36572);
not I_1993 (I36594,I36555);
nand I_1994 (I36243,I36594,I36433);
nor I_1995 (I36625,I64378,I64372);
not I_1996 (I36642,I36625);
nor I_1997 (I36659,I36594,I36642);
nor I_1998 (I36676,I36300,I36659);
DFFARX1 I_1999 (I36676,I2683,I36266,I36252,);
nor I_2000 (I36707,I36360,I36642);
nor I_2001 (I36240,I36555,I36707);
nor I_2002 (I36249,I36490,I36625);
nor I_2003 (I36237,I36360,I36625);
not I_2004 (I36793,I2690);
DFFARX1 I_2005 (I174742,I2683,I36793,I36819,);
not I_2006 (I36827,I36819);
nand I_2007 (I36844,I174754,I174739);
and I_2008 (I36861,I36844,I174733);
DFFARX1 I_2009 (I36861,I2683,I36793,I36887,);
DFFARX1 I_2010 (I174748,I2683,I36793,I36904,);
and I_2011 (I36912,I36904,I174736);
nor I_2012 (I36929,I36887,I36912);
DFFARX1 I_2013 (I36929,I2683,I36793,I36761,);
nand I_2014 (I36960,I36904,I174736);
nand I_2015 (I36977,I36827,I36960);
not I_2016 (I36773,I36977);
DFFARX1 I_2017 (I174745,I2683,I36793,I37017,);
DFFARX1 I_2018 (I37017,I2683,I36793,I36782,);
nand I_2019 (I37039,I174751,I174757);
and I_2020 (I37056,I37039,I174733);
DFFARX1 I_2021 (I37056,I2683,I36793,I37082,);
DFFARX1 I_2022 (I37082,I2683,I36793,I37099,);
not I_2023 (I36785,I37099);
not I_2024 (I37121,I37082);
nand I_2025 (I36770,I37121,I36960);
nor I_2026 (I37152,I174736,I174757);
not I_2027 (I37169,I37152);
nor I_2028 (I37186,I37121,I37169);
nor I_2029 (I37203,I36827,I37186);
DFFARX1 I_2030 (I37203,I2683,I36793,I36779,);
nor I_2031 (I37234,I36887,I37169);
nor I_2032 (I36767,I37082,I37234);
nor I_2033 (I36776,I37017,I37152);
nor I_2034 (I36764,I36887,I37152);
not I_2035 (I37320,I2690);
DFFARX1 I_2036 (I201333,I2683,I37320,I37346,);
not I_2037 (I37354,I37346);
nand I_2038 (I37371,I201324,I201342);
and I_2039 (I37388,I37371,I201321);
DFFARX1 I_2040 (I37388,I2683,I37320,I37414,);
DFFARX1 I_2041 (I201324,I2683,I37320,I37431,);
and I_2042 (I37439,I37431,I201327);
nor I_2043 (I37456,I37414,I37439);
DFFARX1 I_2044 (I37456,I2683,I37320,I37288,);
nand I_2045 (I37487,I37431,I201327);
nand I_2046 (I37504,I37354,I37487);
not I_2047 (I37300,I37504);
DFFARX1 I_2048 (I201321,I2683,I37320,I37544,);
DFFARX1 I_2049 (I37544,I2683,I37320,I37309,);
nand I_2050 (I37566,I201339,I201330);
and I_2051 (I37583,I37566,I201345);
DFFARX1 I_2052 (I37583,I2683,I37320,I37609,);
DFFARX1 I_2053 (I37609,I2683,I37320,I37626,);
not I_2054 (I37312,I37626);
not I_2055 (I37648,I37609);
nand I_2056 (I37297,I37648,I37487);
nor I_2057 (I37679,I201336,I201330);
not I_2058 (I37696,I37679);
nor I_2059 (I37713,I37648,I37696);
nor I_2060 (I37730,I37354,I37713);
DFFARX1 I_2061 (I37730,I2683,I37320,I37306,);
nor I_2062 (I37761,I37414,I37696);
nor I_2063 (I37294,I37609,I37761);
nor I_2064 (I37303,I37544,I37679);
nor I_2065 (I37291,I37414,I37679);
not I_2066 (I37847,I2690);
DFFARX1 I_2067 (I258195,I2683,I37847,I37873,);
not I_2068 (I37881,I37873);
nand I_2069 (I37898,I258192,I258207);
and I_2070 (I37915,I37898,I258189);
DFFARX1 I_2071 (I37915,I2683,I37847,I37941,);
DFFARX1 I_2072 (I258186,I2683,I37847,I37958,);
and I_2073 (I37966,I37958,I258186);
nor I_2074 (I37983,I37941,I37966);
DFFARX1 I_2075 (I37983,I2683,I37847,I37815,);
nand I_2076 (I38014,I37958,I258186);
nand I_2077 (I38031,I37881,I38014);
not I_2078 (I37827,I38031);
DFFARX1 I_2079 (I258189,I2683,I37847,I38071,);
DFFARX1 I_2080 (I38071,I2683,I37847,I37836,);
nand I_2081 (I38093,I258201,I258192);
and I_2082 (I38110,I38093,I258204);
DFFARX1 I_2083 (I38110,I2683,I37847,I38136,);
DFFARX1 I_2084 (I38136,I2683,I37847,I38153,);
not I_2085 (I37839,I38153);
not I_2086 (I38175,I38136);
nand I_2087 (I37824,I38175,I38014);
nor I_2088 (I38206,I258198,I258192);
not I_2089 (I38223,I38206);
nor I_2090 (I38240,I38175,I38223);
nor I_2091 (I38257,I37881,I38240);
DFFARX1 I_2092 (I38257,I2683,I37847,I37833,);
nor I_2093 (I38288,I37941,I38223);
nor I_2094 (I37821,I38136,I38288);
nor I_2095 (I37830,I38071,I38206);
nor I_2096 (I37818,I37941,I38206);
not I_2097 (I38374,I2690);
DFFARX1 I_2098 (I122179,I2683,I38374,I38400,);
not I_2099 (I38408,I38400);
nand I_2100 (I38425,I122161,I122176);
and I_2101 (I38442,I38425,I122152);
DFFARX1 I_2102 (I38442,I2683,I38374,I38468,);
DFFARX1 I_2103 (I122155,I2683,I38374,I38485,);
and I_2104 (I38493,I38485,I122170);
nor I_2105 (I38510,I38468,I38493);
DFFARX1 I_2106 (I38510,I2683,I38374,I38342,);
nand I_2107 (I38541,I38485,I122170);
nand I_2108 (I38558,I38408,I38541);
not I_2109 (I38354,I38558);
DFFARX1 I_2110 (I122173,I2683,I38374,I38598,);
DFFARX1 I_2111 (I38598,I2683,I38374,I38363,);
nand I_2112 (I38620,I122152,I122164);
and I_2113 (I38637,I38620,I122158);
DFFARX1 I_2114 (I38637,I2683,I38374,I38663,);
DFFARX1 I_2115 (I38663,I2683,I38374,I38680,);
not I_2116 (I38366,I38680);
not I_2117 (I38702,I38663);
nand I_2118 (I38351,I38702,I38541);
nor I_2119 (I38733,I122167,I122164);
not I_2120 (I38750,I38733);
nor I_2121 (I38767,I38702,I38750);
nor I_2122 (I38784,I38408,I38767);
DFFARX1 I_2123 (I38784,I2683,I38374,I38360,);
nor I_2124 (I38815,I38468,I38750);
nor I_2125 (I38348,I38663,I38815);
nor I_2126 (I38357,I38598,I38733);
nor I_2127 (I38345,I38468,I38733);
not I_2128 (I38901,I2690);
DFFARX1 I_2129 (I376835,I2683,I38901,I38927,);
not I_2130 (I38935,I38927);
nand I_2131 (I38952,I376829,I376850);
and I_2132 (I38969,I38952,I376841);
DFFARX1 I_2133 (I38969,I2683,I38901,I38995,);
DFFARX1 I_2134 (I376832,I2683,I38901,I39012,);
and I_2135 (I39020,I39012,I376844);
nor I_2136 (I39037,I38995,I39020);
DFFARX1 I_2137 (I39037,I2683,I38901,I38869,);
nand I_2138 (I39068,I39012,I376844);
nand I_2139 (I39085,I38935,I39068);
not I_2140 (I38881,I39085);
DFFARX1 I_2141 (I376832,I2683,I38901,I39125,);
DFFARX1 I_2142 (I39125,I2683,I38901,I38890,);
nand I_2143 (I39147,I376853,I376838);
and I_2144 (I39164,I39147,I376829);
DFFARX1 I_2145 (I39164,I2683,I38901,I39190,);
DFFARX1 I_2146 (I39190,I2683,I38901,I39207,);
not I_2147 (I38893,I39207);
not I_2148 (I39229,I39190);
nand I_2149 (I38878,I39229,I39068);
nor I_2150 (I39260,I376847,I376838);
not I_2151 (I39277,I39260);
nor I_2152 (I39294,I39229,I39277);
nor I_2153 (I39311,I38935,I39294);
DFFARX1 I_2154 (I39311,I2683,I38901,I38887,);
nor I_2155 (I39342,I38995,I39277);
nor I_2156 (I38875,I39190,I39342);
nor I_2157 (I38884,I39125,I39260);
nor I_2158 (I38872,I38995,I39260);
not I_2159 (I39428,I2690);
DFFARX1 I_2160 (I233701,I2683,I39428,I39454,);
not I_2161 (I39462,I39454);
nand I_2162 (I39479,I233692,I233710);
and I_2163 (I39496,I39479,I233689);
DFFARX1 I_2164 (I39496,I2683,I39428,I39522,);
DFFARX1 I_2165 (I233692,I2683,I39428,I39539,);
and I_2166 (I39547,I39539,I233695);
nor I_2167 (I39564,I39522,I39547);
DFFARX1 I_2168 (I39564,I2683,I39428,I39396,);
nand I_2169 (I39595,I39539,I233695);
nand I_2170 (I39612,I39462,I39595);
not I_2171 (I39408,I39612);
DFFARX1 I_2172 (I233689,I2683,I39428,I39652,);
DFFARX1 I_2173 (I39652,I2683,I39428,I39417,);
nand I_2174 (I39674,I233707,I233698);
and I_2175 (I39691,I39674,I233713);
DFFARX1 I_2176 (I39691,I2683,I39428,I39717,);
DFFARX1 I_2177 (I39717,I2683,I39428,I39734,);
not I_2178 (I39420,I39734);
not I_2179 (I39756,I39717);
nand I_2180 (I39405,I39756,I39595);
nor I_2181 (I39787,I233704,I233698);
not I_2182 (I39804,I39787);
nor I_2183 (I39821,I39756,I39804);
nor I_2184 (I39838,I39462,I39821);
DFFARX1 I_2185 (I39838,I2683,I39428,I39414,);
nor I_2186 (I39869,I39522,I39804);
nor I_2187 (I39402,I39717,I39869);
nor I_2188 (I39411,I39652,I39787);
nor I_2189 (I39399,I39522,I39787);
not I_2190 (I39955,I2690);
DFFARX1 I_2191 (I263465,I2683,I39955,I39981,);
not I_2192 (I39989,I39981);
nand I_2193 (I40006,I263462,I263477);
and I_2194 (I40023,I40006,I263459);
DFFARX1 I_2195 (I40023,I2683,I39955,I40049,);
DFFARX1 I_2196 (I263456,I2683,I39955,I40066,);
and I_2197 (I40074,I40066,I263456);
nor I_2198 (I40091,I40049,I40074);
DFFARX1 I_2199 (I40091,I2683,I39955,I39923,);
nand I_2200 (I40122,I40066,I263456);
nand I_2201 (I40139,I39989,I40122);
not I_2202 (I39935,I40139);
DFFARX1 I_2203 (I263459,I2683,I39955,I40179,);
DFFARX1 I_2204 (I40179,I2683,I39955,I39944,);
nand I_2205 (I40201,I263471,I263462);
and I_2206 (I40218,I40201,I263474);
DFFARX1 I_2207 (I40218,I2683,I39955,I40244,);
DFFARX1 I_2208 (I40244,I2683,I39955,I40261,);
not I_2209 (I39947,I40261);
not I_2210 (I40283,I40244);
nand I_2211 (I39932,I40283,I40122);
nor I_2212 (I40314,I263468,I263462);
not I_2213 (I40331,I40314);
nor I_2214 (I40348,I40283,I40331);
nor I_2215 (I40365,I39989,I40348);
DFFARX1 I_2216 (I40365,I2683,I39955,I39941,);
nor I_2217 (I40396,I40049,I40331);
nor I_2218 (I39929,I40244,I40396);
nor I_2219 (I39938,I40179,I40314);
nor I_2220 (I39926,I40049,I40314);
not I_2221 (I40482,I2690);
DFFARX1 I_2222 (I209425,I2683,I40482,I40508,);
not I_2223 (I40516,I40508);
nand I_2224 (I40533,I209416,I209434);
and I_2225 (I40550,I40533,I209413);
DFFARX1 I_2226 (I40550,I2683,I40482,I40576,);
DFFARX1 I_2227 (I209416,I2683,I40482,I40593,);
and I_2228 (I40601,I40593,I209419);
nor I_2229 (I40618,I40576,I40601);
DFFARX1 I_2230 (I40618,I2683,I40482,I40450,);
nand I_2231 (I40649,I40593,I209419);
nand I_2232 (I40666,I40516,I40649);
not I_2233 (I40462,I40666);
DFFARX1 I_2234 (I209413,I2683,I40482,I40706,);
DFFARX1 I_2235 (I40706,I2683,I40482,I40471,);
nand I_2236 (I40728,I209431,I209422);
and I_2237 (I40745,I40728,I209437);
DFFARX1 I_2238 (I40745,I2683,I40482,I40771,);
DFFARX1 I_2239 (I40771,I2683,I40482,I40788,);
not I_2240 (I40474,I40788);
not I_2241 (I40810,I40771);
nand I_2242 (I40459,I40810,I40649);
nor I_2243 (I40841,I209428,I209422);
not I_2244 (I40858,I40841);
nor I_2245 (I40875,I40810,I40858);
nor I_2246 (I40892,I40516,I40875);
DFFARX1 I_2247 (I40892,I2683,I40482,I40468,);
nor I_2248 (I40923,I40576,I40858);
nor I_2249 (I40456,I40771,I40923);
nor I_2250 (I40465,I40706,I40841);
nor I_2251 (I40453,I40576,I40841);
not I_2252 (I41009,I2690);
DFFARX1 I_2253 (I84611,I2683,I41009,I41035,);
not I_2254 (I41043,I41035);
nand I_2255 (I41060,I84605,I84599);
and I_2256 (I41077,I41060,I84620);
DFFARX1 I_2257 (I41077,I2683,I41009,I41103,);
DFFARX1 I_2258 (I84617,I2683,I41009,I41120,);
and I_2259 (I41128,I41120,I84614);
nor I_2260 (I41145,I41103,I41128);
DFFARX1 I_2261 (I41145,I2683,I41009,I40977,);
nand I_2262 (I41176,I41120,I84614);
nand I_2263 (I41193,I41043,I41176);
not I_2264 (I40989,I41193);
DFFARX1 I_2265 (I84599,I2683,I41009,I41233,);
DFFARX1 I_2266 (I41233,I2683,I41009,I40998,);
nand I_2267 (I41255,I84602,I84602);
and I_2268 (I41272,I41255,I84623);
DFFARX1 I_2269 (I41272,I2683,I41009,I41298,);
DFFARX1 I_2270 (I41298,I2683,I41009,I41315,);
not I_2271 (I41001,I41315);
not I_2272 (I41337,I41298);
nand I_2273 (I40986,I41337,I41176);
nor I_2274 (I41368,I84608,I84602);
not I_2275 (I41385,I41368);
nor I_2276 (I41402,I41337,I41385);
nor I_2277 (I41419,I41043,I41402);
DFFARX1 I_2278 (I41419,I2683,I41009,I40995,);
nor I_2279 (I41450,I41103,I41385);
nor I_2280 (I40983,I41298,I41450);
nor I_2281 (I40992,I41233,I41368);
nor I_2282 (I40980,I41103,I41368);
not I_2283 (I41536,I2690);
DFFARX1 I_2284 (I307903,I2683,I41536,I41562,);
not I_2285 (I41570,I41562);
nand I_2286 (I41587,I307921,I307915);
and I_2287 (I41604,I41587,I307894);
DFFARX1 I_2288 (I41604,I2683,I41536,I41630,);
DFFARX1 I_2289 (I307912,I2683,I41536,I41647,);
and I_2290 (I41655,I41647,I307897);
nor I_2291 (I41672,I41630,I41655);
DFFARX1 I_2292 (I41672,I2683,I41536,I41504,);
nand I_2293 (I41703,I41647,I307897);
nand I_2294 (I41720,I41570,I41703);
not I_2295 (I41516,I41720);
DFFARX1 I_2296 (I307909,I2683,I41536,I41760,);
DFFARX1 I_2297 (I41760,I2683,I41536,I41525,);
nand I_2298 (I41782,I307918,I307906);
and I_2299 (I41799,I41782,I307900);
DFFARX1 I_2300 (I41799,I2683,I41536,I41825,);
DFFARX1 I_2301 (I41825,I2683,I41536,I41842,);
not I_2302 (I41528,I41842);
not I_2303 (I41864,I41825);
nand I_2304 (I41513,I41864,I41703);
nor I_2305 (I41895,I307894,I307906);
not I_2306 (I41912,I41895);
nor I_2307 (I41929,I41864,I41912);
nor I_2308 (I41946,I41570,I41929);
DFFARX1 I_2309 (I41946,I2683,I41536,I41522,);
nor I_2310 (I41977,I41630,I41912);
nor I_2311 (I41510,I41825,I41977);
nor I_2312 (I41519,I41760,I41895);
nor I_2313 (I41507,I41630,I41895);
not I_2314 (I42063,I2690);
DFFARX1 I_2315 (I119544,I2683,I42063,I42089,);
not I_2316 (I42097,I42089);
nand I_2317 (I42114,I119526,I119541);
and I_2318 (I42131,I42114,I119517);
DFFARX1 I_2319 (I42131,I2683,I42063,I42157,);
DFFARX1 I_2320 (I119520,I2683,I42063,I42174,);
and I_2321 (I42182,I42174,I119535);
nor I_2322 (I42199,I42157,I42182);
DFFARX1 I_2323 (I42199,I2683,I42063,I42031,);
nand I_2324 (I42230,I42174,I119535);
nand I_2325 (I42247,I42097,I42230);
not I_2326 (I42043,I42247);
DFFARX1 I_2327 (I119538,I2683,I42063,I42287,);
DFFARX1 I_2328 (I42287,I2683,I42063,I42052,);
nand I_2329 (I42309,I119517,I119529);
and I_2330 (I42326,I42309,I119523);
DFFARX1 I_2331 (I42326,I2683,I42063,I42352,);
DFFARX1 I_2332 (I42352,I2683,I42063,I42369,);
not I_2333 (I42055,I42369);
not I_2334 (I42391,I42352);
nand I_2335 (I42040,I42391,I42230);
nor I_2336 (I42422,I119532,I119529);
not I_2337 (I42439,I42422);
nor I_2338 (I42456,I42391,I42439);
nor I_2339 (I42473,I42097,I42456);
DFFARX1 I_2340 (I42473,I2683,I42063,I42049,);
nor I_2341 (I42504,I42157,I42439);
nor I_2342 (I42037,I42352,I42504);
nor I_2343 (I42046,I42287,I42422);
nor I_2344 (I42034,I42157,I42422);
not I_2345 (I42590,I2690);
DFFARX1 I_2346 (I243966,I2683,I42590,I42616,);
not I_2347 (I42624,I42616);
nand I_2348 (I42641,I243963,I243978);
and I_2349 (I42658,I42641,I243960);
DFFARX1 I_2350 (I42658,I2683,I42590,I42684,);
DFFARX1 I_2351 (I243957,I2683,I42590,I42701,);
and I_2352 (I42709,I42701,I243957);
nor I_2353 (I42726,I42684,I42709);
DFFARX1 I_2354 (I42726,I2683,I42590,I42558,);
nand I_2355 (I42757,I42701,I243957);
nand I_2356 (I42774,I42624,I42757);
not I_2357 (I42570,I42774);
DFFARX1 I_2358 (I243960,I2683,I42590,I42814,);
DFFARX1 I_2359 (I42814,I2683,I42590,I42579,);
nand I_2360 (I42836,I243972,I243963);
and I_2361 (I42853,I42836,I243975);
DFFARX1 I_2362 (I42853,I2683,I42590,I42879,);
DFFARX1 I_2363 (I42879,I2683,I42590,I42896,);
not I_2364 (I42582,I42896);
not I_2365 (I42918,I42879);
nand I_2366 (I42567,I42918,I42757);
nor I_2367 (I42949,I243969,I243963);
not I_2368 (I42966,I42949);
nor I_2369 (I42983,I42918,I42966);
nor I_2370 (I43000,I42624,I42983);
DFFARX1 I_2371 (I43000,I2683,I42590,I42576,);
nor I_2372 (I43031,I42684,I42966);
nor I_2373 (I42564,I42879,I43031);
nor I_2374 (I42573,I42814,I42949);
nor I_2375 (I42561,I42684,I42949);
not I_2376 (I43117,I2690);
DFFARX1 I_2377 (I114801,I2683,I43117,I43143,);
not I_2378 (I43151,I43143);
nand I_2379 (I43168,I114783,I114798);
and I_2380 (I43185,I43168,I114774);
DFFARX1 I_2381 (I43185,I2683,I43117,I43211,);
DFFARX1 I_2382 (I114777,I2683,I43117,I43228,);
and I_2383 (I43236,I43228,I114792);
nor I_2384 (I43253,I43211,I43236);
DFFARX1 I_2385 (I43253,I2683,I43117,I43085,);
nand I_2386 (I43284,I43228,I114792);
nand I_2387 (I43301,I43151,I43284);
not I_2388 (I43097,I43301);
DFFARX1 I_2389 (I114795,I2683,I43117,I43341,);
DFFARX1 I_2390 (I43341,I2683,I43117,I43106,);
nand I_2391 (I43363,I114774,I114786);
and I_2392 (I43380,I43363,I114780);
DFFARX1 I_2393 (I43380,I2683,I43117,I43406,);
DFFARX1 I_2394 (I43406,I2683,I43117,I43423,);
not I_2395 (I43109,I43423);
not I_2396 (I43445,I43406);
nand I_2397 (I43094,I43445,I43284);
nor I_2398 (I43476,I114789,I114786);
not I_2399 (I43493,I43476);
nor I_2400 (I43510,I43445,I43493);
nor I_2401 (I43527,I43151,I43510);
DFFARX1 I_2402 (I43527,I2683,I43117,I43103,);
nor I_2403 (I43558,I43211,I43493);
nor I_2404 (I43091,I43406,I43558);
nor I_2405 (I43100,I43341,I43476);
nor I_2406 (I43088,I43211,I43476);
not I_2407 (I43644,I2690);
DFFARX1 I_2408 (I78066,I2683,I43644,I43670,);
not I_2409 (I43678,I43670);
nand I_2410 (I43695,I78060,I78054);
and I_2411 (I43712,I43695,I78075);
DFFARX1 I_2412 (I43712,I2683,I43644,I43738,);
DFFARX1 I_2413 (I78072,I2683,I43644,I43755,);
and I_2414 (I43763,I43755,I78069);
nor I_2415 (I43780,I43738,I43763);
DFFARX1 I_2416 (I43780,I2683,I43644,I43612,);
nand I_2417 (I43811,I43755,I78069);
nand I_2418 (I43828,I43678,I43811);
not I_2419 (I43624,I43828);
DFFARX1 I_2420 (I78054,I2683,I43644,I43868,);
DFFARX1 I_2421 (I43868,I2683,I43644,I43633,);
nand I_2422 (I43890,I78057,I78057);
and I_2423 (I43907,I43890,I78078);
DFFARX1 I_2424 (I43907,I2683,I43644,I43933,);
DFFARX1 I_2425 (I43933,I2683,I43644,I43950,);
not I_2426 (I43636,I43950);
not I_2427 (I43972,I43933);
nand I_2428 (I43621,I43972,I43811);
nor I_2429 (I44003,I78063,I78057);
not I_2430 (I44020,I44003);
nor I_2431 (I44037,I43972,I44020);
nor I_2432 (I44054,I43678,I44037);
DFFARX1 I_2433 (I44054,I2683,I43644,I43630,);
nor I_2434 (I44085,I43738,I44020);
nor I_2435 (I43618,I43933,I44085);
nor I_2436 (I43627,I43868,I44003);
nor I_2437 (I43615,I43738,I44003);
not I_2438 (I44174,I2690);
DFFARX1 I_2439 (I61418,I2683,I44174,I44200,);
not I_2440 (I44208,I44200);
DFFARX1 I_2441 (I61412,I2683,I44174,I44234,);
not I_2442 (I44242,I61397);
or I_2443 (I44259,I61406,I61397);
nor I_2444 (I44276,I44234,I61406);
nand I_2445 (I44151,I44242,I44276);
nor I_2446 (I44307,I61394,I61406);
nand I_2447 (I44145,I44307,I44242);
not I_2448 (I44338,I61400);
nand I_2449 (I44355,I44242,I44338);
nor I_2450 (I44372,I61403,I61415);
not I_2451 (I44389,I44372);
nor I_2452 (I44406,I44389,I44355);
nor I_2453 (I44423,I44307,I44406);
DFFARX1 I_2454 (I44423,I2683,I44174,I44160,);
nor I_2455 (I44157,I44372,I44259);
DFFARX1 I_2456 (I44372,I2683,I44174,I44163,);
nor I_2457 (I44482,I44338,I61403);
nor I_2458 (I44499,I44482,I61397);
nor I_2459 (I44516,I61409,I61397);
DFFARX1 I_2460 (I44516,I2683,I44174,I44542,);
nor I_2461 (I44142,I44542,I44499);
DFFARX1 I_2462 (I44542,I2683,I44174,I44573,);
nand I_2463 (I44581,I44573,I61394);
nor I_2464 (I44166,I44208,I44581);
not I_2465 (I44612,I44542);
nand I_2466 (I44629,I44612,I61394);
nor I_2467 (I44646,I44208,I44629);
nor I_2468 (I44148,I44234,I44646);
nor I_2469 (I44677,I61409,I61394);
nor I_2470 (I44694,I44234,I44677);
DFFARX1 I_2471 (I44694,I2683,I44174,I44139,);
and I_2472 (I44154,I44307,I61409);
not I_2473 (I44769,I2690);
DFFARX1 I_2474 (I248179,I2683,I44769,I44795,);
not I_2475 (I44803,I44795);
DFFARX1 I_2476 (I248179,I2683,I44769,I44829,);
not I_2477 (I44837,I248176);
or I_2478 (I44854,I248188,I248176);
nor I_2479 (I44871,I44829,I248188);
nand I_2480 (I44746,I44837,I44871);
nor I_2481 (I44902,I248182,I248188);
nand I_2482 (I44740,I44902,I44837);
not I_2483 (I44933,I248194);
nand I_2484 (I44950,I44837,I44933);
nor I_2485 (I44967,I248185,I248173);
not I_2486 (I44984,I44967);
nor I_2487 (I45001,I44984,I44950);
nor I_2488 (I45018,I44902,I45001);
DFFARX1 I_2489 (I45018,I2683,I44769,I44755,);
nor I_2490 (I44752,I44967,I44854);
DFFARX1 I_2491 (I44967,I2683,I44769,I44758,);
nor I_2492 (I45077,I44933,I248185);
nor I_2493 (I45094,I45077,I248176);
nor I_2494 (I45111,I248176,I248173);
DFFARX1 I_2495 (I45111,I2683,I44769,I45137,);
nor I_2496 (I44737,I45137,I45094);
DFFARX1 I_2497 (I45137,I2683,I44769,I45168,);
nand I_2498 (I45176,I45168,I248191);
nor I_2499 (I44761,I44803,I45176);
not I_2500 (I45207,I45137);
nand I_2501 (I45224,I45207,I248191);
nor I_2502 (I45241,I44803,I45224);
nor I_2503 (I44743,I44829,I45241);
nor I_2504 (I45272,I248176,I248182);
nor I_2505 (I45289,I44829,I45272);
DFFARX1 I_2506 (I45289,I2683,I44769,I44734,);
and I_2507 (I44749,I44902,I248176);
not I_2508 (I45364,I2690);
DFFARX1 I_2509 (I329062,I2683,I45364,I45390,);
not I_2510 (I45398,I45390);
DFFARX1 I_2511 (I329059,I2683,I45364,I45424,);
not I_2512 (I45432,I329068);
or I_2513 (I45449,I329059,I329068);
nor I_2514 (I45466,I45424,I329059);
nand I_2515 (I45341,I45432,I45466);
nor I_2516 (I45497,I329071,I329059);
nand I_2517 (I45335,I45497,I45432);
not I_2518 (I45528,I329065);
nand I_2519 (I45545,I45432,I45528);
nor I_2520 (I45562,I329062,I329080);
not I_2521 (I45579,I45562);
nor I_2522 (I45596,I45579,I45545);
nor I_2523 (I45613,I45497,I45596);
DFFARX1 I_2524 (I45613,I2683,I45364,I45350,);
nor I_2525 (I45347,I45562,I45449);
DFFARX1 I_2526 (I45562,I2683,I45364,I45353,);
nor I_2527 (I45672,I45528,I329062);
nor I_2528 (I45689,I45672,I329068);
nor I_2529 (I45706,I329083,I329077);
DFFARX1 I_2530 (I45706,I2683,I45364,I45732,);
nor I_2531 (I45332,I45732,I45689);
DFFARX1 I_2532 (I45732,I2683,I45364,I45763,);
nand I_2533 (I45771,I45763,I329074);
nor I_2534 (I45356,I45398,I45771);
not I_2535 (I45802,I45732);
nand I_2536 (I45819,I45802,I329074);
nor I_2537 (I45836,I45398,I45819);
nor I_2538 (I45338,I45424,I45836);
nor I_2539 (I45867,I329083,I329071);
nor I_2540 (I45884,I45424,I45867);
DFFARX1 I_2541 (I45884,I2683,I45364,I45329,);
and I_2542 (I45344,I45497,I329083);
not I_2543 (I45959,I2690);
DFFARX1 I_2544 (I287874,I2683,I45959,I45985,);
not I_2545 (I45993,I45985);
DFFARX1 I_2546 (I287895,I2683,I45959,I46019,);
not I_2547 (I46027,I287877);
or I_2548 (I46044,I287868,I287877);
nor I_2549 (I46061,I46019,I287868);
nand I_2550 (I45936,I46027,I46061);
nor I_2551 (I46092,I287880,I287868);
nand I_2552 (I45930,I46092,I46027);
not I_2553 (I46123,I287871);
nand I_2554 (I46140,I46027,I46123);
nor I_2555 (I46157,I287889,I287892);
not I_2556 (I46174,I46157);
nor I_2557 (I46191,I46174,I46140);
nor I_2558 (I46208,I46092,I46191);
DFFARX1 I_2559 (I46208,I2683,I45959,I45945,);
nor I_2560 (I45942,I46157,I46044);
DFFARX1 I_2561 (I46157,I2683,I45959,I45948,);
nor I_2562 (I46267,I46123,I287889);
nor I_2563 (I46284,I46267,I287877);
nor I_2564 (I46301,I287883,I287886);
DFFARX1 I_2565 (I46301,I2683,I45959,I46327,);
nor I_2566 (I45927,I46327,I46284);
DFFARX1 I_2567 (I46327,I2683,I45959,I46358,);
nand I_2568 (I46366,I46358,I287868);
nor I_2569 (I45951,I45993,I46366);
not I_2570 (I46397,I46327);
nand I_2571 (I46414,I46397,I287868);
nor I_2572 (I46431,I45993,I46414);
nor I_2573 (I45933,I46019,I46431);
nor I_2574 (I46462,I287883,I287880);
nor I_2575 (I46479,I46019,I46462);
DFFARX1 I_2576 (I46479,I2683,I45959,I45924,);
and I_2577 (I45939,I46092,I287883);
not I_2578 (I46554,I2690);
DFFARX1 I_2579 (I207679,I2683,I46554,I46580,);
not I_2580 (I46588,I46580);
DFFARX1 I_2581 (I207700,I2683,I46554,I46614,);
not I_2582 (I46622,I207679);
or I_2583 (I46639,I207691,I207679);
nor I_2584 (I46656,I46614,I207691);
nand I_2585 (I46531,I46622,I46656);
nor I_2586 (I46687,I207688,I207691);
nand I_2587 (I46525,I46687,I46622);
not I_2588 (I46718,I207697);
nand I_2589 (I46735,I46622,I46718);
nor I_2590 (I46752,I207682,I207682);
not I_2591 (I46769,I46752);
nor I_2592 (I46786,I46769,I46735);
nor I_2593 (I46803,I46687,I46786);
DFFARX1 I_2594 (I46803,I2683,I46554,I46540,);
nor I_2595 (I46537,I46752,I46639);
DFFARX1 I_2596 (I46752,I2683,I46554,I46543,);
nor I_2597 (I46862,I46718,I207682);
nor I_2598 (I46879,I46862,I207679);
nor I_2599 (I46896,I207703,I207685);
DFFARX1 I_2600 (I46896,I2683,I46554,I46922,);
nor I_2601 (I46522,I46922,I46879);
DFFARX1 I_2602 (I46922,I2683,I46554,I46953,);
nand I_2603 (I46961,I46953,I207694);
nor I_2604 (I46546,I46588,I46961);
not I_2605 (I46992,I46922);
nand I_2606 (I47009,I46992,I207694);
nor I_2607 (I47026,I46588,I47009);
nor I_2608 (I46528,I46614,I47026);
nor I_2609 (I47057,I207703,I207688);
nor I_2610 (I47074,I46614,I47057);
DFFARX1 I_2611 (I47074,I2683,I46554,I46519,);
and I_2612 (I46534,I46687,I207703);
not I_2613 (I47149,I2690);
DFFARX1 I_2614 (I352760,I2683,I47149,I47175,);
not I_2615 (I47183,I47175);
DFFARX1 I_2616 (I352757,I2683,I47149,I47209,);
not I_2617 (I47217,I352766);
or I_2618 (I47234,I352757,I352766);
nor I_2619 (I47251,I47209,I352757);
nand I_2620 (I47126,I47217,I47251);
nor I_2621 (I47282,I352769,I352757);
nand I_2622 (I47120,I47282,I47217);
not I_2623 (I47313,I352763);
nand I_2624 (I47330,I47217,I47313);
nor I_2625 (I47347,I352760,I352778);
not I_2626 (I47364,I47347);
nor I_2627 (I47381,I47364,I47330);
nor I_2628 (I47398,I47282,I47381);
DFFARX1 I_2629 (I47398,I2683,I47149,I47135,);
nor I_2630 (I47132,I47347,I47234);
DFFARX1 I_2631 (I47347,I2683,I47149,I47138,);
nor I_2632 (I47457,I47313,I352760);
nor I_2633 (I47474,I47457,I352766);
nor I_2634 (I47491,I352781,I352775);
DFFARX1 I_2635 (I47491,I2683,I47149,I47517,);
nor I_2636 (I47117,I47517,I47474);
DFFARX1 I_2637 (I47517,I2683,I47149,I47548,);
nand I_2638 (I47556,I47548,I352772);
nor I_2639 (I47141,I47183,I47556);
not I_2640 (I47587,I47517);
nand I_2641 (I47604,I47587,I352772);
nor I_2642 (I47621,I47183,I47604);
nor I_2643 (I47123,I47209,I47621);
nor I_2644 (I47652,I352781,I352769);
nor I_2645 (I47669,I47209,I47652);
DFFARX1 I_2646 (I47669,I2683,I47149,I47114,);
and I_2647 (I47129,I47282,I352781);
not I_2648 (I47744,I2690);
DFFARX1 I_2649 (I271078,I2683,I47744,I47770,);
not I_2650 (I47778,I47770);
DFFARX1 I_2651 (I271099,I2683,I47744,I47804,);
not I_2652 (I47812,I271081);
or I_2653 (I47829,I271072,I271081);
nor I_2654 (I47846,I47804,I271072);
nand I_2655 (I47721,I47812,I47846);
nor I_2656 (I47877,I271084,I271072);
nand I_2657 (I47715,I47877,I47812);
not I_2658 (I47908,I271075);
nand I_2659 (I47925,I47812,I47908);
nor I_2660 (I47942,I271093,I271096);
not I_2661 (I47959,I47942);
nor I_2662 (I47976,I47959,I47925);
nor I_2663 (I47993,I47877,I47976);
DFFARX1 I_2664 (I47993,I2683,I47744,I47730,);
nor I_2665 (I47727,I47942,I47829);
DFFARX1 I_2666 (I47942,I2683,I47744,I47733,);
nor I_2667 (I48052,I47908,I271093);
nor I_2668 (I48069,I48052,I271081);
nor I_2669 (I48086,I271087,I271090);
DFFARX1 I_2670 (I48086,I2683,I47744,I48112,);
nor I_2671 (I47712,I48112,I48069);
DFFARX1 I_2672 (I48112,I2683,I47744,I48143,);
nand I_2673 (I48151,I48143,I271072);
nor I_2674 (I47736,I47778,I48151);
not I_2675 (I48182,I48112);
nand I_2676 (I48199,I48182,I271072);
nor I_2677 (I48216,I47778,I48199);
nor I_2678 (I47718,I47804,I48216);
nor I_2679 (I48247,I271087,I271084);
nor I_2680 (I48264,I47804,I48247);
DFFARX1 I_2681 (I48264,I2683,I47744,I47709,);
and I_2682 (I47724,I47877,I271087);
not I_2683 (I48336,I2690);
DFFARX1 I_2684 (I305325,I2683,I48336,I48362,);
DFFARX1 I_2685 (I48362,I2683,I48336,I48379,);
not I_2686 (I48328,I48379);
not I_2687 (I48401,I48362);
DFFARX1 I_2688 (I305334,I2683,I48336,I48427,);
not I_2689 (I48435,I48427);
and I_2690 (I48452,I48401,I305322);
not I_2691 (I48469,I305313);
nand I_2692 (I48486,I48469,I305322);
not I_2693 (I48503,I305319);
nor I_2694 (I48520,I48503,I305337);
nand I_2695 (I48537,I48520,I305310);
nor I_2696 (I48554,I48537,I48486);
DFFARX1 I_2697 (I48554,I2683,I48336,I48304,);
not I_2698 (I48585,I48537);
not I_2699 (I48602,I305337);
nand I_2700 (I48619,I48602,I305322);
nor I_2701 (I48636,I305337,I305313);
nand I_2702 (I48316,I48452,I48636);
nand I_2703 (I48310,I48401,I305337);
nand I_2704 (I48681,I48503,I305316);
DFFARX1 I_2705 (I48681,I2683,I48336,I48325,);
DFFARX1 I_2706 (I48681,I2683,I48336,I48319,);
not I_2707 (I48726,I305316);
nor I_2708 (I48743,I48726,I305328);
and I_2709 (I48760,I48743,I305310);
or I_2710 (I48777,I48760,I305331);
DFFARX1 I_2711 (I48777,I2683,I48336,I48803,);
nand I_2712 (I48811,I48803,I48469);
nor I_2713 (I48313,I48811,I48619);
nor I_2714 (I48307,I48803,I48435);
DFFARX1 I_2715 (I48803,I2683,I48336,I48865,);
not I_2716 (I48873,I48865);
nor I_2717 (I48322,I48873,I48585);
not I_2718 (I48931,I2690);
DFFARX1 I_2719 (I259773,I2683,I48931,I48957,);
DFFARX1 I_2720 (I48957,I2683,I48931,I48974,);
not I_2721 (I48923,I48974);
not I_2722 (I48996,I48957);
DFFARX1 I_2723 (I259767,I2683,I48931,I49022,);
not I_2724 (I49030,I49022);
and I_2725 (I49047,I48996,I259785);
not I_2726 (I49064,I259773);
nand I_2727 (I49081,I49064,I259785);
not I_2728 (I49098,I259767);
nor I_2729 (I49115,I49098,I259779);
nand I_2730 (I49132,I49115,I259770);
nor I_2731 (I49149,I49132,I49081);
DFFARX1 I_2732 (I49149,I2683,I48931,I48899,);
not I_2733 (I49180,I49132);
not I_2734 (I49197,I259779);
nand I_2735 (I49214,I49197,I259785);
nor I_2736 (I49231,I259779,I259773);
nand I_2737 (I48911,I49047,I49231);
nand I_2738 (I48905,I48996,I259779);
nand I_2739 (I49276,I49098,I259782);
DFFARX1 I_2740 (I49276,I2683,I48931,I48920,);
DFFARX1 I_2741 (I49276,I2683,I48931,I48914,);
not I_2742 (I49321,I259782);
nor I_2743 (I49338,I49321,I259788);
and I_2744 (I49355,I49338,I259770);
or I_2745 (I49372,I49355,I259776);
DFFARX1 I_2746 (I49372,I2683,I48931,I49398,);
nand I_2747 (I49406,I49398,I49064);
nor I_2748 (I48908,I49406,I49214);
nor I_2749 (I48902,I49398,I49030);
DFFARX1 I_2750 (I49398,I2683,I48931,I49460,);
not I_2751 (I49468,I49460);
nor I_2752 (I48917,I49468,I49180);
not I_2753 (I49526,I2690);
DFFARX1 I_2754 (I223875,I2683,I49526,I49552,);
DFFARX1 I_2755 (I49552,I2683,I49526,I49569,);
not I_2756 (I49518,I49569);
not I_2757 (I49591,I49552);
DFFARX1 I_2758 (I223872,I2683,I49526,I49617,);
not I_2759 (I49625,I49617);
and I_2760 (I49642,I49591,I223878);
not I_2761 (I49659,I223863);
nand I_2762 (I49676,I49659,I223878);
not I_2763 (I49693,I223866);
nor I_2764 (I49710,I49693,I223887);
nand I_2765 (I49727,I49710,I223884);
nor I_2766 (I49744,I49727,I49676);
DFFARX1 I_2767 (I49744,I2683,I49526,I49494,);
not I_2768 (I49775,I49727);
not I_2769 (I49792,I223887);
nand I_2770 (I49809,I49792,I223878);
nor I_2771 (I49826,I223887,I223863);
nand I_2772 (I49506,I49642,I49826);
nand I_2773 (I49500,I49591,I223887);
nand I_2774 (I49871,I49693,I223863);
DFFARX1 I_2775 (I49871,I2683,I49526,I49515,);
DFFARX1 I_2776 (I49871,I2683,I49526,I49509,);
not I_2777 (I49916,I223863);
nor I_2778 (I49933,I49916,I223869);
and I_2779 (I49950,I49933,I223881);
or I_2780 (I49967,I49950,I223866);
DFFARX1 I_2781 (I49967,I2683,I49526,I49993,);
nand I_2782 (I50001,I49993,I49659);
nor I_2783 (I49503,I50001,I49809);
nor I_2784 (I49497,I49993,I49625);
DFFARX1 I_2785 (I49993,I2683,I49526,I50055,);
not I_2786 (I50063,I50055);
nor I_2787 (I49512,I50063,I49775);
not I_2788 (I50121,I2690);
DFFARX1 I_2789 (I157031,I2683,I50121,I50147,);
DFFARX1 I_2790 (I50147,I2683,I50121,I50164,);
not I_2791 (I50113,I50164);
not I_2792 (I50186,I50147);
DFFARX1 I_2793 (I157025,I2683,I50121,I50212,);
not I_2794 (I50220,I50212);
and I_2795 (I50237,I50186,I157040);
not I_2796 (I50254,I157037);
nand I_2797 (I50271,I50254,I157040);
not I_2798 (I50288,I157028);
nor I_2799 (I50305,I50288,I157019);
nand I_2800 (I50322,I50305,I157022);
nor I_2801 (I50339,I50322,I50271);
DFFARX1 I_2802 (I50339,I2683,I50121,I50089,);
not I_2803 (I50370,I50322);
not I_2804 (I50387,I157019);
nand I_2805 (I50404,I50387,I157040);
nor I_2806 (I50421,I157019,I157037);
nand I_2807 (I50101,I50237,I50421);
nand I_2808 (I50095,I50186,I157019);
nand I_2809 (I50466,I50288,I157043);
DFFARX1 I_2810 (I50466,I2683,I50121,I50110,);
DFFARX1 I_2811 (I50466,I2683,I50121,I50104,);
not I_2812 (I50511,I157043);
nor I_2813 (I50528,I50511,I157034);
and I_2814 (I50545,I50528,I157019);
or I_2815 (I50562,I50545,I157022);
DFFARX1 I_2816 (I50562,I2683,I50121,I50588,);
nand I_2817 (I50596,I50588,I50254);
nor I_2818 (I50098,I50596,I50404);
nor I_2819 (I50092,I50588,I50220);
DFFARX1 I_2820 (I50588,I2683,I50121,I50650,);
not I_2821 (I50658,I50650);
nor I_2822 (I50107,I50658,I50370);
not I_2823 (I50716,I2690);
DFFARX1 I_2824 (I193819,I2683,I50716,I50742,);
DFFARX1 I_2825 (I50742,I2683,I50716,I50759,);
not I_2826 (I50708,I50759);
not I_2827 (I50781,I50742);
DFFARX1 I_2828 (I193816,I2683,I50716,I50807,);
not I_2829 (I50815,I50807);
and I_2830 (I50832,I50781,I193822);
not I_2831 (I50849,I193807);
nand I_2832 (I50866,I50849,I193822);
not I_2833 (I50883,I193810);
nor I_2834 (I50900,I50883,I193831);
nand I_2835 (I50917,I50900,I193828);
nor I_2836 (I50934,I50917,I50866);
DFFARX1 I_2837 (I50934,I2683,I50716,I50684,);
not I_2838 (I50965,I50917);
not I_2839 (I50982,I193831);
nand I_2840 (I50999,I50982,I193822);
nor I_2841 (I51016,I193831,I193807);
nand I_2842 (I50696,I50832,I51016);
nand I_2843 (I50690,I50781,I193831);
nand I_2844 (I51061,I50883,I193807);
DFFARX1 I_2845 (I51061,I2683,I50716,I50705,);
DFFARX1 I_2846 (I51061,I2683,I50716,I50699,);
not I_2847 (I51106,I193807);
nor I_2848 (I51123,I51106,I193813);
and I_2849 (I51140,I51123,I193825);
or I_2850 (I51157,I51140,I193810);
DFFARX1 I_2851 (I51157,I2683,I50716,I51183,);
nand I_2852 (I51191,I51183,I50849);
nor I_2853 (I50693,I51191,I50999);
nor I_2854 (I50687,I51183,I50815);
DFFARX1 I_2855 (I51183,I2683,I50716,I51245,);
not I_2856 (I51253,I51245);
nor I_2857 (I50702,I51253,I50965);
not I_2858 (I51311,I2690);
DFFARX1 I_2859 (I130727,I2683,I51311,I51337,);
DFFARX1 I_2860 (I51337,I2683,I51311,I51354,);
not I_2861 (I51303,I51354);
not I_2862 (I51376,I51337);
DFFARX1 I_2863 (I130715,I2683,I51311,I51402,);
not I_2864 (I51410,I51402);
and I_2865 (I51427,I51376,I130724);
not I_2866 (I51444,I130721);
nand I_2867 (I51461,I51444,I130724);
not I_2868 (I51478,I130712);
nor I_2869 (I51495,I51478,I130718);
nand I_2870 (I51512,I51495,I130703);
nor I_2871 (I51529,I51512,I51461);
DFFARX1 I_2872 (I51529,I2683,I51311,I51279,);
not I_2873 (I51560,I51512);
not I_2874 (I51577,I130718);
nand I_2875 (I51594,I51577,I130724);
nor I_2876 (I51611,I130718,I130721);
nand I_2877 (I51291,I51427,I51611);
nand I_2878 (I51285,I51376,I130718);
nand I_2879 (I51656,I51478,I130703);
DFFARX1 I_2880 (I51656,I2683,I51311,I51300,);
DFFARX1 I_2881 (I51656,I2683,I51311,I51294,);
not I_2882 (I51701,I130703);
nor I_2883 (I51718,I51701,I130709);
and I_2884 (I51735,I51718,I130706);
or I_2885 (I51752,I51735,I130730);
DFFARX1 I_2886 (I51752,I2683,I51311,I51778,);
nand I_2887 (I51786,I51778,I51444);
nor I_2888 (I51288,I51786,I51594);
nor I_2889 (I51282,I51778,I51410);
DFFARX1 I_2890 (I51778,I2683,I51311,I51840,);
not I_2891 (I51848,I51840);
nor I_2892 (I51297,I51848,I51560);
not I_2893 (I51906,I2690);
DFFARX1 I_2894 (I359115,I2683,I51906,I51932,);
DFFARX1 I_2895 (I51932,I2683,I51906,I51949,);
not I_2896 (I51898,I51949);
not I_2897 (I51971,I51932);
DFFARX1 I_2898 (I359115,I2683,I51906,I51997,);
not I_2899 (I52005,I51997);
and I_2900 (I52022,I51971,I359118);
not I_2901 (I52039,I359130);
nand I_2902 (I52056,I52039,I359118);
not I_2903 (I52073,I359136);
nor I_2904 (I52090,I52073,I359127);
nand I_2905 (I52107,I52090,I359133);
nor I_2906 (I52124,I52107,I52056);
DFFARX1 I_2907 (I52124,I2683,I51906,I51874,);
not I_2908 (I52155,I52107);
not I_2909 (I52172,I359127);
nand I_2910 (I52189,I52172,I359118);
nor I_2911 (I52206,I359127,I359130);
nand I_2912 (I51886,I52022,I52206);
nand I_2913 (I51880,I51971,I359127);
nand I_2914 (I52251,I52073,I359124);
DFFARX1 I_2915 (I52251,I2683,I51906,I51895,);
DFFARX1 I_2916 (I52251,I2683,I51906,I51889,);
not I_2917 (I52296,I359124);
nor I_2918 (I52313,I52296,I359121);
and I_2919 (I52330,I52313,I359139);
or I_2920 (I52347,I52330,I359118);
DFFARX1 I_2921 (I52347,I2683,I51906,I52373,);
nand I_2922 (I52381,I52373,I52039);
nor I_2923 (I51883,I52381,I52189);
nor I_2924 (I51877,I52373,I52005);
DFFARX1 I_2925 (I52373,I2683,I51906,I52435,);
not I_2926 (I52443,I52435);
nor I_2927 (I51892,I52443,I52155);
not I_2928 (I52501,I2690);
DFFARX1 I_2929 (I238693,I2683,I52501,I52527,);
DFFARX1 I_2930 (I52527,I2683,I52501,I52544,);
not I_2931 (I52493,I52544);
not I_2932 (I52566,I52527);
DFFARX1 I_2933 (I238687,I2683,I52501,I52592,);
not I_2934 (I52600,I52592);
and I_2935 (I52617,I52566,I238705);
not I_2936 (I52634,I238693);
nand I_2937 (I52651,I52634,I238705);
not I_2938 (I52668,I238687);
nor I_2939 (I52685,I52668,I238699);
nand I_2940 (I52702,I52685,I238690);
nor I_2941 (I52719,I52702,I52651);
DFFARX1 I_2942 (I52719,I2683,I52501,I52469,);
not I_2943 (I52750,I52702);
not I_2944 (I52767,I238699);
nand I_2945 (I52784,I52767,I238705);
nor I_2946 (I52801,I238699,I238693);
nand I_2947 (I52481,I52617,I52801);
nand I_2948 (I52475,I52566,I238699);
nand I_2949 (I52846,I52668,I238702);
DFFARX1 I_2950 (I52846,I2683,I52501,I52490,);
DFFARX1 I_2951 (I52846,I2683,I52501,I52484,);
not I_2952 (I52891,I238702);
nor I_2953 (I52908,I52891,I238708);
and I_2954 (I52925,I52908,I238690);
or I_2955 (I52942,I52925,I238696);
DFFARX1 I_2956 (I52942,I2683,I52501,I52968,);
nand I_2957 (I52976,I52968,I52634);
nor I_2958 (I52478,I52976,I52784);
nor I_2959 (I52472,I52968,I52600);
DFFARX1 I_2960 (I52968,I2683,I52501,I53030,);
not I_2961 (I53038,I53030);
nor I_2962 (I52487,I53038,I52750);
not I_2963 (I53096,I2690);
DFFARX1 I_2964 (I94748,I2683,I53096,I53122,);
DFFARX1 I_2965 (I53122,I2683,I53096,I53139,);
not I_2966 (I53088,I53139);
not I_2967 (I53161,I53122);
DFFARX1 I_2968 (I94763,I2683,I53096,I53187,);
not I_2969 (I53195,I53187);
and I_2970 (I53212,I53161,I94760);
not I_2971 (I53229,I94748);
nand I_2972 (I53246,I53229,I94760);
not I_2973 (I53263,I94757);
nor I_2974 (I53280,I53263,I94772);
nand I_2975 (I53297,I53280,I94769);
nor I_2976 (I53314,I53297,I53246);
DFFARX1 I_2977 (I53314,I2683,I53096,I53064,);
not I_2978 (I53345,I53297);
not I_2979 (I53362,I94772);
nand I_2980 (I53379,I53362,I94760);
nor I_2981 (I53396,I94772,I94748);
nand I_2982 (I53076,I53212,I53396);
nand I_2983 (I53070,I53161,I94772);
nand I_2984 (I53441,I53263,I94766);
DFFARX1 I_2985 (I53441,I2683,I53096,I53085,);
DFFARX1 I_2986 (I53441,I2683,I53096,I53079,);
not I_2987 (I53486,I94766);
nor I_2988 (I53503,I53486,I94754);
and I_2989 (I53520,I53503,I94775);
or I_2990 (I53537,I53520,I94751);
DFFARX1 I_2991 (I53537,I2683,I53096,I53563,);
nand I_2992 (I53571,I53563,I53229);
nor I_2993 (I53073,I53571,I53379);
nor I_2994 (I53067,I53563,I53195);
DFFARX1 I_2995 (I53563,I2683,I53096,I53625,);
not I_2996 (I53633,I53625);
nor I_2997 (I53082,I53633,I53345);
not I_2998 (I53691,I2690);
DFFARX1 I_2999 (I252922,I2683,I53691,I53717,);
DFFARX1 I_3000 (I53717,I2683,I53691,I53734,);
not I_3001 (I53683,I53734);
not I_3002 (I53756,I53717);
DFFARX1 I_3003 (I252916,I2683,I53691,I53782,);
not I_3004 (I53790,I53782);
and I_3005 (I53807,I53756,I252934);
not I_3006 (I53824,I252922);
nand I_3007 (I53841,I53824,I252934);
not I_3008 (I53858,I252916);
nor I_3009 (I53875,I53858,I252928);
nand I_3010 (I53892,I53875,I252919);
nor I_3011 (I53909,I53892,I53841);
DFFARX1 I_3012 (I53909,I2683,I53691,I53659,);
not I_3013 (I53940,I53892);
not I_3014 (I53957,I252928);
nand I_3015 (I53974,I53957,I252934);
nor I_3016 (I53991,I252928,I252922);
nand I_3017 (I53671,I53807,I53991);
nand I_3018 (I53665,I53756,I252928);
nand I_3019 (I54036,I53858,I252931);
DFFARX1 I_3020 (I54036,I2683,I53691,I53680,);
DFFARX1 I_3021 (I54036,I2683,I53691,I53674,);
not I_3022 (I54081,I252931);
nor I_3023 (I54098,I54081,I252937);
and I_3024 (I54115,I54098,I252919);
or I_3025 (I54132,I54115,I252925);
DFFARX1 I_3026 (I54132,I2683,I53691,I54158,);
nand I_3027 (I54166,I54158,I53824);
nor I_3028 (I53668,I54166,I53974);
nor I_3029 (I53662,I54158,I53790);
DFFARX1 I_3030 (I54158,I2683,I53691,I54220,);
not I_3031 (I54228,I54220);
nor I_3032 (I53677,I54228,I53940);
not I_3033 (I54286,I2690);
DFFARX1 I_3034 (I126919,I2683,I54286,I54312,);
DFFARX1 I_3035 (I54312,I2683,I54286,I54329,);
not I_3036 (I54278,I54329);
not I_3037 (I54351,I54312);
DFFARX1 I_3038 (I126907,I2683,I54286,I54377,);
not I_3039 (I54385,I54377);
and I_3040 (I54402,I54351,I126916);
not I_3041 (I54419,I126913);
nand I_3042 (I54436,I54419,I126916);
not I_3043 (I54453,I126904);
nor I_3044 (I54470,I54453,I126910);
nand I_3045 (I54487,I54470,I126895);
nor I_3046 (I54504,I54487,I54436);
DFFARX1 I_3047 (I54504,I2683,I54286,I54254,);
not I_3048 (I54535,I54487);
not I_3049 (I54552,I126910);
nand I_3050 (I54569,I54552,I126916);
nor I_3051 (I54586,I126910,I126913);
nand I_3052 (I54266,I54402,I54586);
nand I_3053 (I54260,I54351,I126910);
nand I_3054 (I54631,I54453,I126895);
DFFARX1 I_3055 (I54631,I2683,I54286,I54275,);
DFFARX1 I_3056 (I54631,I2683,I54286,I54269,);
not I_3057 (I54676,I126895);
nor I_3058 (I54693,I54676,I126901);
and I_3059 (I54710,I54693,I126898);
or I_3060 (I54727,I54710,I126922);
DFFARX1 I_3061 (I54727,I2683,I54286,I54753,);
nand I_3062 (I54761,I54753,I54419);
nor I_3063 (I54263,I54761,I54569);
nor I_3064 (I54257,I54753,I54385);
DFFARX1 I_3065 (I54753,I2683,I54286,I54815,);
not I_3066 (I54823,I54815);
nor I_3067 (I54272,I54823,I54535);
not I_3068 (I54881,I2690);
DFFARX1 I_3069 (I102126,I2683,I54881,I54907,);
DFFARX1 I_3070 (I54907,I2683,I54881,I54924,);
not I_3071 (I54873,I54924);
not I_3072 (I54946,I54907);
DFFARX1 I_3073 (I102141,I2683,I54881,I54972,);
not I_3074 (I54980,I54972);
and I_3075 (I54997,I54946,I102138);
not I_3076 (I55014,I102126);
nand I_3077 (I55031,I55014,I102138);
not I_3078 (I55048,I102135);
nor I_3079 (I55065,I55048,I102150);
nand I_3080 (I55082,I55065,I102147);
nor I_3081 (I55099,I55082,I55031);
DFFARX1 I_3082 (I55099,I2683,I54881,I54849,);
not I_3083 (I55130,I55082);
not I_3084 (I55147,I102150);
nand I_3085 (I55164,I55147,I102138);
nor I_3086 (I55181,I102150,I102126);
nand I_3087 (I54861,I54997,I55181);
nand I_3088 (I54855,I54946,I102150);
nand I_3089 (I55226,I55048,I102144);
DFFARX1 I_3090 (I55226,I2683,I54881,I54870,);
DFFARX1 I_3091 (I55226,I2683,I54881,I54864,);
not I_3092 (I55271,I102144);
nor I_3093 (I55288,I55271,I102132);
and I_3094 (I55305,I55288,I102153);
or I_3095 (I55322,I55305,I102129);
DFFARX1 I_3096 (I55322,I2683,I54881,I55348,);
nand I_3097 (I55356,I55348,I55014);
nor I_3098 (I54858,I55356,I55164);
nor I_3099 (I54852,I55348,I54980);
DFFARX1 I_3100 (I55348,I2683,I54881,I55410,);
not I_3101 (I55418,I55410);
nor I_3102 (I54867,I55418,I55130);
not I_3103 (I55476,I2690);
DFFARX1 I_3104 (I154651,I2683,I55476,I55502,);
DFFARX1 I_3105 (I55502,I2683,I55476,I55519,);
not I_3106 (I55468,I55519);
not I_3107 (I55541,I55502);
DFFARX1 I_3108 (I154645,I2683,I55476,I55567,);
not I_3109 (I55575,I55567);
and I_3110 (I55592,I55541,I154660);
not I_3111 (I55609,I154657);
nand I_3112 (I55626,I55609,I154660);
not I_3113 (I55643,I154648);
nor I_3114 (I55660,I55643,I154639);
nand I_3115 (I55677,I55660,I154642);
nor I_3116 (I55694,I55677,I55626);
DFFARX1 I_3117 (I55694,I2683,I55476,I55444,);
not I_3118 (I55725,I55677);
not I_3119 (I55742,I154639);
nand I_3120 (I55759,I55742,I154660);
nor I_3121 (I55776,I154639,I154657);
nand I_3122 (I55456,I55592,I55776);
nand I_3123 (I55450,I55541,I154639);
nand I_3124 (I55821,I55643,I154663);
DFFARX1 I_3125 (I55821,I2683,I55476,I55465,);
DFFARX1 I_3126 (I55821,I2683,I55476,I55459,);
not I_3127 (I55866,I154663);
nor I_3128 (I55883,I55866,I154654);
and I_3129 (I55900,I55883,I154639);
or I_3130 (I55917,I55900,I154642);
DFFARX1 I_3131 (I55917,I2683,I55476,I55943,);
nand I_3132 (I55951,I55943,I55609);
nor I_3133 (I55453,I55951,I55759);
nor I_3134 (I55447,I55943,I55575);
DFFARX1 I_3135 (I55943,I2683,I55476,I56005,);
not I_3136 (I56013,I56005);
nor I_3137 (I55462,I56013,I55725);
not I_3138 (I56071,I2690);
DFFARX1 I_3139 (I364879,I2683,I56071,I56097,);
DFFARX1 I_3140 (I56097,I2683,I56071,I56114,);
not I_3141 (I56063,I56114);
not I_3142 (I56136,I56097);
DFFARX1 I_3143 (I364864,I2683,I56071,I56162,);
not I_3144 (I56170,I56162);
and I_3145 (I56187,I56136,I364882);
not I_3146 (I56204,I364864);
nand I_3147 (I56221,I56204,I364882);
not I_3148 (I56238,I364885);
nor I_3149 (I56255,I56238,I364876);
nand I_3150 (I56272,I56255,I364873);
nor I_3151 (I56289,I56272,I56221);
DFFARX1 I_3152 (I56289,I2683,I56071,I56039,);
not I_3153 (I56320,I56272);
not I_3154 (I56337,I364876);
nand I_3155 (I56354,I56337,I364882);
nor I_3156 (I56371,I364876,I364864);
nand I_3157 (I56051,I56187,I56371);
nand I_3158 (I56045,I56136,I364876);
nand I_3159 (I56416,I56238,I364870);
DFFARX1 I_3160 (I56416,I2683,I56071,I56060,);
DFFARX1 I_3161 (I56416,I2683,I56071,I56054,);
not I_3162 (I56461,I364870);
nor I_3163 (I56478,I56461,I364861);
and I_3164 (I56495,I56478,I364867);
or I_3165 (I56512,I56495,I364861);
DFFARX1 I_3166 (I56512,I2683,I56071,I56538,);
nand I_3167 (I56546,I56538,I56204);
nor I_3168 (I56048,I56546,I56354);
nor I_3169 (I56042,I56538,I56170);
DFFARX1 I_3170 (I56538,I2683,I56071,I56600,);
not I_3171 (I56608,I56600);
nor I_3172 (I56057,I56608,I56320);
not I_3173 (I56666,I2690);
DFFARX1 I_3174 (I329637,I2683,I56666,I56692,);
DFFARX1 I_3175 (I56692,I2683,I56666,I56709,);
not I_3176 (I56658,I56709);
not I_3177 (I56731,I56692);
DFFARX1 I_3178 (I329637,I2683,I56666,I56757,);
not I_3179 (I56765,I56757);
and I_3180 (I56782,I56731,I329640);
not I_3181 (I56799,I329652);
nand I_3182 (I56816,I56799,I329640);
not I_3183 (I56833,I329658);
nor I_3184 (I56850,I56833,I329649);
nand I_3185 (I56867,I56850,I329655);
nor I_3186 (I56884,I56867,I56816);
DFFARX1 I_3187 (I56884,I2683,I56666,I56634,);
not I_3188 (I56915,I56867);
not I_3189 (I56932,I329649);
nand I_3190 (I56949,I56932,I329640);
nor I_3191 (I56966,I329649,I329652);
nand I_3192 (I56646,I56782,I56966);
nand I_3193 (I56640,I56731,I329649);
nand I_3194 (I57011,I56833,I329646);
DFFARX1 I_3195 (I57011,I2683,I56666,I56655,);
DFFARX1 I_3196 (I57011,I2683,I56666,I56649,);
not I_3197 (I57056,I329646);
nor I_3198 (I57073,I57056,I329643);
and I_3199 (I57090,I57073,I329661);
or I_3200 (I57107,I57090,I329640);
DFFARX1 I_3201 (I57107,I2683,I56666,I57133,);
nand I_3202 (I57141,I57133,I56799);
nor I_3203 (I56643,I57141,I56949);
nor I_3204 (I56637,I57133,I56765);
DFFARX1 I_3205 (I57133,I2683,I56666,I57195,);
not I_3206 (I57203,I57195);
nor I_3207 (I56652,I57203,I56915);
not I_3208 (I57261,I2690);
DFFARX1 I_3209 (I144871,I2683,I57261,I57287,);
DFFARX1 I_3210 (I57287,I2683,I57261,I57304,);
not I_3211 (I57253,I57304);
not I_3212 (I57326,I57287);
DFFARX1 I_3213 (I144859,I2683,I57261,I57352,);
not I_3214 (I57360,I57352);
and I_3215 (I57377,I57326,I144868);
not I_3216 (I57394,I144865);
nand I_3217 (I57411,I57394,I144868);
not I_3218 (I57428,I144856);
nor I_3219 (I57445,I57428,I144862);
nand I_3220 (I57462,I57445,I144847);
nor I_3221 (I57479,I57462,I57411);
DFFARX1 I_3222 (I57479,I2683,I57261,I57229,);
not I_3223 (I57510,I57462);
not I_3224 (I57527,I144862);
nand I_3225 (I57544,I57527,I144868);
nor I_3226 (I57561,I144862,I144865);
nand I_3227 (I57241,I57377,I57561);
nand I_3228 (I57235,I57326,I144862);
nand I_3229 (I57606,I57428,I144847);
DFFARX1 I_3230 (I57606,I2683,I57261,I57250,);
DFFARX1 I_3231 (I57606,I2683,I57261,I57244,);
not I_3232 (I57651,I144847);
nor I_3233 (I57668,I57651,I144853);
and I_3234 (I57685,I57668,I144850);
or I_3235 (I57702,I57685,I144874);
DFFARX1 I_3236 (I57702,I2683,I57261,I57728,);
nand I_3237 (I57736,I57728,I57394);
nor I_3238 (I57238,I57736,I57544);
nor I_3239 (I57232,I57728,I57360);
DFFARX1 I_3240 (I57728,I2683,I57261,I57790,);
not I_3241 (I57798,I57790);
nor I_3242 (I57247,I57798,I57510);
not I_3243 (I57856,I2690);
DFFARX1 I_3244 (I97383,I2683,I57856,I57882,);
DFFARX1 I_3245 (I57882,I2683,I57856,I57899,);
not I_3246 (I57848,I57899);
not I_3247 (I57921,I57882);
DFFARX1 I_3248 (I97398,I2683,I57856,I57947,);
not I_3249 (I57955,I57947);
and I_3250 (I57972,I57921,I97395);
not I_3251 (I57989,I97383);
nand I_3252 (I58006,I57989,I97395);
not I_3253 (I58023,I97392);
nor I_3254 (I58040,I58023,I97407);
nand I_3255 (I58057,I58040,I97404);
nor I_3256 (I58074,I58057,I58006);
DFFARX1 I_3257 (I58074,I2683,I57856,I57824,);
not I_3258 (I58105,I58057);
not I_3259 (I58122,I97407);
nand I_3260 (I58139,I58122,I97395);
nor I_3261 (I58156,I97407,I97383);
nand I_3262 (I57836,I57972,I58156);
nand I_3263 (I57830,I57921,I97407);
nand I_3264 (I58201,I58023,I97401);
DFFARX1 I_3265 (I58201,I2683,I57856,I57845,);
DFFARX1 I_3266 (I58201,I2683,I57856,I57839,);
not I_3267 (I58246,I97401);
nor I_3268 (I58263,I58246,I97389);
and I_3269 (I58280,I58263,I97410);
or I_3270 (I58297,I58280,I97386);
DFFARX1 I_3271 (I58297,I2683,I57856,I58323,);
nand I_3272 (I58331,I58323,I57989);
nor I_3273 (I57833,I58331,I58139);
nor I_3274 (I57827,I58323,I57955);
DFFARX1 I_3275 (I58323,I2683,I57856,I58385,);
not I_3276 (I58393,I58385);
nor I_3277 (I57842,I58393,I58105);
not I_3278 (I58451,I2690);
DFFARX1 I_3279 (I324435,I2683,I58451,I58477,);
DFFARX1 I_3280 (I58477,I2683,I58451,I58494,);
not I_3281 (I58443,I58494);
not I_3282 (I58516,I58477);
DFFARX1 I_3283 (I324435,I2683,I58451,I58542,);
not I_3284 (I58550,I58542);
and I_3285 (I58567,I58516,I324438);
not I_3286 (I58584,I324450);
nand I_3287 (I58601,I58584,I324438);
not I_3288 (I58618,I324456);
nor I_3289 (I58635,I58618,I324447);
nand I_3290 (I58652,I58635,I324453);
nor I_3291 (I58669,I58652,I58601);
DFFARX1 I_3292 (I58669,I2683,I58451,I58419,);
not I_3293 (I58700,I58652);
not I_3294 (I58717,I324447);
nand I_3295 (I58734,I58717,I324438);
nor I_3296 (I58751,I324447,I324450);
nand I_3297 (I58431,I58567,I58751);
nand I_3298 (I58425,I58516,I324447);
nand I_3299 (I58796,I58618,I324444);
DFFARX1 I_3300 (I58796,I2683,I58451,I58440,);
DFFARX1 I_3301 (I58796,I2683,I58451,I58434,);
not I_3302 (I58841,I324444);
nor I_3303 (I58858,I58841,I324441);
and I_3304 (I58875,I58858,I324459);
or I_3305 (I58892,I58875,I324438);
DFFARX1 I_3306 (I58892,I2683,I58451,I58918,);
nand I_3307 (I58926,I58918,I58584);
nor I_3308 (I58428,I58926,I58734);
nor I_3309 (I58422,I58918,I58550);
DFFARX1 I_3310 (I58918,I2683,I58451,I58980,);
not I_3311 (I58988,I58980);
nor I_3312 (I58437,I58988,I58700);
not I_3313 (I59046,I2690);
DFFARX1 I_3314 (I156436,I2683,I59046,I59072,);
DFFARX1 I_3315 (I59072,I2683,I59046,I59089,);
not I_3316 (I59038,I59089);
not I_3317 (I59111,I59072);
DFFARX1 I_3318 (I156430,I2683,I59046,I59137,);
not I_3319 (I59145,I59137);
and I_3320 (I59162,I59111,I156445);
not I_3321 (I59179,I156442);
nand I_3322 (I59196,I59179,I156445);
not I_3323 (I59213,I156433);
nor I_3324 (I59230,I59213,I156424);
nand I_3325 (I59247,I59230,I156427);
nor I_3326 (I59264,I59247,I59196);
DFFARX1 I_3327 (I59264,I2683,I59046,I59014,);
not I_3328 (I59295,I59247);
not I_3329 (I59312,I156424);
nand I_3330 (I59329,I59312,I156445);
nor I_3331 (I59346,I156424,I156442);
nand I_3332 (I59026,I59162,I59346);
nand I_3333 (I59020,I59111,I156424);
nand I_3334 (I59391,I59213,I156448);
DFFARX1 I_3335 (I59391,I2683,I59046,I59035,);
DFFARX1 I_3336 (I59391,I2683,I59046,I59029,);
not I_3337 (I59436,I156448);
nor I_3338 (I59453,I59436,I156439);
and I_3339 (I59470,I59453,I156424);
or I_3340 (I59487,I59470,I156427);
DFFARX1 I_3341 (I59487,I2683,I59046,I59513,);
nand I_3342 (I59521,I59513,I59179);
nor I_3343 (I59023,I59521,I59329);
nor I_3344 (I59017,I59513,I59145);
DFFARX1 I_3345 (I59513,I2683,I59046,I59575,);
not I_3346 (I59583,I59575);
nor I_3347 (I59032,I59583,I59295);
not I_3348 (I59641,I2690);
DFFARX1 I_3349 (I296927,I2683,I59641,I59667,);
DFFARX1 I_3350 (I59667,I2683,I59641,I59684,);
not I_3351 (I59633,I59684);
not I_3352 (I59706,I59667);
DFFARX1 I_3353 (I296936,I2683,I59641,I59732,);
not I_3354 (I59740,I59732);
and I_3355 (I59757,I59706,I296924);
not I_3356 (I59774,I296915);
nand I_3357 (I59791,I59774,I296924);
not I_3358 (I59808,I296921);
nor I_3359 (I59825,I59808,I296939);
nand I_3360 (I59842,I59825,I296912);
nor I_3361 (I59859,I59842,I59791);
DFFARX1 I_3362 (I59859,I2683,I59641,I59609,);
not I_3363 (I59890,I59842);
not I_3364 (I59907,I296939);
nand I_3365 (I59924,I59907,I296924);
nor I_3366 (I59941,I296939,I296915);
nand I_3367 (I59621,I59757,I59941);
nand I_3368 (I59615,I59706,I296939);
nand I_3369 (I59986,I59808,I296918);
DFFARX1 I_3370 (I59986,I2683,I59641,I59630,);
DFFARX1 I_3371 (I59986,I2683,I59641,I59624,);
not I_3372 (I60031,I296918);
nor I_3373 (I60048,I60031,I296930);
and I_3374 (I60065,I60048,I296912);
or I_3375 (I60082,I60065,I296933);
DFFARX1 I_3376 (I60082,I2683,I59641,I60108,);
nand I_3377 (I60116,I60108,I59774);
nor I_3378 (I59618,I60116,I59924);
nor I_3379 (I59612,I60108,I59740);
DFFARX1 I_3380 (I60108,I2683,I59641,I60170,);
not I_3381 (I60178,I60170);
nor I_3382 (I59627,I60178,I59890);
not I_3383 (I60236,I2690);
DFFARX1 I_3384 (I115828,I2683,I60236,I60262,);
DFFARX1 I_3385 (I60262,I2683,I60236,I60279,);
not I_3386 (I60228,I60279);
not I_3387 (I60301,I60262);
DFFARX1 I_3388 (I115843,I2683,I60236,I60327,);
not I_3389 (I60335,I60327);
and I_3390 (I60352,I60301,I115840);
not I_3391 (I60369,I115828);
nand I_3392 (I60386,I60369,I115840);
not I_3393 (I60403,I115837);
nor I_3394 (I60420,I60403,I115852);
nand I_3395 (I60437,I60420,I115849);
nor I_3396 (I60454,I60437,I60386);
DFFARX1 I_3397 (I60454,I2683,I60236,I60204,);
not I_3398 (I60485,I60437);
not I_3399 (I60502,I115852);
nand I_3400 (I60519,I60502,I115840);
nor I_3401 (I60536,I115852,I115828);
nand I_3402 (I60216,I60352,I60536);
nand I_3403 (I60210,I60301,I115852);
nand I_3404 (I60581,I60403,I115846);
DFFARX1 I_3405 (I60581,I2683,I60236,I60225,);
DFFARX1 I_3406 (I60581,I2683,I60236,I60219,);
not I_3407 (I60626,I115846);
nor I_3408 (I60643,I60626,I115834);
and I_3409 (I60660,I60643,I115855);
or I_3410 (I60677,I60660,I115831);
DFFARX1 I_3411 (I60677,I2683,I60236,I60703,);
nand I_3412 (I60711,I60703,I60369);
nor I_3413 (I60213,I60711,I60519);
nor I_3414 (I60207,I60703,I60335);
DFFARX1 I_3415 (I60703,I2683,I60236,I60765,);
not I_3416 (I60773,I60765);
nor I_3417 (I60222,I60773,I60485);
not I_3418 (I60831,I2690);
DFFARX1 I_3419 (I136167,I2683,I60831,I60857,);
DFFARX1 I_3420 (I60857,I2683,I60831,I60874,);
not I_3421 (I60823,I60874);
not I_3422 (I60896,I60857);
DFFARX1 I_3423 (I136155,I2683,I60831,I60922,);
not I_3424 (I60930,I60922);
and I_3425 (I60947,I60896,I136164);
not I_3426 (I60964,I136161);
nand I_3427 (I60981,I60964,I136164);
not I_3428 (I60998,I136152);
nor I_3429 (I61015,I60998,I136158);
nand I_3430 (I61032,I61015,I136143);
nor I_3431 (I61049,I61032,I60981);
DFFARX1 I_3432 (I61049,I2683,I60831,I60799,);
not I_3433 (I61080,I61032);
not I_3434 (I61097,I136158);
nand I_3435 (I61114,I61097,I136164);
nor I_3436 (I61131,I136158,I136161);
nand I_3437 (I60811,I60947,I61131);
nand I_3438 (I60805,I60896,I136158);
nand I_3439 (I61176,I60998,I136143);
DFFARX1 I_3440 (I61176,I2683,I60831,I60820,);
DFFARX1 I_3441 (I61176,I2683,I60831,I60814,);
not I_3442 (I61221,I136143);
nor I_3443 (I61238,I61221,I136149);
and I_3444 (I61255,I61238,I136146);
or I_3445 (I61272,I61255,I136170);
DFFARX1 I_3446 (I61272,I2683,I60831,I61298,);
nand I_3447 (I61306,I61298,I60964);
nor I_3448 (I60808,I61306,I61114);
nor I_3449 (I60802,I61298,I60930);
DFFARX1 I_3450 (I61298,I2683,I60831,I61360,);
not I_3451 (I61368,I61360);
nor I_3452 (I60817,I61368,I61080);
not I_3453 (I61426,I2690);
DFFARX1 I_3454 (I1396,I2683,I61426,I61452,);
DFFARX1 I_3455 (I61452,I2683,I61426,I61469,);
not I_3456 (I61418,I61469);
not I_3457 (I61491,I61452);
DFFARX1 I_3458 (I1836,I2683,I61426,I61517,);
not I_3459 (I61525,I61517);
and I_3460 (I61542,I61491,I1452);
not I_3461 (I61559,I2260);
nand I_3462 (I61576,I61559,I1452);
not I_3463 (I61593,I2556);
nor I_3464 (I61610,I61593,I2292);
nand I_3465 (I61627,I61610,I1964);
nor I_3466 (I61644,I61627,I61576);
DFFARX1 I_3467 (I61644,I2683,I61426,I61394,);
not I_3468 (I61675,I61627);
not I_3469 (I61692,I2292);
nand I_3470 (I61709,I61692,I1452);
nor I_3471 (I61726,I2292,I2260);
nand I_3472 (I61406,I61542,I61726);
nand I_3473 (I61400,I61491,I2292);
nand I_3474 (I61771,I61593,I1668);
DFFARX1 I_3475 (I61771,I2683,I61426,I61415,);
DFFARX1 I_3476 (I61771,I2683,I61426,I61409,);
not I_3477 (I61816,I1668);
nor I_3478 (I61833,I61816,I2652);
and I_3479 (I61850,I61833,I1588);
or I_3480 (I61867,I61850,I1380);
DFFARX1 I_3481 (I61867,I2683,I61426,I61893,);
nand I_3482 (I61901,I61893,I61559);
nor I_3483 (I61403,I61901,I61709);
nor I_3484 (I61397,I61893,I61525);
DFFARX1 I_3485 (I61893,I2683,I61426,I61955,);
not I_3486 (I61963,I61955);
nor I_3487 (I61412,I61963,I61675);
not I_3488 (I62021,I2690);
DFFARX1 I_3489 (I42567,I2683,I62021,I62047,);
DFFARX1 I_3490 (I62047,I2683,I62021,I62064,);
not I_3491 (I62013,I62064);
not I_3492 (I62086,I62047);
DFFARX1 I_3493 (I42561,I2683,I62021,I62112,);
not I_3494 (I62120,I62112);
and I_3495 (I62137,I62086,I42558);
not I_3496 (I62154,I42579);
nand I_3497 (I62171,I62154,I42558);
not I_3498 (I62188,I42573);
nor I_3499 (I62205,I62188,I42564);
nand I_3500 (I62222,I62205,I42570);
nor I_3501 (I62239,I62222,I62171);
DFFARX1 I_3502 (I62239,I2683,I62021,I61989,);
not I_3503 (I62270,I62222);
not I_3504 (I62287,I42564);
nand I_3505 (I62304,I62287,I42558);
nor I_3506 (I62321,I42564,I42579);
nand I_3507 (I62001,I62137,I62321);
nand I_3508 (I61995,I62086,I42564);
nand I_3509 (I62366,I62188,I42558);
DFFARX1 I_3510 (I62366,I2683,I62021,I62010,);
DFFARX1 I_3511 (I62366,I2683,I62021,I62004,);
not I_3512 (I62411,I42558);
nor I_3513 (I62428,I62411,I42576);
and I_3514 (I62445,I62428,I42582);
or I_3515 (I62462,I62445,I42561);
DFFARX1 I_3516 (I62462,I2683,I62021,I62488,);
nand I_3517 (I62496,I62488,I62154);
nor I_3518 (I61998,I62496,I62304);
nor I_3519 (I61992,I62488,I62120);
DFFARX1 I_3520 (I62488,I2683,I62021,I62550,);
not I_3521 (I62558,I62550);
nor I_3522 (I62007,I62558,I62270);
not I_3523 (I62616,I2690);
DFFARX1 I_3524 (I236013,I2683,I62616,I62642,);
DFFARX1 I_3525 (I62642,I2683,I62616,I62659,);
not I_3526 (I62608,I62659);
not I_3527 (I62681,I62642);
DFFARX1 I_3528 (I236010,I2683,I62616,I62707,);
not I_3529 (I62715,I62707);
and I_3530 (I62732,I62681,I236016);
not I_3531 (I62749,I236001);
nand I_3532 (I62766,I62749,I236016);
not I_3533 (I62783,I236004);
nor I_3534 (I62800,I62783,I236025);
nand I_3535 (I62817,I62800,I236022);
nor I_3536 (I62834,I62817,I62766);
DFFARX1 I_3537 (I62834,I2683,I62616,I62584,);
not I_3538 (I62865,I62817);
not I_3539 (I62882,I236025);
nand I_3540 (I62899,I62882,I236016);
nor I_3541 (I62916,I236025,I236001);
nand I_3542 (I62596,I62732,I62916);
nand I_3543 (I62590,I62681,I236025);
nand I_3544 (I62961,I62783,I236001);
DFFARX1 I_3545 (I62961,I2683,I62616,I62605,);
DFFARX1 I_3546 (I62961,I2683,I62616,I62599,);
not I_3547 (I63006,I236001);
nor I_3548 (I63023,I63006,I236007);
and I_3549 (I63040,I63023,I236019);
or I_3550 (I63057,I63040,I236004);
DFFARX1 I_3551 (I63057,I2683,I62616,I63083,);
nand I_3552 (I63091,I63083,I62749);
nor I_3553 (I62593,I63091,I62899);
nor I_3554 (I62587,I63083,I62715);
DFFARX1 I_3555 (I63083,I2683,I62616,I63145,);
not I_3556 (I63153,I63145);
nor I_3557 (I62602,I63153,I62865);
not I_3558 (I63211,I2690);
DFFARX1 I_3559 (I6219,I2683,I63211,I63237,);
DFFARX1 I_3560 (I63237,I2683,I63211,I63254,);
not I_3561 (I63203,I63254);
not I_3562 (I63276,I63237);
DFFARX1 I_3563 (I6195,I2683,I63211,I63302,);
not I_3564 (I63310,I63302);
and I_3565 (I63327,I63276,I6210);
not I_3566 (I63344,I6198);
nand I_3567 (I63361,I63344,I6210);
not I_3568 (I63378,I6201);
nor I_3569 (I63395,I63378,I6213);
nand I_3570 (I63412,I63395,I6204);
nor I_3571 (I63429,I63412,I63361);
DFFARX1 I_3572 (I63429,I2683,I63211,I63179,);
not I_3573 (I63460,I63412);
not I_3574 (I63477,I6213);
nand I_3575 (I63494,I63477,I6210);
nor I_3576 (I63511,I6213,I6198);
nand I_3577 (I63191,I63327,I63511);
nand I_3578 (I63185,I63276,I6213);
nand I_3579 (I63556,I63378,I6207);
DFFARX1 I_3580 (I63556,I2683,I63211,I63200,);
DFFARX1 I_3581 (I63556,I2683,I63211,I63194,);
not I_3582 (I63601,I6207);
nor I_3583 (I63618,I63601,I6198);
and I_3584 (I63635,I63618,I6195);
or I_3585 (I63652,I63635,I6216);
DFFARX1 I_3586 (I63652,I2683,I63211,I63678,);
nand I_3587 (I63686,I63678,I63344);
nor I_3588 (I63188,I63686,I63494);
nor I_3589 (I63182,I63678,I63310);
DFFARX1 I_3590 (I63678,I2683,I63211,I63740,);
not I_3591 (I63748,I63740);
nor I_3592 (I63197,I63748,I63460);
not I_3593 (I63806,I2690);
DFFARX1 I_3594 (I197865,I2683,I63806,I63832,);
DFFARX1 I_3595 (I63832,I2683,I63806,I63849,);
not I_3596 (I63798,I63849);
not I_3597 (I63871,I63832);
DFFARX1 I_3598 (I197862,I2683,I63806,I63897,);
not I_3599 (I63905,I63897);
and I_3600 (I63922,I63871,I197868);
not I_3601 (I63939,I197853);
nand I_3602 (I63956,I63939,I197868);
not I_3603 (I63973,I197856);
nor I_3604 (I63990,I63973,I197877);
nand I_3605 (I64007,I63990,I197874);
nor I_3606 (I64024,I64007,I63956);
DFFARX1 I_3607 (I64024,I2683,I63806,I63774,);
not I_3608 (I64055,I64007);
not I_3609 (I64072,I197877);
nand I_3610 (I64089,I64072,I197868);
nor I_3611 (I64106,I197877,I197853);
nand I_3612 (I63786,I63922,I64106);
nand I_3613 (I63780,I63871,I197877);
nand I_3614 (I64151,I63973,I197853);
DFFARX1 I_3615 (I64151,I2683,I63806,I63795,);
DFFARX1 I_3616 (I64151,I2683,I63806,I63789,);
not I_3617 (I64196,I197853);
nor I_3618 (I64213,I64196,I197859);
and I_3619 (I64230,I64213,I197871);
or I_3620 (I64247,I64230,I197856);
DFFARX1 I_3621 (I64247,I2683,I63806,I64273,);
nand I_3622 (I64281,I64273,I63939);
nor I_3623 (I63783,I64281,I64089);
nor I_3624 (I63777,I64273,I63905);
DFFARX1 I_3625 (I64273,I2683,I63806,I64335,);
not I_3626 (I64343,I64335);
nor I_3627 (I63792,I64343,I64055);
not I_3628 (I64401,I2690);
DFFARX1 I_3629 (I372495,I2683,I64401,I64427,);
DFFARX1 I_3630 (I64427,I2683,I64401,I64444,);
not I_3631 (I64393,I64444);
not I_3632 (I64466,I64427);
DFFARX1 I_3633 (I372480,I2683,I64401,I64492,);
not I_3634 (I64500,I64492);
and I_3635 (I64517,I64466,I372498);
not I_3636 (I64534,I372480);
nand I_3637 (I64551,I64534,I372498);
not I_3638 (I64568,I372501);
nor I_3639 (I64585,I64568,I372492);
nand I_3640 (I64602,I64585,I372489);
nor I_3641 (I64619,I64602,I64551);
DFFARX1 I_3642 (I64619,I2683,I64401,I64369,);
not I_3643 (I64650,I64602);
not I_3644 (I64667,I372492);
nand I_3645 (I64684,I64667,I372498);
nor I_3646 (I64701,I372492,I372480);
nand I_3647 (I64381,I64517,I64701);
nand I_3648 (I64375,I64466,I372492);
nand I_3649 (I64746,I64568,I372486);
DFFARX1 I_3650 (I64746,I2683,I64401,I64390,);
DFFARX1 I_3651 (I64746,I2683,I64401,I64384,);
not I_3652 (I64791,I372486);
nor I_3653 (I64808,I64791,I372477);
and I_3654 (I64825,I64808,I372483);
or I_3655 (I64842,I64825,I372477);
DFFARX1 I_3656 (I64842,I2683,I64401,I64868,);
nand I_3657 (I64876,I64868,I64534);
nor I_3658 (I64378,I64876,I64684);
nor I_3659 (I64372,I64868,I64500);
DFFARX1 I_3660 (I64868,I2683,I64401,I64930,);
not I_3661 (I64938,I64930);
nor I_3662 (I64387,I64938,I64650);
not I_3663 (I64996,I2690);
DFFARX1 I_3664 (I222141,I2683,I64996,I65022,);
DFFARX1 I_3665 (I65022,I2683,I64996,I65039,);
not I_3666 (I64988,I65039);
not I_3667 (I65061,I65022);
DFFARX1 I_3668 (I222138,I2683,I64996,I65087,);
not I_3669 (I65095,I65087);
and I_3670 (I65112,I65061,I222144);
not I_3671 (I65129,I222129);
nand I_3672 (I65146,I65129,I222144);
not I_3673 (I65163,I222132);
nor I_3674 (I65180,I65163,I222153);
nand I_3675 (I65197,I65180,I222150);
nor I_3676 (I65214,I65197,I65146);
DFFARX1 I_3677 (I65214,I2683,I64996,I64964,);
not I_3678 (I65245,I65197);
not I_3679 (I65262,I222153);
nand I_3680 (I65279,I65262,I222144);
nor I_3681 (I65296,I222153,I222129);
nand I_3682 (I64976,I65112,I65296);
nand I_3683 (I64970,I65061,I222153);
nand I_3684 (I65341,I65163,I222129);
DFFARX1 I_3685 (I65341,I2683,I64996,I64985,);
DFFARX1 I_3686 (I65341,I2683,I64996,I64979,);
not I_3687 (I65386,I222129);
nor I_3688 (I65403,I65386,I222135);
and I_3689 (I65420,I65403,I222147);
or I_3690 (I65437,I65420,I222132);
DFFARX1 I_3691 (I65437,I2683,I64996,I65463,);
nand I_3692 (I65471,I65463,I65129);
nor I_3693 (I64973,I65471,I65279);
nor I_3694 (I64967,I65463,I65095);
DFFARX1 I_3695 (I65463,I2683,I64996,I65525,);
not I_3696 (I65533,I65525);
nor I_3697 (I64982,I65533,I65245);
not I_3698 (I65591,I2690);
DFFARX1 I_3699 (I215205,I2683,I65591,I65617,);
DFFARX1 I_3700 (I65617,I2683,I65591,I65634,);
not I_3701 (I65583,I65634);
not I_3702 (I65656,I65617);
DFFARX1 I_3703 (I215202,I2683,I65591,I65682,);
not I_3704 (I65690,I65682);
and I_3705 (I65707,I65656,I215208);
not I_3706 (I65724,I215193);
nand I_3707 (I65741,I65724,I215208);
not I_3708 (I65758,I215196);
nor I_3709 (I65775,I65758,I215217);
nand I_3710 (I65792,I65775,I215214);
nor I_3711 (I65809,I65792,I65741);
DFFARX1 I_3712 (I65809,I2683,I65591,I65559,);
not I_3713 (I65840,I65792);
not I_3714 (I65857,I215217);
nand I_3715 (I65874,I65857,I215208);
nor I_3716 (I65891,I215217,I215193);
nand I_3717 (I65571,I65707,I65891);
nand I_3718 (I65565,I65656,I215217);
nand I_3719 (I65936,I65758,I215193);
DFFARX1 I_3720 (I65936,I2683,I65591,I65580,);
DFFARX1 I_3721 (I65936,I2683,I65591,I65574,);
not I_3722 (I65981,I215193);
nor I_3723 (I65998,I65981,I215199);
and I_3724 (I66015,I65998,I215211);
or I_3725 (I66032,I66015,I215196);
DFFARX1 I_3726 (I66032,I2683,I65591,I66058,);
nand I_3727 (I66066,I66058,I65724);
nor I_3728 (I65568,I66066,I65874);
nor I_3729 (I65562,I66058,I65690);
DFFARX1 I_3730 (I66058,I2683,I65591,I66120,);
not I_3731 (I66128,I66120);
nor I_3732 (I65577,I66128,I65840);
not I_3733 (I66186,I2690);
DFFARX1 I_3734 (I153575,I2683,I66186,I66212,);
DFFARX1 I_3735 (I66212,I2683,I66186,I66229,);
not I_3736 (I66178,I66229);
not I_3737 (I66251,I66212);
DFFARX1 I_3738 (I153563,I2683,I66186,I66277,);
not I_3739 (I66285,I66277);
and I_3740 (I66302,I66251,I153572);
not I_3741 (I66319,I153569);
nand I_3742 (I66336,I66319,I153572);
not I_3743 (I66353,I153560);
nor I_3744 (I66370,I66353,I153566);
nand I_3745 (I66387,I66370,I153551);
nor I_3746 (I66404,I66387,I66336);
DFFARX1 I_3747 (I66404,I2683,I66186,I66154,);
not I_3748 (I66435,I66387);
not I_3749 (I66452,I153566);
nand I_3750 (I66469,I66452,I153572);
nor I_3751 (I66486,I153566,I153569);
nand I_3752 (I66166,I66302,I66486);
nand I_3753 (I66160,I66251,I153566);
nand I_3754 (I66531,I66353,I153551);
DFFARX1 I_3755 (I66531,I2683,I66186,I66175,);
DFFARX1 I_3756 (I66531,I2683,I66186,I66169,);
not I_3757 (I66576,I153551);
nor I_3758 (I66593,I66576,I153557);
and I_3759 (I66610,I66593,I153554);
or I_3760 (I66627,I66610,I153578);
DFFARX1 I_3761 (I66627,I2683,I66186,I66653,);
nand I_3762 (I66661,I66653,I66319);
nor I_3763 (I66163,I66661,I66469);
nor I_3764 (I66157,I66653,I66285);
DFFARX1 I_3765 (I66653,I2683,I66186,I66715,);
not I_3766 (I66723,I66715);
nor I_3767 (I66172,I66723,I66435);
not I_3768 (I66781,I2690);
DFFARX1 I_3769 (I177060,I2683,I66781,I66807,);
DFFARX1 I_3770 (I66807,I2683,I66781,I66824,);
not I_3771 (I66773,I66824);
not I_3772 (I66846,I66807);
DFFARX1 I_3773 (I177051,I2683,I66781,I66872,);
not I_3774 (I66880,I66872);
and I_3775 (I66897,I66846,I177069);
not I_3776 (I66914,I177066);
nand I_3777 (I66931,I66914,I177069);
not I_3778 (I66948,I177045);
nor I_3779 (I66965,I66948,I177048);
nand I_3780 (I66982,I66965,I177057);
nor I_3781 (I66999,I66982,I66931);
DFFARX1 I_3782 (I66999,I2683,I66781,I66749,);
not I_3783 (I67030,I66982);
not I_3784 (I67047,I177048);
nand I_3785 (I67064,I67047,I177069);
nor I_3786 (I67081,I177048,I177066);
nand I_3787 (I66761,I66897,I67081);
nand I_3788 (I66755,I66846,I177048);
nand I_3789 (I67126,I66948,I177063);
DFFARX1 I_3790 (I67126,I2683,I66781,I66770,);
DFFARX1 I_3791 (I67126,I2683,I66781,I66764,);
not I_3792 (I67171,I177063);
nor I_3793 (I67188,I67171,I177045);
and I_3794 (I67205,I67188,I177054);
or I_3795 (I67222,I67205,I177048);
DFFARX1 I_3796 (I67222,I2683,I66781,I67248,);
nand I_3797 (I67256,I67248,I66914);
nor I_3798 (I66758,I67256,I67064);
nor I_3799 (I66752,I67248,I66880);
DFFARX1 I_3800 (I67248,I2683,I66781,I67310,);
not I_3801 (I67318,I67310);
nor I_3802 (I66767,I67318,I67030);
not I_3803 (I67376,I2690);
DFFARX1 I_3804 (I279485,I2683,I67376,I67402,);
DFFARX1 I_3805 (I67402,I2683,I67376,I67419,);
not I_3806 (I67368,I67419);
not I_3807 (I67441,I67402);
DFFARX1 I_3808 (I279494,I2683,I67376,I67467,);
not I_3809 (I67475,I67467);
and I_3810 (I67492,I67441,I279482);
not I_3811 (I67509,I279473);
nand I_3812 (I67526,I67509,I279482);
not I_3813 (I67543,I279479);
nor I_3814 (I67560,I67543,I279497);
nand I_3815 (I67577,I67560,I279470);
nor I_3816 (I67594,I67577,I67526);
DFFARX1 I_3817 (I67594,I2683,I67376,I67344,);
not I_3818 (I67625,I67577);
not I_3819 (I67642,I279497);
nand I_3820 (I67659,I67642,I279482);
nor I_3821 (I67676,I279497,I279473);
nand I_3822 (I67356,I67492,I67676);
nand I_3823 (I67350,I67441,I279497);
nand I_3824 (I67721,I67543,I279476);
DFFARX1 I_3825 (I67721,I2683,I67376,I67365,);
DFFARX1 I_3826 (I67721,I2683,I67376,I67359,);
not I_3827 (I67766,I279476);
nor I_3828 (I67783,I67766,I279488);
and I_3829 (I67800,I67783,I279470);
or I_3830 (I67817,I67800,I279491);
DFFARX1 I_3831 (I67817,I2683,I67376,I67843,);
nand I_3832 (I67851,I67843,I67509);
nor I_3833 (I67353,I67851,I67659);
nor I_3834 (I67347,I67843,I67475);
DFFARX1 I_3835 (I67843,I2683,I67376,I67905,);
not I_3836 (I67913,I67905);
nor I_3837 (I67362,I67913,I67625);
not I_3838 (I67971,I2690);
DFFARX1 I_3839 (I333683,I2683,I67971,I67997,);
DFFARX1 I_3840 (I67997,I2683,I67971,I68014,);
not I_3841 (I67963,I68014);
not I_3842 (I68036,I67997);
DFFARX1 I_3843 (I333683,I2683,I67971,I68062,);
not I_3844 (I68070,I68062);
and I_3845 (I68087,I68036,I333686);
not I_3846 (I68104,I333698);
nand I_3847 (I68121,I68104,I333686);
not I_3848 (I68138,I333704);
nor I_3849 (I68155,I68138,I333695);
nand I_3850 (I68172,I68155,I333701);
nor I_3851 (I68189,I68172,I68121);
DFFARX1 I_3852 (I68189,I2683,I67971,I67939,);
not I_3853 (I68220,I68172);
not I_3854 (I68237,I333695);
nand I_3855 (I68254,I68237,I333686);
nor I_3856 (I68271,I333695,I333698);
nand I_3857 (I67951,I68087,I68271);
nand I_3858 (I67945,I68036,I333695);
nand I_3859 (I68316,I68138,I333692);
DFFARX1 I_3860 (I68316,I2683,I67971,I67960,);
DFFARX1 I_3861 (I68316,I2683,I67971,I67954,);
not I_3862 (I68361,I333692);
nor I_3863 (I68378,I68361,I333689);
and I_3864 (I68395,I68378,I333707);
or I_3865 (I68412,I68395,I333686);
DFFARX1 I_3866 (I68412,I2683,I67971,I68438,);
nand I_3867 (I68446,I68438,I68104);
nor I_3868 (I67948,I68446,I68254);
nor I_3869 (I67942,I68438,I68070);
DFFARX1 I_3870 (I68438,I2683,I67971,I68500,);
not I_3871 (I68508,I68500);
nor I_3872 (I67957,I68508,I68220);
not I_3873 (I68566,I2690);
DFFARX1 I_3874 (I146503,I2683,I68566,I68592,);
DFFARX1 I_3875 (I68592,I2683,I68566,I68609,);
not I_3876 (I68558,I68609);
not I_3877 (I68631,I68592);
DFFARX1 I_3878 (I146491,I2683,I68566,I68657,);
not I_3879 (I68665,I68657);
and I_3880 (I68682,I68631,I146500);
not I_3881 (I68699,I146497);
nand I_3882 (I68716,I68699,I146500);
not I_3883 (I68733,I146488);
nor I_3884 (I68750,I68733,I146494);
nand I_3885 (I68767,I68750,I146479);
nor I_3886 (I68784,I68767,I68716);
DFFARX1 I_3887 (I68784,I2683,I68566,I68534,);
not I_3888 (I68815,I68767);
not I_3889 (I68832,I146494);
nand I_3890 (I68849,I68832,I146500);
nor I_3891 (I68866,I146494,I146497);
nand I_3892 (I68546,I68682,I68866);
nand I_3893 (I68540,I68631,I146494);
nand I_3894 (I68911,I68733,I146479);
DFFARX1 I_3895 (I68911,I2683,I68566,I68555,);
DFFARX1 I_3896 (I68911,I2683,I68566,I68549,);
not I_3897 (I68956,I146479);
nor I_3898 (I68973,I68956,I146485);
and I_3899 (I68990,I68973,I146482);
or I_3900 (I69007,I68990,I146506);
DFFARX1 I_3901 (I69007,I2683,I68566,I69033,);
nand I_3902 (I69041,I69033,I68699);
nor I_3903 (I68543,I69041,I68849);
nor I_3904 (I68537,I69033,I68665);
DFFARX1 I_3905 (I69033,I2683,I68566,I69095,);
not I_3906 (I69103,I69095);
nor I_3907 (I68552,I69103,I68815);
not I_3908 (I69161,I2690);
DFFARX1 I_3909 (I315445,I2683,I69161,I69187,);
DFFARX1 I_3910 (I69187,I2683,I69161,I69204,);
not I_3911 (I69153,I69204);
not I_3912 (I69226,I69187);
DFFARX1 I_3913 (I315454,I2683,I69161,I69252,);
not I_3914 (I69260,I69252);
and I_3915 (I69277,I69226,I315448);
not I_3916 (I69294,I315442);
nand I_3917 (I69311,I69294,I315448);
not I_3918 (I69328,I315457);
nor I_3919 (I69345,I69328,I315445);
nand I_3920 (I69362,I69345,I315451);
nor I_3921 (I69379,I69362,I69311);
DFFARX1 I_3922 (I69379,I2683,I69161,I69129,);
not I_3923 (I69410,I69362);
not I_3924 (I69427,I315445);
nand I_3925 (I69444,I69427,I315448);
nor I_3926 (I69461,I315445,I315442);
nand I_3927 (I69141,I69277,I69461);
nand I_3928 (I69135,I69226,I315445);
nand I_3929 (I69506,I69328,I315448);
DFFARX1 I_3930 (I69506,I2683,I69161,I69150,);
DFFARX1 I_3931 (I69506,I2683,I69161,I69144,);
not I_3932 (I69551,I315448);
nor I_3933 (I69568,I69551,I315463);
and I_3934 (I69585,I69568,I315460);
or I_3935 (I69602,I69585,I315442);
DFFARX1 I_3936 (I69602,I2683,I69161,I69628,);
nand I_3937 (I69636,I69628,I69294);
nor I_3938 (I69138,I69636,I69444);
nor I_3939 (I69132,I69628,I69260);
DFFARX1 I_3940 (I69628,I2683,I69161,I69690,);
not I_3941 (I69698,I69690);
nor I_3942 (I69147,I69698,I69410);
not I_3943 (I69756,I2690);
DFFARX1 I_3944 (I220985,I2683,I69756,I69782,);
DFFARX1 I_3945 (I69782,I2683,I69756,I69799,);
not I_3946 (I69748,I69799);
not I_3947 (I69821,I69782);
DFFARX1 I_3948 (I220982,I2683,I69756,I69847,);
not I_3949 (I69855,I69847);
and I_3950 (I69872,I69821,I220988);
not I_3951 (I69889,I220973);
nand I_3952 (I69906,I69889,I220988);
not I_3953 (I69923,I220976);
nor I_3954 (I69940,I69923,I220997);
nand I_3955 (I69957,I69940,I220994);
nor I_3956 (I69974,I69957,I69906);
DFFARX1 I_3957 (I69974,I2683,I69756,I69724,);
not I_3958 (I70005,I69957);
not I_3959 (I70022,I220997);
nand I_3960 (I70039,I70022,I220988);
nor I_3961 (I70056,I220997,I220973);
nand I_3962 (I69736,I69872,I70056);
nand I_3963 (I69730,I69821,I220997);
nand I_3964 (I70101,I69923,I220973);
DFFARX1 I_3965 (I70101,I2683,I69756,I69745,);
DFFARX1 I_3966 (I70101,I2683,I69756,I69739,);
not I_3967 (I70146,I220973);
nor I_3968 (I70163,I70146,I220979);
and I_3969 (I70180,I70163,I220991);
or I_3970 (I70197,I70180,I220976);
DFFARX1 I_3971 (I70197,I2683,I69756,I70223,);
nand I_3972 (I70231,I70223,I69889);
nor I_3973 (I69733,I70231,I70039);
nor I_3974 (I69727,I70223,I69855);
DFFARX1 I_3975 (I70223,I2683,I69756,I70285,);
not I_3976 (I70293,I70285);
nor I_3977 (I69742,I70293,I70005);
not I_3978 (I70351,I2690);
DFFARX1 I_3979 (I229655,I2683,I70351,I70377,);
DFFARX1 I_3980 (I70377,I2683,I70351,I70394,);
not I_3981 (I70343,I70394);
not I_3982 (I70416,I70377);
DFFARX1 I_3983 (I229652,I2683,I70351,I70442,);
not I_3984 (I70450,I70442);
and I_3985 (I70467,I70416,I229658);
not I_3986 (I70484,I229643);
nand I_3987 (I70501,I70484,I229658);
not I_3988 (I70518,I229646);
nor I_3989 (I70535,I70518,I229667);
nand I_3990 (I70552,I70535,I229664);
nor I_3991 (I70569,I70552,I70501);
DFFARX1 I_3992 (I70569,I2683,I70351,I70319,);
not I_3993 (I70600,I70552);
not I_3994 (I70617,I229667);
nand I_3995 (I70634,I70617,I229658);
nor I_3996 (I70651,I229667,I229643);
nand I_3997 (I70331,I70467,I70651);
nand I_3998 (I70325,I70416,I229667);
nand I_3999 (I70696,I70518,I229643);
DFFARX1 I_4000 (I70696,I2683,I70351,I70340,);
DFFARX1 I_4001 (I70696,I2683,I70351,I70334,);
not I_4002 (I70741,I229643);
nor I_4003 (I70758,I70741,I229649);
and I_4004 (I70775,I70758,I229661);
or I_4005 (I70792,I70775,I229646);
DFFARX1 I_4006 (I70792,I2683,I70351,I70818,);
nand I_4007 (I70826,I70818,I70484);
nor I_4008 (I70328,I70826,I70634);
nor I_4009 (I70322,I70818,I70450);
DFFARX1 I_4010 (I70818,I2683,I70351,I70880,);
not I_4011 (I70888,I70880);
nor I_4012 (I70337,I70888,I70600);
not I_4013 (I70946,I2690);
DFFARX1 I_4014 (I157626,I2683,I70946,I70972,);
DFFARX1 I_4015 (I70972,I2683,I70946,I70989,);
not I_4016 (I70938,I70989);
not I_4017 (I71011,I70972);
DFFARX1 I_4018 (I157620,I2683,I70946,I71037,);
not I_4019 (I71045,I71037);
and I_4020 (I71062,I71011,I157635);
not I_4021 (I71079,I157632);
nand I_4022 (I71096,I71079,I157635);
not I_4023 (I71113,I157623);
nor I_4024 (I71130,I71113,I157614);
nand I_4025 (I71147,I71130,I157617);
nor I_4026 (I71164,I71147,I71096);
DFFARX1 I_4027 (I71164,I2683,I70946,I70914,);
not I_4028 (I71195,I71147);
not I_4029 (I71212,I157614);
nand I_4030 (I71229,I71212,I157635);
nor I_4031 (I71246,I157614,I157632);
nand I_4032 (I70926,I71062,I71246);
nand I_4033 (I70920,I71011,I157614);
nand I_4034 (I71291,I71113,I157638);
DFFARX1 I_4035 (I71291,I2683,I70946,I70935,);
DFFARX1 I_4036 (I71291,I2683,I70946,I70929,);
not I_4037 (I71336,I157638);
nor I_4038 (I71353,I71336,I157629);
and I_4039 (I71370,I71353,I157614);
or I_4040 (I71387,I71370,I157617);
DFFARX1 I_4041 (I71387,I2683,I70946,I71413,);
nand I_4042 (I71421,I71413,I71079);
nor I_4043 (I70923,I71421,I71229);
nor I_4044 (I70917,I71413,I71045);
DFFARX1 I_4045 (I71413,I2683,I70946,I71475,);
not I_4046 (I71483,I71475);
nor I_4047 (I70932,I71483,I71195);
not I_4048 (I71541,I2690);
DFFARX1 I_4049 (I360849,I2683,I71541,I71567,);
DFFARX1 I_4050 (I71567,I2683,I71541,I71584,);
not I_4051 (I71533,I71584);
not I_4052 (I71606,I71567);
DFFARX1 I_4053 (I360849,I2683,I71541,I71632,);
not I_4054 (I71640,I71632);
and I_4055 (I71657,I71606,I360852);
not I_4056 (I71674,I360864);
nand I_4057 (I71691,I71674,I360852);
not I_4058 (I71708,I360870);
nor I_4059 (I71725,I71708,I360861);
nand I_4060 (I71742,I71725,I360867);
nor I_4061 (I71759,I71742,I71691);
DFFARX1 I_4062 (I71759,I2683,I71541,I71509,);
not I_4063 (I71790,I71742);
not I_4064 (I71807,I360861);
nand I_4065 (I71824,I71807,I360852);
nor I_4066 (I71841,I360861,I360864);
nand I_4067 (I71521,I71657,I71841);
nand I_4068 (I71515,I71606,I360861);
nand I_4069 (I71886,I71708,I360858);
DFFARX1 I_4070 (I71886,I2683,I71541,I71530,);
DFFARX1 I_4071 (I71886,I2683,I71541,I71524,);
not I_4072 (I71931,I360858);
nor I_4073 (I71948,I71931,I360855);
and I_4074 (I71965,I71948,I360873);
or I_4075 (I71982,I71965,I360852);
DFFARX1 I_4076 (I71982,I2683,I71541,I72008,);
nand I_4077 (I72016,I72008,I71674);
nor I_4078 (I71518,I72016,I71824);
nor I_4079 (I71512,I72008,I71640);
DFFARX1 I_4080 (I72008,I2683,I71541,I72070,);
not I_4081 (I72078,I72070);
nor I_4082 (I71527,I72078,I71790);
not I_4083 (I72136,I2690);
DFFARX1 I_4084 (I181106,I2683,I72136,I72162,);
DFFARX1 I_4085 (I72162,I2683,I72136,I72179,);
not I_4086 (I72128,I72179);
not I_4087 (I72201,I72162);
DFFARX1 I_4088 (I181097,I2683,I72136,I72227,);
not I_4089 (I72235,I72227);
and I_4090 (I72252,I72201,I181115);
not I_4091 (I72269,I181112);
nand I_4092 (I72286,I72269,I181115);
not I_4093 (I72303,I181091);
nor I_4094 (I72320,I72303,I181094);
nand I_4095 (I72337,I72320,I181103);
nor I_4096 (I72354,I72337,I72286);
DFFARX1 I_4097 (I72354,I2683,I72136,I72104,);
not I_4098 (I72385,I72337);
not I_4099 (I72402,I181094);
nand I_4100 (I72419,I72402,I181115);
nor I_4101 (I72436,I181094,I181112);
nand I_4102 (I72116,I72252,I72436);
nand I_4103 (I72110,I72201,I181094);
nand I_4104 (I72481,I72303,I181109);
DFFARX1 I_4105 (I72481,I2683,I72136,I72125,);
DFFARX1 I_4106 (I72481,I2683,I72136,I72119,);
not I_4107 (I72526,I181109);
nor I_4108 (I72543,I72526,I181091);
and I_4109 (I72560,I72543,I181100);
or I_4110 (I72577,I72560,I181094);
DFFARX1 I_4111 (I72577,I2683,I72136,I72603,);
nand I_4112 (I72611,I72603,I72269);
nor I_4113 (I72113,I72611,I72419);
nor I_4114 (I72107,I72603,I72235);
DFFARX1 I_4115 (I72603,I2683,I72136,I72665,);
not I_4116 (I72673,I72665);
nor I_4117 (I72122,I72673,I72385);
not I_4118 (I72731,I2690);
DFFARX1 I_4119 (I121098,I2683,I72731,I72757,);
DFFARX1 I_4120 (I72757,I2683,I72731,I72774,);
not I_4121 (I72723,I72774);
not I_4122 (I72796,I72757);
DFFARX1 I_4123 (I121113,I2683,I72731,I72822,);
not I_4124 (I72830,I72822);
and I_4125 (I72847,I72796,I121110);
not I_4126 (I72864,I121098);
nand I_4127 (I72881,I72864,I121110);
not I_4128 (I72898,I121107);
nor I_4129 (I72915,I72898,I121122);
nand I_4130 (I72932,I72915,I121119);
nor I_4131 (I72949,I72932,I72881);
DFFARX1 I_4132 (I72949,I2683,I72731,I72699,);
not I_4133 (I72980,I72932);
not I_4134 (I72997,I121122);
nand I_4135 (I73014,I72997,I121110);
nor I_4136 (I73031,I121122,I121098);
nand I_4137 (I72711,I72847,I73031);
nand I_4138 (I72705,I72796,I121122);
nand I_4139 (I73076,I72898,I121116);
DFFARX1 I_4140 (I73076,I2683,I72731,I72720,);
DFFARX1 I_4141 (I73076,I2683,I72731,I72714,);
not I_4142 (I73121,I121116);
nor I_4143 (I73138,I73121,I121104);
and I_4144 (I73155,I73138,I121125);
or I_4145 (I73172,I73155,I121101);
DFFARX1 I_4146 (I73172,I2683,I72731,I73198,);
nand I_4147 (I73206,I73198,I72864);
nor I_4148 (I72708,I73206,I73014);
nor I_4149 (I72702,I73198,I72830);
DFFARX1 I_4150 (I73198,I2683,I72731,I73260,);
not I_4151 (I73268,I73260);
nor I_4152 (I72717,I73268,I72980);
not I_4153 (I73326,I2690);
DFFARX1 I_4154 (I282715,I2683,I73326,I73352,);
DFFARX1 I_4155 (I73352,I2683,I73326,I73369,);
not I_4156 (I73318,I73369);
not I_4157 (I73391,I73352);
DFFARX1 I_4158 (I282724,I2683,I73326,I73417,);
not I_4159 (I73425,I73417);
and I_4160 (I73442,I73391,I282712);
not I_4161 (I73459,I282703);
nand I_4162 (I73476,I73459,I282712);
not I_4163 (I73493,I282709);
nor I_4164 (I73510,I73493,I282727);
nand I_4165 (I73527,I73510,I282700);
nor I_4166 (I73544,I73527,I73476);
DFFARX1 I_4167 (I73544,I2683,I73326,I73294,);
not I_4168 (I73575,I73527);
not I_4169 (I73592,I282727);
nand I_4170 (I73609,I73592,I282712);
nor I_4171 (I73626,I282727,I282703);
nand I_4172 (I73306,I73442,I73626);
nand I_4173 (I73300,I73391,I282727);
nand I_4174 (I73671,I73493,I282706);
DFFARX1 I_4175 (I73671,I2683,I73326,I73315,);
DFFARX1 I_4176 (I73671,I2683,I73326,I73309,);
not I_4177 (I73716,I282706);
nor I_4178 (I73733,I73716,I282718);
and I_4179 (I73750,I73733,I282700);
or I_4180 (I73767,I73750,I282721);
DFFARX1 I_4181 (I73767,I2683,I73326,I73793,);
nand I_4182 (I73801,I73793,I73459);
nor I_4183 (I73303,I73801,I73609);
nor I_4184 (I73297,I73793,I73425);
DFFARX1 I_4185 (I73793,I2683,I73326,I73855,);
not I_4186 (I73863,I73855);
nor I_4187 (I73312,I73863,I73575);
not I_4188 (I73921,I2690);
DFFARX1 I_4189 (I367599,I2683,I73921,I73947,);
DFFARX1 I_4190 (I73947,I2683,I73921,I73964,);
not I_4191 (I73913,I73964);
not I_4192 (I73986,I73947);
DFFARX1 I_4193 (I367584,I2683,I73921,I74012,);
not I_4194 (I74020,I74012);
and I_4195 (I74037,I73986,I367602);
not I_4196 (I74054,I367584);
nand I_4197 (I74071,I74054,I367602);
not I_4198 (I74088,I367605);
nor I_4199 (I74105,I74088,I367596);
nand I_4200 (I74122,I74105,I367593);
nor I_4201 (I74139,I74122,I74071);
DFFARX1 I_4202 (I74139,I2683,I73921,I73889,);
not I_4203 (I74170,I74122);
not I_4204 (I74187,I367596);
nand I_4205 (I74204,I74187,I367602);
nor I_4206 (I74221,I367596,I367584);
nand I_4207 (I73901,I74037,I74221);
nand I_4208 (I73895,I73986,I367596);
nand I_4209 (I74266,I74088,I367590);
DFFARX1 I_4210 (I74266,I2683,I73921,I73910,);
DFFARX1 I_4211 (I74266,I2683,I73921,I73904,);
not I_4212 (I74311,I367590);
nor I_4213 (I74328,I74311,I367581);
and I_4214 (I74345,I74328,I367587);
or I_4215 (I74362,I74345,I367581);
DFFARX1 I_4216 (I74362,I2683,I73921,I74388,);
nand I_4217 (I74396,I74388,I74054);
nor I_4218 (I73898,I74396,I74204);
nor I_4219 (I73892,I74388,I74020);
DFFARX1 I_4220 (I74388,I2683,I73921,I74450,);
not I_4221 (I74458,I74450);
nor I_4222 (I73907,I74458,I74170);
not I_4223 (I74516,I2690);
DFFARX1 I_4224 (I216939,I2683,I74516,I74542,);
DFFARX1 I_4225 (I74542,I2683,I74516,I74559,);
not I_4226 (I74508,I74559);
not I_4227 (I74581,I74542);
DFFARX1 I_4228 (I216936,I2683,I74516,I74607,);
not I_4229 (I74615,I74607);
and I_4230 (I74632,I74581,I216942);
not I_4231 (I74649,I216927);
nand I_4232 (I74666,I74649,I216942);
not I_4233 (I74683,I216930);
nor I_4234 (I74700,I74683,I216951);
nand I_4235 (I74717,I74700,I216948);
nor I_4236 (I74734,I74717,I74666);
DFFARX1 I_4237 (I74734,I2683,I74516,I74484,);
not I_4238 (I74765,I74717);
not I_4239 (I74782,I216951);
nand I_4240 (I74799,I74782,I216942);
nor I_4241 (I74816,I216951,I216927);
nand I_4242 (I74496,I74632,I74816);
nand I_4243 (I74490,I74581,I216951);
nand I_4244 (I74861,I74683,I216927);
DFFARX1 I_4245 (I74861,I2683,I74516,I74505,);
DFFARX1 I_4246 (I74861,I2683,I74516,I74499,);
not I_4247 (I74906,I216927);
nor I_4248 (I74923,I74906,I216933);
and I_4249 (I74940,I74923,I216945);
or I_4250 (I74957,I74940,I216930);
DFFARX1 I_4251 (I74957,I2683,I74516,I74983,);
nand I_4252 (I74991,I74983,I74649);
nor I_4253 (I74493,I74991,I74799);
nor I_4254 (I74487,I74983,I74615);
DFFARX1 I_4255 (I74983,I2683,I74516,I75045,);
not I_4256 (I75053,I75045);
nor I_4257 (I74502,I75053,I74765);
not I_4258 (I75111,I2690);
DFFARX1 I_4259 (I309201,I2683,I75111,I75137,);
DFFARX1 I_4260 (I75137,I2683,I75111,I75154,);
not I_4261 (I75103,I75154);
not I_4262 (I75176,I75137);
DFFARX1 I_4263 (I309210,I2683,I75111,I75202,);
not I_4264 (I75210,I75202);
and I_4265 (I75227,I75176,I309198);
not I_4266 (I75244,I309189);
nand I_4267 (I75261,I75244,I309198);
not I_4268 (I75278,I309195);
nor I_4269 (I75295,I75278,I309213);
nand I_4270 (I75312,I75295,I309186);
nor I_4271 (I75329,I75312,I75261);
DFFARX1 I_4272 (I75329,I2683,I75111,I75079,);
not I_4273 (I75360,I75312);
not I_4274 (I75377,I309213);
nand I_4275 (I75394,I75377,I309198);
nor I_4276 (I75411,I309213,I309189);
nand I_4277 (I75091,I75227,I75411);
nand I_4278 (I75085,I75176,I309213);
nand I_4279 (I75456,I75278,I309192);
DFFARX1 I_4280 (I75456,I2683,I75111,I75100,);
DFFARX1 I_4281 (I75456,I2683,I75111,I75094,);
not I_4282 (I75501,I309192);
nor I_4283 (I75518,I75501,I309204);
and I_4284 (I75535,I75518,I309186);
or I_4285 (I75552,I75535,I309207);
DFFARX1 I_4286 (I75552,I2683,I75111,I75578,);
nand I_4287 (I75586,I75578,I75244);
nor I_4288 (I75088,I75586,I75394);
nor I_4289 (I75082,I75578,I75210);
DFFARX1 I_4290 (I75578,I2683,I75111,I75640,);
not I_4291 (I75648,I75640);
nor I_4292 (I75097,I75648,I75360);
not I_4293 (I75706,I2690);
DFFARX1 I_4294 (I112139,I2683,I75706,I75732,);
DFFARX1 I_4295 (I75732,I2683,I75706,I75749,);
not I_4296 (I75698,I75749);
not I_4297 (I75771,I75732);
DFFARX1 I_4298 (I112154,I2683,I75706,I75797,);
not I_4299 (I75805,I75797);
and I_4300 (I75822,I75771,I112151);
not I_4301 (I75839,I112139);
nand I_4302 (I75856,I75839,I112151);
not I_4303 (I75873,I112148);
nor I_4304 (I75890,I75873,I112163);
nand I_4305 (I75907,I75890,I112160);
nor I_4306 (I75924,I75907,I75856);
DFFARX1 I_4307 (I75924,I2683,I75706,I75674,);
not I_4308 (I75955,I75907);
not I_4309 (I75972,I112163);
nand I_4310 (I75989,I75972,I112151);
nor I_4311 (I76006,I112163,I112139);
nand I_4312 (I75686,I75822,I76006);
nand I_4313 (I75680,I75771,I112163);
nand I_4314 (I76051,I75873,I112157);
DFFARX1 I_4315 (I76051,I2683,I75706,I75695,);
DFFARX1 I_4316 (I76051,I2683,I75706,I75689,);
not I_4317 (I76096,I112157);
nor I_4318 (I76113,I76096,I112145);
and I_4319 (I76130,I76113,I112166);
or I_4320 (I76147,I76130,I112142);
DFFARX1 I_4321 (I76147,I2683,I75706,I76173,);
nand I_4322 (I76181,I76173,I75839);
nor I_4323 (I75683,I76181,I75989);
nor I_4324 (I75677,I76173,I75805);
DFFARX1 I_4325 (I76173,I2683,I75706,I76235,);
not I_4326 (I76243,I76235);
nor I_4327 (I75692,I76243,I75955);
not I_4328 (I76301,I2690);
DFFARX1 I_4329 (I253976,I2683,I76301,I76327,);
DFFARX1 I_4330 (I76327,I2683,I76301,I76344,);
not I_4331 (I76293,I76344);
not I_4332 (I76366,I76327);
DFFARX1 I_4333 (I253970,I2683,I76301,I76392,);
not I_4334 (I76400,I76392);
and I_4335 (I76417,I76366,I253988);
not I_4336 (I76434,I253976);
nand I_4337 (I76451,I76434,I253988);
not I_4338 (I76468,I253970);
nor I_4339 (I76485,I76468,I253982);
nand I_4340 (I76502,I76485,I253973);
nor I_4341 (I76519,I76502,I76451);
DFFARX1 I_4342 (I76519,I2683,I76301,I76269,);
not I_4343 (I76550,I76502);
not I_4344 (I76567,I253982);
nand I_4345 (I76584,I76567,I253988);
nor I_4346 (I76601,I253982,I253976);
nand I_4347 (I76281,I76417,I76601);
nand I_4348 (I76275,I76366,I253982);
nand I_4349 (I76646,I76468,I253985);
DFFARX1 I_4350 (I76646,I2683,I76301,I76290,);
DFFARX1 I_4351 (I76646,I2683,I76301,I76284,);
not I_4352 (I76691,I253985);
nor I_4353 (I76708,I76691,I253991);
and I_4354 (I76725,I76708,I253973);
or I_4355 (I76742,I76725,I253979);
DFFARX1 I_4356 (I76742,I2683,I76301,I76768,);
nand I_4357 (I76776,I76768,I76434);
nor I_4358 (I76278,I76776,I76584);
nor I_4359 (I76272,I76768,I76400);
DFFARX1 I_4360 (I76768,I2683,I76301,I76830,);
not I_4361 (I76838,I76830);
nor I_4362 (I76287,I76838,I76550);
not I_4363 (I76896,I2690);
DFFARX1 I_4364 (I173014,I2683,I76896,I76922,);
DFFARX1 I_4365 (I76922,I2683,I76896,I76939,);
not I_4366 (I76888,I76939);
not I_4367 (I76961,I76922);
DFFARX1 I_4368 (I173005,I2683,I76896,I76987,);
not I_4369 (I76995,I76987);
and I_4370 (I77012,I76961,I173023);
not I_4371 (I77029,I173020);
nand I_4372 (I77046,I77029,I173023);
not I_4373 (I77063,I172999);
nor I_4374 (I77080,I77063,I173002);
nand I_4375 (I77097,I77080,I173011);
nor I_4376 (I77114,I77097,I77046);
DFFARX1 I_4377 (I77114,I2683,I76896,I76864,);
not I_4378 (I77145,I77097);
not I_4379 (I77162,I173002);
nand I_4380 (I77179,I77162,I173023);
nor I_4381 (I77196,I173002,I173020);
nand I_4382 (I76876,I77012,I77196);
nand I_4383 (I76870,I76961,I173002);
nand I_4384 (I77241,I77063,I173017);
DFFARX1 I_4385 (I77241,I2683,I76896,I76885,);
DFFARX1 I_4386 (I77241,I2683,I76896,I76879,);
not I_4387 (I77286,I173017);
nor I_4388 (I77303,I77286,I172999);
and I_4389 (I77320,I77303,I173008);
or I_4390 (I77337,I77320,I173002);
DFFARX1 I_4391 (I77337,I2683,I76896,I77363,);
nand I_4392 (I77371,I77363,I77029);
nor I_4393 (I76873,I77371,I77179);
nor I_4394 (I76867,I77363,I76995);
DFFARX1 I_4395 (I77363,I2683,I76896,I77425,);
not I_4396 (I77433,I77425);
nor I_4397 (I76882,I77433,I77145);
not I_4398 (I77491,I2690);
DFFARX1 I_4399 (I115301,I2683,I77491,I77517,);
DFFARX1 I_4400 (I77517,I2683,I77491,I77534,);
not I_4401 (I77483,I77534);
not I_4402 (I77556,I77517);
DFFARX1 I_4403 (I115316,I2683,I77491,I77582,);
not I_4404 (I77590,I77582);
and I_4405 (I77607,I77556,I115313);
not I_4406 (I77624,I115301);
nand I_4407 (I77641,I77624,I115313);
not I_4408 (I77658,I115310);
nor I_4409 (I77675,I77658,I115325);
nand I_4410 (I77692,I77675,I115322);
nor I_4411 (I77709,I77692,I77641);
DFFARX1 I_4412 (I77709,I2683,I77491,I77459,);
not I_4413 (I77740,I77692);
not I_4414 (I77757,I115325);
nand I_4415 (I77774,I77757,I115313);
nor I_4416 (I77791,I115325,I115301);
nand I_4417 (I77471,I77607,I77791);
nand I_4418 (I77465,I77556,I115325);
nand I_4419 (I77836,I77658,I115319);
DFFARX1 I_4420 (I77836,I2683,I77491,I77480,);
DFFARX1 I_4421 (I77836,I2683,I77491,I77474,);
not I_4422 (I77881,I115319);
nor I_4423 (I77898,I77881,I115307);
and I_4424 (I77915,I77898,I115328);
or I_4425 (I77932,I77915,I115304);
DFFARX1 I_4426 (I77932,I2683,I77491,I77958,);
nand I_4427 (I77966,I77958,I77624);
nor I_4428 (I77468,I77966,I77774);
nor I_4429 (I77462,I77958,I77590);
DFFARX1 I_4430 (I77958,I2683,I77491,I78020,);
not I_4431 (I78028,I78020);
nor I_4432 (I77477,I78028,I77740);
not I_4433 (I78086,I2690);
DFFARX1 I_4434 (I298219,I2683,I78086,I78112,);
DFFARX1 I_4435 (I78112,I2683,I78086,I78129,);
not I_4436 (I78078,I78129);
not I_4437 (I78151,I78112);
DFFARX1 I_4438 (I298228,I2683,I78086,I78177,);
not I_4439 (I78185,I78177);
and I_4440 (I78202,I78151,I298216);
not I_4441 (I78219,I298207);
nand I_4442 (I78236,I78219,I298216);
not I_4443 (I78253,I298213);
nor I_4444 (I78270,I78253,I298231);
nand I_4445 (I78287,I78270,I298204);
nor I_4446 (I78304,I78287,I78236);
DFFARX1 I_4447 (I78304,I2683,I78086,I78054,);
not I_4448 (I78335,I78287);
not I_4449 (I78352,I298231);
nand I_4450 (I78369,I78352,I298216);
nor I_4451 (I78386,I298231,I298207);
nand I_4452 (I78066,I78202,I78386);
nand I_4453 (I78060,I78151,I298231);
nand I_4454 (I78431,I78253,I298210);
DFFARX1 I_4455 (I78431,I2683,I78086,I78075,);
DFFARX1 I_4456 (I78431,I2683,I78086,I78069,);
not I_4457 (I78476,I298210);
nor I_4458 (I78493,I78476,I298222);
and I_4459 (I78510,I78493,I298204);
or I_4460 (I78527,I78510,I298225);
DFFARX1 I_4461 (I78527,I2683,I78086,I78553,);
nand I_4462 (I78561,I78553,I78219);
nor I_4463 (I78063,I78561,I78369);
nor I_4464 (I78057,I78553,I78185);
DFFARX1 I_4465 (I78553,I2683,I78086,I78615,);
not I_4466 (I78623,I78615);
nor I_4467 (I78072,I78623,I78335);
not I_4468 (I78681,I2690);
DFFARX1 I_4469 (I292405,I2683,I78681,I78707,);
DFFARX1 I_4470 (I78707,I2683,I78681,I78724,);
not I_4471 (I78673,I78724);
not I_4472 (I78746,I78707);
DFFARX1 I_4473 (I292414,I2683,I78681,I78772,);
not I_4474 (I78780,I78772);
and I_4475 (I78797,I78746,I292402);
not I_4476 (I78814,I292393);
nand I_4477 (I78831,I78814,I292402);
not I_4478 (I78848,I292399);
nor I_4479 (I78865,I78848,I292417);
nand I_4480 (I78882,I78865,I292390);
nor I_4481 (I78899,I78882,I78831);
DFFARX1 I_4482 (I78899,I2683,I78681,I78649,);
not I_4483 (I78930,I78882);
not I_4484 (I78947,I292417);
nand I_4485 (I78964,I78947,I292402);
nor I_4486 (I78981,I292417,I292393);
nand I_4487 (I78661,I78797,I78981);
nand I_4488 (I78655,I78746,I292417);
nand I_4489 (I79026,I78848,I292396);
DFFARX1 I_4490 (I79026,I2683,I78681,I78670,);
DFFARX1 I_4491 (I79026,I2683,I78681,I78664,);
not I_4492 (I79071,I292396);
nor I_4493 (I79088,I79071,I292408);
and I_4494 (I79105,I79088,I292390);
or I_4495 (I79122,I79105,I292411);
DFFARX1 I_4496 (I79122,I2683,I78681,I79148,);
nand I_4497 (I79156,I79148,I78814);
nor I_4498 (I78658,I79156,I78964);
nor I_4499 (I78652,I79148,I78780);
DFFARX1 I_4500 (I79148,I2683,I78681,I79210,);
not I_4501 (I79218,I79210);
nor I_4502 (I78667,I79218,I78930);
not I_4503 (I79276,I2690);
DFFARX1 I_4504 (I261881,I2683,I79276,I79302,);
DFFARX1 I_4505 (I79302,I2683,I79276,I79319,);
not I_4506 (I79268,I79319);
not I_4507 (I79341,I79302);
DFFARX1 I_4508 (I261875,I2683,I79276,I79367,);
not I_4509 (I79375,I79367);
and I_4510 (I79392,I79341,I261893);
not I_4511 (I79409,I261881);
nand I_4512 (I79426,I79409,I261893);
not I_4513 (I79443,I261875);
nor I_4514 (I79460,I79443,I261887);
nand I_4515 (I79477,I79460,I261878);
nor I_4516 (I79494,I79477,I79426);
DFFARX1 I_4517 (I79494,I2683,I79276,I79244,);
not I_4518 (I79525,I79477);
not I_4519 (I79542,I261887);
nand I_4520 (I79559,I79542,I261893);
nor I_4521 (I79576,I261887,I261881);
nand I_4522 (I79256,I79392,I79576);
nand I_4523 (I79250,I79341,I261887);
nand I_4524 (I79621,I79443,I261890);
DFFARX1 I_4525 (I79621,I2683,I79276,I79265,);
DFFARX1 I_4526 (I79621,I2683,I79276,I79259,);
not I_4527 (I79666,I261890);
nor I_4528 (I79683,I79666,I261896);
and I_4529 (I79700,I79683,I261878);
or I_4530 (I79717,I79700,I261884);
DFFARX1 I_4531 (I79717,I2683,I79276,I79743,);
nand I_4532 (I79751,I79743,I79409);
nor I_4533 (I79253,I79751,I79559);
nor I_4534 (I79247,I79743,I79375);
DFFARX1 I_4535 (I79743,I2683,I79276,I79805,);
not I_4536 (I79813,I79805);
nor I_4537 (I79262,I79813,I79525);
not I_4538 (I79871,I2690);
DFFARX1 I_4539 (I40986,I2683,I79871,I79897,);
DFFARX1 I_4540 (I79897,I2683,I79871,I79914,);
not I_4541 (I79863,I79914);
not I_4542 (I79936,I79897);
DFFARX1 I_4543 (I40980,I2683,I79871,I79962,);
not I_4544 (I79970,I79962);
and I_4545 (I79987,I79936,I40977);
not I_4546 (I80004,I40998);
nand I_4547 (I80021,I80004,I40977);
not I_4548 (I80038,I40992);
nor I_4549 (I80055,I80038,I40983);
nand I_4550 (I80072,I80055,I40989);
nor I_4551 (I80089,I80072,I80021);
DFFARX1 I_4552 (I80089,I2683,I79871,I79839,);
not I_4553 (I80120,I80072);
not I_4554 (I80137,I40983);
nand I_4555 (I80154,I80137,I40977);
nor I_4556 (I80171,I40983,I40998);
nand I_4557 (I79851,I79987,I80171);
nand I_4558 (I79845,I79936,I40983);
nand I_4559 (I80216,I80038,I40977);
DFFARX1 I_4560 (I80216,I2683,I79871,I79860,);
DFFARX1 I_4561 (I80216,I2683,I79871,I79854,);
not I_4562 (I80261,I40977);
nor I_4563 (I80278,I80261,I40995);
and I_4564 (I80295,I80278,I41001);
or I_4565 (I80312,I80295,I40980);
DFFARX1 I_4566 (I80312,I2683,I79871,I80338,);
nand I_4567 (I80346,I80338,I80004);
nor I_4568 (I79848,I80346,I80154);
nor I_4569 (I79842,I80338,I79970);
DFFARX1 I_4570 (I80338,I2683,I79871,I80400,);
not I_4571 (I80408,I80400);
nor I_4572 (I79857,I80408,I80120);
not I_4573 (I80466,I2690);
DFFARX1 I_4574 (I400990,I2683,I80466,I80492,);
DFFARX1 I_4575 (I80492,I2683,I80466,I80509,);
not I_4576 (I80458,I80509);
not I_4577 (I80531,I80492);
DFFARX1 I_4578 (I400981,I2683,I80466,I80557,);
not I_4579 (I80565,I80557);
and I_4580 (I80582,I80531,I400975);
not I_4581 (I80599,I400969);
nand I_4582 (I80616,I80599,I400975);
not I_4583 (I80633,I400996);
nor I_4584 (I80650,I80633,I400969);
nand I_4585 (I80667,I80650,I400993);
nor I_4586 (I80684,I80667,I80616);
DFFARX1 I_4587 (I80684,I2683,I80466,I80434,);
not I_4588 (I80715,I80667);
not I_4589 (I80732,I400969);
nand I_4590 (I80749,I80732,I400975);
nor I_4591 (I80766,I400969,I400969);
nand I_4592 (I80446,I80582,I80766);
nand I_4593 (I80440,I80531,I400969);
nand I_4594 (I80811,I80633,I400978);
DFFARX1 I_4595 (I80811,I2683,I80466,I80455,);
DFFARX1 I_4596 (I80811,I2683,I80466,I80449,);
not I_4597 (I80856,I400978);
nor I_4598 (I80873,I80856,I400984);
and I_4599 (I80890,I80873,I400987);
or I_4600 (I80907,I80890,I400972);
DFFARX1 I_4601 (I80907,I2683,I80466,I80933,);
nand I_4602 (I80941,I80933,I80599);
nor I_4603 (I80443,I80941,I80749);
nor I_4604 (I80437,I80933,I80565);
DFFARX1 I_4605 (I80933,I2683,I80466,I80995,);
not I_4606 (I81003,I80995);
nor I_4607 (I80452,I81003,I80715);
not I_4608 (I81061,I2690);
DFFARX1 I_4609 (I30973,I2683,I81061,I81087,);
DFFARX1 I_4610 (I81087,I2683,I81061,I81104,);
not I_4611 (I81053,I81104);
not I_4612 (I81126,I81087);
DFFARX1 I_4613 (I30967,I2683,I81061,I81152,);
not I_4614 (I81160,I81152);
and I_4615 (I81177,I81126,I30964);
not I_4616 (I81194,I30985);
nand I_4617 (I81211,I81194,I30964);
not I_4618 (I81228,I30979);
nor I_4619 (I81245,I81228,I30970);
nand I_4620 (I81262,I81245,I30976);
nor I_4621 (I81279,I81262,I81211);
DFFARX1 I_4622 (I81279,I2683,I81061,I81029,);
not I_4623 (I81310,I81262);
not I_4624 (I81327,I30970);
nand I_4625 (I81344,I81327,I30964);
nor I_4626 (I81361,I30970,I30985);
nand I_4627 (I81041,I81177,I81361);
nand I_4628 (I81035,I81126,I30970);
nand I_4629 (I81406,I81228,I30964);
DFFARX1 I_4630 (I81406,I2683,I81061,I81050,);
DFFARX1 I_4631 (I81406,I2683,I81061,I81044,);
not I_4632 (I81451,I30964);
nor I_4633 (I81468,I81451,I30982);
and I_4634 (I81485,I81468,I30988);
or I_4635 (I81502,I81485,I30967);
DFFARX1 I_4636 (I81502,I2683,I81061,I81528,);
nand I_4637 (I81536,I81528,I81194);
nor I_4638 (I81038,I81536,I81344);
nor I_4639 (I81032,I81528,I81160);
DFFARX1 I_4640 (I81528,I2683,I81061,I81590,);
not I_4641 (I81598,I81590);
nor I_4642 (I81047,I81598,I81310);
not I_4643 (I81656,I2690);
DFFARX1 I_4644 (I164766,I2683,I81656,I81682,);
DFFARX1 I_4645 (I81682,I2683,I81656,I81699,);
not I_4646 (I81648,I81699);
not I_4647 (I81721,I81682);
DFFARX1 I_4648 (I164760,I2683,I81656,I81747,);
not I_4649 (I81755,I81747);
and I_4650 (I81772,I81721,I164775);
not I_4651 (I81789,I164772);
nand I_4652 (I81806,I81789,I164775);
not I_4653 (I81823,I164763);
nor I_4654 (I81840,I81823,I164754);
nand I_4655 (I81857,I81840,I164757);
nor I_4656 (I81874,I81857,I81806);
DFFARX1 I_4657 (I81874,I2683,I81656,I81624,);
not I_4658 (I81905,I81857);
not I_4659 (I81922,I164754);
nand I_4660 (I81939,I81922,I164775);
nor I_4661 (I81956,I164754,I164772);
nand I_4662 (I81636,I81772,I81956);
nand I_4663 (I81630,I81721,I164754);
nand I_4664 (I82001,I81823,I164778);
DFFARX1 I_4665 (I82001,I2683,I81656,I81645,);
DFFARX1 I_4666 (I82001,I2683,I81656,I81639,);
not I_4667 (I82046,I164778);
nor I_4668 (I82063,I82046,I164769);
and I_4669 (I82080,I82063,I164754);
or I_4670 (I82097,I82080,I164757);
DFFARX1 I_4671 (I82097,I2683,I81656,I82123,);
nand I_4672 (I82131,I82123,I81789);
nor I_4673 (I81633,I82131,I81939);
nor I_4674 (I81627,I82123,I81755);
DFFARX1 I_4675 (I82123,I2683,I81656,I82185,);
not I_4676 (I82193,I82185);
nor I_4677 (I81642,I82193,I81905);
not I_4678 (I82251,I2690);
DFFARX1 I_4679 (I182262,I2683,I82251,I82277,);
DFFARX1 I_4680 (I82277,I2683,I82251,I82294,);
not I_4681 (I82243,I82294);
not I_4682 (I82316,I82277);
DFFARX1 I_4683 (I182253,I2683,I82251,I82342,);
not I_4684 (I82350,I82342);
and I_4685 (I82367,I82316,I182271);
not I_4686 (I82384,I182268);
nand I_4687 (I82401,I82384,I182271);
not I_4688 (I82418,I182247);
nor I_4689 (I82435,I82418,I182250);
nand I_4690 (I82452,I82435,I182259);
nor I_4691 (I82469,I82452,I82401);
DFFARX1 I_4692 (I82469,I2683,I82251,I82219,);
not I_4693 (I82500,I82452);
not I_4694 (I82517,I182250);
nand I_4695 (I82534,I82517,I182271);
nor I_4696 (I82551,I182250,I182268);
nand I_4697 (I82231,I82367,I82551);
nand I_4698 (I82225,I82316,I182250);
nand I_4699 (I82596,I82418,I182265);
DFFARX1 I_4700 (I82596,I2683,I82251,I82240,);
DFFARX1 I_4701 (I82596,I2683,I82251,I82234,);
not I_4702 (I82641,I182265);
nor I_4703 (I82658,I82641,I182247);
and I_4704 (I82675,I82658,I182256);
or I_4705 (I82692,I82675,I182250);
DFFARX1 I_4706 (I82692,I2683,I82251,I82718,);
nand I_4707 (I82726,I82718,I82384);
nor I_4708 (I82228,I82726,I82534);
nor I_4709 (I82222,I82718,I82350);
DFFARX1 I_4710 (I82718,I2683,I82251,I82780,);
not I_4711 (I82788,I82780);
nor I_4712 (I82237,I82788,I82500);
not I_4713 (I82846,I2690);
DFFARX1 I_4714 (I91586,I2683,I82846,I82872,);
DFFARX1 I_4715 (I82872,I2683,I82846,I82889,);
not I_4716 (I82838,I82889);
not I_4717 (I82911,I82872);
DFFARX1 I_4718 (I91601,I2683,I82846,I82937,);
not I_4719 (I82945,I82937);
and I_4720 (I82962,I82911,I91598);
not I_4721 (I82979,I91586);
nand I_4722 (I82996,I82979,I91598);
not I_4723 (I83013,I91595);
nor I_4724 (I83030,I83013,I91610);
nand I_4725 (I83047,I83030,I91607);
nor I_4726 (I83064,I83047,I82996);
DFFARX1 I_4727 (I83064,I2683,I82846,I82814,);
not I_4728 (I83095,I83047);
not I_4729 (I83112,I91610);
nand I_4730 (I83129,I83112,I91598);
nor I_4731 (I83146,I91610,I91586);
nand I_4732 (I82826,I82962,I83146);
nand I_4733 (I82820,I82911,I91610);
nand I_4734 (I83191,I83013,I91604);
DFFARX1 I_4735 (I83191,I2683,I82846,I82835,);
DFFARX1 I_4736 (I83191,I2683,I82846,I82829,);
not I_4737 (I83236,I91604);
nor I_4738 (I83253,I83236,I91592);
and I_4739 (I83270,I83253,I91613);
or I_4740 (I83287,I83270,I91589);
DFFARX1 I_4741 (I83287,I2683,I82846,I83313,);
nand I_4742 (I83321,I83313,I82979);
nor I_4743 (I82823,I83321,I83129);
nor I_4744 (I82817,I83313,I82945);
DFFARX1 I_4745 (I83313,I2683,I82846,I83375,);
not I_4746 (I83383,I83375);
nor I_4747 (I82832,I83383,I83095);
not I_4748 (I83441,I2690);
DFFARX1 I_4749 (I300157,I2683,I83441,I83467,);
DFFARX1 I_4750 (I83467,I2683,I83441,I83484,);
not I_4751 (I83433,I83484);
not I_4752 (I83506,I83467);
DFFARX1 I_4753 (I300166,I2683,I83441,I83532,);
not I_4754 (I83540,I83532);
and I_4755 (I83557,I83506,I300154);
not I_4756 (I83574,I300145);
nand I_4757 (I83591,I83574,I300154);
not I_4758 (I83608,I300151);
nor I_4759 (I83625,I83608,I300169);
nand I_4760 (I83642,I83625,I300142);
nor I_4761 (I83659,I83642,I83591);
DFFARX1 I_4762 (I83659,I2683,I83441,I83409,);
not I_4763 (I83690,I83642);
not I_4764 (I83707,I300169);
nand I_4765 (I83724,I83707,I300154);
nor I_4766 (I83741,I300169,I300145);
nand I_4767 (I83421,I83557,I83741);
nand I_4768 (I83415,I83506,I300169);
nand I_4769 (I83786,I83608,I300148);
DFFARX1 I_4770 (I83786,I2683,I83441,I83430,);
DFFARX1 I_4771 (I83786,I2683,I83441,I83424,);
not I_4772 (I83831,I300148);
nor I_4773 (I83848,I83831,I300160);
and I_4774 (I83865,I83848,I300142);
or I_4775 (I83882,I83865,I300163);
DFFARX1 I_4776 (I83882,I2683,I83441,I83908,);
nand I_4777 (I83916,I83908,I83574);
nor I_4778 (I83418,I83916,I83724);
nor I_4779 (I83412,I83908,I83540);
DFFARX1 I_4780 (I83908,I2683,I83441,I83970,);
not I_4781 (I83978,I83970);
nor I_4782 (I83427,I83978,I83690);
not I_4783 (I84036,I2690);
DFFARX1 I_4784 (I409915,I2683,I84036,I84062,);
DFFARX1 I_4785 (I84062,I2683,I84036,I84079,);
not I_4786 (I84028,I84079);
not I_4787 (I84101,I84062);
DFFARX1 I_4788 (I409906,I2683,I84036,I84127,);
not I_4789 (I84135,I84127);
and I_4790 (I84152,I84101,I409900);
not I_4791 (I84169,I409894);
nand I_4792 (I84186,I84169,I409900);
not I_4793 (I84203,I409921);
nor I_4794 (I84220,I84203,I409894);
nand I_4795 (I84237,I84220,I409918);
nor I_4796 (I84254,I84237,I84186);
DFFARX1 I_4797 (I84254,I2683,I84036,I84004,);
not I_4798 (I84285,I84237);
not I_4799 (I84302,I409894);
nand I_4800 (I84319,I84302,I409900);
nor I_4801 (I84336,I409894,I409894);
nand I_4802 (I84016,I84152,I84336);
nand I_4803 (I84010,I84101,I409894);
nand I_4804 (I84381,I84203,I409903);
DFFARX1 I_4805 (I84381,I2683,I84036,I84025,);
DFFARX1 I_4806 (I84381,I2683,I84036,I84019,);
not I_4807 (I84426,I409903);
nor I_4808 (I84443,I84426,I409909);
and I_4809 (I84460,I84443,I409912);
or I_4810 (I84477,I84460,I409897);
DFFARX1 I_4811 (I84477,I2683,I84036,I84503,);
nand I_4812 (I84511,I84503,I84169);
nor I_4813 (I84013,I84511,I84319);
nor I_4814 (I84007,I84503,I84135);
DFFARX1 I_4815 (I84503,I2683,I84036,I84565,);
not I_4816 (I84573,I84565);
nor I_4817 (I84022,I84573,I84285);
not I_4818 (I84631,I2690);
DFFARX1 I_4819 (I406940,I2683,I84631,I84657,);
DFFARX1 I_4820 (I84657,I2683,I84631,I84674,);
not I_4821 (I84623,I84674);
not I_4822 (I84696,I84657);
DFFARX1 I_4823 (I406931,I2683,I84631,I84722,);
not I_4824 (I84730,I84722);
and I_4825 (I84747,I84696,I406925);
not I_4826 (I84764,I406919);
nand I_4827 (I84781,I84764,I406925);
not I_4828 (I84798,I406946);
nor I_4829 (I84815,I84798,I406919);
nand I_4830 (I84832,I84815,I406943);
nor I_4831 (I84849,I84832,I84781);
DFFARX1 I_4832 (I84849,I2683,I84631,I84599,);
not I_4833 (I84880,I84832);
not I_4834 (I84897,I406919);
nand I_4835 (I84914,I84897,I406925);
nor I_4836 (I84931,I406919,I406919);
nand I_4837 (I84611,I84747,I84931);
nand I_4838 (I84605,I84696,I406919);
nand I_4839 (I84976,I84798,I406928);
DFFARX1 I_4840 (I84976,I2683,I84631,I84620,);
DFFARX1 I_4841 (I84976,I2683,I84631,I84614,);
not I_4842 (I85021,I406928);
nor I_4843 (I85038,I85021,I406934);
and I_4844 (I85055,I85038,I406937);
or I_4845 (I85072,I85055,I406922);
DFFARX1 I_4846 (I85072,I2683,I84631,I85098,);
nand I_4847 (I85106,I85098,I84764);
nor I_4848 (I84608,I85106,I84914);
nor I_4849 (I84602,I85098,I84730);
DFFARX1 I_4850 (I85098,I2683,I84631,I85160,);
not I_4851 (I85168,I85160);
nor I_4852 (I84617,I85168,I84880);
not I_4853 (I85226,I2690);
DFFARX1 I_4854 (I5692,I2683,I85226,I85252,);
DFFARX1 I_4855 (I85252,I2683,I85226,I85269,);
not I_4856 (I85218,I85269);
not I_4857 (I85291,I85252);
DFFARX1 I_4858 (I5668,I2683,I85226,I85317,);
not I_4859 (I85325,I85317);
and I_4860 (I85342,I85291,I5683);
not I_4861 (I85359,I5671);
nand I_4862 (I85376,I85359,I5683);
not I_4863 (I85393,I5674);
nor I_4864 (I85410,I85393,I5686);
nand I_4865 (I85427,I85410,I5677);
nor I_4866 (I85444,I85427,I85376);
DFFARX1 I_4867 (I85444,I2683,I85226,I85194,);
not I_4868 (I85475,I85427);
not I_4869 (I85492,I5686);
nand I_4870 (I85509,I85492,I5683);
nor I_4871 (I85526,I5686,I5671);
nand I_4872 (I85206,I85342,I85526);
nand I_4873 (I85200,I85291,I5686);
nand I_4874 (I85571,I85393,I5680);
DFFARX1 I_4875 (I85571,I2683,I85226,I85215,);
DFFARX1 I_4876 (I85571,I2683,I85226,I85209,);
not I_4877 (I85616,I5680);
nor I_4878 (I85633,I85616,I5671);
and I_4879 (I85650,I85633,I5668);
or I_4880 (I85667,I85650,I5689);
DFFARX1 I_4881 (I85667,I2683,I85226,I85693,);
nand I_4882 (I85701,I85693,I85359);
nor I_4883 (I85203,I85701,I85509);
nor I_4884 (I85197,I85693,I85325);
DFFARX1 I_4885 (I85693,I2683,I85226,I85755,);
not I_4886 (I85763,I85755);
nor I_4887 (I85212,I85763,I85475);
not I_4888 (I85824,I2690);
DFFARX1 I_4889 (I237109,I2683,I85824,I85850,);
nand I_4890 (I85858,I237112,I237106);
and I_4891 (I85875,I85858,I237118);
DFFARX1 I_4892 (I85875,I2683,I85824,I85901,);
nor I_4893 (I85792,I85901,I85850);
not I_4894 (I85923,I85901);
DFFARX1 I_4895 (I237121,I2683,I85824,I85949,);
nand I_4896 (I85957,I85949,I237112);
not I_4897 (I85974,I85957);
DFFARX1 I_4898 (I85974,I2683,I85824,I86000,);
not I_4899 (I85816,I86000);
nor I_4900 (I86022,I85850,I85957);
nor I_4901 (I85798,I85901,I86022);
DFFARX1 I_4902 (I237124,I2683,I85824,I86062,);
DFFARX1 I_4903 (I86062,I2683,I85824,I86079,);
not I_4904 (I86087,I86079);
not I_4905 (I86104,I86062);
nand I_4906 (I85801,I86104,I85923);
nand I_4907 (I86135,I237106,I237115);
and I_4908 (I86152,I86135,I237109);
DFFARX1 I_4909 (I86152,I2683,I85824,I86178,);
nor I_4910 (I86186,I86178,I85850);
DFFARX1 I_4911 (I86186,I2683,I85824,I85789,);
DFFARX1 I_4912 (I86178,I2683,I85824,I85807,);
nor I_4913 (I86231,I237127,I237115);
not I_4914 (I86248,I86231);
nor I_4915 (I85810,I86087,I86248);
nand I_4916 (I85795,I86104,I86248);
nor I_4917 (I85804,I85850,I86231);
DFFARX1 I_4918 (I86231,I2683,I85824,I85813,);
not I_4919 (I86351,I2690);
DFFARX1 I_4920 (I390002,I2683,I86351,I86377,);
nand I_4921 (I86385,I389999,I389990);
and I_4922 (I86402,I86385,I389987);
DFFARX1 I_4923 (I86402,I2683,I86351,I86428,);
nor I_4924 (I86319,I86428,I86377);
not I_4925 (I86450,I86428);
DFFARX1 I_4926 (I389996,I2683,I86351,I86476,);
nand I_4927 (I86484,I86476,I390005);
not I_4928 (I86501,I86484);
DFFARX1 I_4929 (I86501,I2683,I86351,I86527,);
not I_4930 (I86343,I86527);
nor I_4931 (I86549,I86377,I86484);
nor I_4932 (I86325,I86428,I86549);
DFFARX1 I_4933 (I390008,I2683,I86351,I86589,);
DFFARX1 I_4934 (I86589,I2683,I86351,I86606,);
not I_4935 (I86614,I86606);
not I_4936 (I86631,I86589);
nand I_4937 (I86328,I86631,I86450);
nand I_4938 (I86662,I389987,I389993);
and I_4939 (I86679,I86662,I390011);
DFFARX1 I_4940 (I86679,I2683,I86351,I86705,);
nor I_4941 (I86713,I86705,I86377);
DFFARX1 I_4942 (I86713,I2683,I86351,I86316,);
DFFARX1 I_4943 (I86705,I2683,I86351,I86334,);
nor I_4944 (I86758,I389990,I389993);
not I_4945 (I86775,I86758);
nor I_4946 (I86337,I86614,I86775);
nand I_4947 (I86322,I86631,I86775);
nor I_4948 (I86331,I86377,I86758);
DFFARX1 I_4949 (I86758,I2683,I86351,I86340,);
not I_4950 (I86878,I2690);
DFFARX1 I_4951 (I385378,I2683,I86878,I86904,);
nand I_4952 (I86912,I385375,I385366);
and I_4953 (I86929,I86912,I385363);
DFFARX1 I_4954 (I86929,I2683,I86878,I86955,);
nor I_4955 (I86846,I86955,I86904);
not I_4956 (I86977,I86955);
DFFARX1 I_4957 (I385372,I2683,I86878,I87003,);
nand I_4958 (I87011,I87003,I385381);
not I_4959 (I87028,I87011);
DFFARX1 I_4960 (I87028,I2683,I86878,I87054,);
not I_4961 (I86870,I87054);
nor I_4962 (I87076,I86904,I87011);
nor I_4963 (I86852,I86955,I87076);
DFFARX1 I_4964 (I385384,I2683,I86878,I87116,);
DFFARX1 I_4965 (I87116,I2683,I86878,I87133,);
not I_4966 (I87141,I87133);
not I_4967 (I87158,I87116);
nand I_4968 (I86855,I87158,I86977);
nand I_4969 (I87189,I385363,I385369);
and I_4970 (I87206,I87189,I385387);
DFFARX1 I_4971 (I87206,I2683,I86878,I87232,);
nor I_4972 (I87240,I87232,I86904);
DFFARX1 I_4973 (I87240,I2683,I86878,I86843,);
DFFARX1 I_4974 (I87232,I2683,I86878,I86861,);
nor I_4975 (I87285,I385366,I385369);
not I_4976 (I87302,I87285);
nor I_4977 (I86864,I87141,I87302);
nand I_4978 (I86849,I87158,I87302);
nor I_4979 (I86858,I86904,I87285);
DFFARX1 I_4980 (I87285,I2683,I86878,I86867,);
not I_4981 (I87405,I2690);
DFFARX1 I_4982 (I207113,I2683,I87405,I87431,);
nand I_4983 (I87439,I207104,I207119);
and I_4984 (I87456,I87439,I207125);
DFFARX1 I_4985 (I87456,I2683,I87405,I87482,);
nor I_4986 (I87373,I87482,I87431);
not I_4987 (I87504,I87482);
DFFARX1 I_4988 (I207110,I2683,I87405,I87530,);
nand I_4989 (I87538,I87530,I207104);
not I_4990 (I87555,I87538);
DFFARX1 I_4991 (I87555,I2683,I87405,I87581,);
not I_4992 (I87397,I87581);
nor I_4993 (I87603,I87431,I87538);
nor I_4994 (I87379,I87482,I87603);
DFFARX1 I_4995 (I207107,I2683,I87405,I87643,);
DFFARX1 I_4996 (I87643,I2683,I87405,I87660,);
not I_4997 (I87668,I87660);
not I_4998 (I87685,I87643);
nand I_4999 (I87382,I87685,I87504);
nand I_5000 (I87716,I207101,I207116);
and I_5001 (I87733,I87716,I207101);
DFFARX1 I_5002 (I87733,I2683,I87405,I87759,);
nor I_5003 (I87767,I87759,I87431);
DFFARX1 I_5004 (I87767,I2683,I87405,I87370,);
DFFARX1 I_5005 (I87759,I2683,I87405,I87388,);
nor I_5006 (I87812,I207122,I207116);
not I_5007 (I87829,I87812);
nor I_5008 (I87391,I87668,I87829);
nand I_5009 (I87376,I87685,I87829);
nor I_5010 (I87385,I87431,I87812);
DFFARX1 I_5011 (I87812,I2683,I87405,I87394,);
not I_5012 (I87932,I2690);
DFFARX1 I_5013 (I384222,I2683,I87932,I87958,);
nand I_5014 (I87966,I384219,I384210);
and I_5015 (I87983,I87966,I384207);
DFFARX1 I_5016 (I87983,I2683,I87932,I88009,);
nor I_5017 (I87900,I88009,I87958);
not I_5018 (I88031,I88009);
DFFARX1 I_5019 (I384216,I2683,I87932,I88057,);
nand I_5020 (I88065,I88057,I384225);
not I_5021 (I88082,I88065);
DFFARX1 I_5022 (I88082,I2683,I87932,I88108,);
not I_5023 (I87924,I88108);
nor I_5024 (I88130,I87958,I88065);
nor I_5025 (I87906,I88009,I88130);
DFFARX1 I_5026 (I384228,I2683,I87932,I88170,);
DFFARX1 I_5027 (I88170,I2683,I87932,I88187,);
not I_5028 (I88195,I88187);
not I_5029 (I88212,I88170);
nand I_5030 (I87909,I88212,I88031);
nand I_5031 (I88243,I384207,I384213);
and I_5032 (I88260,I88243,I384231);
DFFARX1 I_5033 (I88260,I2683,I87932,I88286,);
nor I_5034 (I88294,I88286,I87958);
DFFARX1 I_5035 (I88294,I2683,I87932,I87897,);
DFFARX1 I_5036 (I88286,I2683,I87932,I87915,);
nor I_5037 (I88339,I384210,I384213);
not I_5038 (I88356,I88339);
nor I_5039 (I87918,I88195,I88356);
nand I_5040 (I87903,I88212,I88356);
nor I_5041 (I87912,I87958,I88339);
DFFARX1 I_5042 (I88339,I2683,I87932,I87921,);
not I_5043 (I88459,I2690);
DFFARX1 I_5044 (I399800,I2683,I88459,I88485,);
nand I_5045 (I88493,I399779,I399779);
and I_5046 (I88510,I88493,I399806);
DFFARX1 I_5047 (I88510,I2683,I88459,I88536,);
nor I_5048 (I88427,I88536,I88485);
not I_5049 (I88558,I88536);
DFFARX1 I_5050 (I399794,I2683,I88459,I88584,);
nand I_5051 (I88592,I88584,I399797);
not I_5052 (I88609,I88592);
DFFARX1 I_5053 (I88609,I2683,I88459,I88635,);
not I_5054 (I88451,I88635);
nor I_5055 (I88657,I88485,I88592);
nor I_5056 (I88433,I88536,I88657);
DFFARX1 I_5057 (I399788,I2683,I88459,I88697,);
DFFARX1 I_5058 (I88697,I2683,I88459,I88714,);
not I_5059 (I88722,I88714);
not I_5060 (I88739,I88697);
nand I_5061 (I88436,I88739,I88558);
nand I_5062 (I88770,I399785,I399782);
and I_5063 (I88787,I88770,I399803);
DFFARX1 I_5064 (I88787,I2683,I88459,I88813,);
nor I_5065 (I88821,I88813,I88485);
DFFARX1 I_5066 (I88821,I2683,I88459,I88424,);
DFFARX1 I_5067 (I88813,I2683,I88459,I88442,);
nor I_5068 (I88866,I399791,I399782);
not I_5069 (I88883,I88866);
nor I_5070 (I88445,I88722,I88883);
nand I_5071 (I88430,I88739,I88883);
nor I_5072 (I88439,I88485,I88866);
DFFARX1 I_5073 (I88866,I2683,I88459,I88448,);
not I_5074 (I88986,I2690);
DFFARX1 I_5075 (I407535,I2683,I88986,I89012,);
nand I_5076 (I89020,I407514,I407514);
and I_5077 (I89037,I89020,I407541);
DFFARX1 I_5078 (I89037,I2683,I88986,I89063,);
nor I_5079 (I88954,I89063,I89012);
not I_5080 (I89085,I89063);
DFFARX1 I_5081 (I407529,I2683,I88986,I89111,);
nand I_5082 (I89119,I89111,I407532);
not I_5083 (I89136,I89119);
DFFARX1 I_5084 (I89136,I2683,I88986,I89162,);
not I_5085 (I88978,I89162);
nor I_5086 (I89184,I89012,I89119);
nor I_5087 (I88960,I89063,I89184);
DFFARX1 I_5088 (I407523,I2683,I88986,I89224,);
DFFARX1 I_5089 (I89224,I2683,I88986,I89241,);
not I_5090 (I89249,I89241);
not I_5091 (I89266,I89224);
nand I_5092 (I88963,I89266,I89085);
nand I_5093 (I89297,I407520,I407517);
and I_5094 (I89314,I89297,I407538);
DFFARX1 I_5095 (I89314,I2683,I88986,I89340,);
nor I_5096 (I89348,I89340,I89012);
DFFARX1 I_5097 (I89348,I2683,I88986,I88951,);
DFFARX1 I_5098 (I89340,I2683,I88986,I88969,);
nor I_5099 (I89393,I407526,I407517);
not I_5100 (I89410,I89393);
nor I_5101 (I88972,I89249,I89410);
nand I_5102 (I88957,I89266,I89410);
nor I_5103 (I88966,I89012,I89393);
DFFARX1 I_5104 (I89393,I2683,I88986,I88975,);
not I_5105 (I89513,I2690);
DFFARX1 I_5106 (I141595,I2683,I89513,I89539,);
nand I_5107 (I89547,I141607,I141586);
and I_5108 (I89564,I89547,I141610);
DFFARX1 I_5109 (I89564,I2683,I89513,I89590,);
nor I_5110 (I89481,I89590,I89539);
not I_5111 (I89612,I89590);
DFFARX1 I_5112 (I141601,I2683,I89513,I89638,);
nand I_5113 (I89646,I89638,I141583);
not I_5114 (I89663,I89646);
DFFARX1 I_5115 (I89663,I2683,I89513,I89689,);
not I_5116 (I89505,I89689);
nor I_5117 (I89711,I89539,I89646);
nor I_5118 (I89487,I89590,I89711);
DFFARX1 I_5119 (I141598,I2683,I89513,I89751,);
DFFARX1 I_5120 (I89751,I2683,I89513,I89768,);
not I_5121 (I89776,I89768);
not I_5122 (I89793,I89751);
nand I_5123 (I89490,I89793,I89612);
nand I_5124 (I89824,I141583,I141589);
and I_5125 (I89841,I89824,I141592);
DFFARX1 I_5126 (I89841,I2683,I89513,I89867,);
nor I_5127 (I89875,I89867,I89539);
DFFARX1 I_5128 (I89875,I2683,I89513,I89478,);
DFFARX1 I_5129 (I89867,I2683,I89513,I89496,);
nor I_5130 (I89920,I141604,I141589);
not I_5131 (I89937,I89920);
nor I_5132 (I89499,I89776,I89937);
nand I_5133 (I89484,I89793,I89937);
nor I_5134 (I89493,I89539,I89920);
DFFARX1 I_5135 (I89920,I2683,I89513,I89502,);
not I_5136 (I90040,I2690);
DFFARX1 I_5137 (I408130,I2683,I90040,I90066,);
nand I_5138 (I90074,I408109,I408109);
and I_5139 (I90091,I90074,I408136);
DFFARX1 I_5140 (I90091,I2683,I90040,I90117,);
nor I_5141 (I90008,I90117,I90066);
not I_5142 (I90139,I90117);
DFFARX1 I_5143 (I408124,I2683,I90040,I90165,);
nand I_5144 (I90173,I90165,I408127);
not I_5145 (I90190,I90173);
DFFARX1 I_5146 (I90190,I2683,I90040,I90216,);
not I_5147 (I90032,I90216);
nor I_5148 (I90238,I90066,I90173);
nor I_5149 (I90014,I90117,I90238);
DFFARX1 I_5150 (I408118,I2683,I90040,I90278,);
DFFARX1 I_5151 (I90278,I2683,I90040,I90295,);
not I_5152 (I90303,I90295);
not I_5153 (I90320,I90278);
nand I_5154 (I90017,I90320,I90139);
nand I_5155 (I90351,I408115,I408112);
and I_5156 (I90368,I90351,I408133);
DFFARX1 I_5157 (I90368,I2683,I90040,I90394,);
nor I_5158 (I90402,I90394,I90066);
DFFARX1 I_5159 (I90402,I2683,I90040,I90005,);
DFFARX1 I_5160 (I90394,I2683,I90040,I90023,);
nor I_5161 (I90447,I408121,I408112);
not I_5162 (I90464,I90447);
nor I_5163 (I90026,I90303,I90464);
nand I_5164 (I90011,I90320,I90464);
nor I_5165 (I90020,I90066,I90447);
DFFARX1 I_5166 (I90447,I2683,I90040,I90029,);
not I_5167 (I90567,I2690);
DFFARX1 I_5168 (I392314,I2683,I90567,I90593,);
nand I_5169 (I90601,I392311,I392302);
and I_5170 (I90618,I90601,I392299);
DFFARX1 I_5171 (I90618,I2683,I90567,I90644,);
nor I_5172 (I90535,I90644,I90593);
not I_5173 (I90666,I90644);
DFFARX1 I_5174 (I392308,I2683,I90567,I90692,);
nand I_5175 (I90700,I90692,I392317);
not I_5176 (I90717,I90700);
DFFARX1 I_5177 (I90717,I2683,I90567,I90743,);
not I_5178 (I90559,I90743);
nor I_5179 (I90765,I90593,I90700);
nor I_5180 (I90541,I90644,I90765);
DFFARX1 I_5181 (I392320,I2683,I90567,I90805,);
DFFARX1 I_5182 (I90805,I2683,I90567,I90822,);
not I_5183 (I90830,I90822);
not I_5184 (I90847,I90805);
nand I_5185 (I90544,I90847,I90666);
nand I_5186 (I90878,I392299,I392305);
and I_5187 (I90895,I90878,I392323);
DFFARX1 I_5188 (I90895,I2683,I90567,I90921,);
nor I_5189 (I90929,I90921,I90593);
DFFARX1 I_5190 (I90929,I2683,I90567,I90532,);
DFFARX1 I_5191 (I90921,I2683,I90567,I90550,);
nor I_5192 (I90974,I392302,I392305);
not I_5193 (I90991,I90974);
nor I_5194 (I90553,I90830,I90991);
nand I_5195 (I90538,I90847,I90991);
nor I_5196 (I90547,I90593,I90974);
DFFARX1 I_5197 (I90974,I2683,I90567,I90556,);
not I_5198 (I91094,I2690);
DFFARX1 I_5199 (I56039,I2683,I91094,I91120,);
nand I_5200 (I91128,I56039,I56045);
and I_5201 (I91145,I91128,I56063);
DFFARX1 I_5202 (I91145,I2683,I91094,I91171,);
nor I_5203 (I91062,I91171,I91120);
not I_5204 (I91193,I91171);
DFFARX1 I_5205 (I56051,I2683,I91094,I91219,);
nand I_5206 (I91227,I91219,I56048);
not I_5207 (I91244,I91227);
DFFARX1 I_5208 (I91244,I2683,I91094,I91270,);
not I_5209 (I91086,I91270);
nor I_5210 (I91292,I91120,I91227);
nor I_5211 (I91068,I91171,I91292);
DFFARX1 I_5212 (I56057,I2683,I91094,I91332,);
DFFARX1 I_5213 (I91332,I2683,I91094,I91349,);
not I_5214 (I91357,I91349);
not I_5215 (I91374,I91332);
nand I_5216 (I91071,I91374,I91193);
nand I_5217 (I91405,I56042,I56042);
and I_5218 (I91422,I91405,I56054);
DFFARX1 I_5219 (I91422,I2683,I91094,I91448,);
nor I_5220 (I91456,I91448,I91120);
DFFARX1 I_5221 (I91456,I2683,I91094,I91059,);
DFFARX1 I_5222 (I91448,I2683,I91094,I91077,);
nor I_5223 (I91501,I56060,I56042);
not I_5224 (I91518,I91501);
nor I_5225 (I91080,I91357,I91518);
nand I_5226 (I91065,I91374,I91518);
nor I_5227 (I91074,I91120,I91501);
DFFARX1 I_5228 (I91501,I2683,I91094,I91083,);
not I_5229 (I91621,I2690);
DFFARX1 I_5230 (I260297,I2683,I91621,I91647,);
nand I_5231 (I91655,I260300,I260294);
and I_5232 (I91672,I91655,I260306);
DFFARX1 I_5233 (I91672,I2683,I91621,I91698,);
nor I_5234 (I91589,I91698,I91647);
not I_5235 (I91720,I91698);
DFFARX1 I_5236 (I260309,I2683,I91621,I91746,);
nand I_5237 (I91754,I91746,I260300);
not I_5238 (I91771,I91754);
DFFARX1 I_5239 (I91771,I2683,I91621,I91797,);
not I_5240 (I91613,I91797);
nor I_5241 (I91819,I91647,I91754);
nor I_5242 (I91595,I91698,I91819);
DFFARX1 I_5243 (I260312,I2683,I91621,I91859,);
DFFARX1 I_5244 (I91859,I2683,I91621,I91876,);
not I_5245 (I91884,I91876);
not I_5246 (I91901,I91859);
nand I_5247 (I91598,I91901,I91720);
nand I_5248 (I91932,I260294,I260303);
and I_5249 (I91949,I91932,I260297);
DFFARX1 I_5250 (I91949,I2683,I91621,I91975,);
nor I_5251 (I91983,I91975,I91647);
DFFARX1 I_5252 (I91983,I2683,I91621,I91586,);
DFFARX1 I_5253 (I91975,I2683,I91621,I91604,);
nor I_5254 (I92028,I260315,I260303);
not I_5255 (I92045,I92028);
nor I_5256 (I91607,I91884,I92045);
nand I_5257 (I91592,I91901,I92045);
nor I_5258 (I91601,I91647,I92028);
DFFARX1 I_5259 (I92028,I2683,I91621,I91610,);
not I_5260 (I92148,I2690);
DFFARX1 I_5261 (I418245,I2683,I92148,I92174,);
nand I_5262 (I92182,I418224,I418224);
and I_5263 (I92199,I92182,I418251);
DFFARX1 I_5264 (I92199,I2683,I92148,I92225,);
nor I_5265 (I92116,I92225,I92174);
not I_5266 (I92247,I92225);
DFFARX1 I_5267 (I418239,I2683,I92148,I92273,);
nand I_5268 (I92281,I92273,I418242);
not I_5269 (I92298,I92281);
DFFARX1 I_5270 (I92298,I2683,I92148,I92324,);
not I_5271 (I92140,I92324);
nor I_5272 (I92346,I92174,I92281);
nor I_5273 (I92122,I92225,I92346);
DFFARX1 I_5274 (I418233,I2683,I92148,I92386,);
DFFARX1 I_5275 (I92386,I2683,I92148,I92403,);
not I_5276 (I92411,I92403);
not I_5277 (I92428,I92386);
nand I_5278 (I92125,I92428,I92247);
nand I_5279 (I92459,I418230,I418227);
and I_5280 (I92476,I92459,I418248);
DFFARX1 I_5281 (I92476,I2683,I92148,I92502,);
nor I_5282 (I92510,I92502,I92174);
DFFARX1 I_5283 (I92510,I2683,I92148,I92113,);
DFFARX1 I_5284 (I92502,I2683,I92148,I92131,);
nor I_5285 (I92555,I418236,I418227);
not I_5286 (I92572,I92555);
nor I_5287 (I92134,I92411,I92572);
nand I_5288 (I92119,I92428,I92572);
nor I_5289 (I92128,I92174,I92555);
DFFARX1 I_5290 (I92555,I2683,I92148,I92137,);
not I_5291 (I92675,I2690);
DFFARX1 I_5292 (I337151,I2683,I92675,I92701,);
nand I_5293 (I92709,I337166,I337151);
and I_5294 (I92726,I92709,I337169);
DFFARX1 I_5295 (I92726,I2683,I92675,I92752,);
nor I_5296 (I92643,I92752,I92701);
not I_5297 (I92774,I92752);
DFFARX1 I_5298 (I337175,I2683,I92675,I92800,);
nand I_5299 (I92808,I92800,I337157);
not I_5300 (I92825,I92808);
DFFARX1 I_5301 (I92825,I2683,I92675,I92851,);
not I_5302 (I92667,I92851);
nor I_5303 (I92873,I92701,I92808);
nor I_5304 (I92649,I92752,I92873);
DFFARX1 I_5305 (I337154,I2683,I92675,I92913,);
DFFARX1 I_5306 (I92913,I2683,I92675,I92930,);
not I_5307 (I92938,I92930);
not I_5308 (I92955,I92913);
nand I_5309 (I92652,I92955,I92774);
nand I_5310 (I92986,I337154,I337160);
and I_5311 (I93003,I92986,I337172);
DFFARX1 I_5312 (I93003,I2683,I92675,I93029,);
nor I_5313 (I93037,I93029,I92701);
DFFARX1 I_5314 (I93037,I2683,I92675,I92640,);
DFFARX1 I_5315 (I93029,I2683,I92675,I92658,);
nor I_5316 (I93082,I337163,I337160);
not I_5317 (I93099,I93082);
nor I_5318 (I92661,I92938,I93099);
nand I_5319 (I92646,I92955,I93099);
nor I_5320 (I92655,I92701,I93082);
DFFARX1 I_5321 (I93082,I2683,I92675,I92664,);
not I_5322 (I93202,I2690);
DFFARX1 I_5323 (I299499,I2683,I93202,I93228,);
nand I_5324 (I93236,I299496,I299514);
and I_5325 (I93253,I93236,I299505);
DFFARX1 I_5326 (I93253,I2683,I93202,I93279,);
nor I_5327 (I93170,I93279,I93228);
not I_5328 (I93301,I93279);
DFFARX1 I_5329 (I299520,I2683,I93202,I93327,);
nand I_5330 (I93335,I93327,I299502);
not I_5331 (I93352,I93335);
DFFARX1 I_5332 (I93352,I2683,I93202,I93378,);
not I_5333 (I93194,I93378);
nor I_5334 (I93400,I93228,I93335);
nor I_5335 (I93176,I93279,I93400);
DFFARX1 I_5336 (I299508,I2683,I93202,I93440,);
DFFARX1 I_5337 (I93440,I2683,I93202,I93457,);
not I_5338 (I93465,I93457);
not I_5339 (I93482,I93440);
nand I_5340 (I93179,I93482,I93301);
nand I_5341 (I93513,I299496,I299523);
and I_5342 (I93530,I93513,I299511);
DFFARX1 I_5343 (I93530,I2683,I93202,I93556,);
nor I_5344 (I93564,I93556,I93228);
DFFARX1 I_5345 (I93564,I2683,I93202,I93167,);
DFFARX1 I_5346 (I93556,I2683,I93202,I93185,);
nor I_5347 (I93609,I299517,I299523);
not I_5348 (I93626,I93609);
nor I_5349 (I93188,I93465,I93626);
nand I_5350 (I93173,I93482,I93626);
nor I_5351 (I93182,I93228,I93609);
DFFARX1 I_5352 (I93609,I2683,I93202,I93191,);
not I_5353 (I93729,I2690);
DFFARX1 I_5354 (I82814,I2683,I93729,I93755,);
nand I_5355 (I93763,I82814,I82820);
and I_5356 (I93780,I93763,I82838);
DFFARX1 I_5357 (I93780,I2683,I93729,I93806,);
nor I_5358 (I93697,I93806,I93755);
not I_5359 (I93828,I93806);
DFFARX1 I_5360 (I82826,I2683,I93729,I93854,);
nand I_5361 (I93862,I93854,I82823);
not I_5362 (I93879,I93862);
DFFARX1 I_5363 (I93879,I2683,I93729,I93905,);
not I_5364 (I93721,I93905);
nor I_5365 (I93927,I93755,I93862);
nor I_5366 (I93703,I93806,I93927);
DFFARX1 I_5367 (I82832,I2683,I93729,I93967,);
DFFARX1 I_5368 (I93967,I2683,I93729,I93984,);
not I_5369 (I93992,I93984);
not I_5370 (I94009,I93967);
nand I_5371 (I93706,I94009,I93828);
nand I_5372 (I94040,I82817,I82817);
and I_5373 (I94057,I94040,I82829);
DFFARX1 I_5374 (I94057,I2683,I93729,I94083,);
nor I_5375 (I94091,I94083,I93755);
DFFARX1 I_5376 (I94091,I2683,I93729,I93694,);
DFFARX1 I_5377 (I94083,I2683,I93729,I93712,);
nor I_5378 (I94136,I82835,I82817);
not I_5379 (I94153,I94136);
nor I_5380 (I93715,I93992,I94153);
nand I_5381 (I93700,I94009,I94153);
nor I_5382 (I93709,I93755,I94136);
DFFARX1 I_5383 (I94136,I2683,I93729,I93718,);
not I_5384 (I94256,I2690);
DFFARX1 I_5385 (I388846,I2683,I94256,I94282,);
nand I_5386 (I94290,I388843,I388834);
and I_5387 (I94307,I94290,I388831);
DFFARX1 I_5388 (I94307,I2683,I94256,I94333,);
nor I_5389 (I94224,I94333,I94282);
not I_5390 (I94355,I94333);
DFFARX1 I_5391 (I388840,I2683,I94256,I94381,);
nand I_5392 (I94389,I94381,I388849);
not I_5393 (I94406,I94389);
DFFARX1 I_5394 (I94406,I2683,I94256,I94432,);
not I_5395 (I94248,I94432);
nor I_5396 (I94454,I94282,I94389);
nor I_5397 (I94230,I94333,I94454);
DFFARX1 I_5398 (I388852,I2683,I94256,I94494,);
DFFARX1 I_5399 (I94494,I2683,I94256,I94511,);
not I_5400 (I94519,I94511);
not I_5401 (I94536,I94494);
nand I_5402 (I94233,I94536,I94355);
nand I_5403 (I94567,I388831,I388837);
and I_5404 (I94584,I94567,I388855);
DFFARX1 I_5405 (I94584,I2683,I94256,I94610,);
nor I_5406 (I94618,I94610,I94282);
DFFARX1 I_5407 (I94618,I2683,I94256,I94221,);
DFFARX1 I_5408 (I94610,I2683,I94256,I94239,);
nor I_5409 (I94663,I388834,I388837);
not I_5410 (I94680,I94663);
nor I_5411 (I94242,I94519,I94680);
nand I_5412 (I94227,I94536,I94680);
nor I_5413 (I94236,I94282,I94663);
DFFARX1 I_5414 (I94663,I2683,I94256,I94245,);
not I_5415 (I94783,I2690);
DFFARX1 I_5416 (I38872,I2683,I94783,I94809,);
nand I_5417 (I94817,I38884,I38893);
and I_5418 (I94834,I94817,I38872);
DFFARX1 I_5419 (I94834,I2683,I94783,I94860,);
nor I_5420 (I94751,I94860,I94809);
not I_5421 (I94882,I94860);
DFFARX1 I_5422 (I38887,I2683,I94783,I94908,);
nand I_5423 (I94916,I94908,I38875);
not I_5424 (I94933,I94916);
DFFARX1 I_5425 (I94933,I2683,I94783,I94959,);
not I_5426 (I94775,I94959);
nor I_5427 (I94981,I94809,I94916);
nor I_5428 (I94757,I94860,I94981);
DFFARX1 I_5429 (I38878,I2683,I94783,I95021,);
DFFARX1 I_5430 (I95021,I2683,I94783,I95038,);
not I_5431 (I95046,I95038);
not I_5432 (I95063,I95021);
nand I_5433 (I94760,I95063,I94882);
nand I_5434 (I95094,I38869,I38869);
and I_5435 (I95111,I95094,I38881);
DFFARX1 I_5436 (I95111,I2683,I94783,I95137,);
nor I_5437 (I95145,I95137,I94809);
DFFARX1 I_5438 (I95145,I2683,I94783,I94748,);
DFFARX1 I_5439 (I95137,I2683,I94783,I94766,);
nor I_5440 (I95190,I38890,I38869);
not I_5441 (I95207,I95190);
nor I_5442 (I94769,I95046,I95207);
nand I_5443 (I94754,I95063,I95207);
nor I_5444 (I94763,I94809,I95190);
DFFARX1 I_5445 (I95190,I2683,I94783,I94772,);
not I_5446 (I95310,I2690);
DFFARX1 I_5447 (I330215,I2683,I95310,I95336,);
nand I_5448 (I95344,I330230,I330215);
and I_5449 (I95361,I95344,I330233);
DFFARX1 I_5450 (I95361,I2683,I95310,I95387,);
nor I_5451 (I95278,I95387,I95336);
not I_5452 (I95409,I95387);
DFFARX1 I_5453 (I330239,I2683,I95310,I95435,);
nand I_5454 (I95443,I95435,I330221);
not I_5455 (I95460,I95443);
DFFARX1 I_5456 (I95460,I2683,I95310,I95486,);
not I_5457 (I95302,I95486);
nor I_5458 (I95508,I95336,I95443);
nor I_5459 (I95284,I95387,I95508);
DFFARX1 I_5460 (I330218,I2683,I95310,I95548,);
DFFARX1 I_5461 (I95548,I2683,I95310,I95565,);
not I_5462 (I95573,I95565);
not I_5463 (I95590,I95548);
nand I_5464 (I95287,I95590,I95409);
nand I_5465 (I95621,I330218,I330224);
and I_5466 (I95638,I95621,I330236);
DFFARX1 I_5467 (I95638,I2683,I95310,I95664,);
nor I_5468 (I95672,I95664,I95336);
DFFARX1 I_5469 (I95672,I2683,I95310,I95275,);
DFFARX1 I_5470 (I95664,I2683,I95310,I95293,);
nor I_5471 (I95717,I330227,I330224);
not I_5472 (I95734,I95717);
nor I_5473 (I95296,I95573,I95734);
nand I_5474 (I95281,I95590,I95734);
nor I_5475 (I95290,I95336,I95717);
DFFARX1 I_5476 (I95717,I2683,I95310,I95299,);
not I_5477 (I95837,I2690);
DFFARX1 I_5478 (I169517,I2683,I95837,I95863,);
nand I_5479 (I95871,I169517,I169529);
and I_5480 (I95888,I95871,I169514);
DFFARX1 I_5481 (I95888,I2683,I95837,I95914,);
nor I_5482 (I95805,I95914,I95863);
not I_5483 (I95936,I95914);
DFFARX1 I_5484 (I169538,I2683,I95837,I95962,);
nand I_5485 (I95970,I95962,I169535);
not I_5486 (I95987,I95970);
DFFARX1 I_5487 (I95987,I2683,I95837,I96013,);
not I_5488 (I95829,I96013);
nor I_5489 (I96035,I95863,I95970);
nor I_5490 (I95811,I95914,I96035);
DFFARX1 I_5491 (I169526,I2683,I95837,I96075,);
DFFARX1 I_5492 (I96075,I2683,I95837,I96092,);
not I_5493 (I96100,I96092);
not I_5494 (I96117,I96075);
nand I_5495 (I95814,I96117,I95936);
nand I_5496 (I96148,I169514,I169523);
and I_5497 (I96165,I96148,I169532);
DFFARX1 I_5498 (I96165,I2683,I95837,I96191,);
nor I_5499 (I96199,I96191,I95863);
DFFARX1 I_5500 (I96199,I2683,I95837,I95802,);
DFFARX1 I_5501 (I96191,I2683,I95837,I95820,);
nor I_5502 (I96244,I169520,I169523);
not I_5503 (I96261,I96244);
nor I_5504 (I95823,I96100,I96261);
nand I_5505 (I95808,I96117,I96261);
nor I_5506 (I95817,I95863,I96244);
DFFARX1 I_5507 (I96244,I2683,I95837,I95826,);
not I_5508 (I96364,I2690);
DFFARX1 I_5509 (I58419,I2683,I96364,I96390,);
nand I_5510 (I96398,I58419,I58425);
and I_5511 (I96415,I96398,I58443);
DFFARX1 I_5512 (I96415,I2683,I96364,I96441,);
nor I_5513 (I96332,I96441,I96390);
not I_5514 (I96463,I96441);
DFFARX1 I_5515 (I58431,I2683,I96364,I96489,);
nand I_5516 (I96497,I96489,I58428);
not I_5517 (I96514,I96497);
DFFARX1 I_5518 (I96514,I2683,I96364,I96540,);
not I_5519 (I96356,I96540);
nor I_5520 (I96562,I96390,I96497);
nor I_5521 (I96338,I96441,I96562);
DFFARX1 I_5522 (I58437,I2683,I96364,I96602,);
DFFARX1 I_5523 (I96602,I2683,I96364,I96619,);
not I_5524 (I96627,I96619);
not I_5525 (I96644,I96602);
nand I_5526 (I96341,I96644,I96463);
nand I_5527 (I96675,I58422,I58422);
and I_5528 (I96692,I96675,I58434);
DFFARX1 I_5529 (I96692,I2683,I96364,I96718,);
nor I_5530 (I96726,I96718,I96390);
DFFARX1 I_5531 (I96726,I2683,I96364,I96329,);
DFFARX1 I_5532 (I96718,I2683,I96364,I96347,);
nor I_5533 (I96771,I58440,I58422);
not I_5534 (I96788,I96771);
nor I_5535 (I96350,I96627,I96788);
nand I_5536 (I96335,I96644,I96788);
nor I_5537 (I96344,I96390,I96771);
DFFARX1 I_5538 (I96771,I2683,I96364,I96353,);
not I_5539 (I96891,I2690);
DFFARX1 I_5540 (I294977,I2683,I96891,I96917,);
nand I_5541 (I96925,I294974,I294992);
and I_5542 (I96942,I96925,I294983);
DFFARX1 I_5543 (I96942,I2683,I96891,I96968,);
nor I_5544 (I96859,I96968,I96917);
not I_5545 (I96990,I96968);
DFFARX1 I_5546 (I294998,I2683,I96891,I97016,);
nand I_5547 (I97024,I97016,I294980);
not I_5548 (I97041,I97024);
DFFARX1 I_5549 (I97041,I2683,I96891,I97067,);
not I_5550 (I96883,I97067);
nor I_5551 (I97089,I96917,I97024);
nor I_5552 (I96865,I96968,I97089);
DFFARX1 I_5553 (I294986,I2683,I96891,I97129,);
DFFARX1 I_5554 (I97129,I2683,I96891,I97146,);
not I_5555 (I97154,I97146);
not I_5556 (I97171,I97129);
nand I_5557 (I96868,I97171,I96990);
nand I_5558 (I97202,I294974,I295001);
and I_5559 (I97219,I97202,I294989);
DFFARX1 I_5560 (I97219,I2683,I96891,I97245,);
nor I_5561 (I97253,I97245,I96917);
DFFARX1 I_5562 (I97253,I2683,I96891,I96856,);
DFFARX1 I_5563 (I97245,I2683,I96891,I96874,);
nor I_5564 (I97298,I294995,I295001);
not I_5565 (I97315,I97298);
nor I_5566 (I96877,I97154,I97315);
nand I_5567 (I96862,I97171,I97315);
nor I_5568 (I96871,I96917,I97298);
DFFARX1 I_5569 (I97298,I2683,I96891,I96880,);
not I_5570 (I97418,I2690);
DFFARX1 I_5571 (I387690,I2683,I97418,I97444,);
nand I_5572 (I97452,I387687,I387678);
and I_5573 (I97469,I97452,I387675);
DFFARX1 I_5574 (I97469,I2683,I97418,I97495,);
nor I_5575 (I97386,I97495,I97444);
not I_5576 (I97517,I97495);
DFFARX1 I_5577 (I387684,I2683,I97418,I97543,);
nand I_5578 (I97551,I97543,I387693);
not I_5579 (I97568,I97551);
DFFARX1 I_5580 (I97568,I2683,I97418,I97594,);
not I_5581 (I97410,I97594);
nor I_5582 (I97616,I97444,I97551);
nor I_5583 (I97392,I97495,I97616);
DFFARX1 I_5584 (I387696,I2683,I97418,I97656,);
DFFARX1 I_5585 (I97656,I2683,I97418,I97673,);
not I_5586 (I97681,I97673);
not I_5587 (I97698,I97656);
nand I_5588 (I97395,I97698,I97517);
nand I_5589 (I97729,I387675,I387681);
and I_5590 (I97746,I97729,I387699);
DFFARX1 I_5591 (I97746,I2683,I97418,I97772,);
nor I_5592 (I97780,I97772,I97444);
DFFARX1 I_5593 (I97780,I2683,I97418,I97383,);
DFFARX1 I_5594 (I97772,I2683,I97418,I97401,);
nor I_5595 (I97825,I387678,I387681);
not I_5596 (I97842,I97825);
nor I_5597 (I97404,I97681,I97842);
nand I_5598 (I97389,I97698,I97842);
nor I_5599 (I97398,I97444,I97825);
DFFARX1 I_5600 (I97825,I2683,I97418,I97407,);
not I_5601 (I97945,I2690);
DFFARX1 I_5602 (I57229,I2683,I97945,I97971,);
nand I_5603 (I97979,I57229,I57235);
and I_5604 (I97996,I97979,I57253);
DFFARX1 I_5605 (I97996,I2683,I97945,I98022,);
nor I_5606 (I97913,I98022,I97971);
not I_5607 (I98044,I98022);
DFFARX1 I_5608 (I57241,I2683,I97945,I98070,);
nand I_5609 (I98078,I98070,I57238);
not I_5610 (I98095,I98078);
DFFARX1 I_5611 (I98095,I2683,I97945,I98121,);
not I_5612 (I97937,I98121);
nor I_5613 (I98143,I97971,I98078);
nor I_5614 (I97919,I98022,I98143);
DFFARX1 I_5615 (I57247,I2683,I97945,I98183,);
DFFARX1 I_5616 (I98183,I2683,I97945,I98200,);
not I_5617 (I98208,I98200);
not I_5618 (I98225,I98183);
nand I_5619 (I97922,I98225,I98044);
nand I_5620 (I98256,I57232,I57232);
and I_5621 (I98273,I98256,I57244);
DFFARX1 I_5622 (I98273,I2683,I97945,I98299,);
nor I_5623 (I98307,I98299,I97971);
DFFARX1 I_5624 (I98307,I2683,I97945,I97910,);
DFFARX1 I_5625 (I98299,I2683,I97945,I97928,);
nor I_5626 (I98352,I57250,I57232);
not I_5627 (I98369,I98352);
nor I_5628 (I97931,I98208,I98369);
nand I_5629 (I97916,I98225,I98369);
nor I_5630 (I97925,I97971,I98352);
DFFARX1 I_5631 (I98352,I2683,I97945,I97934,);
not I_5632 (I98472,I2690);
DFFARX1 I_5633 (I307251,I2683,I98472,I98498,);
nand I_5634 (I98506,I307248,I307266);
and I_5635 (I98523,I98506,I307257);
DFFARX1 I_5636 (I98523,I2683,I98472,I98549,);
nor I_5637 (I98440,I98549,I98498);
not I_5638 (I98571,I98549);
DFFARX1 I_5639 (I307272,I2683,I98472,I98597,);
nand I_5640 (I98605,I98597,I307254);
not I_5641 (I98622,I98605);
DFFARX1 I_5642 (I98622,I2683,I98472,I98648,);
not I_5643 (I98464,I98648);
nor I_5644 (I98670,I98498,I98605);
nor I_5645 (I98446,I98549,I98670);
DFFARX1 I_5646 (I307260,I2683,I98472,I98710,);
DFFARX1 I_5647 (I98710,I2683,I98472,I98727,);
not I_5648 (I98735,I98727);
not I_5649 (I98752,I98710);
nand I_5650 (I98449,I98752,I98571);
nand I_5651 (I98783,I307248,I307275);
and I_5652 (I98800,I98783,I307263);
DFFARX1 I_5653 (I98800,I2683,I98472,I98826,);
nor I_5654 (I98834,I98826,I98498);
DFFARX1 I_5655 (I98834,I2683,I98472,I98437,);
DFFARX1 I_5656 (I98826,I2683,I98472,I98455,);
nor I_5657 (I98879,I307269,I307275);
not I_5658 (I98896,I98879);
nor I_5659 (I98458,I98735,I98896);
nand I_5660 (I98443,I98752,I98896);
nor I_5661 (I98452,I98498,I98879);
DFFARX1 I_5662 (I98879,I2683,I98472,I98461,);
not I_5663 (I98999,I2690);
DFFARX1 I_5664 (I405155,I2683,I98999,I99025,);
nand I_5665 (I99033,I405134,I405134);
and I_5666 (I99050,I99033,I405161);
DFFARX1 I_5667 (I99050,I2683,I98999,I99076,);
nor I_5668 (I98967,I99076,I99025);
not I_5669 (I99098,I99076);
DFFARX1 I_5670 (I405149,I2683,I98999,I99124,);
nand I_5671 (I99132,I99124,I405152);
not I_5672 (I99149,I99132);
DFFARX1 I_5673 (I99149,I2683,I98999,I99175,);
not I_5674 (I98991,I99175);
nor I_5675 (I99197,I99025,I99132);
nor I_5676 (I98973,I99076,I99197);
DFFARX1 I_5677 (I405143,I2683,I98999,I99237,);
DFFARX1 I_5678 (I99237,I2683,I98999,I99254,);
not I_5679 (I99262,I99254);
not I_5680 (I99279,I99237);
nand I_5681 (I98976,I99279,I99098);
nand I_5682 (I99310,I405140,I405137);
and I_5683 (I99327,I99310,I405158);
DFFARX1 I_5684 (I99327,I2683,I98999,I99353,);
nor I_5685 (I99361,I99353,I99025);
DFFARX1 I_5686 (I99361,I2683,I98999,I98964,);
DFFARX1 I_5687 (I99353,I2683,I98999,I98982,);
nor I_5688 (I99406,I405146,I405137);
not I_5689 (I99423,I99406);
nor I_5690 (I98985,I99262,I99423);
nand I_5691 (I98970,I99279,I99423);
nor I_5692 (I98979,I99025,I99406);
DFFARX1 I_5693 (I99406,I2683,I98999,I98988,);
not I_5694 (I99526,I2690);
DFFARX1 I_5695 (I130171,I2683,I99526,I99552,);
nand I_5696 (I99560,I130183,I130162);
and I_5697 (I99577,I99560,I130186);
DFFARX1 I_5698 (I99577,I2683,I99526,I99603,);
nor I_5699 (I99494,I99603,I99552);
not I_5700 (I99625,I99603);
DFFARX1 I_5701 (I130177,I2683,I99526,I99651,);
nand I_5702 (I99659,I99651,I130159);
not I_5703 (I99676,I99659);
DFFARX1 I_5704 (I99676,I2683,I99526,I99702,);
not I_5705 (I99518,I99702);
nor I_5706 (I99724,I99552,I99659);
nor I_5707 (I99500,I99603,I99724);
DFFARX1 I_5708 (I130174,I2683,I99526,I99764,);
DFFARX1 I_5709 (I99764,I2683,I99526,I99781,);
not I_5710 (I99789,I99781);
not I_5711 (I99806,I99764);
nand I_5712 (I99503,I99806,I99625);
nand I_5713 (I99837,I130159,I130165);
and I_5714 (I99854,I99837,I130168);
DFFARX1 I_5715 (I99854,I2683,I99526,I99880,);
nor I_5716 (I99888,I99880,I99552);
DFFARX1 I_5717 (I99888,I2683,I99526,I99491,);
DFFARX1 I_5718 (I99880,I2683,I99526,I99509,);
nor I_5719 (I99933,I130180,I130165);
not I_5720 (I99950,I99933);
nor I_5721 (I99512,I99789,I99950);
nand I_5722 (I99497,I99806,I99950);
nor I_5723 (I99506,I99552,I99933);
DFFARX1 I_5724 (I99933,I2683,I99526,I99515,);
not I_5725 (I100053,I2690);
DFFARX1 I_5726 (I204223,I2683,I100053,I100079,);
nand I_5727 (I100087,I204214,I204229);
and I_5728 (I100104,I100087,I204235);
DFFARX1 I_5729 (I100104,I2683,I100053,I100130,);
nor I_5730 (I100021,I100130,I100079);
not I_5731 (I100152,I100130);
DFFARX1 I_5732 (I204220,I2683,I100053,I100178,);
nand I_5733 (I100186,I100178,I204214);
not I_5734 (I100203,I100186);
DFFARX1 I_5735 (I100203,I2683,I100053,I100229,);
not I_5736 (I100045,I100229);
nor I_5737 (I100251,I100079,I100186);
nor I_5738 (I100027,I100130,I100251);
DFFARX1 I_5739 (I204217,I2683,I100053,I100291,);
DFFARX1 I_5740 (I100291,I2683,I100053,I100308,);
not I_5741 (I100316,I100308);
not I_5742 (I100333,I100291);
nand I_5743 (I100030,I100333,I100152);
nand I_5744 (I100364,I204211,I204226);
and I_5745 (I100381,I100364,I204211);
DFFARX1 I_5746 (I100381,I2683,I100053,I100407,);
nor I_5747 (I100415,I100407,I100079);
DFFARX1 I_5748 (I100415,I2683,I100053,I100018,);
DFFARX1 I_5749 (I100407,I2683,I100053,I100036,);
nor I_5750 (I100460,I204232,I204226);
not I_5751 (I100477,I100460);
nor I_5752 (I100039,I100316,I100477);
nand I_5753 (I100024,I100333,I100477);
nor I_5754 (I100033,I100079,I100460);
DFFARX1 I_5755 (I100460,I2683,I100053,I100042,);
not I_5756 (I100580,I2690);
DFFARX1 I_5757 (I310396,I2683,I100580,I100606,);
nand I_5758 (I100614,I310393,I310396);
and I_5759 (I100631,I100614,I310405);
DFFARX1 I_5760 (I100631,I2683,I100580,I100657,);
nor I_5761 (I100548,I100657,I100606);
not I_5762 (I100679,I100657);
DFFARX1 I_5763 (I310393,I2683,I100580,I100705,);
nand I_5764 (I100713,I100705,I310411);
not I_5765 (I100730,I100713);
DFFARX1 I_5766 (I100730,I2683,I100580,I100756,);
not I_5767 (I100572,I100756);
nor I_5768 (I100778,I100606,I100713);
nor I_5769 (I100554,I100657,I100778);
DFFARX1 I_5770 (I310399,I2683,I100580,I100818,);
DFFARX1 I_5771 (I100818,I2683,I100580,I100835,);
not I_5772 (I100843,I100835);
not I_5773 (I100860,I100818);
nand I_5774 (I100557,I100860,I100679);
nand I_5775 (I100891,I310408,I310414);
and I_5776 (I100908,I100891,I310399);
DFFARX1 I_5777 (I100908,I2683,I100580,I100934,);
nor I_5778 (I100942,I100934,I100606);
DFFARX1 I_5779 (I100942,I2683,I100580,I100545,);
DFFARX1 I_5780 (I100934,I2683,I100580,I100563,);
nor I_5781 (I100987,I310402,I310414);
not I_5782 (I101004,I100987);
nor I_5783 (I100566,I100843,I101004);
nand I_5784 (I100551,I100860,I101004);
nor I_5785 (I100560,I100606,I100987);
DFFARX1 I_5786 (I100987,I2683,I100580,I100569,);
not I_5787 (I101107,I2690);
DFFARX1 I_5788 (I316006,I2683,I101107,I101133,);
nand I_5789 (I101141,I316003,I316006);
and I_5790 (I101158,I101141,I316015);
DFFARX1 I_5791 (I101158,I2683,I101107,I101184,);
nor I_5792 (I101075,I101184,I101133);
not I_5793 (I101206,I101184);
DFFARX1 I_5794 (I316003,I2683,I101107,I101232,);
nand I_5795 (I101240,I101232,I316021);
not I_5796 (I101257,I101240);
DFFARX1 I_5797 (I101257,I2683,I101107,I101283,);
not I_5798 (I101099,I101283);
nor I_5799 (I101305,I101133,I101240);
nor I_5800 (I101081,I101184,I101305);
DFFARX1 I_5801 (I316009,I2683,I101107,I101345,);
DFFARX1 I_5802 (I101345,I2683,I101107,I101362,);
not I_5803 (I101370,I101362);
not I_5804 (I101387,I101345);
nand I_5805 (I101084,I101387,I101206);
nand I_5806 (I101418,I316018,I316024);
and I_5807 (I101435,I101418,I316009);
DFFARX1 I_5808 (I101435,I2683,I101107,I101461,);
nor I_5809 (I101469,I101461,I101133);
DFFARX1 I_5810 (I101469,I2683,I101107,I101072,);
DFFARX1 I_5811 (I101461,I2683,I101107,I101090,);
nor I_5812 (I101514,I316012,I316024);
not I_5813 (I101531,I101514);
nor I_5814 (I101093,I101370,I101531);
nand I_5815 (I101078,I101387,I101531);
nor I_5816 (I101087,I101133,I101514);
DFFARX1 I_5817 (I101514,I2683,I101107,I101096,);
not I_5818 (I101634,I2690);
DFFARX1 I_5819 (I314884,I2683,I101634,I101660,);
nand I_5820 (I101668,I314881,I314884);
and I_5821 (I101685,I101668,I314893);
DFFARX1 I_5822 (I101685,I2683,I101634,I101711,);
nor I_5823 (I101602,I101711,I101660);
not I_5824 (I101733,I101711);
DFFARX1 I_5825 (I314881,I2683,I101634,I101759,);
nand I_5826 (I101767,I101759,I314899);
not I_5827 (I101784,I101767);
DFFARX1 I_5828 (I101784,I2683,I101634,I101810,);
not I_5829 (I101626,I101810);
nor I_5830 (I101832,I101660,I101767);
nor I_5831 (I101608,I101711,I101832);
DFFARX1 I_5832 (I314887,I2683,I101634,I101872,);
DFFARX1 I_5833 (I101872,I2683,I101634,I101889,);
not I_5834 (I101897,I101889);
not I_5835 (I101914,I101872);
nand I_5836 (I101611,I101914,I101733);
nand I_5837 (I101945,I314896,I314902);
and I_5838 (I101962,I101945,I314887);
DFFARX1 I_5839 (I101962,I2683,I101634,I101988,);
nor I_5840 (I101996,I101988,I101660);
DFFARX1 I_5841 (I101996,I2683,I101634,I101599,);
DFFARX1 I_5842 (I101988,I2683,I101634,I101617,);
nor I_5843 (I102041,I314890,I314902);
not I_5844 (I102058,I102041);
nor I_5845 (I101620,I101897,I102058);
nand I_5846 (I101605,I101914,I102058);
nor I_5847 (I101614,I101660,I102041);
DFFARX1 I_5848 (I102041,I2683,I101634,I101623,);
not I_5849 (I102161,I2690);
DFFARX1 I_5850 (I24116,I2683,I102161,I102187,);
nand I_5851 (I102195,I24128,I24137);
and I_5852 (I102212,I102195,I24116);
DFFARX1 I_5853 (I102212,I2683,I102161,I102238,);
nor I_5854 (I102129,I102238,I102187);
not I_5855 (I102260,I102238);
DFFARX1 I_5856 (I24131,I2683,I102161,I102286,);
nand I_5857 (I102294,I102286,I24119);
not I_5858 (I102311,I102294);
DFFARX1 I_5859 (I102311,I2683,I102161,I102337,);
not I_5860 (I102153,I102337);
nor I_5861 (I102359,I102187,I102294);
nor I_5862 (I102135,I102238,I102359);
DFFARX1 I_5863 (I24122,I2683,I102161,I102399,);
DFFARX1 I_5864 (I102399,I2683,I102161,I102416,);
not I_5865 (I102424,I102416);
not I_5866 (I102441,I102399);
nand I_5867 (I102138,I102441,I102260);
nand I_5868 (I102472,I24113,I24113);
and I_5869 (I102489,I102472,I24125);
DFFARX1 I_5870 (I102489,I2683,I102161,I102515,);
nor I_5871 (I102523,I102515,I102187);
DFFARX1 I_5872 (I102523,I2683,I102161,I102126,);
DFFARX1 I_5873 (I102515,I2683,I102161,I102144,);
nor I_5874 (I102568,I24134,I24113);
not I_5875 (I102585,I102568);
nor I_5876 (I102147,I102424,I102585);
nand I_5877 (I102132,I102441,I102585);
nor I_5878 (I102141,I102187,I102568);
DFFARX1 I_5879 (I102568,I2683,I102161,I102150,);
not I_5880 (I102688,I2690);
DFFARX1 I_5881 (I29913,I2683,I102688,I102714,);
nand I_5882 (I102722,I29925,I29934);
and I_5883 (I102739,I102722,I29913);
DFFARX1 I_5884 (I102739,I2683,I102688,I102765,);
nor I_5885 (I102656,I102765,I102714);
not I_5886 (I102787,I102765);
DFFARX1 I_5887 (I29928,I2683,I102688,I102813,);
nand I_5888 (I102821,I102813,I29916);
not I_5889 (I102838,I102821);
DFFARX1 I_5890 (I102838,I2683,I102688,I102864,);
not I_5891 (I102680,I102864);
nor I_5892 (I102886,I102714,I102821);
nor I_5893 (I102662,I102765,I102886);
DFFARX1 I_5894 (I29919,I2683,I102688,I102926,);
DFFARX1 I_5895 (I102926,I2683,I102688,I102943,);
not I_5896 (I102951,I102943);
not I_5897 (I102968,I102926);
nand I_5898 (I102665,I102968,I102787);
nand I_5899 (I102999,I29910,I29910);
and I_5900 (I103016,I102999,I29922);
DFFARX1 I_5901 (I103016,I2683,I102688,I103042,);
nor I_5902 (I103050,I103042,I102714);
DFFARX1 I_5903 (I103050,I2683,I102688,I102653,);
DFFARX1 I_5904 (I103042,I2683,I102688,I102671,);
nor I_5905 (I103095,I29931,I29910);
not I_5906 (I103112,I103095);
nor I_5907 (I102674,I102951,I103112);
nand I_5908 (I102659,I102968,I103112);
nor I_5909 (I102668,I102714,I103095);
DFFARX1 I_5910 (I103095,I2683,I102688,I102677,);
not I_5911 (I103215,I2690);
DFFARX1 I_5912 (I371951,I2683,I103215,I103241,);
nand I_5913 (I103249,I371933,I371957);
and I_5914 (I103266,I103249,I371948);
DFFARX1 I_5915 (I103266,I2683,I103215,I103292,);
nor I_5916 (I103183,I103292,I103241);
not I_5917 (I103314,I103292);
DFFARX1 I_5918 (I371954,I2683,I103215,I103340,);
nand I_5919 (I103348,I103340,I371942);
not I_5920 (I103365,I103348);
DFFARX1 I_5921 (I103365,I2683,I103215,I103391,);
not I_5922 (I103207,I103391);
nor I_5923 (I103413,I103241,I103348);
nor I_5924 (I103189,I103292,I103413);
DFFARX1 I_5925 (I371933,I2683,I103215,I103453,);
DFFARX1 I_5926 (I103453,I2683,I103215,I103470,);
not I_5927 (I103478,I103470);
not I_5928 (I103495,I103453);
nand I_5929 (I103192,I103495,I103314);
nand I_5930 (I103526,I371939,I371936);
and I_5931 (I103543,I103526,I371945);
DFFARX1 I_5932 (I103543,I2683,I103215,I103569,);
nor I_5933 (I103577,I103569,I103241);
DFFARX1 I_5934 (I103577,I2683,I103215,I103180,);
DFFARX1 I_5935 (I103569,I2683,I103215,I103198,);
nor I_5936 (I103622,I371936,I371936);
not I_5937 (I103639,I103622);
nor I_5938 (I103201,I103478,I103639);
nand I_5939 (I103186,I103495,I103639);
nor I_5940 (I103195,I103241,I103622);
DFFARX1 I_5941 (I103622,I2683,I103215,I103204,);
not I_5942 (I103742,I2690);
DFFARX1 I_5943 (I364335,I2683,I103742,I103768,);
nand I_5944 (I103776,I364317,I364341);
and I_5945 (I103793,I103776,I364332);
DFFARX1 I_5946 (I103793,I2683,I103742,I103819,);
nor I_5947 (I103710,I103819,I103768);
not I_5948 (I103841,I103819);
DFFARX1 I_5949 (I364338,I2683,I103742,I103867,);
nand I_5950 (I103875,I103867,I364326);
not I_5951 (I103892,I103875);
DFFARX1 I_5952 (I103892,I2683,I103742,I103918,);
not I_5953 (I103734,I103918);
nor I_5954 (I103940,I103768,I103875);
nor I_5955 (I103716,I103819,I103940);
DFFARX1 I_5956 (I364317,I2683,I103742,I103980,);
DFFARX1 I_5957 (I103980,I2683,I103742,I103997,);
not I_5958 (I104005,I103997);
not I_5959 (I104022,I103980);
nand I_5960 (I103719,I104022,I103841);
nand I_5961 (I104053,I364323,I364320);
and I_5962 (I104070,I104053,I364329);
DFFARX1 I_5963 (I104070,I2683,I103742,I104096,);
nor I_5964 (I104104,I104096,I103768);
DFFARX1 I_5965 (I104104,I2683,I103742,I103707,);
DFFARX1 I_5966 (I104096,I2683,I103742,I103725,);
nor I_5967 (I104149,I364320,I364320);
not I_5968 (I104166,I104149);
nor I_5969 (I103728,I104005,I104166);
nand I_5970 (I103713,I104022,I104166);
nor I_5971 (I103722,I103768,I104149);
DFFARX1 I_5972 (I104149,I2683,I103742,I103731,);
not I_5973 (I104269,I2690);
DFFARX1 I_5974 (I171280,I2683,I104269,I104295,);
nand I_5975 (I104303,I171265,I171268);
and I_5976 (I104320,I104303,I171283);
DFFARX1 I_5977 (I104320,I2683,I104269,I104346,);
nor I_5978 (I104237,I104346,I104295);
not I_5979 (I104368,I104346);
DFFARX1 I_5980 (I171277,I2683,I104269,I104394,);
nand I_5981 (I104402,I104394,I171268);
not I_5982 (I104419,I104402);
DFFARX1 I_5983 (I104419,I2683,I104269,I104445,);
not I_5984 (I104261,I104445);
nor I_5985 (I104467,I104295,I104402);
nor I_5986 (I104243,I104346,I104467);
DFFARX1 I_5987 (I171274,I2683,I104269,I104507,);
DFFARX1 I_5988 (I104507,I2683,I104269,I104524,);
not I_5989 (I104532,I104524);
not I_5990 (I104549,I104507);
nand I_5991 (I104246,I104549,I104368);
nand I_5992 (I104580,I171289,I171265);
and I_5993 (I104597,I104580,I171286);
DFFARX1 I_5994 (I104597,I2683,I104269,I104623,);
nor I_5995 (I104631,I104623,I104295);
DFFARX1 I_5996 (I104631,I2683,I104269,I104234,);
DFFARX1 I_5997 (I104623,I2683,I104269,I104252,);
nor I_5998 (I104676,I171271,I171265);
not I_5999 (I104693,I104676);
nor I_6000 (I104255,I104532,I104693);
nand I_6001 (I104240,I104549,I104693);
nor I_6002 (I104249,I104295,I104676);
DFFARX1 I_6003 (I104676,I2683,I104269,I104258,);
not I_6004 (I104796,I2690);
DFFARX1 I_6005 (I43615,I2683,I104796,I104822,);
nand I_6006 (I104830,I43627,I43636);
and I_6007 (I104847,I104830,I43615);
DFFARX1 I_6008 (I104847,I2683,I104796,I104873,);
nor I_6009 (I104764,I104873,I104822);
not I_6010 (I104895,I104873);
DFFARX1 I_6011 (I43630,I2683,I104796,I104921,);
nand I_6012 (I104929,I104921,I43618);
not I_6013 (I104946,I104929);
DFFARX1 I_6014 (I104946,I2683,I104796,I104972,);
not I_6015 (I104788,I104972);
nor I_6016 (I104994,I104822,I104929);
nor I_6017 (I104770,I104873,I104994);
DFFARX1 I_6018 (I43621,I2683,I104796,I105034,);
DFFARX1 I_6019 (I105034,I2683,I104796,I105051,);
not I_6020 (I105059,I105051);
not I_6021 (I105076,I105034);
nand I_6022 (I104773,I105076,I104895);
nand I_6023 (I105107,I43612,I43612);
and I_6024 (I105124,I105107,I43624);
DFFARX1 I_6025 (I105124,I2683,I104796,I105150,);
nor I_6026 (I105158,I105150,I104822);
DFFARX1 I_6027 (I105158,I2683,I104796,I104761,);
DFFARX1 I_6028 (I105150,I2683,I104796,I104779,);
nor I_6029 (I105203,I43633,I43612);
not I_6030 (I105220,I105203);
nor I_6031 (I104782,I105059,I105220);
nand I_6032 (I104767,I105076,I105220);
nor I_6033 (I104776,I104822,I105203);
DFFARX1 I_6034 (I105203,I2683,I104796,I104785,);
not I_6035 (I105323,I2690);
DFFARX1 I_6036 (I1564,I2683,I105323,I105349,);
nand I_6037 (I105357,I1788,I2364);
and I_6038 (I105374,I105357,I2284);
DFFARX1 I_6039 (I105374,I2683,I105323,I105400,);
nor I_6040 (I105291,I105400,I105349);
not I_6041 (I105422,I105400);
DFFARX1 I_6042 (I2572,I2683,I105323,I105448,);
nand I_6043 (I105456,I105448,I1484);
not I_6044 (I105473,I105456);
DFFARX1 I_6045 (I105473,I2683,I105323,I105499,);
not I_6046 (I105315,I105499);
nor I_6047 (I105521,I105349,I105456);
nor I_6048 (I105297,I105400,I105521);
DFFARX1 I_6049 (I1644,I2683,I105323,I105561,);
DFFARX1 I_6050 (I105561,I2683,I105323,I105578,);
not I_6051 (I105586,I105578);
not I_6052 (I105603,I105561);
nand I_6053 (I105300,I105603,I105422);
nand I_6054 (I105634,I2532,I2356);
and I_6055 (I105651,I105634,I1748);
DFFARX1 I_6056 (I105651,I2683,I105323,I105677,);
nor I_6057 (I105685,I105677,I105349);
DFFARX1 I_6058 (I105685,I2683,I105323,I105288,);
DFFARX1 I_6059 (I105677,I2683,I105323,I105306,);
nor I_6060 (I105730,I2156,I2356);
not I_6061 (I105747,I105730);
nor I_6062 (I105309,I105586,I105747);
nand I_6063 (I105294,I105603,I105747);
nor I_6064 (I105303,I105349,I105730);
DFFARX1 I_6065 (I105730,I2683,I105323,I105312,);
not I_6066 (I105850,I2690);
DFFARX1 I_6067 (I241325,I2683,I105850,I105876,);
nand I_6068 (I105884,I241328,I241322);
and I_6069 (I105901,I105884,I241334);
DFFARX1 I_6070 (I105901,I2683,I105850,I105927,);
nor I_6071 (I105818,I105927,I105876);
not I_6072 (I105949,I105927);
DFFARX1 I_6073 (I241337,I2683,I105850,I105975,);
nand I_6074 (I105983,I105975,I241328);
not I_6075 (I106000,I105983);
DFFARX1 I_6076 (I106000,I2683,I105850,I106026,);
not I_6077 (I105842,I106026);
nor I_6078 (I106048,I105876,I105983);
nor I_6079 (I105824,I105927,I106048);
DFFARX1 I_6080 (I241340,I2683,I105850,I106088,);
DFFARX1 I_6081 (I106088,I2683,I105850,I106105,);
not I_6082 (I106113,I106105);
not I_6083 (I106130,I106088);
nand I_6084 (I105827,I106130,I105949);
nand I_6085 (I106161,I241322,I241331);
and I_6086 (I106178,I106161,I241325);
DFFARX1 I_6087 (I106178,I2683,I105850,I106204,);
nor I_6088 (I106212,I106204,I105876);
DFFARX1 I_6089 (I106212,I2683,I105850,I105815,);
DFFARX1 I_6090 (I106204,I2683,I105850,I105833,);
nor I_6091 (I106257,I241343,I241331);
not I_6092 (I106274,I106257);
nor I_6093 (I105836,I106113,I106274);
nand I_6094 (I105821,I106130,I106274);
nor I_6095 (I105830,I105876,I106257);
DFFARX1 I_6096 (I106257,I2683,I105850,I105839,);
not I_6097 (I106377,I2690);
DFFARX1 I_6098 (I303375,I2683,I106377,I106403,);
nand I_6099 (I106411,I303372,I303390);
and I_6100 (I106428,I106411,I303381);
DFFARX1 I_6101 (I106428,I2683,I106377,I106454,);
nor I_6102 (I106345,I106454,I106403);
not I_6103 (I106476,I106454);
DFFARX1 I_6104 (I303396,I2683,I106377,I106502,);
nand I_6105 (I106510,I106502,I303378);
not I_6106 (I106527,I106510);
DFFARX1 I_6107 (I106527,I2683,I106377,I106553,);
not I_6108 (I106369,I106553);
nor I_6109 (I106575,I106403,I106510);
nor I_6110 (I106351,I106454,I106575);
DFFARX1 I_6111 (I303384,I2683,I106377,I106615,);
DFFARX1 I_6112 (I106615,I2683,I106377,I106632,);
not I_6113 (I106640,I106632);
not I_6114 (I106657,I106615);
nand I_6115 (I106354,I106657,I106476);
nand I_6116 (I106688,I303372,I303399);
and I_6117 (I106705,I106688,I303387);
DFFARX1 I_6118 (I106705,I2683,I106377,I106731,);
nor I_6119 (I106739,I106731,I106403);
DFFARX1 I_6120 (I106739,I2683,I106377,I106342,);
DFFARX1 I_6121 (I106731,I2683,I106377,I106360,);
nor I_6122 (I106784,I303393,I303399);
not I_6123 (I106801,I106784);
nor I_6124 (I106363,I106640,I106801);
nand I_6125 (I106348,I106657,I106801);
nor I_6126 (I106357,I106403,I106784);
DFFARX1 I_6127 (I106784,I2683,I106377,I106366,);
not I_6128 (I106904,I2690);
DFFARX1 I_6129 (I352179,I2683,I106904,I106930,);
nand I_6130 (I106938,I352194,I352179);
and I_6131 (I106955,I106938,I352197);
DFFARX1 I_6132 (I106955,I2683,I106904,I106981,);
nor I_6133 (I106872,I106981,I106930);
not I_6134 (I107003,I106981);
DFFARX1 I_6135 (I352203,I2683,I106904,I107029,);
nand I_6136 (I107037,I107029,I352185);
not I_6137 (I107054,I107037);
DFFARX1 I_6138 (I107054,I2683,I106904,I107080,);
not I_6139 (I106896,I107080);
nor I_6140 (I107102,I106930,I107037);
nor I_6141 (I106878,I106981,I107102);
DFFARX1 I_6142 (I352182,I2683,I106904,I107142,);
DFFARX1 I_6143 (I107142,I2683,I106904,I107159,);
not I_6144 (I107167,I107159);
not I_6145 (I107184,I107142);
nand I_6146 (I106881,I107184,I107003);
nand I_6147 (I107215,I352182,I352188);
and I_6148 (I107232,I107215,I352200);
DFFARX1 I_6149 (I107232,I2683,I106904,I107258,);
nor I_6150 (I107266,I107258,I106930);
DFFARX1 I_6151 (I107266,I2683,I106904,I106869,);
DFFARX1 I_6152 (I107258,I2683,I106904,I106887,);
nor I_6153 (I107311,I352191,I352188);
not I_6154 (I107328,I107311);
nor I_6155 (I106890,I107167,I107328);
nand I_6156 (I106875,I107184,I107328);
nor I_6157 (I106884,I106930,I107311);
DFFARX1 I_6158 (I107311,I2683,I106904,I106893,);
not I_6159 (I107431,I2690);
DFFARX1 I_6160 (I145947,I2683,I107431,I107457,);
nand I_6161 (I107465,I145959,I145938);
and I_6162 (I107482,I107465,I145962);
DFFARX1 I_6163 (I107482,I2683,I107431,I107508,);
nor I_6164 (I107399,I107508,I107457);
not I_6165 (I107530,I107508);
DFFARX1 I_6166 (I145953,I2683,I107431,I107556,);
nand I_6167 (I107564,I107556,I145935);
not I_6168 (I107581,I107564);
DFFARX1 I_6169 (I107581,I2683,I107431,I107607,);
not I_6170 (I107423,I107607);
nor I_6171 (I107629,I107457,I107564);
nor I_6172 (I107405,I107508,I107629);
DFFARX1 I_6173 (I145950,I2683,I107431,I107669,);
DFFARX1 I_6174 (I107669,I2683,I107431,I107686,);
not I_6175 (I107694,I107686);
not I_6176 (I107711,I107669);
nand I_6177 (I107408,I107711,I107530);
nand I_6178 (I107742,I145935,I145941);
and I_6179 (I107759,I107742,I145944);
DFFARX1 I_6180 (I107759,I2683,I107431,I107785,);
nor I_6181 (I107793,I107785,I107457);
DFFARX1 I_6182 (I107793,I2683,I107431,I107396,);
DFFARX1 I_6183 (I107785,I2683,I107431,I107414,);
nor I_6184 (I107838,I145956,I145941);
not I_6185 (I107855,I107838);
nor I_6186 (I107417,I107694,I107855);
nand I_6187 (I107402,I107711,I107855);
nor I_6188 (I107411,I107457,I107838);
DFFARX1 I_6189 (I107838,I2683,I107431,I107420,);
not I_6190 (I107958,I2690);
DFFARX1 I_6191 (I142139,I2683,I107958,I107984,);
nand I_6192 (I107992,I142151,I142130);
and I_6193 (I108009,I107992,I142154);
DFFARX1 I_6194 (I108009,I2683,I107958,I108035,);
nor I_6195 (I107926,I108035,I107984);
not I_6196 (I108057,I108035);
DFFARX1 I_6197 (I142145,I2683,I107958,I108083,);
nand I_6198 (I108091,I108083,I142127);
not I_6199 (I108108,I108091);
DFFARX1 I_6200 (I108108,I2683,I107958,I108134,);
not I_6201 (I107950,I108134);
nor I_6202 (I108156,I107984,I108091);
nor I_6203 (I107932,I108035,I108156);
DFFARX1 I_6204 (I142142,I2683,I107958,I108196,);
DFFARX1 I_6205 (I108196,I2683,I107958,I108213,);
not I_6206 (I108221,I108213);
not I_6207 (I108238,I108196);
nand I_6208 (I107935,I108238,I108057);
nand I_6209 (I108269,I142127,I142133);
and I_6210 (I108286,I108269,I142136);
DFFARX1 I_6211 (I108286,I2683,I107958,I108312,);
nor I_6212 (I108320,I108312,I107984);
DFFARX1 I_6213 (I108320,I2683,I107958,I107923,);
DFFARX1 I_6214 (I108312,I2683,I107958,I107941,);
nor I_6215 (I108365,I142148,I142133);
not I_6216 (I108382,I108365);
nor I_6217 (I107944,I108221,I108382);
nand I_6218 (I107929,I108238,I108382);
nor I_6219 (I107938,I107984,I108365);
DFFARX1 I_6220 (I108365,I2683,I107958,I107947,);
not I_6221 (I108485,I2690);
DFFARX1 I_6222 (I237636,I2683,I108485,I108511,);
nand I_6223 (I108519,I237639,I237633);
and I_6224 (I108536,I108519,I237645);
DFFARX1 I_6225 (I108536,I2683,I108485,I108562,);
nor I_6226 (I108453,I108562,I108511);
not I_6227 (I108584,I108562);
DFFARX1 I_6228 (I237648,I2683,I108485,I108610,);
nand I_6229 (I108618,I108610,I237639);
not I_6230 (I108635,I108618);
DFFARX1 I_6231 (I108635,I2683,I108485,I108661,);
not I_6232 (I108477,I108661);
nor I_6233 (I108683,I108511,I108618);
nor I_6234 (I108459,I108562,I108683);
DFFARX1 I_6235 (I237651,I2683,I108485,I108723,);
DFFARX1 I_6236 (I108723,I2683,I108485,I108740,);
not I_6237 (I108748,I108740);
not I_6238 (I108765,I108723);
nand I_6239 (I108462,I108765,I108584);
nand I_6240 (I108796,I237633,I237642);
and I_6241 (I108813,I108796,I237636);
DFFARX1 I_6242 (I108813,I2683,I108485,I108839,);
nor I_6243 (I108847,I108839,I108511);
DFFARX1 I_6244 (I108847,I2683,I108485,I108450,);
DFFARX1 I_6245 (I108839,I2683,I108485,I108468,);
nor I_6246 (I108892,I237654,I237642);
not I_6247 (I108909,I108892);
nor I_6248 (I108471,I108748,I108909);
nand I_6249 (I108456,I108765,I108909);
nor I_6250 (I108465,I108511,I108892);
DFFARX1 I_6251 (I108892,I2683,I108485,I108474,);
not I_6252 (I109012,I2690);
DFFARX1 I_6253 (I194975,I2683,I109012,I109038,);
nand I_6254 (I109046,I194966,I194981);
and I_6255 (I109063,I109046,I194987);
DFFARX1 I_6256 (I109063,I2683,I109012,I109089,);
nor I_6257 (I108980,I109089,I109038);
not I_6258 (I109111,I109089);
DFFARX1 I_6259 (I194972,I2683,I109012,I109137,);
nand I_6260 (I109145,I109137,I194966);
not I_6261 (I109162,I109145);
DFFARX1 I_6262 (I109162,I2683,I109012,I109188,);
not I_6263 (I109004,I109188);
nor I_6264 (I109210,I109038,I109145);
nor I_6265 (I108986,I109089,I109210);
DFFARX1 I_6266 (I194969,I2683,I109012,I109250,);
DFFARX1 I_6267 (I109250,I2683,I109012,I109267,);
not I_6268 (I109275,I109267);
not I_6269 (I109292,I109250);
nand I_6270 (I108989,I109292,I109111);
nand I_6271 (I109323,I194963,I194978);
and I_6272 (I109340,I109323,I194963);
DFFARX1 I_6273 (I109340,I2683,I109012,I109366,);
nor I_6274 (I109374,I109366,I109038);
DFFARX1 I_6275 (I109374,I2683,I109012,I108977,);
DFFARX1 I_6276 (I109366,I2683,I109012,I108995,);
nor I_6277 (I109419,I194984,I194978);
not I_6278 (I109436,I109419);
nor I_6279 (I108998,I109275,I109436);
nand I_6280 (I108983,I109292,I109436);
nor I_6281 (I108992,I109038,I109419);
DFFARX1 I_6282 (I109419,I2683,I109012,I109001,);
not I_6283 (I109539,I2690);
DFFARX1 I_6284 (I59609,I2683,I109539,I109565,);
nand I_6285 (I109573,I59609,I59615);
and I_6286 (I109590,I109573,I59633);
DFFARX1 I_6287 (I109590,I2683,I109539,I109616,);
nor I_6288 (I109507,I109616,I109565);
not I_6289 (I109638,I109616);
DFFARX1 I_6290 (I59621,I2683,I109539,I109664,);
nand I_6291 (I109672,I109664,I59618);
not I_6292 (I109689,I109672);
DFFARX1 I_6293 (I109689,I2683,I109539,I109715,);
not I_6294 (I109531,I109715);
nor I_6295 (I109737,I109565,I109672);
nor I_6296 (I109513,I109616,I109737);
DFFARX1 I_6297 (I59627,I2683,I109539,I109777,);
DFFARX1 I_6298 (I109777,I2683,I109539,I109794,);
not I_6299 (I109802,I109794);
not I_6300 (I109819,I109777);
nand I_6301 (I109516,I109819,I109638);
nand I_6302 (I109850,I59612,I59612);
and I_6303 (I109867,I109850,I59624);
DFFARX1 I_6304 (I109867,I2683,I109539,I109893,);
nor I_6305 (I109901,I109893,I109565);
DFFARX1 I_6306 (I109901,I2683,I109539,I109504,);
DFFARX1 I_6307 (I109893,I2683,I109539,I109522,);
nor I_6308 (I109946,I59630,I59612);
not I_6309 (I109963,I109946);
nor I_6310 (I109525,I109802,I109963);
nand I_6311 (I109510,I109819,I109963);
nor I_6312 (I109519,I109565,I109946);
DFFARX1 I_6313 (I109946,I2683,I109539,I109528,);
not I_6314 (I110066,I2690);
DFFARX1 I_6315 (I165947,I2683,I110066,I110092,);
nand I_6316 (I110100,I165947,I165959);
and I_6317 (I110117,I110100,I165944);
DFFARX1 I_6318 (I110117,I2683,I110066,I110143,);
nor I_6319 (I110034,I110143,I110092);
not I_6320 (I110165,I110143);
DFFARX1 I_6321 (I165968,I2683,I110066,I110191,);
nand I_6322 (I110199,I110191,I165965);
not I_6323 (I110216,I110199);
DFFARX1 I_6324 (I110216,I2683,I110066,I110242,);
not I_6325 (I110058,I110242);
nor I_6326 (I110264,I110092,I110199);
nor I_6327 (I110040,I110143,I110264);
DFFARX1 I_6328 (I165956,I2683,I110066,I110304,);
DFFARX1 I_6329 (I110304,I2683,I110066,I110321,);
not I_6330 (I110329,I110321);
not I_6331 (I110346,I110304);
nand I_6332 (I110043,I110346,I110165);
nand I_6333 (I110377,I165944,I165953);
and I_6334 (I110394,I110377,I165962);
DFFARX1 I_6335 (I110394,I2683,I110066,I110420,);
nor I_6336 (I110428,I110420,I110092);
DFFARX1 I_6337 (I110428,I2683,I110066,I110031,);
DFFARX1 I_6338 (I110420,I2683,I110066,I110049,);
nor I_6339 (I110473,I165950,I165953);
not I_6340 (I110490,I110473);
nor I_6341 (I110052,I110329,I110490);
nand I_6342 (I110037,I110346,I110490);
nor I_6343 (I110046,I110092,I110473);
DFFARX1 I_6344 (I110473,I2683,I110066,I110055,);
not I_6345 (I110593,I2690);
DFFARX1 I_6346 (I374127,I2683,I110593,I110619,);
nand I_6347 (I110627,I374109,I374133);
and I_6348 (I110644,I110627,I374124);
DFFARX1 I_6349 (I110644,I2683,I110593,I110670,);
nor I_6350 (I110561,I110670,I110619);
not I_6351 (I110692,I110670);
DFFARX1 I_6352 (I374130,I2683,I110593,I110718,);
nand I_6353 (I110726,I110718,I374118);
not I_6354 (I110743,I110726);
DFFARX1 I_6355 (I110743,I2683,I110593,I110769,);
not I_6356 (I110585,I110769);
nor I_6357 (I110791,I110619,I110726);
nor I_6358 (I110567,I110670,I110791);
DFFARX1 I_6359 (I374109,I2683,I110593,I110831,);
DFFARX1 I_6360 (I110831,I2683,I110593,I110848,);
not I_6361 (I110856,I110848);
not I_6362 (I110873,I110831);
nand I_6363 (I110570,I110873,I110692);
nand I_6364 (I110904,I374115,I374112);
and I_6365 (I110921,I110904,I374121);
DFFARX1 I_6366 (I110921,I2683,I110593,I110947,);
nor I_6367 (I110955,I110947,I110619);
DFFARX1 I_6368 (I110955,I2683,I110593,I110558,);
DFFARX1 I_6369 (I110947,I2683,I110593,I110576,);
nor I_6370 (I111000,I374112,I374112);
not I_6371 (I111017,I111000);
nor I_6372 (I110579,I110856,I111017);
nand I_6373 (I110564,I110873,I111017);
nor I_6374 (I110573,I110619,I111000);
DFFARX1 I_6375 (I111000,I2683,I110593,I110582,);
not I_6376 (I111120,I2690);
DFFARX1 I_6377 (I208269,I2683,I111120,I111146,);
nand I_6378 (I111154,I208260,I208275);
and I_6379 (I111171,I111154,I208281);
DFFARX1 I_6380 (I111171,I2683,I111120,I111197,);
nor I_6381 (I111088,I111197,I111146);
not I_6382 (I111219,I111197);
DFFARX1 I_6383 (I208266,I2683,I111120,I111245,);
nand I_6384 (I111253,I111245,I208260);
not I_6385 (I111270,I111253);
DFFARX1 I_6386 (I111270,I2683,I111120,I111296,);
not I_6387 (I111112,I111296);
nor I_6388 (I111318,I111146,I111253);
nor I_6389 (I111094,I111197,I111318);
DFFARX1 I_6390 (I208263,I2683,I111120,I111358,);
DFFARX1 I_6391 (I111358,I2683,I111120,I111375,);
not I_6392 (I111383,I111375);
not I_6393 (I111400,I111358);
nand I_6394 (I111097,I111400,I111219);
nand I_6395 (I111431,I208257,I208272);
and I_6396 (I111448,I111431,I208257);
DFFARX1 I_6397 (I111448,I2683,I111120,I111474,);
nor I_6398 (I111482,I111474,I111146);
DFFARX1 I_6399 (I111482,I2683,I111120,I111085,);
DFFARX1 I_6400 (I111474,I2683,I111120,I111103,);
nor I_6401 (I111527,I208278,I208272);
not I_6402 (I111544,I111527);
nor I_6403 (I111106,I111383,I111544);
nand I_6404 (I111091,I111400,I111544);
nor I_6405 (I111100,I111146,I111527);
DFFARX1 I_6406 (I111527,I2683,I111120,I111109,);
not I_6407 (I111647,I2690);
DFFARX1 I_6408 (I226187,I2683,I111647,I111673,);
nand I_6409 (I111681,I226178,I226193);
and I_6410 (I111698,I111681,I226199);
DFFARX1 I_6411 (I111698,I2683,I111647,I111724,);
nor I_6412 (I111615,I111724,I111673);
not I_6413 (I111746,I111724);
DFFARX1 I_6414 (I226184,I2683,I111647,I111772,);
nand I_6415 (I111780,I111772,I226178);
not I_6416 (I111797,I111780);
DFFARX1 I_6417 (I111797,I2683,I111647,I111823,);
not I_6418 (I111639,I111823);
nor I_6419 (I111845,I111673,I111780);
nor I_6420 (I111621,I111724,I111845);
DFFARX1 I_6421 (I226181,I2683,I111647,I111885,);
DFFARX1 I_6422 (I111885,I2683,I111647,I111902,);
not I_6423 (I111910,I111902);
not I_6424 (I111927,I111885);
nand I_6425 (I111624,I111927,I111746);
nand I_6426 (I111958,I226175,I226190);
and I_6427 (I111975,I111958,I226175);
DFFARX1 I_6428 (I111975,I2683,I111647,I112001,);
nor I_6429 (I112009,I112001,I111673);
DFFARX1 I_6430 (I112009,I2683,I111647,I111612,);
DFFARX1 I_6431 (I112001,I2683,I111647,I111630,);
nor I_6432 (I112054,I226196,I226190);
not I_6433 (I112071,I112054);
nor I_6434 (I111633,I111910,I112071);
nand I_6435 (I111618,I111927,I112071);
nor I_6436 (I111627,I111673,I112054);
DFFARX1 I_6437 (I112054,I2683,I111647,I111636,);
not I_6438 (I112174,I2690);
DFFARX1 I_6439 (I316567,I2683,I112174,I112200,);
nand I_6440 (I112208,I316564,I316567);
and I_6441 (I112225,I112208,I316576);
DFFARX1 I_6442 (I112225,I2683,I112174,I112251,);
nor I_6443 (I112142,I112251,I112200);
not I_6444 (I112273,I112251);
DFFARX1 I_6445 (I316564,I2683,I112174,I112299,);
nand I_6446 (I112307,I112299,I316582);
not I_6447 (I112324,I112307);
DFFARX1 I_6448 (I112324,I2683,I112174,I112350,);
not I_6449 (I112166,I112350);
nor I_6450 (I112372,I112200,I112307);
nor I_6451 (I112148,I112251,I112372);
DFFARX1 I_6452 (I316570,I2683,I112174,I112412,);
DFFARX1 I_6453 (I112412,I2683,I112174,I112429,);
not I_6454 (I112437,I112429);
not I_6455 (I112454,I112412);
nand I_6456 (I112151,I112454,I112273);
nand I_6457 (I112485,I316579,I316585);
and I_6458 (I112502,I112485,I316570);
DFFARX1 I_6459 (I112502,I2683,I112174,I112528,);
nor I_6460 (I112536,I112528,I112200);
DFFARX1 I_6461 (I112536,I2683,I112174,I112139,);
DFFARX1 I_6462 (I112528,I2683,I112174,I112157,);
nor I_6463 (I112581,I316573,I316585);
not I_6464 (I112598,I112581);
nor I_6465 (I112160,I112437,I112598);
nand I_6466 (I112145,I112454,I112598);
nor I_6467 (I112154,I112200,I112581);
DFFARX1 I_6468 (I112581,I2683,I112174,I112163,);
not I_6469 (I112701,I2690);
DFFARX1 I_6470 (I167732,I2683,I112701,I112727,);
nand I_6471 (I112735,I167732,I167744);
and I_6472 (I112752,I112735,I167729);
DFFARX1 I_6473 (I112752,I2683,I112701,I112778,);
nor I_6474 (I112669,I112778,I112727);
not I_6475 (I112800,I112778);
DFFARX1 I_6476 (I167753,I2683,I112701,I112826,);
nand I_6477 (I112834,I112826,I167750);
not I_6478 (I112851,I112834);
DFFARX1 I_6479 (I112851,I2683,I112701,I112877,);
not I_6480 (I112693,I112877);
nor I_6481 (I112899,I112727,I112834);
nor I_6482 (I112675,I112778,I112899);
DFFARX1 I_6483 (I167741,I2683,I112701,I112939,);
DFFARX1 I_6484 (I112939,I2683,I112701,I112956,);
not I_6485 (I112964,I112956);
not I_6486 (I112981,I112939);
nand I_6487 (I112678,I112981,I112800);
nand I_6488 (I113012,I167729,I167738);
and I_6489 (I113029,I113012,I167747);
DFFARX1 I_6490 (I113029,I2683,I112701,I113055,);
nor I_6491 (I113063,I113055,I112727);
DFFARX1 I_6492 (I113063,I2683,I112701,I112666,);
DFFARX1 I_6493 (I113055,I2683,I112701,I112684,);
nor I_6494 (I113108,I167735,I167738);
not I_6495 (I113125,I113108);
nor I_6496 (I112687,I112964,I113125);
nand I_6497 (I112672,I112981,I113125);
nor I_6498 (I112681,I112727,I113108);
DFFARX1 I_6499 (I113108,I2683,I112701,I112690,);
not I_6500 (I113228,I2690);
DFFARX1 I_6501 (I1636,I2683,I113228,I113254,);
nand I_6502 (I113262,I2588,I1908);
and I_6503 (I113279,I113262,I1604);
DFFARX1 I_6504 (I113279,I2683,I113228,I113305,);
nor I_6505 (I113196,I113305,I113254);
not I_6506 (I113327,I113305);
DFFARX1 I_6507 (I2316,I2683,I113228,I113353,);
nand I_6508 (I113361,I113353,I1420);
not I_6509 (I113378,I113361);
DFFARX1 I_6510 (I113378,I2683,I113228,I113404,);
not I_6511 (I113220,I113404);
nor I_6512 (I113426,I113254,I113361);
nor I_6513 (I113202,I113305,I113426);
DFFARX1 I_6514 (I2468,I2683,I113228,I113466,);
DFFARX1 I_6515 (I113466,I2683,I113228,I113483,);
not I_6516 (I113491,I113483);
not I_6517 (I113508,I113466);
nand I_6518 (I113205,I113508,I113327);
nand I_6519 (I113539,I2444,I1516);
and I_6520 (I113556,I113539,I1980);
DFFARX1 I_6521 (I113556,I2683,I113228,I113582,);
nor I_6522 (I113590,I113582,I113254);
DFFARX1 I_6523 (I113590,I2683,I113228,I113193,);
DFFARX1 I_6524 (I113582,I2683,I113228,I113211,);
nor I_6525 (I113635,I1412,I1516);
not I_6526 (I113652,I113635);
nor I_6527 (I113214,I113491,I113652);
nand I_6528 (I113199,I113508,I113652);
nor I_6529 (I113208,I113254,I113635);
DFFARX1 I_6530 (I113635,I2683,I113228,I113217,);
not I_6531 (I113755,I2690);
DFFARX1 I_6532 (I231389,I2683,I113755,I113781,);
nand I_6533 (I113789,I231380,I231395);
and I_6534 (I113806,I113789,I231401);
DFFARX1 I_6535 (I113806,I2683,I113755,I113832,);
nor I_6536 (I113723,I113832,I113781);
not I_6537 (I113854,I113832);
DFFARX1 I_6538 (I231386,I2683,I113755,I113880,);
nand I_6539 (I113888,I113880,I231380);
not I_6540 (I113905,I113888);
DFFARX1 I_6541 (I113905,I2683,I113755,I113931,);
not I_6542 (I113747,I113931);
nor I_6543 (I113953,I113781,I113888);
nor I_6544 (I113729,I113832,I113953);
DFFARX1 I_6545 (I231383,I2683,I113755,I113993,);
DFFARX1 I_6546 (I113993,I2683,I113755,I114010,);
not I_6547 (I114018,I114010);
not I_6548 (I114035,I113993);
nand I_6549 (I113732,I114035,I113854);
nand I_6550 (I114066,I231377,I231392);
and I_6551 (I114083,I114066,I231377);
DFFARX1 I_6552 (I114083,I2683,I113755,I114109,);
nor I_6553 (I114117,I114109,I113781);
DFFARX1 I_6554 (I114117,I2683,I113755,I113720,);
DFFARX1 I_6555 (I114109,I2683,I113755,I113738,);
nor I_6556 (I114162,I231398,I231392);
not I_6557 (I114179,I114162);
nor I_6558 (I113741,I114018,I114179);
nand I_6559 (I113726,I114035,I114179);
nor I_6560 (I113735,I113781,I114162);
DFFARX1 I_6561 (I114162,I2683,I113755,I113744,);
not I_6562 (I114282,I2690);
DFFARX1 I_6563 (I200755,I2683,I114282,I114308,);
nand I_6564 (I114316,I200746,I200761);
and I_6565 (I114333,I114316,I200767);
DFFARX1 I_6566 (I114333,I2683,I114282,I114359,);
nor I_6567 (I114250,I114359,I114308);
not I_6568 (I114381,I114359);
DFFARX1 I_6569 (I200752,I2683,I114282,I114407,);
nand I_6570 (I114415,I114407,I200746);
not I_6571 (I114432,I114415);
DFFARX1 I_6572 (I114432,I2683,I114282,I114458,);
not I_6573 (I114274,I114458);
nor I_6574 (I114480,I114308,I114415);
nor I_6575 (I114256,I114359,I114480);
DFFARX1 I_6576 (I200749,I2683,I114282,I114520,);
DFFARX1 I_6577 (I114520,I2683,I114282,I114537,);
not I_6578 (I114545,I114537);
not I_6579 (I114562,I114520);
nand I_6580 (I114259,I114562,I114381);
nand I_6581 (I114593,I200743,I200758);
and I_6582 (I114610,I114593,I200743);
DFFARX1 I_6583 (I114610,I2683,I114282,I114636,);
nor I_6584 (I114644,I114636,I114308);
DFFARX1 I_6585 (I114644,I2683,I114282,I114247,);
DFFARX1 I_6586 (I114636,I2683,I114282,I114265,);
nor I_6587 (I114689,I200764,I200758);
not I_6588 (I114706,I114689);
nor I_6589 (I114268,I114545,I114706);
nand I_6590 (I114253,I114562,I114706);
nor I_6591 (I114262,I114308,I114689);
DFFARX1 I_6592 (I114689,I2683,I114282,I114271,);
not I_6593 (I114809,I2690);
DFFARX1 I_6594 (I362005,I2683,I114809,I114835,);
nand I_6595 (I114843,I362020,I362005);
and I_6596 (I114860,I114843,I362023);
DFFARX1 I_6597 (I114860,I2683,I114809,I114886,);
nor I_6598 (I114777,I114886,I114835);
not I_6599 (I114908,I114886);
DFFARX1 I_6600 (I362029,I2683,I114809,I114934,);
nand I_6601 (I114942,I114934,I362011);
not I_6602 (I114959,I114942);
DFFARX1 I_6603 (I114959,I2683,I114809,I114985,);
not I_6604 (I114801,I114985);
nor I_6605 (I115007,I114835,I114942);
nor I_6606 (I114783,I114886,I115007);
DFFARX1 I_6607 (I362008,I2683,I114809,I115047,);
DFFARX1 I_6608 (I115047,I2683,I114809,I115064,);
not I_6609 (I115072,I115064);
not I_6610 (I115089,I115047);
nand I_6611 (I114786,I115089,I114908);
nand I_6612 (I115120,I362008,I362014);
and I_6613 (I115137,I115120,I362026);
DFFARX1 I_6614 (I115137,I2683,I114809,I115163,);
nor I_6615 (I115171,I115163,I114835);
DFFARX1 I_6616 (I115171,I2683,I114809,I114774,);
DFFARX1 I_6617 (I115163,I2683,I114809,I114792,);
nor I_6618 (I115216,I362017,I362014);
not I_6619 (I115233,I115216);
nor I_6620 (I114795,I115072,I115233);
nand I_6621 (I114780,I115089,I115233);
nor I_6622 (I114789,I114835,I115216);
DFFARX1 I_6623 (I115216,I2683,I114809,I114798,);
not I_6624 (I115336,I2690);
DFFARX1 I_6625 (I281411,I2683,I115336,I115362,);
nand I_6626 (I115370,I281408,I281426);
and I_6627 (I115387,I115370,I281417);
DFFARX1 I_6628 (I115387,I2683,I115336,I115413,);
nor I_6629 (I115304,I115413,I115362);
not I_6630 (I115435,I115413);
DFFARX1 I_6631 (I281432,I2683,I115336,I115461,);
nand I_6632 (I115469,I115461,I281414);
not I_6633 (I115486,I115469);
DFFARX1 I_6634 (I115486,I2683,I115336,I115512,);
not I_6635 (I115328,I115512);
nor I_6636 (I115534,I115362,I115469);
nor I_6637 (I115310,I115413,I115534);
DFFARX1 I_6638 (I281420,I2683,I115336,I115574,);
DFFARX1 I_6639 (I115574,I2683,I115336,I115591,);
not I_6640 (I115599,I115591);
not I_6641 (I115616,I115574);
nand I_6642 (I115313,I115616,I115435);
nand I_6643 (I115647,I281408,I281435);
and I_6644 (I115664,I115647,I281423);
DFFARX1 I_6645 (I115664,I2683,I115336,I115690,);
nor I_6646 (I115698,I115690,I115362);
DFFARX1 I_6647 (I115698,I2683,I115336,I115301,);
DFFARX1 I_6648 (I115690,I2683,I115336,I115319,);
nor I_6649 (I115743,I281429,I281435);
not I_6650 (I115760,I115743);
nor I_6651 (I115322,I115599,I115760);
nand I_6652 (I115307,I115616,I115760);
nor I_6653 (I115316,I115362,I115743);
DFFARX1 I_6654 (I115743,I2683,I115336,I115325,);
not I_6655 (I115863,I2690);
DFFARX1 I_6656 (I385956,I2683,I115863,I115889,);
nand I_6657 (I115897,I385953,I385944);
and I_6658 (I115914,I115897,I385941);
DFFARX1 I_6659 (I115914,I2683,I115863,I115940,);
nor I_6660 (I115831,I115940,I115889);
not I_6661 (I115962,I115940);
DFFARX1 I_6662 (I385950,I2683,I115863,I115988,);
nand I_6663 (I115996,I115988,I385959);
not I_6664 (I116013,I115996);
DFFARX1 I_6665 (I116013,I2683,I115863,I116039,);
not I_6666 (I115855,I116039);
nor I_6667 (I116061,I115889,I115996);
nor I_6668 (I115837,I115940,I116061);
DFFARX1 I_6669 (I385962,I2683,I115863,I116101,);
DFFARX1 I_6670 (I116101,I2683,I115863,I116118,);
not I_6671 (I116126,I116118);
not I_6672 (I116143,I116101);
nand I_6673 (I115840,I116143,I115962);
nand I_6674 (I116174,I385941,I385947);
and I_6675 (I116191,I116174,I385965);
DFFARX1 I_6676 (I116191,I2683,I115863,I116217,);
nor I_6677 (I116225,I116217,I115889);
DFFARX1 I_6678 (I116225,I2683,I115863,I115828,);
DFFARX1 I_6679 (I116217,I2683,I115863,I115846,);
nor I_6680 (I116270,I385944,I385947);
not I_6681 (I116287,I116270);
nor I_6682 (I115849,I116126,I116287);
nand I_6683 (I115834,I116143,I116287);
nor I_6684 (I115843,I115889,I116270);
DFFARX1 I_6685 (I116270,I2683,I115863,I115852,);
not I_6686 (I116390,I2690);
DFFARX1 I_6687 (I376303,I2683,I116390,I116416,);
nand I_6688 (I116424,I376285,I376309);
and I_6689 (I116441,I116424,I376300);
DFFARX1 I_6690 (I116441,I2683,I116390,I116467,);
nor I_6691 (I116358,I116467,I116416);
not I_6692 (I116489,I116467);
DFFARX1 I_6693 (I376306,I2683,I116390,I116515,);
nand I_6694 (I116523,I116515,I376294);
not I_6695 (I116540,I116523);
DFFARX1 I_6696 (I116540,I2683,I116390,I116566,);
not I_6697 (I116382,I116566);
nor I_6698 (I116588,I116416,I116523);
nor I_6699 (I116364,I116467,I116588);
DFFARX1 I_6700 (I376285,I2683,I116390,I116628,);
DFFARX1 I_6701 (I116628,I2683,I116390,I116645,);
not I_6702 (I116653,I116645);
not I_6703 (I116670,I116628);
nand I_6704 (I116367,I116670,I116489);
nand I_6705 (I116701,I376291,I376288);
and I_6706 (I116718,I116701,I376297);
DFFARX1 I_6707 (I116718,I2683,I116390,I116744,);
nor I_6708 (I116752,I116744,I116416);
DFFARX1 I_6709 (I116752,I2683,I116390,I116355,);
DFFARX1 I_6710 (I116744,I2683,I116390,I116373,);
nor I_6711 (I116797,I376288,I376288);
not I_6712 (I116814,I116797);
nor I_6713 (I116376,I116653,I116814);
nand I_6714 (I116361,I116670,I116814);
nor I_6715 (I116370,I116416,I116797);
DFFARX1 I_6716 (I116797,I2683,I116390,I116379,);
not I_6717 (I116917,I2690);
DFFARX1 I_6718 (I149755,I2683,I116917,I116943,);
nand I_6719 (I116951,I149767,I149746);
and I_6720 (I116968,I116951,I149770);
DFFARX1 I_6721 (I116968,I2683,I116917,I116994,);
nor I_6722 (I116885,I116994,I116943);
not I_6723 (I117016,I116994);
DFFARX1 I_6724 (I149761,I2683,I116917,I117042,);
nand I_6725 (I117050,I117042,I149743);
not I_6726 (I117067,I117050);
DFFARX1 I_6727 (I117067,I2683,I116917,I117093,);
not I_6728 (I116909,I117093);
nor I_6729 (I117115,I116943,I117050);
nor I_6730 (I116891,I116994,I117115);
DFFARX1 I_6731 (I149758,I2683,I116917,I117155,);
DFFARX1 I_6732 (I117155,I2683,I116917,I117172,);
not I_6733 (I117180,I117172);
not I_6734 (I117197,I117155);
nand I_6735 (I116894,I117197,I117016);
nand I_6736 (I117228,I149743,I149749);
and I_6737 (I117245,I117228,I149752);
DFFARX1 I_6738 (I117245,I2683,I116917,I117271,);
nor I_6739 (I117279,I117271,I116943);
DFFARX1 I_6740 (I117279,I2683,I116917,I116882,);
DFFARX1 I_6741 (I117271,I2683,I116917,I116900,);
nor I_6742 (I117324,I149764,I149749);
not I_6743 (I117341,I117324);
nor I_6744 (I116903,I117180,I117341);
nand I_6745 (I116888,I117197,I117341);
nor I_6746 (I116897,I116943,I117324);
DFFARX1 I_6747 (I117324,I2683,I116917,I116906,);
not I_6748 (I117444,I2690);
DFFARX1 I_6749 (I203067,I2683,I117444,I117470,);
nand I_6750 (I117478,I203058,I203073);
and I_6751 (I117495,I117478,I203079);
DFFARX1 I_6752 (I117495,I2683,I117444,I117521,);
nor I_6753 (I117412,I117521,I117470);
not I_6754 (I117543,I117521);
DFFARX1 I_6755 (I203064,I2683,I117444,I117569,);
nand I_6756 (I117577,I117569,I203058);
not I_6757 (I117594,I117577);
DFFARX1 I_6758 (I117594,I2683,I117444,I117620,);
not I_6759 (I117436,I117620);
nor I_6760 (I117642,I117470,I117577);
nor I_6761 (I117418,I117521,I117642);
DFFARX1 I_6762 (I203061,I2683,I117444,I117682,);
DFFARX1 I_6763 (I117682,I2683,I117444,I117699,);
not I_6764 (I117707,I117699);
not I_6765 (I117724,I117682);
nand I_6766 (I117421,I117724,I117543);
nand I_6767 (I117755,I203055,I203070);
and I_6768 (I117772,I117755,I203055);
DFFARX1 I_6769 (I117772,I2683,I117444,I117798,);
nor I_6770 (I117806,I117798,I117470);
DFFARX1 I_6771 (I117806,I2683,I117444,I117409,);
DFFARX1 I_6772 (I117798,I2683,I117444,I117427,);
nor I_6773 (I117851,I203076,I203070);
not I_6774 (I117868,I117851);
nor I_6775 (I117430,I117707,I117868);
nand I_6776 (I117415,I117724,I117868);
nor I_6777 (I117424,I117470,I117851);
DFFARX1 I_6778 (I117851,I2683,I117444,I117433,);
not I_6779 (I117971,I2690);
DFFARX1 I_6780 (I52469,I2683,I117971,I117997,);
nand I_6781 (I118005,I52469,I52475);
and I_6782 (I118022,I118005,I52493);
DFFARX1 I_6783 (I118022,I2683,I117971,I118048,);
nor I_6784 (I117939,I118048,I117997);
not I_6785 (I118070,I118048);
DFFARX1 I_6786 (I52481,I2683,I117971,I118096,);
nand I_6787 (I118104,I118096,I52478);
not I_6788 (I118121,I118104);
DFFARX1 I_6789 (I118121,I2683,I117971,I118147,);
not I_6790 (I117963,I118147);
nor I_6791 (I118169,I117997,I118104);
nor I_6792 (I117945,I118048,I118169);
DFFARX1 I_6793 (I52487,I2683,I117971,I118209,);
DFFARX1 I_6794 (I118209,I2683,I117971,I118226,);
not I_6795 (I118234,I118226);
not I_6796 (I118251,I118209);
nand I_6797 (I117948,I118251,I118070);
nand I_6798 (I118282,I52472,I52472);
and I_6799 (I118299,I118282,I52484);
DFFARX1 I_6800 (I118299,I2683,I117971,I118325,);
nor I_6801 (I118333,I118325,I117997);
DFFARX1 I_6802 (I118333,I2683,I117971,I117936,);
DFFARX1 I_6803 (I118325,I2683,I117971,I117954,);
nor I_6804 (I118378,I52490,I52472);
not I_6805 (I118395,I118378);
nor I_6806 (I117957,I118234,I118395);
nand I_6807 (I117942,I118251,I118395);
nor I_6808 (I117951,I117997,I118378);
DFFARX1 I_6809 (I118378,I2683,I117971,I117960,);
not I_6810 (I118498,I2690);
DFFARX1 I_6811 (I131259,I2683,I118498,I118524,);
nand I_6812 (I118532,I131271,I131250);
and I_6813 (I118549,I118532,I131274);
DFFARX1 I_6814 (I118549,I2683,I118498,I118575,);
nor I_6815 (I118466,I118575,I118524);
not I_6816 (I118597,I118575);
DFFARX1 I_6817 (I131265,I2683,I118498,I118623,);
nand I_6818 (I118631,I118623,I131247);
not I_6819 (I118648,I118631);
DFFARX1 I_6820 (I118648,I2683,I118498,I118674,);
not I_6821 (I118490,I118674);
nor I_6822 (I118696,I118524,I118631);
nor I_6823 (I118472,I118575,I118696);
DFFARX1 I_6824 (I131262,I2683,I118498,I118736,);
DFFARX1 I_6825 (I118736,I2683,I118498,I118753,);
not I_6826 (I118761,I118753);
not I_6827 (I118778,I118736);
nand I_6828 (I118475,I118778,I118597);
nand I_6829 (I118809,I131247,I131253);
and I_6830 (I118826,I118809,I131256);
DFFARX1 I_6831 (I118826,I2683,I118498,I118852,);
nor I_6832 (I118860,I118852,I118524);
DFFARX1 I_6833 (I118860,I2683,I118498,I118463,);
DFFARX1 I_6834 (I118852,I2683,I118498,I118481,);
nor I_6835 (I118905,I131268,I131253);
not I_6836 (I118922,I118905);
nor I_6837 (I118484,I118761,I118922);
nand I_6838 (I118469,I118778,I118922);
nor I_6839 (I118478,I118524,I118905);
DFFARX1 I_6840 (I118905,I2683,I118498,I118487,);
not I_6841 (I119025,I2690);
DFFARX1 I_6842 (I34129,I2683,I119025,I119051,);
nand I_6843 (I119059,I34141,I34150);
and I_6844 (I119076,I119059,I34129);
DFFARX1 I_6845 (I119076,I2683,I119025,I119102,);
nor I_6846 (I118993,I119102,I119051);
not I_6847 (I119124,I119102);
DFFARX1 I_6848 (I34144,I2683,I119025,I119150,);
nand I_6849 (I119158,I119150,I34132);
not I_6850 (I119175,I119158);
DFFARX1 I_6851 (I119175,I2683,I119025,I119201,);
not I_6852 (I119017,I119201);
nor I_6853 (I119223,I119051,I119158);
nor I_6854 (I118999,I119102,I119223);
DFFARX1 I_6855 (I34135,I2683,I119025,I119263,);
DFFARX1 I_6856 (I119263,I2683,I119025,I119280,);
not I_6857 (I119288,I119280);
not I_6858 (I119305,I119263);
nand I_6859 (I119002,I119305,I119124);
nand I_6860 (I119336,I34126,I34126);
and I_6861 (I119353,I119336,I34138);
DFFARX1 I_6862 (I119353,I2683,I119025,I119379,);
nor I_6863 (I119387,I119379,I119051);
DFFARX1 I_6864 (I119387,I2683,I119025,I118990,);
DFFARX1 I_6865 (I119379,I2683,I119025,I119008,);
nor I_6866 (I119432,I34147,I34126);
not I_6867 (I119449,I119432);
nor I_6868 (I119011,I119288,I119449);
nand I_6869 (I118996,I119305,I119449);
nor I_6870 (I119005,I119051,I119432);
DFFARX1 I_6871 (I119432,I2683,I119025,I119014,);
not I_6872 (I119552,I2690);
DFFARX1 I_6873 (I321055,I2683,I119552,I119578,);
nand I_6874 (I119586,I321052,I321055);
and I_6875 (I119603,I119586,I321064);
DFFARX1 I_6876 (I119603,I2683,I119552,I119629,);
nor I_6877 (I119520,I119629,I119578);
not I_6878 (I119651,I119629);
DFFARX1 I_6879 (I321052,I2683,I119552,I119677,);
nand I_6880 (I119685,I119677,I321070);
not I_6881 (I119702,I119685);
DFFARX1 I_6882 (I119702,I2683,I119552,I119728,);
not I_6883 (I119544,I119728);
nor I_6884 (I119750,I119578,I119685);
nor I_6885 (I119526,I119629,I119750);
DFFARX1 I_6886 (I321058,I2683,I119552,I119790,);
DFFARX1 I_6887 (I119790,I2683,I119552,I119807,);
not I_6888 (I119815,I119807);
not I_6889 (I119832,I119790);
nand I_6890 (I119529,I119832,I119651);
nand I_6891 (I119863,I321067,I321073);
and I_6892 (I119880,I119863,I321058);
DFFARX1 I_6893 (I119880,I2683,I119552,I119906,);
nor I_6894 (I119914,I119906,I119578);
DFFARX1 I_6895 (I119914,I2683,I119552,I119517,);
DFFARX1 I_6896 (I119906,I2683,I119552,I119535,);
nor I_6897 (I119959,I321061,I321073);
not I_6898 (I119976,I119959);
nor I_6899 (I119538,I119815,I119976);
nand I_6900 (I119523,I119832,I119976);
nor I_6901 (I119532,I119578,I119959);
DFFARX1 I_6902 (I119959,I2683,I119552,I119541,);
not I_6903 (I120079,I2690);
DFFARX1 I_6904 (I322738,I2683,I120079,I120105,);
nand I_6905 (I120113,I322735,I322738);
and I_6906 (I120130,I120113,I322747);
DFFARX1 I_6907 (I120130,I2683,I120079,I120156,);
nor I_6908 (I120047,I120156,I120105);
not I_6909 (I120178,I120156);
DFFARX1 I_6910 (I322735,I2683,I120079,I120204,);
nand I_6911 (I120212,I120204,I322753);
not I_6912 (I120229,I120212);
DFFARX1 I_6913 (I120229,I2683,I120079,I120255,);
not I_6914 (I120071,I120255);
nor I_6915 (I120277,I120105,I120212);
nor I_6916 (I120053,I120156,I120277);
DFFARX1 I_6917 (I322741,I2683,I120079,I120317,);
DFFARX1 I_6918 (I120317,I2683,I120079,I120334,);
not I_6919 (I120342,I120334);
not I_6920 (I120359,I120317);
nand I_6921 (I120056,I120359,I120178);
nand I_6922 (I120390,I322750,I322756);
and I_6923 (I120407,I120390,I322741);
DFFARX1 I_6924 (I120407,I2683,I120079,I120433,);
nor I_6925 (I120441,I120433,I120105);
DFFARX1 I_6926 (I120441,I2683,I120079,I120044,);
DFFARX1 I_6927 (I120433,I2683,I120079,I120062,);
nor I_6928 (I120486,I322744,I322756);
not I_6929 (I120503,I120486);
nor I_6930 (I120065,I120342,I120503);
nand I_6931 (I120050,I120359,I120503);
nor I_6932 (I120059,I120105,I120486);
DFFARX1 I_6933 (I120486,I2683,I120079,I120068,);
not I_6934 (I120606,I2690);
DFFARX1 I_6935 (I48899,I2683,I120606,I120632,);
nand I_6936 (I120640,I48899,I48905);
and I_6937 (I120657,I120640,I48923);
DFFARX1 I_6938 (I120657,I2683,I120606,I120683,);
nor I_6939 (I120574,I120683,I120632);
not I_6940 (I120705,I120683);
DFFARX1 I_6941 (I48911,I2683,I120606,I120731,);
nand I_6942 (I120739,I120731,I48908);
not I_6943 (I120756,I120739);
DFFARX1 I_6944 (I120756,I2683,I120606,I120782,);
not I_6945 (I120598,I120782);
nor I_6946 (I120804,I120632,I120739);
nor I_6947 (I120580,I120683,I120804);
DFFARX1 I_6948 (I48917,I2683,I120606,I120844,);
DFFARX1 I_6949 (I120844,I2683,I120606,I120861,);
not I_6950 (I120869,I120861);
not I_6951 (I120886,I120844);
nand I_6952 (I120583,I120886,I120705);
nand I_6953 (I120917,I48902,I48902);
and I_6954 (I120934,I120917,I48914);
DFFARX1 I_6955 (I120934,I2683,I120606,I120960,);
nor I_6956 (I120968,I120960,I120632);
DFFARX1 I_6957 (I120968,I2683,I120606,I120571,);
DFFARX1 I_6958 (I120960,I2683,I120606,I120589,);
nor I_6959 (I121013,I48920,I48902);
not I_6960 (I121030,I121013);
nor I_6961 (I120592,I120869,I121030);
nand I_6962 (I120577,I120886,I121030);
nor I_6963 (I120586,I120632,I121013);
DFFARX1 I_6964 (I121013,I2683,I120606,I120595,);
not I_6965 (I121133,I2690);
DFFARX1 I_6966 (I188042,I2683,I121133,I121159,);
nand I_6967 (I121167,I188027,I188030);
and I_6968 (I121184,I121167,I188045);
DFFARX1 I_6969 (I121184,I2683,I121133,I121210,);
nor I_6970 (I121101,I121210,I121159);
not I_6971 (I121232,I121210);
DFFARX1 I_6972 (I188039,I2683,I121133,I121258,);
nand I_6973 (I121266,I121258,I188030);
not I_6974 (I121283,I121266);
DFFARX1 I_6975 (I121283,I2683,I121133,I121309,);
not I_6976 (I121125,I121309);
nor I_6977 (I121331,I121159,I121266);
nor I_6978 (I121107,I121210,I121331);
DFFARX1 I_6979 (I188036,I2683,I121133,I121371,);
DFFARX1 I_6980 (I121371,I2683,I121133,I121388,);
not I_6981 (I121396,I121388);
not I_6982 (I121413,I121371);
nand I_6983 (I121110,I121413,I121232);
nand I_6984 (I121444,I188051,I188027);
and I_6985 (I121461,I121444,I188048);
DFFARX1 I_6986 (I121461,I2683,I121133,I121487,);
nor I_6987 (I121495,I121487,I121159);
DFFARX1 I_6988 (I121495,I2683,I121133,I121098,);
DFFARX1 I_6989 (I121487,I2683,I121133,I121116,);
nor I_6990 (I121540,I188033,I188027);
not I_6991 (I121557,I121540);
nor I_6992 (I121119,I121396,I121557);
nand I_6993 (I121104,I121413,I121557);
nor I_6994 (I121113,I121159,I121540);
DFFARX1 I_6995 (I121540,I2683,I121133,I121122,);
not I_6996 (I121660,I2690);
DFFARX1 I_6997 (I351023,I2683,I121660,I121686,);
nand I_6998 (I121694,I351038,I351023);
and I_6999 (I121711,I121694,I351041);
DFFARX1 I_7000 (I121711,I2683,I121660,I121737,);
nor I_7001 (I121628,I121737,I121686);
not I_7002 (I121759,I121737);
DFFARX1 I_7003 (I351047,I2683,I121660,I121785,);
nand I_7004 (I121793,I121785,I351029);
not I_7005 (I121810,I121793);
DFFARX1 I_7006 (I121810,I2683,I121660,I121836,);
not I_7007 (I121652,I121836);
nor I_7008 (I121858,I121686,I121793);
nor I_7009 (I121634,I121737,I121858);
DFFARX1 I_7010 (I351026,I2683,I121660,I121898,);
DFFARX1 I_7011 (I121898,I2683,I121660,I121915,);
not I_7012 (I121923,I121915);
not I_7013 (I121940,I121898);
nand I_7014 (I121637,I121940,I121759);
nand I_7015 (I121971,I351026,I351032);
and I_7016 (I121988,I121971,I351044);
DFFARX1 I_7017 (I121988,I2683,I121660,I122014,);
nor I_7018 (I122022,I122014,I121686);
DFFARX1 I_7019 (I122022,I2683,I121660,I121625,);
DFFARX1 I_7020 (I122014,I2683,I121660,I121643,);
nor I_7021 (I122067,I351035,I351032);
not I_7022 (I122084,I122067);
nor I_7023 (I121646,I121923,I122084);
nand I_7024 (I121631,I121940,I122084);
nor I_7025 (I121640,I121686,I122067);
DFFARX1 I_7026 (I122067,I2683,I121660,I121649,);
not I_7027 (I122187,I2690);
DFFARX1 I_7028 (I184574,I2683,I122187,I122213,);
nand I_7029 (I122221,I184559,I184562);
and I_7030 (I122238,I122221,I184577);
DFFARX1 I_7031 (I122238,I2683,I122187,I122264,);
nor I_7032 (I122155,I122264,I122213);
not I_7033 (I122286,I122264);
DFFARX1 I_7034 (I184571,I2683,I122187,I122312,);
nand I_7035 (I122320,I122312,I184562);
not I_7036 (I122337,I122320);
DFFARX1 I_7037 (I122337,I2683,I122187,I122363,);
not I_7038 (I122179,I122363);
nor I_7039 (I122385,I122213,I122320);
nor I_7040 (I122161,I122264,I122385);
DFFARX1 I_7041 (I184568,I2683,I122187,I122425,);
DFFARX1 I_7042 (I122425,I2683,I122187,I122442,);
not I_7043 (I122450,I122442);
not I_7044 (I122467,I122425);
nand I_7045 (I122164,I122467,I122286);
nand I_7046 (I122498,I184583,I184559);
and I_7047 (I122515,I122498,I184580);
DFFARX1 I_7048 (I122515,I2683,I122187,I122541,);
nor I_7049 (I122549,I122541,I122213);
DFFARX1 I_7050 (I122549,I2683,I122187,I122152,);
DFFARX1 I_7051 (I122541,I2683,I122187,I122170,);
nor I_7052 (I122594,I184565,I184559);
not I_7053 (I122611,I122594);
nor I_7054 (I122173,I122450,I122611);
nand I_7055 (I122158,I122467,I122611);
nor I_7056 (I122167,I122213,I122594);
DFFARX1 I_7057 (I122594,I2683,I122187,I122176,);
not I_7058 (I122714,I2690);
DFFARX1 I_7059 (I171858,I2683,I122714,I122740,);
nand I_7060 (I122748,I171843,I171846);
and I_7061 (I122765,I122748,I171861);
DFFARX1 I_7062 (I122765,I2683,I122714,I122791,);
nor I_7063 (I122682,I122791,I122740);
not I_7064 (I122813,I122791);
DFFARX1 I_7065 (I171855,I2683,I122714,I122839,);
nand I_7066 (I122847,I122839,I171846);
not I_7067 (I122864,I122847);
DFFARX1 I_7068 (I122864,I2683,I122714,I122890,);
not I_7069 (I122706,I122890);
nor I_7070 (I122912,I122740,I122847);
nor I_7071 (I122688,I122791,I122912);
DFFARX1 I_7072 (I171852,I2683,I122714,I122952,);
DFFARX1 I_7073 (I122952,I2683,I122714,I122969,);
not I_7074 (I122977,I122969);
not I_7075 (I122994,I122952);
nand I_7076 (I122691,I122994,I122813);
nand I_7077 (I123025,I171867,I171843);
and I_7078 (I123042,I123025,I171864);
DFFARX1 I_7079 (I123042,I2683,I122714,I123068,);
nor I_7080 (I123076,I123068,I122740);
DFFARX1 I_7081 (I123076,I2683,I122714,I122679,);
DFFARX1 I_7082 (I123068,I2683,I122714,I122697,);
nor I_7083 (I123121,I171849,I171843);
not I_7084 (I123138,I123121);
nor I_7085 (I122700,I122977,I123138);
nand I_7086 (I122685,I122994,I123138);
nor I_7087 (I122694,I122740,I123121);
DFFARX1 I_7088 (I123121,I2683,I122714,I122703,);
not I_7089 (I123241,I2690);
DFFARX1 I_7090 (I137243,I2683,I123241,I123267,);
nand I_7091 (I123275,I137255,I137234);
and I_7092 (I123292,I123275,I137258);
DFFARX1 I_7093 (I123292,I2683,I123241,I123318,);
nor I_7094 (I123209,I123318,I123267);
not I_7095 (I123340,I123318);
DFFARX1 I_7096 (I137249,I2683,I123241,I123366,);
nand I_7097 (I123374,I123366,I137231);
not I_7098 (I123391,I123374);
DFFARX1 I_7099 (I123391,I2683,I123241,I123417,);
not I_7100 (I123233,I123417);
nor I_7101 (I123439,I123267,I123374);
nor I_7102 (I123215,I123318,I123439);
DFFARX1 I_7103 (I137246,I2683,I123241,I123479,);
DFFARX1 I_7104 (I123479,I2683,I123241,I123496,);
not I_7105 (I123504,I123496);
not I_7106 (I123521,I123479);
nand I_7107 (I123218,I123521,I123340);
nand I_7108 (I123552,I137231,I137237);
and I_7109 (I123569,I123552,I137240);
DFFARX1 I_7110 (I123569,I2683,I123241,I123595,);
nor I_7111 (I123603,I123595,I123267);
DFFARX1 I_7112 (I123603,I2683,I123241,I123206,);
DFFARX1 I_7113 (I123595,I2683,I123241,I123224,);
nor I_7114 (I123648,I137252,I137237);
not I_7115 (I123665,I123648);
nor I_7116 (I123227,I123504,I123665);
nand I_7117 (I123212,I123521,I123665);
nor I_7118 (I123221,I123267,I123648);
DFFARX1 I_7119 (I123648,I2683,I123241,I123230,);
not I_7120 (I123768,I2690);
DFFARX1 I_7121 (I355069,I2683,I123768,I123794,);
nand I_7122 (I123802,I355084,I355069);
and I_7123 (I123819,I123802,I355087);
DFFARX1 I_7124 (I123819,I2683,I123768,I123845,);
nor I_7125 (I123736,I123845,I123794);
not I_7126 (I123867,I123845);
DFFARX1 I_7127 (I355093,I2683,I123768,I123893,);
nand I_7128 (I123901,I123893,I355075);
not I_7129 (I123918,I123901);
DFFARX1 I_7130 (I123918,I2683,I123768,I123944,);
not I_7131 (I123760,I123944);
nor I_7132 (I123966,I123794,I123901);
nor I_7133 (I123742,I123845,I123966);
DFFARX1 I_7134 (I355072,I2683,I123768,I124006,);
DFFARX1 I_7135 (I124006,I2683,I123768,I124023,);
not I_7136 (I124031,I124023);
not I_7137 (I124048,I124006);
nand I_7138 (I123745,I124048,I123867);
nand I_7139 (I124079,I355072,I355078);
and I_7140 (I124096,I124079,I355090);
DFFARX1 I_7141 (I124096,I2683,I123768,I124122,);
nor I_7142 (I124130,I124122,I123794);
DFFARX1 I_7143 (I124130,I2683,I123768,I123733,);
DFFARX1 I_7144 (I124122,I2683,I123768,I123751,);
nor I_7145 (I124175,I355081,I355078);
not I_7146 (I124192,I124175);
nor I_7147 (I123754,I124031,I124192);
nand I_7148 (I123739,I124048,I124192);
nor I_7149 (I123748,I123794,I124175);
DFFARX1 I_7150 (I124175,I2683,I123768,I123757,);
not I_7151 (I124295,I2690);
DFFARX1 I_7152 (I203645,I2683,I124295,I124321,);
nand I_7153 (I124329,I203636,I203651);
and I_7154 (I124346,I124329,I203657);
DFFARX1 I_7155 (I124346,I2683,I124295,I124372,);
nor I_7156 (I124263,I124372,I124321);
not I_7157 (I124394,I124372);
DFFARX1 I_7158 (I203642,I2683,I124295,I124420,);
nand I_7159 (I124428,I124420,I203636);
not I_7160 (I124445,I124428);
DFFARX1 I_7161 (I124445,I2683,I124295,I124471,);
not I_7162 (I124287,I124471);
nor I_7163 (I124493,I124321,I124428);
nor I_7164 (I124269,I124372,I124493);
DFFARX1 I_7165 (I203639,I2683,I124295,I124533,);
DFFARX1 I_7166 (I124533,I2683,I124295,I124550,);
not I_7167 (I124558,I124550);
not I_7168 (I124575,I124533);
nand I_7169 (I124272,I124575,I124394);
nand I_7170 (I124606,I203633,I203648);
and I_7171 (I124623,I124606,I203633);
DFFARX1 I_7172 (I124623,I2683,I124295,I124649,);
nor I_7173 (I124657,I124649,I124321);
DFFARX1 I_7174 (I124657,I2683,I124295,I124260,);
DFFARX1 I_7175 (I124649,I2683,I124295,I124278,);
nor I_7176 (I124702,I203654,I203648);
not I_7177 (I124719,I124702);
nor I_7178 (I124281,I124558,I124719);
nand I_7179 (I124266,I124575,I124719);
nor I_7180 (I124275,I124321,I124702);
DFFARX1 I_7181 (I124702,I2683,I124295,I124284,);
not I_7182 (I124822,I2690);
DFFARX1 I_7183 (I205379,I2683,I124822,I124848,);
nand I_7184 (I124856,I205370,I205385);
and I_7185 (I124873,I124856,I205391);
DFFARX1 I_7186 (I124873,I2683,I124822,I124899,);
nor I_7187 (I124790,I124899,I124848);
not I_7188 (I124921,I124899);
DFFARX1 I_7189 (I205376,I2683,I124822,I124947,);
nand I_7190 (I124955,I124947,I205370);
not I_7191 (I124972,I124955);
DFFARX1 I_7192 (I124972,I2683,I124822,I124998,);
not I_7193 (I124814,I124998);
nor I_7194 (I125020,I124848,I124955);
nor I_7195 (I124796,I124899,I125020);
DFFARX1 I_7196 (I205373,I2683,I124822,I125060,);
DFFARX1 I_7197 (I125060,I2683,I124822,I125077,);
not I_7198 (I125085,I125077);
not I_7199 (I125102,I125060);
nand I_7200 (I124799,I125102,I124921);
nand I_7201 (I125133,I205367,I205382);
and I_7202 (I125150,I125133,I205367);
DFFARX1 I_7203 (I125150,I2683,I124822,I125176,);
nor I_7204 (I125184,I125176,I124848);
DFFARX1 I_7205 (I125184,I2683,I124822,I124787,);
DFFARX1 I_7206 (I125176,I2683,I124822,I124805,);
nor I_7207 (I125229,I205388,I205382);
not I_7208 (I125246,I125229);
nor I_7209 (I124808,I125085,I125246);
nand I_7210 (I124793,I125102,I125246);
nor I_7211 (I124802,I124848,I125229);
DFFARX1 I_7212 (I125229,I2683,I124822,I124811,);
not I_7213 (I125349,I2690);
DFFARX1 I_7214 (I177638,I2683,I125349,I125375,);
nand I_7215 (I125383,I177623,I177626);
and I_7216 (I125400,I125383,I177641);
DFFARX1 I_7217 (I125400,I2683,I125349,I125426,);
nor I_7218 (I125317,I125426,I125375);
not I_7219 (I125448,I125426);
DFFARX1 I_7220 (I177635,I2683,I125349,I125474,);
nand I_7221 (I125482,I125474,I177626);
not I_7222 (I125499,I125482);
DFFARX1 I_7223 (I125499,I2683,I125349,I125525,);
not I_7224 (I125341,I125525);
nor I_7225 (I125547,I125375,I125482);
nor I_7226 (I125323,I125426,I125547);
DFFARX1 I_7227 (I177632,I2683,I125349,I125587,);
DFFARX1 I_7228 (I125587,I2683,I125349,I125604,);
not I_7229 (I125612,I125604);
not I_7230 (I125629,I125587);
nand I_7231 (I125326,I125629,I125448);
nand I_7232 (I125660,I177647,I177623);
and I_7233 (I125677,I125660,I177644);
DFFARX1 I_7234 (I125677,I2683,I125349,I125703,);
nor I_7235 (I125711,I125703,I125375);
DFFARX1 I_7236 (I125711,I2683,I125349,I125314,);
DFFARX1 I_7237 (I125703,I2683,I125349,I125332,);
nor I_7238 (I125756,I177629,I177623);
not I_7239 (I125773,I125756);
nor I_7240 (I125335,I125612,I125773);
nand I_7241 (I125320,I125629,I125773);
nor I_7242 (I125329,I125375,I125756);
DFFARX1 I_7243 (I125756,I2683,I125349,I125338,);
not I_7244 (I125876,I2690);
DFFARX1 I_7245 (I74484,I2683,I125876,I125902,);
nand I_7246 (I125910,I74484,I74490);
and I_7247 (I125927,I125910,I74508);
DFFARX1 I_7248 (I125927,I2683,I125876,I125953,);
nor I_7249 (I125844,I125953,I125902);
not I_7250 (I125975,I125953);
DFFARX1 I_7251 (I74496,I2683,I125876,I126001,);
nand I_7252 (I126009,I126001,I74493);
not I_7253 (I126026,I126009);
DFFARX1 I_7254 (I126026,I2683,I125876,I126052,);
not I_7255 (I125868,I126052);
nor I_7256 (I126074,I125902,I126009);
nor I_7257 (I125850,I125953,I126074);
DFFARX1 I_7258 (I74502,I2683,I125876,I126114,);
DFFARX1 I_7259 (I126114,I2683,I125876,I126131,);
not I_7260 (I126139,I126131);
not I_7261 (I126156,I126114);
nand I_7262 (I125853,I126156,I125975);
nand I_7263 (I126187,I74487,I74487);
and I_7264 (I126204,I126187,I74499);
DFFARX1 I_7265 (I126204,I2683,I125876,I126230,);
nor I_7266 (I126238,I126230,I125902);
DFFARX1 I_7267 (I126238,I2683,I125876,I125841,);
DFFARX1 I_7268 (I126230,I2683,I125876,I125859,);
nor I_7269 (I126283,I74505,I74487);
not I_7270 (I126300,I126283);
nor I_7271 (I125862,I126139,I126300);
nand I_7272 (I125847,I126156,I126300);
nor I_7273 (I125856,I125902,I126283);
DFFARX1 I_7274 (I126283,I2683,I125876,I125865,);
not I_7275 (I126403,I2690);
DFFARX1 I_7276 (I32021,I2683,I126403,I126429,);
nand I_7277 (I126437,I32033,I32042);
and I_7278 (I126454,I126437,I32021);
DFFARX1 I_7279 (I126454,I2683,I126403,I126480,);
nor I_7280 (I126371,I126480,I126429);
not I_7281 (I126502,I126480);
DFFARX1 I_7282 (I32036,I2683,I126403,I126528,);
nand I_7283 (I126536,I126528,I32024);
not I_7284 (I126553,I126536);
DFFARX1 I_7285 (I126553,I2683,I126403,I126579,);
not I_7286 (I126395,I126579);
nor I_7287 (I126601,I126429,I126536);
nor I_7288 (I126377,I126480,I126601);
DFFARX1 I_7289 (I32027,I2683,I126403,I126641,);
DFFARX1 I_7290 (I126641,I2683,I126403,I126658,);
not I_7291 (I126666,I126658);
not I_7292 (I126683,I126641);
nand I_7293 (I126380,I126683,I126502);
nand I_7294 (I126714,I32018,I32018);
and I_7295 (I126731,I126714,I32030);
DFFARX1 I_7296 (I126731,I2683,I126403,I126757,);
nor I_7297 (I126765,I126757,I126429);
DFFARX1 I_7298 (I126765,I2683,I126403,I126368,);
DFFARX1 I_7299 (I126757,I2683,I126403,I126386,);
nor I_7300 (I126810,I32039,I32018);
not I_7301 (I126827,I126810);
nor I_7302 (I126389,I126666,I126827);
nand I_7303 (I126374,I126683,I126827);
nor I_7304 (I126383,I126429,I126810);
DFFARX1 I_7305 (I126810,I2683,I126403,I126392,);
not I_7306 (I126930,I2690);
DFFARX1 I_7307 (I170690,I2683,I126930,I126956,);
DFFARX1 I_7308 (I126956,I2683,I126930,I126973,);
not I_7309 (I126922,I126973);
not I_7310 (I126995,I126956);
nand I_7311 (I127012,I170687,I170708);
and I_7312 (I127029,I127012,I170711);
DFFARX1 I_7313 (I127029,I2683,I126930,I127055,);
not I_7314 (I127063,I127055);
DFFARX1 I_7315 (I170696,I2683,I126930,I127089,);
and I_7316 (I127097,I127089,I170699);
nand I_7317 (I127114,I127089,I170699);
nand I_7318 (I126901,I127063,I127114);
DFFARX1 I_7319 (I170702,I2683,I126930,I127154,);
nor I_7320 (I127162,I127154,I127097);
DFFARX1 I_7321 (I127162,I2683,I126930,I126895,);
nor I_7322 (I126910,I127154,I127055);
nand I_7323 (I127207,I170687,I170693);
and I_7324 (I127224,I127207,I170705);
DFFARX1 I_7325 (I127224,I2683,I126930,I127250,);
nor I_7326 (I126898,I127250,I127154);
not I_7327 (I127272,I127250);
nor I_7328 (I127289,I127272,I127063);
nor I_7329 (I127306,I126995,I127289);
DFFARX1 I_7330 (I127306,I2683,I126930,I126913,);
nor I_7331 (I127337,I127272,I127154);
nor I_7332 (I127354,I170690,I170693);
nor I_7333 (I126904,I127354,I127337);
not I_7334 (I127385,I127354);
nand I_7335 (I126907,I127114,I127385);
DFFARX1 I_7336 (I127354,I2683,I126930,I126919,);
DFFARX1 I_7337 (I127354,I2683,I126930,I126916,);
not I_7338 (I127474,I2690);
DFFARX1 I_7339 (I86864,I2683,I127474,I127500,);
DFFARX1 I_7340 (I127500,I2683,I127474,I127517,);
not I_7341 (I127466,I127517);
not I_7342 (I127539,I127500);
nand I_7343 (I127556,I86843,I86867);
and I_7344 (I127573,I127556,I86870);
DFFARX1 I_7345 (I127573,I2683,I127474,I127599,);
not I_7346 (I127607,I127599);
DFFARX1 I_7347 (I86852,I2683,I127474,I127633,);
and I_7348 (I127641,I127633,I86858);
nand I_7349 (I127658,I127633,I86858);
nand I_7350 (I127445,I127607,I127658);
DFFARX1 I_7351 (I86846,I2683,I127474,I127698,);
nor I_7352 (I127706,I127698,I127641);
DFFARX1 I_7353 (I127706,I2683,I127474,I127439,);
nor I_7354 (I127454,I127698,I127599);
nand I_7355 (I127751,I86855,I86843);
and I_7356 (I127768,I127751,I86849);
DFFARX1 I_7357 (I127768,I2683,I127474,I127794,);
nor I_7358 (I127442,I127794,I127698);
not I_7359 (I127816,I127794);
nor I_7360 (I127833,I127816,I127607);
nor I_7361 (I127850,I127539,I127833);
DFFARX1 I_7362 (I127850,I2683,I127474,I127457,);
nor I_7363 (I127881,I127816,I127698);
nor I_7364 (I127898,I86861,I86843);
nor I_7365 (I127448,I127898,I127881);
not I_7366 (I127929,I127898);
nand I_7367 (I127451,I127658,I127929);
DFFARX1 I_7368 (I127898,I2683,I127474,I127463,);
DFFARX1 I_7369 (I127898,I2683,I127474,I127460,);
not I_7370 (I128018,I2690);
DFFARX1 I_7371 (I111633,I2683,I128018,I128044,);
DFFARX1 I_7372 (I128044,I2683,I128018,I128061,);
not I_7373 (I128010,I128061);
not I_7374 (I128083,I128044);
nand I_7375 (I128100,I111612,I111636);
and I_7376 (I128117,I128100,I111639);
DFFARX1 I_7377 (I128117,I2683,I128018,I128143,);
not I_7378 (I128151,I128143);
DFFARX1 I_7379 (I111621,I2683,I128018,I128177,);
and I_7380 (I128185,I128177,I111627);
nand I_7381 (I128202,I128177,I111627);
nand I_7382 (I127989,I128151,I128202);
DFFARX1 I_7383 (I111615,I2683,I128018,I128242,);
nor I_7384 (I128250,I128242,I128185);
DFFARX1 I_7385 (I128250,I2683,I128018,I127983,);
nor I_7386 (I127998,I128242,I128143);
nand I_7387 (I128295,I111624,I111612);
and I_7388 (I128312,I128295,I111618);
DFFARX1 I_7389 (I128312,I2683,I128018,I128338,);
nor I_7390 (I127986,I128338,I128242);
not I_7391 (I128360,I128338);
nor I_7392 (I128377,I128360,I128151);
nor I_7393 (I128394,I128083,I128377);
DFFARX1 I_7394 (I128394,I2683,I128018,I128001,);
nor I_7395 (I128425,I128360,I128242);
nor I_7396 (I128442,I111630,I111612);
nor I_7397 (I127992,I128442,I128425);
not I_7398 (I128473,I128442);
nand I_7399 (I127995,I128202,I128473);
DFFARX1 I_7400 (I128442,I2683,I128018,I128007,);
DFFARX1 I_7401 (I128442,I2683,I128018,I128004,);
not I_7402 (I128562,I2690);
DFFARX1 I_7403 (I263995,I2683,I128562,I128588,);
DFFARX1 I_7404 (I128588,I2683,I128562,I128605,);
not I_7405 (I128554,I128605);
not I_7406 (I128627,I128588);
nand I_7407 (I128644,I263989,I263986);
and I_7408 (I128661,I128644,I264001);
DFFARX1 I_7409 (I128661,I2683,I128562,I128687,);
not I_7410 (I128695,I128687);
DFFARX1 I_7411 (I263989,I2683,I128562,I128721,);
and I_7412 (I128729,I128721,I263983);
nand I_7413 (I128746,I128721,I263983);
nand I_7414 (I128533,I128695,I128746);
DFFARX1 I_7415 (I263983,I2683,I128562,I128786,);
nor I_7416 (I128794,I128786,I128729);
DFFARX1 I_7417 (I128794,I2683,I128562,I128527,);
nor I_7418 (I128542,I128786,I128687);
nand I_7419 (I128839,I263998,I263992);
and I_7420 (I128856,I128839,I263986);
DFFARX1 I_7421 (I128856,I2683,I128562,I128882,);
nor I_7422 (I128530,I128882,I128786);
not I_7423 (I128904,I128882);
nor I_7424 (I128921,I128904,I128695);
nor I_7425 (I128938,I128627,I128921);
DFFARX1 I_7426 (I128938,I2683,I128562,I128545,);
nor I_7427 (I128969,I128904,I128786);
nor I_7428 (I128986,I264004,I263992);
nor I_7429 (I128536,I128986,I128969);
not I_7430 (I129017,I128986);
nand I_7431 (I128539,I128746,I129017);
DFFARX1 I_7432 (I128986,I2683,I128562,I128551,);
DFFARX1 I_7433 (I128986,I2683,I128562,I128548,);
not I_7434 (I129106,I2690);
DFFARX1 I_7435 (I402186,I2683,I129106,I129132,);
DFFARX1 I_7436 (I129132,I2683,I129106,I129149,);
not I_7437 (I129098,I129149);
not I_7438 (I129171,I129132);
nand I_7439 (I129188,I402162,I402183);
and I_7440 (I129205,I129188,I402180);
DFFARX1 I_7441 (I129205,I2683,I129106,I129231,);
not I_7442 (I129239,I129231);
DFFARX1 I_7443 (I402159,I2683,I129106,I129265,);
and I_7444 (I129273,I129265,I402171);
nand I_7445 (I129290,I129265,I402171);
nand I_7446 (I129077,I129239,I129290);
DFFARX1 I_7447 (I402174,I2683,I129106,I129330,);
nor I_7448 (I129338,I129330,I129273);
DFFARX1 I_7449 (I129338,I2683,I129106,I129071,);
nor I_7450 (I129086,I129330,I129231);
nand I_7451 (I129383,I402177,I402165);
and I_7452 (I129400,I129383,I402168);
DFFARX1 I_7453 (I129400,I2683,I129106,I129426,);
nor I_7454 (I129074,I129426,I129330);
not I_7455 (I129448,I129426);
nor I_7456 (I129465,I129448,I129239);
nor I_7457 (I129482,I129171,I129465);
DFFARX1 I_7458 (I129482,I2683,I129106,I129089,);
nor I_7459 (I129513,I129448,I129330);
nor I_7460 (I129530,I402159,I402165);
nor I_7461 (I129080,I129530,I129513);
not I_7462 (I129561,I129530);
nand I_7463 (I129083,I129290,I129561);
DFFARX1 I_7464 (I129530,I2683,I129106,I129095,);
DFFARX1 I_7465 (I129530,I2683,I129106,I129092,);
not I_7466 (I129650,I2690);
DFFARX1 I_7467 (I122700,I2683,I129650,I129676,);
DFFARX1 I_7468 (I129676,I2683,I129650,I129693,);
not I_7469 (I129642,I129693);
not I_7470 (I129715,I129676);
nand I_7471 (I129732,I122679,I122703);
and I_7472 (I129749,I129732,I122706);
DFFARX1 I_7473 (I129749,I2683,I129650,I129775,);
not I_7474 (I129783,I129775);
DFFARX1 I_7475 (I122688,I2683,I129650,I129809,);
and I_7476 (I129817,I129809,I122694);
nand I_7477 (I129834,I129809,I122694);
nand I_7478 (I129621,I129783,I129834);
DFFARX1 I_7479 (I122682,I2683,I129650,I129874,);
nor I_7480 (I129882,I129874,I129817);
DFFARX1 I_7481 (I129882,I2683,I129650,I129615,);
nor I_7482 (I129630,I129874,I129775);
nand I_7483 (I129927,I122691,I122679);
and I_7484 (I129944,I129927,I122685);
DFFARX1 I_7485 (I129944,I2683,I129650,I129970,);
nor I_7486 (I129618,I129970,I129874);
not I_7487 (I129992,I129970);
nor I_7488 (I130009,I129992,I129783);
nor I_7489 (I130026,I129715,I130009);
DFFARX1 I_7490 (I130026,I2683,I129650,I129633,);
nor I_7491 (I130057,I129992,I129874);
nor I_7492 (I130074,I122697,I122679);
nor I_7493 (I129624,I130074,I130057);
not I_7494 (I130105,I130074);
nand I_7495 (I129627,I129834,I130105);
DFFARX1 I_7496 (I130074,I2683,I129650,I129639,);
DFFARX1 I_7497 (I130074,I2683,I129650,I129636,);
not I_7498 (I130194,I2690);
DFFARX1 I_7499 (I81038,I2683,I130194,I130220,);
DFFARX1 I_7500 (I130220,I2683,I130194,I130237,);
not I_7501 (I130186,I130237);
not I_7502 (I130259,I130220);
nand I_7503 (I130276,I81050,I81029);
and I_7504 (I130293,I130276,I81032);
DFFARX1 I_7505 (I130293,I2683,I130194,I130319,);
not I_7506 (I130327,I130319);
DFFARX1 I_7507 (I81041,I2683,I130194,I130353,);
and I_7508 (I130361,I130353,I81053);
nand I_7509 (I130378,I130353,I81053);
nand I_7510 (I130165,I130327,I130378);
DFFARX1 I_7511 (I81047,I2683,I130194,I130418,);
nor I_7512 (I130426,I130418,I130361);
DFFARX1 I_7513 (I130426,I2683,I130194,I130159,);
nor I_7514 (I130174,I130418,I130319);
nand I_7515 (I130471,I81035,I81032);
and I_7516 (I130488,I130471,I81044);
DFFARX1 I_7517 (I130488,I2683,I130194,I130514,);
nor I_7518 (I130162,I130514,I130418);
not I_7519 (I130536,I130514);
nor I_7520 (I130553,I130536,I130327);
nor I_7521 (I130570,I130259,I130553);
DFFARX1 I_7522 (I130570,I2683,I130194,I130177,);
nor I_7523 (I130601,I130536,I130418);
nor I_7524 (I130618,I81029,I81032);
nor I_7525 (I130168,I130618,I130601);
not I_7526 (I130649,I130618);
nand I_7527 (I130171,I130378,I130649);
DFFARX1 I_7528 (I130618,I2683,I130194,I130183,);
DFFARX1 I_7529 (I130618,I2683,I130194,I130180,);
not I_7530 (I130738,I2690);
DFFARX1 I_7531 (I199012,I2683,I130738,I130764,);
DFFARX1 I_7532 (I130764,I2683,I130738,I130781,);
not I_7533 (I130730,I130781);
not I_7534 (I130803,I130764);
nand I_7535 (I130820,I199033,I199024);
and I_7536 (I130837,I130820,I199012);
DFFARX1 I_7537 (I130837,I2683,I130738,I130863,);
not I_7538 (I130871,I130863);
DFFARX1 I_7539 (I199018,I2683,I130738,I130897,);
and I_7540 (I130905,I130897,I199015);
nand I_7541 (I130922,I130897,I199015);
nand I_7542 (I130709,I130871,I130922);
DFFARX1 I_7543 (I199009,I2683,I130738,I130962,);
nor I_7544 (I130970,I130962,I130905);
DFFARX1 I_7545 (I130970,I2683,I130738,I130703,);
nor I_7546 (I130718,I130962,I130863);
nand I_7547 (I131015,I199009,I199021);
and I_7548 (I131032,I131015,I199030);
DFFARX1 I_7549 (I131032,I2683,I130738,I131058,);
nor I_7550 (I130706,I131058,I130962);
not I_7551 (I131080,I131058);
nor I_7552 (I131097,I131080,I130871);
nor I_7553 (I131114,I130803,I131097);
DFFARX1 I_7554 (I131114,I2683,I130738,I130721,);
nor I_7555 (I131145,I131080,I130962);
nor I_7556 (I131162,I199027,I199021);
nor I_7557 (I130712,I131162,I131145);
not I_7558 (I131193,I131162);
nand I_7559 (I130715,I130922,I131193);
DFFARX1 I_7560 (I131162,I2683,I130738,I130727,);
DFFARX1 I_7561 (I131162,I2683,I130738,I130724,);
not I_7562 (I131282,I2690);
DFFARX1 I_7563 (I53073,I2683,I131282,I131308,);
DFFARX1 I_7564 (I131308,I2683,I131282,I131325,);
not I_7565 (I131274,I131325);
not I_7566 (I131347,I131308);
nand I_7567 (I131364,I53085,I53064);
and I_7568 (I131381,I131364,I53067);
DFFARX1 I_7569 (I131381,I2683,I131282,I131407,);
not I_7570 (I131415,I131407);
DFFARX1 I_7571 (I53076,I2683,I131282,I131441,);
and I_7572 (I131449,I131441,I53088);
nand I_7573 (I131466,I131441,I53088);
nand I_7574 (I131253,I131415,I131466);
DFFARX1 I_7575 (I53082,I2683,I131282,I131506,);
nor I_7576 (I131514,I131506,I131449);
DFFARX1 I_7577 (I131514,I2683,I131282,I131247,);
nor I_7578 (I131262,I131506,I131407);
nand I_7579 (I131559,I53070,I53067);
and I_7580 (I131576,I131559,I53079);
DFFARX1 I_7581 (I131576,I2683,I131282,I131602,);
nor I_7582 (I131250,I131602,I131506);
not I_7583 (I131624,I131602);
nor I_7584 (I131641,I131624,I131415);
nor I_7585 (I131658,I131347,I131641);
DFFARX1 I_7586 (I131658,I2683,I131282,I131265,);
nor I_7587 (I131689,I131624,I131506);
nor I_7588 (I131706,I53064,I53067);
nor I_7589 (I131256,I131706,I131689);
not I_7590 (I131737,I131706);
nand I_7591 (I131259,I131466,I131737);
DFFARX1 I_7592 (I131706,I2683,I131282,I131271,);
DFFARX1 I_7593 (I131706,I2683,I131282,I131268,);
not I_7594 (I131826,I2690);
DFFARX1 I_7595 (I332530,I2683,I131826,I131852,);
DFFARX1 I_7596 (I131852,I2683,I131826,I131869,);
not I_7597 (I131818,I131869);
not I_7598 (I131891,I131852);
nand I_7599 (I131908,I332542,I332530);
and I_7600 (I131925,I131908,I332533);
DFFARX1 I_7601 (I131925,I2683,I131826,I131951,);
not I_7602 (I131959,I131951);
DFFARX1 I_7603 (I332551,I2683,I131826,I131985,);
and I_7604 (I131993,I131985,I332527);
nand I_7605 (I132010,I131985,I332527);
nand I_7606 (I131797,I131959,I132010);
DFFARX1 I_7607 (I332545,I2683,I131826,I132050,);
nor I_7608 (I132058,I132050,I131993);
DFFARX1 I_7609 (I132058,I2683,I131826,I131791,);
nor I_7610 (I131806,I132050,I131951);
nand I_7611 (I132103,I332539,I332536);
and I_7612 (I132120,I132103,I332548);
DFFARX1 I_7613 (I132120,I2683,I131826,I132146,);
nor I_7614 (I131794,I132146,I132050);
not I_7615 (I132168,I132146);
nor I_7616 (I132185,I132168,I131959);
nor I_7617 (I132202,I131891,I132185);
DFFARX1 I_7618 (I132202,I2683,I131826,I131809,);
nor I_7619 (I132233,I132168,I132050);
nor I_7620 (I132250,I332527,I332536);
nor I_7621 (I131800,I132250,I132233);
not I_7622 (I132281,I132250);
nand I_7623 (I131803,I132010,I132281);
DFFARX1 I_7624 (I132250,I2683,I131826,I131815,);
DFFARX1 I_7625 (I132250,I2683,I131826,I131812,);
not I_7626 (I132370,I2690);
DFFARX1 I_7627 (I161187,I2683,I132370,I132396,);
DFFARX1 I_7628 (I132396,I2683,I132370,I132413,);
not I_7629 (I132362,I132413);
not I_7630 (I132435,I132396);
nand I_7631 (I132452,I161190,I161208);
and I_7632 (I132469,I132452,I161196);
DFFARX1 I_7633 (I132469,I2683,I132370,I132495,);
not I_7634 (I132503,I132495);
DFFARX1 I_7635 (I161187,I2683,I132370,I132529,);
and I_7636 (I132537,I132529,I161205);
nand I_7637 (I132554,I132529,I161205);
nand I_7638 (I132341,I132503,I132554);
DFFARX1 I_7639 (I161199,I2683,I132370,I132594,);
nor I_7640 (I132602,I132594,I132537);
DFFARX1 I_7641 (I132602,I2683,I132370,I132335,);
nor I_7642 (I132350,I132594,I132495);
nand I_7643 (I132647,I161202,I161184);
and I_7644 (I132664,I132647,I161193);
DFFARX1 I_7645 (I132664,I2683,I132370,I132690,);
nor I_7646 (I132338,I132690,I132594);
not I_7647 (I132712,I132690);
nor I_7648 (I132729,I132712,I132503);
nor I_7649 (I132746,I132435,I132729);
DFFARX1 I_7650 (I132746,I2683,I132370,I132353,);
nor I_7651 (I132777,I132712,I132594);
nor I_7652 (I132794,I161184,I161184);
nor I_7653 (I132344,I132794,I132777);
not I_7654 (I132825,I132794);
nand I_7655 (I132347,I132554,I132825);
DFFARX1 I_7656 (I132794,I2683,I132370,I132359,);
DFFARX1 I_7657 (I132794,I2683,I132370,I132356,);
not I_7658 (I132914,I2690);
DFFARX1 I_7659 (I248712,I2683,I132914,I132940,);
DFFARX1 I_7660 (I132940,I2683,I132914,I132957,);
not I_7661 (I132906,I132957);
not I_7662 (I132979,I132940);
nand I_7663 (I132996,I248706,I248703);
and I_7664 (I133013,I132996,I248718);
DFFARX1 I_7665 (I133013,I2683,I132914,I133039,);
not I_7666 (I133047,I133039);
DFFARX1 I_7667 (I248706,I2683,I132914,I133073,);
and I_7668 (I133081,I133073,I248700);
nand I_7669 (I133098,I133073,I248700);
nand I_7670 (I132885,I133047,I133098);
DFFARX1 I_7671 (I248700,I2683,I132914,I133138,);
nor I_7672 (I133146,I133138,I133081);
DFFARX1 I_7673 (I133146,I2683,I132914,I132879,);
nor I_7674 (I132894,I133138,I133039);
nand I_7675 (I133191,I248715,I248709);
and I_7676 (I133208,I133191,I248703);
DFFARX1 I_7677 (I133208,I2683,I132914,I133234,);
nor I_7678 (I132882,I133234,I133138);
not I_7679 (I133256,I133234);
nor I_7680 (I133273,I133256,I133047);
nor I_7681 (I133290,I132979,I133273);
DFFARX1 I_7682 (I133290,I2683,I132914,I132897,);
nor I_7683 (I133321,I133256,I133138);
nor I_7684 (I133338,I248721,I248709);
nor I_7685 (I132888,I133338,I133321);
not I_7686 (I133369,I133338);
nand I_7687 (I132891,I133098,I133369);
DFFARX1 I_7688 (I133338,I2683,I132914,I132903,);
DFFARX1 I_7689 (I133338,I2683,I132914,I132900,);
not I_7690 (I133458,I2690);
DFFARX1 I_7691 (I325016,I2683,I133458,I133484,);
DFFARX1 I_7692 (I133484,I2683,I133458,I133501,);
not I_7693 (I133450,I133501);
not I_7694 (I133523,I133484);
nand I_7695 (I133540,I325028,I325016);
and I_7696 (I133557,I133540,I325019);
DFFARX1 I_7697 (I133557,I2683,I133458,I133583,);
not I_7698 (I133591,I133583);
DFFARX1 I_7699 (I325037,I2683,I133458,I133617,);
and I_7700 (I133625,I133617,I325013);
nand I_7701 (I133642,I133617,I325013);
nand I_7702 (I133429,I133591,I133642);
DFFARX1 I_7703 (I325031,I2683,I133458,I133682,);
nor I_7704 (I133690,I133682,I133625);
DFFARX1 I_7705 (I133690,I2683,I133458,I133423,);
nor I_7706 (I133438,I133682,I133583);
nand I_7707 (I133735,I325025,I325022);
and I_7708 (I133752,I133735,I325034);
DFFARX1 I_7709 (I133752,I2683,I133458,I133778,);
nor I_7710 (I133426,I133778,I133682);
not I_7711 (I133800,I133778);
nor I_7712 (I133817,I133800,I133591);
nor I_7713 (I133834,I133523,I133817);
DFFARX1 I_7714 (I133834,I2683,I133458,I133441,);
nor I_7715 (I133865,I133800,I133682);
nor I_7716 (I133882,I325013,I325022);
nor I_7717 (I133432,I133882,I133865);
not I_7718 (I133913,I133882);
nand I_7719 (I133435,I133642,I133913);
DFFARX1 I_7720 (I133882,I2683,I133458,I133447,);
DFFARX1 I_7721 (I133882,I2683,I133458,I133444,);
not I_7722 (I134002,I2690);
DFFARX1 I_7723 (I47721,I2683,I134002,I134028,);
DFFARX1 I_7724 (I134028,I2683,I134002,I134045,);
not I_7725 (I133994,I134045);
not I_7726 (I134067,I134028);
nand I_7727 (I134084,I47730,I47733);
and I_7728 (I134101,I134084,I47712);
DFFARX1 I_7729 (I134101,I2683,I134002,I134127,);
not I_7730 (I134135,I134127);
DFFARX1 I_7731 (I47727,I2683,I134002,I134161,);
and I_7732 (I134169,I134161,I47715);
nand I_7733 (I134186,I134161,I47715);
nand I_7734 (I133973,I134135,I134186);
DFFARX1 I_7735 (I47709,I2683,I134002,I134226,);
nor I_7736 (I134234,I134226,I134169);
DFFARX1 I_7737 (I134234,I2683,I134002,I133967,);
nor I_7738 (I133982,I134226,I134127);
nand I_7739 (I134279,I47724,I47718);
and I_7740 (I134296,I134279,I47709);
DFFARX1 I_7741 (I134296,I2683,I134002,I134322,);
nor I_7742 (I133970,I134322,I134226);
not I_7743 (I134344,I134322);
nor I_7744 (I134361,I134344,I134135);
nor I_7745 (I134378,I134067,I134361);
DFFARX1 I_7746 (I134378,I2683,I134002,I133985,);
nor I_7747 (I134409,I134344,I134226);
nor I_7748 (I134426,I47736,I47718);
nor I_7749 (I133976,I134426,I134409);
not I_7750 (I134457,I134426);
nand I_7751 (I133979,I134186,I134457);
DFFARX1 I_7752 (I134426,I2683,I134002,I133991,);
DFFARX1 I_7753 (I134426,I2683,I134002,I133988,);
not I_7754 (I134546,I2690);
DFFARX1 I_7755 (I321613,I2683,I134546,I134572,);
DFFARX1 I_7756 (I134572,I2683,I134546,I134589,);
not I_7757 (I134538,I134589);
not I_7758 (I134611,I134572);
nand I_7759 (I134628,I321613,I321631);
and I_7760 (I134645,I134628,I321625);
DFFARX1 I_7761 (I134645,I2683,I134546,I134671,);
not I_7762 (I134679,I134671);
DFFARX1 I_7763 (I321619,I2683,I134546,I134705,);
and I_7764 (I134713,I134705,I321628);
nand I_7765 (I134730,I134705,I321628);
nand I_7766 (I134517,I134679,I134730);
DFFARX1 I_7767 (I321616,I2683,I134546,I134770,);
nor I_7768 (I134778,I134770,I134713);
DFFARX1 I_7769 (I134778,I2683,I134546,I134511,);
nor I_7770 (I134526,I134770,I134671);
nand I_7771 (I134823,I321616,I321634);
and I_7772 (I134840,I134823,I321619);
DFFARX1 I_7773 (I134840,I2683,I134546,I134866,);
nor I_7774 (I134514,I134866,I134770);
not I_7775 (I134888,I134866);
nor I_7776 (I134905,I134888,I134679);
nor I_7777 (I134922,I134611,I134905);
DFFARX1 I_7778 (I134922,I2683,I134546,I134529,);
nor I_7779 (I134953,I134888,I134770);
nor I_7780 (I134970,I321622,I321634);
nor I_7781 (I134520,I134970,I134953);
not I_7782 (I135001,I134970);
nand I_7783 (I134523,I134730,I135001);
DFFARX1 I_7784 (I134970,I2683,I134546,I134535,);
DFFARX1 I_7785 (I134970,I2683,I134546,I134532,);
not I_7786 (I135090,I2690);
DFFARX1 I_7787 (I211728,I2683,I135090,I135116,);
DFFARX1 I_7788 (I135116,I2683,I135090,I135133,);
not I_7789 (I135082,I135133);
not I_7790 (I135155,I135116);
nand I_7791 (I135172,I211749,I211740);
and I_7792 (I135189,I135172,I211728);
DFFARX1 I_7793 (I135189,I2683,I135090,I135215,);
not I_7794 (I135223,I135215);
DFFARX1 I_7795 (I211734,I2683,I135090,I135249,);
and I_7796 (I135257,I135249,I211731);
nand I_7797 (I135274,I135249,I211731);
nand I_7798 (I135061,I135223,I135274);
DFFARX1 I_7799 (I211725,I2683,I135090,I135314,);
nor I_7800 (I135322,I135314,I135257);
DFFARX1 I_7801 (I135322,I2683,I135090,I135055,);
nor I_7802 (I135070,I135314,I135215);
nand I_7803 (I135367,I211725,I211737);
and I_7804 (I135384,I135367,I211746);
DFFARX1 I_7805 (I135384,I2683,I135090,I135410,);
nor I_7806 (I135058,I135410,I135314);
not I_7807 (I135432,I135410);
nor I_7808 (I135449,I135432,I135223);
nor I_7809 (I135466,I135155,I135449);
DFFARX1 I_7810 (I135466,I2683,I135090,I135073,);
nor I_7811 (I135497,I135432,I135314);
nor I_7812 (I135514,I211743,I211737);
nor I_7813 (I135064,I135514,I135497);
not I_7814 (I135545,I135514);
nand I_7815 (I135067,I135274,I135545);
DFFARX1 I_7816 (I135514,I2683,I135090,I135079,);
DFFARX1 I_7817 (I135514,I2683,I135090,I135076,);
not I_7818 (I135634,I2690);
DFFARX1 I_7819 (I265576,I2683,I135634,I135660,);
DFFARX1 I_7820 (I135660,I2683,I135634,I135677,);
not I_7821 (I135626,I135677);
not I_7822 (I135699,I135660);
nand I_7823 (I135716,I265570,I265567);
and I_7824 (I135733,I135716,I265582);
DFFARX1 I_7825 (I135733,I2683,I135634,I135759,);
not I_7826 (I135767,I135759);
DFFARX1 I_7827 (I265570,I2683,I135634,I135793,);
and I_7828 (I135801,I135793,I265564);
nand I_7829 (I135818,I135793,I265564);
nand I_7830 (I135605,I135767,I135818);
DFFARX1 I_7831 (I265564,I2683,I135634,I135858,);
nor I_7832 (I135866,I135858,I135801);
DFFARX1 I_7833 (I135866,I2683,I135634,I135599,);
nor I_7834 (I135614,I135858,I135759);
nand I_7835 (I135911,I265579,I265573);
and I_7836 (I135928,I135911,I265567);
DFFARX1 I_7837 (I135928,I2683,I135634,I135954,);
nor I_7838 (I135602,I135954,I135858);
not I_7839 (I135976,I135954);
nor I_7840 (I135993,I135976,I135767);
nor I_7841 (I136010,I135699,I135993);
DFFARX1 I_7842 (I136010,I2683,I135634,I135617,);
nor I_7843 (I136041,I135976,I135858);
nor I_7844 (I136058,I265585,I265573);
nor I_7845 (I135608,I136058,I136041);
not I_7846 (I136089,I136058);
nand I_7847 (I135611,I135818,I136089);
DFFARX1 I_7848 (I136058,I2683,I135634,I135623,);
DFFARX1 I_7849 (I136058,I2683,I135634,I135620,);
not I_7850 (I136178,I2690);
DFFARX1 I_7851 (I196700,I2683,I136178,I136204,);
DFFARX1 I_7852 (I136204,I2683,I136178,I136221,);
not I_7853 (I136170,I136221);
not I_7854 (I136243,I136204);
nand I_7855 (I136260,I196721,I196712);
and I_7856 (I136277,I136260,I196700);
DFFARX1 I_7857 (I136277,I2683,I136178,I136303,);
not I_7858 (I136311,I136303);
DFFARX1 I_7859 (I196706,I2683,I136178,I136337,);
and I_7860 (I136345,I136337,I196703);
nand I_7861 (I136362,I136337,I196703);
nand I_7862 (I136149,I136311,I136362);
DFFARX1 I_7863 (I196697,I2683,I136178,I136402,);
nor I_7864 (I136410,I136402,I136345);
DFFARX1 I_7865 (I136410,I2683,I136178,I136143,);
nor I_7866 (I136158,I136402,I136303);
nand I_7867 (I136455,I196697,I196709);
and I_7868 (I136472,I136455,I196718);
DFFARX1 I_7869 (I136472,I2683,I136178,I136498,);
nor I_7870 (I136146,I136498,I136402);
not I_7871 (I136520,I136498);
nor I_7872 (I136537,I136520,I136311);
nor I_7873 (I136554,I136243,I136537);
DFFARX1 I_7874 (I136554,I2683,I136178,I136161,);
nor I_7875 (I136585,I136520,I136402);
nor I_7876 (I136602,I196715,I196709);
nor I_7877 (I136152,I136602,I136585);
not I_7878 (I136633,I136602);
nand I_7879 (I136155,I136362,I136633);
DFFARX1 I_7880 (I136602,I2683,I136178,I136167,);
DFFARX1 I_7881 (I136602,I2683,I136178,I136164,);
not I_7882 (I136722,I2690);
DFFARX1 I_7883 (I347558,I2683,I136722,I136748,);
DFFARX1 I_7884 (I136748,I2683,I136722,I136765,);
not I_7885 (I136714,I136765);
not I_7886 (I136787,I136748);
nand I_7887 (I136804,I347570,I347558);
and I_7888 (I136821,I136804,I347561);
DFFARX1 I_7889 (I136821,I2683,I136722,I136847,);
not I_7890 (I136855,I136847);
DFFARX1 I_7891 (I347579,I2683,I136722,I136881,);
and I_7892 (I136889,I136881,I347555);
nand I_7893 (I136906,I136881,I347555);
nand I_7894 (I136693,I136855,I136906);
DFFARX1 I_7895 (I347573,I2683,I136722,I136946,);
nor I_7896 (I136954,I136946,I136889);
DFFARX1 I_7897 (I136954,I2683,I136722,I136687,);
nor I_7898 (I136702,I136946,I136847);
nand I_7899 (I136999,I347567,I347564);
and I_7900 (I137016,I136999,I347576);
DFFARX1 I_7901 (I137016,I2683,I136722,I137042,);
nor I_7902 (I136690,I137042,I136946);
not I_7903 (I137064,I137042);
nor I_7904 (I137081,I137064,I136855);
nor I_7905 (I137098,I136787,I137081);
DFFARX1 I_7906 (I137098,I2683,I136722,I136705,);
nor I_7907 (I137129,I137064,I136946);
nor I_7908 (I137146,I347555,I347564);
nor I_7909 (I136696,I137146,I137129);
not I_7910 (I137177,I137146);
nand I_7911 (I136699,I136906,I137177);
DFFARX1 I_7912 (I137146,I2683,I136722,I136711,);
DFFARX1 I_7913 (I137146,I2683,I136722,I136708,);
not I_7914 (I137266,I2690);
DFFARX1 I_7915 (I107417,I2683,I137266,I137292,);
DFFARX1 I_7916 (I137292,I2683,I137266,I137309,);
not I_7917 (I137258,I137309);
not I_7918 (I137331,I137292);
nand I_7919 (I137348,I107396,I107420);
and I_7920 (I137365,I137348,I107423);
DFFARX1 I_7921 (I137365,I2683,I137266,I137391,);
not I_7922 (I137399,I137391);
DFFARX1 I_7923 (I107405,I2683,I137266,I137425,);
and I_7924 (I137433,I137425,I107411);
nand I_7925 (I137450,I137425,I107411);
nand I_7926 (I137237,I137399,I137450);
DFFARX1 I_7927 (I107399,I2683,I137266,I137490,);
nor I_7928 (I137498,I137490,I137433);
DFFARX1 I_7929 (I137498,I2683,I137266,I137231,);
nor I_7930 (I137246,I137490,I137391);
nand I_7931 (I137543,I107408,I107396);
and I_7932 (I137560,I137543,I107402);
DFFARX1 I_7933 (I137560,I2683,I137266,I137586,);
nor I_7934 (I137234,I137586,I137490);
not I_7935 (I137608,I137586);
nor I_7936 (I137625,I137608,I137399);
nor I_7937 (I137642,I137331,I137625);
DFFARX1 I_7938 (I137642,I2683,I137266,I137249,);
nor I_7939 (I137673,I137608,I137490);
nor I_7940 (I137690,I107414,I107396);
nor I_7941 (I137240,I137690,I137673);
not I_7942 (I137721,I137690);
nand I_7943 (I137243,I137450,I137721);
DFFARX1 I_7944 (I137690,I2683,I137266,I137255,);
DFFARX1 I_7945 (I137690,I2683,I137266,I137252,);
not I_7946 (I137810,I2690);
DFFARX1 I_7947 (I174158,I2683,I137810,I137836,);
DFFARX1 I_7948 (I137836,I2683,I137810,I137853,);
not I_7949 (I137802,I137853);
not I_7950 (I137875,I137836);
nand I_7951 (I137892,I174155,I174176);
and I_7952 (I137909,I137892,I174179);
DFFARX1 I_7953 (I137909,I2683,I137810,I137935,);
not I_7954 (I137943,I137935);
DFFARX1 I_7955 (I174164,I2683,I137810,I137969,);
and I_7956 (I137977,I137969,I174167);
nand I_7957 (I137994,I137969,I174167);
nand I_7958 (I137781,I137943,I137994);
DFFARX1 I_7959 (I174170,I2683,I137810,I138034,);
nor I_7960 (I138042,I138034,I137977);
DFFARX1 I_7961 (I138042,I2683,I137810,I137775,);
nor I_7962 (I137790,I138034,I137935);
nand I_7963 (I138087,I174155,I174161);
and I_7964 (I138104,I138087,I174173);
DFFARX1 I_7965 (I138104,I2683,I137810,I138130,);
nor I_7966 (I137778,I138130,I138034);
not I_7967 (I138152,I138130);
nor I_7968 (I138169,I138152,I137943);
nor I_7969 (I138186,I137875,I138169);
DFFARX1 I_7970 (I138186,I2683,I137810,I137793,);
nor I_7971 (I138217,I138152,I138034);
nor I_7972 (I138234,I174158,I174161);
nor I_7973 (I137784,I138234,I138217);
not I_7974 (I138265,I138234);
nand I_7975 (I137787,I137994,I138265);
DFFARX1 I_7976 (I138234,I2683,I137810,I137799,);
DFFARX1 I_7977 (I138234,I2683,I137810,I137796,);
not I_7978 (I138354,I2690);
DFFARX1 I_7979 (I200168,I2683,I138354,I138380,);
DFFARX1 I_7980 (I138380,I2683,I138354,I138397,);
not I_7981 (I138346,I138397);
not I_7982 (I138419,I138380);
nand I_7983 (I138436,I200189,I200180);
and I_7984 (I138453,I138436,I200168);
DFFARX1 I_7985 (I138453,I2683,I138354,I138479,);
not I_7986 (I138487,I138479);
DFFARX1 I_7987 (I200174,I2683,I138354,I138513,);
and I_7988 (I138521,I138513,I200171);
nand I_7989 (I138538,I138513,I200171);
nand I_7990 (I138325,I138487,I138538);
DFFARX1 I_7991 (I200165,I2683,I138354,I138578,);
nor I_7992 (I138586,I138578,I138521);
DFFARX1 I_7993 (I138586,I2683,I138354,I138319,);
nor I_7994 (I138334,I138578,I138479);
nand I_7995 (I138631,I200165,I200177);
and I_7996 (I138648,I138631,I200186);
DFFARX1 I_7997 (I138648,I2683,I138354,I138674,);
nor I_7998 (I138322,I138674,I138578);
not I_7999 (I138696,I138674);
nor I_8000 (I138713,I138696,I138487);
nor I_8001 (I138730,I138419,I138713);
DFFARX1 I_8002 (I138730,I2683,I138354,I138337,);
nor I_8003 (I138761,I138696,I138578);
nor I_8004 (I138778,I200183,I200177);
nor I_8005 (I138328,I138778,I138761);
not I_8006 (I138809,I138778);
nand I_8007 (I138331,I138538,I138809);
DFFARX1 I_8008 (I138778,I2683,I138354,I138343,);
DFFARX1 I_8009 (I138778,I2683,I138354,I138340,);
not I_8010 (I138898,I2690);
DFFARX1 I_8011 (I208838,I2683,I138898,I138924,);
DFFARX1 I_8012 (I138924,I2683,I138898,I138941,);
not I_8013 (I138890,I138941);
not I_8014 (I138963,I138924);
nand I_8015 (I138980,I208859,I208850);
and I_8016 (I138997,I138980,I208838);
DFFARX1 I_8017 (I138997,I2683,I138898,I139023,);
not I_8018 (I139031,I139023);
DFFARX1 I_8019 (I208844,I2683,I138898,I139057,);
and I_8020 (I139065,I139057,I208841);
nand I_8021 (I139082,I139057,I208841);
nand I_8022 (I138869,I139031,I139082);
DFFARX1 I_8023 (I208835,I2683,I138898,I139122,);
nor I_8024 (I139130,I139122,I139065);
DFFARX1 I_8025 (I139130,I2683,I138898,I138863,);
nor I_8026 (I138878,I139122,I139023);
nand I_8027 (I139175,I208835,I208847);
and I_8028 (I139192,I139175,I208856);
DFFARX1 I_8029 (I139192,I2683,I138898,I139218,);
nor I_8030 (I138866,I139218,I139122);
not I_8031 (I139240,I139218);
nor I_8032 (I139257,I139240,I139031);
nor I_8033 (I139274,I138963,I139257);
DFFARX1 I_8034 (I139274,I2683,I138898,I138881,);
nor I_8035 (I139305,I139240,I139122);
nor I_8036 (I139322,I208853,I208847);
nor I_8037 (I138872,I139322,I139305);
not I_8038 (I139353,I139322);
nand I_8039 (I138875,I139082,I139353);
DFFARX1 I_8040 (I139322,I2683,I138898,I138887,);
DFFARX1 I_8041 (I139322,I2683,I138898,I138884,);
not I_8042 (I139442,I2690);
DFFARX1 I_8043 (I19903,I2683,I139442,I139468,);
DFFARX1 I_8044 (I139468,I2683,I139442,I139485,);
not I_8045 (I139434,I139485);
not I_8046 (I139507,I139468);
nand I_8047 (I139524,I19918,I19897);
and I_8048 (I139541,I139524,I19900);
DFFARX1 I_8049 (I139541,I2683,I139442,I139567,);
not I_8050 (I139575,I139567);
DFFARX1 I_8051 (I19906,I2683,I139442,I139601,);
and I_8052 (I139609,I139601,I19900);
nand I_8053 (I139626,I139601,I19900);
nand I_8054 (I139413,I139575,I139626);
DFFARX1 I_8055 (I19915,I2683,I139442,I139666,);
nor I_8056 (I139674,I139666,I139609);
DFFARX1 I_8057 (I139674,I2683,I139442,I139407,);
nor I_8058 (I139422,I139666,I139567);
nand I_8059 (I139719,I19897,I19912);
and I_8060 (I139736,I139719,I19909);
DFFARX1 I_8061 (I139736,I2683,I139442,I139762,);
nor I_8062 (I139410,I139762,I139666);
not I_8063 (I139784,I139762);
nor I_8064 (I139801,I139784,I139575);
nor I_8065 (I139818,I139507,I139801);
DFFARX1 I_8066 (I139818,I2683,I139442,I139425,);
nor I_8067 (I139849,I139784,I139666);
nor I_8068 (I139866,I19921,I19912);
nor I_8069 (I139416,I139866,I139849);
not I_8070 (I139897,I139866);
nand I_8071 (I139419,I139626,I139897);
DFFARX1 I_8072 (I139866,I2683,I139442,I139431,);
DFFARX1 I_8073 (I139866,I2683,I139442,I139428,);
not I_8074 (I139986,I2690);
DFFARX1 I_8075 (I266103,I2683,I139986,I140012,);
DFFARX1 I_8076 (I140012,I2683,I139986,I140029,);
not I_8077 (I139978,I140029);
not I_8078 (I140051,I140012);
nand I_8079 (I140068,I266097,I266094);
and I_8080 (I140085,I140068,I266109);
DFFARX1 I_8081 (I140085,I2683,I139986,I140111,);
not I_8082 (I140119,I140111);
DFFARX1 I_8083 (I266097,I2683,I139986,I140145,);
and I_8084 (I140153,I140145,I266091);
nand I_8085 (I140170,I140145,I266091);
nand I_8086 (I139957,I140119,I140170);
DFFARX1 I_8087 (I266091,I2683,I139986,I140210,);
nor I_8088 (I140218,I140210,I140153);
DFFARX1 I_8089 (I140218,I2683,I139986,I139951,);
nor I_8090 (I139966,I140210,I140111);
nand I_8091 (I140263,I266106,I266100);
and I_8092 (I140280,I140263,I266094);
DFFARX1 I_8093 (I140280,I2683,I139986,I140306,);
nor I_8094 (I139954,I140306,I140210);
not I_8095 (I140328,I140306);
nor I_8096 (I140345,I140328,I140119);
nor I_8097 (I140362,I140051,I140345);
DFFARX1 I_8098 (I140362,I2683,I139986,I139969,);
nor I_8099 (I140393,I140328,I140210);
nor I_8100 (I140410,I266112,I266100);
nor I_8101 (I139960,I140410,I140393);
not I_8102 (I140441,I140410);
nand I_8103 (I139963,I140170,I140441);
DFFARX1 I_8104 (I140410,I2683,I139986,I139975,);
DFFARX1 I_8105 (I140410,I2683,I139986,I139972,);
not I_8106 (I140530,I2690);
DFFARX1 I_8107 (I312637,I2683,I140530,I140556,);
DFFARX1 I_8108 (I140556,I2683,I140530,I140573,);
not I_8109 (I140522,I140573);
not I_8110 (I140595,I140556);
nand I_8111 (I140612,I312637,I312655);
and I_8112 (I140629,I140612,I312649);
DFFARX1 I_8113 (I140629,I2683,I140530,I140655,);
not I_8114 (I140663,I140655);
DFFARX1 I_8115 (I312643,I2683,I140530,I140689,);
and I_8116 (I140697,I140689,I312652);
nand I_8117 (I140714,I140689,I312652);
nand I_8118 (I140501,I140663,I140714);
DFFARX1 I_8119 (I312640,I2683,I140530,I140754,);
nor I_8120 (I140762,I140754,I140697);
DFFARX1 I_8121 (I140762,I2683,I140530,I140495,);
nor I_8122 (I140510,I140754,I140655);
nand I_8123 (I140807,I312640,I312658);
and I_8124 (I140824,I140807,I312643);
DFFARX1 I_8125 (I140824,I2683,I140530,I140850,);
nor I_8126 (I140498,I140850,I140754);
not I_8127 (I140872,I140850);
nor I_8128 (I140889,I140872,I140663);
nor I_8129 (I140906,I140595,I140889);
DFFARX1 I_8130 (I140906,I2683,I140530,I140513,);
nor I_8131 (I140937,I140872,I140754);
nor I_8132 (I140954,I312646,I312658);
nor I_8133 (I140504,I140954,I140937);
not I_8134 (I140985,I140954);
nand I_8135 (I140507,I140714,I140985);
DFFARX1 I_8136 (I140954,I2683,I140530,I140519,);
DFFARX1 I_8137 (I140954,I2683,I140530,I140516,);
not I_8138 (I141074,I2690);
DFFARX1 I_8139 (I272370,I2683,I141074,I141100,);
DFFARX1 I_8140 (I141100,I2683,I141074,I141117,);
not I_8141 (I141066,I141117);
not I_8142 (I141139,I141100);
nand I_8143 (I141156,I272385,I272373);
and I_8144 (I141173,I141156,I272364);
DFFARX1 I_8145 (I141173,I2683,I141074,I141199,);
not I_8146 (I141207,I141199);
DFFARX1 I_8147 (I272376,I2683,I141074,I141233,);
and I_8148 (I141241,I141233,I272367);
nand I_8149 (I141258,I141233,I272367);
nand I_8150 (I141045,I141207,I141258);
DFFARX1 I_8151 (I272382,I2683,I141074,I141298,);
nor I_8152 (I141306,I141298,I141241);
DFFARX1 I_8153 (I141306,I2683,I141074,I141039,);
nor I_8154 (I141054,I141298,I141199);
nand I_8155 (I141351,I272391,I272379);
and I_8156 (I141368,I141351,I272388);
DFFARX1 I_8157 (I141368,I2683,I141074,I141394,);
nor I_8158 (I141042,I141394,I141298);
not I_8159 (I141416,I141394);
nor I_8160 (I141433,I141416,I141207);
nor I_8161 (I141450,I141139,I141433);
DFFARX1 I_8162 (I141450,I2683,I141074,I141057,);
nor I_8163 (I141481,I141416,I141298);
nor I_8164 (I141498,I272364,I272379);
nor I_8165 (I141048,I141498,I141481);
not I_8166 (I141529,I141498);
nand I_8167 (I141051,I141258,I141529);
DFFARX1 I_8168 (I141498,I2683,I141074,I141063,);
DFFARX1 I_8169 (I141498,I2683,I141074,I141060,);
not I_8170 (I141618,I2690);
DFFARX1 I_8171 (I386537,I2683,I141618,I141644,);
DFFARX1 I_8172 (I141644,I2683,I141618,I141661,);
not I_8173 (I141610,I141661);
not I_8174 (I141683,I141644);
nand I_8175 (I141700,I386534,I386531);
and I_8176 (I141717,I141700,I386519);
DFFARX1 I_8177 (I141717,I2683,I141618,I141743,);
not I_8178 (I141751,I141743);
DFFARX1 I_8179 (I386543,I2683,I141618,I141777,);
and I_8180 (I141785,I141777,I386528);
nand I_8181 (I141802,I141777,I386528);
nand I_8182 (I141589,I141751,I141802);
DFFARX1 I_8183 (I386522,I2683,I141618,I141842,);
nor I_8184 (I141850,I141842,I141785);
DFFARX1 I_8185 (I141850,I2683,I141618,I141583,);
nor I_8186 (I141598,I141842,I141743);
nand I_8187 (I141895,I386519,I386525);
and I_8188 (I141912,I141895,I386540);
DFFARX1 I_8189 (I141912,I2683,I141618,I141938,);
nor I_8190 (I141586,I141938,I141842);
not I_8191 (I141960,I141938);
nor I_8192 (I141977,I141960,I141751);
nor I_8193 (I141994,I141683,I141977);
DFFARX1 I_8194 (I141994,I2683,I141618,I141601,);
nor I_8195 (I142025,I141960,I141842);
nor I_8196 (I142042,I386522,I386525);
nor I_8197 (I141592,I142042,I142025);
not I_8198 (I142073,I142042);
nand I_8199 (I141595,I141802,I142073);
DFFARX1 I_8200 (I142042,I2683,I141618,I141607,);
DFFARX1 I_8201 (I142042,I2683,I141618,I141604,);
not I_8202 (I142162,I2690);
DFFARX1 I_8203 (I75088,I2683,I142162,I142188,);
DFFARX1 I_8204 (I142188,I2683,I142162,I142205,);
not I_8205 (I142154,I142205);
not I_8206 (I142227,I142188);
nand I_8207 (I142244,I75100,I75079);
and I_8208 (I142261,I142244,I75082);
DFFARX1 I_8209 (I142261,I2683,I142162,I142287,);
not I_8210 (I142295,I142287);
DFFARX1 I_8211 (I75091,I2683,I142162,I142321,);
and I_8212 (I142329,I142321,I75103);
nand I_8213 (I142346,I142321,I75103);
nand I_8214 (I142133,I142295,I142346);
DFFARX1 I_8215 (I75097,I2683,I142162,I142386,);
nor I_8216 (I142394,I142386,I142329);
DFFARX1 I_8217 (I142394,I2683,I142162,I142127,);
nor I_8218 (I142142,I142386,I142287);
nand I_8219 (I142439,I75085,I75082);
and I_8220 (I142456,I142439,I75094);
DFFARX1 I_8221 (I142456,I2683,I142162,I142482,);
nor I_8222 (I142130,I142482,I142386);
not I_8223 (I142504,I142482);
nor I_8224 (I142521,I142504,I142295);
nor I_8225 (I142538,I142227,I142521);
DFFARX1 I_8226 (I142538,I2683,I142162,I142145,);
nor I_8227 (I142569,I142504,I142386);
nor I_8228 (I142586,I75079,I75082);
nor I_8229 (I142136,I142586,I142569);
not I_8230 (I142617,I142586);
nand I_8231 (I142139,I142346,I142617);
DFFARX1 I_8232 (I142586,I2683,I142162,I142151,);
DFFARX1 I_8233 (I142586,I2683,I142162,I142148,);
not I_8234 (I142706,I2690);
DFFARX1 I_8235 (I176470,I2683,I142706,I142732,);
DFFARX1 I_8236 (I142732,I2683,I142706,I142749,);
not I_8237 (I142698,I142749);
not I_8238 (I142771,I142732);
nand I_8239 (I142788,I176467,I176488);
and I_8240 (I142805,I142788,I176491);
DFFARX1 I_8241 (I142805,I2683,I142706,I142831,);
not I_8242 (I142839,I142831);
DFFARX1 I_8243 (I176476,I2683,I142706,I142865,);
and I_8244 (I142873,I142865,I176479);
nand I_8245 (I142890,I142865,I176479);
nand I_8246 (I142677,I142839,I142890);
DFFARX1 I_8247 (I176482,I2683,I142706,I142930,);
nor I_8248 (I142938,I142930,I142873);
DFFARX1 I_8249 (I142938,I2683,I142706,I142671,);
nor I_8250 (I142686,I142930,I142831);
nand I_8251 (I142983,I176467,I176473);
and I_8252 (I143000,I142983,I176485);
DFFARX1 I_8253 (I143000,I2683,I142706,I143026,);
nor I_8254 (I142674,I143026,I142930);
not I_8255 (I143048,I143026);
nor I_8256 (I143065,I143048,I142839);
nor I_8257 (I143082,I142771,I143065);
DFFARX1 I_8258 (I143082,I2683,I142706,I142689,);
nor I_8259 (I143113,I143048,I142930);
nor I_8260 (I143130,I176470,I176473);
nor I_8261 (I142680,I143130,I143113);
not I_8262 (I143161,I143130);
nand I_8263 (I142683,I142890,I143161);
DFFARX1 I_8264 (I143130,I2683,I142706,I142695,);
DFFARX1 I_8265 (I143130,I2683,I142706,I142692,);
not I_8266 (I143250,I2690);
DFFARX1 I_8267 (I61998,I2683,I143250,I143276,);
DFFARX1 I_8268 (I143276,I2683,I143250,I143293,);
not I_8269 (I143242,I143293);
not I_8270 (I143315,I143276);
nand I_8271 (I143332,I62010,I61989);
and I_8272 (I143349,I143332,I61992);
DFFARX1 I_8273 (I143349,I2683,I143250,I143375,);
not I_8274 (I143383,I143375);
DFFARX1 I_8275 (I62001,I2683,I143250,I143409,);
and I_8276 (I143417,I143409,I62013);
nand I_8277 (I143434,I143409,I62013);
nand I_8278 (I143221,I143383,I143434);
DFFARX1 I_8279 (I62007,I2683,I143250,I143474,);
nor I_8280 (I143482,I143474,I143417);
DFFARX1 I_8281 (I143482,I2683,I143250,I143215,);
nor I_8282 (I143230,I143474,I143375);
nand I_8283 (I143527,I61995,I61992);
and I_8284 (I143544,I143527,I62004);
DFFARX1 I_8285 (I143544,I2683,I143250,I143570,);
nor I_8286 (I143218,I143570,I143474);
not I_8287 (I143592,I143570);
nor I_8288 (I143609,I143592,I143383);
nor I_8289 (I143626,I143315,I143609);
DFFARX1 I_8290 (I143626,I2683,I143250,I143233,);
nor I_8291 (I143657,I143592,I143474);
nor I_8292 (I143674,I61989,I61992);
nor I_8293 (I143224,I143674,I143657);
not I_8294 (I143705,I143674);
nand I_8295 (I143227,I143434,I143705);
DFFARX1 I_8296 (I143674,I2683,I143250,I143239,);
DFFARX1 I_8297 (I143674,I2683,I143250,I143236,);
not I_8298 (I143794,I2690);
DFFARX1 I_8299 (I212306,I2683,I143794,I143820,);
DFFARX1 I_8300 (I143820,I2683,I143794,I143837,);
not I_8301 (I143786,I143837);
not I_8302 (I143859,I143820);
nand I_8303 (I143876,I212327,I212318);
and I_8304 (I143893,I143876,I212306);
DFFARX1 I_8305 (I143893,I2683,I143794,I143919,);
not I_8306 (I143927,I143919);
DFFARX1 I_8307 (I212312,I2683,I143794,I143953,);
and I_8308 (I143961,I143953,I212309);
nand I_8309 (I143978,I143953,I212309);
nand I_8310 (I143765,I143927,I143978);
DFFARX1 I_8311 (I212303,I2683,I143794,I144018,);
nor I_8312 (I144026,I144018,I143961);
DFFARX1 I_8313 (I144026,I2683,I143794,I143759,);
nor I_8314 (I143774,I144018,I143919);
nand I_8315 (I144071,I212303,I212315);
and I_8316 (I144088,I144071,I212324);
DFFARX1 I_8317 (I144088,I2683,I143794,I144114,);
nor I_8318 (I143762,I144114,I144018);
not I_8319 (I144136,I144114);
nor I_8320 (I144153,I144136,I143927);
nor I_8321 (I144170,I143859,I144153);
DFFARX1 I_8322 (I144170,I2683,I143794,I143777,);
nor I_8323 (I144201,I144136,I144018);
nor I_8324 (I144218,I212321,I212315);
nor I_8325 (I143768,I144218,I144201);
not I_8326 (I144249,I144218);
nand I_8327 (I143771,I143978,I144249);
DFFARX1 I_8328 (I144218,I2683,I143794,I143783,);
DFFARX1 I_8329 (I144218,I2683,I143794,I143780,);
not I_8330 (I144338,I2690);
DFFARX1 I_8331 (I419441,I2683,I144338,I144364,);
DFFARX1 I_8332 (I144364,I2683,I144338,I144381,);
not I_8333 (I144330,I144381);
not I_8334 (I144403,I144364);
nand I_8335 (I144420,I419417,I419438);
and I_8336 (I144437,I144420,I419435);
DFFARX1 I_8337 (I144437,I2683,I144338,I144463,);
not I_8338 (I144471,I144463);
DFFARX1 I_8339 (I419414,I2683,I144338,I144497,);
and I_8340 (I144505,I144497,I419426);
nand I_8341 (I144522,I144497,I419426);
nand I_8342 (I144309,I144471,I144522);
DFFARX1 I_8343 (I419429,I2683,I144338,I144562,);
nor I_8344 (I144570,I144562,I144505);
DFFARX1 I_8345 (I144570,I2683,I144338,I144303,);
nor I_8346 (I144318,I144562,I144463);
nand I_8347 (I144615,I419432,I419420);
and I_8348 (I144632,I144615,I419423);
DFFARX1 I_8349 (I144632,I2683,I144338,I144658,);
nor I_8350 (I144306,I144658,I144562);
not I_8351 (I144680,I144658);
nor I_8352 (I144697,I144680,I144471);
nor I_8353 (I144714,I144403,I144697);
DFFARX1 I_8354 (I144714,I2683,I144338,I144321,);
nor I_8355 (I144745,I144680,I144562);
nor I_8356 (I144762,I419414,I419420);
nor I_8357 (I144312,I144762,I144745);
not I_8358 (I144793,I144762);
nand I_8359 (I144315,I144522,I144793);
DFFARX1 I_8360 (I144762,I2683,I144338,I144327,);
DFFARX1 I_8361 (I144762,I2683,I144338,I144324,);
not I_8362 (I144882,I2690);
DFFARX1 I_8363 (I300794,I2683,I144882,I144908,);
DFFARX1 I_8364 (I144908,I2683,I144882,I144925,);
not I_8365 (I144874,I144925);
not I_8366 (I144947,I144908);
nand I_8367 (I144964,I300809,I300797);
and I_8368 (I144981,I144964,I300788);
DFFARX1 I_8369 (I144981,I2683,I144882,I145007,);
not I_8370 (I145015,I145007);
DFFARX1 I_8371 (I300800,I2683,I144882,I145041,);
and I_8372 (I145049,I145041,I300791);
nand I_8373 (I145066,I145041,I300791);
nand I_8374 (I144853,I145015,I145066);
DFFARX1 I_8375 (I300806,I2683,I144882,I145106,);
nor I_8376 (I145114,I145106,I145049);
DFFARX1 I_8377 (I145114,I2683,I144882,I144847,);
nor I_8378 (I144862,I145106,I145007);
nand I_8379 (I145159,I300815,I300803);
and I_8380 (I145176,I145159,I300812);
DFFARX1 I_8381 (I145176,I2683,I144882,I145202,);
nor I_8382 (I144850,I145202,I145106);
not I_8383 (I145224,I145202);
nor I_8384 (I145241,I145224,I145015);
nor I_8385 (I145258,I144947,I145241);
DFFARX1 I_8386 (I145258,I2683,I144882,I144865,);
nor I_8387 (I145289,I145224,I145106);
nor I_8388 (I145306,I300788,I300803);
nor I_8389 (I144856,I145306,I145289);
not I_8390 (I145337,I145306);
nand I_8391 (I144859,I145066,I145337);
DFFARX1 I_8392 (I145306,I2683,I144882,I144871,);
DFFARX1 I_8393 (I145306,I2683,I144882,I144868,);
not I_8394 (I145426,I2690);
DFFARX1 I_8395 (I6734,I2683,I145426,I145452,);
DFFARX1 I_8396 (I145452,I2683,I145426,I145469,);
not I_8397 (I145418,I145469);
not I_8398 (I145491,I145452);
nand I_8399 (I145508,I6722,I6737);
and I_8400 (I145525,I145508,I6725);
DFFARX1 I_8401 (I145525,I2683,I145426,I145551,);
not I_8402 (I145559,I145551);
DFFARX1 I_8403 (I6746,I2683,I145426,I145585,);
and I_8404 (I145593,I145585,I6740);
nand I_8405 (I145610,I145585,I6740);
nand I_8406 (I145397,I145559,I145610);
DFFARX1 I_8407 (I6743,I2683,I145426,I145650,);
nor I_8408 (I145658,I145650,I145593);
DFFARX1 I_8409 (I145658,I2683,I145426,I145391,);
nor I_8410 (I145406,I145650,I145551);
nand I_8411 (I145703,I6722,I6725);
and I_8412 (I145720,I145703,I6728);
DFFARX1 I_8413 (I145720,I2683,I145426,I145746,);
nor I_8414 (I145394,I145746,I145650);
not I_8415 (I145768,I145746);
nor I_8416 (I145785,I145768,I145559);
nor I_8417 (I145802,I145491,I145785);
DFFARX1 I_8418 (I145802,I2683,I145426,I145409,);
nor I_8419 (I145833,I145768,I145650);
nor I_8420 (I145850,I6731,I6725);
nor I_8421 (I145400,I145850,I145833);
not I_8422 (I145881,I145850);
nand I_8423 (I145403,I145610,I145881);
DFFARX1 I_8424 (I145850,I2683,I145426,I145415,);
DFFARX1 I_8425 (I145850,I2683,I145426,I145412,);
not I_8426 (I145970,I2690);
DFFARX1 I_8427 (I15693,I2683,I145970,I145996,);
DFFARX1 I_8428 (I145996,I2683,I145970,I146013,);
not I_8429 (I145962,I146013);
not I_8430 (I146035,I145996);
nand I_8431 (I146052,I15681,I15696);
and I_8432 (I146069,I146052,I15684);
DFFARX1 I_8433 (I146069,I2683,I145970,I146095,);
not I_8434 (I146103,I146095);
DFFARX1 I_8435 (I15705,I2683,I145970,I146129,);
and I_8436 (I146137,I146129,I15699);
nand I_8437 (I146154,I146129,I15699);
nand I_8438 (I145941,I146103,I146154);
DFFARX1 I_8439 (I15702,I2683,I145970,I146194,);
nor I_8440 (I146202,I146194,I146137);
DFFARX1 I_8441 (I146202,I2683,I145970,I145935,);
nor I_8442 (I145950,I146194,I146095);
nand I_8443 (I146247,I15681,I15684);
and I_8444 (I146264,I146247,I15687);
DFFARX1 I_8445 (I146264,I2683,I145970,I146290,);
nor I_8446 (I145938,I146290,I146194);
not I_8447 (I146312,I146290);
nor I_8448 (I146329,I146312,I146103);
nor I_8449 (I146346,I146035,I146329);
DFFARX1 I_8450 (I146346,I2683,I145970,I145953,);
nor I_8451 (I146377,I146312,I146194);
nor I_8452 (I146394,I15690,I15684);
nor I_8453 (I145944,I146394,I146377);
not I_8454 (I146425,I146394);
nand I_8455 (I145947,I146154,I146425);
DFFARX1 I_8456 (I146394,I2683,I145970,I145959,);
DFFARX1 I_8457 (I146394,I2683,I145970,I145956,);
not I_8458 (I146514,I2690);
DFFARX1 I_8459 (I345824,I2683,I146514,I146540,);
DFFARX1 I_8460 (I146540,I2683,I146514,I146557,);
not I_8461 (I146506,I146557);
not I_8462 (I146579,I146540);
nand I_8463 (I146596,I345836,I345824);
and I_8464 (I146613,I146596,I345827);
DFFARX1 I_8465 (I146613,I2683,I146514,I146639,);
not I_8466 (I146647,I146639);
DFFARX1 I_8467 (I345845,I2683,I146514,I146673,);
and I_8468 (I146681,I146673,I345821);
nand I_8469 (I146698,I146673,I345821);
nand I_8470 (I146485,I146647,I146698);
DFFARX1 I_8471 (I345839,I2683,I146514,I146738,);
nor I_8472 (I146746,I146738,I146681);
DFFARX1 I_8473 (I146746,I2683,I146514,I146479,);
nor I_8474 (I146494,I146738,I146639);
nand I_8475 (I146791,I345833,I345830);
and I_8476 (I146808,I146791,I345842);
DFFARX1 I_8477 (I146808,I2683,I146514,I146834,);
nor I_8478 (I146482,I146834,I146738);
not I_8479 (I146856,I146834);
nor I_8480 (I146873,I146856,I146647);
nor I_8481 (I146890,I146579,I146873);
DFFARX1 I_8482 (I146890,I2683,I146514,I146497,);
nor I_8483 (I146921,I146856,I146738);
nor I_8484 (I146938,I345821,I345830);
nor I_8485 (I146488,I146938,I146921);
not I_8486 (I146969,I146938);
nand I_8487 (I146491,I146698,I146969);
DFFARX1 I_8488 (I146938,I2683,I146514,I146503,);
DFFARX1 I_8489 (I146938,I2683,I146514,I146500,);
not I_8490 (I147058,I2690);
DFFARX1 I_8491 (I287228,I2683,I147058,I147084,);
DFFARX1 I_8492 (I147084,I2683,I147058,I147101,);
not I_8493 (I147050,I147101);
not I_8494 (I147123,I147084);
nand I_8495 (I147140,I287243,I287231);
and I_8496 (I147157,I147140,I287222);
DFFARX1 I_8497 (I147157,I2683,I147058,I147183,);
not I_8498 (I147191,I147183);
DFFARX1 I_8499 (I287234,I2683,I147058,I147217,);
and I_8500 (I147225,I147217,I287225);
nand I_8501 (I147242,I147217,I287225);
nand I_8502 (I147029,I147191,I147242);
DFFARX1 I_8503 (I287240,I2683,I147058,I147282,);
nor I_8504 (I147290,I147282,I147225);
DFFARX1 I_8505 (I147290,I2683,I147058,I147023,);
nor I_8506 (I147038,I147282,I147183);
nand I_8507 (I147335,I287249,I287237);
and I_8508 (I147352,I147335,I287246);
DFFARX1 I_8509 (I147352,I2683,I147058,I147378,);
nor I_8510 (I147026,I147378,I147282);
not I_8511 (I147400,I147378);
nor I_8512 (I147417,I147400,I147191);
nor I_8513 (I147434,I147123,I147417);
DFFARX1 I_8514 (I147434,I2683,I147058,I147041,);
nor I_8515 (I147465,I147400,I147282);
nor I_8516 (I147482,I287222,I287237);
nor I_8517 (I147032,I147482,I147465);
not I_8518 (I147513,I147482);
nand I_8519 (I147035,I147242,I147513);
DFFARX1 I_8520 (I147482,I2683,I147058,I147047,);
DFFARX1 I_8521 (I147482,I2683,I147058,I147044,);
not I_8522 (I147602,I2690);
DFFARX1 I_8523 (I414681,I2683,I147602,I147628,);
DFFARX1 I_8524 (I147628,I2683,I147602,I147645,);
not I_8525 (I147594,I147645);
not I_8526 (I147667,I147628);
nand I_8527 (I147684,I414657,I414678);
and I_8528 (I147701,I147684,I414675);
DFFARX1 I_8529 (I147701,I2683,I147602,I147727,);
not I_8530 (I147735,I147727);
DFFARX1 I_8531 (I414654,I2683,I147602,I147761,);
and I_8532 (I147769,I147761,I414666);
nand I_8533 (I147786,I147761,I414666);
nand I_8534 (I147573,I147735,I147786);
DFFARX1 I_8535 (I414669,I2683,I147602,I147826,);
nor I_8536 (I147834,I147826,I147769);
DFFARX1 I_8537 (I147834,I2683,I147602,I147567,);
nor I_8538 (I147582,I147826,I147727);
nand I_8539 (I147879,I414672,I414660);
and I_8540 (I147896,I147879,I414663);
DFFARX1 I_8541 (I147896,I2683,I147602,I147922,);
nor I_8542 (I147570,I147922,I147826);
not I_8543 (I147944,I147922);
nor I_8544 (I147961,I147944,I147735);
nor I_8545 (I147978,I147667,I147961);
DFFARX1 I_8546 (I147978,I2683,I147602,I147585,);
nor I_8547 (I148009,I147944,I147826);
nor I_8548 (I148026,I414654,I414660);
nor I_8549 (I147576,I148026,I148009);
not I_8550 (I148057,I148026);
nand I_8551 (I147579,I147786,I148057);
DFFARX1 I_8552 (I148026,I2683,I147602,I147591,);
DFFARX1 I_8553 (I148026,I2683,I147602,I147588,);
not I_8554 (I148146,I2690);
DFFARX1 I_8555 (I344668,I2683,I148146,I148172,);
DFFARX1 I_8556 (I148172,I2683,I148146,I148189,);
not I_8557 (I148138,I148189);
not I_8558 (I148211,I148172);
nand I_8559 (I148228,I344680,I344668);
and I_8560 (I148245,I148228,I344671);
DFFARX1 I_8561 (I148245,I2683,I148146,I148271,);
not I_8562 (I148279,I148271);
DFFARX1 I_8563 (I344689,I2683,I148146,I148305,);
and I_8564 (I148313,I148305,I344665);
nand I_8565 (I148330,I148305,I344665);
nand I_8566 (I148117,I148279,I148330);
DFFARX1 I_8567 (I344683,I2683,I148146,I148370,);
nor I_8568 (I148378,I148370,I148313);
DFFARX1 I_8569 (I148378,I2683,I148146,I148111,);
nor I_8570 (I148126,I148370,I148271);
nand I_8571 (I148423,I344677,I344674);
and I_8572 (I148440,I148423,I344686);
DFFARX1 I_8573 (I148440,I2683,I148146,I148466,);
nor I_8574 (I148114,I148466,I148370);
not I_8575 (I148488,I148466);
nor I_8576 (I148505,I148488,I148279);
nor I_8577 (I148522,I148211,I148505);
DFFARX1 I_8578 (I148522,I2683,I148146,I148129,);
nor I_8579 (I148553,I148488,I148370);
nor I_8580 (I148570,I344665,I344674);
nor I_8581 (I148120,I148570,I148553);
not I_8582 (I148601,I148570);
nand I_8583 (I148123,I148330,I148601);
DFFARX1 I_8584 (I148570,I2683,I148146,I148135,);
DFFARX1 I_8585 (I148570,I2683,I148146,I148132,);
not I_8586 (I148690,I2690);
DFFARX1 I_8587 (I304670,I2683,I148690,I148716,);
DFFARX1 I_8588 (I148716,I2683,I148690,I148733,);
not I_8589 (I148682,I148733);
not I_8590 (I148755,I148716);
nand I_8591 (I148772,I304685,I304673);
and I_8592 (I148789,I148772,I304664);
DFFARX1 I_8593 (I148789,I2683,I148690,I148815,);
not I_8594 (I148823,I148815);
DFFARX1 I_8595 (I304676,I2683,I148690,I148849,);
and I_8596 (I148857,I148849,I304667);
nand I_8597 (I148874,I148849,I304667);
nand I_8598 (I148661,I148823,I148874);
DFFARX1 I_8599 (I304682,I2683,I148690,I148914,);
nor I_8600 (I148922,I148914,I148857);
DFFARX1 I_8601 (I148922,I2683,I148690,I148655,);
nor I_8602 (I148670,I148914,I148815);
nand I_8603 (I148967,I304691,I304679);
and I_8604 (I148984,I148967,I304688);
DFFARX1 I_8605 (I148984,I2683,I148690,I149010,);
nor I_8606 (I148658,I149010,I148914);
not I_8607 (I149032,I149010);
nor I_8608 (I149049,I149032,I148823);
nor I_8609 (I149066,I148755,I149049);
DFFARX1 I_8610 (I149066,I2683,I148690,I148673,);
nor I_8611 (I149097,I149032,I148914);
nor I_8612 (I149114,I304664,I304679);
nor I_8613 (I148664,I149114,I149097);
not I_8614 (I149145,I149114);
nand I_8615 (I148667,I148874,I149145);
DFFARX1 I_8616 (I149114,I2683,I148690,I148679,);
DFFARX1 I_8617 (I149114,I2683,I148690,I148676,);
not I_8618 (I149234,I2690);
DFFARX1 I_8619 (I267157,I2683,I149234,I149260,);
DFFARX1 I_8620 (I149260,I2683,I149234,I149277,);
not I_8621 (I149226,I149277);
not I_8622 (I149299,I149260);
nand I_8623 (I149316,I267151,I267148);
and I_8624 (I149333,I149316,I267163);
DFFARX1 I_8625 (I149333,I2683,I149234,I149359,);
not I_8626 (I149367,I149359);
DFFARX1 I_8627 (I267151,I2683,I149234,I149393,);
and I_8628 (I149401,I149393,I267145);
nand I_8629 (I149418,I149393,I267145);
nand I_8630 (I149205,I149367,I149418);
DFFARX1 I_8631 (I267145,I2683,I149234,I149458,);
nor I_8632 (I149466,I149458,I149401);
DFFARX1 I_8633 (I149466,I2683,I149234,I149199,);
nor I_8634 (I149214,I149458,I149359);
nand I_8635 (I149511,I267160,I267154);
and I_8636 (I149528,I149511,I267148);
DFFARX1 I_8637 (I149528,I2683,I149234,I149554,);
nor I_8638 (I149202,I149554,I149458);
not I_8639 (I149576,I149554);
nor I_8640 (I149593,I149576,I149367);
nor I_8641 (I149610,I149299,I149593);
DFFARX1 I_8642 (I149610,I2683,I149234,I149217,);
nor I_8643 (I149641,I149576,I149458);
nor I_8644 (I149658,I267166,I267154);
nor I_8645 (I149208,I149658,I149641);
not I_8646 (I149689,I149658);
nand I_8647 (I149211,I149418,I149689);
DFFARX1 I_8648 (I149658,I2683,I149234,I149223,);
DFFARX1 I_8649 (I149658,I2683,I149234,I149220,);
not I_8650 (I149778,I2690);
DFFARX1 I_8651 (I268738,I2683,I149778,I149804,);
DFFARX1 I_8652 (I149804,I2683,I149778,I149821,);
not I_8653 (I149770,I149821);
not I_8654 (I149843,I149804);
nand I_8655 (I149860,I268732,I268729);
and I_8656 (I149877,I149860,I268744);
DFFARX1 I_8657 (I149877,I2683,I149778,I149903,);
not I_8658 (I149911,I149903);
DFFARX1 I_8659 (I268732,I2683,I149778,I149937,);
and I_8660 (I149945,I149937,I268726);
nand I_8661 (I149962,I149937,I268726);
nand I_8662 (I149749,I149911,I149962);
DFFARX1 I_8663 (I268726,I2683,I149778,I150002,);
nor I_8664 (I150010,I150002,I149945);
DFFARX1 I_8665 (I150010,I2683,I149778,I149743,);
nor I_8666 (I149758,I150002,I149903);
nand I_8667 (I150055,I268741,I268735);
and I_8668 (I150072,I150055,I268729);
DFFARX1 I_8669 (I150072,I2683,I149778,I150098,);
nor I_8670 (I149746,I150098,I150002);
not I_8671 (I150120,I150098);
nor I_8672 (I150137,I150120,I149911);
nor I_8673 (I150154,I149843,I150137);
DFFARX1 I_8674 (I150154,I2683,I149778,I149761,);
nor I_8675 (I150185,I150120,I150002);
nor I_8676 (I150202,I268747,I268735);
nor I_8677 (I149752,I150202,I150185);
not I_8678 (I150233,I150202);
nand I_8679 (I149755,I149962,I150233);
DFFARX1 I_8680 (I150202,I2683,I149778,I149767,);
DFFARX1 I_8681 (I150202,I2683,I149778,I149764,);
not I_8682 (I150322,I2690);
DFFARX1 I_8683 (I260833,I2683,I150322,I150348,);
DFFARX1 I_8684 (I150348,I2683,I150322,I150365,);
not I_8685 (I150314,I150365);
not I_8686 (I150387,I150348);
nand I_8687 (I150404,I260827,I260824);
and I_8688 (I150421,I150404,I260839);
DFFARX1 I_8689 (I150421,I2683,I150322,I150447,);
not I_8690 (I150455,I150447);
DFFARX1 I_8691 (I260827,I2683,I150322,I150481,);
and I_8692 (I150489,I150481,I260821);
nand I_8693 (I150506,I150481,I260821);
nand I_8694 (I150293,I150455,I150506);
DFFARX1 I_8695 (I260821,I2683,I150322,I150546,);
nor I_8696 (I150554,I150546,I150489);
DFFARX1 I_8697 (I150554,I2683,I150322,I150287,);
nor I_8698 (I150302,I150546,I150447);
nand I_8699 (I150599,I260836,I260830);
and I_8700 (I150616,I150599,I260824);
DFFARX1 I_8701 (I150616,I2683,I150322,I150642,);
nor I_8702 (I150290,I150642,I150546);
not I_8703 (I150664,I150642);
nor I_8704 (I150681,I150664,I150455);
nor I_8705 (I150698,I150387,I150681);
DFFARX1 I_8706 (I150698,I2683,I150322,I150305,);
nor I_8707 (I150729,I150664,I150546);
nor I_8708 (I150746,I260842,I260830);
nor I_8709 (I150296,I150746,I150729);
not I_8710 (I150777,I150746);
nand I_8711 (I150299,I150506,I150777);
DFFARX1 I_8712 (I150746,I2683,I150322,I150311,);
DFFARX1 I_8713 (I150746,I2683,I150322,I150308,);
not I_8714 (I150866,I2690);
DFFARX1 I_8715 (I278830,I2683,I150866,I150892,);
DFFARX1 I_8716 (I150892,I2683,I150866,I150909,);
not I_8717 (I150858,I150909);
not I_8718 (I150931,I150892);
nand I_8719 (I150948,I278845,I278833);
and I_8720 (I150965,I150948,I278824);
DFFARX1 I_8721 (I150965,I2683,I150866,I150991,);
not I_8722 (I150999,I150991);
DFFARX1 I_8723 (I278836,I2683,I150866,I151025,);
and I_8724 (I151033,I151025,I278827);
nand I_8725 (I151050,I151025,I278827);
nand I_8726 (I150837,I150999,I151050);
DFFARX1 I_8727 (I278842,I2683,I150866,I151090,);
nor I_8728 (I151098,I151090,I151033);
DFFARX1 I_8729 (I151098,I2683,I150866,I150831,);
nor I_8730 (I150846,I151090,I150991);
nand I_8731 (I151143,I278851,I278839);
and I_8732 (I151160,I151143,I278848);
DFFARX1 I_8733 (I151160,I2683,I150866,I151186,);
nor I_8734 (I150834,I151186,I151090);
not I_8735 (I151208,I151186);
nor I_8736 (I151225,I151208,I150999);
nor I_8737 (I151242,I150931,I151225);
DFFARX1 I_8738 (I151242,I2683,I150866,I150849,);
nor I_8739 (I151273,I151208,I151090);
nor I_8740 (I151290,I278824,I278839);
nor I_8741 (I150840,I151290,I151273);
not I_8742 (I151321,I151290);
nand I_8743 (I150843,I151050,I151321);
DFFARX1 I_8744 (I151290,I2683,I150866,I150855,);
DFFARX1 I_8745 (I151290,I2683,I150866,I150852,);
not I_8746 (I151410,I2690);
DFFARX1 I_8747 (I411111,I2683,I151410,I151436,);
DFFARX1 I_8748 (I151436,I2683,I151410,I151453,);
not I_8749 (I151402,I151453);
not I_8750 (I151475,I151436);
nand I_8751 (I151492,I411087,I411108);
and I_8752 (I151509,I151492,I411105);
DFFARX1 I_8753 (I151509,I2683,I151410,I151535,);
not I_8754 (I151543,I151535);
DFFARX1 I_8755 (I411084,I2683,I151410,I151569,);
and I_8756 (I151577,I151569,I411096);
nand I_8757 (I151594,I151569,I411096);
nand I_8758 (I151381,I151543,I151594);
DFFARX1 I_8759 (I411099,I2683,I151410,I151634,);
nor I_8760 (I151642,I151634,I151577);
DFFARX1 I_8761 (I151642,I2683,I151410,I151375,);
nor I_8762 (I151390,I151634,I151535);
nand I_8763 (I151687,I411102,I411090);
and I_8764 (I151704,I151687,I411093);
DFFARX1 I_8765 (I151704,I2683,I151410,I151730,);
nor I_8766 (I151378,I151730,I151634);
not I_8767 (I151752,I151730);
nor I_8768 (I151769,I151752,I151543);
nor I_8769 (I151786,I151475,I151769);
DFFARX1 I_8770 (I151786,I2683,I151410,I151393,);
nor I_8771 (I151817,I151752,I151634);
nor I_8772 (I151834,I411084,I411090);
nor I_8773 (I151384,I151834,I151817);
not I_8774 (I151865,I151834);
nand I_8775 (I151387,I151594,I151865);
DFFARX1 I_8776 (I151834,I2683,I151410,I151399,);
DFFARX1 I_8777 (I151834,I2683,I151410,I151396,);
not I_8778 (I151954,I2690);
DFFARX1 I_8779 (I108998,I2683,I151954,I151980,);
DFFARX1 I_8780 (I151980,I2683,I151954,I151997,);
not I_8781 (I151946,I151997);
not I_8782 (I152019,I151980);
nand I_8783 (I152036,I108977,I109001);
and I_8784 (I152053,I152036,I109004);
DFFARX1 I_8785 (I152053,I2683,I151954,I152079,);
not I_8786 (I152087,I152079);
DFFARX1 I_8787 (I108986,I2683,I151954,I152113,);
and I_8788 (I152121,I152113,I108992);
nand I_8789 (I152138,I152113,I108992);
nand I_8790 (I151925,I152087,I152138);
DFFARX1 I_8791 (I108980,I2683,I151954,I152178,);
nor I_8792 (I152186,I152178,I152121);
DFFARX1 I_8793 (I152186,I2683,I151954,I151919,);
nor I_8794 (I151934,I152178,I152079);
nand I_8795 (I152231,I108989,I108977);
and I_8796 (I152248,I152231,I108983);
DFFARX1 I_8797 (I152248,I2683,I151954,I152274,);
nor I_8798 (I151922,I152274,I152178);
not I_8799 (I152296,I152274);
nor I_8800 (I152313,I152296,I152087);
nor I_8801 (I152330,I152019,I152313);
DFFARX1 I_8802 (I152330,I2683,I151954,I151937,);
nor I_8803 (I152361,I152296,I152178);
nor I_8804 (I152378,I108995,I108977);
nor I_8805 (I151928,I152378,I152361);
not I_8806 (I152409,I152378);
nand I_8807 (I151931,I152138,I152409);
DFFARX1 I_8808 (I152378,I2683,I151954,I151943,);
DFFARX1 I_8809 (I152378,I2683,I151954,I151940,);
not I_8810 (I152498,I2690);
DFFARX1 I_8811 (I181672,I2683,I152498,I152524,);
DFFARX1 I_8812 (I152524,I2683,I152498,I152541,);
not I_8813 (I152490,I152541);
not I_8814 (I152563,I152524);
nand I_8815 (I152580,I181669,I181690);
and I_8816 (I152597,I152580,I181693);
DFFARX1 I_8817 (I152597,I2683,I152498,I152623,);
not I_8818 (I152631,I152623);
DFFARX1 I_8819 (I181678,I2683,I152498,I152657,);
and I_8820 (I152665,I152657,I181681);
nand I_8821 (I152682,I152657,I181681);
nand I_8822 (I152469,I152631,I152682);
DFFARX1 I_8823 (I181684,I2683,I152498,I152722,);
nor I_8824 (I152730,I152722,I152665);
DFFARX1 I_8825 (I152730,I2683,I152498,I152463,);
nor I_8826 (I152478,I152722,I152623);
nand I_8827 (I152775,I181669,I181675);
and I_8828 (I152792,I152775,I181687);
DFFARX1 I_8829 (I152792,I2683,I152498,I152818,);
nor I_8830 (I152466,I152818,I152722);
not I_8831 (I152840,I152818);
nor I_8832 (I152857,I152840,I152631);
nor I_8833 (I152874,I152563,I152857);
DFFARX1 I_8834 (I152874,I2683,I152498,I152481,);
nor I_8835 (I152905,I152840,I152722);
nor I_8836 (I152922,I181672,I181675);
nor I_8837 (I152472,I152922,I152905);
not I_8838 (I152953,I152922);
nand I_8839 (I152475,I152682,I152953);
DFFARX1 I_8840 (I152922,I2683,I152498,I152487,);
DFFARX1 I_8841 (I152922,I2683,I152498,I152484,);
not I_8842 (I153042,I2690);
DFFARX1 I_8843 (I79253,I2683,I153042,I153068,);
DFFARX1 I_8844 (I153068,I2683,I153042,I153085,);
not I_8845 (I153034,I153085);
not I_8846 (I153107,I153068);
nand I_8847 (I153124,I79265,I79244);
and I_8848 (I153141,I153124,I79247);
DFFARX1 I_8849 (I153141,I2683,I153042,I153167,);
not I_8850 (I153175,I153167);
DFFARX1 I_8851 (I79256,I2683,I153042,I153201,);
and I_8852 (I153209,I153201,I79268);
nand I_8853 (I153226,I153201,I79268);
nand I_8854 (I153013,I153175,I153226);
DFFARX1 I_8855 (I79262,I2683,I153042,I153266,);
nor I_8856 (I153274,I153266,I153209);
DFFARX1 I_8857 (I153274,I2683,I153042,I153007,);
nor I_8858 (I153022,I153266,I153167);
nand I_8859 (I153319,I79250,I79247);
and I_8860 (I153336,I153319,I79259);
DFFARX1 I_8861 (I153336,I2683,I153042,I153362,);
nor I_8862 (I153010,I153362,I153266);
not I_8863 (I153384,I153362);
nor I_8864 (I153401,I153384,I153175);
nor I_8865 (I153418,I153107,I153401);
DFFARX1 I_8866 (I153418,I2683,I153042,I153025,);
nor I_8867 (I153449,I153384,I153266);
nor I_8868 (I153466,I79244,I79247);
nor I_8869 (I153016,I153466,I153449);
not I_8870 (I153497,I153466);
nand I_8871 (I153019,I153226,I153497);
DFFARX1 I_8872 (I153466,I2683,I153042,I153031,);
DFFARX1 I_8873 (I153466,I2683,I153042,I153028,);
not I_8874 (I153586,I2690);
DFFARX1 I_8875 (I33078,I2683,I153586,I153612,);
DFFARX1 I_8876 (I153612,I2683,I153586,I153629,);
not I_8877 (I153578,I153629);
not I_8878 (I153651,I153612);
nand I_8879 (I153668,I33093,I33072);
and I_8880 (I153685,I153668,I33075);
DFFARX1 I_8881 (I153685,I2683,I153586,I153711,);
not I_8882 (I153719,I153711);
DFFARX1 I_8883 (I33081,I2683,I153586,I153745,);
and I_8884 (I153753,I153745,I33075);
nand I_8885 (I153770,I153745,I33075);
nand I_8886 (I153557,I153719,I153770);
DFFARX1 I_8887 (I33090,I2683,I153586,I153810,);
nor I_8888 (I153818,I153810,I153753);
DFFARX1 I_8889 (I153818,I2683,I153586,I153551,);
nor I_8890 (I153566,I153810,I153711);
nand I_8891 (I153863,I33072,I33087);
and I_8892 (I153880,I153863,I33084);
DFFARX1 I_8893 (I153880,I2683,I153586,I153906,);
nor I_8894 (I153554,I153906,I153810);
not I_8895 (I153928,I153906);
nor I_8896 (I153945,I153928,I153719);
nor I_8897 (I153962,I153651,I153945);
DFFARX1 I_8898 (I153962,I2683,I153586,I153569,);
nor I_8899 (I153993,I153928,I153810);
nor I_8900 (I154010,I33096,I33087);
nor I_8901 (I153560,I154010,I153993);
not I_8902 (I154041,I154010);
nand I_8903 (I153563,I153770,I154041);
DFFARX1 I_8904 (I154010,I2683,I153586,I153575,);
DFFARX1 I_8905 (I154010,I2683,I153586,I153572,);
not I_8906 (I154130,I2690);
DFFARX1 I_8907 (I356228,I2683,I154130,I154156,);
DFFARX1 I_8908 (I154156,I2683,I154130,I154173,);
not I_8909 (I154122,I154173);
not I_8910 (I154195,I154156);
nand I_8911 (I154212,I356240,I356228);
and I_8912 (I154229,I154212,I356231);
DFFARX1 I_8913 (I154229,I2683,I154130,I154255,);
not I_8914 (I154263,I154255);
DFFARX1 I_8915 (I356249,I2683,I154130,I154289,);
and I_8916 (I154297,I154289,I356225);
nand I_8917 (I154314,I154289,I356225);
nand I_8918 (I154101,I154263,I154314);
DFFARX1 I_8919 (I356243,I2683,I154130,I154354,);
nor I_8920 (I154362,I154354,I154297);
DFFARX1 I_8921 (I154362,I2683,I154130,I154095,);
nor I_8922 (I154110,I154354,I154255);
nand I_8923 (I154407,I356237,I356234);
and I_8924 (I154424,I154407,I356246);
DFFARX1 I_8925 (I154424,I2683,I154130,I154450,);
nor I_8926 (I154098,I154450,I154354);
not I_8927 (I154472,I154450);
nor I_8928 (I154489,I154472,I154263);
nor I_8929 (I154506,I154195,I154489);
DFFARX1 I_8930 (I154506,I2683,I154130,I154113,);
nor I_8931 (I154537,I154472,I154354);
nor I_8932 (I154554,I356225,I356234);
nor I_8933 (I154104,I154554,I154537);
not I_8934 (I154585,I154554);
nand I_8935 (I154107,I154314,I154585);
DFFARX1 I_8936 (I154554,I2683,I154130,I154119,);
DFFARX1 I_8937 (I154554,I2683,I154130,I154116,);
not I_8938 (I154671,I2690);
DFFARX1 I_8939 (I358555,I2683,I154671,I154697,);
DFFARX1 I_8940 (I154697,I2683,I154671,I154714,);
not I_8941 (I154663,I154714);
DFFARX1 I_8942 (I358537,I2683,I154671,I154745,);
not I_8943 (I154753,I358543);
nor I_8944 (I154770,I154697,I154753);
not I_8945 (I154787,I358558);
not I_8946 (I154804,I358549);
nand I_8947 (I154821,I154804,I358558);
nor I_8948 (I154838,I154753,I154821);
nor I_8949 (I154855,I154745,I154838);
DFFARX1 I_8950 (I154804,I2683,I154671,I154660,);
nor I_8951 (I154886,I358549,I358561);
nand I_8952 (I154903,I154886,I358540);
nor I_8953 (I154920,I154903,I154787);
nand I_8954 (I154645,I154920,I358543);
DFFARX1 I_8955 (I154903,I2683,I154671,I154657,);
nand I_8956 (I154965,I154787,I358549);
nor I_8957 (I154982,I154787,I358549);
nand I_8958 (I154651,I154770,I154982);
not I_8959 (I155013,I358546);
nor I_8960 (I155030,I155013,I154965);
DFFARX1 I_8961 (I155030,I2683,I154671,I154639,);
nor I_8962 (I155061,I155013,I358552);
and I_8963 (I155078,I155061,I358537);
or I_8964 (I155095,I155078,I358540);
DFFARX1 I_8965 (I155095,I2683,I154671,I155121,);
nor I_8966 (I155129,I155121,I154745);
nor I_8967 (I154648,I154697,I155129);
not I_8968 (I155160,I155121);
nor I_8969 (I155177,I155160,I154855);
DFFARX1 I_8970 (I155177,I2683,I154671,I154654,);
nand I_8971 (I155208,I155160,I154787);
nor I_8972 (I154642,I155013,I155208);
not I_8973 (I155266,I2690);
DFFARX1 I_8974 (I403349,I2683,I155266,I155292,);
DFFARX1 I_8975 (I155292,I2683,I155266,I155309,);
not I_8976 (I155258,I155309);
DFFARX1 I_8977 (I403355,I2683,I155266,I155340,);
not I_8978 (I155348,I403370);
nor I_8979 (I155365,I155292,I155348);
not I_8980 (I155382,I403361);
not I_8981 (I155399,I403358);
nand I_8982 (I155416,I155399,I403361);
nor I_8983 (I155433,I155348,I155416);
nor I_8984 (I155450,I155340,I155433);
DFFARX1 I_8985 (I155399,I2683,I155266,I155255,);
nor I_8986 (I155481,I403358,I403349);
nand I_8987 (I155498,I155481,I403373);
nor I_8988 (I155515,I155498,I155382);
nand I_8989 (I155240,I155515,I403370);
DFFARX1 I_8990 (I155498,I2683,I155266,I155252,);
nand I_8991 (I155560,I155382,I403358);
nor I_8992 (I155577,I155382,I403358);
nand I_8993 (I155246,I155365,I155577);
not I_8994 (I155608,I403367);
nor I_8995 (I155625,I155608,I155560);
DFFARX1 I_8996 (I155625,I2683,I155266,I155234,);
nor I_8997 (I155656,I155608,I403352);
and I_8998 (I155673,I155656,I403364);
or I_8999 (I155690,I155673,I403376);
DFFARX1 I_9000 (I155690,I2683,I155266,I155716,);
nor I_9001 (I155724,I155716,I155340);
nor I_9002 (I155243,I155292,I155724);
not I_9003 (I155755,I155716);
nor I_9004 (I155772,I155755,I155450);
DFFARX1 I_9005 (I155772,I2683,I155266,I155249,);
nand I_9006 (I155803,I155755,I155382);
nor I_9007 (I155237,I155608,I155803);
not I_9008 (I155861,I2690);
DFFARX1 I_9009 (I72104,I2683,I155861,I155887,);
DFFARX1 I_9010 (I155887,I2683,I155861,I155904,);
not I_9011 (I155853,I155904);
DFFARX1 I_9012 (I72128,I2683,I155861,I155935,);
not I_9013 (I155943,I72122);
nor I_9014 (I155960,I155887,I155943);
not I_9015 (I155977,I72116);
not I_9016 (I155994,I72113);
nand I_9017 (I156011,I155994,I72116);
nor I_9018 (I156028,I155943,I156011);
nor I_9019 (I156045,I155935,I156028);
DFFARX1 I_9020 (I155994,I2683,I155861,I155850,);
nor I_9021 (I156076,I72113,I72107);
nand I_9022 (I156093,I156076,I72125);
nor I_9023 (I156110,I156093,I155977);
nand I_9024 (I155835,I156110,I72122);
DFFARX1 I_9025 (I156093,I2683,I155861,I155847,);
nand I_9026 (I156155,I155977,I72113);
nor I_9027 (I156172,I155977,I72113);
nand I_9028 (I155841,I155960,I156172);
not I_9029 (I156203,I72119);
nor I_9030 (I156220,I156203,I156155);
DFFARX1 I_9031 (I156220,I2683,I155861,I155829,);
nor I_9032 (I156251,I156203,I72104);
and I_9033 (I156268,I156251,I72110);
or I_9034 (I156285,I156268,I72107);
DFFARX1 I_9035 (I156285,I2683,I155861,I156311,);
nor I_9036 (I156319,I156311,I155935);
nor I_9037 (I155838,I155887,I156319);
not I_9038 (I156350,I156311);
nor I_9039 (I156367,I156350,I156045);
DFFARX1 I_9040 (I156367,I2683,I155861,I155844,);
nand I_9041 (I156398,I156350,I155977);
nor I_9042 (I155832,I156203,I156398);
not I_9043 (I156456,I2690);
DFFARX1 I_9044 (I133967,I2683,I156456,I156482,);
DFFARX1 I_9045 (I156482,I2683,I156456,I156499,);
not I_9046 (I156448,I156499);
DFFARX1 I_9047 (I133991,I2683,I156456,I156530,);
not I_9048 (I156538,I133970);
nor I_9049 (I156555,I156482,I156538);
not I_9050 (I156572,I133976);
not I_9051 (I156589,I133982);
nand I_9052 (I156606,I156589,I133976);
nor I_9053 (I156623,I156538,I156606);
nor I_9054 (I156640,I156530,I156623);
DFFARX1 I_9055 (I156589,I2683,I156456,I156445,);
nor I_9056 (I156671,I133982,I133994);
nand I_9057 (I156688,I156671,I133988);
nor I_9058 (I156705,I156688,I156572);
nand I_9059 (I156430,I156705,I133970);
DFFARX1 I_9060 (I156688,I2683,I156456,I156442,);
nand I_9061 (I156750,I156572,I133982);
nor I_9062 (I156767,I156572,I133982);
nand I_9063 (I156436,I156555,I156767);
not I_9064 (I156798,I133973);
nor I_9065 (I156815,I156798,I156750);
DFFARX1 I_9066 (I156815,I2683,I156456,I156424,);
nor I_9067 (I156846,I156798,I133967);
and I_9068 (I156863,I156846,I133985);
or I_9069 (I156880,I156863,I133979);
DFFARX1 I_9070 (I156880,I2683,I156456,I156906,);
nor I_9071 (I156914,I156906,I156530);
nor I_9072 (I156433,I156482,I156914);
not I_9073 (I156945,I156906);
nor I_9074 (I156962,I156945,I156640);
DFFARX1 I_9075 (I156962,I2683,I156456,I156439,);
nand I_9076 (I156993,I156945,I156572);
nor I_9077 (I156427,I156798,I156993);
not I_9078 (I157051,I2690);
DFFARX1 I_9079 (I293051,I2683,I157051,I157077,);
DFFARX1 I_9080 (I157077,I2683,I157051,I157094,);
not I_9081 (I157043,I157094);
DFFARX1 I_9082 (I293039,I2683,I157051,I157125,);
not I_9083 (I157133,I293036);
nor I_9084 (I157150,I157077,I157133);
not I_9085 (I157167,I293048);
not I_9086 (I157184,I293045);
nand I_9087 (I157201,I157184,I293048);
nor I_9088 (I157218,I157133,I157201);
nor I_9089 (I157235,I157125,I157218);
DFFARX1 I_9090 (I157184,I2683,I157051,I157040,);
nor I_9091 (I157266,I293045,I293054);
nand I_9092 (I157283,I157266,I293057);
nor I_9093 (I157300,I157283,I157167);
nand I_9094 (I157025,I157300,I293036);
DFFARX1 I_9095 (I157283,I2683,I157051,I157037,);
nand I_9096 (I157345,I157167,I293045);
nor I_9097 (I157362,I157167,I293045);
nand I_9098 (I157031,I157150,I157362);
not I_9099 (I157393,I293060);
nor I_9100 (I157410,I157393,I157345);
DFFARX1 I_9101 (I157410,I2683,I157051,I157019,);
nor I_9102 (I157441,I157393,I293063);
and I_9103 (I157458,I157441,I293042);
or I_9104 (I157475,I157458,I293036);
DFFARX1 I_9105 (I157475,I2683,I157051,I157501,);
nor I_9106 (I157509,I157501,I157125);
nor I_9107 (I157028,I157077,I157509);
not I_9108 (I157540,I157501);
nor I_9109 (I157557,I157540,I157235);
DFFARX1 I_9110 (I157557,I2683,I157051,I157034,);
nand I_9111 (I157588,I157540,I157167);
nor I_9112 (I157022,I157393,I157588);
not I_9113 (I157646,I2690);
DFFARX1 I_9114 (I371389,I2683,I157646,I157672,);
DFFARX1 I_9115 (I157672,I2683,I157646,I157689,);
not I_9116 (I157638,I157689);
DFFARX1 I_9117 (I371404,I2683,I157646,I157720,);
not I_9118 (I157728,I371413);
nor I_9119 (I157745,I157672,I157728);
not I_9120 (I157762,I371392);
not I_9121 (I157779,I371398);
nand I_9122 (I157796,I157779,I371392);
nor I_9123 (I157813,I157728,I157796);
nor I_9124 (I157830,I157720,I157813);
DFFARX1 I_9125 (I157779,I2683,I157646,I157635,);
nor I_9126 (I157861,I371398,I371410);
nand I_9127 (I157878,I157861,I371407);
nor I_9128 (I157895,I157878,I157762);
nand I_9129 (I157620,I157895,I371413);
DFFARX1 I_9130 (I157878,I2683,I157646,I157632,);
nand I_9131 (I157940,I157762,I371398);
nor I_9132 (I157957,I157762,I371398);
nand I_9133 (I157626,I157745,I157957);
not I_9134 (I157988,I371389);
nor I_9135 (I158005,I157988,I157940);
DFFARX1 I_9136 (I158005,I2683,I157646,I157614,);
nor I_9137 (I158036,I157988,I371401);
and I_9138 (I158053,I158036,I371395);
or I_9139 (I158070,I158053,I371392);
DFFARX1 I_9140 (I158070,I2683,I157646,I158096,);
nor I_9141 (I158104,I158096,I157720);
nor I_9142 (I157623,I157672,I158104);
not I_9143 (I158135,I158096);
nor I_9144 (I158152,I158135,I157830);
DFFARX1 I_9145 (I158152,I2683,I157646,I157629,);
nand I_9146 (I158183,I158135,I157762);
nor I_9147 (I157617,I157988,I158183);
not I_9148 (I158241,I2690);
DFFARX1 I_9149 (I87912,I2683,I158241,I158267,);
DFFARX1 I_9150 (I158267,I2683,I158241,I158284,);
not I_9151 (I158233,I158284);
DFFARX1 I_9152 (I87900,I2683,I158241,I158315,);
not I_9153 (I158323,I87903);
nor I_9154 (I158340,I158267,I158323);
not I_9155 (I158357,I87906);
not I_9156 (I158374,I87918);
nand I_9157 (I158391,I158374,I87906);
nor I_9158 (I158408,I158323,I158391);
nor I_9159 (I158425,I158315,I158408);
DFFARX1 I_9160 (I158374,I2683,I158241,I158230,);
nor I_9161 (I158456,I87918,I87909);
nand I_9162 (I158473,I158456,I87897);
nor I_9163 (I158490,I158473,I158357);
nand I_9164 (I158215,I158490,I87903);
DFFARX1 I_9165 (I158473,I2683,I158241,I158227,);
nand I_9166 (I158535,I158357,I87918);
nor I_9167 (I158552,I158357,I87918);
nand I_9168 (I158221,I158340,I158552);
not I_9169 (I158583,I87915);
nor I_9170 (I158600,I158583,I158535);
DFFARX1 I_9171 (I158600,I2683,I158241,I158209,);
nor I_9172 (I158631,I158583,I87921);
and I_9173 (I158648,I158631,I87924);
or I_9174 (I158665,I158648,I87897);
DFFARX1 I_9175 (I158665,I2683,I158241,I158691,);
nor I_9176 (I158699,I158691,I158315);
nor I_9177 (I158218,I158267,I158699);
not I_9178 (I158730,I158691);
nor I_9179 (I158747,I158730,I158425);
DFFARX1 I_9180 (I158747,I2683,I158241,I158224,);
nand I_9181 (I158778,I158730,I158357);
nor I_9182 (I158212,I158583,I158778);
not I_9183 (I158836,I2690);
DFFARX1 I_9184 (I212890,I2683,I158836,I158862,);
DFFARX1 I_9185 (I158862,I2683,I158836,I158879,);
not I_9186 (I158828,I158879);
DFFARX1 I_9187 (I212884,I2683,I158836,I158910,);
not I_9188 (I158918,I212881);
nor I_9189 (I158935,I158862,I158918);
not I_9190 (I158952,I212893);
not I_9191 (I158969,I212896);
nand I_9192 (I158986,I158969,I212893);
nor I_9193 (I159003,I158918,I158986);
nor I_9194 (I159020,I158910,I159003);
DFFARX1 I_9195 (I158969,I2683,I158836,I158825,);
nor I_9196 (I159051,I212896,I212905);
nand I_9197 (I159068,I159051,I212899);
nor I_9198 (I159085,I159068,I158952);
nand I_9199 (I158810,I159085,I212881);
DFFARX1 I_9200 (I159068,I2683,I158836,I158822,);
nand I_9201 (I159130,I158952,I212896);
nor I_9202 (I159147,I158952,I212896);
nand I_9203 (I158816,I158935,I159147);
not I_9204 (I159178,I212887);
nor I_9205 (I159195,I159178,I159130);
DFFARX1 I_9206 (I159195,I2683,I158836,I158804,);
nor I_9207 (I159226,I159178,I212902);
and I_9208 (I159243,I159226,I212881);
or I_9209 (I159260,I159243,I212884);
DFFARX1 I_9210 (I159260,I2683,I158836,I159286,);
nor I_9211 (I159294,I159286,I158910);
nor I_9212 (I158813,I158862,I159294);
not I_9213 (I159325,I159286);
nor I_9214 (I159342,I159325,I159020);
DFFARX1 I_9215 (I159342,I2683,I158836,I158819,);
nand I_9216 (I159373,I159325,I158952);
nor I_9217 (I158807,I159178,I159373);
not I_9218 (I159431,I2690);
DFFARX1 I_9219 (I313759,I2683,I159431,I159457,);
DFFARX1 I_9220 (I159457,I2683,I159431,I159474,);
not I_9221 (I159423,I159474);
DFFARX1 I_9222 (I313762,I2683,I159431,I159505,);
not I_9223 (I159513,I313765);
nor I_9224 (I159530,I159457,I159513);
not I_9225 (I159547,I313777);
not I_9226 (I159564,I313768);
nand I_9227 (I159581,I159564,I313777);
nor I_9228 (I159598,I159513,I159581);
nor I_9229 (I159615,I159505,I159598);
DFFARX1 I_9230 (I159564,I2683,I159431,I159420,);
nor I_9231 (I159646,I313768,I313774);
nand I_9232 (I159663,I159646,I313762);
nor I_9233 (I159680,I159663,I159547);
nand I_9234 (I159405,I159680,I313765);
DFFARX1 I_9235 (I159663,I2683,I159431,I159417,);
nand I_9236 (I159725,I159547,I313768);
nor I_9237 (I159742,I159547,I313768);
nand I_9238 (I159411,I159530,I159742);
not I_9239 (I159773,I313765);
nor I_9240 (I159790,I159773,I159725);
DFFARX1 I_9241 (I159790,I2683,I159431,I159399,);
nor I_9242 (I159821,I159773,I313771);
and I_9243 (I159838,I159821,I313759);
or I_9244 (I159855,I159838,I313780);
DFFARX1 I_9245 (I159855,I2683,I159431,I159881,);
nor I_9246 (I159889,I159881,I159505);
nor I_9247 (I159408,I159457,I159889);
not I_9248 (I159920,I159881);
nor I_9249 (I159937,I159920,I159615);
DFFARX1 I_9250 (I159937,I2683,I159431,I159414,);
nand I_9251 (I159968,I159920,I159547);
nor I_9252 (I159402,I159773,I159968);
not I_9253 (I160026,I2690);
DFFARX1 I_9254 (I39405,I2683,I160026,I160052,);
DFFARX1 I_9255 (I160052,I2683,I160026,I160069,);
not I_9256 (I160018,I160069);
DFFARX1 I_9257 (I39417,I2683,I160026,I160100,);
not I_9258 (I160108,I39408);
nor I_9259 (I160125,I160052,I160108);
not I_9260 (I160142,I39399);
not I_9261 (I160159,I39396);
nand I_9262 (I160176,I160159,I39399);
nor I_9263 (I160193,I160108,I160176);
nor I_9264 (I160210,I160100,I160193);
DFFARX1 I_9265 (I160159,I2683,I160026,I160015,);
nor I_9266 (I160241,I39396,I39396);
nand I_9267 (I160258,I160241,I39414);
nor I_9268 (I160275,I160258,I160142);
nand I_9269 (I160000,I160275,I39408);
DFFARX1 I_9270 (I160258,I2683,I160026,I160012,);
nand I_9271 (I160320,I160142,I39396);
nor I_9272 (I160337,I160142,I39396);
nand I_9273 (I160006,I160125,I160337);
not I_9274 (I160368,I39420);
nor I_9275 (I160385,I160368,I160320);
DFFARX1 I_9276 (I160385,I2683,I160026,I159994,);
nor I_9277 (I160416,I160368,I39399);
and I_9278 (I160433,I160416,I39402);
or I_9279 (I160450,I160433,I39411);
DFFARX1 I_9280 (I160450,I2683,I160026,I160476,);
nor I_9281 (I160484,I160476,I160100);
nor I_9282 (I160003,I160052,I160484);
not I_9283 (I160515,I160476);
nor I_9284 (I160532,I160515,I160210);
DFFARX1 I_9285 (I160532,I2683,I160026,I160009,);
nand I_9286 (I160563,I160515,I160142);
nor I_9287 (I159997,I160368,I160563);
not I_9288 (I160621,I2690);
DFFARX1 I_9289 (I382482,I2683,I160621,I160647,);
DFFARX1 I_9290 (I160647,I2683,I160621,I160664,);
not I_9291 (I160613,I160664);
DFFARX1 I_9292 (I382488,I2683,I160621,I160695,);
not I_9293 (I160703,I382476);
nor I_9294 (I160720,I160647,I160703);
not I_9295 (I160737,I382479);
not I_9296 (I160754,I382485);
nand I_9297 (I160771,I160754,I382479);
nor I_9298 (I160788,I160703,I160771);
nor I_9299 (I160805,I160695,I160788);
DFFARX1 I_9300 (I160754,I2683,I160621,I160610,);
nor I_9301 (I160836,I382485,I382476);
nand I_9302 (I160853,I160836,I382494);
nor I_9303 (I160870,I160853,I160737);
nand I_9304 (I160595,I160870,I382476);
DFFARX1 I_9305 (I160853,I2683,I160621,I160607,);
nand I_9306 (I160915,I160737,I382485);
nor I_9307 (I160932,I160737,I382485);
nand I_9308 (I160601,I160720,I160932);
not I_9309 (I160963,I382473);
nor I_9310 (I160980,I160963,I160915);
DFFARX1 I_9311 (I160980,I2683,I160621,I160589,);
nor I_9312 (I161011,I160963,I382497);
and I_9313 (I161028,I161011,I382473);
or I_9314 (I161045,I161028,I382491);
DFFARX1 I_9315 (I161045,I2683,I160621,I161071,);
nor I_9316 (I161079,I161071,I160695);
nor I_9317 (I160598,I160647,I161079);
not I_9318 (I161110,I161071);
nor I_9319 (I161127,I161110,I160805);
DFFARX1 I_9320 (I161127,I2683,I160621,I160604,);
nand I_9321 (I161158,I161110,I160737);
nor I_9322 (I160592,I160963,I161158);
not I_9323 (I161216,I2690);
DFFARX1 I_9324 (I16735,I2683,I161216,I161242,);
DFFARX1 I_9325 (I161242,I2683,I161216,I161259,);
not I_9326 (I161208,I161259);
DFFARX1 I_9327 (I16735,I2683,I161216,I161290,);
not I_9328 (I161298,I16750);
nor I_9329 (I161315,I161242,I161298);
not I_9330 (I161332,I16753);
not I_9331 (I161349,I16744);
nand I_9332 (I161366,I161349,I16753);
nor I_9333 (I161383,I161298,I161366);
nor I_9334 (I161400,I161290,I161383);
DFFARX1 I_9335 (I161349,I2683,I161216,I161205,);
nor I_9336 (I161431,I16744,I16756);
nand I_9337 (I161448,I161431,I16738);
nor I_9338 (I161465,I161448,I161332);
nand I_9339 (I161190,I161465,I16750);
DFFARX1 I_9340 (I161448,I2683,I161216,I161202,);
nand I_9341 (I161510,I161332,I16744);
nor I_9342 (I161527,I161332,I16744);
nand I_9343 (I161196,I161315,I161527);
not I_9344 (I161558,I16738);
nor I_9345 (I161575,I161558,I161510);
DFFARX1 I_9346 (I161575,I2683,I161216,I161184,);
nor I_9347 (I161606,I161558,I16747);
and I_9348 (I161623,I161606,I16741);
or I_9349 (I161640,I161623,I16759);
DFFARX1 I_9350 (I161640,I2683,I161216,I161666,);
nor I_9351 (I161674,I161666,I161290);
nor I_9352 (I161193,I161242,I161674);
not I_9353 (I161705,I161666);
nor I_9354 (I161722,I161705,I161400);
DFFARX1 I_9355 (I161722,I2683,I161216,I161199,);
nand I_9356 (I161753,I161705,I161332);
nor I_9357 (I161187,I161558,I161753);
not I_9358 (I161811,I2690);
DFFARX1 I_9359 (I77459,I2683,I161811,I161837,);
DFFARX1 I_9360 (I161837,I2683,I161811,I161854,);
not I_9361 (I161803,I161854);
DFFARX1 I_9362 (I77483,I2683,I161811,I161885,);
not I_9363 (I161893,I77477);
nor I_9364 (I161910,I161837,I161893);
not I_9365 (I161927,I77471);
not I_9366 (I161944,I77468);
nand I_9367 (I161961,I161944,I77471);
nor I_9368 (I161978,I161893,I161961);
nor I_9369 (I161995,I161885,I161978);
DFFARX1 I_9370 (I161944,I2683,I161811,I161800,);
nor I_9371 (I162026,I77468,I77462);
nand I_9372 (I162043,I162026,I77480);
nor I_9373 (I162060,I162043,I161927);
nand I_9374 (I161785,I162060,I77477);
DFFARX1 I_9375 (I162043,I2683,I161811,I161797,);
nand I_9376 (I162105,I161927,I77468);
nor I_9377 (I162122,I161927,I77468);
nand I_9378 (I161791,I161910,I162122);
not I_9379 (I162153,I77474);
nor I_9380 (I162170,I162153,I162105);
DFFARX1 I_9381 (I162170,I2683,I161811,I161779,);
nor I_9382 (I162201,I162153,I77459);
and I_9383 (I162218,I162201,I77465);
or I_9384 (I162235,I162218,I77462);
DFFARX1 I_9385 (I162235,I2683,I161811,I162261,);
nor I_9386 (I162269,I162261,I161885);
nor I_9387 (I161788,I161837,I162269);
not I_9388 (I162300,I162261);
nor I_9389 (I162317,I162300,I161995);
DFFARX1 I_9390 (I162317,I2683,I161811,I161794,);
nand I_9391 (I162348,I162300,I161927);
nor I_9392 (I161782,I162153,I162348);
not I_9393 (I162406,I2690);
DFFARX1 I_9394 (I249763,I2683,I162406,I162432,);
DFFARX1 I_9395 (I162432,I2683,I162406,I162449,);
not I_9396 (I162398,I162449);
DFFARX1 I_9397 (I249760,I2683,I162406,I162480,);
not I_9398 (I162488,I249760);
nor I_9399 (I162505,I162432,I162488);
not I_9400 (I162522,I249757);
not I_9401 (I162539,I249772);
nand I_9402 (I162556,I162539,I249757);
nor I_9403 (I162573,I162488,I162556);
nor I_9404 (I162590,I162480,I162573);
DFFARX1 I_9405 (I162539,I2683,I162406,I162395,);
nor I_9406 (I162621,I249772,I249766);
nand I_9407 (I162638,I162621,I249754);
nor I_9408 (I162655,I162638,I162522);
nand I_9409 (I162380,I162655,I249760);
DFFARX1 I_9410 (I162638,I2683,I162406,I162392,);
nand I_9411 (I162700,I162522,I249772);
nor I_9412 (I162717,I162522,I249772);
nand I_9413 (I162386,I162505,I162717);
not I_9414 (I162748,I249775);
nor I_9415 (I162765,I162748,I162700);
DFFARX1 I_9416 (I162765,I2683,I162406,I162374,);
nor I_9417 (I162796,I162748,I249754);
and I_9418 (I162813,I162796,I249769);
or I_9419 (I162830,I162813,I249757);
DFFARX1 I_9420 (I162830,I2683,I162406,I162856,);
nor I_9421 (I162864,I162856,I162480);
nor I_9422 (I162383,I162432,I162864);
not I_9423 (I162895,I162856);
nor I_9424 (I162912,I162895,I162590);
DFFARX1 I_9425 (I162912,I2683,I162406,I162389,);
nand I_9426 (I162943,I162895,I162522);
nor I_9427 (I162377,I162748,I162943);
not I_9428 (I163001,I2690);
DFFARX1 I_9429 (I2702,I2683,I163001,I163027,);
DFFARX1 I_9430 (I163027,I2683,I163001,I163044,);
not I_9431 (I162993,I163044);
DFFARX1 I_9432 (I2693,I2683,I163001,I163075,);
not I_9433 (I163083,I2696);
nor I_9434 (I163100,I163027,I163083);
not I_9435 (I163117,I2708);
not I_9436 (I163134,I2693);
nand I_9437 (I163151,I163134,I2708);
nor I_9438 (I163168,I163083,I163151);
nor I_9439 (I163185,I163075,I163168);
DFFARX1 I_9440 (I163134,I2683,I163001,I162990,);
nor I_9441 (I163216,I2693,I2699);
nand I_9442 (I163233,I163216,I2711);
nor I_9443 (I163250,I163233,I163117);
nand I_9444 (I162975,I163250,I2696);
DFFARX1 I_9445 (I163233,I2683,I163001,I162987,);
nand I_9446 (I163295,I163117,I2693);
nor I_9447 (I163312,I163117,I2693);
nand I_9448 (I162981,I163100,I163312);
not I_9449 (I163343,I2714);
nor I_9450 (I163360,I163343,I163295);
DFFARX1 I_9451 (I163360,I2683,I163001,I162969,);
nor I_9452 (I163391,I163343,I2696);
and I_9453 (I163408,I163391,I2705);
or I_9454 (I163425,I163408,I2699);
DFFARX1 I_9455 (I163425,I2683,I163001,I163451,);
nor I_9456 (I163459,I163451,I163075);
nor I_9457 (I162978,I163027,I163459);
not I_9458 (I163490,I163451);
nor I_9459 (I163507,I163490,I163185);
DFFARX1 I_9460 (I163507,I2683,I163001,I162984,);
nand I_9461 (I163538,I163490,I163117);
nor I_9462 (I162972,I163343,I163538);
not I_9463 (I163596,I2690);
DFFARX1 I_9464 (I78649,I2683,I163596,I163622,);
DFFARX1 I_9465 (I163622,I2683,I163596,I163639,);
not I_9466 (I163588,I163639);
DFFARX1 I_9467 (I78673,I2683,I163596,I163670,);
not I_9468 (I163678,I78667);
nor I_9469 (I163695,I163622,I163678);
not I_9470 (I163712,I78661);
not I_9471 (I163729,I78658);
nand I_9472 (I163746,I163729,I78661);
nor I_9473 (I163763,I163678,I163746);
nor I_9474 (I163780,I163670,I163763);
DFFARX1 I_9475 (I163729,I2683,I163596,I163585,);
nor I_9476 (I163811,I78658,I78652);
nand I_9477 (I163828,I163811,I78670);
nor I_9478 (I163845,I163828,I163712);
nand I_9479 (I163570,I163845,I78667);
DFFARX1 I_9480 (I163828,I2683,I163596,I163582,);
nand I_9481 (I163890,I163712,I78658);
nor I_9482 (I163907,I163712,I78658);
nand I_9483 (I163576,I163695,I163907);
not I_9484 (I163938,I78664);
nor I_9485 (I163955,I163938,I163890);
DFFARX1 I_9486 (I163955,I2683,I163596,I163564,);
nor I_9487 (I163986,I163938,I78649);
and I_9488 (I164003,I163986,I78655);
or I_9489 (I164020,I164003,I78652);
DFFARX1 I_9490 (I164020,I2683,I163596,I164046,);
nor I_9491 (I164054,I164046,I163670);
nor I_9492 (I163573,I163622,I164054);
not I_9493 (I164085,I164046);
nor I_9494 (I164102,I164085,I163780);
DFFARX1 I_9495 (I164102,I2683,I163596,I163579,);
nand I_9496 (I164133,I164085,I163712);
nor I_9497 (I163567,I163938,I164133);
not I_9498 (I164191,I2690);
DFFARX1 I_9499 (I314320,I2683,I164191,I164217,);
DFFARX1 I_9500 (I164217,I2683,I164191,I164234,);
not I_9501 (I164183,I164234);
DFFARX1 I_9502 (I314323,I2683,I164191,I164265,);
not I_9503 (I164273,I314326);
nor I_9504 (I164290,I164217,I164273);
not I_9505 (I164307,I314338);
not I_9506 (I164324,I314329);
nand I_9507 (I164341,I164324,I314338);
nor I_9508 (I164358,I164273,I164341);
nor I_9509 (I164375,I164265,I164358);
DFFARX1 I_9510 (I164324,I2683,I164191,I164180,);
nor I_9511 (I164406,I314329,I314335);
nand I_9512 (I164423,I164406,I314323);
nor I_9513 (I164440,I164423,I164307);
nand I_9514 (I164165,I164440,I314326);
DFFARX1 I_9515 (I164423,I2683,I164191,I164177,);
nand I_9516 (I164485,I164307,I314329);
nor I_9517 (I164502,I164307,I314329);
nand I_9518 (I164171,I164290,I164502);
not I_9519 (I164533,I314326);
nor I_9520 (I164550,I164533,I164485);
DFFARX1 I_9521 (I164550,I2683,I164191,I164159,);
nor I_9522 (I164581,I164533,I314332);
and I_9523 (I164598,I164581,I314320);
or I_9524 (I164615,I164598,I314341);
DFFARX1 I_9525 (I164615,I2683,I164191,I164641,);
nor I_9526 (I164649,I164641,I164265);
nor I_9527 (I164168,I164217,I164649);
not I_9528 (I164680,I164641);
nor I_9529 (I164697,I164680,I164375);
DFFARX1 I_9530 (I164697,I2683,I164191,I164174,);
nand I_9531 (I164728,I164680,I164307);
nor I_9532 (I164162,I164533,I164728);
not I_9533 (I164786,I2690);
DFFARX1 I_9534 (I93182,I2683,I164786,I164812,);
DFFARX1 I_9535 (I164812,I2683,I164786,I164829,);
not I_9536 (I164778,I164829);
DFFARX1 I_9537 (I93170,I2683,I164786,I164860,);
not I_9538 (I164868,I93173);
nor I_9539 (I164885,I164812,I164868);
not I_9540 (I164902,I93176);
not I_9541 (I164919,I93188);
nand I_9542 (I164936,I164919,I93176);
nor I_9543 (I164953,I164868,I164936);
nor I_9544 (I164970,I164860,I164953);
DFFARX1 I_9545 (I164919,I2683,I164786,I164775,);
nor I_9546 (I165001,I93188,I93179);
nand I_9547 (I165018,I165001,I93167);
nor I_9548 (I165035,I165018,I164902);
nand I_9549 (I164760,I165035,I93173);
DFFARX1 I_9550 (I165018,I2683,I164786,I164772,);
nand I_9551 (I165080,I164902,I93188);
nor I_9552 (I165097,I164902,I93188);
nand I_9553 (I164766,I164885,I165097);
not I_9554 (I165128,I93185);
nor I_9555 (I165145,I165128,I165080);
DFFARX1 I_9556 (I165145,I2683,I164786,I164754,);
nor I_9557 (I165176,I165128,I93191);
and I_9558 (I165193,I165176,I93194);
or I_9559 (I165210,I165193,I93167);
DFFARX1 I_9560 (I165210,I2683,I164786,I165236,);
nor I_9561 (I165244,I165236,I164860);
nor I_9562 (I164763,I164812,I165244);
not I_9563 (I165275,I165236);
nor I_9564 (I165292,I165275,I164970);
DFFARX1 I_9565 (I165292,I2683,I164786,I164769,);
nand I_9566 (I165323,I165275,I164902);
nor I_9567 (I164757,I165128,I165323);
not I_9568 (I165381,I2690);
DFFARX1 I_9569 (I93709,I2683,I165381,I165407,);
DFFARX1 I_9570 (I165407,I2683,I165381,I165424,);
not I_9571 (I165373,I165424);
DFFARX1 I_9572 (I93697,I2683,I165381,I165455,);
not I_9573 (I165463,I93700);
nor I_9574 (I165480,I165407,I165463);
not I_9575 (I165497,I93703);
not I_9576 (I165514,I93715);
nand I_9577 (I165531,I165514,I93703);
nor I_9578 (I165548,I165463,I165531);
nor I_9579 (I165565,I165455,I165548);
DFFARX1 I_9580 (I165514,I2683,I165381,I165370,);
nor I_9581 (I165596,I93715,I93706);
nand I_9582 (I165613,I165596,I93694);
nor I_9583 (I165630,I165613,I165497);
nand I_9584 (I165355,I165630,I93700);
DFFARX1 I_9585 (I165613,I2683,I165381,I165367,);
nand I_9586 (I165675,I165497,I93715);
nor I_9587 (I165692,I165497,I93715);
nand I_9588 (I165361,I165480,I165692);
not I_9589 (I165723,I93712);
nor I_9590 (I165740,I165723,I165675);
DFFARX1 I_9591 (I165740,I2683,I165381,I165349,);
nor I_9592 (I165771,I165723,I93718);
and I_9593 (I165788,I165771,I93721);
or I_9594 (I165805,I165788,I93694);
DFFARX1 I_9595 (I165805,I2683,I165381,I165831,);
nor I_9596 (I165839,I165831,I165455);
nor I_9597 (I165358,I165407,I165839);
not I_9598 (I165870,I165831);
nor I_9599 (I165887,I165870,I165565);
DFFARX1 I_9600 (I165887,I2683,I165381,I165364,);
nand I_9601 (I165918,I165870,I165497);
nor I_9602 (I165352,I165723,I165918);
not I_9603 (I165976,I2690);
DFFARX1 I_9604 (I333123,I2683,I165976,I166002,);
DFFARX1 I_9605 (I166002,I2683,I165976,I166019,);
not I_9606 (I165968,I166019);
DFFARX1 I_9607 (I333105,I2683,I165976,I166050,);
not I_9608 (I166058,I333111);
nor I_9609 (I166075,I166002,I166058);
not I_9610 (I166092,I333126);
not I_9611 (I166109,I333117);
nand I_9612 (I166126,I166109,I333126);
nor I_9613 (I166143,I166058,I166126);
nor I_9614 (I166160,I166050,I166143);
DFFARX1 I_9615 (I166109,I2683,I165976,I165965,);
nor I_9616 (I166191,I333117,I333129);
nand I_9617 (I166208,I166191,I333108);
nor I_9618 (I166225,I166208,I166092);
nand I_9619 (I165950,I166225,I333111);
DFFARX1 I_9620 (I166208,I2683,I165976,I165962,);
nand I_9621 (I166270,I166092,I333117);
nor I_9622 (I166287,I166092,I333117);
nand I_9623 (I165956,I166075,I166287);
not I_9624 (I166318,I333114);
nor I_9625 (I166335,I166318,I166270);
DFFARX1 I_9626 (I166335,I2683,I165976,I165944,);
nor I_9627 (I166366,I166318,I333120);
and I_9628 (I166383,I166366,I333105);
or I_9629 (I166400,I166383,I333108);
DFFARX1 I_9630 (I166400,I2683,I165976,I166426,);
nor I_9631 (I166434,I166426,I166050);
nor I_9632 (I165953,I166002,I166434);
not I_9633 (I166465,I166426);
nor I_9634 (I166482,I166465,I166160);
DFFARX1 I_9635 (I166482,I2683,I165976,I165959,);
nand I_9636 (I166513,I166465,I166092);
nor I_9637 (I165947,I166318,I166513);
not I_9638 (I166571,I2690);
DFFARX1 I_9639 (I274963,I2683,I166571,I166597,);
DFFARX1 I_9640 (I166597,I2683,I166571,I166614,);
not I_9641 (I166563,I166614);
DFFARX1 I_9642 (I274951,I2683,I166571,I166645,);
not I_9643 (I166653,I274948);
nor I_9644 (I166670,I166597,I166653);
not I_9645 (I166687,I274960);
not I_9646 (I166704,I274957);
nand I_9647 (I166721,I166704,I274960);
nor I_9648 (I166738,I166653,I166721);
nor I_9649 (I166755,I166645,I166738);
DFFARX1 I_9650 (I166704,I2683,I166571,I166560,);
nor I_9651 (I166786,I274957,I274966);
nand I_9652 (I166803,I166786,I274969);
nor I_9653 (I166820,I166803,I166687);
nand I_9654 (I166545,I166820,I274948);
DFFARX1 I_9655 (I166803,I2683,I166571,I166557,);
nand I_9656 (I166865,I166687,I274957);
nor I_9657 (I166882,I166687,I274957);
nand I_9658 (I166551,I166670,I166882);
not I_9659 (I166913,I274972);
nor I_9660 (I166930,I166913,I166865);
DFFARX1 I_9661 (I166930,I2683,I166571,I166539,);
nor I_9662 (I166961,I166913,I274975);
and I_9663 (I166978,I166961,I274954);
or I_9664 (I166995,I166978,I274948);
DFFARX1 I_9665 (I166995,I2683,I166571,I167021,);
nor I_9666 (I167029,I167021,I166645);
nor I_9667 (I166548,I166597,I167029);
not I_9668 (I167060,I167021);
nor I_9669 (I167077,I167060,I166755);
DFFARX1 I_9670 (I167077,I2683,I166571,I166554,);
nand I_9671 (I167108,I167060,I166687);
nor I_9672 (I166542,I166913,I167108);
not I_9673 (I167166,I2690);
DFFARX1 I_9674 (I12519,I2683,I167166,I167192,);
DFFARX1 I_9675 (I167192,I2683,I167166,I167209,);
not I_9676 (I167158,I167209);
DFFARX1 I_9677 (I12519,I2683,I167166,I167240,);
not I_9678 (I167248,I12534);
nor I_9679 (I167265,I167192,I167248);
not I_9680 (I167282,I12537);
not I_9681 (I167299,I12528);
nand I_9682 (I167316,I167299,I12537);
nor I_9683 (I167333,I167248,I167316);
nor I_9684 (I167350,I167240,I167333);
DFFARX1 I_9685 (I167299,I2683,I167166,I167155,);
nor I_9686 (I167381,I12528,I12540);
nand I_9687 (I167398,I167381,I12522);
nor I_9688 (I167415,I167398,I167282);
nand I_9689 (I167140,I167415,I12534);
DFFARX1 I_9690 (I167398,I2683,I167166,I167152,);
nand I_9691 (I167460,I167282,I12528);
nor I_9692 (I167477,I167282,I12528);
nand I_9693 (I167146,I167265,I167477);
not I_9694 (I167508,I12522);
nor I_9695 (I167525,I167508,I167460);
DFFARX1 I_9696 (I167525,I2683,I167166,I167134,);
nor I_9697 (I167556,I167508,I12531);
and I_9698 (I167573,I167556,I12525);
or I_9699 (I167590,I167573,I12543);
DFFARX1 I_9700 (I167590,I2683,I167166,I167616,);
nor I_9701 (I167624,I167616,I167240);
nor I_9702 (I167143,I167192,I167624);
not I_9703 (I167655,I167616);
nor I_9704 (I167672,I167655,I167350);
DFFARX1 I_9705 (I167672,I2683,I167166,I167149,);
nand I_9706 (I167703,I167655,I167282);
nor I_9707 (I167137,I167508,I167703);
not I_9708 (I167761,I2690);
DFFARX1 I_9709 (I267681,I2683,I167761,I167787,);
DFFARX1 I_9710 (I167787,I2683,I167761,I167804,);
not I_9711 (I167753,I167804);
DFFARX1 I_9712 (I267678,I2683,I167761,I167835,);
not I_9713 (I167843,I267678);
nor I_9714 (I167860,I167787,I167843);
not I_9715 (I167877,I267675);
not I_9716 (I167894,I267690);
nand I_9717 (I167911,I167894,I267675);
nor I_9718 (I167928,I167843,I167911);
nor I_9719 (I167945,I167835,I167928);
DFFARX1 I_9720 (I167894,I2683,I167761,I167750,);
nor I_9721 (I167976,I267690,I267684);
nand I_9722 (I167993,I167976,I267672);
nor I_9723 (I168010,I167993,I167877);
nand I_9724 (I167735,I168010,I267678);
DFFARX1 I_9725 (I167993,I2683,I167761,I167747,);
nand I_9726 (I168055,I167877,I267690);
nor I_9727 (I168072,I167877,I267690);
nand I_9728 (I167741,I167860,I168072);
not I_9729 (I168103,I267693);
nor I_9730 (I168120,I168103,I168055);
DFFARX1 I_9731 (I168120,I2683,I167761,I167729,);
nor I_9732 (I168151,I168103,I267672);
and I_9733 (I168168,I168151,I267687);
or I_9734 (I168185,I168168,I267675);
DFFARX1 I_9735 (I168185,I2683,I167761,I168211,);
nor I_9736 (I168219,I168211,I167835);
nor I_9737 (I167738,I167787,I168219);
not I_9738 (I168250,I168211);
nor I_9739 (I168267,I168250,I167945);
DFFARX1 I_9740 (I168267,I2683,I167761,I167744,);
nand I_9741 (I168298,I168250,I167877);
nor I_9742 (I167732,I168103,I168298);
not I_9743 (I168356,I2690);
DFFARX1 I_9744 (I88439,I2683,I168356,I168382,);
DFFARX1 I_9745 (I168382,I2683,I168356,I168399,);
not I_9746 (I168348,I168399);
DFFARX1 I_9747 (I88427,I2683,I168356,I168430,);
not I_9748 (I168438,I88430);
nor I_9749 (I168455,I168382,I168438);
not I_9750 (I168472,I88433);
not I_9751 (I168489,I88445);
nand I_9752 (I168506,I168489,I88433);
nor I_9753 (I168523,I168438,I168506);
nor I_9754 (I168540,I168430,I168523);
DFFARX1 I_9755 (I168489,I2683,I168356,I168345,);
nor I_9756 (I168571,I88445,I88436);
nand I_9757 (I168588,I168571,I88424);
nor I_9758 (I168605,I168588,I168472);
nand I_9759 (I168330,I168605,I88430);
DFFARX1 I_9760 (I168588,I2683,I168356,I168342,);
nand I_9761 (I168650,I168472,I88445);
nor I_9762 (I168667,I168472,I88445);
nand I_9763 (I168336,I168455,I168667);
not I_9764 (I168698,I88442);
nor I_9765 (I168715,I168698,I168650);
DFFARX1 I_9766 (I168715,I2683,I168356,I168324,);
nor I_9767 (I168746,I168698,I88448);
and I_9768 (I168763,I168746,I88451);
or I_9769 (I168780,I168763,I88424);
DFFARX1 I_9770 (I168780,I2683,I168356,I168806,);
nor I_9771 (I168814,I168806,I168430);
nor I_9772 (I168333,I168382,I168814);
not I_9773 (I168845,I168806);
nor I_9774 (I168862,I168845,I168540);
DFFARX1 I_9775 (I168862,I2683,I168356,I168339,);
nand I_9776 (I168893,I168845,I168472);
nor I_9777 (I168327,I168698,I168893);
not I_9778 (I168951,I2690);
DFFARX1 I_9779 (I195550,I2683,I168951,I168977,);
DFFARX1 I_9780 (I168977,I2683,I168951,I168994,);
not I_9781 (I168943,I168994);
DFFARX1 I_9782 (I195544,I2683,I168951,I169025,);
not I_9783 (I169033,I195541);
nor I_9784 (I169050,I168977,I169033);
not I_9785 (I169067,I195553);
not I_9786 (I169084,I195556);
nand I_9787 (I169101,I169084,I195553);
nor I_9788 (I169118,I169033,I169101);
nor I_9789 (I169135,I169025,I169118);
DFFARX1 I_9790 (I169084,I2683,I168951,I168940,);
nor I_9791 (I169166,I195556,I195565);
nand I_9792 (I169183,I169166,I195559);
nor I_9793 (I169200,I169183,I169067);
nand I_9794 (I168925,I169200,I195541);
DFFARX1 I_9795 (I169183,I2683,I168951,I168937,);
nand I_9796 (I169245,I169067,I195556);
nor I_9797 (I169262,I169067,I195556);
nand I_9798 (I168931,I169050,I169262);
not I_9799 (I169293,I195547);
nor I_9800 (I169310,I169293,I169245);
DFFARX1 I_9801 (I169310,I2683,I168951,I168919,);
nor I_9802 (I169341,I169293,I195562);
and I_9803 (I169358,I169341,I195541);
or I_9804 (I169375,I169358,I195544);
DFFARX1 I_9805 (I169375,I2683,I168951,I169401,);
nor I_9806 (I169409,I169401,I169025);
nor I_9807 (I168928,I168977,I169409);
not I_9808 (I169440,I169401);
nor I_9809 (I169457,I169440,I169135);
DFFARX1 I_9810 (I169457,I2683,I168951,I168934,);
nand I_9811 (I169488,I169440,I169067);
nor I_9812 (I168922,I169293,I169488);
not I_9813 (I169546,I2690);
DFFARX1 I_9814 (I88966,I2683,I169546,I169572,);
DFFARX1 I_9815 (I169572,I2683,I169546,I169589,);
not I_9816 (I169538,I169589);
DFFARX1 I_9817 (I88954,I2683,I169546,I169620,);
not I_9818 (I169628,I88957);
nor I_9819 (I169645,I169572,I169628);
not I_9820 (I169662,I88960);
not I_9821 (I169679,I88972);
nand I_9822 (I169696,I169679,I88960);
nor I_9823 (I169713,I169628,I169696);
nor I_9824 (I169730,I169620,I169713);
DFFARX1 I_9825 (I169679,I2683,I169546,I169535,);
nor I_9826 (I169761,I88972,I88963);
nand I_9827 (I169778,I169761,I88951);
nor I_9828 (I169795,I169778,I169662);
nand I_9829 (I169520,I169795,I88957);
DFFARX1 I_9830 (I169778,I2683,I169546,I169532,);
nand I_9831 (I169840,I169662,I88972);
nor I_9832 (I169857,I169662,I88972);
nand I_9833 (I169526,I169645,I169857);
not I_9834 (I169888,I88969);
nor I_9835 (I169905,I169888,I169840);
DFFARX1 I_9836 (I169905,I2683,I169546,I169514,);
nor I_9837 (I169936,I169888,I88975);
and I_9838 (I169953,I169936,I88978);
or I_9839 (I169970,I169953,I88951);
DFFARX1 I_9840 (I169970,I2683,I169546,I169996,);
nor I_9841 (I170004,I169996,I169620);
nor I_9842 (I169523,I169572,I170004);
not I_9843 (I170035,I169996);
nor I_9844 (I170052,I170035,I169730);
DFFARX1 I_9845 (I170052,I2683,I169546,I169529,);
nand I_9846 (I170083,I170035,I169662);
nor I_9847 (I169517,I169888,I170083);
not I_9848 (I170141,I2690);
DFFARX1 I_9849 (I265043,I2683,I170141,I170167,);
not I_9850 (I170175,I170167);
DFFARX1 I_9851 (I265043,I2683,I170141,I170201,);
not I_9852 (I170209,I265040);
nand I_9853 (I170226,I170209,I265055);
not I_9854 (I170243,I170226);
nor I_9855 (I170260,I170243,I265049);
nor I_9856 (I170277,I170175,I170260);
DFFARX1 I_9857 (I170277,I2683,I170141,I170127,);
not I_9858 (I170308,I265049);
nand I_9859 (I170325,I170308,I170243);
and I_9860 (I170342,I170308,I265046);
nand I_9861 (I170359,I170342,I265037);
nor I_9862 (I170124,I170359,I170308);
and I_9863 (I170115,I170201,I170359);
not I_9864 (I170404,I170359);
nand I_9865 (I170118,I170201,I170404);
nor I_9866 (I170112,I170167,I170359);
not I_9867 (I170449,I265058);
nor I_9868 (I170466,I170449,I265046);
nand I_9869 (I170483,I170466,I170308);
nor I_9870 (I170121,I170226,I170483);
nor I_9871 (I170514,I170449,I265037);
and I_9872 (I170531,I170514,I265040);
or I_9873 (I170548,I170531,I265052);
DFFARX1 I_9874 (I170548,I2683,I170141,I170574,);
nor I_9875 (I170582,I170574,I170325);
DFFARX1 I_9876 (I170582,I2683,I170141,I170109,);
DFFARX1 I_9877 (I170574,I2683,I170141,I170133,);
not I_9878 (I170627,I170574);
nor I_9879 (I170644,I170627,I170201);
nor I_9880 (I170661,I170466,I170644);
DFFARX1 I_9881 (I170661,I2683,I170141,I170130,);
not I_9882 (I170719,I2690);
DFFARX1 I_9883 (I337729,I2683,I170719,I170745,);
not I_9884 (I170753,I170745);
DFFARX1 I_9885 (I337735,I2683,I170719,I170779,);
not I_9886 (I170787,I337729);
nand I_9887 (I170804,I170787,I337732);
not I_9888 (I170821,I170804);
nor I_9889 (I170838,I170821,I337750);
nor I_9890 (I170855,I170753,I170838);
DFFARX1 I_9891 (I170855,I2683,I170719,I170705,);
not I_9892 (I170886,I337750);
nand I_9893 (I170903,I170886,I170821);
and I_9894 (I170920,I170886,I337753);
nand I_9895 (I170937,I170920,I337732);
nor I_9896 (I170702,I170937,I170886);
and I_9897 (I170693,I170779,I170937);
not I_9898 (I170982,I170937);
nand I_9899 (I170696,I170779,I170982);
nor I_9900 (I170690,I170745,I170937);
not I_9901 (I171027,I337738);
nor I_9902 (I171044,I171027,I337753);
nand I_9903 (I171061,I171044,I170886);
nor I_9904 (I170699,I170804,I171061);
nor I_9905 (I171092,I171027,I337744);
and I_9906 (I171109,I171092,I337741);
or I_9907 (I171126,I171109,I337747);
DFFARX1 I_9908 (I171126,I2683,I170719,I171152,);
nor I_9909 (I171160,I171152,I170903);
DFFARX1 I_9910 (I171160,I2683,I170719,I170687,);
DFFARX1 I_9911 (I171152,I2683,I170719,I170711,);
not I_9912 (I171205,I171152);
nor I_9913 (I171222,I171205,I170779);
nor I_9914 (I171239,I171044,I171222);
DFFARX1 I_9915 (I171239,I2683,I170719,I170708,);
not I_9916 (I171297,I2690);
DFFARX1 I_9917 (I149211,I2683,I171297,I171323,);
not I_9918 (I171331,I171323);
DFFARX1 I_9919 (I149223,I2683,I171297,I171357,);
not I_9920 (I171365,I149199);
nand I_9921 (I171382,I171365,I149226);
not I_9922 (I171399,I171382);
nor I_9923 (I171416,I171399,I149214);
nor I_9924 (I171433,I171331,I171416);
DFFARX1 I_9925 (I171433,I2683,I171297,I171283,);
not I_9926 (I171464,I149214);
nand I_9927 (I171481,I171464,I171399);
and I_9928 (I171498,I171464,I149199);
nand I_9929 (I171515,I171498,I149202);
nor I_9930 (I171280,I171515,I171464);
and I_9931 (I171271,I171357,I171515);
not I_9932 (I171560,I171515);
nand I_9933 (I171274,I171357,I171560);
nor I_9934 (I171268,I171323,I171515);
not I_9935 (I171605,I149208);
nor I_9936 (I171622,I171605,I149199);
nand I_9937 (I171639,I171622,I171464);
nor I_9938 (I171277,I171382,I171639);
nor I_9939 (I171670,I171605,I149217);
and I_9940 (I171687,I171670,I149205);
or I_9941 (I171704,I171687,I149220);
DFFARX1 I_9942 (I171704,I2683,I171297,I171730,);
nor I_9943 (I171738,I171730,I171481);
DFFARX1 I_9944 (I171738,I2683,I171297,I171265,);
DFFARX1 I_9945 (I171730,I2683,I171297,I171289,);
not I_9946 (I171783,I171730);
nor I_9947 (I171800,I171783,I171357);
nor I_9948 (I171817,I171622,I171800);
DFFARX1 I_9949 (I171817,I2683,I171297,I171286,);
not I_9950 (I171875,I2690);
DFFARX1 I_9951 (I16211,I2683,I171875,I171901,);
not I_9952 (I171909,I171901);
DFFARX1 I_9953 (I16214,I2683,I171875,I171935,);
not I_9954 (I171943,I16208);
nand I_9955 (I171960,I171943,I16232);
not I_9956 (I171977,I171960);
nor I_9957 (I171994,I171977,I16211);
nor I_9958 (I172011,I171909,I171994);
DFFARX1 I_9959 (I172011,I2683,I171875,I171861,);
not I_9960 (I172042,I16211);
nand I_9961 (I172059,I172042,I171977);
and I_9962 (I172076,I172042,I16226);
nand I_9963 (I172093,I172076,I16220);
nor I_9964 (I171858,I172093,I172042);
and I_9965 (I171849,I171935,I172093);
not I_9966 (I172138,I172093);
nand I_9967 (I171852,I171935,I172138);
nor I_9968 (I171846,I171901,I172093);
not I_9969 (I172183,I16229);
nor I_9970 (I172200,I172183,I16226);
nand I_9971 (I172217,I172200,I172042);
nor I_9972 (I171855,I171960,I172217);
nor I_9973 (I172248,I172183,I16208);
and I_9974 (I172265,I172248,I16217);
or I_9975 (I172282,I172265,I16223);
DFFARX1 I_9976 (I172282,I2683,I171875,I172308,);
nor I_9977 (I172316,I172308,I172059);
DFFARX1 I_9978 (I172316,I2683,I171875,I171843,);
DFFARX1 I_9979 (I172308,I2683,I171875,I171867,);
not I_9980 (I172361,I172308);
nor I_9981 (I172378,I172361,I171935);
nor I_9982 (I172395,I172200,I172378);
DFFARX1 I_9983 (I172395,I2683,I171875,I171864,);
not I_9984 (I172453,I2690);
DFFARX1 I_9985 (I213459,I2683,I172453,I172479,);
not I_9986 (I172487,I172479);
DFFARX1 I_9987 (I213471,I2683,I172453,I172513,);
not I_9988 (I172521,I213462);
nand I_9989 (I172538,I172521,I213465);
not I_9990 (I172555,I172538);
nor I_9991 (I172572,I172555,I213468);
nor I_9992 (I172589,I172487,I172572);
DFFARX1 I_9993 (I172589,I2683,I172453,I172439,);
not I_9994 (I172620,I213468);
nand I_9995 (I172637,I172620,I172555);
and I_9996 (I172654,I172620,I213462);
nand I_9997 (I172671,I172654,I213474);
nor I_9998 (I172436,I172671,I172620);
and I_9999 (I172427,I172513,I172671);
not I_10000 (I172716,I172671);
nand I_10001 (I172430,I172513,I172716);
nor I_10002 (I172424,I172479,I172671);
not I_10003 (I172761,I213480);
nor I_10004 (I172778,I172761,I213462);
nand I_10005 (I172795,I172778,I172620);
nor I_10006 (I172433,I172538,I172795);
nor I_10007 (I172826,I172761,I213459);
and I_10008 (I172843,I172826,I213477);
or I_10009 (I172860,I172843,I213483);
DFFARX1 I_10010 (I172860,I2683,I172453,I172886,);
nor I_10011 (I172894,I172886,I172637);
DFFARX1 I_10012 (I172894,I2683,I172453,I172421,);
DFFARX1 I_10013 (I172886,I2683,I172453,I172445,);
not I_10014 (I172939,I172886);
nor I_10015 (I172956,I172939,I172513);
nor I_10016 (I172973,I172778,I172956);
DFFARX1 I_10017 (I172973,I2683,I172453,I172442,);
not I_10018 (I173031,I2690);
DFFARX1 I_10019 (I41528,I2683,I173031,I173057,);
not I_10020 (I173065,I173057);
DFFARX1 I_10021 (I41507,I2683,I173031,I173091,);
not I_10022 (I173099,I41504);
nand I_10023 (I173116,I173099,I41519);
not I_10024 (I173133,I173116);
nor I_10025 (I173150,I173133,I41507);
nor I_10026 (I173167,I173065,I173150);
DFFARX1 I_10027 (I173167,I2683,I173031,I173017,);
not I_10028 (I173198,I41507);
nand I_10029 (I173215,I173198,I173133);
and I_10030 (I173232,I173198,I41510);
nand I_10031 (I173249,I173232,I41525);
nor I_10032 (I173014,I173249,I173198);
and I_10033 (I173005,I173091,I173249);
not I_10034 (I173294,I173249);
nand I_10035 (I173008,I173091,I173294);
nor I_10036 (I173002,I173057,I173249);
not I_10037 (I173339,I41516);
nor I_10038 (I173356,I173339,I41510);
nand I_10039 (I173373,I173356,I173198);
nor I_10040 (I173011,I173116,I173373);
nor I_10041 (I173404,I173339,I41504);
and I_10042 (I173421,I173404,I41513);
or I_10043 (I173438,I173421,I41522);
DFFARX1 I_10044 (I173438,I2683,I173031,I173464,);
nor I_10045 (I173472,I173464,I173215);
DFFARX1 I_10046 (I173472,I2683,I173031,I172999,);
DFFARX1 I_10047 (I173464,I2683,I173031,I173023,);
not I_10048 (I173517,I173464);
nor I_10049 (I173534,I173517,I173091);
nor I_10050 (I173551,I173356,I173534);
DFFARX1 I_10051 (I173551,I2683,I173031,I173020,);
not I_10052 (I173609,I2690);
DFFARX1 I_10053 (I141051,I2683,I173609,I173635,);
not I_10054 (I173643,I173635);
DFFARX1 I_10055 (I141063,I2683,I173609,I173669,);
not I_10056 (I173677,I141039);
nand I_10057 (I173694,I173677,I141066);
not I_10058 (I173711,I173694);
nor I_10059 (I173728,I173711,I141054);
nor I_10060 (I173745,I173643,I173728);
DFFARX1 I_10061 (I173745,I2683,I173609,I173595,);
not I_10062 (I173776,I141054);
nand I_10063 (I173793,I173776,I173711);
and I_10064 (I173810,I173776,I141039);
nand I_10065 (I173827,I173810,I141042);
nor I_10066 (I173592,I173827,I173776);
and I_10067 (I173583,I173669,I173827);
not I_10068 (I173872,I173827);
nand I_10069 (I173586,I173669,I173872);
nor I_10070 (I173580,I173635,I173827);
not I_10071 (I173917,I141048);
nor I_10072 (I173934,I173917,I141039);
nand I_10073 (I173951,I173934,I173776);
nor I_10074 (I173589,I173694,I173951);
nor I_10075 (I173982,I173917,I141057);
and I_10076 (I173999,I173982,I141045);
or I_10077 (I174016,I173999,I141060);
DFFARX1 I_10078 (I174016,I2683,I173609,I174042,);
nor I_10079 (I174050,I174042,I173793);
DFFARX1 I_10080 (I174050,I2683,I173609,I173577,);
DFFARX1 I_10081 (I174042,I2683,I173609,I173601,);
not I_10082 (I174095,I174042);
nor I_10083 (I174112,I174095,I173669);
nor I_10084 (I174129,I173934,I174112);
DFFARX1 I_10085 (I174129,I2683,I173609,I173598,);
not I_10086 (I174187,I2690);
DFFARX1 I_10087 (I159402,I2683,I174187,I174213,);
not I_10088 (I174221,I174213);
DFFARX1 I_10089 (I159414,I2683,I174187,I174247,);
not I_10090 (I174255,I159420);
nand I_10091 (I174272,I174255,I159411);
not I_10092 (I174289,I174272);
nor I_10093 (I174306,I174289,I159417);
nor I_10094 (I174323,I174221,I174306);
DFFARX1 I_10095 (I174323,I2683,I174187,I174173,);
not I_10096 (I174354,I159417);
nand I_10097 (I174371,I174354,I174289);
and I_10098 (I174388,I174354,I159408);
nand I_10099 (I174405,I174388,I159399);
nor I_10100 (I174170,I174405,I174354);
and I_10101 (I174161,I174247,I174405);
not I_10102 (I174450,I174405);
nand I_10103 (I174164,I174247,I174450);
nor I_10104 (I174158,I174213,I174405);
not I_10105 (I174495,I159405);
nor I_10106 (I174512,I174495,I159408);
nand I_10107 (I174529,I174512,I174354);
nor I_10108 (I174167,I174272,I174529);
nor I_10109 (I174560,I174495,I159402);
and I_10110 (I174577,I174560,I159399);
or I_10111 (I174594,I174577,I159423);
DFFARX1 I_10112 (I174594,I2683,I174187,I174620,);
nor I_10113 (I174628,I174620,I174371);
DFFARX1 I_10114 (I174628,I2683,I174187,I174155,);
DFFARX1 I_10115 (I174620,I2683,I174187,I174179,);
not I_10116 (I174673,I174620);
nor I_10117 (I174690,I174673,I174247);
nor I_10118 (I174707,I174512,I174690);
DFFARX1 I_10119 (I174707,I2683,I174187,I174176,);
not I_10120 (I174765,I2690);
DFFARX1 I_10121 (I412274,I2683,I174765,I174791,);
not I_10122 (I174799,I174791);
DFFARX1 I_10123 (I412274,I2683,I174765,I174825,);
not I_10124 (I174833,I412298);
nand I_10125 (I174850,I174833,I412280);
not I_10126 (I174867,I174850);
nor I_10127 (I174884,I174867,I412295);
nor I_10128 (I174901,I174799,I174884);
DFFARX1 I_10129 (I174901,I2683,I174765,I174751,);
not I_10130 (I174932,I412295);
nand I_10131 (I174949,I174932,I174867);
and I_10132 (I174966,I174932,I412277);
nand I_10133 (I174983,I174966,I412286);
nor I_10134 (I174748,I174983,I174932);
and I_10135 (I174739,I174825,I174983);
not I_10136 (I175028,I174983);
nand I_10137 (I174742,I174825,I175028);
nor I_10138 (I174736,I174791,I174983);
not I_10139 (I175073,I412283);
nor I_10140 (I175090,I175073,I412277);
nand I_10141 (I175107,I175090,I174932);
nor I_10142 (I174745,I174850,I175107);
nor I_10143 (I175138,I175073,I412292);
and I_10144 (I175155,I175138,I412301);
or I_10145 (I175172,I175155,I412289);
DFFARX1 I_10146 (I175172,I2683,I174765,I175198,);
nor I_10147 (I175206,I175198,I174949);
DFFARX1 I_10148 (I175206,I2683,I174765,I174733,);
DFFARX1 I_10149 (I175198,I2683,I174765,I174757,);
not I_10150 (I175251,I175198);
nor I_10151 (I175268,I175251,I174825);
nor I_10152 (I175285,I175090,I175268);
DFFARX1 I_10153 (I175285,I2683,I174765,I174754,);
not I_10154 (I175343,I2690);
DFFARX1 I_10155 (I357381,I2683,I175343,I175369,);
not I_10156 (I175377,I175369);
DFFARX1 I_10157 (I357387,I2683,I175343,I175403,);
not I_10158 (I175411,I357381);
nand I_10159 (I175428,I175411,I357384);
not I_10160 (I175445,I175428);
nor I_10161 (I175462,I175445,I357402);
nor I_10162 (I175479,I175377,I175462);
DFFARX1 I_10163 (I175479,I2683,I175343,I175329,);
not I_10164 (I175510,I357402);
nand I_10165 (I175527,I175510,I175445);
and I_10166 (I175544,I175510,I357405);
nand I_10167 (I175561,I175544,I357384);
nor I_10168 (I175326,I175561,I175510);
and I_10169 (I175317,I175403,I175561);
not I_10170 (I175606,I175561);
nand I_10171 (I175320,I175403,I175606);
nor I_10172 (I175314,I175369,I175561);
not I_10173 (I175651,I357390);
nor I_10174 (I175668,I175651,I357405);
nand I_10175 (I175685,I175668,I175510);
nor I_10176 (I175323,I175428,I175685);
nor I_10177 (I175716,I175651,I357396);
and I_10178 (I175733,I175716,I357393);
or I_10179 (I175750,I175733,I357399);
DFFARX1 I_10180 (I175750,I2683,I175343,I175776,);
nor I_10181 (I175784,I175776,I175527);
DFFARX1 I_10182 (I175784,I2683,I175343,I175311,);
DFFARX1 I_10183 (I175776,I2683,I175343,I175335,);
not I_10184 (I175829,I175776);
nor I_10185 (I175846,I175829,I175403);
nor I_10186 (I175863,I175668,I175846);
DFFARX1 I_10187 (I175863,I2683,I175343,I175332,);
not I_10188 (I175921,I2690);
DFFARX1 I_10189 (I66169,I2683,I175921,I175947,);
not I_10190 (I175955,I175947);
DFFARX1 I_10191 (I66154,I2683,I175921,I175981,);
not I_10192 (I175989,I66172);
nand I_10193 (I176006,I175989,I66157);
not I_10194 (I176023,I176006);
nor I_10195 (I176040,I176023,I66154);
nor I_10196 (I176057,I175955,I176040);
DFFARX1 I_10197 (I176057,I2683,I175921,I175907,);
not I_10198 (I176088,I66154);
nand I_10199 (I176105,I176088,I176023);
and I_10200 (I176122,I176088,I66157);
nand I_10201 (I176139,I176122,I66178);
nor I_10202 (I175904,I176139,I176088);
and I_10203 (I175895,I175981,I176139);
not I_10204 (I176184,I176139);
nand I_10205 (I175898,I175981,I176184);
nor I_10206 (I175892,I175947,I176139);
not I_10207 (I176229,I66166);
nor I_10208 (I176246,I176229,I66157);
nand I_10209 (I176263,I176246,I176088);
nor I_10210 (I175901,I176006,I176263);
nor I_10211 (I176294,I176229,I66160);
and I_10212 (I176311,I176294,I66175);
or I_10213 (I176328,I176311,I66163);
DFFARX1 I_10214 (I176328,I2683,I175921,I176354,);
nor I_10215 (I176362,I176354,I176105);
DFFARX1 I_10216 (I176362,I2683,I175921,I175889,);
DFFARX1 I_10217 (I176354,I2683,I175921,I175913,);
not I_10218 (I176407,I176354);
nor I_10219 (I176424,I176407,I175981);
nor I_10220 (I176441,I176246,I176424);
DFFARX1 I_10221 (I176441,I2683,I175921,I175910,);
not I_10222 (I176499,I2690);
DFFARX1 I_10223 (I85209,I2683,I176499,I176525,);
not I_10224 (I176533,I176525);
DFFARX1 I_10225 (I85194,I2683,I176499,I176559,);
not I_10226 (I176567,I85212);
nand I_10227 (I176584,I176567,I85197);
not I_10228 (I176601,I176584);
nor I_10229 (I176618,I176601,I85194);
nor I_10230 (I176635,I176533,I176618);
DFFARX1 I_10231 (I176635,I2683,I176499,I176485,);
not I_10232 (I176666,I85194);
nand I_10233 (I176683,I176666,I176601);
and I_10234 (I176700,I176666,I85197);
nand I_10235 (I176717,I176700,I85218);
nor I_10236 (I176482,I176717,I176666);
and I_10237 (I176473,I176559,I176717);
not I_10238 (I176762,I176717);
nand I_10239 (I176476,I176559,I176762);
nor I_10240 (I176470,I176525,I176717);
not I_10241 (I176807,I85206);
nor I_10242 (I176824,I176807,I85197);
nand I_10243 (I176841,I176824,I176666);
nor I_10244 (I176479,I176584,I176841);
nor I_10245 (I176872,I176807,I85200);
and I_10246 (I176889,I176872,I85215);
or I_10247 (I176906,I176889,I85203);
DFFARX1 I_10248 (I176906,I2683,I176499,I176932,);
nor I_10249 (I176940,I176932,I176683);
DFFARX1 I_10250 (I176940,I2683,I176499,I176467,);
DFFARX1 I_10251 (I176932,I2683,I176499,I176491,);
not I_10252 (I176985,I176932);
nor I_10253 (I177002,I176985,I176559);
nor I_10254 (I177019,I176824,I177002);
DFFARX1 I_10255 (I177019,I2683,I176499,I176488,);
not I_10256 (I177077,I2690);
DFFARX1 I_10257 (I369775,I2683,I177077,I177103,);
not I_10258 (I177111,I177103);
DFFARX1 I_10259 (I369769,I2683,I177077,I177137,);
not I_10260 (I177145,I369778);
nand I_10261 (I177162,I177145,I369757);
not I_10262 (I177179,I177162);
nor I_10263 (I177196,I177179,I369766);
nor I_10264 (I177213,I177111,I177196);
DFFARX1 I_10265 (I177213,I2683,I177077,I177063,);
not I_10266 (I177244,I369766);
nand I_10267 (I177261,I177244,I177179);
and I_10268 (I177278,I177244,I369781);
nand I_10269 (I177295,I177278,I369760);
nor I_10270 (I177060,I177295,I177244);
and I_10271 (I177051,I177137,I177295);
not I_10272 (I177340,I177295);
nand I_10273 (I177054,I177137,I177340);
nor I_10274 (I177048,I177103,I177295);
not I_10275 (I177385,I369763);
nor I_10276 (I177402,I177385,I369781);
nand I_10277 (I177419,I177402,I177244);
nor I_10278 (I177057,I177162,I177419);
nor I_10279 (I177450,I177385,I369772);
and I_10280 (I177467,I177450,I369760);
or I_10281 (I177484,I177467,I369757);
DFFARX1 I_10282 (I177484,I2683,I177077,I177510,);
nor I_10283 (I177518,I177510,I177261);
DFFARX1 I_10284 (I177518,I2683,I177077,I177045,);
DFFARX1 I_10285 (I177510,I2683,I177077,I177069,);
not I_10286 (I177563,I177510);
nor I_10287 (I177580,I177563,I177137);
nor I_10288 (I177597,I177402,I177580);
DFFARX1 I_10289 (I177597,I2683,I177077,I177066,);
not I_10290 (I177655,I2690);
DFFARX1 I_10291 (I375215,I2683,I177655,I177681,);
not I_10292 (I177689,I177681);
DFFARX1 I_10293 (I375209,I2683,I177655,I177715,);
not I_10294 (I177723,I375218);
nand I_10295 (I177740,I177723,I375197);
not I_10296 (I177757,I177740);
nor I_10297 (I177774,I177757,I375206);
nor I_10298 (I177791,I177689,I177774);
DFFARX1 I_10299 (I177791,I2683,I177655,I177641,);
not I_10300 (I177822,I375206);
nand I_10301 (I177839,I177822,I177757);
and I_10302 (I177856,I177822,I375221);
nand I_10303 (I177873,I177856,I375200);
nor I_10304 (I177638,I177873,I177822);
and I_10305 (I177629,I177715,I177873);
not I_10306 (I177918,I177873);
nand I_10307 (I177632,I177715,I177918);
nor I_10308 (I177626,I177681,I177873);
not I_10309 (I177963,I375203);
nor I_10310 (I177980,I177963,I375221);
nand I_10311 (I177997,I177980,I177822);
nor I_10312 (I177635,I177740,I177997);
nor I_10313 (I178028,I177963,I375212);
and I_10314 (I178045,I178028,I375200);
or I_10315 (I178062,I178045,I375197);
DFFARX1 I_10316 (I178062,I2683,I177655,I178088,);
nor I_10317 (I178096,I178088,I177839);
DFFARX1 I_10318 (I178096,I2683,I177655,I177623,);
DFFARX1 I_10319 (I178088,I2683,I177655,I177647,);
not I_10320 (I178141,I178088);
nor I_10321 (I178158,I178141,I177715);
nor I_10322 (I178175,I177980,I178158);
DFFARX1 I_10323 (I178175,I2683,I177655,I177644,);
not I_10324 (I178233,I2690);
DFFARX1 I_10325 (I243436,I2683,I178233,I178259,);
not I_10326 (I178267,I178259);
DFFARX1 I_10327 (I243436,I2683,I178233,I178293,);
not I_10328 (I178301,I243433);
nand I_10329 (I178318,I178301,I243448);
not I_10330 (I178335,I178318);
nor I_10331 (I178352,I178335,I243442);
nor I_10332 (I178369,I178267,I178352);
DFFARX1 I_10333 (I178369,I2683,I178233,I178219,);
not I_10334 (I178400,I243442);
nand I_10335 (I178417,I178400,I178335);
and I_10336 (I178434,I178400,I243439);
nand I_10337 (I178451,I178434,I243430);
nor I_10338 (I178216,I178451,I178400);
and I_10339 (I178207,I178293,I178451);
not I_10340 (I178496,I178451);
nand I_10341 (I178210,I178293,I178496);
nor I_10342 (I178204,I178259,I178451);
not I_10343 (I178541,I243451);
nor I_10344 (I178558,I178541,I243439);
nand I_10345 (I178575,I178558,I178400);
nor I_10346 (I178213,I178318,I178575);
nor I_10347 (I178606,I178541,I243430);
and I_10348 (I178623,I178606,I243433);
or I_10349 (I178640,I178623,I243445);
DFFARX1 I_10350 (I178640,I2683,I178233,I178666,);
nor I_10351 (I178674,I178666,I178417);
DFFARX1 I_10352 (I178674,I2683,I178233,I178201,);
DFFARX1 I_10353 (I178666,I2683,I178233,I178225,);
not I_10354 (I178719,I178666);
nor I_10355 (I178736,I178719,I178293);
nor I_10356 (I178753,I178558,I178736);
DFFARX1 I_10357 (I178753,I2683,I178233,I178222,);
not I_10358 (I178811,I2690);
DFFARX1 I_10359 (I67954,I2683,I178811,I178837,);
not I_10360 (I178845,I178837);
DFFARX1 I_10361 (I67939,I2683,I178811,I178871,);
not I_10362 (I178879,I67957);
nand I_10363 (I178896,I178879,I67942);
not I_10364 (I178913,I178896);
nor I_10365 (I178930,I178913,I67939);
nor I_10366 (I178947,I178845,I178930);
DFFARX1 I_10367 (I178947,I2683,I178811,I178797,);
not I_10368 (I178978,I67939);
nand I_10369 (I178995,I178978,I178913);
and I_10370 (I179012,I178978,I67942);
nand I_10371 (I179029,I179012,I67963);
nor I_10372 (I178794,I179029,I178978);
and I_10373 (I178785,I178871,I179029);
not I_10374 (I179074,I179029);
nand I_10375 (I178788,I178871,I179074);
nor I_10376 (I178782,I178837,I179029);
not I_10377 (I179119,I67951);
nor I_10378 (I179136,I179119,I67942);
nand I_10379 (I179153,I179136,I178978);
nor I_10380 (I178791,I178896,I179153);
nor I_10381 (I179184,I179119,I67945);
and I_10382 (I179201,I179184,I67960);
or I_10383 (I179218,I179201,I67948);
DFFARX1 I_10384 (I179218,I2683,I178811,I179244,);
nor I_10385 (I179252,I179244,I178995);
DFFARX1 I_10386 (I179252,I2683,I178811,I178779,);
DFFARX1 I_10387 (I179244,I2683,I178811,I178803,);
not I_10388 (I179297,I179244);
nor I_10389 (I179314,I179297,I178871);
nor I_10390 (I179331,I179136,I179314);
DFFARX1 I_10391 (I179331,I2683,I178811,I178800,);
not I_10392 (I179389,I2690);
DFFARX1 I_10393 (I151387,I2683,I179389,I179415,);
not I_10394 (I179423,I179415);
DFFARX1 I_10395 (I151399,I2683,I179389,I179449,);
not I_10396 (I179457,I151375);
nand I_10397 (I179474,I179457,I151402);
not I_10398 (I179491,I179474);
nor I_10399 (I179508,I179491,I151390);
nor I_10400 (I179525,I179423,I179508);
DFFARX1 I_10401 (I179525,I2683,I179389,I179375,);
not I_10402 (I179556,I151390);
nand I_10403 (I179573,I179556,I179491);
and I_10404 (I179590,I179556,I151375);
nand I_10405 (I179607,I179590,I151378);
nor I_10406 (I179372,I179607,I179556);
and I_10407 (I179363,I179449,I179607);
not I_10408 (I179652,I179607);
nand I_10409 (I179366,I179449,I179652);
nor I_10410 (I179360,I179415,I179607);
not I_10411 (I179697,I151384);
nor I_10412 (I179714,I179697,I151375);
nand I_10413 (I179731,I179714,I179556);
nor I_10414 (I179369,I179474,I179731);
nor I_10415 (I179762,I179697,I151393);
and I_10416 (I179779,I179762,I151381);
or I_10417 (I179796,I179779,I151396);
DFFARX1 I_10418 (I179796,I2683,I179389,I179822,);
nor I_10419 (I179830,I179822,I179573);
DFFARX1 I_10420 (I179830,I2683,I179389,I179357,);
DFFARX1 I_10421 (I179822,I2683,I179389,I179381,);
not I_10422 (I179875,I179822);
nor I_10423 (I179892,I179875,I179449);
nor I_10424 (I179909,I179714,I179892);
DFFARX1 I_10425 (I179909,I2683,I179389,I179378,);
not I_10426 (I179967,I2690);
DFFARX1 I_10427 (I112672,I2683,I179967,I179993,);
not I_10428 (I180001,I179993);
DFFARX1 I_10429 (I112687,I2683,I179967,I180027,);
not I_10430 (I180035,I112690);
nand I_10431 (I180052,I180035,I112669);
not I_10432 (I180069,I180052);
nor I_10433 (I180086,I180069,I112693);
nor I_10434 (I180103,I180001,I180086);
DFFARX1 I_10435 (I180103,I2683,I179967,I179953,);
not I_10436 (I180134,I112693);
nand I_10437 (I180151,I180134,I180069);
and I_10438 (I180168,I180134,I112675);
nand I_10439 (I180185,I180168,I112666);
nor I_10440 (I179950,I180185,I180134);
and I_10441 (I179941,I180027,I180185);
not I_10442 (I180230,I180185);
nand I_10443 (I179944,I180027,I180230);
nor I_10444 (I179938,I179993,I180185);
not I_10445 (I180275,I112666);
nor I_10446 (I180292,I180275,I112675);
nand I_10447 (I180309,I180292,I180134);
nor I_10448 (I179947,I180052,I180309);
nor I_10449 (I180340,I180275,I112681);
and I_10450 (I180357,I180340,I112684);
or I_10451 (I180374,I180357,I112678);
DFFARX1 I_10452 (I180374,I2683,I179967,I180400,);
nor I_10453 (I180408,I180400,I180151);
DFFARX1 I_10454 (I180408,I2683,I179967,I179935,);
DFFARX1 I_10455 (I180400,I2683,I179967,I179959,);
not I_10456 (I180453,I180400);
nor I_10457 (I180470,I180453,I180027);
nor I_10458 (I180487,I180292,I180470);
DFFARX1 I_10459 (I180487,I2683,I179967,I179956,);
not I_10460 (I180545,I2690);
DFFARX1 I_10461 (I76284,I2683,I180545,I180571,);
not I_10462 (I180579,I180571);
DFFARX1 I_10463 (I76269,I2683,I180545,I180605,);
not I_10464 (I180613,I76287);
nand I_10465 (I180630,I180613,I76272);
not I_10466 (I180647,I180630);
nor I_10467 (I180664,I180647,I76269);
nor I_10468 (I180681,I180579,I180664);
DFFARX1 I_10469 (I180681,I2683,I180545,I180531,);
not I_10470 (I180712,I76269);
nand I_10471 (I180729,I180712,I180647);
and I_10472 (I180746,I180712,I76272);
nand I_10473 (I180763,I180746,I76293);
nor I_10474 (I180528,I180763,I180712);
and I_10475 (I180519,I180605,I180763);
not I_10476 (I180808,I180763);
nand I_10477 (I180522,I180605,I180808);
nor I_10478 (I180516,I180571,I180763);
not I_10479 (I180853,I76281);
nor I_10480 (I180870,I180853,I76272);
nand I_10481 (I180887,I180870,I180712);
nor I_10482 (I180525,I180630,I180887);
nor I_10483 (I180918,I180853,I76275);
and I_10484 (I180935,I180918,I76290);
or I_10485 (I180952,I180935,I76278);
DFFARX1 I_10486 (I180952,I2683,I180545,I180978,);
nor I_10487 (I180986,I180978,I180729);
DFFARX1 I_10488 (I180986,I2683,I180545,I180513,);
DFFARX1 I_10489 (I180978,I2683,I180545,I180537,);
not I_10490 (I181031,I180978);
nor I_10491 (I181048,I181031,I180605);
nor I_10492 (I181065,I180870,I181048);
DFFARX1 I_10493 (I181065,I2683,I180545,I180534,);
not I_10494 (I181123,I2690);
DFFARX1 I_10495 (I405729,I2683,I181123,I181149,);
not I_10496 (I181157,I181149);
DFFARX1 I_10497 (I405729,I2683,I181123,I181183,);
not I_10498 (I181191,I405753);
nand I_10499 (I181208,I181191,I405735);
not I_10500 (I181225,I181208);
nor I_10501 (I181242,I181225,I405750);
nor I_10502 (I181259,I181157,I181242);
DFFARX1 I_10503 (I181259,I2683,I181123,I181109,);
not I_10504 (I181290,I405750);
nand I_10505 (I181307,I181290,I181225);
and I_10506 (I181324,I181290,I405732);
nand I_10507 (I181341,I181324,I405741);
nor I_10508 (I181106,I181341,I181290);
and I_10509 (I181097,I181183,I181341);
not I_10510 (I181386,I181341);
nand I_10511 (I181100,I181183,I181386);
nor I_10512 (I181094,I181149,I181341);
not I_10513 (I181431,I405738);
nor I_10514 (I181448,I181431,I405732);
nand I_10515 (I181465,I181448,I181290);
nor I_10516 (I181103,I181208,I181465);
nor I_10517 (I181496,I181431,I405747);
and I_10518 (I181513,I181496,I405756);
or I_10519 (I181530,I181513,I405744);
DFFARX1 I_10520 (I181530,I2683,I181123,I181556,);
nor I_10521 (I181564,I181556,I181307);
DFFARX1 I_10522 (I181564,I2683,I181123,I181091,);
DFFARX1 I_10523 (I181556,I2683,I181123,I181115,);
not I_10524 (I181609,I181556);
nor I_10525 (I181626,I181609,I181183);
nor I_10526 (I181643,I181448,I181626);
DFFARX1 I_10527 (I181643,I2683,I181123,I181112,);
not I_10528 (I181701,I2690);
DFFARX1 I_10529 (I214615,I2683,I181701,I181727,);
not I_10530 (I181735,I181727);
DFFARX1 I_10531 (I214627,I2683,I181701,I181761,);
not I_10532 (I181769,I214618);
nand I_10533 (I181786,I181769,I214621);
not I_10534 (I181803,I181786);
nor I_10535 (I181820,I181803,I214624);
nor I_10536 (I181837,I181735,I181820);
DFFARX1 I_10537 (I181837,I2683,I181701,I181687,);
not I_10538 (I181868,I214624);
nand I_10539 (I181885,I181868,I181803);
and I_10540 (I181902,I181868,I214618);
nand I_10541 (I181919,I181902,I214630);
nor I_10542 (I181684,I181919,I181868);
and I_10543 (I181675,I181761,I181919);
not I_10544 (I181964,I181919);
nand I_10545 (I181678,I181761,I181964);
nor I_10546 (I181672,I181727,I181919);
not I_10547 (I182009,I214636);
nor I_10548 (I182026,I182009,I214618);
nand I_10549 (I182043,I182026,I181868);
nor I_10550 (I181681,I181786,I182043);
nor I_10551 (I182074,I182009,I214615);
and I_10552 (I182091,I182074,I214633);
or I_10553 (I182108,I182091,I214639);
DFFARX1 I_10554 (I182108,I2683,I181701,I182134,);
nor I_10555 (I182142,I182134,I181885);
DFFARX1 I_10556 (I182142,I2683,I181701,I181669,);
DFFARX1 I_10557 (I182134,I2683,I181701,I181693,);
not I_10558 (I182187,I182134);
nor I_10559 (I182204,I182187,I181761);
nor I_10560 (I182221,I182026,I182204);
DFFARX1 I_10561 (I182221,I2683,I181701,I181690,);
not I_10562 (I182279,I2690);
DFFARX1 I_10563 (I105821,I2683,I182279,I182305,);
not I_10564 (I182313,I182305);
DFFARX1 I_10565 (I105836,I2683,I182279,I182339,);
not I_10566 (I182347,I105839);
nand I_10567 (I182364,I182347,I105818);
not I_10568 (I182381,I182364);
nor I_10569 (I182398,I182381,I105842);
nor I_10570 (I182415,I182313,I182398);
DFFARX1 I_10571 (I182415,I2683,I182279,I182265,);
not I_10572 (I182446,I105842);
nand I_10573 (I182463,I182446,I182381);
and I_10574 (I182480,I182446,I105824);
nand I_10575 (I182497,I182480,I105815);
nor I_10576 (I182262,I182497,I182446);
and I_10577 (I182253,I182339,I182497);
not I_10578 (I182542,I182497);
nand I_10579 (I182256,I182339,I182542);
nor I_10580 (I182250,I182305,I182497);
not I_10581 (I182587,I105815);
nor I_10582 (I182604,I182587,I105824);
nand I_10583 (I182621,I182604,I182446);
nor I_10584 (I182259,I182364,I182621);
nor I_10585 (I182652,I182587,I105830);
and I_10586 (I182669,I182652,I105833);
or I_10587 (I182686,I182669,I105827);
DFFARX1 I_10588 (I182686,I2683,I182279,I182712,);
nor I_10589 (I182720,I182712,I182463);
DFFARX1 I_10590 (I182720,I2683,I182279,I182247,);
DFFARX1 I_10591 (I182712,I2683,I182279,I182271,);
not I_10592 (I182765,I182712);
nor I_10593 (I182782,I182765,I182339);
nor I_10594 (I182799,I182604,I182782);
DFFARX1 I_10595 (I182799,I2683,I182279,I182268,);
not I_10596 (I182857,I2690);
DFFARX1 I_10597 (I123739,I2683,I182857,I182883,);
not I_10598 (I182891,I182883);
DFFARX1 I_10599 (I123754,I2683,I182857,I182917,);
not I_10600 (I182925,I123757);
nand I_10601 (I182942,I182925,I123736);
not I_10602 (I182959,I182942);
nor I_10603 (I182976,I182959,I123760);
nor I_10604 (I182993,I182891,I182976);
DFFARX1 I_10605 (I182993,I2683,I182857,I182843,);
not I_10606 (I183024,I123760);
nand I_10607 (I183041,I183024,I182959);
and I_10608 (I183058,I183024,I123742);
nand I_10609 (I183075,I183058,I123733);
nor I_10610 (I182840,I183075,I183024);
and I_10611 (I182831,I182917,I183075);
not I_10612 (I183120,I183075);
nand I_10613 (I182834,I182917,I183120);
nor I_10614 (I182828,I182883,I183075);
not I_10615 (I183165,I123733);
nor I_10616 (I183182,I183165,I123742);
nand I_10617 (I183199,I183182,I183024);
nor I_10618 (I182837,I182942,I183199);
nor I_10619 (I183230,I183165,I123748);
and I_10620 (I183247,I183230,I123751);
or I_10621 (I183264,I183247,I123745);
DFFARX1 I_10622 (I183264,I2683,I182857,I183290,);
nor I_10623 (I183298,I183290,I183041);
DFFARX1 I_10624 (I183298,I2683,I182857,I182825,);
DFFARX1 I_10625 (I183290,I2683,I182857,I182849,);
not I_10626 (I183343,I183290);
nor I_10627 (I183360,I183343,I182917);
nor I_10628 (I183377,I183182,I183360);
DFFARX1 I_10629 (I183377,I2683,I182857,I182846,);
not I_10630 (I183435,I2690);
DFFARX1 I_10631 (I20448,I2683,I183435,I183461,);
not I_10632 (I183469,I183461);
DFFARX1 I_10633 (I20427,I2683,I183435,I183495,);
not I_10634 (I183503,I20424);
nand I_10635 (I183520,I183503,I20439);
not I_10636 (I183537,I183520);
nor I_10637 (I183554,I183537,I20427);
nor I_10638 (I183571,I183469,I183554);
DFFARX1 I_10639 (I183571,I2683,I183435,I183421,);
not I_10640 (I183602,I20427);
nand I_10641 (I183619,I183602,I183537);
and I_10642 (I183636,I183602,I20430);
nand I_10643 (I183653,I183636,I20445);
nor I_10644 (I183418,I183653,I183602);
and I_10645 (I183409,I183495,I183653);
not I_10646 (I183698,I183653);
nand I_10647 (I183412,I183495,I183698);
nor I_10648 (I183406,I183461,I183653);
not I_10649 (I183743,I20436);
nor I_10650 (I183760,I183743,I20430);
nand I_10651 (I183777,I183760,I183602);
nor I_10652 (I183415,I183520,I183777);
nor I_10653 (I183808,I183743,I20424);
and I_10654 (I183825,I183808,I20433);
or I_10655 (I183842,I183825,I20442);
DFFARX1 I_10656 (I183842,I2683,I183435,I183868,);
nor I_10657 (I183876,I183868,I183619);
DFFARX1 I_10658 (I183876,I2683,I183435,I183403,);
DFFARX1 I_10659 (I183868,I2683,I183435,I183427,);
not I_10660 (I183921,I183868);
nor I_10661 (I183938,I183921,I183495);
nor I_10662 (I183955,I183760,I183938);
DFFARX1 I_10663 (I183955,I2683,I183435,I183424,);
not I_10664 (I184013,I2690);
DFFARX1 I_10665 (I142683,I2683,I184013,I184039,);
not I_10666 (I184047,I184039);
DFFARX1 I_10667 (I142695,I2683,I184013,I184073,);
not I_10668 (I184081,I142671);
nand I_10669 (I184098,I184081,I142698);
not I_10670 (I184115,I184098);
nor I_10671 (I184132,I184115,I142686);
nor I_10672 (I184149,I184047,I184132);
DFFARX1 I_10673 (I184149,I2683,I184013,I183999,);
not I_10674 (I184180,I142686);
nand I_10675 (I184197,I184180,I184115);
and I_10676 (I184214,I184180,I142671);
nand I_10677 (I184231,I184214,I142674);
nor I_10678 (I183996,I184231,I184180);
and I_10679 (I183987,I184073,I184231);
not I_10680 (I184276,I184231);
nand I_10681 (I183990,I184073,I184276);
nor I_10682 (I183984,I184039,I184231);
not I_10683 (I184321,I142680);
nor I_10684 (I184338,I184321,I142671);
nand I_10685 (I184355,I184338,I184180);
nor I_10686 (I183993,I184098,I184355);
nor I_10687 (I184386,I184321,I142689);
and I_10688 (I184403,I184386,I142677);
or I_10689 (I184420,I184403,I142692);
DFFARX1 I_10690 (I184420,I2683,I184013,I184446,);
nor I_10691 (I184454,I184446,I184197);
DFFARX1 I_10692 (I184454,I2683,I184013,I183981,);
DFFARX1 I_10693 (I184446,I2683,I184013,I184005,);
not I_10694 (I184499,I184446);
nor I_10695 (I184516,I184499,I184073);
nor I_10696 (I184533,I184338,I184516);
DFFARX1 I_10697 (I184533,I2683,I184013,I184002,);
not I_10698 (I184591,I2690);
DFFARX1 I_10699 (I36258,I2683,I184591,I184617,);
not I_10700 (I184625,I184617);
DFFARX1 I_10701 (I36237,I2683,I184591,I184651,);
not I_10702 (I184659,I36234);
nand I_10703 (I184676,I184659,I36249);
not I_10704 (I184693,I184676);
nor I_10705 (I184710,I184693,I36237);
nor I_10706 (I184727,I184625,I184710);
DFFARX1 I_10707 (I184727,I2683,I184591,I184577,);
not I_10708 (I184758,I36237);
nand I_10709 (I184775,I184758,I184693);
and I_10710 (I184792,I184758,I36240);
nand I_10711 (I184809,I184792,I36255);
nor I_10712 (I184574,I184809,I184758);
and I_10713 (I184565,I184651,I184809);
not I_10714 (I184854,I184809);
nand I_10715 (I184568,I184651,I184854);
nor I_10716 (I184562,I184617,I184809);
not I_10717 (I184899,I36246);
nor I_10718 (I184916,I184899,I36240);
nand I_10719 (I184933,I184916,I184758);
nor I_10720 (I184571,I184676,I184933);
nor I_10721 (I184964,I184899,I36234);
and I_10722 (I184981,I184964,I36243);
or I_10723 (I184998,I184981,I36252);
DFFARX1 I_10724 (I184998,I2683,I184591,I185024,);
nor I_10725 (I185032,I185024,I184775);
DFFARX1 I_10726 (I185032,I2683,I184591,I184559,);
DFFARX1 I_10727 (I185024,I2683,I184591,I184583,);
not I_10728 (I185077,I185024);
nor I_10729 (I185094,I185077,I184651);
nor I_10730 (I185111,I184916,I185094);
DFFARX1 I_10731 (I185111,I2683,I184591,I184580,);
not I_10732 (I185169,I2690);
DFFARX1 I_10733 (I251341,I2683,I185169,I185195,);
not I_10734 (I185203,I185195);
DFFARX1 I_10735 (I251341,I2683,I185169,I185229,);
not I_10736 (I185237,I251338);
nand I_10737 (I185254,I185237,I251353);
not I_10738 (I185271,I185254);
nor I_10739 (I185288,I185271,I251347);
nor I_10740 (I185305,I185203,I185288);
DFFARX1 I_10741 (I185305,I2683,I185169,I185155,);
not I_10742 (I185336,I251347);
nand I_10743 (I185353,I185336,I185271);
and I_10744 (I185370,I185336,I251344);
nand I_10745 (I185387,I185370,I251335);
nor I_10746 (I185152,I185387,I185336);
and I_10747 (I185143,I185229,I185387);
not I_10748 (I185432,I185387);
nand I_10749 (I185146,I185229,I185432);
nor I_10750 (I185140,I185195,I185387);
not I_10751 (I185477,I251356);
nor I_10752 (I185494,I185477,I251344);
nand I_10753 (I185511,I185494,I185336);
nor I_10754 (I185149,I185254,I185511);
nor I_10755 (I185542,I185477,I251335);
and I_10756 (I185559,I185542,I251338);
or I_10757 (I185576,I185559,I251350);
DFFARX1 I_10758 (I185576,I2683,I185169,I185602,);
nor I_10759 (I185610,I185602,I185353);
DFFARX1 I_10760 (I185610,I2683,I185169,I185137,);
DFFARX1 I_10761 (I185602,I2683,I185169,I185161,);
not I_10762 (I185655,I185602);
nor I_10763 (I185672,I185655,I185229);
nor I_10764 (I185689,I185494,I185672);
DFFARX1 I_10765 (I185689,I2683,I185169,I185158,);
not I_10766 (I185747,I2690);
DFFARX1 I_10767 (I161782,I2683,I185747,I185773,);
not I_10768 (I185781,I185773);
DFFARX1 I_10769 (I161794,I2683,I185747,I185807,);
not I_10770 (I185815,I161800);
nand I_10771 (I185832,I185815,I161791);
not I_10772 (I185849,I185832);
nor I_10773 (I185866,I185849,I161797);
nor I_10774 (I185883,I185781,I185866);
DFFARX1 I_10775 (I185883,I2683,I185747,I185733,);
not I_10776 (I185914,I161797);
nand I_10777 (I185931,I185914,I185849);
and I_10778 (I185948,I185914,I161788);
nand I_10779 (I185965,I185948,I161779);
nor I_10780 (I185730,I185965,I185914);
and I_10781 (I185721,I185807,I185965);
not I_10782 (I186010,I185965);
nand I_10783 (I185724,I185807,I186010);
nor I_10784 (I185718,I185773,I185965);
not I_10785 (I186055,I161785);
nor I_10786 (I186072,I186055,I161788);
nand I_10787 (I186089,I186072,I185914);
nor I_10788 (I185727,I185832,I186089);
nor I_10789 (I186120,I186055,I161782);
and I_10790 (I186137,I186120,I161779);
or I_10791 (I186154,I186137,I161803);
DFFARX1 I_10792 (I186154,I2683,I185747,I186180,);
nor I_10793 (I186188,I186180,I185931);
DFFARX1 I_10794 (I186188,I2683,I185747,I185715,);
DFFARX1 I_10795 (I186180,I2683,I185747,I185739,);
not I_10796 (I186233,I186180);
nor I_10797 (I186250,I186233,I185807);
nor I_10798 (I186267,I186072,I186250);
DFFARX1 I_10799 (I186267,I2683,I185747,I185736,);
not I_10800 (I186325,I2690);
DFFARX1 I_10801 (I73309,I2683,I186325,I186351,);
not I_10802 (I186359,I186351);
DFFARX1 I_10803 (I73294,I2683,I186325,I186385,);
not I_10804 (I186393,I73312);
nand I_10805 (I186410,I186393,I73297);
not I_10806 (I186427,I186410);
nor I_10807 (I186444,I186427,I73294);
nor I_10808 (I186461,I186359,I186444);
DFFARX1 I_10809 (I186461,I2683,I186325,I186311,);
not I_10810 (I186492,I73294);
nand I_10811 (I186509,I186492,I186427);
and I_10812 (I186526,I186492,I73297);
nand I_10813 (I186543,I186526,I73318);
nor I_10814 (I186308,I186543,I186492);
and I_10815 (I186299,I186385,I186543);
not I_10816 (I186588,I186543);
nand I_10817 (I186302,I186385,I186588);
nor I_10818 (I186296,I186351,I186543);
not I_10819 (I186633,I73306);
nor I_10820 (I186650,I186633,I73297);
nand I_10821 (I186667,I186650,I186492);
nor I_10822 (I186305,I186410,I186667);
nor I_10823 (I186698,I186633,I73300);
and I_10824 (I186715,I186698,I73315);
or I_10825 (I186732,I186715,I73303);
DFFARX1 I_10826 (I186732,I2683,I186325,I186758,);
nor I_10827 (I186766,I186758,I186509);
DFFARX1 I_10828 (I186766,I2683,I186325,I186293,);
DFFARX1 I_10829 (I186758,I2683,I186325,I186317,);
not I_10830 (I186811,I186758);
nor I_10831 (I186828,I186811,I186385);
nor I_10832 (I186845,I186650,I186828);
DFFARX1 I_10833 (I186845,I2683,I186325,I186314,);
not I_10834 (I186903,I2690);
DFFARX1 I_10835 (I232533,I2683,I186903,I186929,);
not I_10836 (I186937,I186929);
DFFARX1 I_10837 (I232545,I2683,I186903,I186963,);
not I_10838 (I186971,I232536);
nand I_10839 (I186988,I186971,I232539);
not I_10840 (I187005,I186988);
nor I_10841 (I187022,I187005,I232542);
nor I_10842 (I187039,I186937,I187022);
DFFARX1 I_10843 (I187039,I2683,I186903,I186889,);
not I_10844 (I187070,I232542);
nand I_10845 (I187087,I187070,I187005);
and I_10846 (I187104,I187070,I232536);
nand I_10847 (I187121,I187104,I232548);
nor I_10848 (I186886,I187121,I187070);
and I_10849 (I186877,I186963,I187121);
not I_10850 (I187166,I187121);
nand I_10851 (I186880,I186963,I187166);
nor I_10852 (I186874,I186929,I187121);
not I_10853 (I187211,I232554);
nor I_10854 (I187228,I187211,I232536);
nand I_10855 (I187245,I187228,I187070);
nor I_10856 (I186883,I186988,I187245);
nor I_10857 (I187276,I187211,I232533);
and I_10858 (I187293,I187276,I232551);
or I_10859 (I187310,I187293,I232557);
DFFARX1 I_10860 (I187310,I2683,I186903,I187336,);
nor I_10861 (I187344,I187336,I187087);
DFFARX1 I_10862 (I187344,I2683,I186903,I186871,);
DFFARX1 I_10863 (I187336,I2683,I186903,I186895,);
not I_10864 (I187389,I187336);
nor I_10865 (I187406,I187389,I186963);
nor I_10866 (I187423,I187228,I187406);
DFFARX1 I_10867 (I187423,I2683,I186903,I186892,);
not I_10868 (I187481,I2690);
DFFARX1 I_10869 (I44755,I2683,I187481,I187507,);
not I_10870 (I187515,I187507);
DFFARX1 I_10871 (I44734,I2683,I187481,I187541,);
not I_10872 (I187549,I44734);
nand I_10873 (I187566,I187549,I44761);
not I_10874 (I187583,I187566);
nor I_10875 (I187600,I187583,I44737);
nor I_10876 (I187617,I187515,I187600);
DFFARX1 I_10877 (I187617,I2683,I187481,I187467,);
not I_10878 (I187648,I44737);
nand I_10879 (I187665,I187648,I187583);
and I_10880 (I187682,I187648,I44758);
nand I_10881 (I187699,I187682,I44740);
nor I_10882 (I187464,I187699,I187648);
and I_10883 (I187455,I187541,I187699);
not I_10884 (I187744,I187699);
nand I_10885 (I187458,I187541,I187744);
nor I_10886 (I187452,I187507,I187699);
not I_10887 (I187789,I44743);
nor I_10888 (I187806,I187789,I44758);
nand I_10889 (I187823,I187806,I187648);
nor I_10890 (I187461,I187566,I187823);
nor I_10891 (I187854,I187789,I44749);
and I_10892 (I187871,I187854,I44746);
or I_10893 (I187888,I187871,I44752);
DFFARX1 I_10894 (I187888,I2683,I187481,I187914,);
nor I_10895 (I187922,I187914,I187665);
DFFARX1 I_10896 (I187922,I2683,I187481,I187449,);
DFFARX1 I_10897 (I187914,I2683,I187481,I187473,);
not I_10898 (I187967,I187914);
nor I_10899 (I187984,I187967,I187541);
nor I_10900 (I188001,I187806,I187984);
DFFARX1 I_10901 (I188001,I2683,I187481,I187470,);
not I_10902 (I188059,I2690);
DFFARX1 I_10903 (I346977,I2683,I188059,I188085,);
not I_10904 (I188093,I188085);
DFFARX1 I_10905 (I346983,I2683,I188059,I188119,);
not I_10906 (I188127,I346977);
nand I_10907 (I188144,I188127,I346980);
not I_10908 (I188161,I188144);
nor I_10909 (I188178,I188161,I346998);
nor I_10910 (I188195,I188093,I188178);
DFFARX1 I_10911 (I188195,I2683,I188059,I188045,);
not I_10912 (I188226,I346998);
nand I_10913 (I188243,I188226,I188161);
and I_10914 (I188260,I188226,I347001);
nand I_10915 (I188277,I188260,I346980);
nor I_10916 (I188042,I188277,I188226);
and I_10917 (I188033,I188119,I188277);
not I_10918 (I188322,I188277);
nand I_10919 (I188036,I188119,I188322);
nor I_10920 (I188030,I188085,I188277);
not I_10921 (I188367,I346986);
nor I_10922 (I188384,I188367,I347001);
nand I_10923 (I188401,I188384,I188226);
nor I_10924 (I188039,I188144,I188401);
nor I_10925 (I188432,I188367,I346992);
and I_10926 (I188449,I188432,I346989);
or I_10927 (I188466,I188449,I346995);
DFFARX1 I_10928 (I188466,I2683,I188059,I188492,);
nor I_10929 (I188500,I188492,I188243);
DFFARX1 I_10930 (I188500,I2683,I188059,I188027,);
DFFARX1 I_10931 (I188492,I2683,I188059,I188051,);
not I_10932 (I188545,I188492);
nor I_10933 (I188562,I188545,I188119);
nor I_10934 (I188579,I188384,I188562);
DFFARX1 I_10935 (I188579,I2683,I188059,I188048,);
not I_10936 (I188637,I2690);
DFFARX1 I_10937 (I168922,I2683,I188637,I188663,);
not I_10938 (I188671,I188663);
DFFARX1 I_10939 (I168934,I2683,I188637,I188697,);
not I_10940 (I188705,I168940);
nand I_10941 (I188722,I188705,I168931);
not I_10942 (I188739,I188722);
nor I_10943 (I188756,I188739,I168937);
nor I_10944 (I188773,I188671,I188756);
DFFARX1 I_10945 (I188773,I2683,I188637,I188623,);
not I_10946 (I188804,I168937);
nand I_10947 (I188821,I188804,I188739);
and I_10948 (I188838,I188804,I168928);
nand I_10949 (I188855,I188838,I168919);
nor I_10950 (I188620,I188855,I188804);
and I_10951 (I188611,I188697,I188855);
not I_10952 (I188900,I188855);
nand I_10953 (I188614,I188697,I188900);
nor I_10954 (I188608,I188663,I188855);
not I_10955 (I188945,I168925);
nor I_10956 (I188962,I188945,I168928);
nand I_10957 (I188979,I188962,I188804);
nor I_10958 (I188617,I188722,I188979);
nor I_10959 (I189010,I188945,I168922);
and I_10960 (I189027,I189010,I168919);
or I_10961 (I189044,I189027,I168943);
DFFARX1 I_10962 (I189044,I2683,I188637,I189070,);
nor I_10963 (I189078,I189070,I188821);
DFFARX1 I_10964 (I189078,I2683,I188637,I188605,);
DFFARX1 I_10965 (I189070,I2683,I188637,I188629,);
not I_10966 (I189123,I189070);
nor I_10967 (I189140,I189123,I188697);
nor I_10968 (I189157,I188962,I189140);
DFFARX1 I_10969 (I189157,I2683,I188637,I188626,);
not I_10970 (I189215,I2690);
DFFARX1 I_10971 (I282060,I2683,I189215,I189241,);
not I_10972 (I189249,I189241);
DFFARX1 I_10973 (I282057,I2683,I189215,I189275,);
not I_10974 (I189283,I282054);
nand I_10975 (I189300,I189283,I282081);
not I_10976 (I189317,I189300);
nor I_10977 (I189334,I189317,I282069);
nor I_10978 (I189351,I189249,I189334);
DFFARX1 I_10979 (I189351,I2683,I189215,I189201,);
not I_10980 (I189382,I282069);
nand I_10981 (I189399,I189382,I189317);
and I_10982 (I189416,I189382,I282075);
nand I_10983 (I189433,I189416,I282066);
nor I_10984 (I189198,I189433,I189382);
and I_10985 (I189189,I189275,I189433);
not I_10986 (I189478,I189433);
nand I_10987 (I189192,I189275,I189478);
nor I_10988 (I189186,I189241,I189433);
not I_10989 (I189523,I282063);
nor I_10990 (I189540,I189523,I282075);
nand I_10991 (I189557,I189540,I189382);
nor I_10992 (I189195,I189300,I189557);
nor I_10993 (I189588,I189523,I282078);
and I_10994 (I189605,I189588,I282072);
or I_10995 (I189622,I189605,I282054);
DFFARX1 I_10996 (I189622,I2683,I189215,I189648,);
nor I_10997 (I189656,I189648,I189399);
DFFARX1 I_10998 (I189656,I2683,I189215,I189183,);
DFFARX1 I_10999 (I189648,I2683,I189215,I189207,);
not I_11000 (I189701,I189648);
nor I_11001 (I189718,I189701,I189275);
nor I_11002 (I189735,I189540,I189718);
DFFARX1 I_11003 (I189735,I2683,I189215,I189204,);
not I_11004 (I189793,I2690);
DFFARX1 I_11005 (I2028,I2683,I189793,I189819,);
not I_11006 (I189827,I189819);
DFFARX1 I_11007 (I2380,I2683,I189793,I189853,);
not I_11008 (I189861,I1924);
nand I_11009 (I189878,I189861,I1612);
not I_11010 (I189895,I189878);
nor I_11011 (I189912,I189895,I2628);
nor I_11012 (I189929,I189827,I189912);
DFFARX1 I_11013 (I189929,I2683,I189793,I189779,);
not I_11014 (I189960,I2628);
nand I_11015 (I189977,I189960,I189895);
and I_11016 (I189994,I189960,I1740);
nand I_11017 (I190011,I189994,I1972);
nor I_11018 (I189776,I190011,I189960);
and I_11019 (I189767,I189853,I190011);
not I_11020 (I190056,I190011);
nand I_11021 (I189770,I189853,I190056);
nor I_11022 (I189764,I189819,I190011);
not I_11023 (I190101,I2140);
nor I_11024 (I190118,I190101,I1740);
nand I_11025 (I190135,I190118,I189960);
nor I_11026 (I189773,I189878,I190135);
nor I_11027 (I190166,I190101,I2244);
and I_11028 (I190183,I190166,I1428);
or I_11029 (I190200,I190183,I2268);
DFFARX1 I_11030 (I190200,I2683,I189793,I190226,);
nor I_11031 (I190234,I190226,I189977);
DFFARX1 I_11032 (I190234,I2683,I189793,I189761,);
DFFARX1 I_11033 (I190226,I2683,I189793,I189785,);
not I_11034 (I190279,I190226);
nor I_11035 (I190296,I190279,I189853);
nor I_11036 (I190313,I190118,I190296);
DFFARX1 I_11037 (I190313,I2683,I189793,I189782,);
not I_11038 (I190371,I2690);
DFFARX1 I_11039 (I339463,I2683,I190371,I190397,);
not I_11040 (I190405,I190397);
DFFARX1 I_11041 (I339469,I2683,I190371,I190431,);
not I_11042 (I190439,I339463);
nand I_11043 (I190456,I190439,I339466);
not I_11044 (I190473,I190456);
nor I_11045 (I190490,I190473,I339484);
nor I_11046 (I190507,I190405,I190490);
DFFARX1 I_11047 (I190507,I2683,I190371,I190357,);
not I_11048 (I190538,I339484);
nand I_11049 (I190555,I190538,I190473);
and I_11050 (I190572,I190538,I339487);
nand I_11051 (I190589,I190572,I339466);
nor I_11052 (I190354,I190589,I190538);
and I_11053 (I190345,I190431,I190589);
not I_11054 (I190634,I190589);
nand I_11055 (I190348,I190431,I190634);
nor I_11056 (I190342,I190397,I190589);
not I_11057 (I190679,I339472);
nor I_11058 (I190696,I190679,I339487);
nand I_11059 (I190713,I190696,I190538);
nor I_11060 (I190351,I190456,I190713);
nor I_11061 (I190744,I190679,I339478);
and I_11062 (I190761,I190744,I339475);
or I_11063 (I190778,I190761,I339481);
DFFARX1 I_11064 (I190778,I2683,I190371,I190804,);
nor I_11065 (I190812,I190804,I190555);
DFFARX1 I_11066 (I190812,I2683,I190371,I190339,);
DFFARX1 I_11067 (I190804,I2683,I190371,I190363,);
not I_11068 (I190857,I190804);
nor I_11069 (I190874,I190857,I190431);
nor I_11070 (I190891,I190696,I190874);
DFFARX1 I_11071 (I190891,I2683,I190371,I190360,);
not I_11072 (I190949,I2690);
DFFARX1 I_11073 (I313219,I2683,I190949,I190975,);
not I_11074 (I190983,I190975);
DFFARX1 I_11075 (I313210,I2683,I190949,I191009,);
not I_11076 (I191017,I313204);
nand I_11077 (I191034,I191017,I313216);
not I_11078 (I191051,I191034);
nor I_11079 (I191068,I191051,I313207);
nor I_11080 (I191085,I190983,I191068);
DFFARX1 I_11081 (I191085,I2683,I190949,I190935,);
not I_11082 (I191116,I313207);
nand I_11083 (I191133,I191116,I191051);
and I_11084 (I191150,I191116,I313213);
nand I_11085 (I191167,I191150,I313198);
nor I_11086 (I190932,I191167,I191116);
and I_11087 (I190923,I191009,I191167);
not I_11088 (I191212,I191167);
nand I_11089 (I190926,I191009,I191212);
nor I_11090 (I190920,I190975,I191167);
not I_11091 (I191257,I313198);
nor I_11092 (I191274,I191257,I313213);
nand I_11093 (I191291,I191274,I191116);
nor I_11094 (I190929,I191034,I191291);
nor I_11095 (I191322,I191257,I313201);
and I_11096 (I191339,I191322,I313204);
or I_11097 (I191356,I191339,I313201);
DFFARX1 I_11098 (I191356,I2683,I190949,I191382,);
nor I_11099 (I191390,I191382,I191133);
DFFARX1 I_11100 (I191390,I2683,I190949,I190917,);
DFFARX1 I_11101 (I191382,I2683,I190949,I190941,);
not I_11102 (I191435,I191382);
nor I_11103 (I191452,I191435,I191009);
nor I_11104 (I191469,I191274,I191452);
DFFARX1 I_11105 (I191469,I2683,I190949,I190938,);
not I_11106 (I191527,I2690);
DFFARX1 I_11107 (I118469,I2683,I191527,I191553,);
not I_11108 (I191561,I191553);
DFFARX1 I_11109 (I118484,I2683,I191527,I191587,);
not I_11110 (I191595,I118487);
nand I_11111 (I191612,I191595,I118466);
not I_11112 (I191629,I191612);
nor I_11113 (I191646,I191629,I118490);
nor I_11114 (I191663,I191561,I191646);
DFFARX1 I_11115 (I191663,I2683,I191527,I191513,);
not I_11116 (I191694,I118490);
nand I_11117 (I191711,I191694,I191629);
and I_11118 (I191728,I191694,I118472);
nand I_11119 (I191745,I191728,I118463);
nor I_11120 (I191510,I191745,I191694);
and I_11121 (I191501,I191587,I191745);
not I_11122 (I191790,I191745);
nand I_11123 (I191504,I191587,I191790);
nor I_11124 (I191498,I191553,I191745);
not I_11125 (I191835,I118463);
nor I_11126 (I191852,I191835,I118472);
nand I_11127 (I191869,I191852,I191694);
nor I_11128 (I191507,I191612,I191869);
nor I_11129 (I191900,I191835,I118478);
and I_11130 (I191917,I191900,I118481);
or I_11131 (I191934,I191917,I118475);
DFFARX1 I_11132 (I191934,I2683,I191527,I191960,);
nor I_11133 (I191968,I191960,I191711);
DFFARX1 I_11134 (I191968,I2683,I191527,I191495,);
DFFARX1 I_11135 (I191960,I2683,I191527,I191519,);
not I_11136 (I192013,I191960);
nor I_11137 (I192030,I192013,I191587);
nor I_11138 (I192047,I191852,I192030);
DFFARX1 I_11139 (I192047,I2683,I191527,I191516,);
not I_11140 (I192105,I2690);
DFFARX1 I_11141 (I335417,I2683,I192105,I192131,);
not I_11142 (I192139,I192131);
DFFARX1 I_11143 (I335423,I2683,I192105,I192165,);
not I_11144 (I192173,I335417);
nand I_11145 (I192190,I192173,I335420);
not I_11146 (I192207,I192190);
nor I_11147 (I192224,I192207,I335438);
nor I_11148 (I192241,I192139,I192224);
DFFARX1 I_11149 (I192241,I2683,I192105,I192091,);
not I_11150 (I192272,I335438);
nand I_11151 (I192289,I192272,I192207);
and I_11152 (I192306,I192272,I335441);
nand I_11153 (I192323,I192306,I335420);
nor I_11154 (I192088,I192323,I192272);
and I_11155 (I192079,I192165,I192323);
not I_11156 (I192368,I192323);
nand I_11157 (I192082,I192165,I192368);
nor I_11158 (I192076,I192131,I192323);
not I_11159 (I192413,I335426);
nor I_11160 (I192430,I192413,I335441);
nand I_11161 (I192447,I192430,I192272);
nor I_11162 (I192085,I192190,I192447);
nor I_11163 (I192478,I192413,I335432);
and I_11164 (I192495,I192478,I335429);
or I_11165 (I192512,I192495,I335435);
DFFARX1 I_11166 (I192512,I2683,I192105,I192538,);
nor I_11167 (I192546,I192538,I192289);
DFFARX1 I_11168 (I192546,I2683,I192105,I192073,);
DFFARX1 I_11169 (I192538,I2683,I192105,I192097,);
not I_11170 (I192591,I192538);
nor I_11171 (I192608,I192591,I192165);
nor I_11172 (I192625,I192430,I192608);
DFFARX1 I_11173 (I192625,I2683,I192105,I192094,);
not I_11174 (I192683,I2690);
DFFARX1 I_11175 (I325591,I2683,I192683,I192709,);
not I_11176 (I192717,I192709);
DFFARX1 I_11177 (I325597,I2683,I192683,I192743,);
not I_11178 (I192751,I325591);
nand I_11179 (I192768,I192751,I325594);
not I_11180 (I192785,I192768);
nor I_11181 (I192802,I192785,I325612);
nor I_11182 (I192819,I192717,I192802);
DFFARX1 I_11183 (I192819,I2683,I192683,I192669,);
not I_11184 (I192850,I325612);
nand I_11185 (I192867,I192850,I192785);
and I_11186 (I192884,I192850,I325615);
nand I_11187 (I192901,I192884,I325594);
nor I_11188 (I192666,I192901,I192850);
and I_11189 (I192657,I192743,I192901);
not I_11190 (I192946,I192901);
nand I_11191 (I192660,I192743,I192946);
nor I_11192 (I192654,I192709,I192901);
not I_11193 (I192991,I325600);
nor I_11194 (I193008,I192991,I325615);
nand I_11195 (I193025,I193008,I192850);
nor I_11196 (I192663,I192768,I193025);
nor I_11197 (I193056,I192991,I325606);
and I_11198 (I193073,I193056,I325603);
or I_11199 (I193090,I193073,I325609);
DFFARX1 I_11200 (I193090,I2683,I192683,I193116,);
nor I_11201 (I193124,I193116,I192867);
DFFARX1 I_11202 (I193124,I2683,I192683,I192651,);
DFFARX1 I_11203 (I193116,I2683,I192683,I192675,);
not I_11204 (I193169,I193116);
nor I_11205 (I193186,I193169,I192743);
nor I_11206 (I193203,I193008,I193186);
DFFARX1 I_11207 (I193203,I2683,I192683,I192672,);
not I_11208 (I193261,I2690);
DFFARX1 I_11209 (I9360,I2683,I193261,I193287,);
not I_11210 (I193295,I193287);
DFFARX1 I_11211 (I9363,I2683,I193261,I193321,);
not I_11212 (I193329,I9357);
nand I_11213 (I193346,I193329,I9381);
not I_11214 (I193363,I193346);
nor I_11215 (I193380,I193363,I9360);
nor I_11216 (I193397,I193295,I193380);
DFFARX1 I_11217 (I193397,I2683,I193261,I193247,);
not I_11218 (I193428,I9360);
nand I_11219 (I193445,I193428,I193363);
and I_11220 (I193462,I193428,I9375);
nand I_11221 (I193479,I193462,I9369);
nor I_11222 (I193244,I193479,I193428);
and I_11223 (I193235,I193321,I193479);
not I_11224 (I193524,I193479);
nand I_11225 (I193238,I193321,I193524);
nor I_11226 (I193232,I193287,I193479);
not I_11227 (I193569,I9378);
nor I_11228 (I193586,I193569,I9375);
nand I_11229 (I193603,I193586,I193428);
nor I_11230 (I193241,I193346,I193603);
nor I_11231 (I193634,I193569,I9357);
and I_11232 (I193651,I193634,I9366);
or I_11233 (I193668,I193651,I9372);
DFFARX1 I_11234 (I193668,I2683,I193261,I193694,);
nor I_11235 (I193702,I193694,I193445);
DFFARX1 I_11236 (I193702,I2683,I193261,I193229,);
DFFARX1 I_11237 (I193694,I2683,I193261,I193253,);
not I_11238 (I193747,I193694);
nor I_11239 (I193764,I193747,I193321);
nor I_11240 (I193781,I193586,I193764);
DFFARX1 I_11241 (I193781,I2683,I193261,I193250,);
not I_11242 (I193839,I2690);
DFFARX1 I_11243 (I363757,I2683,I193839,I193865,);
not I_11244 (I193873,I193865);
nand I_11245 (I193890,I363739,I363751);
and I_11246 (I193907,I193890,I363754);
DFFARX1 I_11247 (I193907,I2683,I193839,I193933,);
not I_11248 (I193941,I363748);
DFFARX1 I_11249 (I363745,I2683,I193839,I193967,);
not I_11250 (I193975,I193967);
nor I_11251 (I193992,I193975,I193873);
and I_11252 (I194009,I193992,I363748);
nor I_11253 (I194026,I193975,I193941);
nor I_11254 (I193822,I193933,I194026);
DFFARX1 I_11255 (I363763,I2683,I193839,I194066,);
nor I_11256 (I194074,I194066,I193933);
not I_11257 (I194091,I194074);
not I_11258 (I194108,I194066);
nor I_11259 (I194125,I194108,I194009);
DFFARX1 I_11260 (I194125,I2683,I193839,I193825,);
nand I_11261 (I194156,I363742,I363742);
and I_11262 (I194173,I194156,I363739);
DFFARX1 I_11263 (I194173,I2683,I193839,I194199,);
nor I_11264 (I194207,I194199,I194066);
DFFARX1 I_11265 (I194207,I2683,I193839,I193807,);
nand I_11266 (I194238,I194199,I194108);
nand I_11267 (I193816,I194091,I194238);
not I_11268 (I194269,I194199);
nor I_11269 (I194286,I194269,I194009);
DFFARX1 I_11270 (I194286,I2683,I193839,I193828,);
nor I_11271 (I194317,I363760,I363742);
or I_11272 (I193819,I194066,I194317);
nor I_11273 (I193810,I194199,I194317);
or I_11274 (I193813,I193933,I194317);
DFFARX1 I_11275 (I194317,I2683,I193839,I193831,);
not I_11276 (I194417,I2690);
DFFARX1 I_11277 (I2612,I2683,I194417,I194443,);
not I_11278 (I194451,I194443);
nand I_11279 (I194468,I2388,I2132);
and I_11280 (I194485,I194468,I2500);
DFFARX1 I_11281 (I194485,I2683,I194417,I194511,);
not I_11282 (I194519,I1500);
DFFARX1 I_11283 (I2516,I2683,I194417,I194545,);
not I_11284 (I194553,I194545);
nor I_11285 (I194570,I194553,I194451);
and I_11286 (I194587,I194570,I1500);
nor I_11287 (I194604,I194553,I194519);
nor I_11288 (I194400,I194511,I194604);
DFFARX1 I_11289 (I1772,I2683,I194417,I194644,);
nor I_11290 (I194652,I194644,I194511);
not I_11291 (I194669,I194652);
not I_11292 (I194686,I194644);
nor I_11293 (I194703,I194686,I194587);
DFFARX1 I_11294 (I194703,I2683,I194417,I194403,);
nand I_11295 (I194734,I1948,I1436);
and I_11296 (I194751,I194734,I1660);
DFFARX1 I_11297 (I194751,I2683,I194417,I194777,);
nor I_11298 (I194785,I194777,I194644);
DFFARX1 I_11299 (I194785,I2683,I194417,I194385,);
nand I_11300 (I194816,I194777,I194686);
nand I_11301 (I194394,I194669,I194816);
not I_11302 (I194847,I194777);
nor I_11303 (I194864,I194847,I194587);
DFFARX1 I_11304 (I194864,I2683,I194417,I194406,);
nor I_11305 (I194895,I1812,I1436);
or I_11306 (I194397,I194644,I194895);
nor I_11307 (I194388,I194777,I194895);
or I_11308 (I194391,I194511,I194895);
DFFARX1 I_11309 (I194895,I2683,I194417,I194409,);
not I_11310 (I194995,I2690);
DFFARX1 I_11311 (I37818,I2683,I194995,I195021,);
not I_11312 (I195029,I195021);
nand I_11313 (I195046,I37827,I37836);
and I_11314 (I195063,I195046,I37815);
DFFARX1 I_11315 (I195063,I2683,I194995,I195089,);
not I_11316 (I195097,I37818);
DFFARX1 I_11317 (I37833,I2683,I194995,I195123,);
not I_11318 (I195131,I195123);
nor I_11319 (I195148,I195131,I195029);
and I_11320 (I195165,I195148,I37818);
nor I_11321 (I195182,I195131,I195097);
nor I_11322 (I194978,I195089,I195182);
DFFARX1 I_11323 (I37824,I2683,I194995,I195222,);
nor I_11324 (I195230,I195222,I195089);
not I_11325 (I195247,I195230);
not I_11326 (I195264,I195222);
nor I_11327 (I195281,I195264,I195165);
DFFARX1 I_11328 (I195281,I2683,I194995,I194981,);
nand I_11329 (I195312,I37839,I37815);
and I_11330 (I195329,I195312,I37821);
DFFARX1 I_11331 (I195329,I2683,I194995,I195355,);
nor I_11332 (I195363,I195355,I195222);
DFFARX1 I_11333 (I195363,I2683,I194995,I194963,);
nand I_11334 (I195394,I195355,I195264);
nand I_11335 (I194972,I195247,I195394);
not I_11336 (I195425,I195355);
nor I_11337 (I195442,I195425,I195165);
DFFARX1 I_11338 (I195442,I2683,I194995,I194984,);
nor I_11339 (I195473,I37830,I37815);
or I_11340 (I194975,I195222,I195473);
nor I_11341 (I194966,I195355,I195473);
or I_11342 (I194969,I195089,I195473);
DFFARX1 I_11343 (I195473,I2683,I194995,I194987,);
not I_11344 (I195573,I2690);
DFFARX1 I_11345 (I117433,I2683,I195573,I195599,);
not I_11346 (I195607,I195599);
nand I_11347 (I195624,I117436,I117412);
and I_11348 (I195641,I195624,I117409);
DFFARX1 I_11349 (I195641,I2683,I195573,I195667,);
not I_11350 (I195675,I117415);
DFFARX1 I_11351 (I117409,I2683,I195573,I195701,);
not I_11352 (I195709,I195701);
nor I_11353 (I195726,I195709,I195607);
and I_11354 (I195743,I195726,I117415);
nor I_11355 (I195760,I195709,I195675);
nor I_11356 (I195556,I195667,I195760);
DFFARX1 I_11357 (I117418,I2683,I195573,I195800,);
nor I_11358 (I195808,I195800,I195667);
not I_11359 (I195825,I195808);
not I_11360 (I195842,I195800);
nor I_11361 (I195859,I195842,I195743);
DFFARX1 I_11362 (I195859,I2683,I195573,I195559,);
nand I_11363 (I195890,I117421,I117430);
and I_11364 (I195907,I195890,I117427);
DFFARX1 I_11365 (I195907,I2683,I195573,I195933,);
nor I_11366 (I195941,I195933,I195800);
DFFARX1 I_11367 (I195941,I2683,I195573,I195541,);
nand I_11368 (I195972,I195933,I195842);
nand I_11369 (I195550,I195825,I195972);
not I_11370 (I196003,I195933);
nor I_11371 (I196020,I196003,I195743);
DFFARX1 I_11372 (I196020,I2683,I195573,I195562,);
nor I_11373 (I196051,I117424,I117430);
or I_11374 (I195553,I195800,I196051);
nor I_11375 (I195544,I195933,I196051);
or I_11376 (I195547,I195667,I196051);
DFFARX1 I_11377 (I196051,I2683,I195573,I195565,);
not I_11378 (I196151,I2690);
DFFARX1 I_11379 (I8315,I2683,I196151,I196177,);
not I_11380 (I196185,I196177);
nand I_11381 (I196202,I8312,I8303);
and I_11382 (I196219,I196202,I8303);
DFFARX1 I_11383 (I196219,I2683,I196151,I196245,);
not I_11384 (I196253,I8306);
DFFARX1 I_11385 (I8321,I2683,I196151,I196279,);
not I_11386 (I196287,I196279);
nor I_11387 (I196304,I196287,I196185);
and I_11388 (I196321,I196304,I8306);
nor I_11389 (I196338,I196287,I196253);
nor I_11390 (I196134,I196245,I196338);
DFFARX1 I_11391 (I8306,I2683,I196151,I196378,);
nor I_11392 (I196386,I196378,I196245);
not I_11393 (I196403,I196386);
not I_11394 (I196420,I196378);
nor I_11395 (I196437,I196420,I196321);
DFFARX1 I_11396 (I196437,I2683,I196151,I196137,);
nand I_11397 (I196468,I8324,I8309);
and I_11398 (I196485,I196468,I8327);
DFFARX1 I_11399 (I196485,I2683,I196151,I196511,);
nor I_11400 (I196519,I196511,I196378);
DFFARX1 I_11401 (I196519,I2683,I196151,I196119,);
nand I_11402 (I196550,I196511,I196420);
nand I_11403 (I196128,I196403,I196550);
not I_11404 (I196581,I196511);
nor I_11405 (I196598,I196581,I196321);
DFFARX1 I_11406 (I196598,I2683,I196151,I196140,);
nor I_11407 (I196629,I8318,I8309);
or I_11408 (I196131,I196378,I196629);
nor I_11409 (I196122,I196511,I196629);
or I_11410 (I196125,I196245,I196629);
DFFARX1 I_11411 (I196629,I2683,I196151,I196143,);
not I_11412 (I196729,I2690);
DFFARX1 I_11413 (I273034,I2683,I196729,I196755,);
not I_11414 (I196763,I196755);
nand I_11415 (I196780,I273010,I273025);
and I_11416 (I196797,I196780,I273037);
DFFARX1 I_11417 (I196797,I2683,I196729,I196823,);
not I_11418 (I196831,I273022);
DFFARX1 I_11419 (I273013,I2683,I196729,I196857,);
not I_11420 (I196865,I196857);
nor I_11421 (I196882,I196865,I196763);
and I_11422 (I196899,I196882,I273022);
nor I_11423 (I196916,I196865,I196831);
nor I_11424 (I196712,I196823,I196916);
DFFARX1 I_11425 (I273010,I2683,I196729,I196956,);
nor I_11426 (I196964,I196956,I196823);
not I_11427 (I196981,I196964);
not I_11428 (I196998,I196956);
nor I_11429 (I197015,I196998,I196899);
DFFARX1 I_11430 (I197015,I2683,I196729,I196715,);
nand I_11431 (I197046,I273028,I273019);
and I_11432 (I197063,I197046,I273031);
DFFARX1 I_11433 (I197063,I2683,I196729,I197089,);
nor I_11434 (I197097,I197089,I196956);
DFFARX1 I_11435 (I197097,I2683,I196729,I196697,);
nand I_11436 (I197128,I197089,I196998);
nand I_11437 (I196706,I196981,I197128);
not I_11438 (I197159,I197089);
nor I_11439 (I197176,I197159,I196899);
DFFARX1 I_11440 (I197176,I2683,I196729,I196718,);
nor I_11441 (I197207,I273016,I273019);
or I_11442 (I196709,I196956,I197207);
nor I_11443 (I196700,I197089,I197207);
or I_11444 (I196703,I196823,I197207);
DFFARX1 I_11445 (I197207,I2683,I196729,I196721,);
not I_11446 (I197307,I2690);
DFFARX1 I_11447 (I113744,I2683,I197307,I197333,);
not I_11448 (I197341,I197333);
nand I_11449 (I197358,I113747,I113723);
and I_11450 (I197375,I197358,I113720);
DFFARX1 I_11451 (I197375,I2683,I197307,I197401,);
not I_11452 (I197409,I113726);
DFFARX1 I_11453 (I113720,I2683,I197307,I197435,);
not I_11454 (I197443,I197435);
nor I_11455 (I197460,I197443,I197341);
and I_11456 (I197477,I197460,I113726);
nor I_11457 (I197494,I197443,I197409);
nor I_11458 (I197290,I197401,I197494);
DFFARX1 I_11459 (I113729,I2683,I197307,I197534,);
nor I_11460 (I197542,I197534,I197401);
not I_11461 (I197559,I197542);
not I_11462 (I197576,I197534);
nor I_11463 (I197593,I197576,I197477);
DFFARX1 I_11464 (I197593,I2683,I197307,I197293,);
nand I_11465 (I197624,I113732,I113741);
and I_11466 (I197641,I197624,I113738);
DFFARX1 I_11467 (I197641,I2683,I197307,I197667,);
nor I_11468 (I197675,I197667,I197534);
DFFARX1 I_11469 (I197675,I2683,I197307,I197275,);
nand I_11470 (I197706,I197667,I197576);
nand I_11471 (I197284,I197559,I197706);
not I_11472 (I197737,I197667);
nor I_11473 (I197754,I197737,I197477);
DFFARX1 I_11474 (I197754,I2683,I197307,I197296,);
nor I_11475 (I197785,I113735,I113741);
or I_11476 (I197287,I197534,I197785);
nor I_11477 (I197278,I197667,I197785);
or I_11478 (I197281,I197401,I197785);
DFFARX1 I_11479 (I197785,I2683,I197307,I197299,);
not I_11480 (I197885,I2690);
DFFARX1 I_11481 (I145400,I2683,I197885,I197911,);
not I_11482 (I197919,I197911);
nand I_11483 (I197936,I145391,I145409);
and I_11484 (I197953,I197936,I145412);
DFFARX1 I_11485 (I197953,I2683,I197885,I197979,);
not I_11486 (I197987,I145406);
DFFARX1 I_11487 (I145394,I2683,I197885,I198013,);
not I_11488 (I198021,I198013);
nor I_11489 (I198038,I198021,I197919);
and I_11490 (I198055,I198038,I145406);
nor I_11491 (I198072,I198021,I197987);
nor I_11492 (I197868,I197979,I198072);
DFFARX1 I_11493 (I145403,I2683,I197885,I198112,);
nor I_11494 (I198120,I198112,I197979);
not I_11495 (I198137,I198120);
not I_11496 (I198154,I198112);
nor I_11497 (I198171,I198154,I198055);
DFFARX1 I_11498 (I198171,I2683,I197885,I197871,);
nand I_11499 (I198202,I145418,I145415);
and I_11500 (I198219,I198202,I145397);
DFFARX1 I_11501 (I198219,I2683,I197885,I198245,);
nor I_11502 (I198253,I198245,I198112);
DFFARX1 I_11503 (I198253,I2683,I197885,I197853,);
nand I_11504 (I198284,I198245,I198154);
nand I_11505 (I197862,I198137,I198284);
not I_11506 (I198315,I198245);
nor I_11507 (I198332,I198315,I198055);
DFFARX1 I_11508 (I198332,I2683,I197885,I197874,);
nor I_11509 (I198363,I145391,I145415);
or I_11510 (I197865,I198112,I198363);
nor I_11511 (I197856,I198245,I198363);
or I_11512 (I197859,I197979,I198363);
DFFARX1 I_11513 (I198363,I2683,I197885,I197877,);
not I_11514 (I198463,I2690);
DFFARX1 I_11515 (I360289,I2683,I198463,I198489,);
not I_11516 (I198497,I198489);
nand I_11517 (I198514,I360271,I360283);
and I_11518 (I198531,I198514,I360286);
DFFARX1 I_11519 (I198531,I2683,I198463,I198557,);
not I_11520 (I198565,I360280);
DFFARX1 I_11521 (I360277,I2683,I198463,I198591,);
not I_11522 (I198599,I198591);
nor I_11523 (I198616,I198599,I198497);
and I_11524 (I198633,I198616,I360280);
nor I_11525 (I198650,I198599,I198565);
nor I_11526 (I198446,I198557,I198650);
DFFARX1 I_11527 (I360295,I2683,I198463,I198690,);
nor I_11528 (I198698,I198690,I198557);
not I_11529 (I198715,I198698);
not I_11530 (I198732,I198690);
nor I_11531 (I198749,I198732,I198633);
DFFARX1 I_11532 (I198749,I2683,I198463,I198449,);
nand I_11533 (I198780,I360274,I360274);
and I_11534 (I198797,I198780,I360271);
DFFARX1 I_11535 (I198797,I2683,I198463,I198823,);
nor I_11536 (I198831,I198823,I198690);
DFFARX1 I_11537 (I198831,I2683,I198463,I198431,);
nand I_11538 (I198862,I198823,I198732);
nand I_11539 (I198440,I198715,I198862);
not I_11540 (I198893,I198823);
nor I_11541 (I198910,I198893,I198633);
DFFARX1 I_11542 (I198910,I2683,I198463,I198452,);
nor I_11543 (I198941,I360292,I360274);
or I_11544 (I198443,I198690,I198941);
nor I_11545 (I198434,I198823,I198941);
or I_11546 (I198437,I198557,I198941);
DFFARX1 I_11547 (I198941,I2683,I198463,I198455,);
not I_11548 (I199041,I2690);
DFFARX1 I_11549 (I166539,I2683,I199041,I199067,);
not I_11550 (I199075,I199067);
nand I_11551 (I199092,I166554,I166539);
and I_11552 (I199109,I199092,I166542);
DFFARX1 I_11553 (I199109,I2683,I199041,I199135,);
not I_11554 (I199143,I166542);
DFFARX1 I_11555 (I166551,I2683,I199041,I199169,);
not I_11556 (I199177,I199169);
nor I_11557 (I199194,I199177,I199075);
and I_11558 (I199211,I199194,I166542);
nor I_11559 (I199228,I199177,I199143);
nor I_11560 (I199024,I199135,I199228);
DFFARX1 I_11561 (I166545,I2683,I199041,I199268,);
nor I_11562 (I199276,I199268,I199135);
not I_11563 (I199293,I199276);
not I_11564 (I199310,I199268);
nor I_11565 (I199327,I199310,I199211);
DFFARX1 I_11566 (I199327,I2683,I199041,I199027,);
nand I_11567 (I199358,I166548,I166557);
and I_11568 (I199375,I199358,I166563);
DFFARX1 I_11569 (I199375,I2683,I199041,I199401,);
nor I_11570 (I199409,I199401,I199268);
DFFARX1 I_11571 (I199409,I2683,I199041,I199009,);
nand I_11572 (I199440,I199401,I199310);
nand I_11573 (I199018,I199293,I199440);
not I_11574 (I199471,I199401);
nor I_11575 (I199488,I199471,I199211);
DFFARX1 I_11576 (I199488,I2683,I199041,I199030,);
nor I_11577 (I199519,I166560,I166557);
or I_11578 (I199021,I199268,I199519);
nor I_11579 (I199012,I199401,I199519);
or I_11580 (I199015,I199135,I199519);
DFFARX1 I_11581 (I199519,I2683,I199041,I199033,);
not I_11582 (I199619,I2690);
DFFARX1 I_11583 (I370845,I2683,I199619,I199645,);
not I_11584 (I199653,I199645);
nand I_11585 (I199670,I370848,I370857);
and I_11586 (I199687,I199670,I370860);
DFFARX1 I_11587 (I199687,I2683,I199619,I199713,);
not I_11588 (I199721,I370869);
DFFARX1 I_11589 (I370851,I2683,I199619,I199747,);
not I_11590 (I199755,I199747);
nor I_11591 (I199772,I199755,I199653);
and I_11592 (I199789,I199772,I370869);
nor I_11593 (I199806,I199755,I199721);
nor I_11594 (I199602,I199713,I199806);
DFFARX1 I_11595 (I370848,I2683,I199619,I199846,);
nor I_11596 (I199854,I199846,I199713);
not I_11597 (I199871,I199854);
not I_11598 (I199888,I199846);
nor I_11599 (I199905,I199888,I199789);
DFFARX1 I_11600 (I199905,I2683,I199619,I199605,);
nand I_11601 (I199936,I370866,I370845);
and I_11602 (I199953,I199936,I370863);
DFFARX1 I_11603 (I199953,I2683,I199619,I199979,);
nor I_11604 (I199987,I199979,I199846);
DFFARX1 I_11605 (I199987,I2683,I199619,I199587,);
nand I_11606 (I200018,I199979,I199888);
nand I_11607 (I199596,I199871,I200018);
not I_11608 (I200049,I199979);
nor I_11609 (I200066,I200049,I199789);
DFFARX1 I_11610 (I200066,I2683,I199619,I199608,);
nor I_11611 (I200097,I370854,I370845);
or I_11612 (I199599,I199846,I200097);
nor I_11613 (I199590,I199979,I200097);
or I_11614 (I199593,I199713,I200097);
DFFARX1 I_11615 (I200097,I2683,I199619,I199611,);
not I_11616 (I200197,I2690);
DFFARX1 I_11617 (I2492,I2683,I200197,I200223,);
not I_11618 (I200231,I200223);
nand I_11619 (I200248,I1548,I2332);
and I_11620 (I200265,I200248,I1892);
DFFARX1 I_11621 (I200265,I2683,I200197,I200291,);
not I_11622 (I200299,I1852);
DFFARX1 I_11623 (I2188,I2683,I200197,I200325,);
not I_11624 (I200333,I200325);
nor I_11625 (I200350,I200333,I200231);
and I_11626 (I200367,I200350,I1852);
nor I_11627 (I200384,I200333,I200299);
nor I_11628 (I200180,I200291,I200384);
DFFARX1 I_11629 (I2676,I2683,I200197,I200424,);
nor I_11630 (I200432,I200424,I200291);
not I_11631 (I200449,I200432);
not I_11632 (I200466,I200424);
nor I_11633 (I200483,I200466,I200367);
DFFARX1 I_11634 (I200483,I2683,I200197,I200183,);
nand I_11635 (I200514,I2164,I1732);
and I_11636 (I200531,I200514,I2004);
DFFARX1 I_11637 (I200531,I2683,I200197,I200557,);
nor I_11638 (I200565,I200557,I200424);
DFFARX1 I_11639 (I200565,I2683,I200197,I200165,);
nand I_11640 (I200596,I200557,I200466);
nand I_11641 (I200174,I200449,I200596);
not I_11642 (I200627,I200557);
nor I_11643 (I200644,I200627,I200367);
DFFARX1 I_11644 (I200644,I2683,I200197,I200186,);
nor I_11645 (I200675,I2172,I1732);
or I_11646 (I200177,I200424,I200675);
nor I_11647 (I200168,I200557,I200675);
or I_11648 (I200171,I200291,I200675);
DFFARX1 I_11649 (I200675,I2683,I200197,I200189,);
not I_11650 (I200775,I2690);
DFFARX1 I_11651 (I308564,I2683,I200775,I200801,);
not I_11652 (I200809,I200801);
nand I_11653 (I200826,I308540,I308555);
and I_11654 (I200843,I200826,I308567);
DFFARX1 I_11655 (I200843,I2683,I200775,I200869,);
not I_11656 (I200877,I308552);
DFFARX1 I_11657 (I308543,I2683,I200775,I200903,);
not I_11658 (I200911,I200903);
nor I_11659 (I200928,I200911,I200809);
and I_11660 (I200945,I200928,I308552);
nor I_11661 (I200962,I200911,I200877);
nor I_11662 (I200758,I200869,I200962);
DFFARX1 I_11663 (I308540,I2683,I200775,I201002,);
nor I_11664 (I201010,I201002,I200869);
not I_11665 (I201027,I201010);
not I_11666 (I201044,I201002);
nor I_11667 (I201061,I201044,I200945);
DFFARX1 I_11668 (I201061,I2683,I200775,I200761,);
nand I_11669 (I201092,I308558,I308549);
and I_11670 (I201109,I201092,I308561);
DFFARX1 I_11671 (I201109,I2683,I200775,I201135,);
nor I_11672 (I201143,I201135,I201002);
DFFARX1 I_11673 (I201143,I2683,I200775,I200743,);
nand I_11674 (I201174,I201135,I201044);
nand I_11675 (I200752,I201027,I201174);
not I_11676 (I201205,I201135);
nor I_11677 (I201222,I201205,I200945);
DFFARX1 I_11678 (I201222,I2683,I200775,I200764,);
nor I_11679 (I201253,I308546,I308549);
or I_11680 (I200755,I201002,I201253);
nor I_11681 (I200746,I201135,I201253);
or I_11682 (I200749,I200869,I201253);
DFFARX1 I_11683 (I201253,I2683,I200775,I200767,);
not I_11684 (I201353,I2690);
DFFARX1 I_11685 (I103731,I2683,I201353,I201379,);
not I_11686 (I201387,I201379);
nand I_11687 (I201404,I103734,I103710);
and I_11688 (I201421,I201404,I103707);
DFFARX1 I_11689 (I201421,I2683,I201353,I201447,);
not I_11690 (I201455,I103713);
DFFARX1 I_11691 (I103707,I2683,I201353,I201481,);
not I_11692 (I201489,I201481);
nor I_11693 (I201506,I201489,I201387);
and I_11694 (I201523,I201506,I103713);
nor I_11695 (I201540,I201489,I201455);
nor I_11696 (I201336,I201447,I201540);
DFFARX1 I_11697 (I103716,I2683,I201353,I201580,);
nor I_11698 (I201588,I201580,I201447);
not I_11699 (I201605,I201588);
not I_11700 (I201622,I201580);
nor I_11701 (I201639,I201622,I201523);
DFFARX1 I_11702 (I201639,I2683,I201353,I201339,);
nand I_11703 (I201670,I103719,I103728);
and I_11704 (I201687,I201670,I103725);
DFFARX1 I_11705 (I201687,I2683,I201353,I201713,);
nor I_11706 (I201721,I201713,I201580);
DFFARX1 I_11707 (I201721,I2683,I201353,I201321,);
nand I_11708 (I201752,I201713,I201622);
nand I_11709 (I201330,I201605,I201752);
not I_11710 (I201783,I201713);
nor I_11711 (I201800,I201783,I201523);
DFFARX1 I_11712 (I201800,I2683,I201353,I201342,);
nor I_11713 (I201831,I103722,I103728);
or I_11714 (I201333,I201580,I201831);
nor I_11715 (I201324,I201713,I201831);
or I_11716 (I201327,I201447,I201831);
DFFARX1 I_11717 (I201831,I2683,I201353,I201345,);
not I_11718 (I201931,I2690);
DFFARX1 I_11719 (I179357,I2683,I201931,I201957,);
not I_11720 (I201965,I201957);
nand I_11721 (I201982,I179366,I179375);
and I_11722 (I201999,I201982,I179381);
DFFARX1 I_11723 (I201999,I2683,I201931,I202025,);
not I_11724 (I202033,I179378);
DFFARX1 I_11725 (I179363,I2683,I201931,I202059,);
not I_11726 (I202067,I202059);
nor I_11727 (I202084,I202067,I201965);
and I_11728 (I202101,I202084,I179378);
nor I_11729 (I202118,I202067,I202033);
nor I_11730 (I201914,I202025,I202118);
DFFARX1 I_11731 (I179372,I2683,I201931,I202158,);
nor I_11732 (I202166,I202158,I202025);
not I_11733 (I202183,I202166);
not I_11734 (I202200,I202158);
nor I_11735 (I202217,I202200,I202101);
DFFARX1 I_11736 (I202217,I2683,I201931,I201917,);
nand I_11737 (I202248,I179369,I179360);
and I_11738 (I202265,I202248,I179357);
DFFARX1 I_11739 (I202265,I2683,I201931,I202291,);
nor I_11740 (I202299,I202291,I202158);
DFFARX1 I_11741 (I202299,I2683,I201931,I201899,);
nand I_11742 (I202330,I202291,I202200);
nand I_11743 (I201908,I202183,I202330);
not I_11744 (I202361,I202291);
nor I_11745 (I202378,I202361,I202101);
DFFARX1 I_11746 (I202378,I2683,I201931,I201920,);
nor I_11747 (I202409,I179360,I179360);
or I_11748 (I201911,I202158,I202409);
nor I_11749 (I201902,I202291,I202409);
or I_11750 (I201905,I202025,I202409);
DFFARX1 I_11751 (I202409,I2683,I201931,I201923,);
not I_11752 (I202509,I2690);
DFFARX1 I_11753 (I381895,I2683,I202509,I202535,);
not I_11754 (I202543,I202535);
nand I_11755 (I202560,I381919,I381901);
and I_11756 (I202577,I202560,I381907);
DFFARX1 I_11757 (I202577,I2683,I202509,I202603,);
not I_11758 (I202611,I381913);
DFFARX1 I_11759 (I381898,I2683,I202509,I202637,);
not I_11760 (I202645,I202637);
nor I_11761 (I202662,I202645,I202543);
and I_11762 (I202679,I202662,I381913);
nor I_11763 (I202696,I202645,I202611);
nor I_11764 (I202492,I202603,I202696);
DFFARX1 I_11765 (I381910,I2683,I202509,I202736,);
nor I_11766 (I202744,I202736,I202603);
not I_11767 (I202761,I202744);
not I_11768 (I202778,I202736);
nor I_11769 (I202795,I202778,I202679);
DFFARX1 I_11770 (I202795,I2683,I202509,I202495,);
nand I_11771 (I202826,I381916,I381904);
and I_11772 (I202843,I202826,I381898);
DFFARX1 I_11773 (I202843,I2683,I202509,I202869,);
nor I_11774 (I202877,I202869,I202736);
DFFARX1 I_11775 (I202877,I2683,I202509,I202477,);
nand I_11776 (I202908,I202869,I202778);
nand I_11777 (I202486,I202761,I202908);
not I_11778 (I202939,I202869);
nor I_11779 (I202956,I202939,I202679);
DFFARX1 I_11780 (I202956,I2683,I202509,I202498,);
nor I_11781 (I202987,I381895,I381904);
or I_11782 (I202489,I202736,I202987);
nor I_11783 (I202480,I202869,I202987);
or I_11784 (I202483,I202603,I202987);
DFFARX1 I_11785 (I202987,I2683,I202509,I202501,);
not I_11786 (I203087,I2690);
DFFARX1 I_11787 (I409326,I2683,I203087,I203113,);
not I_11788 (I203121,I203113);
nand I_11789 (I203138,I409311,I409299);
and I_11790 (I203155,I203138,I409314);
DFFARX1 I_11791 (I203155,I2683,I203087,I203181,);
not I_11792 (I203189,I409299);
DFFARX1 I_11793 (I409317,I2683,I203087,I203215,);
not I_11794 (I203223,I203215);
nor I_11795 (I203240,I203223,I203121);
and I_11796 (I203257,I203240,I409299);
nor I_11797 (I203274,I203223,I203189);
nor I_11798 (I203070,I203181,I203274);
DFFARX1 I_11799 (I409305,I2683,I203087,I203314,);
nor I_11800 (I203322,I203314,I203181);
not I_11801 (I203339,I203322);
not I_11802 (I203356,I203314);
nor I_11803 (I203373,I203356,I203257);
DFFARX1 I_11804 (I203373,I2683,I203087,I203073,);
nand I_11805 (I203404,I409302,I409308);
and I_11806 (I203421,I203404,I409323);
DFFARX1 I_11807 (I203421,I2683,I203087,I203447,);
nor I_11808 (I203455,I203447,I203314);
DFFARX1 I_11809 (I203455,I2683,I203087,I203055,);
nand I_11810 (I203486,I203447,I203356);
nand I_11811 (I203064,I203339,I203486);
not I_11812 (I203517,I203447);
nor I_11813 (I203534,I203517,I203257);
DFFARX1 I_11814 (I203534,I2683,I203087,I203076,);
nor I_11815 (I203565,I409320,I409308);
or I_11816 (I203067,I203314,I203565);
nor I_11817 (I203058,I203447,I203565);
or I_11818 (I203061,I203181,I203565);
DFFARX1 I_11819 (I203565,I2683,I203087,I203079,);
not I_11820 (I203665,I2690);
DFFARX1 I_11821 (I2508,I2683,I203665,I203691,);
not I_11822 (I203699,I203691);
nand I_11823 (I203716,I2204,I1716);
and I_11824 (I203733,I203716,I2436);
DFFARX1 I_11825 (I203733,I2683,I203665,I203759,);
not I_11826 (I203767,I2660);
DFFARX1 I_11827 (I1596,I2683,I203665,I203793,);
not I_11828 (I203801,I203793);
nor I_11829 (I203818,I203801,I203699);
and I_11830 (I203835,I203818,I2660);
nor I_11831 (I203852,I203801,I203767);
nor I_11832 (I203648,I203759,I203852);
DFFARX1 I_11833 (I1916,I2683,I203665,I203892,);
nor I_11834 (I203900,I203892,I203759);
not I_11835 (I203917,I203900);
not I_11836 (I203934,I203892);
nor I_11837 (I203951,I203934,I203835);
DFFARX1 I_11838 (I203951,I2683,I203665,I203651,);
nand I_11839 (I203982,I1492,I2196);
and I_11840 (I203999,I203982,I1724);
DFFARX1 I_11841 (I203999,I2683,I203665,I204025,);
nor I_11842 (I204033,I204025,I203892);
DFFARX1 I_11843 (I204033,I2683,I203665,I203633,);
nand I_11844 (I204064,I204025,I203934);
nand I_11845 (I203642,I203917,I204064);
not I_11846 (I204095,I204025);
nor I_11847 (I204112,I204095,I203835);
DFFARX1 I_11848 (I204112,I2683,I203665,I203654,);
nor I_11849 (I204143,I2460,I2196);
or I_11850 (I203645,I203892,I204143);
nor I_11851 (I203636,I204025,I204143);
or I_11852 (I203639,I203759,I204143);
DFFARX1 I_11853 (I204143,I2683,I203665,I203657,);
not I_11854 (I204243,I2690);
DFFARX1 I_11855 (I90556,I2683,I204243,I204269,);
not I_11856 (I204277,I204269);
nand I_11857 (I204294,I90559,I90535);
and I_11858 (I204311,I204294,I90532);
DFFARX1 I_11859 (I204311,I2683,I204243,I204337,);
not I_11860 (I204345,I90538);
DFFARX1 I_11861 (I90532,I2683,I204243,I204371,);
not I_11862 (I204379,I204371);
nor I_11863 (I204396,I204379,I204277);
and I_11864 (I204413,I204396,I90538);
nor I_11865 (I204430,I204379,I204345);
nor I_11866 (I204226,I204337,I204430);
DFFARX1 I_11867 (I90541,I2683,I204243,I204470,);
nor I_11868 (I204478,I204470,I204337);
not I_11869 (I204495,I204478);
not I_11870 (I204512,I204470);
nor I_11871 (I204529,I204512,I204413);
DFFARX1 I_11872 (I204529,I2683,I204243,I204229,);
nand I_11873 (I204560,I90544,I90553);
and I_11874 (I204577,I204560,I90550);
DFFARX1 I_11875 (I204577,I2683,I204243,I204603,);
nor I_11876 (I204611,I204603,I204470);
DFFARX1 I_11877 (I204611,I2683,I204243,I204211,);
nand I_11878 (I204642,I204603,I204512);
nand I_11879 (I204220,I204495,I204642);
not I_11880 (I204673,I204603);
nor I_11881 (I204690,I204673,I204413);
DFFARX1 I_11882 (I204690,I2683,I204243,I204232,);
nor I_11883 (I204721,I90547,I90553);
or I_11884 (I204223,I204470,I204721);
nor I_11885 (I204214,I204603,I204721);
or I_11886 (I204217,I204337,I204721);
DFFARX1 I_11887 (I204721,I2683,I204243,I204235,);
not I_11888 (I204821,I2690);
DFFARX1 I_11889 (I349307,I2683,I204821,I204847,);
not I_11890 (I204855,I204847);
nand I_11891 (I204872,I349289,I349301);
and I_11892 (I204889,I204872,I349304);
DFFARX1 I_11893 (I204889,I2683,I204821,I204915,);
not I_11894 (I204923,I349298);
DFFARX1 I_11895 (I349295,I2683,I204821,I204949,);
not I_11896 (I204957,I204949);
nor I_11897 (I204974,I204957,I204855);
and I_11898 (I204991,I204974,I349298);
nor I_11899 (I205008,I204957,I204923);
nor I_11900 (I204804,I204915,I205008);
DFFARX1 I_11901 (I349313,I2683,I204821,I205048,);
nor I_11902 (I205056,I205048,I204915);
not I_11903 (I205073,I205056);
not I_11904 (I205090,I205048);
nor I_11905 (I205107,I205090,I204991);
DFFARX1 I_11906 (I205107,I2683,I204821,I204807,);
nand I_11907 (I205138,I349292,I349292);
and I_11908 (I205155,I205138,I349289);
DFFARX1 I_11909 (I205155,I2683,I204821,I205181,);
nor I_11910 (I205189,I205181,I205048);
DFFARX1 I_11911 (I205189,I2683,I204821,I204789,);
nand I_11912 (I205220,I205181,I205090);
nand I_11913 (I204798,I205073,I205220);
not I_11914 (I205251,I205181);
nor I_11915 (I205268,I205251,I204991);
DFFARX1 I_11916 (I205268,I2683,I204821,I204810,);
nor I_11917 (I205299,I349310,I349292);
or I_11918 (I204801,I205048,I205299);
nor I_11919 (I204792,I205181,I205299);
or I_11920 (I204795,I204915,I205299);
DFFARX1 I_11921 (I205299,I2683,I204821,I204813,);
not I_11922 (I205399,I2690);
DFFARX1 I_11923 (I10423,I2683,I205399,I205425,);
not I_11924 (I205433,I205425);
nand I_11925 (I205450,I10420,I10411);
and I_11926 (I205467,I205450,I10411);
DFFARX1 I_11927 (I205467,I2683,I205399,I205493,);
not I_11928 (I205501,I10414);
DFFARX1 I_11929 (I10429,I2683,I205399,I205527,);
not I_11930 (I205535,I205527);
nor I_11931 (I205552,I205535,I205433);
and I_11932 (I205569,I205552,I10414);
nor I_11933 (I205586,I205535,I205501);
nor I_11934 (I205382,I205493,I205586);
DFFARX1 I_11935 (I10414,I2683,I205399,I205626,);
nor I_11936 (I205634,I205626,I205493);
not I_11937 (I205651,I205634);
not I_11938 (I205668,I205626);
nor I_11939 (I205685,I205668,I205569);
DFFARX1 I_11940 (I205685,I2683,I205399,I205385,);
nand I_11941 (I205716,I10432,I10417);
and I_11942 (I205733,I205716,I10435);
DFFARX1 I_11943 (I205733,I2683,I205399,I205759,);
nor I_11944 (I205767,I205759,I205626);
DFFARX1 I_11945 (I205767,I2683,I205399,I205367,);
nand I_11946 (I205798,I205759,I205668);
nand I_11947 (I205376,I205651,I205798);
not I_11948 (I205829,I205759);
nor I_11949 (I205846,I205829,I205569);
DFFARX1 I_11950 (I205846,I2683,I205399,I205388,);
nor I_11951 (I205877,I10426,I10417);
or I_11952 (I205379,I205626,I205877);
nor I_11953 (I205370,I205759,I205877);
or I_11954 (I205373,I205493,I205877);
DFFARX1 I_11955 (I205877,I2683,I205399,I205391,);
not I_11956 (I205977,I2690);
DFFARX1 I_11957 (I383051,I2683,I205977,I206003,);
not I_11958 (I206011,I206003);
nand I_11959 (I206028,I383075,I383057);
and I_11960 (I206045,I206028,I383063);
DFFARX1 I_11961 (I206045,I2683,I205977,I206071,);
not I_11962 (I206079,I383069);
DFFARX1 I_11963 (I383054,I2683,I205977,I206105,);
not I_11964 (I206113,I206105);
nor I_11965 (I206130,I206113,I206011);
and I_11966 (I206147,I206130,I383069);
nor I_11967 (I206164,I206113,I206079);
nor I_11968 (I205960,I206071,I206164);
DFFARX1 I_11969 (I383066,I2683,I205977,I206204,);
nor I_11970 (I206212,I206204,I206071);
not I_11971 (I206229,I206212);
not I_11972 (I206246,I206204);
nor I_11973 (I206263,I206246,I206147);
DFFARX1 I_11974 (I206263,I2683,I205977,I205963,);
nand I_11975 (I206294,I383072,I383060);
and I_11976 (I206311,I206294,I383054);
DFFARX1 I_11977 (I206311,I2683,I205977,I206337,);
nor I_11978 (I206345,I206337,I206204);
DFFARX1 I_11979 (I206345,I2683,I205977,I205945,);
nand I_11980 (I206376,I206337,I206246);
nand I_11981 (I205954,I206229,I206376);
not I_11982 (I206407,I206337);
nor I_11983 (I206424,I206407,I206147);
DFFARX1 I_11984 (I206424,I2683,I205977,I205966,);
nor I_11985 (I206455,I383051,I383060);
or I_11986 (I205957,I206204,I206455);
nor I_11987 (I205948,I206337,I206455);
or I_11988 (I205951,I206071,I206455);
DFFARX1 I_11989 (I206455,I2683,I205977,I205969,);
not I_11990 (I206555,I2690);
DFFARX1 I_11991 (I165349,I2683,I206555,I206581,);
not I_11992 (I206589,I206581);
nand I_11993 (I206606,I165364,I165349);
and I_11994 (I206623,I206606,I165352);
DFFARX1 I_11995 (I206623,I2683,I206555,I206649,);
not I_11996 (I206657,I165352);
DFFARX1 I_11997 (I165361,I2683,I206555,I206683,);
not I_11998 (I206691,I206683);
nor I_11999 (I206708,I206691,I206589);
and I_12000 (I206725,I206708,I165352);
nor I_12001 (I206742,I206691,I206657);
nor I_12002 (I206538,I206649,I206742);
DFFARX1 I_12003 (I165355,I2683,I206555,I206782,);
nor I_12004 (I206790,I206782,I206649);
not I_12005 (I206807,I206790);
not I_12006 (I206824,I206782);
nor I_12007 (I206841,I206824,I206725);
DFFARX1 I_12008 (I206841,I2683,I206555,I206541,);
nand I_12009 (I206872,I165358,I165367);
and I_12010 (I206889,I206872,I165373);
DFFARX1 I_12011 (I206889,I2683,I206555,I206915,);
nor I_12012 (I206923,I206915,I206782);
DFFARX1 I_12013 (I206923,I2683,I206555,I206523,);
nand I_12014 (I206954,I206915,I206824);
nand I_12015 (I206532,I206807,I206954);
not I_12016 (I206985,I206915);
nor I_12017 (I207002,I206985,I206725);
DFFARX1 I_12018 (I207002,I2683,I206555,I206544,);
nor I_12019 (I207033,I165370,I165367);
or I_12020 (I206535,I206782,I207033);
nor I_12021 (I206526,I206915,I207033);
or I_12022 (I206529,I206649,I207033);
DFFARX1 I_12023 (I207033,I2683,I206555,I206547,);
not I_12024 (I207133,I2690);
DFFARX1 I_12025 (I1572,I2683,I207133,I207159,);
not I_12026 (I207167,I207159);
nand I_12027 (I207184,I2044,I1556);
and I_12028 (I207201,I207184,I2228);
DFFARX1 I_12029 (I207201,I2683,I207133,I207227,);
not I_12030 (I207235,I1468);
DFFARX1 I_12031 (I1932,I2683,I207133,I207261,);
not I_12032 (I207269,I207261);
nor I_12033 (I207286,I207269,I207167);
and I_12034 (I207303,I207286,I1468);
nor I_12035 (I207320,I207269,I207235);
nor I_12036 (I207116,I207227,I207320);
DFFARX1 I_12037 (I2148,I2683,I207133,I207360,);
nor I_12038 (I207368,I207360,I207227);
not I_12039 (I207385,I207368);
not I_12040 (I207402,I207360);
nor I_12041 (I207419,I207402,I207303);
DFFARX1 I_12042 (I207419,I2683,I207133,I207119,);
nand I_12043 (I207450,I1372,I1692);
and I_12044 (I207467,I207450,I2340);
DFFARX1 I_12045 (I207467,I2683,I207133,I207493,);
nor I_12046 (I207501,I207493,I207360);
DFFARX1 I_12047 (I207501,I2683,I207133,I207101,);
nand I_12048 (I207532,I207493,I207402);
nand I_12049 (I207110,I207385,I207532);
not I_12050 (I207563,I207493);
nor I_12051 (I207580,I207563,I207303);
DFFARX1 I_12052 (I207580,I2683,I207133,I207122,);
nor I_12053 (I207611,I1580,I1692);
or I_12054 (I207113,I207360,I207611);
nor I_12055 (I207104,I207493,I207611);
or I_12056 (I207107,I207227,I207611);
DFFARX1 I_12057 (I207611,I2683,I207133,I207125,);
not I_12058 (I207711,I2690);
DFFARX1 I_12059 (I114271,I2683,I207711,I207737,);
not I_12060 (I207745,I207737);
nand I_12061 (I207762,I114274,I114250);
and I_12062 (I207779,I207762,I114247);
DFFARX1 I_12063 (I207779,I2683,I207711,I207805,);
not I_12064 (I207813,I114253);
DFFARX1 I_12065 (I114247,I2683,I207711,I207839,);
not I_12066 (I207847,I207839);
nor I_12067 (I207864,I207847,I207745);
and I_12068 (I207881,I207864,I114253);
nor I_12069 (I207898,I207847,I207813);
nor I_12070 (I207694,I207805,I207898);
DFFARX1 I_12071 (I114256,I2683,I207711,I207938,);
nor I_12072 (I207946,I207938,I207805);
not I_12073 (I207963,I207946);
not I_12074 (I207980,I207938);
nor I_12075 (I207997,I207980,I207881);
DFFARX1 I_12076 (I207997,I2683,I207711,I207697,);
nand I_12077 (I208028,I114259,I114268);
and I_12078 (I208045,I208028,I114265);
DFFARX1 I_12079 (I208045,I2683,I207711,I208071,);
nor I_12080 (I208079,I208071,I207938);
DFFARX1 I_12081 (I208079,I2683,I207711,I207679,);
nand I_12082 (I208110,I208071,I207980);
nand I_12083 (I207688,I207963,I208110);
not I_12084 (I208141,I208071);
nor I_12085 (I208158,I208141,I207881);
DFFARX1 I_12086 (I208158,I2683,I207711,I207700,);
nor I_12087 (I208189,I114262,I114268);
or I_12088 (I207691,I207938,I208189);
nor I_12089 (I207682,I208071,I208189);
or I_12090 (I207685,I207805,I208189);
DFFARX1 I_12091 (I208189,I2683,I207711,I207703,);
not I_12092 (I208289,I2690);
DFFARX1 I_12093 (I126392,I2683,I208289,I208315,);
not I_12094 (I208323,I208315);
nand I_12095 (I208340,I126395,I126371);
and I_12096 (I208357,I208340,I126368);
DFFARX1 I_12097 (I208357,I2683,I208289,I208383,);
not I_12098 (I208391,I126374);
DFFARX1 I_12099 (I126368,I2683,I208289,I208417,);
not I_12100 (I208425,I208417);
nor I_12101 (I208442,I208425,I208323);
and I_12102 (I208459,I208442,I126374);
nor I_12103 (I208476,I208425,I208391);
nor I_12104 (I208272,I208383,I208476);
DFFARX1 I_12105 (I126377,I2683,I208289,I208516,);
nor I_12106 (I208524,I208516,I208383);
not I_12107 (I208541,I208524);
not I_12108 (I208558,I208516);
nor I_12109 (I208575,I208558,I208459);
DFFARX1 I_12110 (I208575,I2683,I208289,I208275,);
nand I_12111 (I208606,I126380,I126389);
and I_12112 (I208623,I208606,I126386);
DFFARX1 I_12113 (I208623,I2683,I208289,I208649,);
nor I_12114 (I208657,I208649,I208516);
DFFARX1 I_12115 (I208657,I2683,I208289,I208257,);
nand I_12116 (I208688,I208649,I208558);
nand I_12117 (I208266,I208541,I208688);
not I_12118 (I208719,I208649);
nor I_12119 (I208736,I208719,I208459);
DFFARX1 I_12120 (I208736,I2683,I208289,I208278,);
nor I_12121 (I208767,I126383,I126389);
or I_12122 (I208269,I208516,I208767);
nor I_12123 (I208260,I208649,I208767);
or I_12124 (I208263,I208383,I208767);
DFFARX1 I_12125 (I208767,I2683,I208289,I208281,);
not I_12126 (I208867,I2690);
DFFARX1 I_12127 (I359711,I2683,I208867,I208893,);
not I_12128 (I208901,I208893);
nand I_12129 (I208918,I359693,I359705);
and I_12130 (I208935,I208918,I359708);
DFFARX1 I_12131 (I208935,I2683,I208867,I208961,);
not I_12132 (I208969,I359702);
DFFARX1 I_12133 (I359699,I2683,I208867,I208995,);
not I_12134 (I209003,I208995);
nor I_12135 (I209020,I209003,I208901);
and I_12136 (I209037,I209020,I359702);
nor I_12137 (I209054,I209003,I208969);
nor I_12138 (I208850,I208961,I209054);
DFFARX1 I_12139 (I359717,I2683,I208867,I209094,);
nor I_12140 (I209102,I209094,I208961);
not I_12141 (I209119,I209102);
not I_12142 (I209136,I209094);
nor I_12143 (I209153,I209136,I209037);
DFFARX1 I_12144 (I209153,I2683,I208867,I208853,);
nand I_12145 (I209184,I359696,I359696);
and I_12146 (I209201,I209184,I359693);
DFFARX1 I_12147 (I209201,I2683,I208867,I209227,);
nor I_12148 (I209235,I209227,I209094);
DFFARX1 I_12149 (I209235,I2683,I208867,I208835,);
nand I_12150 (I209266,I209227,I209136);
nand I_12151 (I208844,I209119,I209266);
not I_12152 (I209297,I209227);
nor I_12153 (I209314,I209297,I209037);
DFFARX1 I_12154 (I209314,I2683,I208867,I208856,);
nor I_12155 (I209345,I359714,I359696);
or I_12156 (I208847,I209094,I209345);
nor I_12157 (I208838,I209227,I209345);
or I_12158 (I208841,I208961,I209345);
DFFARX1 I_12159 (I209345,I2683,I208867,I208859,);
not I_12160 (I209445,I2690);
DFFARX1 I_12161 (I125338,I2683,I209445,I209471,);
not I_12162 (I209479,I209471);
nand I_12163 (I209496,I125341,I125317);
and I_12164 (I209513,I209496,I125314);
DFFARX1 I_12165 (I209513,I2683,I209445,I209539,);
not I_12166 (I209547,I125320);
DFFARX1 I_12167 (I125314,I2683,I209445,I209573,);
not I_12168 (I209581,I209573);
nor I_12169 (I209598,I209581,I209479);
and I_12170 (I209615,I209598,I125320);
nor I_12171 (I209632,I209581,I209547);
nor I_12172 (I209428,I209539,I209632);
DFFARX1 I_12173 (I125323,I2683,I209445,I209672,);
nor I_12174 (I209680,I209672,I209539);
not I_12175 (I209697,I209680);
not I_12176 (I209714,I209672);
nor I_12177 (I209731,I209714,I209615);
DFFARX1 I_12178 (I209731,I2683,I209445,I209431,);
nand I_12179 (I209762,I125326,I125335);
and I_12180 (I209779,I209762,I125332);
DFFARX1 I_12181 (I209779,I2683,I209445,I209805,);
nor I_12182 (I209813,I209805,I209672);
DFFARX1 I_12183 (I209813,I2683,I209445,I209413,);
nand I_12184 (I209844,I209805,I209714);
nand I_12185 (I209422,I209697,I209844);
not I_12186 (I209875,I209805);
nor I_12187 (I209892,I209875,I209615);
DFFARX1 I_12188 (I209892,I2683,I209445,I209434,);
nor I_12189 (I209923,I125329,I125335);
or I_12190 (I209425,I209672,I209923);
nor I_12191 (I209416,I209805,I209923);
or I_12192 (I209419,I209539,I209923);
DFFARX1 I_12193 (I209923,I2683,I209445,I209437,);
not I_12194 (I210023,I2690);
DFFARX1 I_12195 (I391721,I2683,I210023,I210049,);
not I_12196 (I210057,I210049);
nand I_12197 (I210074,I391745,I391727);
and I_12198 (I210091,I210074,I391733);
DFFARX1 I_12199 (I210091,I2683,I210023,I210117,);
not I_12200 (I210125,I391739);
DFFARX1 I_12201 (I391724,I2683,I210023,I210151,);
not I_12202 (I210159,I210151);
nor I_12203 (I210176,I210159,I210057);
and I_12204 (I210193,I210176,I391739);
nor I_12205 (I210210,I210159,I210125);
nor I_12206 (I210006,I210117,I210210);
DFFARX1 I_12207 (I391736,I2683,I210023,I210250,);
nor I_12208 (I210258,I210250,I210117);
not I_12209 (I210275,I210258);
not I_12210 (I210292,I210250);
nor I_12211 (I210309,I210292,I210193);
DFFARX1 I_12212 (I210309,I2683,I210023,I210009,);
nand I_12213 (I210340,I391742,I391730);
and I_12214 (I210357,I210340,I391724);
DFFARX1 I_12215 (I210357,I2683,I210023,I210383,);
nor I_12216 (I210391,I210383,I210250);
DFFARX1 I_12217 (I210391,I2683,I210023,I209991,);
nand I_12218 (I210422,I210383,I210292);
nand I_12219 (I210000,I210275,I210422);
not I_12220 (I210453,I210383);
nor I_12221 (I210470,I210453,I210193);
DFFARX1 I_12222 (I210470,I2683,I210023,I210012,);
nor I_12223 (I210501,I391721,I391730);
or I_12224 (I210003,I210250,I210501);
nor I_12225 (I209994,I210383,I210501);
or I_12226 (I209997,I210117,I210501);
DFFARX1 I_12227 (I210501,I2683,I210023,I210015,);
not I_12228 (I210601,I2690);
DFFARX1 I_12229 (I148664,I2683,I210601,I210627,);
not I_12230 (I210635,I210627);
nand I_12231 (I210652,I148655,I148673);
and I_12232 (I210669,I210652,I148676);
DFFARX1 I_12233 (I210669,I2683,I210601,I210695,);
not I_12234 (I210703,I148670);
DFFARX1 I_12235 (I148658,I2683,I210601,I210729,);
not I_12236 (I210737,I210729);
nor I_12237 (I210754,I210737,I210635);
and I_12238 (I210771,I210754,I148670);
nor I_12239 (I210788,I210737,I210703);
nor I_12240 (I210584,I210695,I210788);
DFFARX1 I_12241 (I148667,I2683,I210601,I210828,);
nor I_12242 (I210836,I210828,I210695);
not I_12243 (I210853,I210836);
not I_12244 (I210870,I210828);
nor I_12245 (I210887,I210870,I210771);
DFFARX1 I_12246 (I210887,I2683,I210601,I210587,);
nand I_12247 (I210918,I148682,I148679);
and I_12248 (I210935,I210918,I148661);
DFFARX1 I_12249 (I210935,I2683,I210601,I210961,);
nor I_12250 (I210969,I210961,I210828);
DFFARX1 I_12251 (I210969,I2683,I210601,I210569,);
nand I_12252 (I211000,I210961,I210870);
nand I_12253 (I210578,I210853,I211000);
not I_12254 (I211031,I210961);
nor I_12255 (I211048,I211031,I210771);
DFFARX1 I_12256 (I211048,I2683,I210601,I210590,);
nor I_12257 (I211079,I148655,I148679);
or I_12258 (I210581,I210828,I211079);
nor I_12259 (I210572,I210961,I211079);
or I_12260 (I210575,I210695,I211079);
DFFARX1 I_12261 (I211079,I2683,I210601,I210593,);
not I_12262 (I211179,I2690);
DFFARX1 I_12263 (I87394,I2683,I211179,I211205,);
not I_12264 (I211213,I211205);
nand I_12265 (I211230,I87397,I87373);
and I_12266 (I211247,I211230,I87370);
DFFARX1 I_12267 (I211247,I2683,I211179,I211273,);
not I_12268 (I211281,I87376);
DFFARX1 I_12269 (I87370,I2683,I211179,I211307,);
not I_12270 (I211315,I211307);
nor I_12271 (I211332,I211315,I211213);
and I_12272 (I211349,I211332,I87376);
nor I_12273 (I211366,I211315,I211281);
nor I_12274 (I211162,I211273,I211366);
DFFARX1 I_12275 (I87379,I2683,I211179,I211406,);
nor I_12276 (I211414,I211406,I211273);
not I_12277 (I211431,I211414);
not I_12278 (I211448,I211406);
nor I_12279 (I211465,I211448,I211349);
DFFARX1 I_12280 (I211465,I2683,I211179,I211165,);
nand I_12281 (I211496,I87382,I87391);
and I_12282 (I211513,I211496,I87388);
DFFARX1 I_12283 (I211513,I2683,I211179,I211539,);
nor I_12284 (I211547,I211539,I211406);
DFFARX1 I_12285 (I211547,I2683,I211179,I211147,);
nand I_12286 (I211578,I211539,I211448);
nand I_12287 (I211156,I211431,I211578);
not I_12288 (I211609,I211539);
nor I_12289 (I211626,I211609,I211349);
DFFARX1 I_12290 (I211626,I2683,I211179,I211168,);
nor I_12291 (I211657,I87385,I87391);
or I_12292 (I211159,I211406,I211657);
nor I_12293 (I211150,I211539,I211657);
or I_12294 (I211153,I211273,I211657);
DFFARX1 I_12295 (I211657,I2683,I211179,I211171,);
not I_12296 (I211757,I2690);
DFFARX1 I_12297 (I250296,I2683,I211757,I211783,);
not I_12298 (I211791,I211783);
nand I_12299 (I211808,I250284,I250302);
and I_12300 (I211825,I211808,I250299);
DFFARX1 I_12301 (I211825,I2683,I211757,I211851,);
not I_12302 (I211859,I250290);
DFFARX1 I_12303 (I250287,I2683,I211757,I211885,);
not I_12304 (I211893,I211885);
nor I_12305 (I211910,I211893,I211791);
and I_12306 (I211927,I211910,I250290);
nor I_12307 (I211944,I211893,I211859);
nor I_12308 (I211740,I211851,I211944);
DFFARX1 I_12309 (I250281,I2683,I211757,I211984,);
nor I_12310 (I211992,I211984,I211851);
not I_12311 (I212009,I211992);
not I_12312 (I212026,I211984);
nor I_12313 (I212043,I212026,I211927);
DFFARX1 I_12314 (I212043,I2683,I211757,I211743,);
nand I_12315 (I212074,I250281,I250284);
and I_12316 (I212091,I212074,I250287);
DFFARX1 I_12317 (I212091,I2683,I211757,I212117,);
nor I_12318 (I212125,I212117,I211984);
DFFARX1 I_12319 (I212125,I2683,I211757,I211725,);
nand I_12320 (I212156,I212117,I212026);
nand I_12321 (I211734,I212009,I212156);
not I_12322 (I212187,I212117);
nor I_12323 (I212204,I212187,I211927);
DFFARX1 I_12324 (I212204,I2683,I211757,I211746,);
nor I_12325 (I212235,I250293,I250284);
or I_12326 (I211737,I211984,I212235);
nor I_12327 (I211728,I212117,I212235);
or I_12328 (I211731,I211851,I212235);
DFFARX1 I_12329 (I212235,I2683,I211757,I211749,);
not I_12330 (I212335,I2690);
DFFARX1 I_12331 (I268214,I2683,I212335,I212361,);
not I_12332 (I212369,I212361);
nand I_12333 (I212386,I268202,I268220);
and I_12334 (I212403,I212386,I268217);
DFFARX1 I_12335 (I212403,I2683,I212335,I212429,);
not I_12336 (I212437,I268208);
DFFARX1 I_12337 (I268205,I2683,I212335,I212463,);
not I_12338 (I212471,I212463);
nor I_12339 (I212488,I212471,I212369);
and I_12340 (I212505,I212488,I268208);
nor I_12341 (I212522,I212471,I212437);
nor I_12342 (I212318,I212429,I212522);
DFFARX1 I_12343 (I268199,I2683,I212335,I212562,);
nor I_12344 (I212570,I212562,I212429);
not I_12345 (I212587,I212570);
not I_12346 (I212604,I212562);
nor I_12347 (I212621,I212604,I212505);
DFFARX1 I_12348 (I212621,I2683,I212335,I212321,);
nand I_12349 (I212652,I268199,I268202);
and I_12350 (I212669,I212652,I268205);
DFFARX1 I_12351 (I212669,I2683,I212335,I212695,);
nor I_12352 (I212703,I212695,I212562);
DFFARX1 I_12353 (I212703,I2683,I212335,I212303,);
nand I_12354 (I212734,I212695,I212604);
nand I_12355 (I212312,I212587,I212734);
not I_12356 (I212765,I212695);
nor I_12357 (I212782,I212765,I212505);
DFFARX1 I_12358 (I212782,I2683,I212335,I212324,);
nor I_12359 (I212813,I268211,I268202);
or I_12360 (I212315,I212562,I212813);
nor I_12361 (I212306,I212695,I212813);
or I_12362 (I212309,I212429,I212813);
DFFARX1 I_12363 (I212813,I2683,I212335,I212327,);
not I_12364 (I212913,I2690);
DFFARX1 I_12365 (I414086,I2683,I212913,I212939,);
not I_12366 (I212947,I212939);
nand I_12367 (I212964,I414071,I414059);
and I_12368 (I212981,I212964,I414074);
DFFARX1 I_12369 (I212981,I2683,I212913,I213007,);
not I_12370 (I213015,I414059);
DFFARX1 I_12371 (I414077,I2683,I212913,I213041,);
not I_12372 (I213049,I213041);
nor I_12373 (I213066,I213049,I212947);
and I_12374 (I213083,I213066,I414059);
nor I_12375 (I213100,I213049,I213015);
nor I_12376 (I212896,I213007,I213100);
DFFARX1 I_12377 (I414065,I2683,I212913,I213140,);
nor I_12378 (I213148,I213140,I213007);
not I_12379 (I213165,I213148);
not I_12380 (I213182,I213140);
nor I_12381 (I213199,I213182,I213083);
DFFARX1 I_12382 (I213199,I2683,I212913,I212899,);
nand I_12383 (I213230,I414062,I414068);
and I_12384 (I213247,I213230,I414083);
DFFARX1 I_12385 (I213247,I2683,I212913,I213273,);
nor I_12386 (I213281,I213273,I213140);
DFFARX1 I_12387 (I213281,I2683,I212913,I212881,);
nand I_12388 (I213312,I213273,I213182);
nand I_12389 (I212890,I213165,I213312);
not I_12390 (I213343,I213273);
nor I_12391 (I213360,I213343,I213083);
DFFARX1 I_12392 (I213360,I2683,I212913,I212902,);
nor I_12393 (I213391,I414080,I414068);
or I_12394 (I212893,I213140,I213391);
nor I_12395 (I212884,I213273,I213391);
or I_12396 (I212887,I213007,I213391);
DFFARX1 I_12397 (I213391,I2683,I212913,I212905,);
not I_12398 (I213491,I2690);
DFFARX1 I_12399 (I23589,I2683,I213491,I213517,);
not I_12400 (I213525,I213517);
nand I_12401 (I213542,I23598,I23607);
and I_12402 (I213559,I213542,I23586);
DFFARX1 I_12403 (I213559,I2683,I213491,I213585,);
not I_12404 (I213593,I23589);
DFFARX1 I_12405 (I23604,I2683,I213491,I213619,);
not I_12406 (I213627,I213619);
nor I_12407 (I213644,I213627,I213525);
and I_12408 (I213661,I213644,I23589);
nor I_12409 (I213678,I213627,I213593);
nor I_12410 (I213474,I213585,I213678);
DFFARX1 I_12411 (I23595,I2683,I213491,I213718,);
nor I_12412 (I213726,I213718,I213585);
not I_12413 (I213743,I213726);
not I_12414 (I213760,I213718);
nor I_12415 (I213777,I213760,I213661);
DFFARX1 I_12416 (I213777,I2683,I213491,I213477,);
nand I_12417 (I213808,I23610,I23586);
and I_12418 (I213825,I213808,I23592);
DFFARX1 I_12419 (I213825,I2683,I213491,I213851,);
nor I_12420 (I213859,I213851,I213718);
DFFARX1 I_12421 (I213859,I2683,I213491,I213459,);
nand I_12422 (I213890,I213851,I213760);
nand I_12423 (I213468,I213743,I213890);
not I_12424 (I213921,I213851);
nor I_12425 (I213938,I213921,I213661);
DFFARX1 I_12426 (I213938,I2683,I213491,I213480,);
nor I_12427 (I213969,I23601,I23586);
or I_12428 (I213471,I213718,I213969);
nor I_12429 (I213462,I213851,I213969);
or I_12430 (I213465,I213585,I213969);
DFFARX1 I_12431 (I213969,I2683,I213491,I213483,);
not I_12432 (I214069,I2690);
DFFARX1 I_12433 (I103204,I2683,I214069,I214095,);
not I_12434 (I214103,I214095);
nand I_12435 (I214120,I103207,I103183);
and I_12436 (I214137,I214120,I103180);
DFFARX1 I_12437 (I214137,I2683,I214069,I214163,);
not I_12438 (I214171,I103186);
DFFARX1 I_12439 (I103180,I2683,I214069,I214197,);
not I_12440 (I214205,I214197);
nor I_12441 (I214222,I214205,I214103);
and I_12442 (I214239,I214222,I103186);
nor I_12443 (I214256,I214205,I214171);
nor I_12444 (I214052,I214163,I214256);
DFFARX1 I_12445 (I103189,I2683,I214069,I214296,);
nor I_12446 (I214304,I214296,I214163);
not I_12447 (I214321,I214304);
not I_12448 (I214338,I214296);
nor I_12449 (I214355,I214338,I214239);
DFFARX1 I_12450 (I214355,I2683,I214069,I214055,);
nand I_12451 (I214386,I103192,I103201);
and I_12452 (I214403,I214386,I103198);
DFFARX1 I_12453 (I214403,I2683,I214069,I214429,);
nor I_12454 (I214437,I214429,I214296);
DFFARX1 I_12455 (I214437,I2683,I214069,I214037,);
nand I_12456 (I214468,I214429,I214338);
nand I_12457 (I214046,I214321,I214468);
not I_12458 (I214499,I214429);
nor I_12459 (I214516,I214499,I214239);
DFFARX1 I_12460 (I214516,I2683,I214069,I214058,);
nor I_12461 (I214547,I103195,I103201);
or I_12462 (I214049,I214296,I214547);
nor I_12463 (I214040,I214429,I214547);
or I_12464 (I214043,I214163,I214547);
DFFARX1 I_12465 (I214547,I2683,I214069,I214061,);
not I_12466 (I214647,I2690);
DFFARX1 I_12467 (I101623,I2683,I214647,I214673,);
not I_12468 (I214681,I214673);
nand I_12469 (I214698,I101626,I101602);
and I_12470 (I214715,I214698,I101599);
DFFARX1 I_12471 (I214715,I2683,I214647,I214741,);
not I_12472 (I214749,I101605);
DFFARX1 I_12473 (I101599,I2683,I214647,I214775,);
not I_12474 (I214783,I214775);
nor I_12475 (I214800,I214783,I214681);
and I_12476 (I214817,I214800,I101605);
nor I_12477 (I214834,I214783,I214749);
nor I_12478 (I214630,I214741,I214834);
DFFARX1 I_12479 (I101608,I2683,I214647,I214874,);
nor I_12480 (I214882,I214874,I214741);
not I_12481 (I214899,I214882);
not I_12482 (I214916,I214874);
nor I_12483 (I214933,I214916,I214817);
DFFARX1 I_12484 (I214933,I2683,I214647,I214633,);
nand I_12485 (I214964,I101611,I101620);
and I_12486 (I214981,I214964,I101617);
DFFARX1 I_12487 (I214981,I2683,I214647,I215007,);
nor I_12488 (I215015,I215007,I214874);
DFFARX1 I_12489 (I215015,I2683,I214647,I214615,);
nand I_12490 (I215046,I215007,I214916);
nand I_12491 (I214624,I214899,I215046);
not I_12492 (I215077,I215007);
nor I_12493 (I215094,I215077,I214817);
DFFARX1 I_12494 (I215094,I2683,I214647,I214636,);
nor I_12495 (I215125,I101614,I101620);
or I_12496 (I214627,I214874,I215125);
nor I_12497 (I214618,I215007,I215125);
or I_12498 (I214621,I214741,I215125);
DFFARX1 I_12499 (I215125,I2683,I214647,I214639,);
not I_12500 (I215225,I2690);
DFFARX1 I_12501 (I185715,I2683,I215225,I215251,);
not I_12502 (I215259,I215251);
nand I_12503 (I215276,I185724,I185733);
and I_12504 (I215293,I215276,I185739);
DFFARX1 I_12505 (I215293,I2683,I215225,I215319,);
not I_12506 (I215327,I185736);
DFFARX1 I_12507 (I185721,I2683,I215225,I215353,);
not I_12508 (I215361,I215353);
nor I_12509 (I215378,I215361,I215259);
and I_12510 (I215395,I215378,I185736);
nor I_12511 (I215412,I215361,I215327);
nor I_12512 (I215208,I215319,I215412);
DFFARX1 I_12513 (I185730,I2683,I215225,I215452,);
nor I_12514 (I215460,I215452,I215319);
not I_12515 (I215477,I215460);
not I_12516 (I215494,I215452);
nor I_12517 (I215511,I215494,I215395);
DFFARX1 I_12518 (I215511,I2683,I215225,I215211,);
nand I_12519 (I215542,I185727,I185718);
and I_12520 (I215559,I215542,I185715);
DFFARX1 I_12521 (I215559,I2683,I215225,I215585,);
nor I_12522 (I215593,I215585,I215452);
DFFARX1 I_12523 (I215593,I2683,I215225,I215193,);
nand I_12524 (I215624,I215585,I215494);
nand I_12525 (I215202,I215477,I215624);
not I_12526 (I215655,I215585);
nor I_12527 (I215672,I215655,I215395);
DFFARX1 I_12528 (I215672,I2683,I215225,I215214,);
nor I_12529 (I215703,I185718,I185718);
or I_12530 (I215205,I215452,I215703);
nor I_12531 (I215196,I215585,I215703);
or I_12532 (I215199,I215319,I215703);
DFFARX1 I_12533 (I215703,I2683,I215225,I215217,);
not I_12534 (I215803,I2690);
DFFARX1 I_12535 (I69724,I2683,I215803,I215829,);
not I_12536 (I215837,I215829);
nand I_12537 (I215854,I69727,I69748);
and I_12538 (I215871,I215854,I69736);
DFFARX1 I_12539 (I215871,I2683,I215803,I215897,);
not I_12540 (I215905,I69733);
DFFARX1 I_12541 (I69724,I2683,I215803,I215931,);
not I_12542 (I215939,I215931);
nor I_12543 (I215956,I215939,I215837);
and I_12544 (I215973,I215956,I69733);
nor I_12545 (I215990,I215939,I215905);
nor I_12546 (I215786,I215897,I215990);
DFFARX1 I_12547 (I69742,I2683,I215803,I216030,);
nor I_12548 (I216038,I216030,I215897);
not I_12549 (I216055,I216038);
not I_12550 (I216072,I216030);
nor I_12551 (I216089,I216072,I215973);
DFFARX1 I_12552 (I216089,I2683,I215803,I215789,);
nand I_12553 (I216120,I69727,I69730);
and I_12554 (I216137,I216120,I69739);
DFFARX1 I_12555 (I216137,I2683,I215803,I216163,);
nor I_12556 (I216171,I216163,I216030);
DFFARX1 I_12557 (I216171,I2683,I215803,I215771,);
nand I_12558 (I216202,I216163,I216072);
nand I_12559 (I215780,I216055,I216202);
not I_12560 (I216233,I216163);
nor I_12561 (I216250,I216233,I215973);
DFFARX1 I_12562 (I216250,I2683,I215803,I215792,);
nor I_12563 (I216281,I69745,I69730);
or I_12564 (I215783,I216030,I216281);
nor I_12565 (I215774,I216163,I216281);
or I_12566 (I215777,I215897,I216281);
DFFARX1 I_12567 (I216281,I2683,I215803,I215795,);
not I_12568 (I216381,I2690);
DFFARX1 I_12569 (I398616,I2683,I216381,I216407,);
not I_12570 (I216415,I216407);
nand I_12571 (I216432,I398601,I398589);
and I_12572 (I216449,I216432,I398604);
DFFARX1 I_12573 (I216449,I2683,I216381,I216475,);
not I_12574 (I216483,I398589);
DFFARX1 I_12575 (I398607,I2683,I216381,I216509,);
not I_12576 (I216517,I216509);
nor I_12577 (I216534,I216517,I216415);
and I_12578 (I216551,I216534,I398589);
nor I_12579 (I216568,I216517,I216483);
nor I_12580 (I216364,I216475,I216568);
DFFARX1 I_12581 (I398595,I2683,I216381,I216608,);
nor I_12582 (I216616,I216608,I216475);
not I_12583 (I216633,I216616);
not I_12584 (I216650,I216608);
nor I_12585 (I216667,I216650,I216551);
DFFARX1 I_12586 (I216667,I2683,I216381,I216367,);
nand I_12587 (I216698,I398592,I398598);
and I_12588 (I216715,I216698,I398613);
DFFARX1 I_12589 (I216715,I2683,I216381,I216741,);
nor I_12590 (I216749,I216741,I216608);
DFFARX1 I_12591 (I216749,I2683,I216381,I216349,);
nand I_12592 (I216780,I216741,I216650);
nand I_12593 (I216358,I216633,I216780);
not I_12594 (I216811,I216741);
nor I_12595 (I216828,I216811,I216551);
DFFARX1 I_12596 (I216828,I2683,I216381,I216370,);
nor I_12597 (I216859,I398610,I398598);
or I_12598 (I216361,I216608,I216859);
nor I_12599 (I216352,I216741,I216859);
or I_12600 (I216355,I216475,I216859);
DFFARX1 I_12601 (I216859,I2683,I216381,I216373,);
not I_12602 (I216959,I2690);
DFFARX1 I_12603 (I152472,I2683,I216959,I216985,);
not I_12604 (I216993,I216985);
nand I_12605 (I217010,I152463,I152481);
and I_12606 (I217027,I217010,I152484);
DFFARX1 I_12607 (I217027,I2683,I216959,I217053,);
not I_12608 (I217061,I152478);
DFFARX1 I_12609 (I152466,I2683,I216959,I217087,);
not I_12610 (I217095,I217087);
nor I_12611 (I217112,I217095,I216993);
and I_12612 (I217129,I217112,I152478);
nor I_12613 (I217146,I217095,I217061);
nor I_12614 (I216942,I217053,I217146);
DFFARX1 I_12615 (I152475,I2683,I216959,I217186,);
nor I_12616 (I217194,I217186,I217053);
not I_12617 (I217211,I217194);
not I_12618 (I217228,I217186);
nor I_12619 (I217245,I217228,I217129);
DFFARX1 I_12620 (I217245,I2683,I216959,I216945,);
nand I_12621 (I217276,I152490,I152487);
and I_12622 (I217293,I217276,I152469);
DFFARX1 I_12623 (I217293,I2683,I216959,I217319,);
nor I_12624 (I217327,I217319,I217186);
DFFARX1 I_12625 (I217327,I2683,I216959,I216927,);
nand I_12626 (I217358,I217319,I217228);
nand I_12627 (I216936,I217211,I217358);
not I_12628 (I217389,I217319);
nor I_12629 (I217406,I217389,I217129);
DFFARX1 I_12630 (I217406,I2683,I216959,I216948,);
nor I_12631 (I217437,I152463,I152487);
or I_12632 (I216939,I217186,I217437);
nor I_12633 (I216930,I217319,I217437);
or I_12634 (I216933,I217053,I217437);
DFFARX1 I_12635 (I217437,I2683,I216959,I216951,);
not I_12636 (I217537,I2690);
DFFARX1 I_12637 (I355665,I2683,I217537,I217563,);
not I_12638 (I217571,I217563);
nand I_12639 (I217588,I355647,I355659);
and I_12640 (I217605,I217588,I355662);
DFFARX1 I_12641 (I217605,I2683,I217537,I217631,);
not I_12642 (I217639,I355656);
DFFARX1 I_12643 (I355653,I2683,I217537,I217665,);
not I_12644 (I217673,I217665);
nor I_12645 (I217690,I217673,I217571);
and I_12646 (I217707,I217690,I355656);
nor I_12647 (I217724,I217673,I217639);
nor I_12648 (I217520,I217631,I217724);
DFFARX1 I_12649 (I355671,I2683,I217537,I217764,);
nor I_12650 (I217772,I217764,I217631);
not I_12651 (I217789,I217772);
not I_12652 (I217806,I217764);
nor I_12653 (I217823,I217806,I217707);
DFFARX1 I_12654 (I217823,I2683,I217537,I217523,);
nand I_12655 (I217854,I355650,I355650);
and I_12656 (I217871,I217854,I355647);
DFFARX1 I_12657 (I217871,I2683,I217537,I217897,);
nor I_12658 (I217905,I217897,I217764);
DFFARX1 I_12659 (I217905,I2683,I217537,I217505,);
nand I_12660 (I217936,I217897,I217806);
nand I_12661 (I217514,I217789,I217936);
not I_12662 (I217967,I217897);
nor I_12663 (I217984,I217967,I217707);
DFFARX1 I_12664 (I217984,I2683,I217537,I217526,);
nor I_12665 (I218015,I355668,I355650);
or I_12666 (I217517,I217764,I218015);
nor I_12667 (I217508,I217897,I218015);
or I_12668 (I217511,I217631,I218015);
DFFARX1 I_12669 (I218015,I2683,I217537,I217529,);
not I_12670 (I218115,I2690);
DFFARX1 I_12671 (I3294,I2683,I218115,I218141,);
not I_12672 (I218149,I218141);
nand I_12673 (I218166,I3297,I3309);
and I_12674 (I218183,I218166,I3288);
DFFARX1 I_12675 (I218183,I2683,I218115,I218209,);
not I_12676 (I218217,I3288);
DFFARX1 I_12677 (I3291,I2683,I218115,I218243,);
not I_12678 (I218251,I218243);
nor I_12679 (I218268,I218251,I218149);
and I_12680 (I218285,I218268,I3288);
nor I_12681 (I218302,I218251,I218217);
nor I_12682 (I218098,I218209,I218302);
DFFARX1 I_12683 (I3303,I2683,I218115,I218342,);
nor I_12684 (I218350,I218342,I218209);
not I_12685 (I218367,I218350);
not I_12686 (I218384,I218342);
nor I_12687 (I218401,I218384,I218285);
DFFARX1 I_12688 (I218401,I2683,I218115,I218101,);
nand I_12689 (I218432,I3306,I3291);
and I_12690 (I218449,I218432,I3300);
DFFARX1 I_12691 (I218449,I2683,I218115,I218475,);
nor I_12692 (I218483,I218475,I218342);
DFFARX1 I_12693 (I218483,I2683,I218115,I218083,);
nand I_12694 (I218514,I218475,I218384);
nand I_12695 (I218092,I218367,I218514);
not I_12696 (I218545,I218475);
nor I_12697 (I218562,I218545,I218285);
DFFARX1 I_12698 (I218562,I2683,I218115,I218104,);
nor I_12699 (I218593,I3294,I3291);
or I_12700 (I218095,I218342,I218593);
nor I_12701 (I218086,I218475,I218593);
or I_12702 (I218089,I218209,I218593);
DFFARX1 I_12703 (I218593,I2683,I218115,I218107,);
not I_12704 (I218693,I2690);
DFFARX1 I_12705 (I134520,I2683,I218693,I218719,);
not I_12706 (I218727,I218719);
nand I_12707 (I218744,I134511,I134529);
and I_12708 (I218761,I218744,I134532);
DFFARX1 I_12709 (I218761,I2683,I218693,I218787,);
not I_12710 (I218795,I134526);
DFFARX1 I_12711 (I134514,I2683,I218693,I218821,);
not I_12712 (I218829,I218821);
nor I_12713 (I218846,I218829,I218727);
and I_12714 (I218863,I218846,I134526);
nor I_12715 (I218880,I218829,I218795);
nor I_12716 (I218676,I218787,I218880);
DFFARX1 I_12717 (I134523,I2683,I218693,I218920,);
nor I_12718 (I218928,I218920,I218787);
not I_12719 (I218945,I218928);
not I_12720 (I218962,I218920);
nor I_12721 (I218979,I218962,I218863);
DFFARX1 I_12722 (I218979,I2683,I218693,I218679,);
nand I_12723 (I219010,I134538,I134535);
and I_12724 (I219027,I219010,I134517);
DFFARX1 I_12725 (I219027,I2683,I218693,I219053,);
nor I_12726 (I219061,I219053,I218920);
DFFARX1 I_12727 (I219061,I2683,I218693,I218661,);
nand I_12728 (I219092,I219053,I218962);
nand I_12729 (I218670,I218945,I219092);
not I_12730 (I219123,I219053);
nor I_12731 (I219140,I219123,I218863);
DFFARX1 I_12732 (I219140,I2683,I218693,I218682,);
nor I_12733 (I219171,I134511,I134535);
or I_12734 (I218673,I218920,I219171);
nor I_12735 (I218664,I219053,I219171);
or I_12736 (I218667,I218787,I219171);
DFFARX1 I_12737 (I219171,I2683,I218693,I218685,);
not I_12738 (I219271,I2690);
DFFARX1 I_12739 (I70914,I2683,I219271,I219297,);
not I_12740 (I219305,I219297);
nand I_12741 (I219322,I70917,I70938);
and I_12742 (I219339,I219322,I70926);
DFFARX1 I_12743 (I219339,I2683,I219271,I219365,);
not I_12744 (I219373,I70923);
DFFARX1 I_12745 (I70914,I2683,I219271,I219399,);
not I_12746 (I219407,I219399);
nor I_12747 (I219424,I219407,I219305);
and I_12748 (I219441,I219424,I70923);
nor I_12749 (I219458,I219407,I219373);
nor I_12750 (I219254,I219365,I219458);
DFFARX1 I_12751 (I70932,I2683,I219271,I219498,);
nor I_12752 (I219506,I219498,I219365);
not I_12753 (I219523,I219506);
not I_12754 (I219540,I219498);
nor I_12755 (I219557,I219540,I219441);
DFFARX1 I_12756 (I219557,I2683,I219271,I219257,);
nand I_12757 (I219588,I70917,I70920);
and I_12758 (I219605,I219588,I70929);
DFFARX1 I_12759 (I219605,I2683,I219271,I219631,);
nor I_12760 (I219639,I219631,I219498);
DFFARX1 I_12761 (I219639,I2683,I219271,I219239,);
nand I_12762 (I219670,I219631,I219540);
nand I_12763 (I219248,I219523,I219670);
not I_12764 (I219701,I219631);
nor I_12765 (I219718,I219701,I219441);
DFFARX1 I_12766 (I219718,I2683,I219271,I219260,);
nor I_12767 (I219749,I70935,I70920);
or I_12768 (I219251,I219498,I219749);
nor I_12769 (I219242,I219631,I219749);
or I_12770 (I219245,I219365,I219749);
DFFARX1 I_12771 (I219749,I2683,I219271,I219263,);
not I_12772 (I219849,I2690);
DFFARX1 I_12773 (I249242,I2683,I219849,I219875,);
not I_12774 (I219883,I219875);
nand I_12775 (I219900,I249230,I249248);
and I_12776 (I219917,I219900,I249245);
DFFARX1 I_12777 (I219917,I2683,I219849,I219943,);
not I_12778 (I219951,I249236);
DFFARX1 I_12779 (I249233,I2683,I219849,I219977,);
not I_12780 (I219985,I219977);
nor I_12781 (I220002,I219985,I219883);
and I_12782 (I220019,I220002,I249236);
nor I_12783 (I220036,I219985,I219951);
nor I_12784 (I219832,I219943,I220036);
DFFARX1 I_12785 (I249227,I2683,I219849,I220076,);
nor I_12786 (I220084,I220076,I219943);
not I_12787 (I220101,I220084);
not I_12788 (I220118,I220076);
nor I_12789 (I220135,I220118,I220019);
DFFARX1 I_12790 (I220135,I2683,I219849,I219835,);
nand I_12791 (I220166,I249227,I249230);
and I_12792 (I220183,I220166,I249233);
DFFARX1 I_12793 (I220183,I2683,I219849,I220209,);
nor I_12794 (I220217,I220209,I220076);
DFFARX1 I_12795 (I220217,I2683,I219849,I219817,);
nand I_12796 (I220248,I220209,I220118);
nand I_12797 (I219826,I220101,I220248);
not I_12798 (I220279,I220209);
nor I_12799 (I220296,I220279,I220019);
DFFARX1 I_12800 (I220296,I2683,I219849,I219838,);
nor I_12801 (I220327,I249239,I249230);
or I_12802 (I219829,I220076,I220327);
nor I_12803 (I219820,I220209,I220327);
or I_12804 (I219823,I219943,I220327);
DFFARX1 I_12805 (I220327,I2683,I219849,I219841,);
not I_12806 (I220427,I2690);
DFFARX1 I_12807 (I284662,I2683,I220427,I220453,);
not I_12808 (I220461,I220453);
nand I_12809 (I220478,I284638,I284653);
and I_12810 (I220495,I220478,I284665);
DFFARX1 I_12811 (I220495,I2683,I220427,I220521,);
not I_12812 (I220529,I284650);
DFFARX1 I_12813 (I284641,I2683,I220427,I220555,);
not I_12814 (I220563,I220555);
nor I_12815 (I220580,I220563,I220461);
and I_12816 (I220597,I220580,I284650);
nor I_12817 (I220614,I220563,I220529);
nor I_12818 (I220410,I220521,I220614);
DFFARX1 I_12819 (I284638,I2683,I220427,I220654,);
nor I_12820 (I220662,I220654,I220521);
not I_12821 (I220679,I220662);
not I_12822 (I220696,I220654);
nor I_12823 (I220713,I220696,I220597);
DFFARX1 I_12824 (I220713,I2683,I220427,I220413,);
nand I_12825 (I220744,I284656,I284647);
and I_12826 (I220761,I220744,I284659);
DFFARX1 I_12827 (I220761,I2683,I220427,I220787,);
nor I_12828 (I220795,I220787,I220654);
DFFARX1 I_12829 (I220795,I2683,I220427,I220395,);
nand I_12830 (I220826,I220787,I220696);
nand I_12831 (I220404,I220679,I220826);
not I_12832 (I220857,I220787);
nor I_12833 (I220874,I220857,I220597);
DFFARX1 I_12834 (I220874,I2683,I220427,I220416,);
nor I_12835 (I220905,I284644,I284647);
or I_12836 (I220407,I220654,I220905);
nor I_12837 (I220398,I220787,I220905);
or I_12838 (I220401,I220521,I220905);
DFFARX1 I_12839 (I220905,I2683,I220427,I220419,);
not I_12840 (I221005,I2690);
DFFARX1 I_12841 (I363179,I2683,I221005,I221031,);
not I_12842 (I221039,I221031);
nand I_12843 (I221056,I363161,I363173);
and I_12844 (I221073,I221056,I363176);
DFFARX1 I_12845 (I221073,I2683,I221005,I221099,);
not I_12846 (I221107,I363170);
DFFARX1 I_12847 (I363167,I2683,I221005,I221133,);
not I_12848 (I221141,I221133);
nor I_12849 (I221158,I221141,I221039);
and I_12850 (I221175,I221158,I363170);
nor I_12851 (I221192,I221141,I221107);
nor I_12852 (I220988,I221099,I221192);
DFFARX1 I_12853 (I363185,I2683,I221005,I221232,);
nor I_12854 (I221240,I221232,I221099);
not I_12855 (I221257,I221240);
not I_12856 (I221274,I221232);
nor I_12857 (I221291,I221274,I221175);
DFFARX1 I_12858 (I221291,I2683,I221005,I220991,);
nand I_12859 (I221322,I363164,I363164);
and I_12860 (I221339,I221322,I363161);
DFFARX1 I_12861 (I221339,I2683,I221005,I221365,);
nor I_12862 (I221373,I221365,I221232);
DFFARX1 I_12863 (I221373,I2683,I221005,I220973,);
nand I_12864 (I221404,I221365,I221274);
nand I_12865 (I220982,I221257,I221404);
not I_12866 (I221435,I221365);
nor I_12867 (I221452,I221435,I221175);
DFFARX1 I_12868 (I221452,I2683,I221005,I220994,);
nor I_12869 (I221483,I363182,I363164);
or I_12870 (I220985,I221232,I221483);
nor I_12871 (I220976,I221365,I221483);
or I_12872 (I220979,I221099,I221483);
DFFARX1 I_12873 (I221483,I2683,I221005,I220997,);
not I_12874 (I221583,I2690);
DFFARX1 I_12875 (I38345,I2683,I221583,I221609,);
not I_12876 (I221617,I221609);
nand I_12877 (I221634,I38354,I38363);
and I_12878 (I221651,I221634,I38342);
DFFARX1 I_12879 (I221651,I2683,I221583,I221677,);
not I_12880 (I221685,I38345);
DFFARX1 I_12881 (I38360,I2683,I221583,I221711,);
not I_12882 (I221719,I221711);
nor I_12883 (I221736,I221719,I221617);
and I_12884 (I221753,I221736,I38345);
nor I_12885 (I221770,I221719,I221685);
nor I_12886 (I221566,I221677,I221770);
DFFARX1 I_12887 (I38351,I2683,I221583,I221810,);
nor I_12888 (I221818,I221810,I221677);
not I_12889 (I221835,I221818);
not I_12890 (I221852,I221810);
nor I_12891 (I221869,I221852,I221753);
DFFARX1 I_12892 (I221869,I2683,I221583,I221569,);
nand I_12893 (I221900,I38366,I38342);
and I_12894 (I221917,I221900,I38348);
DFFARX1 I_12895 (I221917,I2683,I221583,I221943,);
nor I_12896 (I221951,I221943,I221810);
DFFARX1 I_12897 (I221951,I2683,I221583,I221551,);
nand I_12898 (I221982,I221943,I221852);
nand I_12899 (I221560,I221835,I221982);
not I_12900 (I222013,I221943);
nor I_12901 (I222030,I222013,I221753);
DFFARX1 I_12902 (I222030,I2683,I221583,I221572,);
nor I_12903 (I222061,I38357,I38342);
or I_12904 (I221563,I221810,I222061);
nor I_12905 (I221554,I221943,I222061);
or I_12906 (I221557,I221677,I222061);
DFFARX1 I_12907 (I222061,I2683,I221583,I221575,);
not I_12908 (I222161,I2690);
DFFARX1 I_12909 (I251877,I2683,I222161,I222187,);
not I_12910 (I222195,I222187);
nand I_12911 (I222212,I251865,I251883);
and I_12912 (I222229,I222212,I251880);
DFFARX1 I_12913 (I222229,I2683,I222161,I222255,);
not I_12914 (I222263,I251871);
DFFARX1 I_12915 (I251868,I2683,I222161,I222289,);
not I_12916 (I222297,I222289);
nor I_12917 (I222314,I222297,I222195);
and I_12918 (I222331,I222314,I251871);
nor I_12919 (I222348,I222297,I222263);
nor I_12920 (I222144,I222255,I222348);
DFFARX1 I_12921 (I251862,I2683,I222161,I222388,);
nor I_12922 (I222396,I222388,I222255);
not I_12923 (I222413,I222396);
not I_12924 (I222430,I222388);
nor I_12925 (I222447,I222430,I222331);
DFFARX1 I_12926 (I222447,I2683,I222161,I222147,);
nand I_12927 (I222478,I251862,I251865);
and I_12928 (I222495,I222478,I251868);
DFFARX1 I_12929 (I222495,I2683,I222161,I222521,);
nor I_12930 (I222529,I222521,I222388);
DFFARX1 I_12931 (I222529,I2683,I222161,I222129,);
nand I_12932 (I222560,I222521,I222430);
nand I_12933 (I222138,I222413,I222560);
not I_12934 (I222591,I222521);
nor I_12935 (I222608,I222591,I222331);
DFFARX1 I_12936 (I222608,I2683,I222161,I222150,);
nor I_12937 (I222639,I251874,I251865);
or I_12938 (I222141,I222388,I222639);
nor I_12939 (I222132,I222521,I222639);
or I_12940 (I222135,I222255,I222639);
DFFARX1 I_12941 (I222639,I2683,I222161,I222153,);
not I_12942 (I222739,I2690);
DFFARX1 I_12943 (I132344,I2683,I222739,I222765,);
not I_12944 (I222773,I222765);
nand I_12945 (I222790,I132335,I132353);
and I_12946 (I222807,I222790,I132356);
DFFARX1 I_12947 (I222807,I2683,I222739,I222833,);
not I_12948 (I222841,I132350);
DFFARX1 I_12949 (I132338,I2683,I222739,I222867,);
not I_12950 (I222875,I222867);
nor I_12951 (I222892,I222875,I222773);
and I_12952 (I222909,I222892,I132350);
nor I_12953 (I222926,I222875,I222841);
nor I_12954 (I222722,I222833,I222926);
DFFARX1 I_12955 (I132347,I2683,I222739,I222966,);
nor I_12956 (I222974,I222966,I222833);
not I_12957 (I222991,I222974);
not I_12958 (I223008,I222966);
nor I_12959 (I223025,I223008,I222909);
DFFARX1 I_12960 (I223025,I2683,I222739,I222725,);
nand I_12961 (I223056,I132362,I132359);
and I_12962 (I223073,I223056,I132341);
DFFARX1 I_12963 (I223073,I2683,I222739,I223099,);
nor I_12964 (I223107,I223099,I222966);
DFFARX1 I_12965 (I223107,I2683,I222739,I222707,);
nand I_12966 (I223138,I223099,I223008);
nand I_12967 (I222716,I222991,I223138);
not I_12968 (I223169,I223099);
nor I_12969 (I223186,I223169,I222909);
DFFARX1 I_12970 (I223186,I2683,I222739,I222728,);
nor I_12971 (I223217,I132335,I132359);
or I_12972 (I222719,I222966,I223217);
nor I_12973 (I222710,I223099,I223217);
or I_12974 (I222713,I222833,I223217);
DFFARX1 I_12975 (I223217,I2683,I222739,I222731,);
not I_12976 (I223317,I2690);
DFFARX1 I_12977 (I138872,I2683,I223317,I223343,);
not I_12978 (I223351,I223343);
nand I_12979 (I223368,I138863,I138881);
and I_12980 (I223385,I223368,I138884);
DFFARX1 I_12981 (I223385,I2683,I223317,I223411,);
not I_12982 (I223419,I138878);
DFFARX1 I_12983 (I138866,I2683,I223317,I223445,);
not I_12984 (I223453,I223445);
nor I_12985 (I223470,I223453,I223351);
and I_12986 (I223487,I223470,I138878);
nor I_12987 (I223504,I223453,I223419);
nor I_12988 (I223300,I223411,I223504);
DFFARX1 I_12989 (I138875,I2683,I223317,I223544,);
nor I_12990 (I223552,I223544,I223411);
not I_12991 (I223569,I223552);
not I_12992 (I223586,I223544);
nor I_12993 (I223603,I223586,I223487);
DFFARX1 I_12994 (I223603,I2683,I223317,I223303,);
nand I_12995 (I223634,I138890,I138887);
and I_12996 (I223651,I223634,I138869);
DFFARX1 I_12997 (I223651,I2683,I223317,I223677,);
nor I_12998 (I223685,I223677,I223544);
DFFARX1 I_12999 (I223685,I2683,I223317,I223285,);
nand I_13000 (I223716,I223677,I223586);
nand I_13001 (I223294,I223569,I223716);
not I_13002 (I223747,I223677);
nor I_13003 (I223764,I223747,I223487);
DFFARX1 I_13004 (I223764,I2683,I223317,I223306,);
nor I_13005 (I223795,I138863,I138887);
or I_13006 (I223297,I223544,I223795);
nor I_13007 (I223288,I223677,I223795);
or I_13008 (I223291,I223411,I223795);
DFFARX1 I_13009 (I223795,I2683,I223317,I223309,);
not I_13010 (I223895,I2690);
DFFARX1 I_13011 (I288538,I2683,I223895,I223921,);
not I_13012 (I223929,I223921);
nand I_13013 (I223946,I288514,I288529);
and I_13014 (I223963,I223946,I288541);
DFFARX1 I_13015 (I223963,I2683,I223895,I223989,);
not I_13016 (I223997,I288526);
DFFARX1 I_13017 (I288517,I2683,I223895,I224023,);
not I_13018 (I224031,I224023);
nor I_13019 (I224048,I224031,I223929);
and I_13020 (I224065,I224048,I288526);
nor I_13021 (I224082,I224031,I223997);
nor I_13022 (I223878,I223989,I224082);
DFFARX1 I_13023 (I288514,I2683,I223895,I224122,);
nor I_13024 (I224130,I224122,I223989);
not I_13025 (I224147,I224130);
not I_13026 (I224164,I224122);
nor I_13027 (I224181,I224164,I224065);
DFFARX1 I_13028 (I224181,I2683,I223895,I223881,);
nand I_13029 (I224212,I288532,I288523);
and I_13030 (I224229,I224212,I288535);
DFFARX1 I_13031 (I224229,I2683,I223895,I224255,);
nor I_13032 (I224263,I224255,I224122);
DFFARX1 I_13033 (I224263,I2683,I223895,I223863,);
nand I_13034 (I224294,I224255,I224164);
nand I_13035 (I223872,I224147,I224294);
not I_13036 (I224325,I224255);
nor I_13037 (I224342,I224325,I224065);
DFFARX1 I_13038 (I224342,I2683,I223895,I223884,);
nor I_13039 (I224373,I288520,I288523);
or I_13040 (I223875,I224122,I224373);
nor I_13041 (I223866,I224255,I224373);
or I_13042 (I223869,I223989,I224373);
DFFARX1 I_13043 (I224373,I2683,I223895,I223887,);
not I_13044 (I224473,I2690);
DFFARX1 I_13045 (I186871,I2683,I224473,I224499,);
not I_13046 (I224507,I224499);
nand I_13047 (I224524,I186880,I186889);
and I_13048 (I224541,I224524,I186895);
DFFARX1 I_13049 (I224541,I2683,I224473,I224567,);
not I_13050 (I224575,I186892);
DFFARX1 I_13051 (I186877,I2683,I224473,I224601,);
not I_13052 (I224609,I224601);
nor I_13053 (I224626,I224609,I224507);
and I_13054 (I224643,I224626,I186892);
nor I_13055 (I224660,I224609,I224575);
nor I_13056 (I224456,I224567,I224660);
DFFARX1 I_13057 (I186886,I2683,I224473,I224700,);
nor I_13058 (I224708,I224700,I224567);
not I_13059 (I224725,I224708);
not I_13060 (I224742,I224700);
nor I_13061 (I224759,I224742,I224643);
DFFARX1 I_13062 (I224759,I2683,I224473,I224459,);
nand I_13063 (I224790,I186883,I186874);
and I_13064 (I224807,I224790,I186871);
DFFARX1 I_13065 (I224807,I2683,I224473,I224833,);
nor I_13066 (I224841,I224833,I224700);
DFFARX1 I_13067 (I224841,I2683,I224473,I224441,);
nand I_13068 (I224872,I224833,I224742);
nand I_13069 (I224450,I224725,I224872);
not I_13070 (I224903,I224833);
nor I_13071 (I224920,I224903,I224643);
DFFARX1 I_13072 (I224920,I2683,I224473,I224462,);
nor I_13073 (I224951,I186874,I186874);
or I_13074 (I224453,I224700,I224951);
nor I_13075 (I224444,I224833,I224951);
or I_13076 (I224447,I224567,I224951);
DFFARX1 I_13077 (I224951,I2683,I224473,I224465,);
not I_13078 (I225051,I2690);
DFFARX1 I_13079 (I35710,I2683,I225051,I225077,);
not I_13080 (I225085,I225077);
nand I_13081 (I225102,I35719,I35728);
and I_13082 (I225119,I225102,I35707);
DFFARX1 I_13083 (I225119,I2683,I225051,I225145,);
not I_13084 (I225153,I35710);
DFFARX1 I_13085 (I35725,I2683,I225051,I225179,);
not I_13086 (I225187,I225179);
nor I_13087 (I225204,I225187,I225085);
and I_13088 (I225221,I225204,I35710);
nor I_13089 (I225238,I225187,I225153);
nor I_13090 (I225034,I225145,I225238);
DFFARX1 I_13091 (I35716,I2683,I225051,I225278,);
nor I_13092 (I225286,I225278,I225145);
not I_13093 (I225303,I225286);
not I_13094 (I225320,I225278);
nor I_13095 (I225337,I225320,I225221);
DFFARX1 I_13096 (I225337,I2683,I225051,I225037,);
nand I_13097 (I225368,I35731,I35707);
and I_13098 (I225385,I225368,I35713);
DFFARX1 I_13099 (I225385,I2683,I225051,I225411,);
nor I_13100 (I225419,I225411,I225278);
DFFARX1 I_13101 (I225419,I2683,I225051,I225019,);
nand I_13102 (I225450,I225411,I225320);
nand I_13103 (I225028,I225303,I225450);
not I_13104 (I225481,I225411);
nor I_13105 (I225498,I225481,I225221);
DFFARX1 I_13106 (I225498,I2683,I225051,I225040,);
nor I_13107 (I225529,I35722,I35707);
or I_13108 (I225031,I225278,I225529);
nor I_13109 (I225022,I225411,I225529);
or I_13110 (I225025,I225145,I225529);
DFFARX1 I_13111 (I225529,I2683,I225051,I225043,);
not I_13112 (I225629,I2690);
DFFARX1 I_13113 (I276264,I2683,I225629,I225655,);
not I_13114 (I225663,I225655);
nand I_13115 (I225680,I276240,I276255);
and I_13116 (I225697,I225680,I276267);
DFFARX1 I_13117 (I225697,I2683,I225629,I225723,);
not I_13118 (I225731,I276252);
DFFARX1 I_13119 (I276243,I2683,I225629,I225757,);
not I_13120 (I225765,I225757);
nor I_13121 (I225782,I225765,I225663);
and I_13122 (I225799,I225782,I276252);
nor I_13123 (I225816,I225765,I225731);
nor I_13124 (I225612,I225723,I225816);
DFFARX1 I_13125 (I276240,I2683,I225629,I225856,);
nor I_13126 (I225864,I225856,I225723);
not I_13127 (I225881,I225864);
not I_13128 (I225898,I225856);
nor I_13129 (I225915,I225898,I225799);
DFFARX1 I_13130 (I225915,I2683,I225629,I225615,);
nand I_13131 (I225946,I276258,I276249);
and I_13132 (I225963,I225946,I276261);
DFFARX1 I_13133 (I225963,I2683,I225629,I225989,);
nor I_13134 (I225997,I225989,I225856);
DFFARX1 I_13135 (I225997,I2683,I225629,I225597,);
nand I_13136 (I226028,I225989,I225898);
nand I_13137 (I225606,I225881,I226028);
not I_13138 (I226059,I225989);
nor I_13139 (I226076,I226059,I225799);
DFFARX1 I_13140 (I226076,I2683,I225629,I225618,);
nor I_13141 (I226107,I276246,I276249);
or I_13142 (I225609,I225856,I226107);
nor I_13143 (I225600,I225989,I226107);
or I_13144 (I225603,I225723,I226107);
DFFARX1 I_13145 (I226107,I2683,I225629,I225621,);
not I_13146 (I226207,I2690);
DFFARX1 I_13147 (I2348,I2683,I226207,I226233,);
not I_13148 (I226241,I226233);
nand I_13149 (I226258,I2372,I1996);
and I_13150 (I226275,I226258,I1884);
DFFARX1 I_13151 (I226275,I2683,I226207,I226301,);
not I_13152 (I226309,I2668);
DFFARX1 I_13153 (I1540,I2683,I226207,I226335,);
not I_13154 (I226343,I226335);
nor I_13155 (I226360,I226343,I226241);
and I_13156 (I226377,I226360,I2668);
nor I_13157 (I226394,I226343,I226309);
nor I_13158 (I226190,I226301,I226394);
DFFARX1 I_13159 (I2068,I2683,I226207,I226434,);
nor I_13160 (I226442,I226434,I226301);
not I_13161 (I226459,I226442);
not I_13162 (I226476,I226434);
nor I_13163 (I226493,I226476,I226377);
DFFARX1 I_13164 (I226493,I2683,I226207,I226193,);
nand I_13165 (I226524,I2100,I2236);
and I_13166 (I226541,I226524,I2428);
DFFARX1 I_13167 (I226541,I2683,I226207,I226567,);
nor I_13168 (I226575,I226567,I226434);
DFFARX1 I_13169 (I226575,I2683,I226207,I226175,);
nand I_13170 (I226606,I226567,I226476);
nand I_13171 (I226184,I226459,I226606);
not I_13172 (I226637,I226567);
nor I_13173 (I226654,I226637,I226377);
DFFARX1 I_13174 (I226654,I2683,I226207,I226196,);
nor I_13175 (I226685,I2604,I2236);
or I_13176 (I226187,I226434,I226685);
nor I_13177 (I226178,I226567,I226685);
or I_13178 (I226181,I226301,I226685);
DFFARX1 I_13179 (I226685,I2683,I226207,I226199,);
not I_13180 (I226785,I2690);
DFFARX1 I_13181 (I239756,I2683,I226785,I226811,);
not I_13182 (I226819,I226811);
nand I_13183 (I226836,I239744,I239762);
and I_13184 (I226853,I226836,I239759);
DFFARX1 I_13185 (I226853,I2683,I226785,I226879,);
not I_13186 (I226887,I239750);
DFFARX1 I_13187 (I239747,I2683,I226785,I226913,);
not I_13188 (I226921,I226913);
nor I_13189 (I226938,I226921,I226819);
and I_13190 (I226955,I226938,I239750);
nor I_13191 (I226972,I226921,I226887);
nor I_13192 (I226768,I226879,I226972);
DFFARX1 I_13193 (I239741,I2683,I226785,I227012,);
nor I_13194 (I227020,I227012,I226879);
not I_13195 (I227037,I227020);
not I_13196 (I227054,I227012);
nor I_13197 (I227071,I227054,I226955);
DFFARX1 I_13198 (I227071,I2683,I226785,I226771,);
nand I_13199 (I227102,I239741,I239744);
and I_13200 (I227119,I227102,I239747);
DFFARX1 I_13201 (I227119,I2683,I226785,I227145,);
nor I_13202 (I227153,I227145,I227012);
DFFARX1 I_13203 (I227153,I2683,I226785,I226753,);
nand I_13204 (I227184,I227145,I227054);
nand I_13205 (I226762,I227037,I227184);
not I_13206 (I227215,I227145);
nor I_13207 (I227232,I227215,I226955);
DFFARX1 I_13208 (I227232,I2683,I226785,I226774,);
nor I_13209 (I227263,I239753,I239744);
or I_13210 (I226765,I227012,I227263);
nor I_13211 (I226756,I227145,I227263);
or I_13212 (I226759,I226879,I227263);
DFFARX1 I_13213 (I227263,I2683,I226785,I226777,);
not I_13214 (I227363,I2690);
DFFARX1 I_13215 (I280140,I2683,I227363,I227389,);
not I_13216 (I227397,I227389);
nand I_13217 (I227414,I280116,I280131);
and I_13218 (I227431,I227414,I280143);
DFFARX1 I_13219 (I227431,I2683,I227363,I227457,);
not I_13220 (I227465,I280128);
DFFARX1 I_13221 (I280119,I2683,I227363,I227491,);
not I_13222 (I227499,I227491);
nor I_13223 (I227516,I227499,I227397);
and I_13224 (I227533,I227516,I280128);
nor I_13225 (I227550,I227499,I227465);
nor I_13226 (I227346,I227457,I227550);
DFFARX1 I_13227 (I280116,I2683,I227363,I227590,);
nor I_13228 (I227598,I227590,I227457);
not I_13229 (I227615,I227598);
not I_13230 (I227632,I227590);
nor I_13231 (I227649,I227632,I227533);
DFFARX1 I_13232 (I227649,I2683,I227363,I227349,);
nand I_13233 (I227680,I280134,I280125);
and I_13234 (I227697,I227680,I280137);
DFFARX1 I_13235 (I227697,I2683,I227363,I227723,);
nor I_13236 (I227731,I227723,I227590);
DFFARX1 I_13237 (I227731,I2683,I227363,I227331,);
nand I_13238 (I227762,I227723,I227632);
nand I_13239 (I227340,I227615,I227762);
not I_13240 (I227793,I227723);
nor I_13241 (I227810,I227793,I227533);
DFFARX1 I_13242 (I227810,I2683,I227363,I227352,);
nor I_13243 (I227841,I280122,I280125);
or I_13244 (I227343,I227590,I227841);
nor I_13245 (I227334,I227723,I227841);
or I_13246 (I227337,I227457,I227841);
DFFARX1 I_13247 (I227841,I2683,I227363,I227355,);
not I_13248 (I227941,I2690);
DFFARX1 I_13249 (I256093,I2683,I227941,I227967,);
not I_13250 (I227975,I227967);
nand I_13251 (I227992,I256081,I256099);
and I_13252 (I228009,I227992,I256096);
DFFARX1 I_13253 (I228009,I2683,I227941,I228035,);
not I_13254 (I228043,I256087);
DFFARX1 I_13255 (I256084,I2683,I227941,I228069,);
not I_13256 (I228077,I228069);
nor I_13257 (I228094,I228077,I227975);
and I_13258 (I228111,I228094,I256087);
nor I_13259 (I228128,I228077,I228043);
nor I_13260 (I227924,I228035,I228128);
DFFARX1 I_13261 (I256078,I2683,I227941,I228168,);
nor I_13262 (I228176,I228168,I228035);
not I_13263 (I228193,I228176);
not I_13264 (I228210,I228168);
nor I_13265 (I228227,I228210,I228111);
DFFARX1 I_13266 (I228227,I2683,I227941,I227927,);
nand I_13267 (I228258,I256078,I256081);
and I_13268 (I228275,I228258,I256084);
DFFARX1 I_13269 (I228275,I2683,I227941,I228301,);
nor I_13270 (I228309,I228301,I228168);
DFFARX1 I_13271 (I228309,I2683,I227941,I227909,);
nand I_13272 (I228340,I228301,I228210);
nand I_13273 (I227918,I228193,I228340);
not I_13274 (I228371,I228301);
nor I_13275 (I228388,I228371,I228111);
DFFARX1 I_13276 (I228388,I2683,I227941,I227930,);
nor I_13277 (I228419,I256090,I256081);
or I_13278 (I227921,I228168,I228419);
nor I_13279 (I227912,I228301,I228419);
or I_13280 (I227915,I228035,I228419);
DFFARX1 I_13281 (I228419,I2683,I227941,I227933,);
not I_13282 (I228519,I2690);
DFFARX1 I_13283 (I236594,I2683,I228519,I228545,);
not I_13284 (I228553,I228545);
nand I_13285 (I228570,I236582,I236600);
and I_13286 (I228587,I228570,I236597);
DFFARX1 I_13287 (I228587,I2683,I228519,I228613,);
not I_13288 (I228621,I236588);
DFFARX1 I_13289 (I236585,I2683,I228519,I228647,);
not I_13290 (I228655,I228647);
nor I_13291 (I228672,I228655,I228553);
and I_13292 (I228689,I228672,I236588);
nor I_13293 (I228706,I228655,I228621);
nor I_13294 (I228502,I228613,I228706);
DFFARX1 I_13295 (I236579,I2683,I228519,I228746,);
nor I_13296 (I228754,I228746,I228613);
not I_13297 (I228771,I228754);
not I_13298 (I228788,I228746);
nor I_13299 (I228805,I228788,I228689);
DFFARX1 I_13300 (I228805,I2683,I228519,I228505,);
nand I_13301 (I228836,I236579,I236582);
and I_13302 (I228853,I228836,I236585);
DFFARX1 I_13303 (I228853,I2683,I228519,I228879,);
nor I_13304 (I228887,I228879,I228746);
DFFARX1 I_13305 (I228887,I2683,I228519,I228487,);
nand I_13306 (I228918,I228879,I228788);
nand I_13307 (I228496,I228771,I228918);
not I_13308 (I228949,I228879);
nor I_13309 (I228966,I228949,I228689);
DFFARX1 I_13310 (I228966,I2683,I228519,I228508,);
nor I_13311 (I228997,I236591,I236582);
or I_13312 (I228499,I228746,I228997);
nor I_13313 (I228490,I228879,I228997);
or I_13314 (I228493,I228613,I228997);
DFFARX1 I_13315 (I228997,I2683,I228519,I228511,);
not I_13316 (I229097,I2690);
DFFARX1 I_13317 (I2012,I2683,I229097,I229123,);
not I_13318 (I229131,I229123);
nand I_13319 (I229148,I1796,I1364);
and I_13320 (I229165,I229148,I1460);
DFFARX1 I_13321 (I229165,I2683,I229097,I229191,);
not I_13322 (I229199,I2116);
DFFARX1 I_13323 (I1844,I2683,I229097,I229225,);
not I_13324 (I229233,I229225);
nor I_13325 (I229250,I229233,I229131);
and I_13326 (I229267,I229250,I2116);
nor I_13327 (I229284,I229233,I229199);
nor I_13328 (I229080,I229191,I229284);
DFFARX1 I_13329 (I2620,I2683,I229097,I229324,);
nor I_13330 (I229332,I229324,I229191);
not I_13331 (I229349,I229332);
not I_13332 (I229366,I229324);
nor I_13333 (I229383,I229366,I229267);
DFFARX1 I_13334 (I229383,I2683,I229097,I229083,);
nand I_13335 (I229414,I2396,I2124);
and I_13336 (I229431,I229414,I2548);
DFFARX1 I_13337 (I229431,I2683,I229097,I229457,);
nor I_13338 (I229465,I229457,I229324);
DFFARX1 I_13339 (I229465,I2683,I229097,I229065,);
nand I_13340 (I229496,I229457,I229366);
nand I_13341 (I229074,I229349,I229496);
not I_13342 (I229527,I229457);
nor I_13343 (I229544,I229527,I229267);
DFFARX1 I_13344 (I229544,I2683,I229097,I229086,);
nor I_13345 (I229575,I2180,I2124);
or I_13346 (I229077,I229324,I229575);
nor I_13347 (I229068,I229457,I229575);
or I_13348 (I229071,I229191,I229575);
DFFARX1 I_13349 (I229575,I2683,I229097,I229089,);
not I_13350 (I229675,I2690);
DFFARX1 I_13351 (I416466,I2683,I229675,I229701,);
not I_13352 (I229709,I229701);
nand I_13353 (I229726,I416451,I416439);
and I_13354 (I229743,I229726,I416454);
DFFARX1 I_13355 (I229743,I2683,I229675,I229769,);
not I_13356 (I229777,I416439);
DFFARX1 I_13357 (I416457,I2683,I229675,I229803,);
not I_13358 (I229811,I229803);
nor I_13359 (I229828,I229811,I229709);
and I_13360 (I229845,I229828,I416439);
nor I_13361 (I229862,I229811,I229777);
nor I_13362 (I229658,I229769,I229862);
DFFARX1 I_13363 (I416445,I2683,I229675,I229902,);
nor I_13364 (I229910,I229902,I229769);
not I_13365 (I229927,I229910);
not I_13366 (I229944,I229902);
nor I_13367 (I229961,I229944,I229845);
DFFARX1 I_13368 (I229961,I2683,I229675,I229661,);
nand I_13369 (I229992,I416442,I416448);
and I_13370 (I230009,I229992,I416463);
DFFARX1 I_13371 (I230009,I2683,I229675,I230035,);
nor I_13372 (I230043,I230035,I229902);
DFFARX1 I_13373 (I230043,I2683,I229675,I229643,);
nand I_13374 (I230074,I230035,I229944);
nand I_13375 (I229652,I229927,I230074);
not I_13376 (I230105,I230035);
nor I_13377 (I230122,I230105,I229845);
DFFARX1 I_13378 (I230122,I2683,I229675,I229664,);
nor I_13379 (I230153,I416460,I416448);
or I_13380 (I229655,I229902,I230153);
nor I_13381 (I229646,I230035,I230153);
or I_13382 (I229649,I229769,I230153);
DFFARX1 I_13383 (I230153,I2683,I229675,I229667,);
not I_13384 (I230253,I2690);
DFFARX1 I_13385 (I79839,I2683,I230253,I230279,);
not I_13386 (I230287,I230279);
nand I_13387 (I230304,I79842,I79863);
and I_13388 (I230321,I230304,I79851);
DFFARX1 I_13389 (I230321,I2683,I230253,I230347,);
not I_13390 (I230355,I79848);
DFFARX1 I_13391 (I79839,I2683,I230253,I230381,);
not I_13392 (I230389,I230381);
nor I_13393 (I230406,I230389,I230287);
and I_13394 (I230423,I230406,I79848);
nor I_13395 (I230440,I230389,I230355);
nor I_13396 (I230236,I230347,I230440);
DFFARX1 I_13397 (I79857,I2683,I230253,I230480,);
nor I_13398 (I230488,I230480,I230347);
not I_13399 (I230505,I230488);
not I_13400 (I230522,I230480);
nor I_13401 (I230539,I230522,I230423);
DFFARX1 I_13402 (I230539,I2683,I230253,I230239,);
nand I_13403 (I230570,I79842,I79845);
and I_13404 (I230587,I230570,I79854);
DFFARX1 I_13405 (I230587,I2683,I230253,I230613,);
nor I_13406 (I230621,I230613,I230480);
DFFARX1 I_13407 (I230621,I2683,I230253,I230221,);
nand I_13408 (I230652,I230613,I230522);
nand I_13409 (I230230,I230505,I230652);
not I_13410 (I230683,I230613);
nor I_13411 (I230700,I230683,I230423);
DFFARX1 I_13412 (I230700,I2683,I230253,I230242,);
nor I_13413 (I230731,I79860,I79845);
or I_13414 (I230233,I230480,I230731);
nor I_13415 (I230224,I230613,I230731);
or I_13416 (I230227,I230347,I230731);
DFFARX1 I_13417 (I230731,I2683,I230253,I230245,);
not I_13418 (I230831,I2690);
DFFARX1 I_13419 (I274326,I2683,I230831,I230857,);
not I_13420 (I230865,I230857);
nand I_13421 (I230882,I274302,I274317);
and I_13422 (I230899,I230882,I274329);
DFFARX1 I_13423 (I230899,I2683,I230831,I230925,);
not I_13424 (I230933,I274314);
DFFARX1 I_13425 (I274305,I2683,I230831,I230959,);
not I_13426 (I230967,I230959);
nor I_13427 (I230984,I230967,I230865);
and I_13428 (I231001,I230984,I274314);
nor I_13429 (I231018,I230967,I230933);
nor I_13430 (I230814,I230925,I231018);
DFFARX1 I_13431 (I274302,I2683,I230831,I231058,);
nor I_13432 (I231066,I231058,I230925);
not I_13433 (I231083,I231066);
not I_13434 (I231100,I231058);
nor I_13435 (I231117,I231100,I231001);
DFFARX1 I_13436 (I231117,I2683,I230831,I230817,);
nand I_13437 (I231148,I274320,I274311);
and I_13438 (I231165,I231148,I274323);
DFFARX1 I_13439 (I231165,I2683,I230831,I231191,);
nor I_13440 (I231199,I231191,I231058);
DFFARX1 I_13441 (I231199,I2683,I230831,I230799,);
nand I_13442 (I231230,I231191,I231100);
nand I_13443 (I230808,I231083,I231230);
not I_13444 (I231261,I231191);
nor I_13445 (I231278,I231261,I231001);
DFFARX1 I_13446 (I231278,I2683,I230831,I230820,);
nor I_13447 (I231309,I274308,I274311);
or I_13448 (I230811,I231058,I231309);
nor I_13449 (I230802,I231191,I231309);
or I_13450 (I230805,I230925,I231309);
DFFARX1 I_13451 (I231309,I2683,I230831,I230823,);
not I_13452 (I231409,I2690);
DFFARX1 I_13453 (I22535,I2683,I231409,I231435,);
not I_13454 (I231443,I231435);
nand I_13455 (I231460,I22544,I22553);
and I_13456 (I231477,I231460,I22532);
DFFARX1 I_13457 (I231477,I2683,I231409,I231503,);
not I_13458 (I231511,I22535);
DFFARX1 I_13459 (I22550,I2683,I231409,I231537,);
not I_13460 (I231545,I231537);
nor I_13461 (I231562,I231545,I231443);
and I_13462 (I231579,I231562,I22535);
nor I_13463 (I231596,I231545,I231511);
nor I_13464 (I231392,I231503,I231596);
DFFARX1 I_13465 (I22541,I2683,I231409,I231636,);
nor I_13466 (I231644,I231636,I231503);
not I_13467 (I231661,I231644);
not I_13468 (I231678,I231636);
nor I_13469 (I231695,I231678,I231579);
DFFARX1 I_13470 (I231695,I2683,I231409,I231395,);
nand I_13471 (I231726,I22556,I22532);
and I_13472 (I231743,I231726,I22538);
DFFARX1 I_13473 (I231743,I2683,I231409,I231769,);
nor I_13474 (I231777,I231769,I231636);
DFFARX1 I_13475 (I231777,I2683,I231409,I231377,);
nand I_13476 (I231808,I231769,I231678);
nand I_13477 (I231386,I231661,I231808);
not I_13478 (I231839,I231769);
nor I_13479 (I231856,I231839,I231579);
DFFARX1 I_13480 (I231856,I2683,I231409,I231398,);
nor I_13481 (I231887,I22547,I22532);
or I_13482 (I231389,I231636,I231887);
nor I_13483 (I231380,I231769,I231887);
or I_13484 (I231383,I231503,I231887);
DFFARX1 I_13485 (I231887,I2683,I231409,I231401,);
not I_13486 (I231987,I2690);
DFFARX1 I_13487 (I394014,I2683,I231987,I232013,);
not I_13488 (I232021,I232013);
nand I_13489 (I232038,I394002,I394020);
and I_13490 (I232055,I232038,I394011);
DFFARX1 I_13491 (I232055,I2683,I231987,I232081,);
not I_13492 (I232089,I394026);
DFFARX1 I_13493 (I394023,I2683,I231987,I232115,);
not I_13494 (I232123,I232115);
nor I_13495 (I232140,I232123,I232021);
and I_13496 (I232157,I232140,I394026);
nor I_13497 (I232174,I232123,I232089);
nor I_13498 (I231970,I232081,I232174);
DFFARX1 I_13499 (I394005,I2683,I231987,I232214,);
nor I_13500 (I232222,I232214,I232081);
not I_13501 (I232239,I232222);
not I_13502 (I232256,I232214);
nor I_13503 (I232273,I232256,I232157);
DFFARX1 I_13504 (I232273,I2683,I231987,I231973,);
nand I_13505 (I232304,I393999,I393999);
and I_13506 (I232321,I232304,I394008);
DFFARX1 I_13507 (I232321,I2683,I231987,I232347,);
nor I_13508 (I232355,I232347,I232214);
DFFARX1 I_13509 (I232355,I2683,I231987,I231955,);
nand I_13510 (I232386,I232347,I232256);
nand I_13511 (I231964,I232239,I232386);
not I_13512 (I232417,I232347);
nor I_13513 (I232434,I232417,I232157);
DFFARX1 I_13514 (I232434,I2683,I231987,I231976,);
nor I_13515 (I232465,I394017,I393999);
or I_13516 (I231967,I232214,I232465);
nor I_13517 (I231958,I232347,I232465);
or I_13518 (I231961,I232081,I232465);
DFFARX1 I_13519 (I232465,I2683,I231987,I231979,);
not I_13520 (I232565,I2690);
DFFARX1 I_13521 (I5079,I2683,I232565,I232591,);
not I_13522 (I232599,I232591);
nand I_13523 (I232616,I5082,I5094);
and I_13524 (I232633,I232616,I5073);
DFFARX1 I_13525 (I232633,I2683,I232565,I232659,);
not I_13526 (I232667,I5073);
DFFARX1 I_13527 (I5076,I2683,I232565,I232693,);
not I_13528 (I232701,I232693);
nor I_13529 (I232718,I232701,I232599);
and I_13530 (I232735,I232718,I5073);
nor I_13531 (I232752,I232701,I232667);
nor I_13532 (I232548,I232659,I232752);
DFFARX1 I_13533 (I5088,I2683,I232565,I232792,);
nor I_13534 (I232800,I232792,I232659);
not I_13535 (I232817,I232800);
not I_13536 (I232834,I232792);
nor I_13537 (I232851,I232834,I232735);
DFFARX1 I_13538 (I232851,I2683,I232565,I232551,);
nand I_13539 (I232882,I5091,I5076);
and I_13540 (I232899,I232882,I5085);
DFFARX1 I_13541 (I232899,I2683,I232565,I232925,);
nor I_13542 (I232933,I232925,I232792);
DFFARX1 I_13543 (I232933,I2683,I232565,I232533,);
nand I_13544 (I232964,I232925,I232834);
nand I_13545 (I232542,I232817,I232964);
not I_13546 (I232995,I232925);
nor I_13547 (I233012,I232995,I232735);
DFFARX1 I_13548 (I233012,I2683,I232565,I232554,);
nor I_13549 (I233043,I5079,I5076);
or I_13550 (I232545,I232792,I233043);
nor I_13551 (I232536,I232925,I233043);
or I_13552 (I232539,I232659,I233043);
DFFARX1 I_13553 (I233043,I2683,I232565,I232557,);
not I_13554 (I233143,I2690);
DFFARX1 I_13555 (I24643,I2683,I233143,I233169,);
not I_13556 (I233177,I233169);
nand I_13557 (I233194,I24652,I24661);
and I_13558 (I233211,I233194,I24640);
DFFARX1 I_13559 (I233211,I2683,I233143,I233237,);
not I_13560 (I233245,I24643);
DFFARX1 I_13561 (I24658,I2683,I233143,I233271,);
not I_13562 (I233279,I233271);
nor I_13563 (I233296,I233279,I233177);
and I_13564 (I233313,I233296,I24643);
nor I_13565 (I233330,I233279,I233245);
nor I_13566 (I233126,I233237,I233330);
DFFARX1 I_13567 (I24649,I2683,I233143,I233370,);
nor I_13568 (I233378,I233370,I233237);
not I_13569 (I233395,I233378);
not I_13570 (I233412,I233370);
nor I_13571 (I233429,I233412,I233313);
DFFARX1 I_13572 (I233429,I2683,I233143,I233129,);
nand I_13573 (I233460,I24664,I24640);
and I_13574 (I233477,I233460,I24646);
DFFARX1 I_13575 (I233477,I2683,I233143,I233503,);
nor I_13576 (I233511,I233503,I233370);
DFFARX1 I_13577 (I233511,I2683,I233143,I233111,);
nand I_13578 (I233542,I233503,I233412);
nand I_13579 (I233120,I233395,I233542);
not I_13580 (I233573,I233503);
nor I_13581 (I233590,I233573,I233313);
DFFARX1 I_13582 (I233590,I2683,I233143,I233132,);
nor I_13583 (I233621,I24655,I24640);
or I_13584 (I233123,I233370,I233621);
nor I_13585 (I233114,I233503,I233621);
or I_13586 (I233117,I233237,I233621);
DFFARX1 I_13587 (I233621,I2683,I233143,I233135,);
not I_13588 (I233721,I2690);
DFFARX1 I_13589 (I73889,I2683,I233721,I233747,);
not I_13590 (I233755,I233747);
nand I_13591 (I233772,I73892,I73913);
and I_13592 (I233789,I233772,I73901);
DFFARX1 I_13593 (I233789,I2683,I233721,I233815,);
not I_13594 (I233823,I73898);
DFFARX1 I_13595 (I73889,I2683,I233721,I233849,);
not I_13596 (I233857,I233849);
nor I_13597 (I233874,I233857,I233755);
and I_13598 (I233891,I233874,I73898);
nor I_13599 (I233908,I233857,I233823);
nor I_13600 (I233704,I233815,I233908);
DFFARX1 I_13601 (I73907,I2683,I233721,I233948,);
nor I_13602 (I233956,I233948,I233815);
not I_13603 (I233973,I233956);
not I_13604 (I233990,I233948);
nor I_13605 (I234007,I233990,I233891);
DFFARX1 I_13606 (I234007,I2683,I233721,I233707,);
nand I_13607 (I234038,I73892,I73895);
and I_13608 (I234055,I234038,I73904);
DFFARX1 I_13609 (I234055,I2683,I233721,I234081,);
nor I_13610 (I234089,I234081,I233948);
DFFARX1 I_13611 (I234089,I2683,I233721,I233689,);
nand I_13612 (I234120,I234081,I233990);
nand I_13613 (I233698,I233973,I234120);
not I_13614 (I234151,I234081);
nor I_13615 (I234168,I234151,I233891);
DFFARX1 I_13616 (I234168,I2683,I233721,I233710,);
nor I_13617 (I234199,I73910,I73895);
or I_13618 (I233701,I233948,I234199);
nor I_13619 (I233692,I234081,I234199);
or I_13620 (I233695,I233815,I234199);
DFFARX1 I_13621 (I234199,I2683,I233721,I233713,);
not I_13622 (I234299,I2690);
DFFARX1 I_13623 (I140504,I2683,I234299,I234325,);
not I_13624 (I234333,I234325);
nand I_13625 (I234350,I140495,I140513);
and I_13626 (I234367,I234350,I140516);
DFFARX1 I_13627 (I234367,I2683,I234299,I234393,);
not I_13628 (I234401,I140510);
DFFARX1 I_13629 (I140498,I2683,I234299,I234427,);
not I_13630 (I234435,I234427);
nor I_13631 (I234452,I234435,I234333);
and I_13632 (I234469,I234452,I140510);
nor I_13633 (I234486,I234435,I234401);
nor I_13634 (I234282,I234393,I234486);
DFFARX1 I_13635 (I140507,I2683,I234299,I234526,);
nor I_13636 (I234534,I234526,I234393);
not I_13637 (I234551,I234534);
not I_13638 (I234568,I234526);
nor I_13639 (I234585,I234568,I234469);
DFFARX1 I_13640 (I234585,I2683,I234299,I234285,);
nand I_13641 (I234616,I140522,I140519);
and I_13642 (I234633,I234616,I140501);
DFFARX1 I_13643 (I234633,I2683,I234299,I234659,);
nor I_13644 (I234667,I234659,I234526);
DFFARX1 I_13645 (I234667,I2683,I234299,I234267,);
nand I_13646 (I234698,I234659,I234568);
nand I_13647 (I234276,I234551,I234698);
not I_13648 (I234729,I234659);
nor I_13649 (I234746,I234729,I234469);
DFFARX1 I_13650 (I234746,I2683,I234299,I234288,);
nor I_13651 (I234777,I140495,I140519);
or I_13652 (I234279,I234526,I234777);
nor I_13653 (I234270,I234659,I234777);
or I_13654 (I234273,I234393,I234777);
DFFARX1 I_13655 (I234777,I2683,I234299,I234291,);
not I_13656 (I234877,I2690);
DFFARX1 I_13657 (I175889,I2683,I234877,I234903,);
not I_13658 (I234911,I234903);
nand I_13659 (I234928,I175898,I175907);
and I_13660 (I234945,I234928,I175913);
DFFARX1 I_13661 (I234945,I2683,I234877,I234971,);
not I_13662 (I234979,I175910);
DFFARX1 I_13663 (I175895,I2683,I234877,I235005,);
not I_13664 (I235013,I235005);
nor I_13665 (I235030,I235013,I234911);
and I_13666 (I235047,I235030,I175910);
nor I_13667 (I235064,I235013,I234979);
nor I_13668 (I234860,I234971,I235064);
DFFARX1 I_13669 (I175904,I2683,I234877,I235104,);
nor I_13670 (I235112,I235104,I234971);
not I_13671 (I235129,I235112);
not I_13672 (I235146,I235104);
nor I_13673 (I235163,I235146,I235047);
DFFARX1 I_13674 (I235163,I2683,I234877,I234863,);
nand I_13675 (I235194,I175901,I175892);
and I_13676 (I235211,I235194,I175889);
DFFARX1 I_13677 (I235211,I2683,I234877,I235237,);
nor I_13678 (I235245,I235237,I235104);
DFFARX1 I_13679 (I235245,I2683,I234877,I234845,);
nand I_13680 (I235276,I235237,I235146);
nand I_13681 (I234854,I235129,I235276);
not I_13682 (I235307,I235237);
nor I_13683 (I235324,I235307,I235047);
DFFARX1 I_13684 (I235324,I2683,I234877,I234866,);
nor I_13685 (I235355,I175892,I175892);
or I_13686 (I234857,I235104,I235355);
nor I_13687 (I234848,I235237,I235355);
or I_13688 (I234851,I234971,I235355);
DFFARX1 I_13689 (I235355,I2683,I234877,I234869,);
not I_13690 (I235455,I2690);
DFFARX1 I_13691 (I187449,I2683,I235455,I235481,);
not I_13692 (I235489,I235481);
nand I_13693 (I235506,I187458,I187467);
and I_13694 (I235523,I235506,I187473);
DFFARX1 I_13695 (I235523,I2683,I235455,I235549,);
not I_13696 (I235557,I187470);
DFFARX1 I_13697 (I187455,I2683,I235455,I235583,);
not I_13698 (I235591,I235583);
nor I_13699 (I235608,I235591,I235489);
and I_13700 (I235625,I235608,I187470);
nor I_13701 (I235642,I235591,I235557);
nor I_13702 (I235438,I235549,I235642);
DFFARX1 I_13703 (I187464,I2683,I235455,I235682,);
nor I_13704 (I235690,I235682,I235549);
not I_13705 (I235707,I235690);
not I_13706 (I235724,I235682);
nor I_13707 (I235741,I235724,I235625);
DFFARX1 I_13708 (I235741,I2683,I235455,I235441,);
nand I_13709 (I235772,I187461,I187452);
and I_13710 (I235789,I235772,I187449);
DFFARX1 I_13711 (I235789,I2683,I235455,I235815,);
nor I_13712 (I235823,I235815,I235682);
DFFARX1 I_13713 (I235823,I2683,I235455,I235423,);
nand I_13714 (I235854,I235815,I235724);
nand I_13715 (I235432,I235707,I235854);
not I_13716 (I235885,I235815);
nor I_13717 (I235902,I235885,I235625);
DFFARX1 I_13718 (I235902,I2683,I235455,I235444,);
nor I_13719 (I235933,I187452,I187452);
or I_13720 (I235435,I235682,I235933);
nor I_13721 (I235426,I235815,I235933);
or I_13722 (I235429,I235549,I235933);
DFFARX1 I_13723 (I235933,I2683,I235455,I235447,);
not I_13724 (I236033,I2690);
DFFARX1 I_13725 (I21481,I2683,I236033,I236059,);
not I_13726 (I236067,I236059);
nand I_13727 (I236084,I21490,I21499);
and I_13728 (I236101,I236084,I21478);
DFFARX1 I_13729 (I236101,I2683,I236033,I236127,);
not I_13730 (I236135,I21481);
DFFARX1 I_13731 (I21496,I2683,I236033,I236161,);
not I_13732 (I236169,I236161);
nor I_13733 (I236186,I236169,I236067);
and I_13734 (I236203,I236186,I21481);
nor I_13735 (I236220,I236169,I236135);
nor I_13736 (I236016,I236127,I236220);
DFFARX1 I_13737 (I21487,I2683,I236033,I236260,);
nor I_13738 (I236268,I236260,I236127);
not I_13739 (I236285,I236268);
not I_13740 (I236302,I236260);
nor I_13741 (I236319,I236302,I236203);
DFFARX1 I_13742 (I236319,I2683,I236033,I236019,);
nand I_13743 (I236350,I21502,I21478);
and I_13744 (I236367,I236350,I21484);
DFFARX1 I_13745 (I236367,I2683,I236033,I236393,);
nor I_13746 (I236401,I236393,I236260);
DFFARX1 I_13747 (I236401,I2683,I236033,I236001,);
nand I_13748 (I236432,I236393,I236302);
nand I_13749 (I236010,I236285,I236432);
not I_13750 (I236463,I236393);
nor I_13751 (I236480,I236463,I236203);
DFFARX1 I_13752 (I236480,I2683,I236033,I236022,);
nor I_13753 (I236511,I21493,I21478);
or I_13754 (I236013,I236260,I236511);
nor I_13755 (I236004,I236393,I236511);
or I_13756 (I236007,I236127,I236511);
DFFARX1 I_13757 (I236511,I2683,I236033,I236025,);
not I_13758 (I236608,I2690);
DFFARX1 I_13759 (I286579,I2683,I236608,I236634,);
not I_13760 (I236642,I236634);
nand I_13761 (I236659,I286594,I286576);
and I_13762 (I236676,I236659,I286576);
DFFARX1 I_13763 (I236676,I2683,I236608,I236702,);
DFFARX1 I_13764 (I236702,I2683,I236608,I236597,);
DFFARX1 I_13765 (I286585,I2683,I236608,I236733,);
nand I_13766 (I236741,I236733,I286603);
not I_13767 (I236758,I236741);
DFFARX1 I_13768 (I236758,I2683,I236608,I236784,);
not I_13769 (I236792,I236784);
nor I_13770 (I236600,I236642,I236792);
DFFARX1 I_13771 (I286600,I2683,I236608,I236832,);
nor I_13772 (I236591,I236832,I236702);
nor I_13773 (I236582,I236832,I236758);
nand I_13774 (I236868,I286597,I286588);
and I_13775 (I236885,I236868,I286582);
DFFARX1 I_13776 (I236885,I2683,I236608,I236911,);
not I_13777 (I236919,I236911);
nand I_13778 (I236936,I236919,I236832);
nand I_13779 (I236585,I236919,I236741);
nor I_13780 (I236967,I286591,I286588);
and I_13781 (I236984,I236832,I236967);
nor I_13782 (I237001,I236919,I236984);
DFFARX1 I_13783 (I237001,I2683,I236608,I236594,);
nor I_13784 (I237032,I236634,I236967);
DFFARX1 I_13785 (I237032,I2683,I236608,I236579,);
nor I_13786 (I237063,I236911,I236967);
not I_13787 (I237080,I237063);
nand I_13788 (I236588,I237080,I236936);
not I_13789 (I237135,I2690);
DFFARX1 I_13790 (I219239,I2683,I237135,I237161,);
not I_13791 (I237169,I237161);
nand I_13792 (I237186,I219242,I219239);
and I_13793 (I237203,I237186,I219251);
DFFARX1 I_13794 (I237203,I2683,I237135,I237229,);
DFFARX1 I_13795 (I237229,I2683,I237135,I237124,);
DFFARX1 I_13796 (I219248,I2683,I237135,I237260,);
nand I_13797 (I237268,I237260,I219254);
not I_13798 (I237285,I237268);
DFFARX1 I_13799 (I237285,I2683,I237135,I237311,);
not I_13800 (I237319,I237311);
nor I_13801 (I237127,I237169,I237319);
DFFARX1 I_13802 (I219263,I2683,I237135,I237359,);
nor I_13803 (I237118,I237359,I237229);
nor I_13804 (I237109,I237359,I237285);
nand I_13805 (I237395,I219257,I219245);
and I_13806 (I237412,I237395,I219242);
DFFARX1 I_13807 (I237412,I2683,I237135,I237438,);
not I_13808 (I237446,I237438);
nand I_13809 (I237463,I237446,I237359);
nand I_13810 (I237112,I237446,I237268);
nor I_13811 (I237494,I219260,I219245);
and I_13812 (I237511,I237359,I237494);
nor I_13813 (I237528,I237446,I237511);
DFFARX1 I_13814 (I237528,I2683,I237135,I237121,);
nor I_13815 (I237559,I237161,I237494);
DFFARX1 I_13816 (I237559,I2683,I237135,I237106,);
nor I_13817 (I237590,I237438,I237494);
not I_13818 (I237607,I237590);
nand I_13819 (I237115,I237607,I237463);
not I_13820 (I237662,I2690);
DFFARX1 I_13821 (I28353,I2683,I237662,I237688,);
not I_13822 (I237696,I237688);
nand I_13823 (I237713,I28329,I28338);
and I_13824 (I237730,I237713,I28332);
DFFARX1 I_13825 (I237730,I2683,I237662,I237756,);
DFFARX1 I_13826 (I237756,I2683,I237662,I237651,);
DFFARX1 I_13827 (I28350,I2683,I237662,I237787,);
nand I_13828 (I237795,I237787,I28341);
not I_13829 (I237812,I237795);
DFFARX1 I_13830 (I237812,I2683,I237662,I237838,);
not I_13831 (I237846,I237838);
nor I_13832 (I237654,I237696,I237846);
DFFARX1 I_13833 (I28335,I2683,I237662,I237886,);
nor I_13834 (I237645,I237886,I237756);
nor I_13835 (I237636,I237886,I237812);
nand I_13836 (I237922,I28347,I28344);
and I_13837 (I237939,I237922,I28332);
DFFARX1 I_13838 (I237939,I2683,I237662,I237965,);
not I_13839 (I237973,I237965);
nand I_13840 (I237990,I237973,I237886);
nand I_13841 (I237639,I237973,I237795);
nor I_13842 (I238021,I28329,I28344);
and I_13843 (I238038,I237886,I238021);
nor I_13844 (I238055,I237973,I238038);
DFFARX1 I_13845 (I238055,I2683,I237662,I237648,);
nor I_13846 (I238086,I237688,I238021);
DFFARX1 I_13847 (I238086,I2683,I237662,I237633,);
nor I_13848 (I238117,I237965,I238021);
not I_13849 (I238134,I238117);
nand I_13850 (I237642,I238134,I237990);
not I_13851 (I238189,I2690);
DFFARX1 I_13852 (I158215,I2683,I238189,I238215,);
not I_13853 (I238223,I238215);
nand I_13854 (I238240,I158233,I158224);
and I_13855 (I238257,I238240,I158227);
DFFARX1 I_13856 (I238257,I2683,I238189,I238283,);
DFFARX1 I_13857 (I238283,I2683,I238189,I238178,);
DFFARX1 I_13858 (I158221,I2683,I238189,I238314,);
nand I_13859 (I238322,I238314,I158212);
not I_13860 (I238339,I238322);
DFFARX1 I_13861 (I238339,I2683,I238189,I238365,);
not I_13862 (I238373,I238365);
nor I_13863 (I238181,I238223,I238373);
DFFARX1 I_13864 (I158218,I2683,I238189,I238413,);
nor I_13865 (I238172,I238413,I238283);
nor I_13866 (I238163,I238413,I238339);
nand I_13867 (I238449,I158212,I158209);
and I_13868 (I238466,I238449,I158230);
DFFARX1 I_13869 (I238466,I2683,I238189,I238492,);
not I_13870 (I238500,I238492);
nand I_13871 (I238517,I238500,I238413);
nand I_13872 (I238166,I238500,I238322);
nor I_13873 (I238548,I158209,I158209);
and I_13874 (I238565,I238413,I238548);
nor I_13875 (I238582,I238500,I238565);
DFFARX1 I_13876 (I238582,I2683,I238189,I238175,);
nor I_13877 (I238613,I238215,I238548);
DFFARX1 I_13878 (I238613,I2683,I238189,I238160,);
nor I_13879 (I238644,I238492,I238548);
not I_13880 (I238661,I238644);
nand I_13881 (I238169,I238661,I238517);
not I_13882 (I238716,I2690);
DFFARX1 I_13883 (I311524,I2683,I238716,I238742,);
not I_13884 (I238750,I238742);
nand I_13885 (I238767,I311533,I311521);
and I_13886 (I238784,I238767,I311518);
DFFARX1 I_13887 (I238784,I2683,I238716,I238810,);
DFFARX1 I_13888 (I238810,I2683,I238716,I238705,);
DFFARX1 I_13889 (I311518,I2683,I238716,I238841,);
nand I_13890 (I238849,I238841,I311515);
not I_13891 (I238866,I238849);
DFFARX1 I_13892 (I238866,I2683,I238716,I238892,);
not I_13893 (I238900,I238892);
nor I_13894 (I238708,I238750,I238900);
DFFARX1 I_13895 (I311521,I2683,I238716,I238940,);
nor I_13896 (I238699,I238940,I238810);
nor I_13897 (I238690,I238940,I238866);
nand I_13898 (I238976,I311536,I311527);
and I_13899 (I238993,I238976,I311530);
DFFARX1 I_13900 (I238993,I2683,I238716,I239019,);
not I_13901 (I239027,I239019);
nand I_13902 (I239044,I239027,I238940);
nand I_13903 (I238693,I239027,I238849);
nor I_13904 (I239075,I311515,I311527);
and I_13905 (I239092,I238940,I239075);
nor I_13906 (I239109,I239027,I239092);
DFFARX1 I_13907 (I239109,I2683,I238716,I238702,);
nor I_13908 (I239140,I238742,I239075);
DFFARX1 I_13909 (I239140,I2683,I238716,I238687,);
nor I_13910 (I239171,I239019,I239075);
not I_13911 (I239188,I239171);
nand I_13912 (I238696,I239188,I239044);
not I_13913 (I239243,I2690);
DFFARX1 I_13914 (I60805,I2683,I239243,I239269,);
not I_13915 (I239277,I239269);
nand I_13916 (I239294,I60802,I60820);
and I_13917 (I239311,I239294,I60811);
DFFARX1 I_13918 (I239311,I2683,I239243,I239337,);
DFFARX1 I_13919 (I239337,I2683,I239243,I239232,);
DFFARX1 I_13920 (I60817,I2683,I239243,I239368,);
nand I_13921 (I239376,I239368,I60814);
not I_13922 (I239393,I239376);
DFFARX1 I_13923 (I239393,I2683,I239243,I239419,);
not I_13924 (I239427,I239419);
nor I_13925 (I239235,I239277,I239427);
DFFARX1 I_13926 (I60808,I2683,I239243,I239467,);
nor I_13927 (I239226,I239467,I239337);
nor I_13928 (I239217,I239467,I239393);
nand I_13929 (I239503,I60799,I60823);
and I_13930 (I239520,I239503,I60802);
DFFARX1 I_13931 (I239520,I2683,I239243,I239546,);
not I_13932 (I239554,I239546);
nand I_13933 (I239571,I239554,I239467);
nand I_13934 (I239220,I239554,I239376);
nor I_13935 (I239602,I60799,I60823);
and I_13936 (I239619,I239467,I239602);
nor I_13937 (I239636,I239554,I239619);
DFFARX1 I_13938 (I239636,I2683,I239243,I239229,);
nor I_13939 (I239667,I239269,I239602);
DFFARX1 I_13940 (I239667,I2683,I239243,I239214,);
nor I_13941 (I239698,I239546,I239602);
not I_13942 (I239715,I239698);
nand I_13943 (I239223,I239715,I239571);
not I_13944 (I239770,I2690);
DFFARX1 I_13945 (I283349,I2683,I239770,I239796,);
not I_13946 (I239804,I239796);
nand I_13947 (I239821,I283364,I283346);
and I_13948 (I239838,I239821,I283346);
DFFARX1 I_13949 (I239838,I2683,I239770,I239864,);
DFFARX1 I_13950 (I239864,I2683,I239770,I239759,);
DFFARX1 I_13951 (I283355,I2683,I239770,I239895,);
nand I_13952 (I239903,I239895,I283373);
not I_13953 (I239920,I239903);
DFFARX1 I_13954 (I239920,I2683,I239770,I239946,);
not I_13955 (I239954,I239946);
nor I_13956 (I239762,I239804,I239954);
DFFARX1 I_13957 (I283370,I2683,I239770,I239994,);
nor I_13958 (I239753,I239994,I239864);
nor I_13959 (I239744,I239994,I239920);
nand I_13960 (I240030,I283367,I283358);
and I_13961 (I240047,I240030,I283352);
DFFARX1 I_13962 (I240047,I2683,I239770,I240073,);
not I_13963 (I240081,I240073);
nand I_13964 (I240098,I240081,I239994);
nand I_13965 (I239747,I240081,I239903);
nor I_13966 (I240129,I283361,I283358);
and I_13967 (I240146,I239994,I240129);
nor I_13968 (I240163,I240081,I240146);
DFFARX1 I_13969 (I240163,I2683,I239770,I239756,);
nor I_13970 (I240194,I239796,I240129);
DFFARX1 I_13971 (I240194,I2683,I239770,I239741,);
nor I_13972 (I240225,I240073,I240129);
not I_13973 (I240242,I240225);
nand I_13974 (I239750,I240242,I240098);
not I_13975 (I240297,I2690);
DFFARX1 I_13976 (I4493,I2683,I240297,I240323,);
not I_13977 (I240331,I240323);
nand I_13978 (I240348,I4499,I4481);
and I_13979 (I240365,I240348,I4490);
DFFARX1 I_13980 (I240365,I2683,I240297,I240391,);
DFFARX1 I_13981 (I240391,I2683,I240297,I240286,);
DFFARX1 I_13982 (I4481,I2683,I240297,I240422,);
nand I_13983 (I240430,I240422,I4484);
not I_13984 (I240447,I240430);
DFFARX1 I_13985 (I240447,I2683,I240297,I240473,);
not I_13986 (I240481,I240473);
nor I_13987 (I240289,I240331,I240481);
DFFARX1 I_13988 (I4484,I2683,I240297,I240521,);
nor I_13989 (I240280,I240521,I240391);
nor I_13990 (I240271,I240521,I240447);
nand I_13991 (I240557,I4487,I4496);
and I_13992 (I240574,I240557,I4478);
DFFARX1 I_13993 (I240574,I2683,I240297,I240600,);
not I_13994 (I240608,I240600);
nand I_13995 (I240625,I240608,I240521);
nand I_13996 (I240274,I240608,I240430);
nor I_13997 (I240656,I4478,I4496);
and I_13998 (I240673,I240521,I240656);
nor I_13999 (I240690,I240608,I240673);
DFFARX1 I_14000 (I240690,I2683,I240297,I240283,);
nor I_14001 (I240721,I240323,I240656);
DFFARX1 I_14002 (I240721,I2683,I240297,I240268,);
nor I_14003 (I240752,I240600,I240656);
not I_14004 (I240769,I240752);
nand I_14005 (I240277,I240769,I240625);
not I_14006 (I240824,I2690);
DFFARX1 I_14007 (I189776,I2683,I240824,I240850,);
not I_14008 (I240858,I240850);
nand I_14009 (I240875,I189761,I189782);
and I_14010 (I240892,I240875,I189770);
DFFARX1 I_14011 (I240892,I2683,I240824,I240918,);
DFFARX1 I_14012 (I240918,I2683,I240824,I240813,);
DFFARX1 I_14013 (I189764,I2683,I240824,I240949,);
nand I_14014 (I240957,I240949,I189773);
not I_14015 (I240974,I240957);
DFFARX1 I_14016 (I240974,I2683,I240824,I241000,);
not I_14017 (I241008,I241000);
nor I_14018 (I240816,I240858,I241008);
DFFARX1 I_14019 (I189779,I2683,I240824,I241048,);
nor I_14020 (I240807,I241048,I240918);
nor I_14021 (I240798,I241048,I240974);
nand I_14022 (I241084,I189761,I189764);
and I_14023 (I241101,I241084,I189785);
DFFARX1 I_14024 (I241101,I2683,I240824,I241127,);
not I_14025 (I241135,I241127);
nand I_14026 (I241152,I241135,I241048);
nand I_14027 (I240801,I241135,I240957);
nor I_14028 (I241183,I189767,I189764);
and I_14029 (I241200,I241048,I241183);
nor I_14030 (I241217,I241135,I241200);
DFFARX1 I_14031 (I241217,I2683,I240824,I240810,);
nor I_14032 (I241248,I240850,I241183);
DFFARX1 I_14033 (I241248,I2683,I240824,I240795,);
nor I_14034 (I241279,I241127,I241183);
not I_14035 (I241296,I241279);
nand I_14036 (I240804,I241296,I241152);
not I_14037 (I241351,I2690);
DFFARX1 I_14038 (I380757,I2683,I241351,I241377,);
not I_14039 (I241385,I241377);
nand I_14040 (I241402,I380739,I380742);
and I_14041 (I241419,I241402,I380754);
DFFARX1 I_14042 (I241419,I2683,I241351,I241445,);
DFFARX1 I_14043 (I241445,I2683,I241351,I241340,);
DFFARX1 I_14044 (I380763,I2683,I241351,I241476,);
nand I_14045 (I241484,I241476,I380748);
not I_14046 (I241501,I241484);
DFFARX1 I_14047 (I241501,I2683,I241351,I241527,);
not I_14048 (I241535,I241527);
nor I_14049 (I241343,I241385,I241535);
DFFARX1 I_14050 (I380760,I2683,I241351,I241575,);
nor I_14051 (I241334,I241575,I241445);
nor I_14052 (I241325,I241575,I241501);
nand I_14053 (I241611,I380751,I380745);
and I_14054 (I241628,I241611,I380739);
DFFARX1 I_14055 (I241628,I2683,I241351,I241654,);
not I_14056 (I241662,I241654);
nand I_14057 (I241679,I241662,I241575);
nand I_14058 (I241328,I241662,I241484);
nor I_14059 (I241710,I380742,I380745);
and I_14060 (I241727,I241575,I241710);
nor I_14061 (I241744,I241662,I241727);
DFFARX1 I_14062 (I241744,I2683,I241351,I241337,);
nor I_14063 (I241775,I241377,I241710);
DFFARX1 I_14064 (I241775,I2683,I241351,I241322,);
nor I_14065 (I241806,I241654,I241710);
not I_14066 (I241823,I241806);
nand I_14067 (I241331,I241823,I241679);
not I_14068 (I241878,I2690);
DFFARX1 I_14069 (I402769,I2683,I241878,I241904,);
not I_14070 (I241912,I241904);
nand I_14071 (I241929,I402766,I402775);
and I_14072 (I241946,I241929,I402754);
DFFARX1 I_14073 (I241946,I2683,I241878,I241972,);
DFFARX1 I_14074 (I241972,I2683,I241878,I241867,);
DFFARX1 I_14075 (I402757,I2683,I241878,I242003,);
nand I_14076 (I242011,I242003,I402772);
not I_14077 (I242028,I242011);
DFFARX1 I_14078 (I242028,I2683,I241878,I242054,);
not I_14079 (I242062,I242054);
nor I_14080 (I241870,I241912,I242062);
DFFARX1 I_14081 (I402778,I2683,I241878,I242102,);
nor I_14082 (I241861,I242102,I241972);
nor I_14083 (I241852,I242102,I242028);
nand I_14084 (I242138,I402760,I402781);
and I_14085 (I242155,I242138,I402763);
DFFARX1 I_14086 (I242155,I2683,I241878,I242181,);
not I_14087 (I242189,I242181);
nand I_14088 (I242206,I242189,I242102);
nand I_14089 (I241855,I242189,I242011);
nor I_14090 (I242237,I402754,I402781);
and I_14091 (I242254,I242102,I242237);
nor I_14092 (I242271,I242189,I242254);
DFFARX1 I_14093 (I242271,I2683,I241878,I241864,);
nor I_14094 (I242302,I241904,I242237);
DFFARX1 I_14095 (I242302,I2683,I241878,I241849,);
nor I_14096 (I242333,I242181,I242237);
not I_14097 (I242350,I242333);
nand I_14098 (I241858,I242350,I242206);
not I_14099 (I242405,I2690);
DFFARX1 I_14100 (I56640,I2683,I242405,I242431,);
not I_14101 (I242439,I242431);
nand I_14102 (I242456,I56637,I56655);
and I_14103 (I242473,I242456,I56646);
DFFARX1 I_14104 (I242473,I2683,I242405,I242499,);
DFFARX1 I_14105 (I242499,I2683,I242405,I242394,);
DFFARX1 I_14106 (I56652,I2683,I242405,I242530,);
nand I_14107 (I242538,I242530,I56649);
not I_14108 (I242555,I242538);
DFFARX1 I_14109 (I242555,I2683,I242405,I242581,);
not I_14110 (I242589,I242581);
nor I_14111 (I242397,I242439,I242589);
DFFARX1 I_14112 (I56643,I2683,I242405,I242629,);
nor I_14113 (I242388,I242629,I242499);
nor I_14114 (I242379,I242629,I242555);
nand I_14115 (I242665,I56634,I56658);
and I_14116 (I242682,I242665,I56637);
DFFARX1 I_14117 (I242682,I2683,I242405,I242708,);
not I_14118 (I242716,I242708);
nand I_14119 (I242733,I242716,I242629);
nand I_14120 (I242382,I242716,I242538);
nor I_14121 (I242764,I56634,I56658);
and I_14122 (I242781,I242629,I242764);
nor I_14123 (I242798,I242716,I242781);
DFFARX1 I_14124 (I242798,I2683,I242405,I242391,);
nor I_14125 (I242829,I242431,I242764);
DFFARX1 I_14126 (I242829,I2683,I242405,I242376,);
nor I_14127 (I242860,I242708,I242764);
not I_14128 (I242877,I242860);
nand I_14129 (I242385,I242877,I242733);
not I_14130 (I242932,I2690);
DFFARX1 I_14131 (I357977,I2683,I242932,I242958,);
not I_14132 (I242966,I242958);
nand I_14133 (I242983,I357959,I357959);
and I_14134 (I243000,I242983,I357965);
DFFARX1 I_14135 (I243000,I2683,I242932,I243026,);
DFFARX1 I_14136 (I243026,I2683,I242932,I242921,);
DFFARX1 I_14137 (I357962,I2683,I242932,I243057,);
nand I_14138 (I243065,I243057,I357971);
not I_14139 (I243082,I243065);
DFFARX1 I_14140 (I243082,I2683,I242932,I243108,);
not I_14141 (I243116,I243108);
nor I_14142 (I242924,I242966,I243116);
DFFARX1 I_14143 (I357983,I2683,I242932,I243156,);
nor I_14144 (I242915,I243156,I243026);
nor I_14145 (I242906,I243156,I243082);
nand I_14146 (I243192,I357974,I357968);
and I_14147 (I243209,I243192,I357962);
DFFARX1 I_14148 (I243209,I2683,I242932,I243235,);
not I_14149 (I243243,I243235);
nand I_14150 (I243260,I243243,I243156);
nand I_14151 (I242909,I243243,I243065);
nor I_14152 (I243291,I357980,I357968);
and I_14153 (I243308,I243156,I243291);
nor I_14154 (I243325,I243243,I243308);
DFFARX1 I_14155 (I243325,I2683,I242932,I242918,);
nor I_14156 (I243356,I242958,I243291);
DFFARX1 I_14157 (I243356,I2683,I242932,I242903,);
nor I_14158 (I243387,I243235,I243291);
not I_14159 (I243404,I243387);
nand I_14160 (I242912,I243404,I243260);
not I_14161 (I243459,I2690);
DFFARX1 I_14162 (I294331,I2683,I243459,I243485,);
not I_14163 (I243493,I243485);
nand I_14164 (I243510,I294346,I294328);
and I_14165 (I243527,I243510,I294328);
DFFARX1 I_14166 (I243527,I2683,I243459,I243553,);
DFFARX1 I_14167 (I243553,I2683,I243459,I243448,);
DFFARX1 I_14168 (I294337,I2683,I243459,I243584,);
nand I_14169 (I243592,I243584,I294355);
not I_14170 (I243609,I243592);
DFFARX1 I_14171 (I243609,I2683,I243459,I243635,);
not I_14172 (I243643,I243635);
nor I_14173 (I243451,I243493,I243643);
DFFARX1 I_14174 (I294352,I2683,I243459,I243683,);
nor I_14175 (I243442,I243683,I243553);
nor I_14176 (I243433,I243683,I243609);
nand I_14177 (I243719,I294349,I294340);
and I_14178 (I243736,I243719,I294334);
DFFARX1 I_14179 (I243736,I2683,I243459,I243762,);
not I_14180 (I243770,I243762);
nand I_14181 (I243787,I243770,I243683);
nand I_14182 (I243436,I243770,I243592);
nor I_14183 (I243818,I294343,I294340);
and I_14184 (I243835,I243683,I243818);
nor I_14185 (I243852,I243770,I243835);
DFFARX1 I_14186 (I243852,I2683,I243459,I243445,);
nor I_14187 (I243883,I243485,I243818);
DFFARX1 I_14188 (I243883,I2683,I243459,I243430,);
nor I_14189 (I243914,I243762,I243818);
not I_14190 (I243931,I243914);
nand I_14191 (I243439,I243931,I243787);
not I_14192 (I243986,I2690);
DFFARX1 I_14193 (I75680,I2683,I243986,I244012,);
not I_14194 (I244020,I244012);
nand I_14195 (I244037,I75677,I75695);
and I_14196 (I244054,I244037,I75686);
DFFARX1 I_14197 (I244054,I2683,I243986,I244080,);
DFFARX1 I_14198 (I244080,I2683,I243986,I243975,);
DFFARX1 I_14199 (I75692,I2683,I243986,I244111,);
nand I_14200 (I244119,I244111,I75689);
not I_14201 (I244136,I244119);
DFFARX1 I_14202 (I244136,I2683,I243986,I244162,);
not I_14203 (I244170,I244162);
nor I_14204 (I243978,I244020,I244170);
DFFARX1 I_14205 (I75683,I2683,I243986,I244210,);
nor I_14206 (I243969,I244210,I244080);
nor I_14207 (I243960,I244210,I244136);
nand I_14208 (I244246,I75674,I75698);
and I_14209 (I244263,I244246,I75677);
DFFARX1 I_14210 (I244263,I2683,I243986,I244289,);
not I_14211 (I244297,I244289);
nand I_14212 (I244314,I244297,I244210);
nand I_14213 (I243963,I244297,I244119);
nor I_14214 (I244345,I75674,I75698);
and I_14215 (I244362,I244210,I244345);
nor I_14216 (I244379,I244297,I244362);
DFFARX1 I_14217 (I244379,I2683,I243986,I243972,);
nor I_14218 (I244410,I244012,I244345);
DFFARX1 I_14219 (I244410,I2683,I243986,I243957,);
nor I_14220 (I244441,I244289,I244345);
not I_14221 (I244458,I244441);
nand I_14222 (I243966,I244458,I244314);
not I_14223 (I244513,I2690);
DFFARX1 I_14224 (I104770,I2683,I244513,I244539,);
not I_14225 (I244547,I244539);
nand I_14226 (I244564,I104761,I104761);
and I_14227 (I244581,I244564,I104779);
DFFARX1 I_14228 (I244581,I2683,I244513,I244607,);
DFFARX1 I_14229 (I244607,I2683,I244513,I244502,);
DFFARX1 I_14230 (I104782,I2683,I244513,I244638,);
nand I_14231 (I244646,I244638,I104764);
not I_14232 (I244663,I244646);
DFFARX1 I_14233 (I244663,I2683,I244513,I244689,);
not I_14234 (I244697,I244689);
nor I_14235 (I244505,I244547,I244697);
DFFARX1 I_14236 (I104776,I2683,I244513,I244737,);
nor I_14237 (I244496,I244737,I244607);
nor I_14238 (I244487,I244737,I244663);
nand I_14239 (I244773,I104788,I104767);
and I_14240 (I244790,I244773,I104773);
DFFARX1 I_14241 (I244790,I2683,I244513,I244816,);
not I_14242 (I244824,I244816);
nand I_14243 (I244841,I244824,I244737);
nand I_14244 (I244490,I244824,I244646);
nor I_14245 (I244872,I104785,I104767);
and I_14246 (I244889,I244737,I244872);
nor I_14247 (I244906,I244824,I244889);
DFFARX1 I_14248 (I244906,I2683,I244513,I244499,);
nor I_14249 (I244937,I244539,I244872);
DFFARX1 I_14250 (I244937,I2683,I244513,I244484,);
nor I_14251 (I244968,I244816,I244872);
not I_14252 (I244985,I244968);
nand I_14253 (I244493,I244985,I244841);
not I_14254 (I245040,I2690);
DFFARX1 I_14255 (I379601,I2683,I245040,I245066,);
not I_14256 (I245074,I245066);
nand I_14257 (I245091,I379583,I379586);
and I_14258 (I245108,I245091,I379598);
DFFARX1 I_14259 (I245108,I2683,I245040,I245134,);
DFFARX1 I_14260 (I245134,I2683,I245040,I245029,);
DFFARX1 I_14261 (I379607,I2683,I245040,I245165,);
nand I_14262 (I245173,I245165,I379592);
not I_14263 (I245190,I245173);
DFFARX1 I_14264 (I245190,I2683,I245040,I245216,);
not I_14265 (I245224,I245216);
nor I_14266 (I245032,I245074,I245224);
DFFARX1 I_14267 (I379604,I2683,I245040,I245264,);
nor I_14268 (I245023,I245264,I245134);
nor I_14269 (I245014,I245264,I245190);
nand I_14270 (I245300,I379595,I379589);
and I_14271 (I245317,I245300,I379583);
DFFARX1 I_14272 (I245317,I2683,I245040,I245343,);
not I_14273 (I245351,I245343);
nand I_14274 (I245368,I245351,I245264);
nand I_14275 (I245017,I245351,I245173);
nor I_14276 (I245399,I379586,I379589);
and I_14277 (I245416,I245264,I245399);
nor I_14278 (I245433,I245351,I245416);
DFFARX1 I_14279 (I245433,I2683,I245040,I245026,);
nor I_14280 (I245464,I245066,I245399);
DFFARX1 I_14281 (I245464,I2683,I245040,I245011,);
nor I_14282 (I245495,I245343,I245399);
not I_14283 (I245512,I245495);
nand I_14284 (I245020,I245512,I245368);
not I_14285 (I245567,I2690);
DFFARX1 I_14286 (I170124,I2683,I245567,I245593,);
not I_14287 (I245601,I245593);
nand I_14288 (I245618,I170109,I170130);
and I_14289 (I245635,I245618,I170118);
DFFARX1 I_14290 (I245635,I2683,I245567,I245661,);
DFFARX1 I_14291 (I245661,I2683,I245567,I245556,);
DFFARX1 I_14292 (I170112,I2683,I245567,I245692,);
nand I_14293 (I245700,I245692,I170121);
not I_14294 (I245717,I245700);
DFFARX1 I_14295 (I245717,I2683,I245567,I245743,);
not I_14296 (I245751,I245743);
nor I_14297 (I245559,I245601,I245751);
DFFARX1 I_14298 (I170127,I2683,I245567,I245791,);
nor I_14299 (I245550,I245791,I245661);
nor I_14300 (I245541,I245791,I245717);
nand I_14301 (I245827,I170109,I170112);
and I_14302 (I245844,I245827,I170133);
DFFARX1 I_14303 (I245844,I2683,I245567,I245870,);
not I_14304 (I245878,I245870);
nand I_14305 (I245895,I245878,I245791);
nand I_14306 (I245544,I245878,I245700);
nor I_14307 (I245926,I170115,I170112);
and I_14308 (I245943,I245791,I245926);
nor I_14309 (I245960,I245878,I245943);
DFFARX1 I_14310 (I245960,I2683,I245567,I245553,);
nor I_14311 (I245991,I245593,I245926);
DFFARX1 I_14312 (I245991,I2683,I245567,I245538,);
nor I_14313 (I246022,I245870,I245926);
not I_14314 (I246039,I246022);
nand I_14315 (I245547,I246039,I245895);
not I_14316 (I246094,I2690);
DFFARX1 I_14317 (I27299,I2683,I246094,I246120,);
not I_14318 (I246128,I246120);
nand I_14319 (I246145,I27275,I27284);
and I_14320 (I246162,I246145,I27278);
DFFARX1 I_14321 (I246162,I2683,I246094,I246188,);
DFFARX1 I_14322 (I246188,I2683,I246094,I246083,);
DFFARX1 I_14323 (I27296,I2683,I246094,I246219,);
nand I_14324 (I246227,I246219,I27287);
not I_14325 (I246244,I246227);
DFFARX1 I_14326 (I246244,I2683,I246094,I246270,);
not I_14327 (I246278,I246270);
nor I_14328 (I246086,I246128,I246278);
DFFARX1 I_14329 (I27281,I2683,I246094,I246318,);
nor I_14330 (I246077,I246318,I246188);
nor I_14331 (I246068,I246318,I246244);
nand I_14332 (I246354,I27293,I27290);
and I_14333 (I246371,I246354,I27278);
DFFARX1 I_14334 (I246371,I2683,I246094,I246397,);
not I_14335 (I246405,I246397);
nand I_14336 (I246422,I246405,I246318);
nand I_14337 (I246071,I246405,I246227);
nor I_14338 (I246453,I27275,I27290);
and I_14339 (I246470,I246318,I246453);
nor I_14340 (I246487,I246405,I246470);
DFFARX1 I_14341 (I246487,I2683,I246094,I246080,);
nor I_14342 (I246518,I246120,I246453);
DFFARX1 I_14343 (I246518,I2683,I246094,I246065,);
nor I_14344 (I246549,I246397,I246453);
not I_14345 (I246566,I246549);
nand I_14346 (I246074,I246566,I246422);
not I_14347 (I246621,I2690);
DFFARX1 I_14348 (I29407,I2683,I246621,I246647,);
not I_14349 (I246655,I246647);
nand I_14350 (I246672,I29383,I29392);
and I_14351 (I246689,I246672,I29386);
DFFARX1 I_14352 (I246689,I2683,I246621,I246715,);
DFFARX1 I_14353 (I246715,I2683,I246621,I246610,);
DFFARX1 I_14354 (I29404,I2683,I246621,I246746,);
nand I_14355 (I246754,I246746,I29395);
not I_14356 (I246771,I246754);
DFFARX1 I_14357 (I246771,I2683,I246621,I246797,);
not I_14358 (I246805,I246797);
nor I_14359 (I246613,I246655,I246805);
DFFARX1 I_14360 (I29389,I2683,I246621,I246845,);
nor I_14361 (I246604,I246845,I246715);
nor I_14362 (I246595,I246845,I246771);
nand I_14363 (I246881,I29401,I29398);
and I_14364 (I246898,I246881,I29386);
DFFARX1 I_14365 (I246898,I2683,I246621,I246924,);
not I_14366 (I246932,I246924);
nand I_14367 (I246949,I246932,I246845);
nand I_14368 (I246598,I246932,I246754);
nor I_14369 (I246980,I29383,I29398);
and I_14370 (I246997,I246845,I246980);
nor I_14371 (I247014,I246932,I246997);
DFFARX1 I_14372 (I247014,I2683,I246621,I246607,);
nor I_14373 (I247045,I246647,I246980);
DFFARX1 I_14374 (I247045,I2683,I246621,I246592,);
nor I_14375 (I247076,I246924,I246980);
not I_14376 (I247093,I247076);
nand I_14377 (I246601,I247093,I246949);
not I_14378 (I247148,I2690);
DFFARX1 I_14379 (I392883,I2683,I247148,I247174,);
not I_14380 (I247182,I247174);
nand I_14381 (I247199,I392877,I392895);
and I_14382 (I247216,I247199,I392880);
DFFARX1 I_14383 (I247216,I2683,I247148,I247242,);
DFFARX1 I_14384 (I247242,I2683,I247148,I247137,);
DFFARX1 I_14385 (I392901,I2683,I247148,I247273,);
nand I_14386 (I247281,I247273,I392886);
not I_14387 (I247298,I247281);
DFFARX1 I_14388 (I247298,I2683,I247148,I247324,);
not I_14389 (I247332,I247324);
nor I_14390 (I247140,I247182,I247332);
DFFARX1 I_14391 (I392898,I2683,I247148,I247372,);
nor I_14392 (I247131,I247372,I247242);
nor I_14393 (I247122,I247372,I247298);
nand I_14394 (I247408,I392889,I392904);
and I_14395 (I247425,I247408,I392892);
DFFARX1 I_14396 (I247425,I2683,I247148,I247451,);
not I_14397 (I247459,I247451);
nand I_14398 (I247476,I247459,I247372);
nand I_14399 (I247125,I247459,I247281);
nor I_14400 (I247507,I392877,I392904);
and I_14401 (I247524,I247372,I247507);
nor I_14402 (I247541,I247459,I247524);
DFFARX1 I_14403 (I247541,I2683,I247148,I247134,);
nor I_14404 (I247572,I247174,I247507);
DFFARX1 I_14405 (I247572,I2683,I247148,I247119,);
nor I_14406 (I247603,I247451,I247507);
not I_14407 (I247620,I247603);
nand I_14408 (I247128,I247620,I247476);
not I_14409 (I247675,I2690);
DFFARX1 I_14410 (I11474,I2683,I247675,I247701,);
not I_14411 (I247709,I247701);
nand I_14412 (I247726,I11486,I11489);
and I_14413 (I247743,I247726,I11465);
DFFARX1 I_14414 (I247743,I2683,I247675,I247769,);
DFFARX1 I_14415 (I247769,I2683,I247675,I247664,);
DFFARX1 I_14416 (I11483,I2683,I247675,I247800,);
nand I_14417 (I247808,I247800,I11471);
not I_14418 (I247825,I247808);
DFFARX1 I_14419 (I247825,I2683,I247675,I247851,);
not I_14420 (I247859,I247851);
nor I_14421 (I247667,I247709,I247859);
DFFARX1 I_14422 (I11468,I2683,I247675,I247899,);
nor I_14423 (I247658,I247899,I247769);
nor I_14424 (I247649,I247899,I247825);
nand I_14425 (I247935,I11477,I11468);
and I_14426 (I247952,I247935,I11465);
DFFARX1 I_14427 (I247952,I2683,I247675,I247978,);
not I_14428 (I247986,I247978);
nand I_14429 (I248003,I247986,I247899);
nand I_14430 (I247652,I247986,I247808);
nor I_14431 (I248034,I11480,I11468);
and I_14432 (I248051,I247899,I248034);
nor I_14433 (I248068,I247986,I248051);
DFFARX1 I_14434 (I248068,I2683,I247675,I247661,);
nor I_14435 (I248099,I247701,I248034);
DFFARX1 I_14436 (I248099,I2683,I247675,I247646,);
nor I_14437 (I248130,I247978,I248034);
not I_14438 (I248147,I248130);
nand I_14439 (I247655,I248147,I248003);
not I_14440 (I248202,I2690);
DFFARX1 I_14441 (I353931,I2683,I248202,I248228,);
not I_14442 (I248236,I248228);
nand I_14443 (I248253,I353913,I353913);
and I_14444 (I248270,I248253,I353919);
DFFARX1 I_14445 (I248270,I2683,I248202,I248296,);
DFFARX1 I_14446 (I248296,I2683,I248202,I248191,);
DFFARX1 I_14447 (I353916,I2683,I248202,I248327,);
nand I_14448 (I248335,I248327,I353925);
not I_14449 (I248352,I248335);
DFFARX1 I_14450 (I248352,I2683,I248202,I248378,);
not I_14451 (I248386,I248378);
nor I_14452 (I248194,I248236,I248386);
DFFARX1 I_14453 (I353937,I2683,I248202,I248426,);
nor I_14454 (I248185,I248426,I248296);
nor I_14455 (I248176,I248426,I248352);
nand I_14456 (I248462,I353928,I353922);
and I_14457 (I248479,I248462,I353916);
DFFARX1 I_14458 (I248479,I2683,I248202,I248505,);
not I_14459 (I248513,I248505);
nand I_14460 (I248530,I248513,I248426);
nand I_14461 (I248179,I248513,I248335);
nor I_14462 (I248561,I353934,I353922);
and I_14463 (I248578,I248426,I248561);
nor I_14464 (I248595,I248513,I248578);
DFFARX1 I_14465 (I248595,I2683,I248202,I248188,);
nor I_14466 (I248626,I248228,I248561);
DFFARX1 I_14467 (I248626,I2683,I248202,I248173,);
nor I_14468 (I248657,I248505,I248561);
not I_14469 (I248674,I248657);
nand I_14470 (I248182,I248674,I248530);
not I_14471 (I248729,I2690);
DFFARX1 I_14472 (I379023,I2683,I248729,I248755,);
not I_14473 (I248763,I248755);
nand I_14474 (I248780,I379005,I379008);
and I_14475 (I248797,I248780,I379020);
DFFARX1 I_14476 (I248797,I2683,I248729,I248823,);
DFFARX1 I_14477 (I248823,I2683,I248729,I248718,);
DFFARX1 I_14478 (I379029,I2683,I248729,I248854,);
nand I_14479 (I248862,I248854,I379014);
not I_14480 (I248879,I248862);
DFFARX1 I_14481 (I248879,I2683,I248729,I248905,);
not I_14482 (I248913,I248905);
nor I_14483 (I248721,I248763,I248913);
DFFARX1 I_14484 (I379026,I2683,I248729,I248953,);
nor I_14485 (I248712,I248953,I248823);
nor I_14486 (I248703,I248953,I248879);
nand I_14487 (I248989,I379017,I379011);
and I_14488 (I249006,I248989,I379005);
DFFARX1 I_14489 (I249006,I2683,I248729,I249032,);
not I_14490 (I249040,I249032);
nand I_14491 (I249057,I249040,I248953);
nand I_14492 (I248706,I249040,I248862);
nor I_14493 (I249088,I379008,I379011);
and I_14494 (I249105,I248953,I249088);
nor I_14495 (I249122,I249040,I249105);
DFFARX1 I_14496 (I249122,I2683,I248729,I248715,);
nor I_14497 (I249153,I248755,I249088);
DFFARX1 I_14498 (I249153,I2683,I248729,I248700,);
nor I_14499 (I249184,I249032,I249088);
not I_14500 (I249201,I249184);
nand I_14501 (I248709,I249201,I249057);
not I_14502 (I249256,I2690);
DFFARX1 I_14503 (I59020,I2683,I249256,I249282,);
not I_14504 (I249290,I249282);
nand I_14505 (I249307,I59017,I59035);
and I_14506 (I249324,I249307,I59026);
DFFARX1 I_14507 (I249324,I2683,I249256,I249350,);
DFFARX1 I_14508 (I249350,I2683,I249256,I249245,);
DFFARX1 I_14509 (I59032,I2683,I249256,I249381,);
nand I_14510 (I249389,I249381,I59029);
not I_14511 (I249406,I249389);
DFFARX1 I_14512 (I249406,I2683,I249256,I249432,);
not I_14513 (I249440,I249432);
nor I_14514 (I249248,I249290,I249440);
DFFARX1 I_14515 (I59023,I2683,I249256,I249480,);
nor I_14516 (I249239,I249480,I249350);
nor I_14517 (I249230,I249480,I249406);
nand I_14518 (I249516,I59014,I59038);
and I_14519 (I249533,I249516,I59017);
DFFARX1 I_14520 (I249533,I2683,I249256,I249559,);
not I_14521 (I249567,I249559);
nand I_14522 (I249584,I249567,I249480);
nand I_14523 (I249233,I249567,I249389);
nor I_14524 (I249615,I59014,I59038);
and I_14525 (I249632,I249480,I249615);
nor I_14526 (I249649,I249567,I249632);
DFFARX1 I_14527 (I249649,I2683,I249256,I249242,);
nor I_14528 (I249680,I249282,I249615);
DFFARX1 I_14529 (I249680,I2683,I249256,I249227,);
nor I_14530 (I249711,I249559,I249615);
not I_14531 (I249728,I249711);
nand I_14532 (I249236,I249728,I249584);
not I_14533 (I249783,I2690);
DFFARX1 I_14534 (I83415,I2683,I249783,I249809,);
not I_14535 (I249817,I249809);
nand I_14536 (I249834,I83412,I83430);
and I_14537 (I249851,I249834,I83421);
DFFARX1 I_14538 (I249851,I2683,I249783,I249877,);
DFFARX1 I_14539 (I249877,I2683,I249783,I249772,);
DFFARX1 I_14540 (I83427,I2683,I249783,I249908,);
nand I_14541 (I249916,I249908,I83424);
not I_14542 (I249933,I249916);
DFFARX1 I_14543 (I249933,I2683,I249783,I249959,);
not I_14544 (I249967,I249959);
nor I_14545 (I249775,I249817,I249967);
DFFARX1 I_14546 (I83418,I2683,I249783,I250007,);
nor I_14547 (I249766,I250007,I249877);
nor I_14548 (I249757,I250007,I249933);
nand I_14549 (I250043,I83409,I83433);
and I_14550 (I250060,I250043,I83412);
DFFARX1 I_14551 (I250060,I2683,I249783,I250086,);
not I_14552 (I250094,I250086);
nand I_14553 (I250111,I250094,I250007);
nand I_14554 (I249760,I250094,I249916);
nor I_14555 (I250142,I83409,I83433);
and I_14556 (I250159,I250007,I250142);
nor I_14557 (I250176,I250094,I250159);
DFFARX1 I_14558 (I250176,I2683,I249783,I249769,);
nor I_14559 (I250207,I249809,I250142);
DFFARX1 I_14560 (I250207,I2683,I249783,I249754,);
nor I_14561 (I250238,I250086,I250142);
not I_14562 (I250255,I250238);
nand I_14563 (I249763,I250255,I250111);
not I_14564 (I250310,I2690);
DFFARX1 I_14565 (I190354,I2683,I250310,I250336,);
not I_14566 (I250344,I250336);
nand I_14567 (I250361,I190339,I190360);
and I_14568 (I250378,I250361,I190348);
DFFARX1 I_14569 (I250378,I2683,I250310,I250404,);
DFFARX1 I_14570 (I250404,I2683,I250310,I250299,);
DFFARX1 I_14571 (I190342,I2683,I250310,I250435,);
nand I_14572 (I250443,I250435,I190351);
not I_14573 (I250460,I250443);
DFFARX1 I_14574 (I250460,I2683,I250310,I250486,);
not I_14575 (I250494,I250486);
nor I_14576 (I250302,I250344,I250494);
DFFARX1 I_14577 (I190357,I2683,I250310,I250534,);
nor I_14578 (I250293,I250534,I250404);
nor I_14579 (I250284,I250534,I250460);
nand I_14580 (I250570,I190339,I190342);
and I_14581 (I250587,I250570,I190363);
DFFARX1 I_14582 (I250587,I2683,I250310,I250613,);
not I_14583 (I250621,I250613);
nand I_14584 (I250638,I250621,I250534);
nand I_14585 (I250287,I250621,I250443);
nor I_14586 (I250669,I190345,I190342);
and I_14587 (I250686,I250534,I250669);
nor I_14588 (I250703,I250621,I250686);
DFFARX1 I_14589 (I250703,I2683,I250310,I250296,);
nor I_14590 (I250734,I250336,I250669);
DFFARX1 I_14591 (I250734,I2683,I250310,I250281,);
nor I_14592 (I250765,I250613,I250669);
not I_14593 (I250782,I250765);
nand I_14594 (I250290,I250782,I250638);
not I_14595 (I250837,I2690);
DFFARX1 I_14596 (I7258,I2683,I250837,I250863,);
not I_14597 (I250871,I250863);
nand I_14598 (I250888,I7270,I7273);
and I_14599 (I250905,I250888,I7249);
DFFARX1 I_14600 (I250905,I2683,I250837,I250931,);
DFFARX1 I_14601 (I250931,I2683,I250837,I250826,);
DFFARX1 I_14602 (I7267,I2683,I250837,I250962,);
nand I_14603 (I250970,I250962,I7255);
not I_14604 (I250987,I250970);
DFFARX1 I_14605 (I250987,I2683,I250837,I251013,);
not I_14606 (I251021,I251013);
nor I_14607 (I250829,I250871,I251021);
DFFARX1 I_14608 (I7252,I2683,I250837,I251061,);
nor I_14609 (I250820,I251061,I250931);
nor I_14610 (I250811,I251061,I250987);
nand I_14611 (I251097,I7261,I7252);
and I_14612 (I251114,I251097,I7249);
DFFARX1 I_14613 (I251114,I2683,I250837,I251140,);
not I_14614 (I251148,I251140);
nand I_14615 (I251165,I251148,I251061);
nand I_14616 (I250814,I251148,I250970);
nor I_14617 (I251196,I7264,I7252);
and I_14618 (I251213,I251061,I251196);
nor I_14619 (I251230,I251148,I251213);
DFFARX1 I_14620 (I251230,I2683,I250837,I250823,);
nor I_14621 (I251261,I250863,I251196);
DFFARX1 I_14622 (I251261,I2683,I250837,I250808,);
nor I_14623 (I251292,I251140,I251196);
not I_14624 (I251309,I251292);
nand I_14625 (I250817,I251309,I251165);
not I_14626 (I251364,I2690);
DFFARX1 I_14627 (I228487,I2683,I251364,I251390,);
not I_14628 (I251398,I251390);
nand I_14629 (I251415,I228490,I228487);
and I_14630 (I251432,I251415,I228499);
DFFARX1 I_14631 (I251432,I2683,I251364,I251458,);
DFFARX1 I_14632 (I251458,I2683,I251364,I251353,);
DFFARX1 I_14633 (I228496,I2683,I251364,I251489,);
nand I_14634 (I251497,I251489,I228502);
not I_14635 (I251514,I251497);
DFFARX1 I_14636 (I251514,I2683,I251364,I251540,);
not I_14637 (I251548,I251540);
nor I_14638 (I251356,I251398,I251548);
DFFARX1 I_14639 (I228511,I2683,I251364,I251588,);
nor I_14640 (I251347,I251588,I251458);
nor I_14641 (I251338,I251588,I251514);
nand I_14642 (I251624,I228505,I228493);
and I_14643 (I251641,I251624,I228490);
DFFARX1 I_14644 (I251641,I2683,I251364,I251667,);
not I_14645 (I251675,I251667);
nand I_14646 (I251692,I251675,I251588);
nand I_14647 (I251341,I251675,I251497);
nor I_14648 (I251723,I228508,I228493);
and I_14649 (I251740,I251588,I251723);
nor I_14650 (I251757,I251675,I251740);
DFFARX1 I_14651 (I251757,I2683,I251364,I251350,);
nor I_14652 (I251788,I251390,I251723);
DFFARX1 I_14653 (I251788,I2683,I251364,I251335,);
nor I_14654 (I251819,I251667,I251723);
not I_14655 (I251836,I251819);
nand I_14656 (I251344,I251836,I251692);
not I_14657 (I251891,I2690);
DFFARX1 I_14658 (I406339,I2683,I251891,I251917,);
not I_14659 (I251925,I251917);
nand I_14660 (I251942,I406336,I406345);
and I_14661 (I251959,I251942,I406324);
DFFARX1 I_14662 (I251959,I2683,I251891,I251985,);
DFFARX1 I_14663 (I251985,I2683,I251891,I251880,);
DFFARX1 I_14664 (I406327,I2683,I251891,I252016,);
nand I_14665 (I252024,I252016,I406342);
not I_14666 (I252041,I252024);
DFFARX1 I_14667 (I252041,I2683,I251891,I252067,);
not I_14668 (I252075,I252067);
nor I_14669 (I251883,I251925,I252075);
DFFARX1 I_14670 (I406348,I2683,I251891,I252115,);
nor I_14671 (I251874,I252115,I251985);
nor I_14672 (I251865,I252115,I252041);
nand I_14673 (I252151,I406330,I406351);
and I_14674 (I252168,I252151,I406333);
DFFARX1 I_14675 (I252168,I2683,I251891,I252194,);
not I_14676 (I252202,I252194);
nand I_14677 (I252219,I252202,I252115);
nand I_14678 (I251868,I252202,I252024);
nor I_14679 (I252250,I406324,I406351);
and I_14680 (I252267,I252115,I252250);
nor I_14681 (I252284,I252202,I252267);
DFFARX1 I_14682 (I252284,I2683,I251891,I251877,);
nor I_14683 (I252315,I251917,I252250);
DFFARX1 I_14684 (I252315,I2683,I251891,I251862,);
nor I_14685 (I252346,I252194,I252250);
not I_14686 (I252363,I252346);
nand I_14687 (I251871,I252363,I252219);
not I_14688 (I252418,I2690);
DFFARX1 I_14689 (I230799,I2683,I252418,I252444,);
not I_14690 (I252452,I252444);
nand I_14691 (I252469,I230802,I230799);
and I_14692 (I252486,I252469,I230811);
DFFARX1 I_14693 (I252486,I2683,I252418,I252512,);
DFFARX1 I_14694 (I252512,I2683,I252418,I252407,);
DFFARX1 I_14695 (I230808,I2683,I252418,I252543,);
nand I_14696 (I252551,I252543,I230814);
not I_14697 (I252568,I252551);
DFFARX1 I_14698 (I252568,I2683,I252418,I252594,);
not I_14699 (I252602,I252594);
nor I_14700 (I252410,I252452,I252602);
DFFARX1 I_14701 (I230823,I2683,I252418,I252642,);
nor I_14702 (I252401,I252642,I252512);
nor I_14703 (I252392,I252642,I252568);
nand I_14704 (I252678,I230817,I230805);
and I_14705 (I252695,I252678,I230802);
DFFARX1 I_14706 (I252695,I2683,I252418,I252721,);
not I_14707 (I252729,I252721);
nand I_14708 (I252746,I252729,I252642);
nand I_14709 (I252395,I252729,I252551);
nor I_14710 (I252777,I230820,I230805);
and I_14711 (I252794,I252642,I252777);
nor I_14712 (I252811,I252729,I252794);
DFFARX1 I_14713 (I252811,I2683,I252418,I252404,);
nor I_14714 (I252842,I252444,I252777);
DFFARX1 I_14715 (I252842,I2683,I252418,I252389,);
nor I_14716 (I252873,I252721,I252777);
not I_14717 (I252890,I252873);
nand I_14718 (I252398,I252890,I252746);
not I_14719 (I252945,I2690);
DFFARX1 I_14720 (I384803,I2683,I252945,I252971,);
not I_14721 (I252979,I252971);
nand I_14722 (I252996,I384785,I384788);
and I_14723 (I253013,I252996,I384800);
DFFARX1 I_14724 (I253013,I2683,I252945,I253039,);
DFFARX1 I_14725 (I253039,I2683,I252945,I252934,);
DFFARX1 I_14726 (I384809,I2683,I252945,I253070,);
nand I_14727 (I253078,I253070,I384794);
not I_14728 (I253095,I253078);
DFFARX1 I_14729 (I253095,I2683,I252945,I253121,);
not I_14730 (I253129,I253121);
nor I_14731 (I252937,I252979,I253129);
DFFARX1 I_14732 (I384806,I2683,I252945,I253169,);
nor I_14733 (I252928,I253169,I253039);
nor I_14734 (I252919,I253169,I253095);
nand I_14735 (I253205,I384797,I384791);
and I_14736 (I253222,I253205,I384785);
DFFARX1 I_14737 (I253222,I2683,I252945,I253248,);
not I_14738 (I253256,I253248);
nand I_14739 (I253273,I253256,I253169);
nand I_14740 (I252922,I253256,I253078);
nor I_14741 (I253304,I384788,I384791);
and I_14742 (I253321,I253169,I253304);
nor I_14743 (I253338,I253256,I253321);
DFFARX1 I_14744 (I253338,I2683,I252945,I252931,);
nor I_14745 (I253369,I252971,I253304);
DFFARX1 I_14746 (I253369,I2683,I252945,I252916,);
nor I_14747 (I253400,I253248,I253304);
not I_14748 (I253417,I253400);
nand I_14749 (I252925,I253417,I253273);
not I_14750 (I253472,I2690);
DFFARX1 I_14751 (I101081,I2683,I253472,I253498,);
not I_14752 (I253506,I253498);
nand I_14753 (I253523,I101072,I101072);
and I_14754 (I253540,I253523,I101090);
DFFARX1 I_14755 (I253540,I2683,I253472,I253566,);
DFFARX1 I_14756 (I253566,I2683,I253472,I253461,);
DFFARX1 I_14757 (I101093,I2683,I253472,I253597,);
nand I_14758 (I253605,I253597,I101075);
not I_14759 (I253622,I253605);
DFFARX1 I_14760 (I253622,I2683,I253472,I253648,);
not I_14761 (I253656,I253648);
nor I_14762 (I253464,I253506,I253656);
DFFARX1 I_14763 (I101087,I2683,I253472,I253696,);
nor I_14764 (I253455,I253696,I253566);
nor I_14765 (I253446,I253696,I253622);
nand I_14766 (I253732,I101099,I101078);
and I_14767 (I253749,I253732,I101084);
DFFARX1 I_14768 (I253749,I2683,I253472,I253775,);
not I_14769 (I253783,I253775);
nand I_14770 (I253800,I253783,I253696);
nand I_14771 (I253449,I253783,I253605);
nor I_14772 (I253831,I101096,I101078);
and I_14773 (I253848,I253696,I253831);
nor I_14774 (I253865,I253783,I253848);
DFFARX1 I_14775 (I253865,I2683,I253472,I253458,);
nor I_14776 (I253896,I253498,I253831);
DFFARX1 I_14777 (I253896,I2683,I253472,I253443,);
nor I_14778 (I253927,I253775,I253831);
not I_14779 (I253944,I253927);
nand I_14780 (I253452,I253944,I253800);
not I_14781 (I253999,I2690);
DFFARX1 I_14782 (I102662,I2683,I253999,I254025,);
not I_14783 (I254033,I254025);
nand I_14784 (I254050,I102653,I102653);
and I_14785 (I254067,I254050,I102671);
DFFARX1 I_14786 (I254067,I2683,I253999,I254093,);
DFFARX1 I_14787 (I254093,I2683,I253999,I253988,);
DFFARX1 I_14788 (I102674,I2683,I253999,I254124,);
nand I_14789 (I254132,I254124,I102656);
not I_14790 (I254149,I254132);
DFFARX1 I_14791 (I254149,I2683,I253999,I254175,);
not I_14792 (I254183,I254175);
nor I_14793 (I253991,I254033,I254183);
DFFARX1 I_14794 (I102668,I2683,I253999,I254223,);
nor I_14795 (I253982,I254223,I254093);
nor I_14796 (I253973,I254223,I254149);
nand I_14797 (I254259,I102680,I102659);
and I_14798 (I254276,I254259,I102665);
DFFARX1 I_14799 (I254276,I2683,I253999,I254302,);
not I_14800 (I254310,I254302);
nand I_14801 (I254327,I254310,I254223);
nand I_14802 (I253976,I254310,I254132);
nor I_14803 (I254358,I102677,I102659);
and I_14804 (I254375,I254223,I254358);
nor I_14805 (I254392,I254310,I254375);
DFFARX1 I_14806 (I254392,I2683,I253999,I253985,);
nor I_14807 (I254423,I254025,I254358);
DFFARX1 I_14808 (I254423,I2683,I253999,I253970,);
nor I_14809 (I254454,I254302,I254358);
not I_14810 (I254471,I254454);
nand I_14811 (I253979,I254471,I254327);
not I_14812 (I254526,I2690);
DFFARX1 I_14813 (I15163,I2683,I254526,I254552,);
not I_14814 (I254560,I254552);
nand I_14815 (I254577,I15175,I15178);
and I_14816 (I254594,I254577,I15154);
DFFARX1 I_14817 (I254594,I2683,I254526,I254620,);
DFFARX1 I_14818 (I254620,I2683,I254526,I254515,);
DFFARX1 I_14819 (I15172,I2683,I254526,I254651,);
nand I_14820 (I254659,I254651,I15160);
not I_14821 (I254676,I254659);
DFFARX1 I_14822 (I254676,I2683,I254526,I254702,);
not I_14823 (I254710,I254702);
nor I_14824 (I254518,I254560,I254710);
DFFARX1 I_14825 (I15157,I2683,I254526,I254750,);
nor I_14826 (I254509,I254750,I254620);
nor I_14827 (I254500,I254750,I254676);
nand I_14828 (I254786,I15166,I15157);
and I_14829 (I254803,I254786,I15154);
DFFARX1 I_14830 (I254803,I2683,I254526,I254829,);
not I_14831 (I254837,I254829);
nand I_14832 (I254854,I254837,I254750);
nand I_14833 (I254503,I254837,I254659);
nor I_14834 (I254885,I15169,I15157);
and I_14835 (I254902,I254750,I254885);
nor I_14836 (I254919,I254837,I254902);
DFFARX1 I_14837 (I254919,I2683,I254526,I254512,);
nor I_14838 (I254950,I254552,I254885);
DFFARX1 I_14839 (I254950,I2683,I254526,I254497,);
nor I_14840 (I254981,I254829,I254885);
not I_14841 (I254998,I254981);
nand I_14842 (I254506,I254998,I254854);
not I_14843 (I255053,I2690);
DFFARX1 I_14844 (I366505,I2683,I255053,I255079,);
not I_14845 (I255087,I255079);
nand I_14846 (I255104,I366511,I366493);
and I_14847 (I255121,I255104,I366502);
DFFARX1 I_14848 (I255121,I2683,I255053,I255147,);
DFFARX1 I_14849 (I255147,I2683,I255053,I255042,);
DFFARX1 I_14850 (I366508,I2683,I255053,I255178,);
nand I_14851 (I255186,I255178,I366496);
not I_14852 (I255203,I255186);
DFFARX1 I_14853 (I255203,I2683,I255053,I255229,);
not I_14854 (I255237,I255229);
nor I_14855 (I255045,I255087,I255237);
DFFARX1 I_14856 (I366514,I2683,I255053,I255277,);
nor I_14857 (I255036,I255277,I255147);
nor I_14858 (I255027,I255277,I255203);
nand I_14859 (I255313,I366493,I366499);
and I_14860 (I255330,I255313,I366517);
DFFARX1 I_14861 (I255330,I2683,I255053,I255356,);
not I_14862 (I255364,I255356);
nand I_14863 (I255381,I255364,I255277);
nand I_14864 (I255030,I255364,I255186);
nor I_14865 (I255412,I366496,I366499);
and I_14866 (I255429,I255277,I255412);
nor I_14867 (I255446,I255364,I255429);
DFFARX1 I_14868 (I255446,I2683,I255053,I255039,);
nor I_14869 (I255477,I255079,I255412);
DFFARX1 I_14870 (I255477,I2683,I255053,I255024,);
nor I_14871 (I255508,I255356,I255412);
not I_14872 (I255525,I255508);
nand I_14873 (I255033,I255525,I255381);
not I_14874 (I255580,I2690);
DFFARX1 I_14875 (I331389,I2683,I255580,I255606,);
not I_14876 (I255614,I255606);
nand I_14877 (I255631,I331371,I331371);
and I_14878 (I255648,I255631,I331377);
DFFARX1 I_14879 (I255648,I2683,I255580,I255674,);
DFFARX1 I_14880 (I255674,I2683,I255580,I255569,);
DFFARX1 I_14881 (I331374,I2683,I255580,I255705,);
nand I_14882 (I255713,I255705,I331383);
not I_14883 (I255730,I255713);
DFFARX1 I_14884 (I255730,I2683,I255580,I255756,);
not I_14885 (I255764,I255756);
nor I_14886 (I255572,I255614,I255764);
DFFARX1 I_14887 (I331395,I2683,I255580,I255804,);
nor I_14888 (I255563,I255804,I255674);
nor I_14889 (I255554,I255804,I255730);
nand I_14890 (I255840,I331386,I331380);
and I_14891 (I255857,I255840,I331374);
DFFARX1 I_14892 (I255857,I2683,I255580,I255883,);
not I_14893 (I255891,I255883);
nand I_14894 (I255908,I255891,I255804);
nand I_14895 (I255557,I255891,I255713);
nor I_14896 (I255939,I331392,I331380);
and I_14897 (I255956,I255804,I255939);
nor I_14898 (I255973,I255891,I255956);
DFFARX1 I_14899 (I255973,I2683,I255580,I255566,);
nor I_14900 (I256004,I255606,I255939);
DFFARX1 I_14901 (I256004,I2683,I255580,I255551,);
nor I_14902 (I256035,I255883,I255939);
not I_14903 (I256052,I256035);
nand I_14904 (I255560,I256052,I255908);
not I_14905 (I256107,I2690);
DFFARX1 I_14906 (I50095,I2683,I256107,I256133,);
not I_14907 (I256141,I256133);
nand I_14908 (I256158,I50092,I50110);
and I_14909 (I256175,I256158,I50101);
DFFARX1 I_14910 (I256175,I2683,I256107,I256201,);
DFFARX1 I_14911 (I256201,I2683,I256107,I256096,);
DFFARX1 I_14912 (I50107,I2683,I256107,I256232,);
nand I_14913 (I256240,I256232,I50104);
not I_14914 (I256257,I256240);
DFFARX1 I_14915 (I256257,I2683,I256107,I256283,);
not I_14916 (I256291,I256283);
nor I_14917 (I256099,I256141,I256291);
DFFARX1 I_14918 (I50098,I2683,I256107,I256331,);
nor I_14919 (I256090,I256331,I256201);
nor I_14920 (I256081,I256331,I256257);
nand I_14921 (I256367,I50089,I50113);
and I_14922 (I256384,I256367,I50092);
DFFARX1 I_14923 (I256384,I2683,I256107,I256410,);
not I_14924 (I256418,I256410);
nand I_14925 (I256435,I256418,I256331);
nand I_14926 (I256084,I256418,I256240);
nor I_14927 (I256466,I50089,I50113);
and I_14928 (I256483,I256331,I256466);
nor I_14929 (I256500,I256418,I256483);
DFFARX1 I_14930 (I256500,I2683,I256107,I256093,);
nor I_14931 (I256531,I256133,I256466);
DFFARX1 I_14932 (I256531,I2683,I256107,I256078,);
nor I_14933 (I256562,I256410,I256466);
not I_14934 (I256579,I256562);
nand I_14935 (I256087,I256579,I256435);
not I_14936 (I256634,I2690);
DFFARX1 I_14937 (I338903,I2683,I256634,I256660,);
not I_14938 (I256668,I256660);
nand I_14939 (I256685,I338885,I338885);
and I_14940 (I256702,I256685,I338891);
DFFARX1 I_14941 (I256702,I2683,I256634,I256728,);
DFFARX1 I_14942 (I256728,I2683,I256634,I256623,);
DFFARX1 I_14943 (I338888,I2683,I256634,I256759,);
nand I_14944 (I256767,I256759,I338897);
not I_14945 (I256784,I256767);
DFFARX1 I_14946 (I256784,I2683,I256634,I256810,);
not I_14947 (I256818,I256810);
nor I_14948 (I256626,I256668,I256818);
DFFARX1 I_14949 (I338909,I2683,I256634,I256858,);
nor I_14950 (I256617,I256858,I256728);
nor I_14951 (I256608,I256858,I256784);
nand I_14952 (I256894,I338900,I338894);
and I_14953 (I256911,I256894,I338888);
DFFARX1 I_14954 (I256911,I2683,I256634,I256937,);
not I_14955 (I256945,I256937);
nand I_14956 (I256962,I256945,I256858);
nand I_14957 (I256611,I256945,I256767);
nor I_14958 (I256993,I338906,I338894);
and I_14959 (I257010,I256858,I256993);
nor I_14960 (I257027,I256945,I257010);
DFFARX1 I_14961 (I257027,I2683,I256634,I256620,);
nor I_14962 (I257058,I256660,I256993);
DFFARX1 I_14963 (I257058,I2683,I256634,I256605,);
nor I_14964 (I257089,I256937,I256993);
not I_14965 (I257106,I257089);
nand I_14966 (I256614,I257106,I256962);
not I_14967 (I257161,I2690);
DFFARX1 I_14968 (I204789,I2683,I257161,I257187,);
not I_14969 (I257195,I257187);
nand I_14970 (I257212,I204792,I204789);
and I_14971 (I257229,I257212,I204801);
DFFARX1 I_14972 (I257229,I2683,I257161,I257255,);
DFFARX1 I_14973 (I257255,I2683,I257161,I257150,);
DFFARX1 I_14974 (I204798,I2683,I257161,I257286,);
nand I_14975 (I257294,I257286,I204804);
not I_14976 (I257311,I257294);
DFFARX1 I_14977 (I257311,I2683,I257161,I257337,);
not I_14978 (I257345,I257337);
nor I_14979 (I257153,I257195,I257345);
DFFARX1 I_14980 (I204813,I2683,I257161,I257385,);
nor I_14981 (I257144,I257385,I257255);
nor I_14982 (I257135,I257385,I257311);
nand I_14983 (I257421,I204807,I204795);
and I_14984 (I257438,I257421,I204792);
DFFARX1 I_14985 (I257438,I2683,I257161,I257464,);
not I_14986 (I257472,I257464);
nand I_14987 (I257489,I257472,I257385);
nand I_14988 (I257138,I257472,I257294);
nor I_14989 (I257520,I204810,I204795);
and I_14990 (I257537,I257385,I257520);
nor I_14991 (I257554,I257472,I257537);
DFFARX1 I_14992 (I257554,I2683,I257161,I257147,);
nor I_14993 (I257585,I257187,I257520);
DFFARX1 I_14994 (I257585,I2683,I257161,I257132,);
nor I_14995 (I257616,I257464,I257520);
not I_14996 (I257633,I257616);
nand I_14997 (I257141,I257633,I257489);
not I_14998 (I257688,I2690);
DFFARX1 I_14999 (I296269,I2683,I257688,I257714,);
not I_15000 (I257722,I257714);
nand I_15001 (I257739,I296284,I296266);
and I_15002 (I257756,I257739,I296266);
DFFARX1 I_15003 (I257756,I2683,I257688,I257782,);
DFFARX1 I_15004 (I257782,I2683,I257688,I257677,);
DFFARX1 I_15005 (I296275,I2683,I257688,I257813,);
nand I_15006 (I257821,I257813,I296293);
not I_15007 (I257838,I257821);
DFFARX1 I_15008 (I257838,I2683,I257688,I257864,);
not I_15009 (I257872,I257864);
nor I_15010 (I257680,I257722,I257872);
DFFARX1 I_15011 (I296290,I2683,I257688,I257912,);
nor I_15012 (I257671,I257912,I257782);
nor I_15013 (I257662,I257912,I257838);
nand I_15014 (I257948,I296287,I296278);
and I_15015 (I257965,I257948,I296272);
DFFARX1 I_15016 (I257965,I2683,I257688,I257991,);
not I_15017 (I257999,I257991);
nand I_15018 (I258016,I257999,I257912);
nand I_15019 (I257665,I257999,I257821);
nor I_15020 (I258047,I296281,I296278);
and I_15021 (I258064,I257912,I258047);
nor I_15022 (I258081,I257999,I258064);
DFFARX1 I_15023 (I258081,I2683,I257688,I257674,);
nor I_15024 (I258112,I257714,I258047);
DFFARX1 I_15025 (I258112,I2683,I257688,I257659,);
nor I_15026 (I258143,I257991,I258047);
not I_15027 (I258160,I258143);
nand I_15028 (I257668,I258160,I258016);
not I_15029 (I258215,I2690);
DFFARX1 I_15030 (I110567,I2683,I258215,I258241,);
not I_15031 (I258249,I258241);
nand I_15032 (I258266,I110558,I110558);
and I_15033 (I258283,I258266,I110576);
DFFARX1 I_15034 (I258283,I2683,I258215,I258309,);
DFFARX1 I_15035 (I258309,I2683,I258215,I258204,);
DFFARX1 I_15036 (I110579,I2683,I258215,I258340,);
nand I_15037 (I258348,I258340,I110561);
not I_15038 (I258365,I258348);
DFFARX1 I_15039 (I258365,I2683,I258215,I258391,);
not I_15040 (I258399,I258391);
nor I_15041 (I258207,I258249,I258399);
DFFARX1 I_15042 (I110573,I2683,I258215,I258439,);
nor I_15043 (I258198,I258439,I258309);
nor I_15044 (I258189,I258439,I258365);
nand I_15045 (I258475,I110585,I110564);
and I_15046 (I258492,I258475,I110570);
DFFARX1 I_15047 (I258492,I2683,I258215,I258518,);
not I_15048 (I258526,I258518);
nand I_15049 (I258543,I258526,I258439);
nand I_15050 (I258192,I258526,I258348);
nor I_15051 (I258574,I110582,I110564);
and I_15052 (I258591,I258439,I258574);
nor I_15053 (I258608,I258526,I258591);
DFFARX1 I_15054 (I258608,I2683,I258215,I258201,);
nor I_15055 (I258639,I258241,I258574);
DFFARX1 I_15056 (I258639,I2683,I258215,I258186,);
nor I_15057 (I258670,I258518,I258574);
not I_15058 (I258687,I258670);
nand I_15059 (I258195,I258687,I258543);
not I_15060 (I258742,I2690);
DFFARX1 I_15061 (I123215,I2683,I258742,I258768,);
not I_15062 (I258776,I258768);
nand I_15063 (I258793,I123206,I123206);
and I_15064 (I258810,I258793,I123224);
DFFARX1 I_15065 (I258810,I2683,I258742,I258836,);
DFFARX1 I_15066 (I258836,I2683,I258742,I258731,);
DFFARX1 I_15067 (I123227,I2683,I258742,I258867,);
nand I_15068 (I258875,I258867,I123209);
not I_15069 (I258892,I258875);
DFFARX1 I_15070 (I258892,I2683,I258742,I258918,);
not I_15071 (I258926,I258918);
nor I_15072 (I258734,I258776,I258926);
DFFARX1 I_15073 (I123221,I2683,I258742,I258966,);
nor I_15074 (I258725,I258966,I258836);
nor I_15075 (I258716,I258966,I258892);
nand I_15076 (I259002,I123233,I123212);
and I_15077 (I259019,I259002,I123218);
DFFARX1 I_15078 (I259019,I2683,I258742,I259045,);
not I_15079 (I259053,I259045);
nand I_15080 (I259070,I259053,I258966);
nand I_15081 (I258719,I259053,I258875);
nor I_15082 (I259101,I123230,I123212);
and I_15083 (I259118,I258966,I259101);
nor I_15084 (I259135,I259053,I259118);
DFFARX1 I_15085 (I259135,I2683,I258742,I258728,);
nor I_15086 (I259166,I258768,I259101);
DFFARX1 I_15087 (I259166,I2683,I258742,I258713,);
nor I_15088 (I259197,I259045,I259101);
not I_15089 (I259214,I259197);
nand I_15090 (I258722,I259214,I259070);
not I_15091 (I259269,I2690);
DFFARX1 I_15092 (I68540,I2683,I259269,I259295,);
not I_15093 (I259303,I259295);
nand I_15094 (I259320,I68537,I68555);
and I_15095 (I259337,I259320,I68546);
DFFARX1 I_15096 (I259337,I2683,I259269,I259363,);
DFFARX1 I_15097 (I259363,I2683,I259269,I259258,);
DFFARX1 I_15098 (I68552,I2683,I259269,I259394,);
nand I_15099 (I259402,I259394,I68549);
not I_15100 (I259419,I259402);
DFFARX1 I_15101 (I259419,I2683,I259269,I259445,);
not I_15102 (I259453,I259445);
nor I_15103 (I259261,I259303,I259453);
DFFARX1 I_15104 (I68543,I2683,I259269,I259493,);
nor I_15105 (I259252,I259493,I259363);
nor I_15106 (I259243,I259493,I259419);
nand I_15107 (I259529,I68534,I68558);
and I_15108 (I259546,I259529,I68537);
DFFARX1 I_15109 (I259546,I2683,I259269,I259572,);
not I_15110 (I259580,I259572);
nand I_15111 (I259597,I259580,I259493);
nand I_15112 (I259246,I259580,I259402);
nor I_15113 (I259628,I68534,I68558);
and I_15114 (I259645,I259493,I259628);
nor I_15115 (I259662,I259580,I259645);
DFFARX1 I_15116 (I259662,I2683,I259269,I259255,);
nor I_15117 (I259693,I259295,I259628);
DFFARX1 I_15118 (I259693,I2683,I259269,I259240,);
nor I_15119 (I259724,I259572,I259628);
not I_15120 (I259741,I259724);
nand I_15121 (I259249,I259741,I259597);
not I_15122 (I259796,I2690);
DFFARX1 I_15123 (I343527,I2683,I259796,I259822,);
not I_15124 (I259830,I259822);
nand I_15125 (I259847,I343509,I343509);
and I_15126 (I259864,I259847,I343515);
DFFARX1 I_15127 (I259864,I2683,I259796,I259890,);
DFFARX1 I_15128 (I259890,I2683,I259796,I259785,);
DFFARX1 I_15129 (I343512,I2683,I259796,I259921,);
nand I_15130 (I259929,I259921,I343521);
not I_15131 (I259946,I259929);
DFFARX1 I_15132 (I259946,I2683,I259796,I259972,);
not I_15133 (I259980,I259972);
nor I_15134 (I259788,I259830,I259980);
DFFARX1 I_15135 (I343533,I2683,I259796,I260020,);
nor I_15136 (I259779,I260020,I259890);
nor I_15137 (I259770,I260020,I259946);
nand I_15138 (I260056,I343524,I343518);
and I_15139 (I260073,I260056,I343512);
DFFARX1 I_15140 (I260073,I2683,I259796,I260099,);
not I_15141 (I260107,I260099);
nand I_15142 (I260124,I260107,I260020);
nand I_15143 (I259773,I260107,I259929);
nor I_15144 (I260155,I343530,I343518);
and I_15145 (I260172,I260020,I260155);
nor I_15146 (I260189,I260107,I260172);
DFFARX1 I_15147 (I260189,I2683,I259796,I259782,);
nor I_15148 (I260220,I259822,I260155);
DFFARX1 I_15149 (I260220,I2683,I259796,I259767,);
nor I_15150 (I260251,I260099,I260155);
not I_15151 (I260268,I260251);
nand I_15152 (I259776,I260268,I260124);
not I_15153 (I260323,I2690);
DFFARX1 I_15154 (I216349,I2683,I260323,I260349,);
not I_15155 (I260357,I260349);
nand I_15156 (I260374,I216352,I216349);
and I_15157 (I260391,I260374,I216361);
DFFARX1 I_15158 (I260391,I2683,I260323,I260417,);
DFFARX1 I_15159 (I260417,I2683,I260323,I260312,);
DFFARX1 I_15160 (I216358,I2683,I260323,I260448,);
nand I_15161 (I260456,I260448,I216364);
not I_15162 (I260473,I260456);
DFFARX1 I_15163 (I260473,I2683,I260323,I260499,);
not I_15164 (I260507,I260499);
nor I_15165 (I260315,I260357,I260507);
DFFARX1 I_15166 (I216373,I2683,I260323,I260547,);
nor I_15167 (I260306,I260547,I260417);
nor I_15168 (I260297,I260547,I260473);
nand I_15169 (I260583,I216367,I216355);
and I_15170 (I260600,I260583,I216352);
DFFARX1 I_15171 (I260600,I2683,I260323,I260626,);
not I_15172 (I260634,I260626);
nand I_15173 (I260651,I260634,I260547);
nand I_15174 (I260300,I260634,I260456);
nor I_15175 (I260682,I216370,I216355);
and I_15176 (I260699,I260547,I260682);
nor I_15177 (I260716,I260634,I260699);
DFFARX1 I_15178 (I260716,I2683,I260323,I260309,);
nor I_15179 (I260747,I260349,I260682);
DFFARX1 I_15180 (I260747,I2683,I260323,I260294,);
nor I_15181 (I260778,I260626,I260682);
not I_15182 (I260795,I260778);
nand I_15183 (I260303,I260795,I260651);
not I_15184 (I260850,I2690);
DFFARX1 I_15185 (I66755,I2683,I260850,I260876,);
not I_15186 (I260884,I260876);
nand I_15187 (I260901,I66752,I66770);
and I_15188 (I260918,I260901,I66761);
DFFARX1 I_15189 (I260918,I2683,I260850,I260944,);
DFFARX1 I_15190 (I260944,I2683,I260850,I260839,);
DFFARX1 I_15191 (I66767,I2683,I260850,I260975,);
nand I_15192 (I260983,I260975,I66764);
not I_15193 (I261000,I260983);
DFFARX1 I_15194 (I261000,I2683,I260850,I261026,);
not I_15195 (I261034,I261026);
nor I_15196 (I260842,I260884,I261034);
DFFARX1 I_15197 (I66758,I2683,I260850,I261074,);
nor I_15198 (I260833,I261074,I260944);
nor I_15199 (I260824,I261074,I261000);
nand I_15200 (I261110,I66749,I66773);
and I_15201 (I261127,I261110,I66752);
DFFARX1 I_15202 (I261127,I2683,I260850,I261153,);
not I_15203 (I261161,I261153);
nand I_15204 (I261178,I261161,I261074);
nand I_15205 (I260827,I261161,I260983);
nor I_15206 (I261209,I66749,I66773);
and I_15207 (I261226,I261074,I261209);
nor I_15208 (I261243,I261161,I261226);
DFFARX1 I_15209 (I261243,I2683,I260850,I260836,);
nor I_15210 (I261274,I260876,I261209);
DFFARX1 I_15211 (I261274,I2683,I260850,I260821,);
nor I_15212 (I261305,I261153,I261209);
not I_15213 (I261322,I261305);
nand I_15214 (I260830,I261322,I261178);
not I_15215 (I261377,I2690);
DFFARX1 I_15216 (I217505,I2683,I261377,I261403,);
not I_15217 (I261411,I261403);
nand I_15218 (I261428,I217508,I217505);
and I_15219 (I261445,I261428,I217517);
DFFARX1 I_15220 (I261445,I2683,I261377,I261471,);
DFFARX1 I_15221 (I261471,I2683,I261377,I261366,);
DFFARX1 I_15222 (I217514,I2683,I261377,I261502,);
nand I_15223 (I261510,I261502,I217520);
not I_15224 (I261527,I261510);
DFFARX1 I_15225 (I261527,I2683,I261377,I261553,);
not I_15226 (I261561,I261553);
nor I_15227 (I261369,I261411,I261561);
DFFARX1 I_15228 (I217529,I2683,I261377,I261601,);
nor I_15229 (I261360,I261601,I261471);
nor I_15230 (I261351,I261601,I261527);
nand I_15231 (I261637,I217523,I217511);
and I_15232 (I261654,I261637,I217508);
DFFARX1 I_15233 (I261654,I2683,I261377,I261680,);
not I_15234 (I261688,I261680);
nand I_15235 (I261705,I261688,I261601);
nand I_15236 (I261354,I261688,I261510);
nor I_15237 (I261736,I217526,I217511);
and I_15238 (I261753,I261601,I261736);
nor I_15239 (I261770,I261688,I261753);
DFFARX1 I_15240 (I261770,I2683,I261377,I261363,);
nor I_15241 (I261801,I261403,I261736);
DFFARX1 I_15242 (I261801,I2683,I261377,I261348,);
nor I_15243 (I261832,I261680,I261736);
not I_15244 (I261849,I261832);
nand I_15245 (I261357,I261849,I261705);
not I_15246 (I261904,I2690);
DFFARX1 I_15247 (I222707,I2683,I261904,I261930,);
not I_15248 (I261938,I261930);
nand I_15249 (I261955,I222710,I222707);
and I_15250 (I261972,I261955,I222719);
DFFARX1 I_15251 (I261972,I2683,I261904,I261998,);
DFFARX1 I_15252 (I261998,I2683,I261904,I261893,);
DFFARX1 I_15253 (I222716,I2683,I261904,I262029,);
nand I_15254 (I262037,I262029,I222722);
not I_15255 (I262054,I262037);
DFFARX1 I_15256 (I262054,I2683,I261904,I262080,);
not I_15257 (I262088,I262080);
nor I_15258 (I261896,I261938,I262088);
DFFARX1 I_15259 (I222731,I2683,I261904,I262128,);
nor I_15260 (I261887,I262128,I261998);
nor I_15261 (I261878,I262128,I262054);
nand I_15262 (I262164,I222725,I222713);
and I_15263 (I262181,I262164,I222710);
DFFARX1 I_15264 (I262181,I2683,I261904,I262207,);
not I_15265 (I262215,I262207);
nand I_15266 (I262232,I262215,I262128);
nand I_15267 (I261881,I262215,I262037);
nor I_15268 (I262263,I222728,I222713);
and I_15269 (I262280,I262128,I262263);
nor I_15270 (I262297,I262215,I262280);
DFFARX1 I_15271 (I262297,I2683,I261904,I261890,);
nor I_15272 (I262328,I261930,I262263);
DFFARX1 I_15273 (I262328,I2683,I261904,I261875,);
nor I_15274 (I262359,I262207,I262263);
not I_15275 (I262376,I262359);
nand I_15276 (I261884,I262376,I262232);
not I_15277 (I262431,I2690);
DFFARX1 I_15278 (I155835,I2683,I262431,I262457,);
not I_15279 (I262465,I262457);
nand I_15280 (I262482,I155853,I155844);
and I_15281 (I262499,I262482,I155847);
DFFARX1 I_15282 (I262499,I2683,I262431,I262525,);
DFFARX1 I_15283 (I262525,I2683,I262431,I262420,);
DFFARX1 I_15284 (I155841,I2683,I262431,I262556,);
nand I_15285 (I262564,I262556,I155832);
not I_15286 (I262581,I262564);
DFFARX1 I_15287 (I262581,I2683,I262431,I262607,);
not I_15288 (I262615,I262607);
nor I_15289 (I262423,I262465,I262615);
DFFARX1 I_15290 (I155838,I2683,I262431,I262655,);
nor I_15291 (I262414,I262655,I262525);
nor I_15292 (I262405,I262655,I262581);
nand I_15293 (I262691,I155832,I155829);
and I_15294 (I262708,I262691,I155850);
DFFARX1 I_15295 (I262708,I2683,I262431,I262734,);
not I_15296 (I262742,I262734);
nand I_15297 (I262759,I262742,I262655);
nand I_15298 (I262408,I262742,I262564);
nor I_15299 (I262790,I155829,I155829);
and I_15300 (I262807,I262655,I262790);
nor I_15301 (I262824,I262742,I262807);
DFFARX1 I_15302 (I262824,I2683,I262431,I262417,);
nor I_15303 (I262855,I262457,I262790);
DFFARX1 I_15304 (I262855,I2683,I262431,I262402,);
nor I_15305 (I262886,I262734,I262790);
not I_15306 (I262903,I262886);
nand I_15307 (I262411,I262903,I262759);
not I_15308 (I262958,I2690);
DFFARX1 I_15309 (I381335,I2683,I262958,I262984,);
not I_15310 (I262992,I262984);
nand I_15311 (I263009,I381317,I381320);
and I_15312 (I263026,I263009,I381332);
DFFARX1 I_15313 (I263026,I2683,I262958,I263052,);
DFFARX1 I_15314 (I263052,I2683,I262958,I262947,);
DFFARX1 I_15315 (I381341,I2683,I262958,I263083,);
nand I_15316 (I263091,I263083,I381326);
not I_15317 (I263108,I263091);
DFFARX1 I_15318 (I263108,I2683,I262958,I263134,);
not I_15319 (I263142,I263134);
nor I_15320 (I262950,I262992,I263142);
DFFARX1 I_15321 (I381338,I2683,I262958,I263182,);
nor I_15322 (I262941,I263182,I263052);
nor I_15323 (I262932,I263182,I263108);
nand I_15324 (I263218,I381329,I381323);
and I_15325 (I263235,I263218,I381317);
DFFARX1 I_15326 (I263235,I2683,I262958,I263261,);
not I_15327 (I263269,I263261);
nand I_15328 (I263286,I263269,I263182);
nand I_15329 (I262935,I263269,I263091);
nor I_15330 (I263317,I381320,I381323);
and I_15331 (I263334,I263182,I263317);
nor I_15332 (I263351,I263269,I263334);
DFFARX1 I_15333 (I263351,I2683,I262958,I262944,);
nor I_15334 (I263382,I262984,I263317);
DFFARX1 I_15335 (I263382,I2683,I262958,I262929,);
nor I_15336 (I263413,I263261,I263317);
not I_15337 (I263430,I263413);
nand I_15338 (I262938,I263430,I263286);
not I_15339 (I263485,I2690);
DFFARX1 I_15340 (I124269,I2683,I263485,I263511,);
not I_15341 (I263519,I263511);
nand I_15342 (I263536,I124260,I124260);
and I_15343 (I263553,I263536,I124278);
DFFARX1 I_15344 (I263553,I2683,I263485,I263579,);
DFFARX1 I_15345 (I263579,I2683,I263485,I263474,);
DFFARX1 I_15346 (I124281,I2683,I263485,I263610,);
nand I_15347 (I263618,I263610,I124263);
not I_15348 (I263635,I263618);
DFFARX1 I_15349 (I263635,I2683,I263485,I263661,);
not I_15350 (I263669,I263661);
nor I_15351 (I263477,I263519,I263669);
DFFARX1 I_15352 (I124275,I2683,I263485,I263709,);
nor I_15353 (I263468,I263709,I263579);
nor I_15354 (I263459,I263709,I263635);
nand I_15355 (I263745,I124287,I124266);
and I_15356 (I263762,I263745,I124272);
DFFARX1 I_15357 (I263762,I2683,I263485,I263788,);
not I_15358 (I263796,I263788);
nand I_15359 (I263813,I263796,I263709);
nand I_15360 (I263462,I263796,I263618);
nor I_15361 (I263844,I124284,I124266);
and I_15362 (I263861,I263709,I263844);
nor I_15363 (I263878,I263796,I263861);
DFFARX1 I_15364 (I263878,I2683,I263485,I263471,);
nor I_15365 (I263909,I263511,I263844);
DFFARX1 I_15366 (I263909,I2683,I263485,I263456,);
nor I_15367 (I263940,I263788,I263844);
not I_15368 (I263957,I263940);
nand I_15369 (I263465,I263957,I263813);
not I_15370 (I264012,I2690);
DFFARX1 I_15371 (I17271,I2683,I264012,I264038,);
not I_15372 (I264046,I264038);
nand I_15373 (I264063,I17283,I17286);
and I_15374 (I264080,I264063,I17262);
DFFARX1 I_15375 (I264080,I2683,I264012,I264106,);
DFFARX1 I_15376 (I264106,I2683,I264012,I264001,);
DFFARX1 I_15377 (I17280,I2683,I264012,I264137,);
nand I_15378 (I264145,I264137,I17268);
not I_15379 (I264162,I264145);
DFFARX1 I_15380 (I264162,I2683,I264012,I264188,);
not I_15381 (I264196,I264188);
nor I_15382 (I264004,I264046,I264196);
DFFARX1 I_15383 (I17265,I2683,I264012,I264236,);
nor I_15384 (I263995,I264236,I264106);
nor I_15385 (I263986,I264236,I264162);
nand I_15386 (I264272,I17274,I17265);
and I_15387 (I264289,I264272,I17262);
DFFARX1 I_15388 (I264289,I2683,I264012,I264315,);
not I_15389 (I264323,I264315);
nand I_15390 (I264340,I264323,I264236);
nand I_15391 (I263989,I264323,I264145);
nor I_15392 (I264371,I17277,I17265);
and I_15393 (I264388,I264236,I264371);
nor I_15394 (I264405,I264323,I264388);
DFFARX1 I_15395 (I264405,I2683,I264012,I263998,);
nor I_15396 (I264436,I264038,I264371);
DFFARX1 I_15397 (I264436,I2683,I264012,I263983,);
nor I_15398 (I264467,I264315,I264371);
not I_15399 (I264484,I264467);
nand I_15400 (I263992,I264484,I264340);
not I_15401 (I264539,I2690);
DFFARX1 I_15402 (I135061,I2683,I264539,I264565,);
not I_15403 (I264573,I264565);
nand I_15404 (I264590,I135058,I135067);
and I_15405 (I264607,I264590,I135076);
DFFARX1 I_15406 (I264607,I2683,I264539,I264633,);
DFFARX1 I_15407 (I264633,I2683,I264539,I264528,);
DFFARX1 I_15408 (I135079,I2683,I264539,I264664,);
nand I_15409 (I264672,I264664,I135082);
not I_15410 (I264689,I264672);
DFFARX1 I_15411 (I264689,I2683,I264539,I264715,);
not I_15412 (I264723,I264715);
nor I_15413 (I264531,I264573,I264723);
DFFARX1 I_15414 (I135055,I2683,I264539,I264763,);
nor I_15415 (I264522,I264763,I264633);
nor I_15416 (I264513,I264763,I264689);
nand I_15417 (I264799,I135070,I135073);
and I_15418 (I264816,I264799,I135064);
DFFARX1 I_15419 (I264816,I2683,I264539,I264842,);
not I_15420 (I264850,I264842);
nand I_15421 (I264867,I264850,I264763);
nand I_15422 (I264516,I264850,I264672);
nor I_15423 (I264898,I135055,I135073);
and I_15424 (I264915,I264763,I264898);
nor I_15425 (I264932,I264850,I264915);
DFFARX1 I_15426 (I264932,I2683,I264539,I264525,);
nor I_15427 (I264963,I264565,I264898);
DFFARX1 I_15428 (I264963,I2683,I264539,I264510,);
nor I_15429 (I264994,I264842,I264898);
not I_15430 (I265011,I264994);
nand I_15431 (I264519,I265011,I264867);
not I_15432 (I265066,I2690);
DFFARX1 I_15433 (I113202,I2683,I265066,I265092,);
not I_15434 (I265100,I265092);
nand I_15435 (I265117,I113193,I113193);
and I_15436 (I265134,I265117,I113211);
DFFARX1 I_15437 (I265134,I2683,I265066,I265160,);
DFFARX1 I_15438 (I265160,I2683,I265066,I265055,);
DFFARX1 I_15439 (I113214,I2683,I265066,I265191,);
nand I_15440 (I265199,I265191,I113196);
not I_15441 (I265216,I265199);
DFFARX1 I_15442 (I265216,I2683,I265066,I265242,);
not I_15443 (I265250,I265242);
nor I_15444 (I265058,I265100,I265250);
DFFARX1 I_15445 (I113208,I2683,I265066,I265290,);
nor I_15446 (I265049,I265290,I265160);
nor I_15447 (I265040,I265290,I265216);
nand I_15448 (I265326,I113220,I113199);
and I_15449 (I265343,I265326,I113205);
DFFARX1 I_15450 (I265343,I2683,I265066,I265369,);
not I_15451 (I265377,I265369);
nand I_15452 (I265394,I265377,I265290);
nand I_15453 (I265043,I265377,I265199);
nor I_15454 (I265425,I113217,I113199);
and I_15455 (I265442,I265290,I265425);
nor I_15456 (I265459,I265377,I265442);
DFFARX1 I_15457 (I265459,I2683,I265066,I265052,);
nor I_15458 (I265490,I265092,I265425);
DFFARX1 I_15459 (I265490,I2683,I265066,I265037,);
nor I_15460 (I265521,I265369,I265425);
not I_15461 (I265538,I265521);
nand I_15462 (I265046,I265538,I265394);
not I_15463 (I265593,I2690);
DFFARX1 I_15464 (I107932,I2683,I265593,I265619,);
not I_15465 (I265627,I265619);
nand I_15466 (I265644,I107923,I107923);
and I_15467 (I265661,I265644,I107941);
DFFARX1 I_15468 (I265661,I2683,I265593,I265687,);
DFFARX1 I_15469 (I265687,I2683,I265593,I265582,);
DFFARX1 I_15470 (I107944,I2683,I265593,I265718,);
nand I_15471 (I265726,I265718,I107926);
not I_15472 (I265743,I265726);
DFFARX1 I_15473 (I265743,I2683,I265593,I265769,);
not I_15474 (I265777,I265769);
nor I_15475 (I265585,I265627,I265777);
DFFARX1 I_15476 (I107938,I2683,I265593,I265817,);
nor I_15477 (I265576,I265817,I265687);
nor I_15478 (I265567,I265817,I265743);
nand I_15479 (I265853,I107950,I107929);
and I_15480 (I265870,I265853,I107935);
DFFARX1 I_15481 (I265870,I2683,I265593,I265896,);
not I_15482 (I265904,I265896);
nand I_15483 (I265921,I265904,I265817);
nand I_15484 (I265570,I265904,I265726);
nor I_15485 (I265952,I107947,I107929);
and I_15486 (I265969,I265817,I265952);
nor I_15487 (I265986,I265904,I265969);
DFFARX1 I_15488 (I265986,I2683,I265593,I265579,);
nor I_15489 (I266017,I265619,I265952);
DFFARX1 I_15490 (I266017,I2683,I265593,I265564,);
nor I_15491 (I266048,I265896,I265952);
not I_15492 (I266065,I266048);
nand I_15493 (I265573,I266065,I265921);
not I_15494 (I266120,I2690);
DFFARX1 I_15495 (I336013,I2683,I266120,I266146,);
not I_15496 (I266154,I266146);
nand I_15497 (I266171,I335995,I335995);
and I_15498 (I266188,I266171,I336001);
DFFARX1 I_15499 (I266188,I2683,I266120,I266214,);
DFFARX1 I_15500 (I266214,I2683,I266120,I266109,);
DFFARX1 I_15501 (I335998,I2683,I266120,I266245,);
nand I_15502 (I266253,I266245,I336007);
not I_15503 (I266270,I266253);
DFFARX1 I_15504 (I266270,I2683,I266120,I266296,);
not I_15505 (I266304,I266296);
nor I_15506 (I266112,I266154,I266304);
DFFARX1 I_15507 (I336019,I2683,I266120,I266344,);
nor I_15508 (I266103,I266344,I266214);
nor I_15509 (I266094,I266344,I266270);
nand I_15510 (I266380,I336010,I336004);
and I_15511 (I266397,I266380,I335998);
DFFARX1 I_15512 (I266397,I2683,I266120,I266423,);
not I_15513 (I266431,I266423);
nand I_15514 (I266448,I266431,I266344);
nand I_15515 (I266097,I266431,I266253);
nor I_15516 (I266479,I336016,I336004);
and I_15517 (I266496,I266344,I266479);
nor I_15518 (I266513,I266431,I266496);
DFFARX1 I_15519 (I266513,I2683,I266120,I266106,);
nor I_15520 (I266544,I266146,I266479);
DFFARX1 I_15521 (I266544,I2683,I266120,I266091,);
nor I_15522 (I266575,I266423,I266479);
not I_15523 (I266592,I266575);
nand I_15524 (I266100,I266592,I266448);
not I_15525 (I266647,I2690);
DFFARX1 I_15526 (I40474,I2683,I266647,I266673,);
not I_15527 (I266681,I266673);
nand I_15528 (I266698,I40450,I40459);
and I_15529 (I266715,I266698,I40453);
DFFARX1 I_15530 (I266715,I2683,I266647,I266741,);
DFFARX1 I_15531 (I266741,I2683,I266647,I266636,);
DFFARX1 I_15532 (I40471,I2683,I266647,I266772,);
nand I_15533 (I266780,I266772,I40462);
not I_15534 (I266797,I266780);
DFFARX1 I_15535 (I266797,I2683,I266647,I266823,);
not I_15536 (I266831,I266823);
nor I_15537 (I266639,I266681,I266831);
DFFARX1 I_15538 (I40456,I2683,I266647,I266871,);
nor I_15539 (I266630,I266871,I266741);
nor I_15540 (I266621,I266871,I266797);
nand I_15541 (I266907,I40468,I40465);
and I_15542 (I266924,I266907,I40453);
DFFARX1 I_15543 (I266924,I2683,I266647,I266950,);
not I_15544 (I266958,I266950);
nand I_15545 (I266975,I266958,I266871);
nand I_15546 (I266624,I266958,I266780);
nor I_15547 (I267006,I40450,I40465);
and I_15548 (I267023,I266871,I267006);
nor I_15549 (I267040,I266958,I267023);
DFFARX1 I_15550 (I267040,I2683,I266647,I266633,);
nor I_15551 (I267071,I266673,I267006);
DFFARX1 I_15552 (I267071,I2683,I266647,I266618,);
nor I_15553 (I267102,I266950,I267006);
not I_15554 (I267119,I267102);
nand I_15555 (I266627,I267119,I266975);
not I_15556 (I267174,I2690);
DFFARX1 I_15557 (I65565,I2683,I267174,I267200,);
not I_15558 (I267208,I267200);
nand I_15559 (I267225,I65562,I65580);
and I_15560 (I267242,I267225,I65571);
DFFARX1 I_15561 (I267242,I2683,I267174,I267268,);
DFFARX1 I_15562 (I267268,I2683,I267174,I267163,);
DFFARX1 I_15563 (I65577,I2683,I267174,I267299,);
nand I_15564 (I267307,I267299,I65574);
not I_15565 (I267324,I267307);
DFFARX1 I_15566 (I267324,I2683,I267174,I267350,);
not I_15567 (I267358,I267350);
nor I_15568 (I267166,I267208,I267358);
DFFARX1 I_15569 (I65568,I2683,I267174,I267398,);
nor I_15570 (I267157,I267398,I267268);
nor I_15571 (I267148,I267398,I267324);
nand I_15572 (I267434,I65559,I65583);
and I_15573 (I267451,I267434,I65562);
DFFARX1 I_15574 (I267451,I2683,I267174,I267477,);
not I_15575 (I267485,I267477);
nand I_15576 (I267502,I267485,I267398);
nand I_15577 (I267151,I267485,I267307);
nor I_15578 (I267533,I65559,I65583);
and I_15579 (I267550,I267398,I267533);
nor I_15580 (I267567,I267485,I267550);
DFFARX1 I_15581 (I267567,I2683,I267174,I267160,);
nor I_15582 (I267598,I267200,I267533);
DFFARX1 I_15583 (I267598,I2683,I267174,I267145,);
nor I_15584 (I267629,I267477,I267533);
not I_15585 (I267646,I267629);
nand I_15586 (I267154,I267646,I267502);
not I_15587 (I267701,I2690);
DFFARX1 I_15588 (I143765,I2683,I267701,I267727,);
not I_15589 (I267735,I267727);
nand I_15590 (I267752,I143762,I143771);
and I_15591 (I267769,I267752,I143780);
DFFARX1 I_15592 (I267769,I2683,I267701,I267795,);
DFFARX1 I_15593 (I267795,I2683,I267701,I267690,);
DFFARX1 I_15594 (I143783,I2683,I267701,I267826,);
nand I_15595 (I267834,I267826,I143786);
not I_15596 (I267851,I267834);
DFFARX1 I_15597 (I267851,I2683,I267701,I267877,);
not I_15598 (I267885,I267877);
nor I_15599 (I267693,I267735,I267885);
DFFARX1 I_15600 (I143759,I2683,I267701,I267925,);
nor I_15601 (I267684,I267925,I267795);
nor I_15602 (I267675,I267925,I267851);
nand I_15603 (I267961,I143774,I143777);
and I_15604 (I267978,I267961,I143768);
DFFARX1 I_15605 (I267978,I2683,I267701,I268004,);
not I_15606 (I268012,I268004);
nand I_15607 (I268029,I268012,I267925);
nand I_15608 (I267678,I268012,I267834);
nor I_15609 (I268060,I143759,I143777);
and I_15610 (I268077,I267925,I268060);
nor I_15611 (I268094,I268012,I268077);
DFFARX1 I_15612 (I268094,I2683,I267701,I267687,);
nor I_15613 (I268125,I267727,I268060);
DFFARX1 I_15614 (I268125,I2683,I267701,I267672,);
nor I_15615 (I268156,I268004,I268060);
not I_15616 (I268173,I268156);
nand I_15617 (I267681,I268173,I268029);
not I_15618 (I268228,I2690);
DFFARX1 I_15619 (I18867,I2683,I268228,I268254,);
not I_15620 (I268262,I268254);
nand I_15621 (I268279,I18843,I18852);
and I_15622 (I268296,I268279,I18846);
DFFARX1 I_15623 (I268296,I2683,I268228,I268322,);
DFFARX1 I_15624 (I268322,I2683,I268228,I268217,);
DFFARX1 I_15625 (I18864,I2683,I268228,I268353,);
nand I_15626 (I268361,I268353,I18855);
not I_15627 (I268378,I268361);
DFFARX1 I_15628 (I268378,I2683,I268228,I268404,);
not I_15629 (I268412,I268404);
nor I_15630 (I268220,I268262,I268412);
DFFARX1 I_15631 (I18849,I2683,I268228,I268452,);
nor I_15632 (I268211,I268452,I268322);
nor I_15633 (I268202,I268452,I268378);
nand I_15634 (I268488,I18861,I18858);
and I_15635 (I268505,I268488,I18846);
DFFARX1 I_15636 (I268505,I2683,I268228,I268531,);
not I_15637 (I268539,I268531);
nand I_15638 (I268556,I268539,I268452);
nand I_15639 (I268205,I268539,I268361);
nor I_15640 (I268587,I18843,I18858);
and I_15641 (I268604,I268452,I268587);
nor I_15642 (I268621,I268539,I268604);
DFFARX1 I_15643 (I268621,I2683,I268228,I268214,);
nor I_15644 (I268652,I268254,I268587);
DFFARX1 I_15645 (I268652,I2683,I268228,I268199,);
nor I_15646 (I268683,I268531,I268587);
not I_15647 (I268700,I268683);
nand I_15648 (I268208,I268700,I268556);
not I_15649 (I268755,I2690);
DFFARX1 I_15650 (I51285,I2683,I268755,I268781,);
not I_15651 (I268789,I268781);
nand I_15652 (I268806,I51282,I51300);
and I_15653 (I268823,I268806,I51291);
DFFARX1 I_15654 (I268823,I2683,I268755,I268849,);
DFFARX1 I_15655 (I268849,I2683,I268755,I268744,);
DFFARX1 I_15656 (I51297,I2683,I268755,I268880,);
nand I_15657 (I268888,I268880,I51294);
not I_15658 (I268905,I268888);
DFFARX1 I_15659 (I268905,I2683,I268755,I268931,);
not I_15660 (I268939,I268931);
nor I_15661 (I268747,I268789,I268939);
DFFARX1 I_15662 (I51288,I2683,I268755,I268979,);
nor I_15663 (I268738,I268979,I268849);
nor I_15664 (I268729,I268979,I268905);
nand I_15665 (I269015,I51279,I51303);
and I_15666 (I269032,I269015,I51282);
DFFARX1 I_15667 (I269032,I2683,I268755,I269058,);
not I_15668 (I269066,I269058);
nand I_15669 (I269083,I269066,I268979);
nand I_15670 (I268732,I269066,I268888);
nor I_15671 (I269114,I51279,I51303);
and I_15672 (I269131,I268979,I269114);
nor I_15673 (I269148,I269066,I269131);
DFFARX1 I_15674 (I269148,I2683,I268755,I268741,);
nor I_15675 (I269179,I268781,I269114);
DFFARX1 I_15676 (I269179,I2683,I268755,I268726,);
nor I_15677 (I269210,I269058,I269114);
not I_15678 (I269227,I269210);
nand I_15679 (I268735,I269227,I269083);
not I_15680 (I269282,I2690);
DFFARX1 I_15681 (I144309,I2683,I269282,I269308,);
not I_15682 (I269316,I269308);
nand I_15683 (I269333,I144306,I144315);
and I_15684 (I269350,I269333,I144324);
DFFARX1 I_15685 (I269350,I2683,I269282,I269376,);
DFFARX1 I_15686 (I269376,I2683,I269282,I269271,);
DFFARX1 I_15687 (I144327,I2683,I269282,I269407,);
nand I_15688 (I269415,I269407,I144330);
not I_15689 (I269432,I269415);
DFFARX1 I_15690 (I269432,I2683,I269282,I269458,);
not I_15691 (I269466,I269458);
nor I_15692 (I269274,I269316,I269466);
DFFARX1 I_15693 (I144303,I2683,I269282,I269506,);
nor I_15694 (I269265,I269506,I269376);
nor I_15695 (I269256,I269506,I269432);
nand I_15696 (I269542,I144318,I144321);
and I_15697 (I269559,I269542,I144312);
DFFARX1 I_15698 (I269559,I2683,I269282,I269585,);
not I_15699 (I269593,I269585);
nand I_15700 (I269610,I269593,I269506);
nand I_15701 (I269259,I269593,I269415);
nor I_15702 (I269641,I144303,I144321);
and I_15703 (I269658,I269506,I269641);
nor I_15704 (I269675,I269593,I269658);
DFFARX1 I_15705 (I269675,I2683,I269282,I269268,);
nor I_15706 (I269706,I269308,I269641);
DFFARX1 I_15707 (I269706,I2683,I269282,I269253,);
nor I_15708 (I269737,I269585,I269641);
not I_15709 (I269754,I269737);
nand I_15710 (I269262,I269754,I269610);
not I_15711 (I269815,I2690);
DFFARX1 I_15712 (I229071,I2683,I269815,I269841,);
DFFARX1 I_15713 (I229065,I2683,I269815,I269858,);
not I_15714 (I269866,I269858);
not I_15715 (I269883,I229080);
nor I_15716 (I269900,I269883,I229065);
not I_15717 (I269917,I229074);
nor I_15718 (I269934,I269900,I229083);
nor I_15719 (I269951,I269858,I269934);
DFFARX1 I_15720 (I269951,I2683,I269815,I269801,);
nor I_15721 (I269982,I229083,I229065);
nand I_15722 (I269999,I269982,I229080);
DFFARX1 I_15723 (I269999,I2683,I269815,I269804,);
nor I_15724 (I270030,I269917,I229083);
nand I_15725 (I270047,I270030,I229068);
nor I_15726 (I270064,I269841,I270047);
DFFARX1 I_15727 (I270064,I2683,I269815,I269780,);
not I_15728 (I270095,I270047);
nand I_15729 (I269792,I269858,I270095);
DFFARX1 I_15730 (I270047,I2683,I269815,I270135,);
not I_15731 (I270143,I270135);
not I_15732 (I270160,I229083);
not I_15733 (I270177,I229077);
nor I_15734 (I270194,I270177,I229074);
nor I_15735 (I269807,I270143,I270194);
nor I_15736 (I270225,I270177,I229086);
and I_15737 (I270242,I270225,I229089);
or I_15738 (I270259,I270242,I229068);
DFFARX1 I_15739 (I270259,I2683,I269815,I270285,);
nor I_15740 (I269795,I270285,I269841);
not I_15741 (I270307,I270285);
and I_15742 (I270324,I270307,I269841);
nor I_15743 (I269789,I269866,I270324);
nand I_15744 (I270355,I270307,I269917);
nor I_15745 (I269783,I270177,I270355);
nand I_15746 (I269786,I270307,I270095);
nand I_15747 (I270400,I269917,I229077);
nor I_15748 (I269798,I270160,I270400);
not I_15749 (I270461,I2690);
DFFARX1 I_15750 (I110031,I2683,I270461,I270487,);
DFFARX1 I_15751 (I110037,I2683,I270461,I270504,);
not I_15752 (I270512,I270504);
not I_15753 (I270529,I110058);
nor I_15754 (I270546,I270529,I110046);
not I_15755 (I270563,I110055);
nor I_15756 (I270580,I270546,I110040);
nor I_15757 (I270597,I270504,I270580);
DFFARX1 I_15758 (I270597,I2683,I270461,I270447,);
nor I_15759 (I270628,I110040,I110046);
nand I_15760 (I270645,I270628,I110058);
DFFARX1 I_15761 (I270645,I2683,I270461,I270450,);
nor I_15762 (I270676,I270563,I110040);
nand I_15763 (I270693,I270676,I110031);
nor I_15764 (I270710,I270487,I270693);
DFFARX1 I_15765 (I270710,I2683,I270461,I270426,);
not I_15766 (I270741,I270693);
nand I_15767 (I270438,I270504,I270741);
DFFARX1 I_15768 (I270693,I2683,I270461,I270781,);
not I_15769 (I270789,I270781);
not I_15770 (I270806,I110040);
not I_15771 (I270823,I110043);
nor I_15772 (I270840,I270823,I110055);
nor I_15773 (I270453,I270789,I270840);
nor I_15774 (I270871,I270823,I110052);
and I_15775 (I270888,I270871,I110034);
or I_15776 (I270905,I270888,I110049);
DFFARX1 I_15777 (I270905,I2683,I270461,I270931,);
nor I_15778 (I270441,I270931,I270487);
not I_15779 (I270953,I270931);
and I_15780 (I270970,I270953,I270487);
nor I_15781 (I270435,I270512,I270970);
nand I_15782 (I271001,I270953,I270563);
nor I_15783 (I270429,I270823,I271001);
nand I_15784 (I270432,I270953,I270741);
nand I_15785 (I271046,I270563,I110043);
nor I_15786 (I270444,I270806,I271046);
not I_15787 (I271107,I2690);
DFFARX1 I_15788 (I162377,I2683,I271107,I271133,);
DFFARX1 I_15789 (I162389,I2683,I271107,I271150,);
not I_15790 (I271158,I271150);
not I_15791 (I271175,I162374);
nor I_15792 (I271192,I271175,I162392);
not I_15793 (I271209,I162398);
nor I_15794 (I271226,I271192,I162380);
nor I_15795 (I271243,I271150,I271226);
DFFARX1 I_15796 (I271243,I2683,I271107,I271093,);
nor I_15797 (I271274,I162380,I162392);
nand I_15798 (I271291,I271274,I162374);
DFFARX1 I_15799 (I271291,I2683,I271107,I271096,);
nor I_15800 (I271322,I271209,I162380);
nand I_15801 (I271339,I271322,I162383);
nor I_15802 (I271356,I271133,I271339);
DFFARX1 I_15803 (I271356,I2683,I271107,I271072,);
not I_15804 (I271387,I271339);
nand I_15805 (I271084,I271150,I271387);
DFFARX1 I_15806 (I271339,I2683,I271107,I271427,);
not I_15807 (I271435,I271427);
not I_15808 (I271452,I162380);
not I_15809 (I271469,I162386);
nor I_15810 (I271486,I271469,I162398);
nor I_15811 (I271099,I271435,I271486);
nor I_15812 (I271517,I271469,I162395);
and I_15813 (I271534,I271517,I162374);
or I_15814 (I271551,I271534,I162377);
DFFARX1 I_15815 (I271551,I2683,I271107,I271577,);
nor I_15816 (I271087,I271577,I271133);
not I_15817 (I271599,I271577);
and I_15818 (I271616,I271599,I271133);
nor I_15819 (I271081,I271158,I271616);
nand I_15820 (I271647,I271599,I271209);
nor I_15821 (I271075,I271469,I271647);
nand I_15822 (I271078,I271599,I271387);
nand I_15823 (I271692,I271209,I162386);
nor I_15824 (I271090,I271452,I271692);
not I_15825 (I271753,I2690);
DFFARX1 I_15826 (I186296,I2683,I271753,I271779,);
DFFARX1 I_15827 (I186308,I2683,I271753,I271796,);
not I_15828 (I271804,I271796);
not I_15829 (I271821,I186317);
nor I_15830 (I271838,I271821,I186293);
not I_15831 (I271855,I186311);
nor I_15832 (I271872,I271838,I186305);
nor I_15833 (I271889,I271796,I271872);
DFFARX1 I_15834 (I271889,I2683,I271753,I271739,);
nor I_15835 (I271920,I186305,I186293);
nand I_15836 (I271937,I271920,I186317);
DFFARX1 I_15837 (I271937,I2683,I271753,I271742,);
nor I_15838 (I271968,I271855,I186305);
nand I_15839 (I271985,I271968,I186299);
nor I_15840 (I272002,I271779,I271985);
DFFARX1 I_15841 (I272002,I2683,I271753,I271718,);
not I_15842 (I272033,I271985);
nand I_15843 (I271730,I271796,I272033);
DFFARX1 I_15844 (I271985,I2683,I271753,I272073,);
not I_15845 (I272081,I272073);
not I_15846 (I272098,I186305);
not I_15847 (I272115,I186314);
nor I_15848 (I272132,I272115,I186311);
nor I_15849 (I271745,I272081,I272132);
nor I_15850 (I272163,I272115,I186296);
and I_15851 (I272180,I272163,I186293);
or I_15852 (I272197,I272180,I186302);
DFFARX1 I_15853 (I272197,I2683,I271753,I272223,);
nor I_15854 (I271733,I272223,I271779);
not I_15855 (I272245,I272223);
and I_15856 (I272262,I272245,I271779);
nor I_15857 (I271727,I271804,I272262);
nand I_15858 (I272293,I272245,I271855);
nor I_15859 (I271721,I272115,I272293);
nand I_15860 (I271724,I272245,I272033);
nand I_15861 (I272338,I271855,I186314);
nor I_15862 (I271736,I272098,I272338);
not I_15863 (I272399,I2690);
DFFARX1 I_15864 (I264516,I2683,I272399,I272425,);
DFFARX1 I_15865 (I264513,I2683,I272399,I272442,);
not I_15866 (I272450,I272442);
not I_15867 (I272467,I264513);
nor I_15868 (I272484,I272467,I264516);
not I_15869 (I272501,I264528);
nor I_15870 (I272518,I272484,I264522);
nor I_15871 (I272535,I272442,I272518);
DFFARX1 I_15872 (I272535,I2683,I272399,I272385,);
nor I_15873 (I272566,I264522,I264516);
nand I_15874 (I272583,I272566,I264513);
DFFARX1 I_15875 (I272583,I2683,I272399,I272388,);
nor I_15876 (I272614,I272501,I264522);
nand I_15877 (I272631,I272614,I264510);
nor I_15878 (I272648,I272425,I272631);
DFFARX1 I_15879 (I272648,I2683,I272399,I272364,);
not I_15880 (I272679,I272631);
nand I_15881 (I272376,I272442,I272679);
DFFARX1 I_15882 (I272631,I2683,I272399,I272719,);
not I_15883 (I272727,I272719);
not I_15884 (I272744,I264522);
not I_15885 (I272761,I264519);
nor I_15886 (I272778,I272761,I264528);
nor I_15887 (I272391,I272727,I272778);
nor I_15888 (I272809,I272761,I264525);
and I_15889 (I272826,I272809,I264531);
or I_15890 (I272843,I272826,I264510);
DFFARX1 I_15891 (I272843,I2683,I272399,I272869,);
nor I_15892 (I272379,I272869,I272425);
not I_15893 (I272891,I272869);
and I_15894 (I272908,I272891,I272425);
nor I_15895 (I272373,I272450,I272908);
nand I_15896 (I272939,I272891,I272501);
nor I_15897 (I272367,I272761,I272939);
nand I_15898 (I272370,I272891,I272679);
nand I_15899 (I272984,I272501,I264519);
nor I_15900 (I272382,I272744,I272984);
not I_15901 (I273045,I2690);
DFFARX1 I_15902 (I334279,I2683,I273045,I273071,);
DFFARX1 I_15903 (I334261,I2683,I273045,I273088,);
not I_15904 (I273096,I273088);
not I_15905 (I273113,I334270);
nor I_15906 (I273130,I273113,I334282);
not I_15907 (I273147,I334264);
nor I_15908 (I273164,I273130,I334273);
nor I_15909 (I273181,I273088,I273164);
DFFARX1 I_15910 (I273181,I2683,I273045,I273031,);
nor I_15911 (I273212,I334273,I334282);
nand I_15912 (I273229,I273212,I334270);
DFFARX1 I_15913 (I273229,I2683,I273045,I273034,);
nor I_15914 (I273260,I273147,I334273);
nand I_15915 (I273277,I273260,I334285);
nor I_15916 (I273294,I273071,I273277);
DFFARX1 I_15917 (I273294,I2683,I273045,I273010,);
not I_15918 (I273325,I273277);
nand I_15919 (I273022,I273088,I273325);
DFFARX1 I_15920 (I273277,I2683,I273045,I273365,);
not I_15921 (I273373,I273365);
not I_15922 (I273390,I334273);
not I_15923 (I273407,I334261);
nor I_15924 (I273424,I273407,I334264);
nor I_15925 (I273037,I273373,I273424);
nor I_15926 (I273455,I273407,I334267);
and I_15927 (I273472,I273455,I334276);
or I_15928 (I273489,I273472,I334264);
DFFARX1 I_15929 (I273489,I2683,I273045,I273515,);
nor I_15930 (I273025,I273515,I273071);
not I_15931 (I273537,I273515);
and I_15932 (I273554,I273537,I273071);
nor I_15933 (I273019,I273096,I273554);
nand I_15934 (I273585,I273537,I273147);
nor I_15935 (I273013,I273407,I273585);
nand I_15936 (I273016,I273537,I273325);
nand I_15937 (I273630,I273147,I334261);
nor I_15938 (I273028,I273390,I273630);
not I_15939 (I273691,I2690);
DFFARX1 I_15940 (I120044,I2683,I273691,I273717,);
DFFARX1 I_15941 (I120050,I2683,I273691,I273734,);
not I_15942 (I273742,I273734);
not I_15943 (I273759,I120071);
nor I_15944 (I273776,I273759,I120059);
not I_15945 (I273793,I120068);
nor I_15946 (I273810,I273776,I120053);
nor I_15947 (I273827,I273734,I273810);
DFFARX1 I_15948 (I273827,I2683,I273691,I273677,);
nor I_15949 (I273858,I120053,I120059);
nand I_15950 (I273875,I273858,I120071);
DFFARX1 I_15951 (I273875,I2683,I273691,I273680,);
nor I_15952 (I273906,I273793,I120053);
nand I_15953 (I273923,I273906,I120044);
nor I_15954 (I273940,I273717,I273923);
DFFARX1 I_15955 (I273940,I2683,I273691,I273656,);
not I_15956 (I273971,I273923);
nand I_15957 (I273668,I273734,I273971);
DFFARX1 I_15958 (I273923,I2683,I273691,I274011,);
not I_15959 (I274019,I274011);
not I_15960 (I274036,I120053);
not I_15961 (I274053,I120056);
nor I_15962 (I274070,I274053,I120068);
nor I_15963 (I273683,I274019,I274070);
nor I_15964 (I274101,I274053,I120065);
and I_15965 (I274118,I274101,I120047);
or I_15966 (I274135,I274118,I120062);
DFFARX1 I_15967 (I274135,I2683,I273691,I274161,);
nor I_15968 (I273671,I274161,I273717);
not I_15969 (I274183,I274161);
and I_15970 (I274200,I274183,I273717);
nor I_15971 (I273665,I273742,I274200);
nand I_15972 (I274231,I274183,I273793);
nor I_15973 (I273659,I274053,I274231);
nand I_15974 (I273662,I274183,I273971);
nand I_15975 (I274276,I273793,I120056);
nor I_15976 (I273674,I274036,I274276);
not I_15977 (I274337,I2690);
DFFARX1 I_15978 (I189186,I2683,I274337,I274363,);
DFFARX1 I_15979 (I189198,I2683,I274337,I274380,);
not I_15980 (I274388,I274380);
not I_15981 (I274405,I189207);
nor I_15982 (I274422,I274405,I189183);
not I_15983 (I274439,I189201);
nor I_15984 (I274456,I274422,I189195);
nor I_15985 (I274473,I274380,I274456);
DFFARX1 I_15986 (I274473,I2683,I274337,I274323,);
nor I_15987 (I274504,I189195,I189183);
nand I_15988 (I274521,I274504,I189207);
DFFARX1 I_15989 (I274521,I2683,I274337,I274326,);
nor I_15990 (I274552,I274439,I189195);
nand I_15991 (I274569,I274552,I189189);
nor I_15992 (I274586,I274363,I274569);
DFFARX1 I_15993 (I274586,I2683,I274337,I274302,);
not I_15994 (I274617,I274569);
nand I_15995 (I274314,I274380,I274617);
DFFARX1 I_15996 (I274569,I2683,I274337,I274657,);
not I_15997 (I274665,I274657);
not I_15998 (I274682,I189195);
not I_15999 (I274699,I189204);
nor I_16000 (I274716,I274699,I189201);
nor I_16001 (I274329,I274665,I274716);
nor I_16002 (I274747,I274699,I189186);
and I_16003 (I274764,I274747,I189183);
or I_16004 (I274781,I274764,I189192);
DFFARX1 I_16005 (I274781,I2683,I274337,I274807,);
nor I_16006 (I274317,I274807,I274363);
not I_16007 (I274829,I274807);
and I_16008 (I274846,I274829,I274363);
nor I_16009 (I274311,I274388,I274846);
nand I_16010 (I274877,I274829,I274439);
nor I_16011 (I274305,I274699,I274877);
nand I_16012 (I274308,I274829,I274617);
nand I_16013 (I274922,I274439,I189204);
nor I_16014 (I274320,I274682,I274922);
not I_16015 (I274983,I2690);
DFFARX1 I_16016 (I162972,I2683,I274983,I275009,);
DFFARX1 I_16017 (I162984,I2683,I274983,I275026,);
not I_16018 (I275034,I275026);
not I_16019 (I275051,I162969);
nor I_16020 (I275068,I275051,I162987);
not I_16021 (I275085,I162993);
nor I_16022 (I275102,I275068,I162975);
nor I_16023 (I275119,I275026,I275102);
DFFARX1 I_16024 (I275119,I2683,I274983,I274969,);
nor I_16025 (I275150,I162975,I162987);
nand I_16026 (I275167,I275150,I162969);
DFFARX1 I_16027 (I275167,I2683,I274983,I274972,);
nor I_16028 (I275198,I275085,I162975);
nand I_16029 (I275215,I275198,I162978);
nor I_16030 (I275232,I275009,I275215);
DFFARX1 I_16031 (I275232,I2683,I274983,I274948,);
not I_16032 (I275263,I275215);
nand I_16033 (I274960,I275026,I275263);
DFFARX1 I_16034 (I275215,I2683,I274983,I275303,);
not I_16035 (I275311,I275303);
not I_16036 (I275328,I162975);
not I_16037 (I275345,I162981);
nor I_16038 (I275362,I275345,I162993);
nor I_16039 (I274975,I275311,I275362);
nor I_16040 (I275393,I275345,I162990);
and I_16041 (I275410,I275393,I162969);
or I_16042 (I275427,I275410,I162972);
DFFARX1 I_16043 (I275427,I2683,I274983,I275453,);
nor I_16044 (I274963,I275453,I275009);
not I_16045 (I275475,I275453);
and I_16046 (I275492,I275475,I275009);
nor I_16047 (I274957,I275034,I275492);
nand I_16048 (I275523,I275475,I275085);
nor I_16049 (I274951,I275345,I275523);
nand I_16050 (I274954,I275475,I275263);
nand I_16051 (I275568,I275085,I162981);
nor I_16052 (I274966,I275328,I275568);
not I_16053 (I275629,I2690);
DFFARX1 I_16054 (I403944,I2683,I275629,I275655,);
DFFARX1 I_16055 (I403968,I2683,I275629,I275672,);
not I_16056 (I275680,I275672);
not I_16057 (I275697,I403950);
nor I_16058 (I275714,I275697,I403959);
not I_16059 (I275731,I403944);
nor I_16060 (I275748,I275714,I403965);
nor I_16061 (I275765,I275672,I275748);
DFFARX1 I_16062 (I275765,I2683,I275629,I275615,);
nor I_16063 (I275796,I403965,I403959);
nand I_16064 (I275813,I275796,I403950);
DFFARX1 I_16065 (I275813,I2683,I275629,I275618,);
nor I_16066 (I275844,I275731,I403965);
nand I_16067 (I275861,I275844,I403962);
nor I_16068 (I275878,I275655,I275861);
DFFARX1 I_16069 (I275878,I2683,I275629,I275594,);
not I_16070 (I275909,I275861);
nand I_16071 (I275606,I275672,I275909);
DFFARX1 I_16072 (I275861,I2683,I275629,I275949,);
not I_16073 (I275957,I275949);
not I_16074 (I275974,I403965);
not I_16075 (I275991,I403956);
nor I_16076 (I276008,I275991,I403944);
nor I_16077 (I275621,I275957,I276008);
nor I_16078 (I276039,I275991,I403947);
and I_16079 (I276056,I276039,I403971);
or I_16080 (I276073,I276056,I403953);
DFFARX1 I_16081 (I276073,I2683,I275629,I276099,);
nor I_16082 (I275609,I276099,I275655);
not I_16083 (I276121,I276099);
and I_16084 (I276138,I276121,I275655);
nor I_16085 (I275603,I275680,I276138);
nand I_16086 (I276169,I276121,I275731);
nor I_16087 (I275597,I275991,I276169);
nand I_16088 (I275600,I276121,I275909);
nand I_16089 (I276214,I275731,I403956);
nor I_16090 (I275612,I275974,I276214);
not I_16091 (I276275,I2690);
DFFARX1 I_16092 (I9884,I2683,I276275,I276301,);
DFFARX1 I_16093 (I9890,I2683,I276275,I276318,);
not I_16094 (I276326,I276318);
not I_16095 (I276343,I9884);
nor I_16096 (I276360,I276343,I9896);
not I_16097 (I276377,I9908);
nor I_16098 (I276394,I276360,I9902);
nor I_16099 (I276411,I276318,I276394);
DFFARX1 I_16100 (I276411,I2683,I276275,I276261,);
nor I_16101 (I276442,I9902,I9896);
nand I_16102 (I276459,I276442,I9884);
DFFARX1 I_16103 (I276459,I2683,I276275,I276264,);
nor I_16104 (I276490,I276377,I9902);
nand I_16105 (I276507,I276490,I9887);
nor I_16106 (I276524,I276301,I276507);
DFFARX1 I_16107 (I276524,I2683,I276275,I276240,);
not I_16108 (I276555,I276507);
nand I_16109 (I276252,I276318,I276555);
DFFARX1 I_16110 (I276507,I2683,I276275,I276595,);
not I_16111 (I276603,I276595);
not I_16112 (I276620,I9902);
not I_16113 (I276637,I9887);
nor I_16114 (I276654,I276637,I9908);
nor I_16115 (I276267,I276603,I276654);
nor I_16116 (I276685,I276637,I9905);
and I_16117 (I276702,I276685,I9899);
or I_16118 (I276719,I276702,I9893);
DFFARX1 I_16119 (I276719,I2683,I276275,I276745,);
nor I_16120 (I276255,I276745,I276301);
not I_16121 (I276767,I276745);
and I_16122 (I276784,I276767,I276301);
nor I_16123 (I276249,I276326,I276784);
nand I_16124 (I276815,I276767,I276377);
nor I_16125 (I276243,I276637,I276815);
nand I_16126 (I276246,I276767,I276555);
nand I_16127 (I276860,I276377,I9887);
nor I_16128 (I276258,I276620,I276860);
not I_16129 (I276921,I2690);
DFFARX1 I_16130 (I96329,I2683,I276921,I276947,);
DFFARX1 I_16131 (I96335,I2683,I276921,I276964,);
not I_16132 (I276972,I276964);
not I_16133 (I276989,I96356);
nor I_16134 (I277006,I276989,I96344);
not I_16135 (I277023,I96353);
nor I_16136 (I277040,I277006,I96338);
nor I_16137 (I277057,I276964,I277040);
DFFARX1 I_16138 (I277057,I2683,I276921,I276907,);
nor I_16139 (I277088,I96338,I96344);
nand I_16140 (I277105,I277088,I96356);
DFFARX1 I_16141 (I277105,I2683,I276921,I276910,);
nor I_16142 (I277136,I277023,I96338);
nand I_16143 (I277153,I277136,I96329);
nor I_16144 (I277170,I276947,I277153);
DFFARX1 I_16145 (I277170,I2683,I276921,I276886,);
not I_16146 (I277201,I277153);
nand I_16147 (I276898,I276964,I277201);
DFFARX1 I_16148 (I277153,I2683,I276921,I277241,);
not I_16149 (I277249,I277241);
not I_16150 (I277266,I96338);
not I_16151 (I277283,I96341);
nor I_16152 (I277300,I277283,I96353);
nor I_16153 (I276913,I277249,I277300);
nor I_16154 (I277331,I277283,I96350);
and I_16155 (I277348,I277331,I96332);
or I_16156 (I277365,I277348,I96347);
DFFARX1 I_16157 (I277365,I2683,I276921,I277391,);
nor I_16158 (I276901,I277391,I276947);
not I_16159 (I277413,I277391);
and I_16160 (I277430,I277413,I276947);
nor I_16161 (I276895,I276972,I277430);
nand I_16162 (I277461,I277413,I277023);
nor I_16163 (I276889,I277283,I277461);
nand I_16164 (I276892,I277413,I277201);
nand I_16165 (I277506,I277023,I96341);
nor I_16166 (I276904,I277266,I277506);
not I_16167 (I277567,I2690);
DFFARX1 I_16168 (I129621,I2683,I277567,I277593,);
DFFARX1 I_16169 (I129618,I2683,I277567,I277610,);
not I_16170 (I277618,I277610);
not I_16171 (I277635,I129633);
nor I_16172 (I277652,I277635,I129636);
not I_16173 (I277669,I129624);
nor I_16174 (I277686,I277652,I129630);
nor I_16175 (I277703,I277610,I277686);
DFFARX1 I_16176 (I277703,I2683,I277567,I277553,);
nor I_16177 (I277734,I129630,I129636);
nand I_16178 (I277751,I277734,I129633);
DFFARX1 I_16179 (I277751,I2683,I277567,I277556,);
nor I_16180 (I277782,I277669,I129630);
nand I_16181 (I277799,I277782,I129642);
nor I_16182 (I277816,I277593,I277799);
DFFARX1 I_16183 (I277816,I2683,I277567,I277532,);
not I_16184 (I277847,I277799);
nand I_16185 (I277544,I277610,I277847);
DFFARX1 I_16186 (I277799,I2683,I277567,I277887,);
not I_16187 (I277895,I277887);
not I_16188 (I277912,I129630);
not I_16189 (I277929,I129615);
nor I_16190 (I277946,I277929,I129624);
nor I_16191 (I277559,I277895,I277946);
nor I_16192 (I277977,I277929,I129627);
and I_16193 (I277994,I277977,I129615);
or I_16194 (I278011,I277994,I129639);
DFFARX1 I_16195 (I278011,I2683,I277567,I278037,);
nor I_16196 (I277547,I278037,I277593);
not I_16197 (I278059,I278037);
and I_16198 (I278076,I278059,I277593);
nor I_16199 (I277541,I277618,I278076);
nand I_16200 (I278107,I278059,I277669);
nor I_16201 (I277535,I277929,I278107);
nand I_16202 (I277538,I278059,I277847);
nand I_16203 (I278152,I277669,I129615);
nor I_16204 (I277550,I277912,I278152);
not I_16205 (I278213,I2690);
DFFARX1 I_16206 (I22005,I2683,I278213,I278239,);
DFFARX1 I_16207 (I22011,I2683,I278213,I278256,);
not I_16208 (I278264,I278256);
not I_16209 (I278281,I22029);
nor I_16210 (I278298,I278281,I22008);
not I_16211 (I278315,I22014);
nor I_16212 (I278332,I278298,I22020);
nor I_16213 (I278349,I278256,I278332);
DFFARX1 I_16214 (I278349,I2683,I278213,I278199,);
nor I_16215 (I278380,I22020,I22008);
nand I_16216 (I278397,I278380,I22029);
DFFARX1 I_16217 (I278397,I2683,I278213,I278202,);
nor I_16218 (I278428,I278315,I22020);
nand I_16219 (I278445,I278428,I22026);
nor I_16220 (I278462,I278239,I278445);
DFFARX1 I_16221 (I278462,I2683,I278213,I278178,);
not I_16222 (I278493,I278445);
nand I_16223 (I278190,I278256,I278493);
DFFARX1 I_16224 (I278445,I2683,I278213,I278533,);
not I_16225 (I278541,I278533);
not I_16226 (I278558,I22020);
not I_16227 (I278575,I22008);
nor I_16228 (I278592,I278575,I22014);
nor I_16229 (I278205,I278541,I278592);
nor I_16230 (I278623,I278575,I22017);
and I_16231 (I278640,I278623,I22005);
or I_16232 (I278657,I278640,I22023);
DFFARX1 I_16233 (I278657,I2683,I278213,I278683,);
nor I_16234 (I278193,I278683,I278239);
not I_16235 (I278705,I278683);
and I_16236 (I278722,I278705,I278239);
nor I_16237 (I278187,I278264,I278722);
nand I_16238 (I278753,I278705,I278315);
nor I_16239 (I278181,I278575,I278753);
nand I_16240 (I278184,I278705,I278493);
nand I_16241 (I278798,I278315,I22008);
nor I_16242 (I278196,I278558,I278798);
not I_16243 (I278859,I2690);
DFFARX1 I_16244 (I201905,I2683,I278859,I278885,);
DFFARX1 I_16245 (I201899,I2683,I278859,I278902,);
not I_16246 (I278910,I278902);
not I_16247 (I278927,I201914);
nor I_16248 (I278944,I278927,I201899);
not I_16249 (I278961,I201908);
nor I_16250 (I278978,I278944,I201917);
nor I_16251 (I278995,I278902,I278978);
DFFARX1 I_16252 (I278995,I2683,I278859,I278845,);
nor I_16253 (I279026,I201917,I201899);
nand I_16254 (I279043,I279026,I201914);
DFFARX1 I_16255 (I279043,I2683,I278859,I278848,);
nor I_16256 (I279074,I278961,I201917);
nand I_16257 (I279091,I279074,I201902);
nor I_16258 (I279108,I278885,I279091);
DFFARX1 I_16259 (I279108,I2683,I278859,I278824,);
not I_16260 (I279139,I279091);
nand I_16261 (I278836,I278902,I279139);
DFFARX1 I_16262 (I279091,I2683,I278859,I279179,);
not I_16263 (I279187,I279179);
not I_16264 (I279204,I201917);
not I_16265 (I279221,I201911);
nor I_16266 (I279238,I279221,I201908);
nor I_16267 (I278851,I279187,I279238);
nor I_16268 (I279269,I279221,I201920);
and I_16269 (I279286,I279269,I201923);
or I_16270 (I279303,I279286,I201902);
DFFARX1 I_16271 (I279303,I2683,I278859,I279329,);
nor I_16272 (I278839,I279329,I278885);
not I_16273 (I279351,I279329);
and I_16274 (I279368,I279351,I278885);
nor I_16275 (I278833,I278910,I279368);
nand I_16276 (I279399,I279351,I278961);
nor I_16277 (I278827,I279221,I279399);
nand I_16278 (I278830,I279351,I279139);
nand I_16279 (I279444,I278961,I201911);
nor I_16280 (I278842,I279204,I279444);
not I_16281 (I279505,I2690);
DFFARX1 I_16282 (I98964,I2683,I279505,I279531,);
DFFARX1 I_16283 (I98970,I2683,I279505,I279548,);
not I_16284 (I279556,I279548);
not I_16285 (I279573,I98991);
nor I_16286 (I279590,I279573,I98979);
not I_16287 (I279607,I98988);
nor I_16288 (I279624,I279590,I98973);
nor I_16289 (I279641,I279548,I279624);
DFFARX1 I_16290 (I279641,I2683,I279505,I279491,);
nor I_16291 (I279672,I98973,I98979);
nand I_16292 (I279689,I279672,I98991);
DFFARX1 I_16293 (I279689,I2683,I279505,I279494,);
nor I_16294 (I279720,I279607,I98973);
nand I_16295 (I279737,I279720,I98964);
nor I_16296 (I279754,I279531,I279737);
DFFARX1 I_16297 (I279754,I2683,I279505,I279470,);
not I_16298 (I279785,I279737);
nand I_16299 (I279482,I279548,I279785);
DFFARX1 I_16300 (I279737,I2683,I279505,I279825,);
not I_16301 (I279833,I279825);
not I_16302 (I279850,I98973);
not I_16303 (I279867,I98976);
nor I_16304 (I279884,I279867,I98988);
nor I_16305 (I279497,I279833,I279884);
nor I_16306 (I279915,I279867,I98985);
and I_16307 (I279932,I279915,I98967);
or I_16308 (I279949,I279932,I98982);
DFFARX1 I_16309 (I279949,I2683,I279505,I279975,);
nor I_16310 (I279485,I279975,I279531);
not I_16311 (I279997,I279975);
and I_16312 (I280014,I279997,I279531);
nor I_16313 (I279479,I279556,I280014);
nand I_16314 (I280045,I279997,I279607);
nor I_16315 (I279473,I279867,I280045);
nand I_16316 (I279476,I279997,I279785);
nand I_16317 (I280090,I279607,I98976);
nor I_16318 (I279488,I279850,I280090);
not I_16319 (I280151,I2690);
DFFARX1 I_16320 (I49500,I2683,I280151,I280177,);
DFFARX1 I_16321 (I49512,I2683,I280151,I280194,);
not I_16322 (I280202,I280194);
not I_16323 (I280219,I49518);
nor I_16324 (I280236,I280219,I49503);
not I_16325 (I280253,I49494);
nor I_16326 (I280270,I280236,I49515);
nor I_16327 (I280287,I280194,I280270);
DFFARX1 I_16328 (I280287,I2683,I280151,I280137,);
nor I_16329 (I280318,I49515,I49503);
nand I_16330 (I280335,I280318,I49518);
DFFARX1 I_16331 (I280335,I2683,I280151,I280140,);
nor I_16332 (I280366,I280253,I49515);
nand I_16333 (I280383,I280366,I49497);
nor I_16334 (I280400,I280177,I280383);
DFFARX1 I_16335 (I280400,I2683,I280151,I280116,);
not I_16336 (I280431,I280383);
nand I_16337 (I280128,I280194,I280431);
DFFARX1 I_16338 (I280383,I2683,I280151,I280471,);
not I_16339 (I280479,I280471);
not I_16340 (I280496,I49515);
not I_16341 (I280513,I49506);
nor I_16342 (I280530,I280513,I49494);
nor I_16343 (I280143,I280479,I280530);
nor I_16344 (I280561,I280513,I49509);
and I_16345 (I280578,I280561,I49497);
or I_16346 (I280595,I280578,I49494);
DFFARX1 I_16347 (I280595,I2683,I280151,I280621,);
nor I_16348 (I280131,I280621,I280177);
not I_16349 (I280643,I280621);
and I_16350 (I280660,I280643,I280177);
nor I_16351 (I280125,I280202,I280660);
nand I_16352 (I280691,I280643,I280253);
nor I_16353 (I280119,I280513,I280691);
nand I_16354 (I280122,I280643,I280431);
nand I_16355 (I280736,I280253,I49506);
nor I_16356 (I280134,I280496,I280736);
not I_16357 (I280797,I2690);
DFFARX1 I_16358 (I378479,I2683,I280797,I280823,);
DFFARX1 I_16359 (I378485,I2683,I280797,I280840,);
not I_16360 (I280848,I280840);
not I_16361 (I280865,I378482);
nor I_16362 (I280882,I280865,I378461);
not I_16363 (I280899,I378464);
nor I_16364 (I280916,I280882,I378470);
nor I_16365 (I280933,I280840,I280916);
DFFARX1 I_16366 (I280933,I2683,I280797,I280783,);
nor I_16367 (I280964,I378470,I378461);
nand I_16368 (I280981,I280964,I378482);
DFFARX1 I_16369 (I280981,I2683,I280797,I280786,);
nor I_16370 (I281012,I280899,I378470);
nand I_16371 (I281029,I281012,I378464);
nor I_16372 (I281046,I280823,I281029);
DFFARX1 I_16373 (I281046,I2683,I280797,I280762,);
not I_16374 (I281077,I281029);
nand I_16375 (I280774,I280840,I281077);
DFFARX1 I_16376 (I281029,I2683,I280797,I281117,);
not I_16377 (I281125,I281117);
not I_16378 (I281142,I378470);
not I_16379 (I281159,I378473);
nor I_16380 (I281176,I281159,I378464);
nor I_16381 (I280789,I281125,I281176);
nor I_16382 (I281207,I281159,I378461);
and I_16383 (I281224,I281207,I378467);
or I_16384 (I281241,I281224,I378476);
DFFARX1 I_16385 (I281241,I2683,I280797,I281267,);
nor I_16386 (I280777,I281267,I280823);
not I_16387 (I281289,I281267);
and I_16388 (I281306,I281289,I280823);
nor I_16389 (I280771,I280848,I281306);
nand I_16390 (I281337,I281289,I280899);
nor I_16391 (I280765,I281159,I281337);
nand I_16392 (I280768,I281289,I281077);
nand I_16393 (I281382,I280899,I378473);
nor I_16394 (I280780,I281142,I281382);
not I_16395 (I281443,I2690);
DFFARX1 I_16396 (I259246,I2683,I281443,I281469,);
DFFARX1 I_16397 (I259243,I2683,I281443,I281486,);
not I_16398 (I281494,I281486);
not I_16399 (I281511,I259243);
nor I_16400 (I281528,I281511,I259246);
not I_16401 (I281545,I259258);
nor I_16402 (I281562,I281528,I259252);
nor I_16403 (I281579,I281486,I281562);
DFFARX1 I_16404 (I281579,I2683,I281443,I281429,);
nor I_16405 (I281610,I259252,I259246);
nand I_16406 (I281627,I281610,I259243);
DFFARX1 I_16407 (I281627,I2683,I281443,I281432,);
nor I_16408 (I281658,I281545,I259252);
nand I_16409 (I281675,I281658,I259240);
nor I_16410 (I281692,I281469,I281675);
DFFARX1 I_16411 (I281692,I2683,I281443,I281408,);
not I_16412 (I281723,I281675);
nand I_16413 (I281420,I281486,I281723);
DFFARX1 I_16414 (I281675,I2683,I281443,I281763,);
not I_16415 (I281771,I281763);
not I_16416 (I281788,I259252);
not I_16417 (I281805,I259249);
nor I_16418 (I281822,I281805,I259258);
nor I_16419 (I281435,I281771,I281822);
nor I_16420 (I281853,I281805,I259255);
and I_16421 (I281870,I281853,I259261);
or I_16422 (I281887,I281870,I259240);
DFFARX1 I_16423 (I281887,I2683,I281443,I281913,);
nor I_16424 (I281423,I281913,I281469);
not I_16425 (I281935,I281913);
and I_16426 (I281952,I281935,I281469);
nor I_16427 (I281417,I281494,I281952);
nand I_16428 (I281983,I281935,I281545);
nor I_16429 (I281411,I281805,I281983);
nand I_16430 (I281414,I281935,I281723);
nand I_16431 (I282028,I281545,I259249);
nor I_16432 (I281426,I281788,I282028);
not I_16433 (I282089,I2690);
DFFARX1 I_16434 (I121625,I2683,I282089,I282115,);
DFFARX1 I_16435 (I121631,I2683,I282089,I282132,);
not I_16436 (I282140,I282132);
not I_16437 (I282157,I121652);
nor I_16438 (I282174,I282157,I121640);
not I_16439 (I282191,I121649);
nor I_16440 (I282208,I282174,I121634);
nor I_16441 (I282225,I282132,I282208);
DFFARX1 I_16442 (I282225,I2683,I282089,I282075,);
nor I_16443 (I282256,I121634,I121640);
nand I_16444 (I282273,I282256,I121652);
DFFARX1 I_16445 (I282273,I2683,I282089,I282078,);
nor I_16446 (I282304,I282191,I121634);
nand I_16447 (I282321,I282304,I121625);
nor I_16448 (I282338,I282115,I282321);
DFFARX1 I_16449 (I282338,I2683,I282089,I282054,);
not I_16450 (I282369,I282321);
nand I_16451 (I282066,I282132,I282369);
DFFARX1 I_16452 (I282321,I2683,I282089,I282409,);
not I_16453 (I282417,I282409);
not I_16454 (I282434,I121634);
not I_16455 (I282451,I121637);
nor I_16456 (I282468,I282451,I121649);
nor I_16457 (I282081,I282417,I282468);
nor I_16458 (I282499,I282451,I121646);
and I_16459 (I282516,I282499,I121628);
or I_16460 (I282533,I282516,I121643);
DFFARX1 I_16461 (I282533,I2683,I282089,I282559,);
nor I_16462 (I282069,I282559,I282115);
not I_16463 (I282581,I282559);
and I_16464 (I282598,I282581,I282115);
nor I_16465 (I282063,I282140,I282598);
nand I_16466 (I282629,I282581,I282191);
nor I_16467 (I282057,I282451,I282629);
nand I_16468 (I282060,I282581,I282369);
nand I_16469 (I282674,I282191,I121637);
nor I_16470 (I282072,I282434,I282674);
not I_16471 (I282735,I2690);
DFFARX1 I_16472 (I95275,I2683,I282735,I282761,);
DFFARX1 I_16473 (I95281,I2683,I282735,I282778,);
not I_16474 (I282786,I282778);
not I_16475 (I282803,I95302);
nor I_16476 (I282820,I282803,I95290);
not I_16477 (I282837,I95299);
nor I_16478 (I282854,I282820,I95284);
nor I_16479 (I282871,I282778,I282854);
DFFARX1 I_16480 (I282871,I2683,I282735,I282721,);
nor I_16481 (I282902,I95284,I95290);
nand I_16482 (I282919,I282902,I95302);
DFFARX1 I_16483 (I282919,I2683,I282735,I282724,);
nor I_16484 (I282950,I282837,I95284);
nand I_16485 (I282967,I282950,I95275);
nor I_16486 (I282984,I282761,I282967);
DFFARX1 I_16487 (I282984,I2683,I282735,I282700,);
not I_16488 (I283015,I282967);
nand I_16489 (I282712,I282778,I283015);
DFFARX1 I_16490 (I282967,I2683,I282735,I283055,);
not I_16491 (I283063,I283055);
not I_16492 (I283080,I95284);
not I_16493 (I283097,I95287);
nor I_16494 (I283114,I283097,I95299);
nor I_16495 (I282727,I283063,I283114);
nor I_16496 (I283145,I283097,I95296);
and I_16497 (I283162,I283145,I95278);
or I_16498 (I283179,I283162,I95293);
DFFARX1 I_16499 (I283179,I2683,I282735,I283205,);
nor I_16500 (I282715,I283205,I282761);
not I_16501 (I283227,I283205);
and I_16502 (I283244,I283227,I282761);
nor I_16503 (I282709,I282786,I283244);
nand I_16504 (I283275,I283227,I282837);
nor I_16505 (I282703,I283097,I283275);
nand I_16506 (I282706,I283227,I283015);
nand I_16507 (I283320,I282837,I95287);
nor I_16508 (I282718,I283080,I283320);
not I_16509 (I283381,I2690);
DFFARX1 I_16510 (I96856,I2683,I283381,I283407,);
DFFARX1 I_16511 (I96862,I2683,I283381,I283424,);
not I_16512 (I283432,I283424);
not I_16513 (I283449,I96883);
nor I_16514 (I283466,I283449,I96871);
not I_16515 (I283483,I96880);
nor I_16516 (I283500,I283466,I96865);
nor I_16517 (I283517,I283424,I283500);
DFFARX1 I_16518 (I283517,I2683,I283381,I283367,);
nor I_16519 (I283548,I96865,I96871);
nand I_16520 (I283565,I283548,I96883);
DFFARX1 I_16521 (I283565,I2683,I283381,I283370,);
nor I_16522 (I283596,I283483,I96865);
nand I_16523 (I283613,I283596,I96856);
nor I_16524 (I283630,I283407,I283613);
DFFARX1 I_16525 (I283630,I2683,I283381,I283346,);
not I_16526 (I283661,I283613);
nand I_16527 (I283358,I283424,I283661);
DFFARX1 I_16528 (I283613,I2683,I283381,I283701,);
not I_16529 (I283709,I283701);
not I_16530 (I283726,I96865);
not I_16531 (I283743,I96868);
nor I_16532 (I283760,I283743,I96880);
nor I_16533 (I283373,I283709,I283760);
nor I_16534 (I283791,I283743,I96877);
and I_16535 (I283808,I283791,I96859);
or I_16536 (I283825,I283808,I96874);
DFFARX1 I_16537 (I283825,I2683,I283381,I283851,);
nor I_16538 (I283361,I283851,I283407);
not I_16539 (I283873,I283851);
and I_16540 (I283890,I283873,I283407);
nor I_16541 (I283355,I283432,I283890);
nand I_16542 (I283921,I283873,I283483);
nor I_16543 (I283349,I283743,I283921);
nand I_16544 (I283352,I283873,I283661);
nand I_16545 (I283966,I283483,I96868);
nor I_16546 (I283364,I283726,I283966);
not I_16547 (I284027,I2690);
DFFARX1 I_16548 (I368143,I2683,I284027,I284053,);
DFFARX1 I_16549 (I368149,I2683,I284027,I284070,);
not I_16550 (I284078,I284070);
not I_16551 (I284095,I368146);
nor I_16552 (I284112,I284095,I368125);
not I_16553 (I284129,I368128);
nor I_16554 (I284146,I284112,I368134);
nor I_16555 (I284163,I284070,I284146);
DFFARX1 I_16556 (I284163,I2683,I284027,I284013,);
nor I_16557 (I284194,I368134,I368125);
nand I_16558 (I284211,I284194,I368146);
DFFARX1 I_16559 (I284211,I2683,I284027,I284016,);
nor I_16560 (I284242,I284129,I368134);
nand I_16561 (I284259,I284242,I368128);
nor I_16562 (I284276,I284053,I284259);
DFFARX1 I_16563 (I284276,I2683,I284027,I283992,);
not I_16564 (I284307,I284259);
nand I_16565 (I284004,I284070,I284307);
DFFARX1 I_16566 (I284259,I2683,I284027,I284347,);
not I_16567 (I284355,I284347);
not I_16568 (I284372,I368134);
not I_16569 (I284389,I368137);
nor I_16570 (I284406,I284389,I368128);
nor I_16571 (I284019,I284355,I284406);
nor I_16572 (I284437,I284389,I368125);
and I_16573 (I284454,I284437,I368131);
or I_16574 (I284471,I284454,I368140);
DFFARX1 I_16575 (I284471,I2683,I284027,I284497,);
nor I_16576 (I284007,I284497,I284053);
not I_16577 (I284519,I284497);
and I_16578 (I284536,I284519,I284053);
nor I_16579 (I284001,I284078,I284536);
nand I_16580 (I284567,I284519,I284129);
nor I_16581 (I283995,I284389,I284567);
nand I_16582 (I283998,I284519,I284307);
nand I_16583 (I284612,I284129,I368137);
nor I_16584 (I284010,I284372,I284612);
not I_16585 (I284673,I2690);
DFFARX1 I_16586 (I178782,I2683,I284673,I284699,);
DFFARX1 I_16587 (I178794,I2683,I284673,I284716,);
not I_16588 (I284724,I284716);
not I_16589 (I284741,I178803);
nor I_16590 (I284758,I284741,I178779);
not I_16591 (I284775,I178797);
nor I_16592 (I284792,I284758,I178791);
nor I_16593 (I284809,I284716,I284792);
DFFARX1 I_16594 (I284809,I2683,I284673,I284659,);
nor I_16595 (I284840,I178791,I178779);
nand I_16596 (I284857,I284840,I178803);
DFFARX1 I_16597 (I284857,I2683,I284673,I284662,);
nor I_16598 (I284888,I284775,I178791);
nand I_16599 (I284905,I284888,I178785);
nor I_16600 (I284922,I284699,I284905);
DFFARX1 I_16601 (I284922,I2683,I284673,I284638,);
not I_16602 (I284953,I284905);
nand I_16603 (I284650,I284716,I284953);
DFFARX1 I_16604 (I284905,I2683,I284673,I284993,);
not I_16605 (I285001,I284993);
not I_16606 (I285018,I178791);
not I_16607 (I285035,I178800);
nor I_16608 (I285052,I285035,I178797);
nor I_16609 (I284665,I285001,I285052);
nor I_16610 (I285083,I285035,I178782);
and I_16611 (I285100,I285083,I178779);
or I_16612 (I285117,I285100,I178788);
DFFARX1 I_16613 (I285117,I2683,I284673,I285143,);
nor I_16614 (I284653,I285143,I284699);
not I_16615 (I285165,I285143);
and I_16616 (I285182,I285165,I284699);
nor I_16617 (I284647,I284724,I285182);
nand I_16618 (I285213,I285165,I284775);
nor I_16619 (I284641,I285035,I285213);
nand I_16620 (I284644,I285165,I284953);
nand I_16621 (I285258,I284775,I178800);
nor I_16622 (I284656,I285018,I285258);
not I_16623 (I285319,I2690);
DFFARX1 I_16624 (I255557,I2683,I285319,I285345,);
DFFARX1 I_16625 (I255554,I2683,I285319,I285362,);
not I_16626 (I285370,I285362);
not I_16627 (I285387,I255554);
nor I_16628 (I285404,I285387,I255557);
not I_16629 (I285421,I255569);
nor I_16630 (I285438,I285404,I255563);
nor I_16631 (I285455,I285362,I285438);
DFFARX1 I_16632 (I285455,I2683,I285319,I285305,);
nor I_16633 (I285486,I255563,I255557);
nand I_16634 (I285503,I285486,I255554);
DFFARX1 I_16635 (I285503,I2683,I285319,I285308,);
nor I_16636 (I285534,I285421,I255563);
nand I_16637 (I285551,I285534,I255551);
nor I_16638 (I285568,I285345,I285551);
DFFARX1 I_16639 (I285568,I2683,I285319,I285284,);
not I_16640 (I285599,I285551);
nand I_16641 (I285296,I285362,I285599);
DFFARX1 I_16642 (I285551,I2683,I285319,I285639,);
not I_16643 (I285647,I285639);
not I_16644 (I285664,I255563);
not I_16645 (I285681,I255560);
nor I_16646 (I285698,I285681,I255569);
nor I_16647 (I285311,I285647,I285698);
nor I_16648 (I285729,I285681,I255566);
and I_16649 (I285746,I285729,I255572);
or I_16650 (I285763,I285746,I255551);
DFFARX1 I_16651 (I285763,I2683,I285319,I285789,);
nor I_16652 (I285299,I285789,I285345);
not I_16653 (I285811,I285789);
and I_16654 (I285828,I285811,I285345);
nor I_16655 (I285293,I285370,I285828);
nand I_16656 (I285859,I285811,I285421);
nor I_16657 (I285287,I285681,I285859);
nand I_16658 (I285290,I285811,I285599);
nand I_16659 (I285904,I285421,I255560);
nor I_16660 (I285302,I285664,I285904);
not I_16661 (I285965,I2690);
DFFARX1 I_16662 (I317686,I2683,I285965,I285991,);
DFFARX1 I_16663 (I317689,I2683,I285965,I286008,);
not I_16664 (I286016,I286008);
not I_16665 (I286033,I317686);
nor I_16666 (I286050,I286033,I317698);
not I_16667 (I286067,I317707);
nor I_16668 (I286084,I286050,I317695);
nor I_16669 (I286101,I286008,I286084);
DFFARX1 I_16670 (I286101,I2683,I285965,I285951,);
nor I_16671 (I286132,I317695,I317698);
nand I_16672 (I286149,I286132,I317686);
DFFARX1 I_16673 (I286149,I2683,I285965,I285954,);
nor I_16674 (I286180,I286067,I317695);
nand I_16675 (I286197,I286180,I317701);
nor I_16676 (I286214,I285991,I286197);
DFFARX1 I_16677 (I286214,I2683,I285965,I285930,);
not I_16678 (I286245,I286197);
nand I_16679 (I285942,I286008,I286245);
DFFARX1 I_16680 (I286197,I2683,I285965,I286285,);
not I_16681 (I286293,I286285);
not I_16682 (I286310,I317695);
not I_16683 (I286327,I317692);
nor I_16684 (I286344,I286327,I317707);
nor I_16685 (I285957,I286293,I286344);
nor I_16686 (I286375,I286327,I317704);
and I_16687 (I286392,I286375,I317692);
or I_16688 (I286409,I286392,I317689);
DFFARX1 I_16689 (I286409,I2683,I285965,I286435,);
nor I_16690 (I285945,I286435,I285991);
not I_16691 (I286457,I286435);
and I_16692 (I286474,I286457,I285991);
nor I_16693 (I285939,I286016,I286474);
nand I_16694 (I286505,I286457,I286067);
nor I_16695 (I285933,I286327,I286505);
nand I_16696 (I285936,I286457,I286245);
nand I_16697 (I286550,I286067,I317692);
nor I_16698 (I285948,I286310,I286550);
not I_16699 (I286611,I2690);
DFFARX1 I_16700 (I226759,I2683,I286611,I286637,);
DFFARX1 I_16701 (I226753,I2683,I286611,I286654,);
not I_16702 (I286662,I286654);
not I_16703 (I286679,I226768);
nor I_16704 (I286696,I286679,I226753);
not I_16705 (I286713,I226762);
nor I_16706 (I286730,I286696,I226771);
nor I_16707 (I286747,I286654,I286730);
DFFARX1 I_16708 (I286747,I2683,I286611,I286597,);
nor I_16709 (I286778,I226771,I226753);
nand I_16710 (I286795,I286778,I226768);
DFFARX1 I_16711 (I286795,I2683,I286611,I286600,);
nor I_16712 (I286826,I286713,I226771);
nand I_16713 (I286843,I286826,I226756);
nor I_16714 (I286860,I286637,I286843);
DFFARX1 I_16715 (I286860,I2683,I286611,I286576,);
not I_16716 (I286891,I286843);
nand I_16717 (I286588,I286654,I286891);
DFFARX1 I_16718 (I286843,I2683,I286611,I286931,);
not I_16719 (I286939,I286931);
not I_16720 (I286956,I226771);
not I_16721 (I286973,I226765);
nor I_16722 (I286990,I286973,I226762);
nor I_16723 (I286603,I286939,I286990);
nor I_16724 (I287021,I286973,I226774);
and I_16725 (I287038,I287021,I226777);
or I_16726 (I287055,I287038,I226756);
DFFARX1 I_16727 (I287055,I2683,I286611,I287081,);
nor I_16728 (I286591,I287081,I286637);
not I_16729 (I287103,I287081);
and I_16730 (I287120,I287103,I286637);
nor I_16731 (I286585,I286662,I287120);
nand I_16732 (I287151,I287103,I286713);
nor I_16733 (I286579,I286973,I287151);
nand I_16734 (I286582,I287103,I286891);
nand I_16735 (I287196,I286713,I226765);
nor I_16736 (I286594,I286956,I287196);
not I_16737 (I287257,I2690);
DFFARX1 I_16738 (I109504,I2683,I287257,I287283,);
DFFARX1 I_16739 (I109510,I2683,I287257,I287300,);
not I_16740 (I287308,I287300);
not I_16741 (I287325,I109531);
nor I_16742 (I287342,I287325,I109519);
not I_16743 (I287359,I109528);
nor I_16744 (I287376,I287342,I109513);
nor I_16745 (I287393,I287300,I287376);
DFFARX1 I_16746 (I287393,I2683,I287257,I287243,);
nor I_16747 (I287424,I109513,I109519);
nand I_16748 (I287441,I287424,I109531);
DFFARX1 I_16749 (I287441,I2683,I287257,I287246,);
nor I_16750 (I287472,I287359,I109513);
nand I_16751 (I287489,I287472,I109504);
nor I_16752 (I287506,I287283,I287489);
DFFARX1 I_16753 (I287506,I2683,I287257,I287222,);
not I_16754 (I287537,I287489);
nand I_16755 (I287234,I287300,I287537);
DFFARX1 I_16756 (I287489,I2683,I287257,I287577,);
not I_16757 (I287585,I287577);
not I_16758 (I287602,I109513);
not I_16759 (I287619,I109516);
nor I_16760 (I287636,I287619,I109528);
nor I_16761 (I287249,I287585,I287636);
nor I_16762 (I287667,I287619,I109525);
and I_16763 (I287684,I287667,I109507);
or I_16764 (I287701,I287684,I109522);
DFFARX1 I_16765 (I287701,I2683,I287257,I287727,);
nor I_16766 (I287237,I287727,I287283);
not I_16767 (I287749,I287727);
and I_16768 (I287766,I287749,I287283);
nor I_16769 (I287231,I287308,I287766);
nand I_16770 (I287797,I287749,I287359);
nor I_16771 (I287225,I287619,I287797);
nand I_16772 (I287228,I287749,I287537);
nand I_16773 (I287842,I287359,I109516);
nor I_16774 (I287240,I287602,I287842);
not I_16775 (I287903,I2690);
DFFARX1 I_16776 (I346417,I2683,I287903,I287929,);
DFFARX1 I_16777 (I346399,I2683,I287903,I287946,);
not I_16778 (I287954,I287946);
not I_16779 (I287971,I346408);
nor I_16780 (I287988,I287971,I346420);
not I_16781 (I288005,I346402);
nor I_16782 (I288022,I287988,I346411);
nor I_16783 (I288039,I287946,I288022);
DFFARX1 I_16784 (I288039,I2683,I287903,I287889,);
nor I_16785 (I288070,I346411,I346420);
nand I_16786 (I288087,I288070,I346408);
DFFARX1 I_16787 (I288087,I2683,I287903,I287892,);
nor I_16788 (I288118,I288005,I346411);
nand I_16789 (I288135,I288118,I346423);
nor I_16790 (I288152,I287929,I288135);
DFFARX1 I_16791 (I288152,I2683,I287903,I287868,);
not I_16792 (I288183,I288135);
nand I_16793 (I287880,I287946,I288183);
DFFARX1 I_16794 (I288135,I2683,I287903,I288223,);
not I_16795 (I288231,I288223);
not I_16796 (I288248,I346411);
not I_16797 (I288265,I346399);
nor I_16798 (I288282,I288265,I346402);
nor I_16799 (I287895,I288231,I288282);
nor I_16800 (I288313,I288265,I346405);
and I_16801 (I288330,I288313,I346414);
or I_16802 (I288347,I288330,I346402);
DFFARX1 I_16803 (I288347,I2683,I287903,I288373,);
nor I_16804 (I287883,I288373,I287929);
not I_16805 (I288395,I288373);
and I_16806 (I288412,I288395,I287929);
nor I_16807 (I287877,I287954,I288412);
nand I_16808 (I288443,I288395,I288005);
nor I_16809 (I287871,I288265,I288443);
nand I_16810 (I287874,I288395,I288183);
nand I_16811 (I288488,I288005,I346399);
nor I_16812 (I287886,I288248,I288488);
not I_16813 (I288549,I2690);
DFFARX1 I_16814 (I211153,I2683,I288549,I288575,);
DFFARX1 I_16815 (I211147,I2683,I288549,I288592,);
not I_16816 (I288600,I288592);
not I_16817 (I288617,I211162);
nor I_16818 (I288634,I288617,I211147);
not I_16819 (I288651,I211156);
nor I_16820 (I288668,I288634,I211165);
nor I_16821 (I288685,I288592,I288668);
DFFARX1 I_16822 (I288685,I2683,I288549,I288535,);
nor I_16823 (I288716,I211165,I211147);
nand I_16824 (I288733,I288716,I211162);
DFFARX1 I_16825 (I288733,I2683,I288549,I288538,);
nor I_16826 (I288764,I288651,I211165);
nand I_16827 (I288781,I288764,I211150);
nor I_16828 (I288798,I288575,I288781);
DFFARX1 I_16829 (I288798,I2683,I288549,I288514,);
not I_16830 (I288829,I288781);
nand I_16831 (I288526,I288592,I288829);
DFFARX1 I_16832 (I288781,I2683,I288549,I288869,);
not I_16833 (I288877,I288869);
not I_16834 (I288894,I211165);
not I_16835 (I288911,I211159);
nor I_16836 (I288928,I288911,I211156);
nor I_16837 (I288541,I288877,I288928);
nor I_16838 (I288959,I288911,I211168);
and I_16839 (I288976,I288959,I211171);
or I_16840 (I288993,I288976,I211150);
DFFARX1 I_16841 (I288993,I2683,I288549,I289019,);
nor I_16842 (I288529,I289019,I288575);
not I_16843 (I289041,I289019);
and I_16844 (I289058,I289041,I288575);
nor I_16845 (I288523,I288600,I289058);
nand I_16846 (I289089,I289041,I288651);
nor I_16847 (I288517,I288911,I289089);
nand I_16848 (I288520,I289041,I288829);
nand I_16849 (I289134,I288651,I211159);
nor I_16850 (I288532,I288894,I289134);
not I_16851 (I289195,I2690);
DFFARX1 I_16852 (I100545,I2683,I289195,I289221,);
DFFARX1 I_16853 (I100551,I2683,I289195,I289238,);
not I_16854 (I289246,I289238);
not I_16855 (I289263,I100572);
nor I_16856 (I289280,I289263,I100560);
not I_16857 (I289297,I100569);
nor I_16858 (I289314,I289280,I100554);
nor I_16859 (I289331,I289238,I289314);
DFFARX1 I_16860 (I289331,I2683,I289195,I289181,);
nor I_16861 (I289362,I100554,I100560);
nand I_16862 (I289379,I289362,I100572);
DFFARX1 I_16863 (I289379,I2683,I289195,I289184,);
nor I_16864 (I289410,I289297,I100554);
nand I_16865 (I289427,I289410,I100545);
nor I_16866 (I289444,I289221,I289427);
DFFARX1 I_16867 (I289444,I2683,I289195,I289160,);
not I_16868 (I289475,I289427);
nand I_16869 (I289172,I289238,I289475);
DFFARX1 I_16870 (I289427,I2683,I289195,I289515,);
not I_16871 (I289523,I289515);
not I_16872 (I289540,I100554);
not I_16873 (I289557,I100557);
nor I_16874 (I289574,I289557,I100569);
nor I_16875 (I289187,I289523,I289574);
nor I_16876 (I289605,I289557,I100566);
and I_16877 (I289622,I289605,I100548);
or I_16878 (I289639,I289622,I100563);
DFFARX1 I_16879 (I289639,I2683,I289195,I289665,);
nor I_16880 (I289175,I289665,I289221);
not I_16881 (I289687,I289665);
and I_16882 (I289704,I289687,I289221);
nor I_16883 (I289169,I289246,I289704);
nand I_16884 (I289735,I289687,I289297);
nor I_16885 (I289163,I289557,I289735);
nand I_16886 (I289166,I289687,I289475);
nand I_16887 (I289780,I289297,I100557);
nor I_16888 (I289178,I289540,I289780);
not I_16889 (I289841,I2690);
DFFARX1 I_16890 (I23059,I2683,I289841,I289867,);
DFFARX1 I_16891 (I23065,I2683,I289841,I289884,);
not I_16892 (I289892,I289884);
not I_16893 (I289909,I23083);
nor I_16894 (I289926,I289909,I23062);
not I_16895 (I289943,I23068);
nor I_16896 (I289960,I289926,I23074);
nor I_16897 (I289977,I289884,I289960);
DFFARX1 I_16898 (I289977,I2683,I289841,I289827,);
nor I_16899 (I290008,I23074,I23062);
nand I_16900 (I290025,I290008,I23083);
DFFARX1 I_16901 (I290025,I2683,I289841,I289830,);
nor I_16902 (I290056,I289943,I23074);
nand I_16903 (I290073,I290056,I23080);
nor I_16904 (I290090,I289867,I290073);
DFFARX1 I_16905 (I290090,I2683,I289841,I289806,);
not I_16906 (I290121,I290073);
nand I_16907 (I289818,I289884,I290121);
DFFARX1 I_16908 (I290073,I2683,I289841,I290161,);
not I_16909 (I290169,I290161);
not I_16910 (I290186,I23074);
not I_16911 (I290203,I23062);
nor I_16912 (I290220,I290203,I23068);
nor I_16913 (I289833,I290169,I290220);
nor I_16914 (I290251,I290203,I23071);
and I_16915 (I290268,I290251,I23059);
or I_16916 (I290285,I290268,I23077);
DFFARX1 I_16917 (I290285,I2683,I289841,I290311,);
nor I_16918 (I289821,I290311,I289867);
not I_16919 (I290333,I290311);
and I_16920 (I290350,I290333,I289867);
nor I_16921 (I289815,I289892,I290350);
nand I_16922 (I290381,I290333,I289943);
nor I_16923 (I289809,I290203,I290381);
nand I_16924 (I289812,I290333,I290121);
nand I_16925 (I290426,I289943,I23062);
nor I_16926 (I289824,I290186,I290426);
not I_16927 (I290487,I2690);
DFFARX1 I_16928 (I395697,I2683,I290487,I290513,);
DFFARX1 I_16929 (I395694,I2683,I290487,I290530,);
not I_16930 (I290538,I290530);
not I_16931 (I290555,I395691);
nor I_16932 (I290572,I290555,I395682);
not I_16933 (I290589,I395703);
nor I_16934 (I290606,I290572,I395682);
nor I_16935 (I290623,I290530,I290606);
DFFARX1 I_16936 (I290623,I2683,I290487,I290473,);
nor I_16937 (I290654,I395682,I395682);
nand I_16938 (I290671,I290654,I395691);
DFFARX1 I_16939 (I290671,I2683,I290487,I290476,);
nor I_16940 (I290702,I290589,I395682);
nand I_16941 (I290719,I290702,I395706);
nor I_16942 (I290736,I290513,I290719);
DFFARX1 I_16943 (I290736,I2683,I290487,I290452,);
not I_16944 (I290767,I290719);
nand I_16945 (I290464,I290530,I290767);
DFFARX1 I_16946 (I290719,I2683,I290487,I290807,);
not I_16947 (I290815,I290807);
not I_16948 (I290832,I395682);
not I_16949 (I290849,I395685);
nor I_16950 (I290866,I290849,I395703);
nor I_16951 (I290479,I290815,I290866);
nor I_16952 (I290897,I290849,I395688);
and I_16953 (I290914,I290897,I395709);
or I_16954 (I290931,I290914,I395700);
DFFARX1 I_16955 (I290931,I2683,I290487,I290957,);
nor I_16956 (I290467,I290957,I290513);
not I_16957 (I290979,I290957);
and I_16958 (I290996,I290979,I290513);
nor I_16959 (I290461,I290538,I290996);
nand I_16960 (I291027,I290979,I290589);
nor I_16961 (I290455,I290849,I291027);
nand I_16962 (I290458,I290979,I290767);
nand I_16963 (I291072,I290589,I395685);
nor I_16964 (I290470,I290832,I291072);
not I_16965 (I291133,I2690);
DFFARX1 I_16966 (I138325,I2683,I291133,I291159,);
DFFARX1 I_16967 (I138322,I2683,I291133,I291176,);
not I_16968 (I291184,I291176);
not I_16969 (I291201,I138337);
nor I_16970 (I291218,I291201,I138340);
not I_16971 (I291235,I138328);
nor I_16972 (I291252,I291218,I138334);
nor I_16973 (I291269,I291176,I291252);
DFFARX1 I_16974 (I291269,I2683,I291133,I291119,);
nor I_16975 (I291300,I138334,I138340);
nand I_16976 (I291317,I291300,I138337);
DFFARX1 I_16977 (I291317,I2683,I291133,I291122,);
nor I_16978 (I291348,I291235,I138334);
nand I_16979 (I291365,I291348,I138346);
nor I_16980 (I291382,I291159,I291365);
DFFARX1 I_16981 (I291382,I2683,I291133,I291098,);
not I_16982 (I291413,I291365);
nand I_16983 (I291110,I291176,I291413);
DFFARX1 I_16984 (I291365,I2683,I291133,I291453,);
not I_16985 (I291461,I291453);
not I_16986 (I291478,I138334);
not I_16987 (I291495,I138319);
nor I_16988 (I291512,I291495,I138328);
nor I_16989 (I291125,I291461,I291512);
nor I_16990 (I291543,I291495,I138331);
and I_16991 (I291560,I291543,I138319);
or I_16992 (I291577,I291560,I138343);
DFFARX1 I_16993 (I291577,I2683,I291133,I291603,);
nor I_16994 (I291113,I291603,I291159);
not I_16995 (I291625,I291603);
and I_16996 (I291642,I291625,I291159);
nor I_16997 (I291107,I291184,I291642);
nand I_16998 (I291673,I291625,I291235);
nor I_16999 (I291101,I291495,I291673);
nand I_17000 (I291104,I291625,I291413);
nand I_17001 (I291718,I291235,I138319);
nor I_17002 (I291116,I291478,I291718);
not I_17003 (I291779,I2690);
DFFARX1 I_17004 (I139957,I2683,I291779,I291805,);
DFFARX1 I_17005 (I139954,I2683,I291779,I291822,);
not I_17006 (I291830,I291822);
not I_17007 (I291847,I139969);
nor I_17008 (I291864,I291847,I139972);
not I_17009 (I291881,I139960);
nor I_17010 (I291898,I291864,I139966);
nor I_17011 (I291915,I291822,I291898);
DFFARX1 I_17012 (I291915,I2683,I291779,I291765,);
nor I_17013 (I291946,I139966,I139972);
nand I_17014 (I291963,I291946,I139969);
DFFARX1 I_17015 (I291963,I2683,I291779,I291768,);
nor I_17016 (I291994,I291881,I139966);
nand I_17017 (I292011,I291994,I139978);
nor I_17018 (I292028,I291805,I292011);
DFFARX1 I_17019 (I292028,I2683,I291779,I291744,);
not I_17020 (I292059,I292011);
nand I_17021 (I291756,I291822,I292059);
DFFARX1 I_17022 (I292011,I2683,I291779,I292099,);
not I_17023 (I292107,I292099);
not I_17024 (I292124,I139966);
not I_17025 (I292141,I139951);
nor I_17026 (I292158,I292141,I139960);
nor I_17027 (I291771,I292107,I292158);
nor I_17028 (I292189,I292141,I139963);
and I_17029 (I292206,I292189,I139951);
or I_17030 (I292223,I292206,I139975);
DFFARX1 I_17031 (I292223,I2683,I291779,I292249,);
nor I_17032 (I291759,I292249,I291805);
not I_17033 (I292271,I292249);
and I_17034 (I292288,I292271,I291805);
nor I_17035 (I291753,I291830,I292288);
nand I_17036 (I292319,I292271,I291881);
nor I_17037 (I291747,I292141,I292319);
nand I_17038 (I291750,I292271,I292059);
nand I_17039 (I292364,I291881,I139951);
nor I_17040 (I291762,I292124,I292364);
not I_17041 (I292425,I2690);
DFFARX1 I_17042 (I54855,I2683,I292425,I292451,);
DFFARX1 I_17043 (I54867,I2683,I292425,I292468,);
not I_17044 (I292476,I292468);
not I_17045 (I292493,I54873);
nor I_17046 (I292510,I292493,I54858);
not I_17047 (I292527,I54849);
nor I_17048 (I292544,I292510,I54870);
nor I_17049 (I292561,I292468,I292544);
DFFARX1 I_17050 (I292561,I2683,I292425,I292411,);
nor I_17051 (I292592,I54870,I54858);
nand I_17052 (I292609,I292592,I54873);
DFFARX1 I_17053 (I292609,I2683,I292425,I292414,);
nor I_17054 (I292640,I292527,I54870);
nand I_17055 (I292657,I292640,I54852);
nor I_17056 (I292674,I292451,I292657);
DFFARX1 I_17057 (I292674,I2683,I292425,I292390,);
not I_17058 (I292705,I292657);
nand I_17059 (I292402,I292468,I292705);
DFFARX1 I_17060 (I292657,I2683,I292425,I292745,);
not I_17061 (I292753,I292745);
not I_17062 (I292770,I54870);
not I_17063 (I292787,I54861);
nor I_17064 (I292804,I292787,I54849);
nor I_17065 (I292417,I292753,I292804);
nor I_17066 (I292835,I292787,I54864);
and I_17067 (I292852,I292835,I54852);
or I_17068 (I292869,I292852,I54849);
DFFARX1 I_17069 (I292869,I2683,I292425,I292895,);
nor I_17070 (I292405,I292895,I292451);
not I_17071 (I292917,I292895);
and I_17072 (I292934,I292917,I292451);
nor I_17073 (I292399,I292476,I292934);
nand I_17074 (I292965,I292917,I292527);
nor I_17075 (I292393,I292787,I292965);
nand I_17076 (I292396,I292917,I292705);
nand I_17077 (I293010,I292527,I54861);
nor I_17078 (I292408,I292770,I293010);
not I_17079 (I293071,I2690);
DFFARX1 I_17080 (I150293,I2683,I293071,I293097,);
DFFARX1 I_17081 (I150290,I2683,I293071,I293114,);
not I_17082 (I293122,I293114);
not I_17083 (I293139,I150305);
nor I_17084 (I293156,I293139,I150308);
not I_17085 (I293173,I150296);
nor I_17086 (I293190,I293156,I150302);
nor I_17087 (I293207,I293114,I293190);
DFFARX1 I_17088 (I293207,I2683,I293071,I293057,);
nor I_17089 (I293238,I150302,I150308);
nand I_17090 (I293255,I293238,I150305);
DFFARX1 I_17091 (I293255,I2683,I293071,I293060,);
nor I_17092 (I293286,I293173,I150302);
nand I_17093 (I293303,I293286,I150314);
nor I_17094 (I293320,I293097,I293303);
DFFARX1 I_17095 (I293320,I2683,I293071,I293036,);
not I_17096 (I293351,I293303);
nand I_17097 (I293048,I293114,I293351);
DFFARX1 I_17098 (I293303,I2683,I293071,I293391,);
not I_17099 (I293399,I293391);
not I_17100 (I293416,I150302);
not I_17101 (I293433,I150287);
nor I_17102 (I293450,I293433,I150296);
nor I_17103 (I293063,I293399,I293450);
nor I_17104 (I293481,I293433,I150299);
and I_17105 (I293498,I293481,I150287);
or I_17106 (I293515,I293498,I150311);
DFFARX1 I_17107 (I293515,I2683,I293071,I293541,);
nor I_17108 (I293051,I293541,I293097);
not I_17109 (I293563,I293541);
and I_17110 (I293580,I293563,I293097);
nor I_17111 (I293045,I293122,I293580);
nand I_17112 (I293611,I293563,I293173);
nor I_17113 (I293039,I293433,I293611);
nand I_17114 (I293042,I293563,I293351);
nand I_17115 (I293656,I293173,I150287);
nor I_17116 (I293054,I293416,I293656);
not I_17117 (I293717,I2690);
DFFARX1 I_17118 (I17789,I2683,I293717,I293743,);
DFFARX1 I_17119 (I17795,I2683,I293717,I293760,);
not I_17120 (I293768,I293760);
not I_17121 (I293785,I17789);
nor I_17122 (I293802,I293785,I17801);
not I_17123 (I293819,I17813);
nor I_17124 (I293836,I293802,I17807);
nor I_17125 (I293853,I293760,I293836);
DFFARX1 I_17126 (I293853,I2683,I293717,I293703,);
nor I_17127 (I293884,I17807,I17801);
nand I_17128 (I293901,I293884,I17789);
DFFARX1 I_17129 (I293901,I2683,I293717,I293706,);
nor I_17130 (I293932,I293819,I17807);
nand I_17131 (I293949,I293932,I17792);
nor I_17132 (I293966,I293743,I293949);
DFFARX1 I_17133 (I293966,I2683,I293717,I293682,);
not I_17134 (I293997,I293949);
nand I_17135 (I293694,I293760,I293997);
DFFARX1 I_17136 (I293949,I2683,I293717,I294037,);
not I_17137 (I294045,I294037);
not I_17138 (I294062,I17807);
not I_17139 (I294079,I17792);
nor I_17140 (I294096,I294079,I17813);
nor I_17141 (I293709,I294045,I294096);
nor I_17142 (I294127,I294079,I17810);
and I_17143 (I294144,I294127,I17804);
or I_17144 (I294161,I294144,I17798);
DFFARX1 I_17145 (I294161,I2683,I293717,I294187,);
nor I_17146 (I293697,I294187,I293743);
not I_17147 (I294209,I294187);
and I_17148 (I294226,I294209,I293743);
nor I_17149 (I293691,I293768,I294226);
nand I_17150 (I294257,I294209,I293819);
nor I_17151 (I293685,I294079,I294257);
nand I_17152 (I293688,I294209,I293997);
nand I_17153 (I294302,I293819,I17792);
nor I_17154 (I293700,I294062,I294302);
not I_17155 (I294363,I2690);
DFFARX1 I_17156 (I341793,I2683,I294363,I294389,);
DFFARX1 I_17157 (I341775,I2683,I294363,I294406,);
not I_17158 (I294414,I294406);
not I_17159 (I294431,I341784);
nor I_17160 (I294448,I294431,I341796);
not I_17161 (I294465,I341778);
nor I_17162 (I294482,I294448,I341787);
nor I_17163 (I294499,I294406,I294482);
DFFARX1 I_17164 (I294499,I2683,I294363,I294349,);
nor I_17165 (I294530,I341787,I341796);
nand I_17166 (I294547,I294530,I341784);
DFFARX1 I_17167 (I294547,I2683,I294363,I294352,);
nor I_17168 (I294578,I294465,I341787);
nand I_17169 (I294595,I294578,I341799);
nor I_17170 (I294612,I294389,I294595);
DFFARX1 I_17171 (I294612,I2683,I294363,I294328,);
not I_17172 (I294643,I294595);
nand I_17173 (I294340,I294406,I294643);
DFFARX1 I_17174 (I294595,I2683,I294363,I294683,);
not I_17175 (I294691,I294683);
not I_17176 (I294708,I341787);
not I_17177 (I294725,I341775);
nor I_17178 (I294742,I294725,I341778);
nor I_17179 (I294355,I294691,I294742);
nor I_17180 (I294773,I294725,I341781);
and I_17181 (I294790,I294773,I341790);
or I_17182 (I294807,I294790,I341778);
DFFARX1 I_17183 (I294807,I2683,I294363,I294833,);
nor I_17184 (I294343,I294833,I294389);
not I_17185 (I294855,I294833);
and I_17186 (I294872,I294855,I294389);
nor I_17187 (I294337,I294414,I294872);
nand I_17188 (I294903,I294855,I294465);
nor I_17189 (I294331,I294725,I294903);
nand I_17190 (I294334,I294855,I294643);
nand I_17191 (I294948,I294465,I341775);
nor I_17192 (I294346,I294708,I294948);
not I_17193 (I295009,I2690);
DFFARX1 I_17194 (I319930,I2683,I295009,I295035,);
DFFARX1 I_17195 (I319933,I2683,I295009,I295052,);
not I_17196 (I295060,I295052);
not I_17197 (I295077,I319930);
nor I_17198 (I295094,I295077,I319942);
not I_17199 (I295111,I319951);
nor I_17200 (I295128,I295094,I319939);
nor I_17201 (I295145,I295052,I295128);
DFFARX1 I_17202 (I295145,I2683,I295009,I294995,);
nor I_17203 (I295176,I319939,I319942);
nand I_17204 (I295193,I295176,I319930);
DFFARX1 I_17205 (I295193,I2683,I295009,I294998,);
nor I_17206 (I295224,I295111,I319939);
nand I_17207 (I295241,I295224,I319945);
nor I_17208 (I295258,I295035,I295241);
DFFARX1 I_17209 (I295258,I2683,I295009,I294974,);
not I_17210 (I295289,I295241);
nand I_17211 (I294986,I295052,I295289);
DFFARX1 I_17212 (I295241,I2683,I295009,I295329,);
not I_17213 (I295337,I295329);
not I_17214 (I295354,I319939);
not I_17215 (I295371,I319936);
nor I_17216 (I295388,I295371,I319951);
nor I_17217 (I295001,I295337,I295388);
nor I_17218 (I295419,I295371,I319948);
and I_17219 (I295436,I295419,I319936);
or I_17220 (I295453,I295436,I319933);
DFFARX1 I_17221 (I295453,I2683,I295009,I295479,);
nor I_17222 (I294989,I295479,I295035);
not I_17223 (I295501,I295479);
and I_17224 (I295518,I295501,I295035);
nor I_17225 (I294983,I295060,I295518);
nand I_17226 (I295549,I295501,I295111);
nor I_17227 (I294977,I295371,I295549);
nand I_17228 (I294980,I295501,I295289);
nand I_17229 (I295594,I295111,I319936);
nor I_17230 (I294992,I295354,I295594);
not I_17231 (I295655,I2690);
DFFARX1 I_17232 (I25694,I2683,I295655,I295681,);
DFFARX1 I_17233 (I25700,I2683,I295655,I295698,);
not I_17234 (I295706,I295698);
not I_17235 (I295723,I25718);
nor I_17236 (I295740,I295723,I25697);
not I_17237 (I295757,I25703);
nor I_17238 (I295774,I295740,I25709);
nor I_17239 (I295791,I295698,I295774);
DFFARX1 I_17240 (I295791,I2683,I295655,I295641,);
nor I_17241 (I295822,I25709,I25697);
nand I_17242 (I295839,I295822,I25718);
DFFARX1 I_17243 (I295839,I2683,I295655,I295644,);
nor I_17244 (I295870,I295757,I25709);
nand I_17245 (I295887,I295870,I25715);
nor I_17246 (I295904,I295681,I295887);
DFFARX1 I_17247 (I295904,I2683,I295655,I295620,);
not I_17248 (I295935,I295887);
nand I_17249 (I295632,I295698,I295935);
DFFARX1 I_17250 (I295887,I2683,I295655,I295975,);
not I_17251 (I295983,I295975);
not I_17252 (I296000,I25709);
not I_17253 (I296017,I25697);
nor I_17254 (I296034,I296017,I25703);
nor I_17255 (I295647,I295983,I296034);
nor I_17256 (I296065,I296017,I25706);
and I_17257 (I296082,I296065,I25694);
or I_17258 (I296099,I296082,I25712);
DFFARX1 I_17259 (I296099,I2683,I295655,I296125,);
nor I_17260 (I295635,I296125,I295681);
not I_17261 (I296147,I296125);
and I_17262 (I296164,I296147,I295681);
nor I_17263 (I295629,I295706,I296164);
nand I_17264 (I296195,I296147,I295757);
nor I_17265 (I295623,I296017,I296195);
nand I_17266 (I295626,I296147,I295935);
nand I_17267 (I296240,I295757,I25697);
nor I_17268 (I295638,I296000,I296240);
not I_17269 (I296301,I2690);
DFFARX1 I_17270 (I209997,I2683,I296301,I296327,);
DFFARX1 I_17271 (I209991,I2683,I296301,I296344,);
not I_17272 (I296352,I296344);
not I_17273 (I296369,I210006);
nor I_17274 (I296386,I296369,I209991);
not I_17275 (I296403,I210000);
nor I_17276 (I296420,I296386,I210009);
nor I_17277 (I296437,I296344,I296420);
DFFARX1 I_17278 (I296437,I2683,I296301,I296287,);
nor I_17279 (I296468,I210009,I209991);
nand I_17280 (I296485,I296468,I210006);
DFFARX1 I_17281 (I296485,I2683,I296301,I296290,);
nor I_17282 (I296516,I296403,I210009);
nand I_17283 (I296533,I296516,I209994);
nor I_17284 (I296550,I296327,I296533);
DFFARX1 I_17285 (I296550,I2683,I296301,I296266,);
not I_17286 (I296581,I296533);
nand I_17287 (I296278,I296344,I296581);
DFFARX1 I_17288 (I296533,I2683,I296301,I296621,);
not I_17289 (I296629,I296621);
not I_17290 (I296646,I210009);
not I_17291 (I296663,I210003);
nor I_17292 (I296680,I296663,I210000);
nor I_17293 (I296293,I296629,I296680);
nor I_17294 (I296711,I296663,I210012);
and I_17295 (I296728,I296711,I210015);
or I_17296 (I296745,I296728,I209994);
DFFARX1 I_17297 (I296745,I2683,I296301,I296771,);
nor I_17298 (I296281,I296771,I296327);
not I_17299 (I296793,I296771);
and I_17300 (I296810,I296793,I296327);
nor I_17301 (I296275,I296352,I296810);
nand I_17302 (I296841,I296793,I296403);
nor I_17303 (I296269,I296663,I296841);
nand I_17304 (I296272,I296793,I296581);
nand I_17305 (I296886,I296403,I210003);
nor I_17306 (I296284,I296646,I296886);
not I_17307 (I296947,I2690);
DFFARX1 I_17308 (I36761,I2683,I296947,I296973,);
DFFARX1 I_17309 (I36767,I2683,I296947,I296990,);
not I_17310 (I296998,I296990);
not I_17311 (I297015,I36785);
nor I_17312 (I297032,I297015,I36764);
not I_17313 (I297049,I36770);
nor I_17314 (I297066,I297032,I36776);
nor I_17315 (I297083,I296990,I297066);
DFFARX1 I_17316 (I297083,I2683,I296947,I296933,);
nor I_17317 (I297114,I36776,I36764);
nand I_17318 (I297131,I297114,I36785);
DFFARX1 I_17319 (I297131,I2683,I296947,I296936,);
nor I_17320 (I297162,I297049,I36776);
nand I_17321 (I297179,I297162,I36782);
nor I_17322 (I297196,I296973,I297179);
DFFARX1 I_17323 (I297196,I2683,I296947,I296912,);
not I_17324 (I297227,I297179);
nand I_17325 (I296924,I296990,I297227);
DFFARX1 I_17326 (I297179,I2683,I296947,I297267,);
not I_17327 (I297275,I297267);
not I_17328 (I297292,I36776);
not I_17329 (I297309,I36764);
nor I_17330 (I297326,I297309,I36770);
nor I_17331 (I296939,I297275,I297326);
nor I_17332 (I297357,I297309,I36773);
and I_17333 (I297374,I297357,I36761);
or I_17334 (I297391,I297374,I36779);
DFFARX1 I_17335 (I297391,I2683,I296947,I297417,);
nor I_17336 (I296927,I297417,I296973);
not I_17337 (I297439,I297417);
and I_17338 (I297456,I297439,I296973);
nor I_17339 (I296921,I296998,I297456);
nand I_17340 (I297487,I297439,I297049);
nor I_17341 (I296915,I297309,I297487);
nand I_17342 (I296918,I297439,I297227);
nand I_17343 (I297532,I297049,I36764);
nor I_17344 (I296930,I297292,I297532);
not I_17345 (I297593,I2690);
DFFARX1 I_17346 (I334857,I2683,I297593,I297619,);
DFFARX1 I_17347 (I334839,I2683,I297593,I297636,);
not I_17348 (I297644,I297636);
not I_17349 (I297661,I334848);
nor I_17350 (I297678,I297661,I334860);
not I_17351 (I297695,I334842);
nor I_17352 (I297712,I297678,I334851);
nor I_17353 (I297729,I297636,I297712);
DFFARX1 I_17354 (I297729,I2683,I297593,I297579,);
nor I_17355 (I297760,I334851,I334860);
nand I_17356 (I297777,I297760,I334848);
DFFARX1 I_17357 (I297777,I2683,I297593,I297582,);
nor I_17358 (I297808,I297695,I334851);
nand I_17359 (I297825,I297808,I334863);
nor I_17360 (I297842,I297619,I297825);
DFFARX1 I_17361 (I297842,I2683,I297593,I297558,);
not I_17362 (I297873,I297825);
nand I_17363 (I297570,I297636,I297873);
DFFARX1 I_17364 (I297825,I2683,I297593,I297913,);
not I_17365 (I297921,I297913);
not I_17366 (I297938,I334851);
not I_17367 (I297955,I334839);
nor I_17368 (I297972,I297955,I334842);
nor I_17369 (I297585,I297921,I297972);
nor I_17370 (I298003,I297955,I334845);
and I_17371 (I298020,I298003,I334854);
or I_17372 (I298037,I298020,I334842);
DFFARX1 I_17373 (I298037,I2683,I297593,I298063,);
nor I_17374 (I297573,I298063,I297619);
not I_17375 (I298085,I298063);
and I_17376 (I298102,I298085,I297619);
nor I_17377 (I297567,I297644,I298102);
nand I_17378 (I298133,I298085,I297695);
nor I_17379 (I297561,I297955,I298133);
nand I_17380 (I297564,I298085,I297873);
nand I_17381 (I298178,I297695,I334839);
nor I_17382 (I297576,I297938,I298178);
not I_17383 (I298239,I2690);
DFFARX1 I_17384 (I320491,I2683,I298239,I298265,);
DFFARX1 I_17385 (I320494,I2683,I298239,I298282,);
not I_17386 (I298290,I298282);
not I_17387 (I298307,I320491);
nor I_17388 (I298324,I298307,I320503);
not I_17389 (I298341,I320512);
nor I_17390 (I298358,I298324,I320500);
nor I_17391 (I298375,I298282,I298358);
DFFARX1 I_17392 (I298375,I2683,I298239,I298225,);
nor I_17393 (I298406,I320500,I320503);
nand I_17394 (I298423,I298406,I320491);
DFFARX1 I_17395 (I298423,I2683,I298239,I298228,);
nor I_17396 (I298454,I298341,I320500);
nand I_17397 (I298471,I298454,I320506);
nor I_17398 (I298488,I298265,I298471);
DFFARX1 I_17399 (I298488,I2683,I298239,I298204,);
not I_17400 (I298519,I298471);
nand I_17401 (I298216,I298282,I298519);
DFFARX1 I_17402 (I298471,I2683,I298239,I298559,);
not I_17403 (I298567,I298559);
not I_17404 (I298584,I320500);
not I_17405 (I298601,I320497);
nor I_17406 (I298618,I298601,I320512);
nor I_17407 (I298231,I298567,I298618);
nor I_17408 (I298649,I298601,I320509);
and I_17409 (I298666,I298649,I320497);
or I_17410 (I298683,I298666,I320494);
DFFARX1 I_17411 (I298683,I2683,I298239,I298709,);
nor I_17412 (I298219,I298709,I298265);
not I_17413 (I298731,I298709);
and I_17414 (I298748,I298731,I298265);
nor I_17415 (I298213,I298290,I298748);
nand I_17416 (I298779,I298731,I298341);
nor I_17417 (I298207,I298601,I298779);
nand I_17418 (I298210,I298731,I298519);
nand I_17419 (I298824,I298341,I320497);
nor I_17420 (I298222,I298584,I298824);
not I_17421 (I298885,I2690);
DFFARX1 I_17422 (I400374,I2683,I298885,I298911,);
DFFARX1 I_17423 (I400398,I2683,I298885,I298928,);
not I_17424 (I298936,I298928);
not I_17425 (I298953,I400380);
nor I_17426 (I298970,I298953,I400389);
not I_17427 (I298987,I400374);
nor I_17428 (I299004,I298970,I400395);
nor I_17429 (I299021,I298928,I299004);
DFFARX1 I_17430 (I299021,I2683,I298885,I298871,);
nor I_17431 (I299052,I400395,I400389);
nand I_17432 (I299069,I299052,I400380);
DFFARX1 I_17433 (I299069,I2683,I298885,I298874,);
nor I_17434 (I299100,I298987,I400395);
nand I_17435 (I299117,I299100,I400392);
nor I_17436 (I299134,I298911,I299117);
DFFARX1 I_17437 (I299134,I2683,I298885,I298850,);
not I_17438 (I299165,I299117);
nand I_17439 (I298862,I298928,I299165);
DFFARX1 I_17440 (I299117,I2683,I298885,I299205,);
not I_17441 (I299213,I299205);
not I_17442 (I299230,I400395);
not I_17443 (I299247,I400386);
nor I_17444 (I299264,I299247,I400374);
nor I_17445 (I298877,I299213,I299264);
nor I_17446 (I299295,I299247,I400377);
and I_17447 (I299312,I299295,I400401);
or I_17448 (I299329,I299312,I400383);
DFFARX1 I_17449 (I299329,I2683,I298885,I299355,);
nor I_17450 (I298865,I299355,I298911);
not I_17451 (I299377,I299355);
and I_17452 (I299394,I299377,I298911);
nor I_17453 (I298859,I298936,I299394);
nand I_17454 (I299425,I299377,I298987);
nor I_17455 (I298853,I299247,I299425);
nand I_17456 (I298856,I299377,I299165);
nand I_17457 (I299470,I298987,I400386);
nor I_17458 (I298868,I299230,I299470);
not I_17459 (I299531,I2690);
DFFARX1 I_17460 (I47132,I2683,I299531,I299557,);
DFFARX1 I_17461 (I47135,I2683,I299531,I299574,);
not I_17462 (I299582,I299574);
not I_17463 (I299599,I47120);
nor I_17464 (I299616,I299599,I47114);
not I_17465 (I299633,I47123);
nor I_17466 (I299650,I299616,I47138);
nor I_17467 (I299667,I299574,I299650);
DFFARX1 I_17468 (I299667,I2683,I299531,I299517,);
nor I_17469 (I299698,I47138,I47114);
nand I_17470 (I299715,I299698,I47120);
DFFARX1 I_17471 (I299715,I2683,I299531,I299520,);
nor I_17472 (I299746,I299633,I47138);
nand I_17473 (I299763,I299746,I47141);
nor I_17474 (I299780,I299557,I299763);
DFFARX1 I_17475 (I299780,I2683,I299531,I299496,);
not I_17476 (I299811,I299763);
nand I_17477 (I299508,I299574,I299811);
DFFARX1 I_17478 (I299763,I2683,I299531,I299851,);
not I_17479 (I299859,I299851);
not I_17480 (I299876,I47138);
not I_17481 (I299893,I47117);
nor I_17482 (I299910,I299893,I47123);
nor I_17483 (I299523,I299859,I299910);
nor I_17484 (I299941,I299893,I47126);
and I_17485 (I299958,I299941,I47114);
or I_17486 (I299975,I299958,I47129);
DFFARX1 I_17487 (I299975,I2683,I299531,I300001,);
nor I_17488 (I299511,I300001,I299557);
not I_17489 (I300023,I300001);
and I_17490 (I300040,I300023,I299557);
nor I_17491 (I299505,I299582,I300040);
nand I_17492 (I300071,I300023,I299633);
nor I_17493 (I299499,I299893,I300071);
nand I_17494 (I299502,I300023,I299811);
nand I_17495 (I300116,I299633,I47117);
nor I_17496 (I299514,I299876,I300116);
not I_17497 (I300177,I2690);
DFFARX1 I_17498 (I3886,I2683,I300177,I300203,);
DFFARX1 I_17499 (I3883,I2683,I300177,I300220,);
not I_17500 (I300228,I300220);
not I_17501 (I300245,I3895);
nor I_17502 (I300262,I300245,I3892);
not I_17503 (I300279,I3901);
nor I_17504 (I300296,I300262,I3898);
nor I_17505 (I300313,I300220,I300296);
DFFARX1 I_17506 (I300313,I2683,I300177,I300163,);
nor I_17507 (I300344,I3898,I3892);
nand I_17508 (I300361,I300344,I3895);
DFFARX1 I_17509 (I300361,I2683,I300177,I300166,);
nor I_17510 (I300392,I300279,I3898);
nand I_17511 (I300409,I300392,I3889);
nor I_17512 (I300426,I300203,I300409);
DFFARX1 I_17513 (I300426,I2683,I300177,I300142,);
not I_17514 (I300457,I300409);
nand I_17515 (I300154,I300220,I300457);
DFFARX1 I_17516 (I300409,I2683,I300177,I300497,);
not I_17517 (I300505,I300497);
not I_17518 (I300522,I3898);
not I_17519 (I300539,I3889);
nor I_17520 (I300556,I300539,I3901);
nor I_17521 (I300169,I300505,I300556);
nor I_17522 (I300587,I300539,I3883);
and I_17523 (I300604,I300587,I3904);
or I_17524 (I300621,I300604,I3886);
DFFARX1 I_17525 (I300621,I2683,I300177,I300647,);
nor I_17526 (I300157,I300647,I300203);
not I_17527 (I300669,I300647);
and I_17528 (I300686,I300669,I300203);
nor I_17529 (I300151,I300228,I300686);
nand I_17530 (I300717,I300669,I300279);
nor I_17531 (I300145,I300539,I300717);
nand I_17532 (I300148,I300669,I300457);
nand I_17533 (I300762,I300279,I3889);
nor I_17534 (I300160,I300522,I300762);
not I_17535 (I300823,I2690);
DFFARX1 I_17536 (I19370,I2683,I300823,I300849,);
DFFARX1 I_17537 (I19376,I2683,I300823,I300866,);
not I_17538 (I300874,I300866);
not I_17539 (I300891,I19394);
nor I_17540 (I300908,I300891,I19373);
not I_17541 (I300925,I19379);
nor I_17542 (I300942,I300908,I19385);
nor I_17543 (I300959,I300866,I300942);
DFFARX1 I_17544 (I300959,I2683,I300823,I300809,);
nor I_17545 (I300990,I19385,I19373);
nand I_17546 (I301007,I300990,I19394);
DFFARX1 I_17547 (I301007,I2683,I300823,I300812,);
nor I_17548 (I301038,I300925,I19385);
nand I_17549 (I301055,I301038,I19391);
nor I_17550 (I301072,I300849,I301055);
DFFARX1 I_17551 (I301072,I2683,I300823,I300788,);
not I_17552 (I301103,I301055);
nand I_17553 (I300800,I300866,I301103);
DFFARX1 I_17554 (I301055,I2683,I300823,I301143,);
not I_17555 (I301151,I301143);
not I_17556 (I301168,I19385);
not I_17557 (I301185,I19373);
nor I_17558 (I301202,I301185,I19379);
nor I_17559 (I300815,I301151,I301202);
nor I_17560 (I301233,I301185,I19382);
and I_17561 (I301250,I301233,I19370);
or I_17562 (I301267,I301250,I19388);
DFFARX1 I_17563 (I301267,I2683,I300823,I301293,);
nor I_17564 (I300803,I301293,I300849);
not I_17565 (I301315,I301293);
and I_17566 (I301332,I301315,I300849);
nor I_17567 (I300797,I300874,I301332);
nand I_17568 (I301363,I301315,I300925);
nor I_17569 (I300791,I301185,I301363);
nand I_17570 (I300794,I301315,I301103);
nand I_17571 (I301408,I300925,I19373);
nor I_17572 (I300806,I301168,I301408);
not I_17573 (I301469,I2690);
DFFARX1 I_17574 (I391152,I2683,I301469,I301495,);
DFFARX1 I_17575 (I391146,I2683,I301469,I301512,);
not I_17576 (I301520,I301512);
not I_17577 (I301537,I391155);
nor I_17578 (I301554,I301537,I391167);
not I_17579 (I301571,I391149);
nor I_17580 (I301588,I301554,I391146);
nor I_17581 (I301605,I301512,I301588);
DFFARX1 I_17582 (I301605,I2683,I301469,I301455,);
nor I_17583 (I301636,I391146,I391167);
nand I_17584 (I301653,I301636,I391155);
DFFARX1 I_17585 (I301653,I2683,I301469,I301458,);
nor I_17586 (I301684,I301571,I391146);
nand I_17587 (I301701,I301684,I391143);
nor I_17588 (I301718,I301495,I301701);
DFFARX1 I_17589 (I301718,I2683,I301469,I301434,);
not I_17590 (I301749,I301701);
nand I_17591 (I301446,I301512,I301749);
DFFARX1 I_17592 (I301701,I2683,I301469,I301789,);
not I_17593 (I301797,I301789);
not I_17594 (I301814,I391146);
not I_17595 (I301831,I391164);
nor I_17596 (I301848,I301831,I391149);
nor I_17597 (I301461,I301797,I301848);
nor I_17598 (I301879,I301831,I391158);
and I_17599 (I301896,I301879,I391143);
or I_17600 (I301913,I301896,I391161);
DFFARX1 I_17601 (I301913,I2683,I301469,I301939,);
nor I_17602 (I301449,I301939,I301495);
not I_17603 (I301961,I301939);
and I_17604 (I301978,I301961,I301495);
nor I_17605 (I301443,I301520,I301978);
nand I_17606 (I302009,I301961,I301571);
nor I_17607 (I301437,I301831,I302009);
nand I_17608 (I301440,I301961,I301749);
nand I_17609 (I302054,I301571,I391164);
nor I_17610 (I301452,I301814,I302054);
not I_17611 (I302115,I2690);
DFFARX1 I_17612 (I310954,I2683,I302115,I302141,);
DFFARX1 I_17613 (I310957,I2683,I302115,I302158,);
not I_17614 (I302166,I302158);
not I_17615 (I302183,I310954);
nor I_17616 (I302200,I302183,I310966);
not I_17617 (I302217,I310975);
nor I_17618 (I302234,I302200,I310963);
nor I_17619 (I302251,I302158,I302234);
DFFARX1 I_17620 (I302251,I2683,I302115,I302101,);
nor I_17621 (I302282,I310963,I310966);
nand I_17622 (I302299,I302282,I310954);
DFFARX1 I_17623 (I302299,I2683,I302115,I302104,);
nor I_17624 (I302330,I302217,I310963);
nand I_17625 (I302347,I302330,I310969);
nor I_17626 (I302364,I302141,I302347);
DFFARX1 I_17627 (I302364,I2683,I302115,I302080,);
not I_17628 (I302395,I302347);
nand I_17629 (I302092,I302158,I302395);
DFFARX1 I_17630 (I302347,I2683,I302115,I302435,);
not I_17631 (I302443,I302435);
not I_17632 (I302460,I310963);
not I_17633 (I302477,I310960);
nor I_17634 (I302494,I302477,I310975);
nor I_17635 (I302107,I302443,I302494);
nor I_17636 (I302525,I302477,I310972);
and I_17637 (I302542,I302525,I310960);
or I_17638 (I302559,I302542,I310957);
DFFARX1 I_17639 (I302559,I2683,I302115,I302585,);
nor I_17640 (I302095,I302585,I302141);
not I_17641 (I302607,I302585);
and I_17642 (I302624,I302607,I302141);
nor I_17643 (I302089,I302166,I302624);
nand I_17644 (I302655,I302607,I302217);
nor I_17645 (I302083,I302477,I302655);
nand I_17646 (I302086,I302607,I302395);
nand I_17647 (I302700,I302217,I310960);
nor I_17648 (I302098,I302460,I302700);
not I_17649 (I302761,I2690);
DFFARX1 I_17650 (I178204,I2683,I302761,I302787,);
DFFARX1 I_17651 (I178216,I2683,I302761,I302804,);
not I_17652 (I302812,I302804);
not I_17653 (I302829,I178225);
nor I_17654 (I302846,I302829,I178201);
not I_17655 (I302863,I178219);
nor I_17656 (I302880,I302846,I178213);
nor I_17657 (I302897,I302804,I302880);
DFFARX1 I_17658 (I302897,I2683,I302761,I302747,);
nor I_17659 (I302928,I178213,I178201);
nand I_17660 (I302945,I302928,I178225);
DFFARX1 I_17661 (I302945,I2683,I302761,I302750,);
nor I_17662 (I302976,I302863,I178213);
nand I_17663 (I302993,I302976,I178207);
nor I_17664 (I303010,I302787,I302993);
DFFARX1 I_17665 (I303010,I2683,I302761,I302726,);
not I_17666 (I303041,I302993);
nand I_17667 (I302738,I302804,I303041);
DFFARX1 I_17668 (I302993,I2683,I302761,I303081,);
not I_17669 (I303089,I303081);
not I_17670 (I303106,I178213);
not I_17671 (I303123,I178222);
nor I_17672 (I303140,I303123,I178219);
nor I_17673 (I302753,I303089,I303140);
nor I_17674 (I303171,I303123,I178204);
and I_17675 (I303188,I303171,I178201);
or I_17676 (I303205,I303188,I178210);
DFFARX1 I_17677 (I303205,I2683,I302761,I303231,);
nor I_17678 (I302741,I303231,I302787);
not I_17679 (I303253,I303231);
and I_17680 (I303270,I303253,I302787);
nor I_17681 (I302735,I302812,I303270);
nand I_17682 (I303301,I303253,I302863);
nor I_17683 (I302729,I303123,I303301);
nand I_17684 (I302732,I303253,I303041);
nand I_17685 (I303346,I302863,I178222);
nor I_17686 (I302744,I303106,I303346);
not I_17687 (I303407,I2690);
DFFARX1 I_17688 (I369231,I2683,I303407,I303433,);
DFFARX1 I_17689 (I369237,I2683,I303407,I303450,);
not I_17690 (I303458,I303450);
not I_17691 (I303475,I369234);
nor I_17692 (I303492,I303475,I369213);
not I_17693 (I303509,I369216);
nor I_17694 (I303526,I303492,I369222);
nor I_17695 (I303543,I303450,I303526);
DFFARX1 I_17696 (I303543,I2683,I303407,I303393,);
nor I_17697 (I303574,I369222,I369213);
nand I_17698 (I303591,I303574,I369234);
DFFARX1 I_17699 (I303591,I2683,I303407,I303396,);
nor I_17700 (I303622,I303509,I369222);
nand I_17701 (I303639,I303622,I369216);
nor I_17702 (I303656,I303433,I303639);
DFFARX1 I_17703 (I303656,I2683,I303407,I303372,);
not I_17704 (I303687,I303639);
nand I_17705 (I303384,I303450,I303687);
DFFARX1 I_17706 (I303639,I2683,I303407,I303727,);
not I_17707 (I303735,I303727);
not I_17708 (I303752,I369222);
not I_17709 (I303769,I369225);
nor I_17710 (I303786,I303769,I369216);
nor I_17711 (I303399,I303735,I303786);
nor I_17712 (I303817,I303769,I369213);
and I_17713 (I303834,I303817,I369219);
or I_17714 (I303851,I303834,I369228);
DFFARX1 I_17715 (I303851,I2683,I303407,I303877,);
nor I_17716 (I303387,I303877,I303433);
not I_17717 (I303899,I303877);
and I_17718 (I303916,I303899,I303433);
nor I_17719 (I303381,I303458,I303916);
nand I_17720 (I303947,I303899,I303509);
nor I_17721 (I303375,I303769,I303947);
nand I_17722 (I303378,I303899,I303687);
nand I_17723 (I303992,I303509,I369225);
nor I_17724 (I303390,I303752,I303992);
not I_17725 (I304053,I2690);
DFFARX1 I_17726 (I99491,I2683,I304053,I304079,);
DFFARX1 I_17727 (I99497,I2683,I304053,I304096,);
not I_17728 (I304104,I304096);
not I_17729 (I304121,I99518);
nor I_17730 (I304138,I304121,I99506);
not I_17731 (I304155,I99515);
nor I_17732 (I304172,I304138,I99500);
nor I_17733 (I304189,I304096,I304172);
DFFARX1 I_17734 (I304189,I2683,I304053,I304039,);
nor I_17735 (I304220,I99500,I99506);
nand I_17736 (I304237,I304220,I99518);
DFFARX1 I_17737 (I304237,I2683,I304053,I304042,);
nor I_17738 (I304268,I304155,I99500);
nand I_17739 (I304285,I304268,I99491);
nor I_17740 (I304302,I304079,I304285);
DFFARX1 I_17741 (I304302,I2683,I304053,I304018,);
not I_17742 (I304333,I304285);
nand I_17743 (I304030,I304096,I304333);
DFFARX1 I_17744 (I304285,I2683,I304053,I304373,);
not I_17745 (I304381,I304373);
not I_17746 (I304398,I99500);
not I_17747 (I304415,I99503);
nor I_17748 (I304432,I304415,I99515);
nor I_17749 (I304045,I304381,I304432);
nor I_17750 (I304463,I304415,I99512);
and I_17751 (I304480,I304463,I99494);
or I_17752 (I304497,I304480,I99509);
DFFARX1 I_17753 (I304497,I2683,I304053,I304523,);
nor I_17754 (I304033,I304523,I304079);
not I_17755 (I304545,I304523);
and I_17756 (I304562,I304545,I304079);
nor I_17757 (I304027,I304104,I304562);
nand I_17758 (I304593,I304545,I304155);
nor I_17759 (I304021,I304415,I304593);
nand I_17760 (I304024,I304545,I304333);
nand I_17761 (I304638,I304155,I99503);
nor I_17762 (I304036,I304398,I304638);
not I_17763 (I304699,I2690);
DFFARX1 I_17764 (I143221,I2683,I304699,I304725,);
DFFARX1 I_17765 (I143218,I2683,I304699,I304742,);
not I_17766 (I304750,I304742);
not I_17767 (I304767,I143233);
nor I_17768 (I304784,I304767,I143236);
not I_17769 (I304801,I143224);
nor I_17770 (I304818,I304784,I143230);
nor I_17771 (I304835,I304742,I304818);
DFFARX1 I_17772 (I304835,I2683,I304699,I304685,);
nor I_17773 (I304866,I143230,I143236);
nand I_17774 (I304883,I304866,I143233);
DFFARX1 I_17775 (I304883,I2683,I304699,I304688,);
nor I_17776 (I304914,I304801,I143230);
nand I_17777 (I304931,I304914,I143242);
nor I_17778 (I304948,I304725,I304931);
DFFARX1 I_17779 (I304948,I2683,I304699,I304664,);
not I_17780 (I304979,I304931);
nand I_17781 (I304676,I304742,I304979);
DFFARX1 I_17782 (I304931,I2683,I304699,I305019,);
not I_17783 (I305027,I305019);
not I_17784 (I305044,I143230);
not I_17785 (I305061,I143215);
nor I_17786 (I305078,I305061,I143224);
nor I_17787 (I304691,I305027,I305078);
nor I_17788 (I305109,I305061,I143227);
and I_17789 (I305126,I305109,I143215);
or I_17790 (I305143,I305126,I143239);
DFFARX1 I_17791 (I305143,I2683,I304699,I305169,);
nor I_17792 (I304679,I305169,I304725);
not I_17793 (I305191,I305169);
and I_17794 (I305208,I305191,I304725);
nor I_17795 (I304673,I304750,I305208);
nand I_17796 (I305239,I305191,I304801);
nor I_17797 (I304667,I305061,I305239);
nand I_17798 (I304670,I305191,I304979);
nand I_17799 (I305284,I304801,I143215);
nor I_17800 (I304682,I305044,I305284);
not I_17801 (I305345,I2690);
DFFARX1 I_17802 (I365423,I2683,I305345,I305371,);
DFFARX1 I_17803 (I365429,I2683,I305345,I305388,);
not I_17804 (I305396,I305388);
not I_17805 (I305413,I365426);
nor I_17806 (I305430,I305413,I365405);
not I_17807 (I305447,I365408);
nor I_17808 (I305464,I305430,I365414);
nor I_17809 (I305481,I305388,I305464);
DFFARX1 I_17810 (I305481,I2683,I305345,I305331,);
nor I_17811 (I305512,I365414,I365405);
nand I_17812 (I305529,I305512,I365426);
DFFARX1 I_17813 (I305529,I2683,I305345,I305334,);
nor I_17814 (I305560,I305447,I365414);
nand I_17815 (I305577,I305560,I365408);
nor I_17816 (I305594,I305371,I305577);
DFFARX1 I_17817 (I305594,I2683,I305345,I305310,);
not I_17818 (I305625,I305577);
nand I_17819 (I305322,I305388,I305625);
DFFARX1 I_17820 (I305577,I2683,I305345,I305665,);
not I_17821 (I305673,I305665);
not I_17822 (I305690,I365414);
not I_17823 (I305707,I365417);
nor I_17824 (I305724,I305707,I365408);
nor I_17825 (I305337,I305673,I305724);
nor I_17826 (I305755,I305707,I365405);
and I_17827 (I305772,I305755,I365411);
or I_17828 (I305789,I305772,I365420);
DFFARX1 I_17829 (I305789,I2683,I305345,I305815,);
nor I_17830 (I305325,I305815,I305371);
not I_17831 (I305837,I305815);
and I_17832 (I305854,I305837,I305371);
nor I_17833 (I305319,I305396,I305854);
nand I_17834 (I305885,I305837,I305447);
nor I_17835 (I305313,I305707,I305885);
nand I_17836 (I305316,I305837,I305625);
nand I_17837 (I305930,I305447,I365417);
nor I_17838 (I305328,I305690,I305930);
not I_17839 (I305991,I2690);
DFFARX1 I_17840 (I86316,I2683,I305991,I306017,);
DFFARX1 I_17841 (I86322,I2683,I305991,I306034,);
not I_17842 (I306042,I306034);
not I_17843 (I306059,I86343);
nor I_17844 (I306076,I306059,I86331);
not I_17845 (I306093,I86340);
nor I_17846 (I306110,I306076,I86325);
nor I_17847 (I306127,I306034,I306110);
DFFARX1 I_17848 (I306127,I2683,I305991,I305977,);
nor I_17849 (I306158,I86325,I86331);
nand I_17850 (I306175,I306158,I86343);
DFFARX1 I_17851 (I306175,I2683,I305991,I305980,);
nor I_17852 (I306206,I306093,I86325);
nand I_17853 (I306223,I306206,I86316);
nor I_17854 (I306240,I306017,I306223);
DFFARX1 I_17855 (I306240,I2683,I305991,I305956,);
not I_17856 (I306271,I306223);
nand I_17857 (I305968,I306034,I306271);
DFFARX1 I_17858 (I306223,I2683,I305991,I306311,);
not I_17859 (I306319,I306311);
not I_17860 (I306336,I86325);
not I_17861 (I306353,I86328);
nor I_17862 (I306370,I306353,I86340);
nor I_17863 (I305983,I306319,I306370);
nor I_17864 (I306401,I306353,I86337);
and I_17865 (I306418,I306401,I86319);
or I_17866 (I306435,I306418,I86334);
DFFARX1 I_17867 (I306435,I2683,I305991,I306461,);
nor I_17868 (I305971,I306461,I306017);
not I_17869 (I306483,I306461);
and I_17870 (I306500,I306483,I306017);
nor I_17871 (I305965,I306042,I306500);
nand I_17872 (I306531,I306483,I306093);
nor I_17873 (I305959,I306353,I306531);
nand I_17874 (I305962,I306483,I306271);
nand I_17875 (I306576,I306093,I86328);
nor I_17876 (I305974,I306336,I306576);
not I_17877 (I306637,I2690);
DFFARX1 I_17878 (I350463,I2683,I306637,I306663,);
DFFARX1 I_17879 (I350445,I2683,I306637,I306680,);
not I_17880 (I306688,I306680);
not I_17881 (I306705,I350454);
nor I_17882 (I306722,I306705,I350466);
not I_17883 (I306739,I350448);
nor I_17884 (I306756,I306722,I350457);
nor I_17885 (I306773,I306680,I306756);
DFFARX1 I_17886 (I306773,I2683,I306637,I306623,);
nor I_17887 (I306804,I350457,I350466);
nand I_17888 (I306821,I306804,I350454);
DFFARX1 I_17889 (I306821,I2683,I306637,I306626,);
nor I_17890 (I306852,I306739,I350457);
nand I_17891 (I306869,I306852,I350469);
nor I_17892 (I306886,I306663,I306869);
DFFARX1 I_17893 (I306886,I2683,I306637,I306602,);
not I_17894 (I306917,I306869);
nand I_17895 (I306614,I306680,I306917);
DFFARX1 I_17896 (I306869,I2683,I306637,I306957,);
not I_17897 (I306965,I306957);
not I_17898 (I306982,I350457);
not I_17899 (I306999,I350445);
nor I_17900 (I307016,I306999,I350448);
nor I_17901 (I306629,I306965,I307016);
nor I_17902 (I307047,I306999,I350451);
and I_17903 (I307064,I307047,I350460);
or I_17904 (I307081,I307064,I350448);
DFFARX1 I_17905 (I307081,I2683,I306637,I307107,);
nor I_17906 (I306617,I307107,I306663);
not I_17907 (I307129,I307107);
and I_17908 (I307146,I307129,I306663);
nor I_17909 (I306611,I306688,I307146);
nand I_17910 (I307177,I307129,I306739);
nor I_17911 (I306605,I306999,I307177);
nand I_17912 (I306608,I307129,I306917);
nand I_17913 (I307222,I306739,I350445);
nor I_17914 (I306620,I306982,I307222);
not I_17915 (I307283,I2690);
DFFARX1 I_17916 (I377391,I2683,I307283,I307309,);
DFFARX1 I_17917 (I377397,I2683,I307283,I307326,);
not I_17918 (I307334,I307326);
not I_17919 (I307351,I377394);
nor I_17920 (I307368,I307351,I377373);
not I_17921 (I307385,I377376);
nor I_17922 (I307402,I307368,I377382);
nor I_17923 (I307419,I307326,I307402);
DFFARX1 I_17924 (I307419,I2683,I307283,I307269,);
nor I_17925 (I307450,I377382,I377373);
nand I_17926 (I307467,I307450,I377394);
DFFARX1 I_17927 (I307467,I2683,I307283,I307272,);
nor I_17928 (I307498,I307385,I377382);
nand I_17929 (I307515,I307498,I377376);
nor I_17930 (I307532,I307309,I307515);
DFFARX1 I_17931 (I307532,I2683,I307283,I307248,);
not I_17932 (I307563,I307515);
nand I_17933 (I307260,I307326,I307563);
DFFARX1 I_17934 (I307515,I2683,I307283,I307603,);
not I_17935 (I307611,I307603);
not I_17936 (I307628,I377382);
not I_17937 (I307645,I377385);
nor I_17938 (I307662,I307645,I377376);
nor I_17939 (I307275,I307611,I307662);
nor I_17940 (I307693,I307645,I377373);
and I_17941 (I307710,I307693,I377379);
or I_17942 (I307727,I307710,I377388);
DFFARX1 I_17943 (I307727,I2683,I307283,I307753,);
nor I_17944 (I307263,I307753,I307309);
not I_17945 (I307775,I307753);
and I_17946 (I307792,I307775,I307309);
nor I_17947 (I307257,I307334,I307792);
nand I_17948 (I307823,I307775,I307385);
nor I_17949 (I307251,I307645,I307823);
nand I_17950 (I307254,I307775,I307563);
nand I_17951 (I307868,I307385,I377385);
nor I_17952 (I307266,I307628,I307868);
not I_17953 (I307929,I2690);
DFFARX1 I_17954 (I1508,I2683,I307929,I307955,);
DFFARX1 I_17955 (I2484,I2683,I307929,I307972,);
not I_17956 (I307980,I307972);
not I_17957 (I307997,I1876);
nor I_17958 (I308014,I307997,I2020);
not I_17959 (I308031,I2452);
nor I_17960 (I308048,I308014,I1764);
nor I_17961 (I308065,I307972,I308048);
DFFARX1 I_17962 (I308065,I2683,I307929,I307915,);
nor I_17963 (I308096,I1764,I2020);
nand I_17964 (I308113,I308096,I1876);
DFFARX1 I_17965 (I308113,I2683,I307929,I307918,);
nor I_17966 (I308144,I308031,I1764);
nand I_17967 (I308161,I308144,I2252);
nor I_17968 (I308178,I307955,I308161);
DFFARX1 I_17969 (I308178,I2683,I307929,I307894,);
not I_17970 (I308209,I308161);
nand I_17971 (I307906,I307972,I308209);
DFFARX1 I_17972 (I308161,I2683,I307929,I308249,);
not I_17973 (I308257,I308249);
not I_17974 (I308274,I1764);
not I_17975 (I308291,I2036);
nor I_17976 (I308308,I308291,I2452);
nor I_17977 (I307921,I308257,I308308);
nor I_17978 (I308339,I308291,I2596);
and I_17979 (I308356,I308339,I2476);
or I_17980 (I308373,I308356,I1988);
DFFARX1 I_17981 (I308373,I2683,I307929,I308399,);
nor I_17982 (I307909,I308399,I307955);
not I_17983 (I308421,I308399);
and I_17984 (I308438,I308421,I307955);
nor I_17985 (I307903,I307980,I308438);
nand I_17986 (I308469,I308421,I308031);
nor I_17987 (I307897,I308291,I308469);
nand I_17988 (I307900,I308421,I308209);
nand I_17989 (I308514,I308031,I2036);
nor I_17990 (I307912,I308274,I308514);
not I_17991 (I308575,I2690);
DFFARX1 I_17992 (I13573,I2683,I308575,I308601,);
DFFARX1 I_17993 (I13579,I2683,I308575,I308618,);
not I_17994 (I308626,I308618);
not I_17995 (I308643,I13573);
nor I_17996 (I308660,I308643,I13585);
not I_17997 (I308677,I13597);
nor I_17998 (I308694,I308660,I13591);
nor I_17999 (I308711,I308618,I308694);
DFFARX1 I_18000 (I308711,I2683,I308575,I308561,);
nor I_18001 (I308742,I13591,I13585);
nand I_18002 (I308759,I308742,I13573);
DFFARX1 I_18003 (I308759,I2683,I308575,I308564,);
nor I_18004 (I308790,I308677,I13591);
nand I_18005 (I308807,I308790,I13576);
nor I_18006 (I308824,I308601,I308807);
DFFARX1 I_18007 (I308824,I2683,I308575,I308540,);
not I_18008 (I308855,I308807);
nand I_18009 (I308552,I308618,I308855);
DFFARX1 I_18010 (I308807,I2683,I308575,I308895,);
not I_18011 (I308903,I308895);
not I_18012 (I308920,I13591);
not I_18013 (I308937,I13576);
nor I_18014 (I308954,I308937,I13597);
nor I_18015 (I308567,I308903,I308954);
nor I_18016 (I308985,I308937,I13594);
and I_18017 (I309002,I308985,I13588);
or I_18018 (I309019,I309002,I13582);
DFFARX1 I_18019 (I309019,I2683,I308575,I309045,);
nor I_18020 (I308555,I309045,I308601);
not I_18021 (I309067,I309045);
and I_18022 (I309084,I309067,I308601);
nor I_18023 (I308549,I308626,I309084);
nand I_18024 (I309115,I309067,I308677);
nor I_18025 (I308543,I308937,I309115);
nand I_18026 (I308546,I309067,I308855);
nand I_18027 (I309160,I308677,I13576);
nor I_18028 (I308558,I308920,I309160);
not I_18029 (I309221,I2690);
DFFARX1 I_18030 (I133429,I2683,I309221,I309247,);
DFFARX1 I_18031 (I133426,I2683,I309221,I309264,);
not I_18032 (I309272,I309264);
not I_18033 (I309289,I133441);
nor I_18034 (I309306,I309289,I133444);
not I_18035 (I309323,I133432);
nor I_18036 (I309340,I309306,I133438);
nor I_18037 (I309357,I309264,I309340);
DFFARX1 I_18038 (I309357,I2683,I309221,I309207,);
nor I_18039 (I309388,I133438,I133444);
nand I_18040 (I309405,I309388,I133441);
DFFARX1 I_18041 (I309405,I2683,I309221,I309210,);
nor I_18042 (I309436,I309323,I133438);
nand I_18043 (I309453,I309436,I133450);
nor I_18044 (I309470,I309247,I309453);
DFFARX1 I_18045 (I309470,I2683,I309221,I309186,);
not I_18046 (I309501,I309453);
nand I_18047 (I309198,I309264,I309501);
DFFARX1 I_18048 (I309453,I2683,I309221,I309541,);
not I_18049 (I309549,I309541);
not I_18050 (I309566,I133438);
not I_18051 (I309583,I133423);
nor I_18052 (I309600,I309583,I133432);
nor I_18053 (I309213,I309549,I309600);
nor I_18054 (I309631,I309583,I133435);
and I_18055 (I309648,I309631,I133423);
or I_18056 (I309665,I309648,I133447);
DFFARX1 I_18057 (I309665,I2683,I309221,I309691,);
nor I_18058 (I309201,I309691,I309247);
not I_18059 (I309713,I309691);
and I_18060 (I309730,I309713,I309247);
nor I_18061 (I309195,I309272,I309730);
nand I_18062 (I309761,I309713,I309323);
nor I_18063 (I309189,I309583,I309761);
nand I_18064 (I309192,I309713,I309501);
nand I_18065 (I309806,I309323,I133423);
nor I_18066 (I309204,I309566,I309806);
not I_18067 (I309861,I2690);
DFFARX1 I_18068 (I51877,I2683,I309861,I309887,);
DFFARX1 I_18069 (I309887,I2683,I309861,I309904,);
not I_18070 (I309853,I309904);
not I_18071 (I309926,I309887);
DFFARX1 I_18072 (I51892,I2683,I309861,I309952,);
nand I_18073 (I309960,I309952,I51874);
not I_18074 (I309977,I51874);
not I_18075 (I309994,I51883);
nand I_18076 (I310011,I51889,I51880);
and I_18077 (I310028,I51889,I51880);
not I_18078 (I310045,I51877);
nand I_18079 (I310062,I310045,I309994);
nor I_18080 (I309835,I310062,I309960);
nor I_18081 (I310093,I309977,I310062);
nand I_18082 (I309838,I310028,I310093);
not I_18083 (I310124,I51874);
nor I_18084 (I310141,I310124,I51889);
nor I_18085 (I310158,I310141,I51877);
nor I_18086 (I310175,I309926,I310158);
DFFARX1 I_18087 (I310175,I2683,I309861,I309847,);
not I_18088 (I310206,I310141);
DFFARX1 I_18089 (I310206,I2683,I309861,I309850,);
and I_18090 (I309844,I309952,I310141);
nor I_18091 (I310251,I310124,I51898);
and I_18092 (I310268,I310251,I51895);
or I_18093 (I310285,I310268,I51886);
DFFARX1 I_18094 (I310285,I2683,I309861,I310311,);
nor I_18095 (I310319,I310311,I310045);
DFFARX1 I_18096 (I310319,I2683,I309861,I309832,);
nand I_18097 (I310350,I310311,I309952);
nand I_18098 (I310367,I310045,I310350);
nor I_18099 (I309841,I310367,I310011);
not I_18100 (I310422,I2690);
DFFARX1 I_18101 (I417644,I2683,I310422,I310448,);
DFFARX1 I_18102 (I310448,I2683,I310422,I310465,);
not I_18103 (I310414,I310465);
not I_18104 (I310487,I310448);
DFFARX1 I_18105 (I417638,I2683,I310422,I310513,);
nand I_18106 (I310521,I310513,I417629);
not I_18107 (I310538,I417629);
not I_18108 (I310555,I417656);
nand I_18109 (I310572,I417641,I417650);
and I_18110 (I310589,I417641,I417650);
not I_18111 (I310606,I417635);
nand I_18112 (I310623,I310606,I310555);
nor I_18113 (I310396,I310623,I310521);
nor I_18114 (I310654,I310538,I310623);
nand I_18115 (I310399,I310589,I310654);
not I_18116 (I310685,I417653);
nor I_18117 (I310702,I310685,I417641);
nor I_18118 (I310719,I310702,I417635);
nor I_18119 (I310736,I310487,I310719);
DFFARX1 I_18120 (I310736,I2683,I310422,I310408,);
not I_18121 (I310767,I310702);
DFFARX1 I_18122 (I310767,I2683,I310422,I310411,);
and I_18123 (I310405,I310513,I310702);
nor I_18124 (I310812,I310685,I417647);
and I_18125 (I310829,I310812,I417629);
or I_18126 (I310846,I310829,I417632);
DFFARX1 I_18127 (I310846,I2683,I310422,I310872,);
nor I_18128 (I310880,I310872,I310606);
DFFARX1 I_18129 (I310880,I2683,I310422,I310393,);
nand I_18130 (I310911,I310872,I310513);
nand I_18131 (I310928,I310606,I310911);
nor I_18132 (I310402,I310928,I310572);
not I_18133 (I310983,I2690);
DFFARX1 I_18134 (I221554,I2683,I310983,I311009,);
DFFARX1 I_18135 (I311009,I2683,I310983,I311026,);
not I_18136 (I310975,I311026);
not I_18137 (I311048,I311009);
DFFARX1 I_18138 (I221566,I2683,I310983,I311074,);
nand I_18139 (I311082,I311074,I221575);
not I_18140 (I311099,I221575);
not I_18141 (I311116,I221557);
nand I_18142 (I311133,I221560,I221551);
and I_18143 (I311150,I221560,I221551);
not I_18144 (I311167,I221569);
nand I_18145 (I311184,I311167,I311116);
nor I_18146 (I310957,I311184,I311082);
nor I_18147 (I311215,I311099,I311184);
nand I_18148 (I310960,I311150,I311215);
not I_18149 (I311246,I221572);
nor I_18150 (I311263,I311246,I221560);
nor I_18151 (I311280,I311263,I221569);
nor I_18152 (I311297,I311048,I311280);
DFFARX1 I_18153 (I311297,I2683,I310983,I310969,);
not I_18154 (I311328,I311263);
DFFARX1 I_18155 (I311328,I2683,I310983,I310972,);
and I_18156 (I310966,I311074,I311263);
nor I_18157 (I311373,I311246,I221551);
and I_18158 (I311390,I311373,I221563);
or I_18159 (I311407,I311390,I221554);
DFFARX1 I_18160 (I311407,I2683,I310983,I311433,);
nor I_18161 (I311441,I311433,I311167);
DFFARX1 I_18162 (I311441,I2683,I310983,I310954,);
nand I_18163 (I311472,I311433,I311074);
nand I_18164 (I311489,I311167,I311472);
nor I_18165 (I310963,I311489,I311133);
not I_18166 (I311544,I2690);
DFFARX1 I_18167 (I105309,I2683,I311544,I311570,);
DFFARX1 I_18168 (I311570,I2683,I311544,I311587,);
not I_18169 (I311536,I311587);
not I_18170 (I311609,I311570);
DFFARX1 I_18171 (I105306,I2683,I311544,I311635,);
nand I_18172 (I311643,I311635,I105300);
not I_18173 (I311660,I105300);
not I_18174 (I311677,I105297);
nand I_18175 (I311694,I105291,I105288);
and I_18176 (I311711,I105291,I105288);
not I_18177 (I311728,I105303);
nand I_18178 (I311745,I311728,I311677);
nor I_18179 (I311518,I311745,I311643);
nor I_18180 (I311776,I311660,I311745);
nand I_18181 (I311521,I311711,I311776);
not I_18182 (I311807,I105315);
nor I_18183 (I311824,I311807,I105291);
nor I_18184 (I311841,I311824,I105303);
nor I_18185 (I311858,I311609,I311841);
DFFARX1 I_18186 (I311858,I2683,I311544,I311530,);
not I_18187 (I311889,I311824);
DFFARX1 I_18188 (I311889,I2683,I311544,I311533,);
and I_18189 (I311527,I311635,I311824);
nor I_18190 (I311934,I311807,I105312);
and I_18191 (I311951,I311934,I105288);
or I_18192 (I311968,I311951,I105294);
DFFARX1 I_18193 (I311968,I2683,I311544,I311994,);
nor I_18194 (I312002,I311994,I311728);
DFFARX1 I_18195 (I312002,I2683,I311544,I311515,);
nand I_18196 (I312033,I311994,I311635);
nand I_18197 (I312050,I311728,I312033);
nor I_18198 (I311524,I312050,I311694);
not I_18199 (I312105,I2690);
DFFARX1 I_18200 (I92661,I2683,I312105,I312131,);
DFFARX1 I_18201 (I312131,I2683,I312105,I312148,);
not I_18202 (I312097,I312148);
not I_18203 (I312170,I312131);
DFFARX1 I_18204 (I92658,I2683,I312105,I312196,);
nand I_18205 (I312204,I312196,I92652);
not I_18206 (I312221,I92652);
not I_18207 (I312238,I92649);
nand I_18208 (I312255,I92643,I92640);
and I_18209 (I312272,I92643,I92640);
not I_18210 (I312289,I92655);
nand I_18211 (I312306,I312289,I312238);
nor I_18212 (I312079,I312306,I312204);
nor I_18213 (I312337,I312221,I312306);
nand I_18214 (I312082,I312272,I312337);
not I_18215 (I312368,I92667);
nor I_18216 (I312385,I312368,I92643);
nor I_18217 (I312402,I312385,I92655);
nor I_18218 (I312419,I312170,I312402);
DFFARX1 I_18219 (I312419,I2683,I312105,I312091,);
not I_18220 (I312450,I312385);
DFFARX1 I_18221 (I312450,I2683,I312105,I312094,);
and I_18222 (I312088,I312196,I312385);
nor I_18223 (I312495,I312368,I92664);
and I_18224 (I312512,I312495,I92640);
or I_18225 (I312529,I312512,I92646);
DFFARX1 I_18226 (I312529,I2683,I312105,I312555,);
nor I_18227 (I312563,I312555,I312289);
DFFARX1 I_18228 (I312563,I2683,I312105,I312076,);
nand I_18229 (I312594,I312555,I312196);
nand I_18230 (I312611,I312289,I312594);
nor I_18231 (I312085,I312611,I312255);
not I_18232 (I312666,I2690);
DFFARX1 I_18233 (I2212,I2683,I312666,I312692,);
DFFARX1 I_18234 (I312692,I2683,I312666,I312709,);
not I_18235 (I312658,I312709);
not I_18236 (I312731,I312692);
DFFARX1 I_18237 (I1780,I2683,I312666,I312757,);
nand I_18238 (I312765,I312757,I2580);
not I_18239 (I312782,I2580);
not I_18240 (I312799,I2564);
nand I_18241 (I312816,I1860,I1676);
and I_18242 (I312833,I1860,I1676);
not I_18243 (I312850,I2052);
nand I_18244 (I312867,I312850,I312799);
nor I_18245 (I312640,I312867,I312765);
nor I_18246 (I312898,I312782,I312867);
nand I_18247 (I312643,I312833,I312898);
not I_18248 (I312929,I2404);
nor I_18249 (I312946,I312929,I1860);
nor I_18250 (I312963,I312946,I2052);
nor I_18251 (I312980,I312731,I312963);
DFFARX1 I_18252 (I312980,I2683,I312666,I312652,);
not I_18253 (I313011,I312946);
DFFARX1 I_18254 (I313011,I2683,I312666,I312655,);
and I_18255 (I312649,I312757,I312946);
nor I_18256 (I313056,I312929,I1388);
and I_18257 (I313073,I313056,I1708);
or I_18258 (I313090,I313073,I1524);
DFFARX1 I_18259 (I313090,I2683,I312666,I313116,);
nor I_18260 (I313124,I313116,I312850);
DFFARX1 I_18261 (I313124,I2683,I312666,I312637,);
nand I_18262 (I313155,I313116,I312757);
nand I_18263 (I313172,I312850,I313155);
nor I_18264 (I312646,I313172,I312816);
not I_18265 (I313227,I2690);
DFFARX1 I_18266 (I365955,I2683,I313227,I313253,);
DFFARX1 I_18267 (I313253,I2683,I313227,I313270,);
not I_18268 (I313219,I313270);
not I_18269 (I313292,I313253);
DFFARX1 I_18270 (I365961,I2683,I313227,I313318,);
nand I_18271 (I313326,I313318,I365970);
not I_18272 (I313343,I365970);
not I_18273 (I313360,I365949);
nand I_18274 (I313377,I365952,I365952);
and I_18275 (I313394,I365952,I365952);
not I_18276 (I313411,I365964);
nand I_18277 (I313428,I313411,I313360);
nor I_18278 (I313201,I313428,I313326);
nor I_18279 (I313459,I313343,I313428);
nand I_18280 (I313204,I313394,I313459);
not I_18281 (I313490,I365958);
nor I_18282 (I313507,I313490,I365952);
nor I_18283 (I313524,I313507,I365964);
nor I_18284 (I313541,I313292,I313524);
DFFARX1 I_18285 (I313541,I2683,I313227,I313213,);
not I_18286 (I313572,I313507);
DFFARX1 I_18287 (I313572,I2683,I313227,I313216,);
and I_18288 (I313210,I313318,I313507);
nor I_18289 (I313617,I313490,I365973);
and I_18290 (I313634,I313617,I365949);
or I_18291 (I313651,I313634,I365967);
DFFARX1 I_18292 (I313651,I2683,I313227,I313677,);
nor I_18293 (I313685,I313677,I313411);
DFFARX1 I_18294 (I313685,I2683,I313227,I313198,);
nand I_18295 (I313716,I313677,I313318);
nand I_18296 (I313733,I313411,I313716);
nor I_18297 (I313207,I313733,I313377);
not I_18298 (I313788,I2690);
DFFARX1 I_18299 (I218086,I2683,I313788,I313814,);
DFFARX1 I_18300 (I313814,I2683,I313788,I313831,);
not I_18301 (I313780,I313831);
not I_18302 (I313853,I313814);
DFFARX1 I_18303 (I218098,I2683,I313788,I313879,);
nand I_18304 (I313887,I313879,I218107);
not I_18305 (I313904,I218107);
not I_18306 (I313921,I218089);
nand I_18307 (I313938,I218092,I218083);
and I_18308 (I313955,I218092,I218083);
not I_18309 (I313972,I218101);
nand I_18310 (I313989,I313972,I313921);
nor I_18311 (I313762,I313989,I313887);
nor I_18312 (I314020,I313904,I313989);
nand I_18313 (I313765,I313955,I314020);
not I_18314 (I314051,I218104);
nor I_18315 (I314068,I314051,I218092);
nor I_18316 (I314085,I314068,I218101);
nor I_18317 (I314102,I313853,I314085);
DFFARX1 I_18318 (I314102,I2683,I313788,I313774,);
not I_18319 (I314133,I314068);
DFFARX1 I_18320 (I314133,I2683,I313788,I313777,);
and I_18321 (I313771,I313879,I314068);
nor I_18322 (I314178,I314051,I218083);
and I_18323 (I314195,I314178,I218095);
or I_18324 (I314212,I314195,I218086);
DFFARX1 I_18325 (I314212,I2683,I313788,I314238,);
nor I_18326 (I314246,I314238,I313972);
DFFARX1 I_18327 (I314246,I2683,I313788,I313759,);
nand I_18328 (I314277,I314238,I313879);
nand I_18329 (I314294,I313972,I314277);
nor I_18330 (I313768,I314294,I313938);
not I_18331 (I314349,I2690);
DFFARX1 I_18332 (I20963,I2683,I314349,I314375,);
DFFARX1 I_18333 (I314375,I2683,I314349,I314392,);
not I_18334 (I314341,I314392);
not I_18335 (I314414,I314375);
DFFARX1 I_18336 (I20951,I2683,I314349,I314440,);
nand I_18337 (I314448,I314440,I20966);
not I_18338 (I314465,I20966);
not I_18339 (I314482,I20954);
nand I_18340 (I314499,I20975,I20969);
and I_18341 (I314516,I20975,I20969);
not I_18342 (I314533,I20957);
nand I_18343 (I314550,I314533,I314482);
nor I_18344 (I314323,I314550,I314448);
nor I_18345 (I314581,I314465,I314550);
nand I_18346 (I314326,I314516,I314581);
not I_18347 (I314612,I20960);
nor I_18348 (I314629,I314612,I20975);
nor I_18349 (I314646,I314629,I20957);
nor I_18350 (I314663,I314414,I314646);
DFFARX1 I_18351 (I314663,I2683,I314349,I314335,);
not I_18352 (I314694,I314629);
DFFARX1 I_18353 (I314694,I2683,I314349,I314338,);
and I_18354 (I314332,I314440,I314629);
nor I_18355 (I314739,I314612,I20954);
and I_18356 (I314756,I314739,I20951);
or I_18357 (I314773,I314756,I20972);
DFFARX1 I_18358 (I314773,I2683,I314349,I314799,);
nor I_18359 (I314807,I314799,I314533);
DFFARX1 I_18360 (I314807,I2683,I314349,I314320,);
nand I_18361 (I314838,I314799,I314440);
nand I_18362 (I314855,I314533,I314838);
nor I_18363 (I314329,I314855,I314499);
not I_18364 (I314910,I2690);
DFFARX1 I_18365 (I108471,I2683,I314910,I314936,);
DFFARX1 I_18366 (I314936,I2683,I314910,I314953,);
not I_18367 (I314902,I314953);
not I_18368 (I314975,I314936);
DFFARX1 I_18369 (I108468,I2683,I314910,I315001,);
nand I_18370 (I315009,I315001,I108462);
not I_18371 (I315026,I108462);
not I_18372 (I315043,I108459);
nand I_18373 (I315060,I108453,I108450);
and I_18374 (I315077,I108453,I108450);
not I_18375 (I315094,I108465);
nand I_18376 (I315111,I315094,I315043);
nor I_18377 (I314884,I315111,I315009);
nor I_18378 (I315142,I315026,I315111);
nand I_18379 (I314887,I315077,I315142);
not I_18380 (I315173,I108477);
nor I_18381 (I315190,I315173,I108453);
nor I_18382 (I315207,I315190,I108465);
nor I_18383 (I315224,I314975,I315207);
DFFARX1 I_18384 (I315224,I2683,I314910,I314896,);
not I_18385 (I315255,I315190);
DFFARX1 I_18386 (I315255,I2683,I314910,I314899,);
and I_18387 (I314893,I315001,I315190);
nor I_18388 (I315300,I315173,I108474);
and I_18389 (I315317,I315300,I108450);
or I_18390 (I315334,I315317,I108456);
DFFARX1 I_18391 (I315334,I2683,I314910,I315360,);
nor I_18392 (I315368,I315360,I315094);
DFFARX1 I_18393 (I315368,I2683,I314910,I314881,);
nand I_18394 (I315399,I315360,I315001);
nand I_18395 (I315416,I315094,I315399);
nor I_18396 (I314890,I315416,I315060);
not I_18397 (I315471,I2690);
DFFARX1 I_18398 (I136711,I2683,I315471,I315497,);
DFFARX1 I_18399 (I315497,I2683,I315471,I315514,);
not I_18400 (I315463,I315514);
not I_18401 (I315536,I315497);
DFFARX1 I_18402 (I136699,I2683,I315471,I315562,);
nand I_18403 (I315570,I315562,I136705);
not I_18404 (I315587,I136705);
not I_18405 (I315604,I136702);
nand I_18406 (I315621,I136690,I136687);
and I_18407 (I315638,I136690,I136687);
not I_18408 (I315655,I136714);
nand I_18409 (I315672,I315655,I315604);
nor I_18410 (I315445,I315672,I315570);
nor I_18411 (I315703,I315587,I315672);
nand I_18412 (I315448,I315638,I315703);
not I_18413 (I315734,I136687);
nor I_18414 (I315751,I315734,I136690);
nor I_18415 (I315768,I315751,I136714);
nor I_18416 (I315785,I315536,I315768);
DFFARX1 I_18417 (I315785,I2683,I315471,I315457,);
not I_18418 (I315816,I315751);
DFFARX1 I_18419 (I315816,I2683,I315471,I315460,);
and I_18420 (I315454,I315562,I315751);
nor I_18421 (I315861,I315734,I136696);
and I_18422 (I315878,I315861,I136693);
or I_18423 (I315895,I315878,I136708);
DFFARX1 I_18424 (I315895,I2683,I315471,I315921,);
nor I_18425 (I315929,I315921,I315655);
DFFARX1 I_18426 (I315929,I2683,I315471,I315442,);
nand I_18427 (I315960,I315921,I315562);
nand I_18428 (I315977,I315655,I315960);
nor I_18429 (I315451,I315977,I315621);
not I_18430 (I316032,I2690);
DFFARX1 I_18431 (I62587,I2683,I316032,I316058,);
DFFARX1 I_18432 (I316058,I2683,I316032,I316075,);
not I_18433 (I316024,I316075);
not I_18434 (I316097,I316058);
DFFARX1 I_18435 (I62602,I2683,I316032,I316123,);
nand I_18436 (I316131,I316123,I62584);
not I_18437 (I316148,I62584);
not I_18438 (I316165,I62593);
nand I_18439 (I316182,I62599,I62590);
and I_18440 (I316199,I62599,I62590);
not I_18441 (I316216,I62587);
nand I_18442 (I316233,I316216,I316165);
nor I_18443 (I316006,I316233,I316131);
nor I_18444 (I316264,I316148,I316233);
nand I_18445 (I316009,I316199,I316264);
not I_18446 (I316295,I62584);
nor I_18447 (I316312,I316295,I62599);
nor I_18448 (I316329,I316312,I62587);
nor I_18449 (I316346,I316097,I316329);
DFFARX1 I_18450 (I316346,I2683,I316032,I316018,);
not I_18451 (I316377,I316312);
DFFARX1 I_18452 (I316377,I2683,I316032,I316021,);
and I_18453 (I316015,I316123,I316312);
nor I_18454 (I316422,I316295,I62608);
and I_18455 (I316439,I316422,I62605);
or I_18456 (I316456,I316439,I62596);
DFFARX1 I_18457 (I316456,I2683,I316032,I316482,);
nor I_18458 (I316490,I316482,I316216);
DFFARX1 I_18459 (I316490,I2683,I316032,I316003,);
nand I_18460 (I316521,I316482,I316123);
nand I_18461 (I316538,I316216,I316521);
nor I_18462 (I316012,I316538,I316182);
not I_18463 (I316593,I2690);
DFFARX1 I_18464 (I413479,I2683,I316593,I316619,);
DFFARX1 I_18465 (I316619,I2683,I316593,I316636,);
not I_18466 (I316585,I316636);
not I_18467 (I316658,I316619);
DFFARX1 I_18468 (I413473,I2683,I316593,I316684,);
nand I_18469 (I316692,I316684,I413464);
not I_18470 (I316709,I413464);
not I_18471 (I316726,I413491);
nand I_18472 (I316743,I413476,I413485);
and I_18473 (I316760,I413476,I413485);
not I_18474 (I316777,I413470);
nand I_18475 (I316794,I316777,I316726);
nor I_18476 (I316567,I316794,I316692);
nor I_18477 (I316825,I316709,I316794);
nand I_18478 (I316570,I316760,I316825);
not I_18479 (I316856,I413488);
nor I_18480 (I316873,I316856,I413476);
nor I_18481 (I316890,I316873,I413470);
nor I_18482 (I316907,I316658,I316890);
DFFARX1 I_18483 (I316907,I2683,I316593,I316579,);
not I_18484 (I316938,I316873);
DFFARX1 I_18485 (I316938,I2683,I316593,I316582,);
and I_18486 (I316576,I316684,I316873);
nor I_18487 (I316983,I316856,I413482);
and I_18488 (I317000,I316983,I413464);
or I_18489 (I317017,I317000,I413467);
DFFARX1 I_18490 (I317017,I2683,I316593,I317043,);
nor I_18491 (I317051,I317043,I316777);
DFFARX1 I_18492 (I317051,I2683,I316593,I316564,);
nand I_18493 (I317082,I317043,I316684);
nand I_18494 (I317099,I316777,I317082);
nor I_18495 (I316573,I317099,I316743);
not I_18496 (I317154,I2690);
DFFARX1 I_18497 (I55447,I2683,I317154,I317180,);
DFFARX1 I_18498 (I317180,I2683,I317154,I317197,);
not I_18499 (I317146,I317197);
not I_18500 (I317219,I317180);
DFFARX1 I_18501 (I55462,I2683,I317154,I317245,);
nand I_18502 (I317253,I317245,I55444);
not I_18503 (I317270,I55444);
not I_18504 (I317287,I55453);
nand I_18505 (I317304,I55459,I55450);
and I_18506 (I317321,I55459,I55450);
not I_18507 (I317338,I55447);
nand I_18508 (I317355,I317338,I317287);
nor I_18509 (I317128,I317355,I317253);
nor I_18510 (I317386,I317270,I317355);
nand I_18511 (I317131,I317321,I317386);
not I_18512 (I317417,I55444);
nor I_18513 (I317434,I317417,I55459);
nor I_18514 (I317451,I317434,I55447);
nor I_18515 (I317468,I317219,I317451);
DFFARX1 I_18516 (I317468,I2683,I317154,I317140,);
not I_18517 (I317499,I317434);
DFFARX1 I_18518 (I317499,I2683,I317154,I317143,);
and I_18519 (I317137,I317245,I317434);
nor I_18520 (I317544,I317417,I55468);
and I_18521 (I317561,I317544,I55465);
or I_18522 (I317578,I317561,I55456);
DFFARX1 I_18523 (I317578,I2683,I317154,I317604,);
nor I_18524 (I317612,I317604,I317338);
DFFARX1 I_18525 (I317612,I2683,I317154,I317125,);
nand I_18526 (I317643,I317604,I317245);
nand I_18527 (I317660,I317338,I317643);
nor I_18528 (I317134,I317660,I317304);
not I_18529 (I317715,I2690);
DFFARX1 I_18530 (I193229,I2683,I317715,I317741,);
DFFARX1 I_18531 (I317741,I2683,I317715,I317758,);
not I_18532 (I317707,I317758);
not I_18533 (I317780,I317741);
DFFARX1 I_18534 (I193244,I2683,I317715,I317806,);
nand I_18535 (I317814,I317806,I193235);
not I_18536 (I317831,I193235);
not I_18537 (I317848,I193241);
nand I_18538 (I317865,I193238,I193247);
and I_18539 (I317882,I193238,I193247);
not I_18540 (I317899,I193232);
nand I_18541 (I317916,I317899,I317848);
nor I_18542 (I317689,I317916,I317814);
nor I_18543 (I317947,I317831,I317916);
nand I_18544 (I317692,I317882,I317947);
not I_18545 (I317978,I193229);
nor I_18546 (I317995,I317978,I193238);
nor I_18547 (I318012,I317995,I193232);
nor I_18548 (I318029,I317780,I318012);
DFFARX1 I_18549 (I318029,I2683,I317715,I317701,);
not I_18550 (I318060,I317995);
DFFARX1 I_18551 (I318060,I2683,I317715,I317704,);
and I_18552 (I317698,I317806,I317995);
nor I_18553 (I318105,I317978,I193253);
and I_18554 (I318122,I318105,I193232);
or I_18555 (I318139,I318122,I193250);
DFFARX1 I_18556 (I318139,I2683,I317715,I318165,);
nor I_18557 (I318173,I318165,I317899);
DFFARX1 I_18558 (I318173,I2683,I317715,I317686,);
nand I_18559 (I318204,I318165,I317806);
nand I_18560 (I318221,I317899,I318204);
nor I_18561 (I317695,I318221,I317865);
not I_18562 (I318276,I2690);
DFFARX1 I_18563 (I327340,I2683,I318276,I318302,);
DFFARX1 I_18564 (I318302,I2683,I318276,I318319,);
not I_18565 (I318268,I318319);
not I_18566 (I318341,I318302);
DFFARX1 I_18567 (I327331,I2683,I318276,I318367,);
nand I_18568 (I318375,I318367,I327328);
not I_18569 (I318392,I327328);
not I_18570 (I318409,I327337);
nand I_18571 (I318426,I327346,I327328);
and I_18572 (I318443,I327346,I327328);
not I_18573 (I318460,I327325);
nand I_18574 (I318477,I318460,I318409);
nor I_18575 (I318250,I318477,I318375);
nor I_18576 (I318508,I318392,I318477);
nand I_18577 (I318253,I318443,I318508);
not I_18578 (I318539,I327334);
nor I_18579 (I318556,I318539,I327346);
nor I_18580 (I318573,I318556,I327325);
nor I_18581 (I318590,I318341,I318573);
DFFARX1 I_18582 (I318590,I2683,I318276,I318262,);
not I_18583 (I318621,I318556);
DFFARX1 I_18584 (I318621,I2683,I318276,I318265,);
and I_18585 (I318259,I318367,I318556);
nor I_18586 (I318666,I318539,I327349);
and I_18587 (I318683,I318666,I327325);
or I_18588 (I318700,I318683,I327343);
DFFARX1 I_18589 (I318700,I2683,I318276,I318726,);
nor I_18590 (I318734,I318726,I318460);
DFFARX1 I_18591 (I318734,I2683,I318276,I318247,);
nand I_18592 (I318765,I318726,I318367);
nand I_18593 (I318782,I318460,I318765);
nor I_18594 (I318256,I318782,I318426);
not I_18595 (I318837,I2690);
DFFARX1 I_18596 (I341212,I2683,I318837,I318863,);
DFFARX1 I_18597 (I318863,I2683,I318837,I318880,);
not I_18598 (I318829,I318880);
not I_18599 (I318902,I318863);
DFFARX1 I_18600 (I341203,I2683,I318837,I318928,);
nand I_18601 (I318936,I318928,I341200);
not I_18602 (I318953,I341200);
not I_18603 (I318970,I341209);
nand I_18604 (I318987,I341218,I341200);
and I_18605 (I319004,I341218,I341200);
not I_18606 (I319021,I341197);
nand I_18607 (I319038,I319021,I318970);
nor I_18608 (I318811,I319038,I318936);
nor I_18609 (I319069,I318953,I319038);
nand I_18610 (I318814,I319004,I319069);
not I_18611 (I319100,I341206);
nor I_18612 (I319117,I319100,I341218);
nor I_18613 (I319134,I319117,I341197);
nor I_18614 (I319151,I318902,I319134);
DFFARX1 I_18615 (I319151,I2683,I318837,I318823,);
not I_18616 (I319182,I319117);
DFFARX1 I_18617 (I319182,I2683,I318837,I318826,);
and I_18618 (I318820,I318928,I319117);
nor I_18619 (I319227,I319100,I341221);
and I_18620 (I319244,I319227,I341197);
or I_18621 (I319261,I319244,I341215);
DFFARX1 I_18622 (I319261,I2683,I318837,I319287,);
nor I_18623 (I319295,I319287,I319021);
DFFARX1 I_18624 (I319295,I2683,I318837,I318808,);
nand I_18625 (I319326,I319287,I318928);
nand I_18626 (I319343,I319021,I319326);
nor I_18627 (I318817,I319343,I318987);
not I_18628 (I319398,I2690);
DFFARX1 I_18629 (I253452,I2683,I319398,I319424,);
DFFARX1 I_18630 (I319424,I2683,I319398,I319441,);
not I_18631 (I319390,I319441);
not I_18632 (I319463,I319424);
DFFARX1 I_18633 (I253449,I2683,I319398,I319489,);
nand I_18634 (I319497,I319489,I253464);
not I_18635 (I319514,I253464);
not I_18636 (I319531,I253461);
nand I_18637 (I319548,I253458,I253446);
and I_18638 (I319565,I253458,I253446);
not I_18639 (I319582,I253443);
nand I_18640 (I319599,I319582,I319531);
nor I_18641 (I319372,I319599,I319497);
nor I_18642 (I319630,I319514,I319599);
nand I_18643 (I319375,I319565,I319630);
not I_18644 (I319661,I253449);
nor I_18645 (I319678,I319661,I253458);
nor I_18646 (I319695,I319678,I253443);
nor I_18647 (I319712,I319463,I319695);
DFFARX1 I_18648 (I319712,I2683,I319398,I319384,);
not I_18649 (I319743,I319678);
DFFARX1 I_18650 (I319743,I2683,I319398,I319387,);
and I_18651 (I319381,I319489,I319678);
nor I_18652 (I319788,I319661,I253455);
and I_18653 (I319805,I319788,I253443);
or I_18654 (I319822,I319805,I253446);
DFFARX1 I_18655 (I319822,I2683,I319398,I319848,);
nor I_18656 (I319856,I319848,I319582);
DFFARX1 I_18657 (I319856,I2683,I319398,I319369,);
nand I_18658 (I319887,I319848,I319489);
nand I_18659 (I319904,I319582,I319887);
nor I_18660 (I319378,I319904,I319548);
not I_18661 (I319959,I2690);
DFFARX1 I_18662 (I106890,I2683,I319959,I319985,);
DFFARX1 I_18663 (I319985,I2683,I319959,I320002,);
not I_18664 (I319951,I320002);
not I_18665 (I320024,I319985);
DFFARX1 I_18666 (I106887,I2683,I319959,I320050,);
nand I_18667 (I320058,I320050,I106881);
not I_18668 (I320075,I106881);
not I_18669 (I320092,I106878);
nand I_18670 (I320109,I106872,I106869);
and I_18671 (I320126,I106872,I106869);
not I_18672 (I320143,I106884);
nand I_18673 (I320160,I320143,I320092);
nor I_18674 (I319933,I320160,I320058);
nor I_18675 (I320191,I320075,I320160);
nand I_18676 (I319936,I320126,I320191);
not I_18677 (I320222,I106896);
nor I_18678 (I320239,I320222,I106872);
nor I_18679 (I320256,I320239,I106884);
nor I_18680 (I320273,I320024,I320256);
DFFARX1 I_18681 (I320273,I2683,I319959,I319945,);
not I_18682 (I320304,I320239);
DFFARX1 I_18683 (I320304,I2683,I319959,I319948,);
and I_18684 (I319942,I320050,I320239);
nor I_18685 (I320349,I320222,I106893);
and I_18686 (I320366,I320349,I106869);
or I_18687 (I320383,I320366,I106875);
DFFARX1 I_18688 (I320383,I2683,I319959,I320409,);
nor I_18689 (I320417,I320409,I320143);
DFFARX1 I_18690 (I320417,I2683,I319959,I319930,);
nand I_18691 (I320448,I320409,I320050);
nand I_18692 (I320465,I320143,I320448);
nor I_18693 (I319939,I320465,I320109);
not I_18694 (I320520,I2690);
DFFARX1 I_18695 (I351616,I2683,I320520,I320546,);
DFFARX1 I_18696 (I320546,I2683,I320520,I320563,);
not I_18697 (I320512,I320563);
not I_18698 (I320585,I320546);
DFFARX1 I_18699 (I351607,I2683,I320520,I320611,);
nand I_18700 (I320619,I320611,I351604);
not I_18701 (I320636,I351604);
not I_18702 (I320653,I351613);
nand I_18703 (I320670,I351622,I351604);
and I_18704 (I320687,I351622,I351604);
not I_18705 (I320704,I351601);
nand I_18706 (I320721,I320704,I320653);
nor I_18707 (I320494,I320721,I320619);
nor I_18708 (I320752,I320636,I320721);
nand I_18709 (I320497,I320687,I320752);
not I_18710 (I320783,I351610);
nor I_18711 (I320800,I320783,I351622);
nor I_18712 (I320817,I320800,I351601);
nor I_18713 (I320834,I320585,I320817);
DFFARX1 I_18714 (I320834,I2683,I320520,I320506,);
not I_18715 (I320865,I320800);
DFFARX1 I_18716 (I320865,I2683,I320520,I320509,);
and I_18717 (I320503,I320611,I320800);
nor I_18718 (I320910,I320783,I351625);
and I_18719 (I320927,I320910,I351601);
or I_18720 (I320944,I320927,I351619);
DFFARX1 I_18721 (I320944,I2683,I320520,I320970,);
nor I_18722 (I320978,I320970,I320704);
DFFARX1 I_18723 (I320978,I2683,I320520,I320491,);
nand I_18724 (I321009,I320970,I320611);
nand I_18725 (I321026,I320704,I321009);
nor I_18726 (I320500,I321026,I320670);
not I_18727 (I321081,I2690);
DFFARX1 I_18728 (I63777,I2683,I321081,I321107,);
DFFARX1 I_18729 (I321107,I2683,I321081,I321124,);
not I_18730 (I321073,I321124);
not I_18731 (I321146,I321107);
DFFARX1 I_18732 (I63792,I2683,I321081,I321172,);
nand I_18733 (I321180,I321172,I63774);
not I_18734 (I321197,I63774);
not I_18735 (I321214,I63783);
nand I_18736 (I321231,I63789,I63780);
and I_18737 (I321248,I63789,I63780);
not I_18738 (I321265,I63777);
nand I_18739 (I321282,I321265,I321214);
nor I_18740 (I321055,I321282,I321180);
nor I_18741 (I321313,I321197,I321282);
nand I_18742 (I321058,I321248,I321313);
not I_18743 (I321344,I63774);
nor I_18744 (I321361,I321344,I63789);
nor I_18745 (I321378,I321361,I63777);
nor I_18746 (I321395,I321146,I321378);
DFFARX1 I_18747 (I321395,I2683,I321081,I321067,);
not I_18748 (I321426,I321361);
DFFARX1 I_18749 (I321426,I2683,I321081,I321070,);
and I_18750 (I321064,I321172,I321361);
nor I_18751 (I321471,I321344,I63798);
and I_18752 (I321488,I321471,I63795);
or I_18753 (I321505,I321488,I63786);
DFFARX1 I_18754 (I321505,I2683,I321081,I321531,);
nor I_18755 (I321539,I321531,I321265);
DFFARX1 I_18756 (I321539,I2683,I321081,I321052,);
nand I_18757 (I321570,I321531,I321172);
nand I_18758 (I321587,I321265,I321570);
nor I_18759 (I321061,I321587,I321231);
not I_18760 (I321642,I2690);
DFFARX1 I_18761 (I240804,I2683,I321642,I321668,);
DFFARX1 I_18762 (I321668,I2683,I321642,I321685,);
not I_18763 (I321634,I321685);
not I_18764 (I321707,I321668);
DFFARX1 I_18765 (I240801,I2683,I321642,I321733,);
nand I_18766 (I321741,I321733,I240816);
not I_18767 (I321758,I240816);
not I_18768 (I321775,I240813);
nand I_18769 (I321792,I240810,I240798);
and I_18770 (I321809,I240810,I240798);
not I_18771 (I321826,I240795);
nand I_18772 (I321843,I321826,I321775);
nor I_18773 (I321616,I321843,I321741);
nor I_18774 (I321874,I321758,I321843);
nand I_18775 (I321619,I321809,I321874);
not I_18776 (I321905,I240801);
nor I_18777 (I321922,I321905,I240810);
nor I_18778 (I321939,I321922,I240795);
nor I_18779 (I321956,I321707,I321939);
DFFARX1 I_18780 (I321956,I2683,I321642,I321628,);
not I_18781 (I321987,I321922);
DFFARX1 I_18782 (I321987,I2683,I321642,I321631,);
and I_18783 (I321625,I321733,I321922);
nor I_18784 (I322032,I321905,I240807);
and I_18785 (I322049,I322032,I240795);
or I_18786 (I322066,I322049,I240798);
DFFARX1 I_18787 (I322066,I2683,I321642,I322092,);
nor I_18788 (I322100,I322092,I321826);
DFFARX1 I_18789 (I322100,I2683,I321642,I321613,);
nand I_18790 (I322131,I322092,I321733);
nand I_18791 (I322148,I321826,I322131);
nor I_18792 (I321622,I322148,I321792);
not I_18793 (I322203,I2690);
DFFARX1 I_18794 (I10956,I2683,I322203,I322229,);
DFFARX1 I_18795 (I322229,I2683,I322203,I322246,);
not I_18796 (I322195,I322246);
not I_18797 (I322268,I322229);
DFFARX1 I_18798 (I10941,I2683,I322203,I322294,);
nand I_18799 (I322302,I322294,I10953);
not I_18800 (I322319,I10953);
not I_18801 (I322336,I10959);
nand I_18802 (I322353,I10947,I10938);
and I_18803 (I322370,I10947,I10938);
not I_18804 (I322387,I10944);
nand I_18805 (I322404,I322387,I322336);
nor I_18806 (I322177,I322404,I322302);
nor I_18807 (I322435,I322319,I322404);
nand I_18808 (I322180,I322370,I322435);
not I_18809 (I322466,I10950);
nor I_18810 (I322483,I322466,I10947);
nor I_18811 (I322500,I322483,I10944);
nor I_18812 (I322517,I322268,I322500);
DFFARX1 I_18813 (I322517,I2683,I322203,I322189,);
not I_18814 (I322548,I322483);
DFFARX1 I_18815 (I322548,I2683,I322203,I322192,);
and I_18816 (I322186,I322294,I322483);
nor I_18817 (I322593,I322466,I10938);
and I_18818 (I322610,I322593,I10962);
or I_18819 (I322627,I322610,I10941);
DFFARX1 I_18820 (I322627,I2683,I322203,I322653,);
nor I_18821 (I322661,I322653,I322387);
DFFARX1 I_18822 (I322661,I2683,I322203,I322174,);
nand I_18823 (I322692,I322653,I322294);
nand I_18824 (I322709,I322387,I322692);
nor I_18825 (I322183,I322709,I322353);
not I_18826 (I322764,I2690);
DFFARX1 I_18827 (I199590,I2683,I322764,I322790,);
DFFARX1 I_18828 (I322790,I2683,I322764,I322807,);
not I_18829 (I322756,I322807);
not I_18830 (I322829,I322790);
DFFARX1 I_18831 (I199602,I2683,I322764,I322855,);
nand I_18832 (I322863,I322855,I199611);
not I_18833 (I322880,I199611);
not I_18834 (I322897,I199593);
nand I_18835 (I322914,I199596,I199587);
and I_18836 (I322931,I199596,I199587);
not I_18837 (I322948,I199605);
nand I_18838 (I322965,I322948,I322897);
nor I_18839 (I322738,I322965,I322863);
nor I_18840 (I322996,I322880,I322965);
nand I_18841 (I322741,I322931,I322996);
not I_18842 (I323027,I199608);
nor I_18843 (I323044,I323027,I199596);
nor I_18844 (I323061,I323044,I199605);
nor I_18845 (I323078,I322829,I323061);
DFFARX1 I_18846 (I323078,I2683,I322764,I322750,);
not I_18847 (I323109,I323044);
DFFARX1 I_18848 (I323109,I2683,I322764,I322753,);
and I_18849 (I322747,I322855,I323044);
nor I_18850 (I323154,I323027,I199587);
and I_18851 (I323171,I323154,I199599);
or I_18852 (I323188,I323171,I199590);
DFFARX1 I_18853 (I323188,I2683,I322764,I323214,);
nor I_18854 (I323222,I323214,I322948);
DFFARX1 I_18855 (I323222,I2683,I322764,I322735,);
nand I_18856 (I323253,I323214,I322855);
nand I_18857 (I323270,I322948,I323253);
nor I_18858 (I322744,I323270,I322914);
not I_18859 (I323325,I2690);
DFFARX1 I_18860 (I340056,I2683,I323325,I323351,);
DFFARX1 I_18861 (I323351,I2683,I323325,I323368,);
not I_18862 (I323317,I323368);
not I_18863 (I323390,I323351);
DFFARX1 I_18864 (I340047,I2683,I323325,I323416,);
nand I_18865 (I323424,I323416,I340044);
not I_18866 (I323441,I340044);
not I_18867 (I323458,I340053);
nand I_18868 (I323475,I340062,I340044);
and I_18869 (I323492,I340062,I340044);
not I_18870 (I323509,I340041);
nand I_18871 (I323526,I323509,I323458);
nor I_18872 (I323299,I323526,I323424);
nor I_18873 (I323557,I323441,I323526);
nand I_18874 (I323302,I323492,I323557);
not I_18875 (I323588,I340050);
nor I_18876 (I323605,I323588,I340062);
nor I_18877 (I323622,I323605,I340041);
nor I_18878 (I323639,I323390,I323622);
DFFARX1 I_18879 (I323639,I2683,I323325,I323311,);
not I_18880 (I323670,I323605);
DFFARX1 I_18881 (I323670,I2683,I323325,I323314,);
and I_18882 (I323308,I323416,I323605);
nor I_18883 (I323715,I323588,I340065);
and I_18884 (I323732,I323715,I340041);
or I_18885 (I323749,I323732,I340059);
DFFARX1 I_18886 (I323749,I2683,I323325,I323775,);
nor I_18887 (I323783,I323775,I323509);
DFFARX1 I_18888 (I323783,I2683,I323325,I323296,);
nand I_18889 (I323814,I323775,I323416);
nand I_18890 (I323831,I323509,I323814);
nor I_18891 (I323305,I323831,I323475);
not I_18892 (I323889,I2690);
DFFARX1 I_18893 (I223300,I2683,I323889,I323915,);
and I_18894 (I323923,I323915,I223288);
DFFARX1 I_18895 (I323923,I2683,I323889,I323872,);
DFFARX1 I_18896 (I223291,I2683,I323889,I323963,);
not I_18897 (I323971,I223285);
not I_18898 (I323988,I223309);
nand I_18899 (I324005,I323988,I323971);
nor I_18900 (I323860,I323963,I324005);
DFFARX1 I_18901 (I324005,I2683,I323889,I324045,);
not I_18902 (I323881,I324045);
not I_18903 (I324067,I223297);
nand I_18904 (I324084,I323988,I324067);
DFFARX1 I_18905 (I324084,I2683,I323889,I324110,);
not I_18906 (I324118,I324110);
not I_18907 (I324135,I223306);
nand I_18908 (I324152,I324135,I223303);
and I_18909 (I324169,I323971,I324152);
nor I_18910 (I324186,I324084,I324169);
DFFARX1 I_18911 (I324186,I2683,I323889,I323857,);
DFFARX1 I_18912 (I324169,I2683,I323889,I323878,);
nor I_18913 (I324231,I223306,I223294);
nor I_18914 (I323869,I324084,I324231);
or I_18915 (I324262,I223306,I223294);
nor I_18916 (I324279,I223285,I223288);
DFFARX1 I_18917 (I324279,I2683,I323889,I324305,);
not I_18918 (I324313,I324305);
nor I_18919 (I323875,I324313,I324118);
nand I_18920 (I324344,I324313,I323963);
not I_18921 (I324361,I223285);
nand I_18922 (I324378,I324361,I324067);
nand I_18923 (I324395,I324313,I324378);
nand I_18924 (I323866,I324395,I324344);
nand I_18925 (I323863,I324378,I324262);
not I_18926 (I324467,I2690);
DFFARX1 I_18927 (I273662,I2683,I324467,I324493,);
and I_18928 (I324501,I324493,I273656);
DFFARX1 I_18929 (I324501,I2683,I324467,I324450,);
DFFARX1 I_18930 (I273674,I2683,I324467,I324541,);
not I_18931 (I324549,I273665);
not I_18932 (I324566,I273677);
nand I_18933 (I324583,I324566,I324549);
nor I_18934 (I324438,I324541,I324583);
DFFARX1 I_18935 (I324583,I2683,I324467,I324623,);
not I_18936 (I324459,I324623);
not I_18937 (I324645,I273683);
nand I_18938 (I324662,I324566,I324645);
DFFARX1 I_18939 (I324662,I2683,I324467,I324688,);
not I_18940 (I324696,I324688);
not I_18941 (I324713,I273659);
nand I_18942 (I324730,I324713,I273680);
and I_18943 (I324747,I324549,I324730);
nor I_18944 (I324764,I324662,I324747);
DFFARX1 I_18945 (I324764,I2683,I324467,I324435,);
DFFARX1 I_18946 (I324747,I2683,I324467,I324456,);
nor I_18947 (I324809,I273659,I273671);
nor I_18948 (I324447,I324662,I324809);
or I_18949 (I324840,I273659,I273671);
nor I_18950 (I324857,I273656,I273668);
DFFARX1 I_18951 (I324857,I2683,I324467,I324883,);
not I_18952 (I324891,I324883);
nor I_18953 (I324453,I324891,I324696);
nand I_18954 (I324922,I324891,I324541);
not I_18955 (I324939,I273656);
nand I_18956 (I324956,I324939,I324645);
nand I_18957 (I324973,I324891,I324956);
nand I_18958 (I324444,I324973,I324922);
nand I_18959 (I324441,I324956,I324840);
not I_18960 (I325045,I2690);
DFFARX1 I_18961 (I124814,I2683,I325045,I325071,);
and I_18962 (I325079,I325071,I124799);
DFFARX1 I_18963 (I325079,I2683,I325045,I325028,);
DFFARX1 I_18964 (I124805,I2683,I325045,I325119,);
not I_18965 (I325127,I124787);
not I_18966 (I325144,I124808);
nand I_18967 (I325161,I325144,I325127);
nor I_18968 (I325016,I325119,I325161);
DFFARX1 I_18969 (I325161,I2683,I325045,I325201,);
not I_18970 (I325037,I325201);
not I_18971 (I325223,I124811);
nand I_18972 (I325240,I325144,I325223);
DFFARX1 I_18973 (I325240,I2683,I325045,I325266,);
not I_18974 (I325274,I325266);
not I_18975 (I325291,I124802);
nand I_18976 (I325308,I325291,I124790);
and I_18977 (I325325,I325127,I325308);
nor I_18978 (I325342,I325240,I325325);
DFFARX1 I_18979 (I325342,I2683,I325045,I325013,);
DFFARX1 I_18980 (I325325,I2683,I325045,I325034,);
nor I_18981 (I325387,I124802,I124796);
nor I_18982 (I325025,I325240,I325387);
or I_18983 (I325418,I124802,I124796);
nor I_18984 (I325435,I124793,I124787);
DFFARX1 I_18985 (I325435,I2683,I325045,I325461,);
not I_18986 (I325469,I325461);
nor I_18987 (I325031,I325469,I325274);
nand I_18988 (I325500,I325469,I325119);
not I_18989 (I325517,I124793);
nand I_18990 (I325534,I325517,I325223);
nand I_18991 (I325551,I325469,I325534);
nand I_18992 (I325022,I325551,I325500);
nand I_18993 (I325019,I325534,I325418);
not I_18994 (I325623,I2690);
DFFARX1 I_18995 (I393438,I2683,I325623,I325649,);
and I_18996 (I325657,I325649,I393465);
DFFARX1 I_18997 (I325657,I2683,I325623,I325606,);
DFFARX1 I_18998 (I393447,I2683,I325623,I325697,);
not I_18999 (I325705,I393456);
not I_19000 (I325722,I393459);
nand I_19001 (I325739,I325722,I325705);
nor I_19002 (I325594,I325697,I325739);
DFFARX1 I_19003 (I325739,I2683,I325623,I325779,);
not I_19004 (I325615,I325779);
not I_19005 (I325801,I393453);
nand I_19006 (I325818,I325722,I325801);
DFFARX1 I_19007 (I325818,I2683,I325623,I325844,);
not I_19008 (I325852,I325844);
not I_19009 (I325869,I393441);
nand I_19010 (I325886,I325869,I393444);
and I_19011 (I325903,I325705,I325886);
nor I_19012 (I325920,I325818,I325903);
DFFARX1 I_19013 (I325920,I2683,I325623,I325591,);
DFFARX1 I_19014 (I325903,I2683,I325623,I325612,);
nor I_19015 (I325965,I393441,I393462);
nor I_19016 (I325603,I325818,I325965);
or I_19017 (I325996,I393441,I393462);
nor I_19018 (I326013,I393450,I393438);
DFFARX1 I_19019 (I326013,I2683,I325623,I326039,);
not I_19020 (I326047,I326039);
nor I_19021 (I325609,I326047,I325852);
nand I_19022 (I326078,I326047,I325697);
not I_19023 (I326095,I393450);
nand I_19024 (I326112,I326095,I325801);
nand I_19025 (I326129,I326047,I326112);
nand I_19026 (I325600,I326129,I326078);
nand I_19027 (I325597,I326112,I325996);
not I_19028 (I326201,I2690);
DFFARX1 I_19029 (I318250,I2683,I326201,I326227,);
and I_19030 (I326235,I326227,I318247);
DFFARX1 I_19031 (I326235,I2683,I326201,I326184,);
DFFARX1 I_19032 (I318253,I2683,I326201,I326275,);
not I_19033 (I326283,I318256);
not I_19034 (I326300,I318250);
nand I_19035 (I326317,I326300,I326283);
nor I_19036 (I326172,I326275,I326317);
DFFARX1 I_19037 (I326317,I2683,I326201,I326357,);
not I_19038 (I326193,I326357);
not I_19039 (I326379,I318265);
nand I_19040 (I326396,I326300,I326379);
DFFARX1 I_19041 (I326396,I2683,I326201,I326422,);
not I_19042 (I326430,I326422);
not I_19043 (I326447,I318262);
nand I_19044 (I326464,I326447,I318268);
and I_19045 (I326481,I326283,I326464);
nor I_19046 (I326498,I326396,I326481);
DFFARX1 I_19047 (I326498,I2683,I326201,I326169,);
DFFARX1 I_19048 (I326481,I2683,I326201,I326190,);
nor I_19049 (I326543,I318262,I318247);
nor I_19050 (I326181,I326396,I326543);
or I_19051 (I326574,I318262,I318247);
nor I_19052 (I326591,I318259,I318253);
DFFARX1 I_19053 (I326591,I2683,I326201,I326617,);
not I_19054 (I326625,I326617);
nor I_19055 (I326187,I326625,I326430);
nand I_19056 (I326656,I326625,I326275);
not I_19057 (I326673,I318259);
nand I_19058 (I326690,I326673,I326379);
nand I_19059 (I326707,I326625,I326690);
nand I_19060 (I326178,I326707,I326656);
nand I_19061 (I326175,I326690,I326574);
not I_19062 (I326779,I2690);
DFFARX1 I_19063 (I192666,I2683,I326779,I326805,);
and I_19064 (I326813,I326805,I192654);
DFFARX1 I_19065 (I326813,I2683,I326779,I326762,);
DFFARX1 I_19066 (I192669,I2683,I326779,I326853,);
not I_19067 (I326861,I192660);
not I_19068 (I326878,I192651);
nand I_19069 (I326895,I326878,I326861);
nor I_19070 (I326750,I326853,I326895);
DFFARX1 I_19071 (I326895,I2683,I326779,I326935,);
not I_19072 (I326771,I326935);
not I_19073 (I326957,I192657);
nand I_19074 (I326974,I326878,I326957);
DFFARX1 I_19075 (I326974,I2683,I326779,I327000,);
not I_19076 (I327008,I327000);
not I_19077 (I327025,I192672);
nand I_19078 (I327042,I327025,I192675);
and I_19079 (I327059,I326861,I327042);
nor I_19080 (I327076,I326974,I327059);
DFFARX1 I_19081 (I327076,I2683,I326779,I326747,);
DFFARX1 I_19082 (I327059,I2683,I326779,I326768,);
nor I_19083 (I327121,I192672,I192651);
nor I_19084 (I326759,I326974,I327121);
or I_19085 (I327152,I192672,I192651);
nor I_19086 (I327169,I192663,I192654);
DFFARX1 I_19087 (I327169,I2683,I326779,I327195,);
not I_19088 (I327203,I327195);
nor I_19089 (I326765,I327203,I327008);
nand I_19090 (I327234,I327203,I326853);
not I_19091 (I327251,I192663);
nand I_19092 (I327268,I327251,I326957);
nand I_19093 (I327285,I327203,I327268);
nand I_19094 (I326756,I327285,I327234);
nand I_19095 (I326753,I327268,I327152);
not I_19096 (I327357,I2690);
DFFARX1 I_19097 (I289812,I2683,I327357,I327383,);
and I_19098 (I327391,I327383,I289806);
DFFARX1 I_19099 (I327391,I2683,I327357,I327340,);
DFFARX1 I_19100 (I289824,I2683,I327357,I327431,);
not I_19101 (I327439,I289815);
not I_19102 (I327456,I289827);
nand I_19103 (I327473,I327456,I327439);
nor I_19104 (I327328,I327431,I327473);
DFFARX1 I_19105 (I327473,I2683,I327357,I327513,);
not I_19106 (I327349,I327513);
not I_19107 (I327535,I289833);
nand I_19108 (I327552,I327456,I327535);
DFFARX1 I_19109 (I327552,I2683,I327357,I327578,);
not I_19110 (I327586,I327578);
not I_19111 (I327603,I289809);
nand I_19112 (I327620,I327603,I289830);
and I_19113 (I327637,I327439,I327620);
nor I_19114 (I327654,I327552,I327637);
DFFARX1 I_19115 (I327654,I2683,I327357,I327325,);
DFFARX1 I_19116 (I327637,I2683,I327357,I327346,);
nor I_19117 (I327699,I289809,I289821);
nor I_19118 (I327337,I327552,I327699);
or I_19119 (I327730,I289809,I289821);
nor I_19120 (I327747,I289806,I289818);
DFFARX1 I_19121 (I327747,I2683,I327357,I327773,);
not I_19122 (I327781,I327773);
nor I_19123 (I327343,I327781,I327586);
nand I_19124 (I327812,I327781,I327431);
not I_19125 (I327829,I289806);
nand I_19126 (I327846,I327829,I327535);
nand I_19127 (I327863,I327781,I327846);
nand I_19128 (I327334,I327863,I327812);
nand I_19129 (I327331,I327846,I327730);
not I_19130 (I327935,I2690);
DFFARX1 I_19131 (I261351,I2683,I327935,I327961,);
and I_19132 (I327969,I327961,I261357);
DFFARX1 I_19133 (I327969,I2683,I327935,I327918,);
DFFARX1 I_19134 (I261363,I2683,I327935,I328009,);
not I_19135 (I328017,I261348);
not I_19136 (I328034,I261348);
nand I_19137 (I328051,I328034,I328017);
nor I_19138 (I327906,I328009,I328051);
DFFARX1 I_19139 (I328051,I2683,I327935,I328091,);
not I_19140 (I327927,I328091);
not I_19141 (I328113,I261366);
nand I_19142 (I328130,I328034,I328113);
DFFARX1 I_19143 (I328130,I2683,I327935,I328156,);
not I_19144 (I328164,I328156);
not I_19145 (I328181,I261360);
nand I_19146 (I328198,I328181,I261351);
and I_19147 (I328215,I328017,I328198);
nor I_19148 (I328232,I328130,I328215);
DFFARX1 I_19149 (I328232,I2683,I327935,I327903,);
DFFARX1 I_19150 (I328215,I2683,I327935,I327924,);
nor I_19151 (I328277,I261360,I261369);
nor I_19152 (I327915,I328130,I328277);
or I_19153 (I328308,I261360,I261369);
nor I_19154 (I328325,I261354,I261354);
DFFARX1 I_19155 (I328325,I2683,I327935,I328351,);
not I_19156 (I328359,I328351);
nor I_19157 (I327921,I328359,I328164);
nand I_19158 (I328390,I328359,I328009);
not I_19159 (I328407,I261354);
nand I_19160 (I328424,I328407,I328113);
nand I_19161 (I328441,I328359,I328424);
nand I_19162 (I327912,I328441,I328390);
nand I_19163 (I327909,I328424,I328308);
not I_19164 (I328513,I2690);
DFFARX1 I_19165 (I30461,I2683,I328513,I328539,);
and I_19166 (I328547,I328539,I30437);
DFFARX1 I_19167 (I328547,I2683,I328513,I328496,);
DFFARX1 I_19168 (I30455,I2683,I328513,I328587,);
not I_19169 (I328595,I30443);
not I_19170 (I328612,I30440);
nand I_19171 (I328629,I328612,I328595);
nor I_19172 (I328484,I328587,I328629);
DFFARX1 I_19173 (I328629,I2683,I328513,I328669,);
not I_19174 (I328505,I328669);
not I_19175 (I328691,I30449);
nand I_19176 (I328708,I328612,I328691);
DFFARX1 I_19177 (I328708,I2683,I328513,I328734,);
not I_19178 (I328742,I328734);
not I_19179 (I328759,I30440);
nand I_19180 (I328776,I328759,I30458);
and I_19181 (I328793,I328595,I328776);
nor I_19182 (I328810,I328708,I328793);
DFFARX1 I_19183 (I328810,I2683,I328513,I328481,);
DFFARX1 I_19184 (I328793,I2683,I328513,I328502,);
nor I_19185 (I328855,I30440,I30452);
nor I_19186 (I328493,I328708,I328855);
or I_19187 (I328886,I30440,I30452);
nor I_19188 (I328903,I30446,I30437);
DFFARX1 I_19189 (I328903,I2683,I328513,I328929,);
not I_19190 (I328937,I328929);
nor I_19191 (I328499,I328937,I328742);
nand I_19192 (I328968,I328937,I328587);
not I_19193 (I328985,I30446);
nand I_19194 (I329002,I328985,I328691);
nand I_19195 (I329019,I328937,I329002);
nand I_19196 (I328490,I329019,I328968);
nand I_19197 (I328487,I329002,I328886);
not I_19198 (I329091,I2690);
DFFARX1 I_19199 (I92140,I2683,I329091,I329117,);
and I_19200 (I329125,I329117,I92125);
DFFARX1 I_19201 (I329125,I2683,I329091,I329074,);
DFFARX1 I_19202 (I92131,I2683,I329091,I329165,);
not I_19203 (I329173,I92113);
not I_19204 (I329190,I92134);
nand I_19205 (I329207,I329190,I329173);
nor I_19206 (I329062,I329165,I329207);
DFFARX1 I_19207 (I329207,I2683,I329091,I329247,);
not I_19208 (I329083,I329247);
not I_19209 (I329269,I92137);
nand I_19210 (I329286,I329190,I329269);
DFFARX1 I_19211 (I329286,I2683,I329091,I329312,);
not I_19212 (I329320,I329312);
not I_19213 (I329337,I92128);
nand I_19214 (I329354,I329337,I92116);
and I_19215 (I329371,I329173,I329354);
nor I_19216 (I329388,I329286,I329371);
DFFARX1 I_19217 (I329388,I2683,I329091,I329059,);
DFFARX1 I_19218 (I329371,I2683,I329091,I329080,);
nor I_19219 (I329433,I92128,I92122);
nor I_19220 (I329071,I329286,I329433);
or I_19221 (I329464,I92128,I92122);
nor I_19222 (I329481,I92119,I92113);
DFFARX1 I_19223 (I329481,I2683,I329091,I329507,);
not I_19224 (I329515,I329507);
nor I_19225 (I329077,I329515,I329320);
nand I_19226 (I329546,I329515,I329165);
not I_19227 (I329563,I92119);
nand I_19228 (I329580,I329563,I329269);
nand I_19229 (I329597,I329515,I329580);
nand I_19230 (I329068,I329597,I329546);
nand I_19231 (I329065,I329580,I329464);
not I_19232 (I329669,I2690);
DFFARX1 I_19233 (I390589,I2683,I329669,I329695,);
and I_19234 (I329703,I329695,I390571);
DFFARX1 I_19235 (I329703,I2683,I329669,I329652,);
DFFARX1 I_19236 (I390580,I2683,I329669,I329743,);
not I_19237 (I329751,I390565);
not I_19238 (I329768,I390577);
nand I_19239 (I329785,I329768,I329751);
nor I_19240 (I329640,I329743,I329785);
DFFARX1 I_19241 (I329785,I2683,I329669,I329825,);
not I_19242 (I329661,I329825);
not I_19243 (I329847,I390568);
nand I_19244 (I329864,I329768,I329847);
DFFARX1 I_19245 (I329864,I2683,I329669,I329890,);
not I_19246 (I329898,I329890);
not I_19247 (I329915,I390565);
nand I_19248 (I329932,I329915,I390568);
and I_19249 (I329949,I329751,I329932);
nor I_19250 (I329966,I329864,I329949);
DFFARX1 I_19251 (I329966,I2683,I329669,I329637,);
DFFARX1 I_19252 (I329949,I2683,I329669,I329658,);
nor I_19253 (I330011,I390565,I390586);
nor I_19254 (I329649,I329864,I330011);
or I_19255 (I330042,I390565,I390586);
nor I_19256 (I330059,I390574,I390583);
DFFARX1 I_19257 (I330059,I2683,I329669,I330085,);
not I_19258 (I330093,I330085);
nor I_19259 (I329655,I330093,I329898);
nand I_19260 (I330124,I330093,I329743);
not I_19261 (I330141,I390574);
nand I_19262 (I330158,I330141,I329847);
nand I_19263 (I330175,I330093,I330158);
nand I_19264 (I329646,I330175,I330124);
nand I_19265 (I329643,I330158,I330042);
not I_19266 (I330247,I2690);
DFFARX1 I_19267 (I172436,I2683,I330247,I330273,);
and I_19268 (I330281,I330273,I172424);
DFFARX1 I_19269 (I330281,I2683,I330247,I330230,);
DFFARX1 I_19270 (I172439,I2683,I330247,I330321,);
not I_19271 (I330329,I172430);
not I_19272 (I330346,I172421);
nand I_19273 (I330363,I330346,I330329);
nor I_19274 (I330218,I330321,I330363);
DFFARX1 I_19275 (I330363,I2683,I330247,I330403,);
not I_19276 (I330239,I330403);
not I_19277 (I330425,I172427);
nand I_19278 (I330442,I330346,I330425);
DFFARX1 I_19279 (I330442,I2683,I330247,I330468,);
not I_19280 (I330476,I330468);
not I_19281 (I330493,I172442);
nand I_19282 (I330510,I330493,I172445);
and I_19283 (I330527,I330329,I330510);
nor I_19284 (I330544,I330442,I330527);
DFFARX1 I_19285 (I330544,I2683,I330247,I330215,);
DFFARX1 I_19286 (I330527,I2683,I330247,I330236,);
nor I_19287 (I330589,I172442,I172421);
nor I_19288 (I330227,I330442,I330589);
or I_19289 (I330620,I172442,I172421);
nor I_19290 (I330637,I172433,I172424);
DFFARX1 I_19291 (I330637,I2683,I330247,I330663,);
not I_19292 (I330671,I330663);
nor I_19293 (I330233,I330671,I330476);
nand I_19294 (I330702,I330671,I330321);
not I_19295 (I330719,I172433);
nand I_19296 (I330736,I330719,I330425);
nand I_19297 (I330753,I330671,I330736);
nand I_19298 (I330224,I330753,I330702);
nand I_19299 (I330221,I330736,I330620);
not I_19300 (I330825,I2690);
DFFARX1 I_19301 (I131791,I2683,I330825,I330851,);
and I_19302 (I330859,I330851,I131806);
DFFARX1 I_19303 (I330859,I2683,I330825,I330808,);
DFFARX1 I_19304 (I131809,I2683,I330825,I330899,);
not I_19305 (I330907,I131803);
not I_19306 (I330924,I131818);
nand I_19307 (I330941,I330924,I330907);
nor I_19308 (I330796,I330899,I330941);
DFFARX1 I_19309 (I330941,I2683,I330825,I330981,);
not I_19310 (I330817,I330981);
not I_19311 (I331003,I131794);
nand I_19312 (I331020,I330924,I331003);
DFFARX1 I_19313 (I331020,I2683,I330825,I331046,);
not I_19314 (I331054,I331046);
not I_19315 (I331071,I131797);
nand I_19316 (I331088,I331071,I131791);
and I_19317 (I331105,I330907,I331088);
nor I_19318 (I331122,I331020,I331105);
DFFARX1 I_19319 (I331122,I2683,I330825,I330793,);
DFFARX1 I_19320 (I331105,I2683,I330825,I330814,);
nor I_19321 (I331167,I131797,I131800);
nor I_19322 (I330805,I331020,I331167);
or I_19323 (I331198,I131797,I131800);
nor I_19324 (I331215,I131815,I131812);
DFFARX1 I_19325 (I331215,I2683,I330825,I331241,);
not I_19326 (I331249,I331241);
nor I_19327 (I330811,I331249,I331054);
nand I_19328 (I331280,I331249,I330899);
not I_19329 (I331297,I131815);
nand I_19330 (I331314,I331297,I331003);
nand I_19331 (I331331,I331249,I331314);
nand I_19332 (I330802,I331331,I331280);
nand I_19333 (I330799,I331314,I331198);
not I_19334 (I331403,I2690);
DFFARX1 I_19335 (I14100,I2683,I331403,I331429,);
and I_19336 (I331437,I331429,I14103);
DFFARX1 I_19337 (I331437,I2683,I331403,I331386,);
DFFARX1 I_19338 (I14103,I2683,I331403,I331477,);
not I_19339 (I331485,I14106);
not I_19340 (I331502,I14121);
nand I_19341 (I331519,I331502,I331485);
nor I_19342 (I331374,I331477,I331519);
DFFARX1 I_19343 (I331519,I2683,I331403,I331559,);
not I_19344 (I331395,I331559);
not I_19345 (I331581,I14115);
nand I_19346 (I331598,I331502,I331581);
DFFARX1 I_19347 (I331598,I2683,I331403,I331624,);
not I_19348 (I331632,I331624);
not I_19349 (I331649,I14118);
nand I_19350 (I331666,I331649,I14100);
and I_19351 (I331683,I331485,I331666);
nor I_19352 (I331700,I331598,I331683);
DFFARX1 I_19353 (I331700,I2683,I331403,I331371,);
DFFARX1 I_19354 (I331683,I2683,I331403,I331392,);
nor I_19355 (I331745,I14118,I14112);
nor I_19356 (I331383,I331598,I331745);
or I_19357 (I331776,I14118,I14112);
nor I_19358 (I331793,I14109,I14124);
DFFARX1 I_19359 (I331793,I2683,I331403,I331819,);
not I_19360 (I331827,I331819);
nor I_19361 (I331389,I331827,I331632);
nand I_19362 (I331858,I331827,I331477);
not I_19363 (I331875,I14109);
nand I_19364 (I331892,I331875,I331581);
nand I_19365 (I331909,I331827,I331892);
nand I_19366 (I331380,I331909,I331858);
nand I_19367 (I331377,I331892,I331776);
not I_19368 (I331981,I2690);
DFFARX1 I_19369 (I153007,I2683,I331981,I332007,);
and I_19370 (I332015,I332007,I153022);
DFFARX1 I_19371 (I332015,I2683,I331981,I331964,);
DFFARX1 I_19372 (I153025,I2683,I331981,I332055,);
not I_19373 (I332063,I153019);
not I_19374 (I332080,I153034);
nand I_19375 (I332097,I332080,I332063);
nor I_19376 (I331952,I332055,I332097);
DFFARX1 I_19377 (I332097,I2683,I331981,I332137,);
not I_19378 (I331973,I332137);
not I_19379 (I332159,I153010);
nand I_19380 (I332176,I332080,I332159);
DFFARX1 I_19381 (I332176,I2683,I331981,I332202,);
not I_19382 (I332210,I332202);
not I_19383 (I332227,I153013);
nand I_19384 (I332244,I332227,I153007);
and I_19385 (I332261,I332063,I332244);
nor I_19386 (I332278,I332176,I332261);
DFFARX1 I_19387 (I332278,I2683,I331981,I331949,);
DFFARX1 I_19388 (I332261,I2683,I331981,I331970,);
nor I_19389 (I332323,I153013,I153016);
nor I_19390 (I331961,I332176,I332323);
or I_19391 (I332354,I153013,I153016);
nor I_19392 (I332371,I153031,I153028);
DFFARX1 I_19393 (I332371,I2683,I331981,I332397,);
not I_19394 (I332405,I332397);
nor I_19395 (I331967,I332405,I332210);
nand I_19396 (I332436,I332405,I332055);
not I_19397 (I332453,I153031);
nand I_19398 (I332470,I332453,I332159);
nand I_19399 (I332487,I332405,I332470);
nand I_19400 (I331958,I332487,I332436);
nand I_19401 (I331955,I332470,I332354);
not I_19402 (I332559,I2690);
DFFARX1 I_19403 (I322177,I2683,I332559,I332585,);
and I_19404 (I332593,I332585,I322174);
DFFARX1 I_19405 (I332593,I2683,I332559,I332542,);
DFFARX1 I_19406 (I322180,I2683,I332559,I332633,);
not I_19407 (I332641,I322183);
not I_19408 (I332658,I322177);
nand I_19409 (I332675,I332658,I332641);
nor I_19410 (I332530,I332633,I332675);
DFFARX1 I_19411 (I332675,I2683,I332559,I332715,);
not I_19412 (I332551,I332715);
not I_19413 (I332737,I322192);
nand I_19414 (I332754,I332658,I332737);
DFFARX1 I_19415 (I332754,I2683,I332559,I332780,);
not I_19416 (I332788,I332780);
not I_19417 (I332805,I322189);
nand I_19418 (I332822,I332805,I322195);
and I_19419 (I332839,I332641,I332822);
nor I_19420 (I332856,I332754,I332839);
DFFARX1 I_19421 (I332856,I2683,I332559,I332527,);
DFFARX1 I_19422 (I332839,I2683,I332559,I332548,);
nor I_19423 (I332901,I322189,I322174);
nor I_19424 (I332539,I332754,I332901);
or I_19425 (I332932,I322189,I322174);
nor I_19426 (I332949,I322186,I322180);
DFFARX1 I_19427 (I332949,I2683,I332559,I332975,);
not I_19428 (I332983,I332975);
nor I_19429 (I332545,I332983,I332788);
nand I_19430 (I333014,I332983,I332633);
not I_19431 (I333031,I322186);
nand I_19432 (I333048,I333031,I332737);
nand I_19433 (I333065,I332983,I333048);
nand I_19434 (I332536,I333065,I333014);
nand I_19435 (I332533,I333048,I332932);
not I_19436 (I333137,I2690);
DFFARX1 I_19437 (I301440,I2683,I333137,I333163,);
and I_19438 (I333171,I333163,I301434);
DFFARX1 I_19439 (I333171,I2683,I333137,I333120,);
DFFARX1 I_19440 (I301452,I2683,I333137,I333211,);
not I_19441 (I333219,I301443);
not I_19442 (I333236,I301455);
nand I_19443 (I333253,I333236,I333219);
nor I_19444 (I333108,I333211,I333253);
DFFARX1 I_19445 (I333253,I2683,I333137,I333293,);
not I_19446 (I333129,I333293);
not I_19447 (I333315,I301461);
nand I_19448 (I333332,I333236,I333315);
DFFARX1 I_19449 (I333332,I2683,I333137,I333358,);
not I_19450 (I333366,I333358);
not I_19451 (I333383,I301437);
nand I_19452 (I333400,I333383,I301458);
and I_19453 (I333417,I333219,I333400);
nor I_19454 (I333434,I333332,I333417);
DFFARX1 I_19455 (I333434,I2683,I333137,I333105,);
DFFARX1 I_19456 (I333417,I2683,I333137,I333126,);
nor I_19457 (I333479,I301437,I301449);
nor I_19458 (I333117,I333332,I333479);
or I_19459 (I333510,I301437,I301449);
nor I_19460 (I333527,I301434,I301446);
DFFARX1 I_19461 (I333527,I2683,I333137,I333553,);
not I_19462 (I333561,I333553);
nor I_19463 (I333123,I333561,I333366);
nand I_19464 (I333592,I333561,I333211);
not I_19465 (I333609,I301434);
nand I_19466 (I333626,I333609,I333315);
nand I_19467 (I333643,I333561,I333626);
nand I_19468 (I333114,I333643,I333592);
nand I_19469 (I333111,I333626,I333510);
not I_19470 (I333715,I2690);
DFFARX1 I_19471 (I182840,I2683,I333715,I333741,);
and I_19472 (I333749,I333741,I182828);
DFFARX1 I_19473 (I333749,I2683,I333715,I333698,);
DFFARX1 I_19474 (I182843,I2683,I333715,I333789,);
not I_19475 (I333797,I182834);
not I_19476 (I333814,I182825);
nand I_19477 (I333831,I333814,I333797);
nor I_19478 (I333686,I333789,I333831);
DFFARX1 I_19479 (I333831,I2683,I333715,I333871,);
not I_19480 (I333707,I333871);
not I_19481 (I333893,I182831);
nand I_19482 (I333910,I333814,I333893);
DFFARX1 I_19483 (I333910,I2683,I333715,I333936,);
not I_19484 (I333944,I333936);
not I_19485 (I333961,I182846);
nand I_19486 (I333978,I333961,I182849);
and I_19487 (I333995,I333797,I333978);
nor I_19488 (I334012,I333910,I333995);
DFFARX1 I_19489 (I334012,I2683,I333715,I333683,);
DFFARX1 I_19490 (I333995,I2683,I333715,I333704,);
nor I_19491 (I334057,I182846,I182825);
nor I_19492 (I333695,I333910,I334057);
or I_19493 (I334088,I182846,I182825);
nor I_19494 (I334105,I182837,I182828);
DFFARX1 I_19495 (I334105,I2683,I333715,I334131,);
not I_19496 (I334139,I334131);
nor I_19497 (I333701,I334139,I333944);
nand I_19498 (I334170,I334139,I333789);
not I_19499 (I334187,I182837);
nand I_19500 (I334204,I334187,I333893);
nand I_19501 (I334221,I334139,I334204);
nand I_19502 (I333692,I334221,I334170);
nand I_19503 (I333689,I334204,I334088);
not I_19504 (I334293,I2690);
DFFARX1 I_19505 (I120598,I2683,I334293,I334319,);
and I_19506 (I334327,I334319,I120583);
DFFARX1 I_19507 (I334327,I2683,I334293,I334276,);
DFFARX1 I_19508 (I120589,I2683,I334293,I334367,);
not I_19509 (I334375,I120571);
not I_19510 (I334392,I120592);
nand I_19511 (I334409,I334392,I334375);
nor I_19512 (I334264,I334367,I334409);
DFFARX1 I_19513 (I334409,I2683,I334293,I334449,);
not I_19514 (I334285,I334449);
not I_19515 (I334471,I120595);
nand I_19516 (I334488,I334392,I334471);
DFFARX1 I_19517 (I334488,I2683,I334293,I334514,);
not I_19518 (I334522,I334514);
not I_19519 (I334539,I120586);
nand I_19520 (I334556,I334539,I120574);
and I_19521 (I334573,I334375,I334556);
nor I_19522 (I334590,I334488,I334573);
DFFARX1 I_19523 (I334590,I2683,I334293,I334261,);
DFFARX1 I_19524 (I334573,I2683,I334293,I334282,);
nor I_19525 (I334635,I120586,I120580);
nor I_19526 (I334273,I334488,I334635);
or I_19527 (I334666,I120586,I120580);
nor I_19528 (I334683,I120577,I120571);
DFFARX1 I_19529 (I334683,I2683,I334293,I334709,);
not I_19530 (I334717,I334709);
nor I_19531 (I334279,I334717,I334522);
nand I_19532 (I334748,I334717,I334367);
not I_19533 (I334765,I120577);
nand I_19534 (I334782,I334765,I334471);
nand I_19535 (I334799,I334717,I334782);
nand I_19536 (I334270,I334799,I334748);
nand I_19537 (I334267,I334782,I334666);
not I_19538 (I334871,I2690);
DFFARX1 I_19539 (I257662,I2683,I334871,I334897,);
and I_19540 (I334905,I334897,I257668);
DFFARX1 I_19541 (I334905,I2683,I334871,I334854,);
DFFARX1 I_19542 (I257674,I2683,I334871,I334945,);
not I_19543 (I334953,I257659);
not I_19544 (I334970,I257659);
nand I_19545 (I334987,I334970,I334953);
nor I_19546 (I334842,I334945,I334987);
DFFARX1 I_19547 (I334987,I2683,I334871,I335027,);
not I_19548 (I334863,I335027);
not I_19549 (I335049,I257677);
nand I_19550 (I335066,I334970,I335049);
DFFARX1 I_19551 (I335066,I2683,I334871,I335092,);
not I_19552 (I335100,I335092);
not I_19553 (I335117,I257671);
nand I_19554 (I335134,I335117,I257662);
and I_19555 (I335151,I334953,I335134);
nor I_19556 (I335168,I335066,I335151);
DFFARX1 I_19557 (I335168,I2683,I334871,I334839,);
DFFARX1 I_19558 (I335151,I2683,I334871,I334860,);
nor I_19559 (I335213,I257671,I257680);
nor I_19560 (I334851,I335066,I335213);
or I_19561 (I335244,I257671,I257680);
nor I_19562 (I335261,I257665,I257665);
DFFARX1 I_19563 (I335261,I2683,I334871,I335287,);
not I_19564 (I335295,I335287);
nor I_19565 (I334857,I335295,I335100);
nand I_19566 (I335326,I335295,I334945);
not I_19567 (I335343,I257665);
nand I_19568 (I335360,I335343,I335049);
nand I_19569 (I335377,I335295,I335360);
nand I_19570 (I334848,I335377,I335326);
nand I_19571 (I334845,I335360,I335244);
not I_19572 (I335449,I2690);
DFFARX1 I_19573 (I238163,I2683,I335449,I335475,);
and I_19574 (I335483,I335475,I238169);
DFFARX1 I_19575 (I335483,I2683,I335449,I335432,);
DFFARX1 I_19576 (I238175,I2683,I335449,I335523,);
not I_19577 (I335531,I238160);
not I_19578 (I335548,I238160);
nand I_19579 (I335565,I335548,I335531);
nor I_19580 (I335420,I335523,I335565);
DFFARX1 I_19581 (I335565,I2683,I335449,I335605,);
not I_19582 (I335441,I335605);
not I_19583 (I335627,I238178);
nand I_19584 (I335644,I335548,I335627);
DFFARX1 I_19585 (I335644,I2683,I335449,I335670,);
not I_19586 (I335678,I335670);
not I_19587 (I335695,I238172);
nand I_19588 (I335712,I335695,I238163);
and I_19589 (I335729,I335531,I335712);
nor I_19590 (I335746,I335644,I335729);
DFFARX1 I_19591 (I335746,I2683,I335449,I335417,);
DFFARX1 I_19592 (I335729,I2683,I335449,I335438,);
nor I_19593 (I335791,I238172,I238181);
nor I_19594 (I335429,I335644,I335791);
or I_19595 (I335822,I238172,I238181);
nor I_19596 (I335839,I238166,I238166);
DFFARX1 I_19597 (I335839,I2683,I335449,I335865,);
not I_19598 (I335873,I335865);
nor I_19599 (I335435,I335873,I335678);
nand I_19600 (I335904,I335873,I335523);
not I_19601 (I335921,I238166);
nand I_19602 (I335938,I335921,I335627);
nand I_19603 (I335955,I335873,I335938);
nand I_19604 (I335426,I335955,I335904);
nand I_19605 (I335423,I335938,I335822);
not I_19606 (I336027,I2690);
DFFARX1 I_19607 (I394560,I2683,I336027,I336053,);
and I_19608 (I336061,I336053,I394587);
DFFARX1 I_19609 (I336061,I2683,I336027,I336010,);
DFFARX1 I_19610 (I394569,I2683,I336027,I336101,);
not I_19611 (I336109,I394578);
not I_19612 (I336126,I394581);
nand I_19613 (I336143,I336126,I336109);
nor I_19614 (I335998,I336101,I336143);
DFFARX1 I_19615 (I336143,I2683,I336027,I336183,);
not I_19616 (I336019,I336183);
not I_19617 (I336205,I394575);
nand I_19618 (I336222,I336126,I336205);
DFFARX1 I_19619 (I336222,I2683,I336027,I336248,);
not I_19620 (I336256,I336248);
not I_19621 (I336273,I394563);
nand I_19622 (I336290,I336273,I394566);
and I_19623 (I336307,I336109,I336290);
nor I_19624 (I336324,I336222,I336307);
DFFARX1 I_19625 (I336324,I2683,I336027,I335995,);
DFFARX1 I_19626 (I336307,I2683,I336027,I336016,);
nor I_19627 (I336369,I394563,I394584);
nor I_19628 (I336007,I336222,I336369);
or I_19629 (I336400,I394563,I394584);
nor I_19630 (I336417,I394572,I394560);
DFFARX1 I_19631 (I336417,I2683,I336027,I336443,);
not I_19632 (I336451,I336443);
nor I_19633 (I336013,I336451,I336256);
nand I_19634 (I336482,I336451,I336101);
not I_19635 (I336499,I394572);
nand I_19636 (I336516,I336499,I336205);
nand I_19637 (I336533,I336451,I336516);
nand I_19638 (I336004,I336533,I336482);
nand I_19639 (I336001,I336516,I336400);
not I_19640 (I336605,I2690);
DFFARX1 I_19641 (I91086,I2683,I336605,I336631,);
and I_19642 (I336639,I336631,I91071);
DFFARX1 I_19643 (I336639,I2683,I336605,I336588,);
DFFARX1 I_19644 (I91077,I2683,I336605,I336679,);
not I_19645 (I336687,I91059);
not I_19646 (I336704,I91080);
nand I_19647 (I336721,I336704,I336687);
nor I_19648 (I336576,I336679,I336721);
DFFARX1 I_19649 (I336721,I2683,I336605,I336761,);
not I_19650 (I336597,I336761);
not I_19651 (I336783,I91083);
nand I_19652 (I336800,I336704,I336783);
DFFARX1 I_19653 (I336800,I2683,I336605,I336826,);
not I_19654 (I336834,I336826);
not I_19655 (I336851,I91074);
nand I_19656 (I336868,I336851,I91062);
and I_19657 (I336885,I336687,I336868);
nor I_19658 (I336902,I336800,I336885);
DFFARX1 I_19659 (I336902,I2683,I336605,I336573,);
DFFARX1 I_19660 (I336885,I2683,I336605,I336594,);
nor I_19661 (I336947,I91074,I91068);
nor I_19662 (I336585,I336800,I336947);
or I_19663 (I336978,I91074,I91068);
nor I_19664 (I336995,I91065,I91059);
DFFARX1 I_19665 (I336995,I2683,I336605,I337021,);
not I_19666 (I337029,I337021);
nor I_19667 (I336591,I337029,I336834);
nand I_19668 (I337060,I337029,I336679);
not I_19669 (I337077,I91065);
nand I_19670 (I337094,I337077,I336783);
nand I_19671 (I337111,I337029,I337094);
nand I_19672 (I336582,I337111,I337060);
nand I_19673 (I336579,I337094,I336978);
not I_19674 (I337183,I2690);
DFFARX1 I_19675 (I231970,I2683,I337183,I337209,);
and I_19676 (I337217,I337209,I231958);
DFFARX1 I_19677 (I337217,I2683,I337183,I337166,);
DFFARX1 I_19678 (I231961,I2683,I337183,I337257,);
not I_19679 (I337265,I231955);
not I_19680 (I337282,I231979);
nand I_19681 (I337299,I337282,I337265);
nor I_19682 (I337154,I337257,I337299);
DFFARX1 I_19683 (I337299,I2683,I337183,I337339,);
not I_19684 (I337175,I337339);
not I_19685 (I337361,I231967);
nand I_19686 (I337378,I337282,I337361);
DFFARX1 I_19687 (I337378,I2683,I337183,I337404,);
not I_19688 (I337412,I337404);
not I_19689 (I337429,I231976);
nand I_19690 (I337446,I337429,I231973);
and I_19691 (I337463,I337265,I337446);
nor I_19692 (I337480,I337378,I337463);
DFFARX1 I_19693 (I337480,I2683,I337183,I337151,);
DFFARX1 I_19694 (I337463,I2683,I337183,I337172,);
nor I_19695 (I337525,I231976,I231964);
nor I_19696 (I337163,I337378,I337525);
or I_19697 (I337556,I231976,I231964);
nor I_19698 (I337573,I231955,I231958);
DFFARX1 I_19699 (I337573,I2683,I337183,I337599,);
not I_19700 (I337607,I337599);
nor I_19701 (I337169,I337607,I337412);
nand I_19702 (I337638,I337607,I337257);
not I_19703 (I337655,I231955);
nand I_19704 (I337672,I337655,I337361);
nand I_19705 (I337689,I337607,I337672);
nand I_19706 (I337160,I337689,I337638);
nand I_19707 (I337157,I337672,I337556);
not I_19708 (I337761,I2690);
DFFARX1 I_19709 (I387121,I2683,I337761,I337787,);
and I_19710 (I337795,I337787,I387103);
DFFARX1 I_19711 (I337795,I2683,I337761,I337744,);
DFFARX1 I_19712 (I387112,I2683,I337761,I337835,);
not I_19713 (I337843,I387097);
not I_19714 (I337860,I387109);
nand I_19715 (I337877,I337860,I337843);
nor I_19716 (I337732,I337835,I337877);
DFFARX1 I_19717 (I337877,I2683,I337761,I337917,);
not I_19718 (I337753,I337917);
not I_19719 (I337939,I387100);
nand I_19720 (I337956,I337860,I337939);
DFFARX1 I_19721 (I337956,I2683,I337761,I337982,);
not I_19722 (I337990,I337982);
not I_19723 (I338007,I387097);
nand I_19724 (I338024,I338007,I387100);
and I_19725 (I338041,I337843,I338024);
nor I_19726 (I338058,I337956,I338041);
DFFARX1 I_19727 (I338058,I2683,I337761,I337729,);
DFFARX1 I_19728 (I338041,I2683,I337761,I337750,);
nor I_19729 (I338103,I387097,I387118);
nor I_19730 (I337741,I337956,I338103);
or I_19731 (I338134,I387097,I387118);
nor I_19732 (I338151,I387106,I387115);
DFFARX1 I_19733 (I338151,I2683,I337761,I338177,);
not I_19734 (I338185,I338177);
nor I_19735 (I337747,I338185,I337990);
nand I_19736 (I338216,I338185,I337835);
not I_19737 (I338233,I387106);
nand I_19738 (I338250,I338233,I337939);
nand I_19739 (I338267,I338185,I338250);
nand I_19740 (I337738,I338267,I338216);
nand I_19741 (I337735,I338250,I338134);
not I_19742 (I338339,I2690);
DFFARX1 I_19743 (I2540,I2683,I338339,I338365,);
and I_19744 (I338373,I338365,I1900);
DFFARX1 I_19745 (I338373,I2683,I338339,I338322,);
DFFARX1 I_19746 (I1756,I2683,I338339,I338413,);
not I_19747 (I338421,I2300);
not I_19748 (I338438,I2644);
nand I_19749 (I338455,I338438,I338421);
nor I_19750 (I338310,I338413,I338455);
DFFARX1 I_19751 (I338455,I2683,I338339,I338495,);
not I_19752 (I338331,I338495);
not I_19753 (I338517,I1684);
nand I_19754 (I338534,I338438,I338517);
DFFARX1 I_19755 (I338534,I2683,I338339,I338560,);
not I_19756 (I338568,I338560);
not I_19757 (I338585,I1700);
nand I_19758 (I338602,I338585,I1476);
and I_19759 (I338619,I338421,I338602);
nor I_19760 (I338636,I338534,I338619);
DFFARX1 I_19761 (I338636,I2683,I338339,I338307,);
DFFARX1 I_19762 (I338619,I2683,I338339,I338328,);
nor I_19763 (I338681,I1700,I2420);
nor I_19764 (I338319,I338534,I338681);
or I_19765 (I338712,I1700,I2420);
nor I_19766 (I338729,I2060,I1804);
DFFARX1 I_19767 (I338729,I2683,I338339,I338755,);
not I_19768 (I338763,I338755);
nor I_19769 (I338325,I338763,I338568);
nand I_19770 (I338794,I338763,I338413);
not I_19771 (I338811,I2060);
nand I_19772 (I338828,I338811,I338517);
nand I_19773 (I338845,I338763,I338828);
nand I_19774 (I338316,I338845,I338794);
nand I_19775 (I338313,I338828,I338712);
not I_19776 (I338917,I2690);
DFFARX1 I_19777 (I106369,I2683,I338917,I338943,);
and I_19778 (I338951,I338943,I106354);
DFFARX1 I_19779 (I338951,I2683,I338917,I338900,);
DFFARX1 I_19780 (I106360,I2683,I338917,I338991,);
not I_19781 (I338999,I106342);
not I_19782 (I339016,I106363);
nand I_19783 (I339033,I339016,I338999);
nor I_19784 (I338888,I338991,I339033);
DFFARX1 I_19785 (I339033,I2683,I338917,I339073,);
not I_19786 (I338909,I339073);
not I_19787 (I339095,I106366);
nand I_19788 (I339112,I339016,I339095);
DFFARX1 I_19789 (I339112,I2683,I338917,I339138,);
not I_19790 (I339146,I339138);
not I_19791 (I339163,I106357);
nand I_19792 (I339180,I339163,I106345);
and I_19793 (I339197,I338999,I339180);
nor I_19794 (I339214,I339112,I339197);
DFFARX1 I_19795 (I339214,I2683,I338917,I338885,);
DFFARX1 I_19796 (I339197,I2683,I338917,I338906,);
nor I_19797 (I339259,I106357,I106351);
nor I_19798 (I338897,I339112,I339259);
or I_19799 (I339290,I106357,I106351);
nor I_19800 (I339307,I106348,I106342);
DFFARX1 I_19801 (I339307,I2683,I338917,I339333,);
not I_19802 (I339341,I339333);
nor I_19803 (I338903,I339341,I339146);
nand I_19804 (I339372,I339341,I338991);
not I_19805 (I339389,I106348);
nand I_19806 (I339406,I339389,I339095);
nand I_19807 (I339423,I339341,I339406);
nand I_19808 (I338894,I339423,I339372);
nand I_19809 (I338891,I339406,I339290);
not I_19810 (I339495,I2690);
DFFARX1 I_19811 (I128527,I2683,I339495,I339521,);
and I_19812 (I339529,I339521,I128542);
DFFARX1 I_19813 (I339529,I2683,I339495,I339478,);
DFFARX1 I_19814 (I128545,I2683,I339495,I339569,);
not I_19815 (I339577,I128539);
not I_19816 (I339594,I128554);
nand I_19817 (I339611,I339594,I339577);
nor I_19818 (I339466,I339569,I339611);
DFFARX1 I_19819 (I339611,I2683,I339495,I339651,);
not I_19820 (I339487,I339651);
not I_19821 (I339673,I128530);
nand I_19822 (I339690,I339594,I339673);
DFFARX1 I_19823 (I339690,I2683,I339495,I339716,);
not I_19824 (I339724,I339716);
not I_19825 (I339741,I128533);
nand I_19826 (I339758,I339741,I128527);
and I_19827 (I339775,I339577,I339758);
nor I_19828 (I339792,I339690,I339775);
DFFARX1 I_19829 (I339792,I2683,I339495,I339463,);
DFFARX1 I_19830 (I339775,I2683,I339495,I339484,);
nor I_19831 (I339837,I128533,I128536);
nor I_19832 (I339475,I339690,I339837);
or I_19833 (I339868,I128533,I128536);
nor I_19834 (I339885,I128551,I128548);
DFFARX1 I_19835 (I339885,I2683,I339495,I339911,);
not I_19836 (I339919,I339911);
nor I_19837 (I339481,I339919,I339724);
nand I_19838 (I339950,I339919,I339569);
not I_19839 (I339967,I128551);
nand I_19840 (I339984,I339967,I339673);
nand I_19841 (I340001,I339919,I339984);
nand I_19842 (I339472,I340001,I339950);
nand I_19843 (I339469,I339984,I339868);
not I_19844 (I340073,I2690);
DFFARX1 I_19845 (I375762,I2683,I340073,I340099,);
and I_19846 (I340107,I340099,I375756);
DFFARX1 I_19847 (I340107,I2683,I340073,I340056,);
DFFARX1 I_19848 (I375741,I2683,I340073,I340147,);
not I_19849 (I340155,I375747);
not I_19850 (I340172,I375759);
nand I_19851 (I340189,I340172,I340155);
nor I_19852 (I340044,I340147,I340189);
DFFARX1 I_19853 (I340189,I2683,I340073,I340229,);
not I_19854 (I340065,I340229);
not I_19855 (I340251,I375741);
nand I_19856 (I340268,I340172,I340251);
DFFARX1 I_19857 (I340268,I2683,I340073,I340294,);
not I_19858 (I340302,I340294);
not I_19859 (I340319,I375765);
nand I_19860 (I340336,I340319,I375753);
and I_19861 (I340353,I340155,I340336);
nor I_19862 (I340370,I340268,I340353);
DFFARX1 I_19863 (I340370,I2683,I340073,I340041,);
DFFARX1 I_19864 (I340353,I2683,I340073,I340062,);
nor I_19865 (I340415,I375765,I375744);
nor I_19866 (I340053,I340268,I340415);
or I_19867 (I340446,I375765,I375744);
nor I_19868 (I340463,I375750,I375744);
DFFARX1 I_19869 (I340463,I2683,I340073,I340489,);
not I_19870 (I340497,I340489);
nor I_19871 (I340059,I340497,I340302);
nand I_19872 (I340528,I340497,I340147);
not I_19873 (I340545,I375750);
nand I_19874 (I340562,I340545,I340251);
nand I_19875 (I340579,I340497,I340562);
nand I_19876 (I340050,I340579,I340528);
nand I_19877 (I340047,I340562,I340446);
not I_19878 (I340651,I2690);
DFFARX1 I_19879 (I159997,I2683,I340651,I340677,);
and I_19880 (I340685,I340677,I160012);
DFFARX1 I_19881 (I340685,I2683,I340651,I340634,);
DFFARX1 I_19882 (I160003,I2683,I340651,I340725,);
not I_19883 (I340733,I159997);
not I_19884 (I340750,I160015);
nand I_19885 (I340767,I340750,I340733);
nor I_19886 (I340622,I340725,I340767);
DFFARX1 I_19887 (I340767,I2683,I340651,I340807,);
not I_19888 (I340643,I340807);
not I_19889 (I340829,I160006);
nand I_19890 (I340846,I340750,I340829);
DFFARX1 I_19891 (I340846,I2683,I340651,I340872,);
not I_19892 (I340880,I340872);
not I_19893 (I340897,I160018);
nand I_19894 (I340914,I340897,I159994);
and I_19895 (I340931,I340733,I340914);
nor I_19896 (I340948,I340846,I340931);
DFFARX1 I_19897 (I340948,I2683,I340651,I340619,);
DFFARX1 I_19898 (I340931,I2683,I340651,I340640,);
nor I_19899 (I340993,I160018,I159994);
nor I_19900 (I340631,I340846,I340993);
or I_19901 (I341024,I160018,I159994);
nor I_19902 (I341041,I160000,I160009);
DFFARX1 I_19903 (I341041,I2683,I340651,I341067,);
not I_19904 (I341075,I341067);
nor I_19905 (I340637,I341075,I340880);
nand I_19906 (I341106,I341075,I340725);
not I_19907 (I341123,I160000);
nand I_19908 (I341140,I341123,I340829);
nand I_19909 (I341157,I341075,I341140);
nand I_19910 (I340628,I341157,I341106);
nand I_19911 (I340625,I341140,I341024);
not I_19912 (I341229,I2690);
DFFARX1 I_19913 (I205960,I2683,I341229,I341255,);
and I_19914 (I341263,I341255,I205948);
DFFARX1 I_19915 (I341263,I2683,I341229,I341212,);
DFFARX1 I_19916 (I205951,I2683,I341229,I341303,);
not I_19917 (I341311,I205945);
not I_19918 (I341328,I205969);
nand I_19919 (I341345,I341328,I341311);
nor I_19920 (I341200,I341303,I341345);
DFFARX1 I_19921 (I341345,I2683,I341229,I341385,);
not I_19922 (I341221,I341385);
not I_19923 (I341407,I205957);
nand I_19924 (I341424,I341328,I341407);
DFFARX1 I_19925 (I341424,I2683,I341229,I341450,);
not I_19926 (I341458,I341450);
not I_19927 (I341475,I205966);
nand I_19928 (I341492,I341475,I205963);
and I_19929 (I341509,I341311,I341492);
nor I_19930 (I341526,I341424,I341509);
DFFARX1 I_19931 (I341526,I2683,I341229,I341197,);
DFFARX1 I_19932 (I341509,I2683,I341229,I341218,);
nor I_19933 (I341571,I205966,I205954);
nor I_19934 (I341209,I341424,I341571);
or I_19935 (I341602,I205966,I205954);
nor I_19936 (I341619,I205945,I205948);
DFFARX1 I_19937 (I341619,I2683,I341229,I341645,);
not I_19938 (I341653,I341645);
nor I_19939 (I341215,I341653,I341458);
nand I_19940 (I341684,I341653,I341303);
not I_19941 (I341701,I205945);
nand I_19942 (I341718,I341701,I341407);
nand I_19943 (I341735,I341653,I341718);
nand I_19944 (I341206,I341735,I341684);
nand I_19945 (I341203,I341718,I341602);
not I_19946 (I341807,I2690);
DFFARX1 I_19947 (I45924,I2683,I341807,I341833,);
and I_19948 (I341841,I341833,I45948);
DFFARX1 I_19949 (I341841,I2683,I341807,I341790,);
DFFARX1 I_19950 (I45924,I2683,I341807,I341881,);
not I_19951 (I341889,I45942);
not I_19952 (I341906,I45927);
nand I_19953 (I341923,I341906,I341889);
nor I_19954 (I341778,I341881,I341923);
DFFARX1 I_19955 (I341923,I2683,I341807,I341963,);
not I_19956 (I341799,I341963);
not I_19957 (I341985,I45936);
nand I_19958 (I342002,I341906,I341985);
DFFARX1 I_19959 (I342002,I2683,I341807,I342028,);
not I_19960 (I342036,I342028);
not I_19961 (I342053,I45933);
nand I_19962 (I342070,I342053,I45930);
and I_19963 (I342087,I341889,I342070);
nor I_19964 (I342104,I342002,I342087);
DFFARX1 I_19965 (I342104,I2683,I341807,I341775,);
DFFARX1 I_19966 (I342087,I2683,I341807,I341796,);
nor I_19967 (I342149,I45933,I45939);
nor I_19968 (I341787,I342002,I342149);
or I_19969 (I342180,I45933,I45939);
nor I_19970 (I342197,I45945,I45951);
DFFARX1 I_19971 (I342197,I2683,I341807,I342223,);
not I_19972 (I342231,I342223);
nor I_19973 (I341793,I342231,I342036);
nand I_19974 (I342262,I342231,I341881);
not I_19975 (I342279,I45945);
nand I_19976 (I342296,I342279,I341985);
nand I_19977 (I342313,I342231,I342296);
nand I_19978 (I341784,I342313,I342262);
nand I_19979 (I341781,I342296,I342180);
not I_19980 (I342385,I2690);
DFFARX1 I_19981 (I396243,I2683,I342385,I342411,);
and I_19982 (I342419,I342411,I396270);
DFFARX1 I_19983 (I342419,I2683,I342385,I342368,);
DFFARX1 I_19984 (I396252,I2683,I342385,I342459,);
not I_19985 (I342467,I396261);
not I_19986 (I342484,I396264);
nand I_19987 (I342501,I342484,I342467);
nor I_19988 (I342356,I342459,I342501);
DFFARX1 I_19989 (I342501,I2683,I342385,I342541,);
not I_19990 (I342377,I342541);
not I_19991 (I342563,I396258);
nand I_19992 (I342580,I342484,I342563);
DFFARX1 I_19993 (I342580,I2683,I342385,I342606,);
not I_19994 (I342614,I342606);
not I_19995 (I342631,I396246);
nand I_19996 (I342648,I342631,I396249);
and I_19997 (I342665,I342467,I342648);
nor I_19998 (I342682,I342580,I342665);
DFFARX1 I_19999 (I342682,I2683,I342385,I342353,);
DFFARX1 I_20000 (I342665,I2683,I342385,I342374,);
nor I_20001 (I342727,I396246,I396267);
nor I_20002 (I342365,I342580,I342727);
or I_20003 (I342758,I396246,I396267);
nor I_20004 (I342775,I396255,I396243);
DFFARX1 I_20005 (I342775,I2683,I342385,I342801,);
not I_20006 (I342809,I342801);
nor I_20007 (I342371,I342809,I342614);
nand I_20008 (I342840,I342809,I342459);
not I_20009 (I342857,I396255);
nand I_20010 (I342874,I342857,I342563);
nand I_20011 (I342891,I342809,I342874);
nand I_20012 (I342362,I342891,I342840);
nand I_20013 (I342359,I342874,I342758);
not I_20014 (I342963,I2690);
DFFARX1 I_20015 (I418846,I2683,I342963,I342989,);
and I_20016 (I342997,I342989,I418828);
DFFARX1 I_20017 (I342997,I2683,I342963,I342946,);
DFFARX1 I_20018 (I418819,I2683,I342963,I343037,);
not I_20019 (I343045,I418834);
not I_20020 (I343062,I418822);
nand I_20021 (I343079,I343062,I343045);
nor I_20022 (I342934,I343037,I343079);
DFFARX1 I_20023 (I343079,I2683,I342963,I343119,);
not I_20024 (I342955,I343119);
not I_20025 (I343141,I418831);
nand I_20026 (I343158,I343062,I343141);
DFFARX1 I_20027 (I343158,I2683,I342963,I343184,);
not I_20028 (I343192,I343184);
not I_20029 (I343209,I418840);
nand I_20030 (I343226,I343209,I418819);
and I_20031 (I343243,I343045,I343226);
nor I_20032 (I343260,I343158,I343243);
DFFARX1 I_20033 (I343260,I2683,I342963,I342931,);
DFFARX1 I_20034 (I343243,I2683,I342963,I342952,);
nor I_20035 (I343305,I418840,I418843);
nor I_20036 (I342943,I343158,I343305);
or I_20037 (I343336,I418840,I418843);
nor I_20038 (I343353,I418837,I418825);
DFFARX1 I_20039 (I343353,I2683,I342963,I343379,);
not I_20040 (I343387,I343379);
nor I_20041 (I342949,I343387,I343192);
nand I_20042 (I343418,I343387,I343037);
not I_20043 (I343435,I418837);
nand I_20044 (I343452,I343435,I343141);
nand I_20045 (I343469,I343387,I343452);
nand I_20046 (I342940,I343469,I343418);
nand I_20047 (I342937,I343452,I343336);
not I_20048 (I343541,I2690);
DFFARX1 I_20049 (I417061,I2683,I343541,I343567,);
and I_20050 (I343575,I343567,I417043);
DFFARX1 I_20051 (I343575,I2683,I343541,I343524,);
DFFARX1 I_20052 (I417034,I2683,I343541,I343615,);
not I_20053 (I343623,I417049);
not I_20054 (I343640,I417037);
nand I_20055 (I343657,I343640,I343623);
nor I_20056 (I343512,I343615,I343657);
DFFARX1 I_20057 (I343657,I2683,I343541,I343697,);
not I_20058 (I343533,I343697);
not I_20059 (I343719,I417046);
nand I_20060 (I343736,I343640,I343719);
DFFARX1 I_20061 (I343736,I2683,I343541,I343762,);
not I_20062 (I343770,I343762);
not I_20063 (I343787,I417055);
nand I_20064 (I343804,I343787,I417034);
and I_20065 (I343821,I343623,I343804);
nor I_20066 (I343838,I343736,I343821);
DFFARX1 I_20067 (I343838,I2683,I343541,I343509,);
DFFARX1 I_20068 (I343821,I2683,I343541,I343530,);
nor I_20069 (I343883,I417055,I417058);
nor I_20070 (I343521,I343736,I343883);
or I_20071 (I343914,I417055,I417058);
nor I_20072 (I343931,I417052,I417040);
DFFARX1 I_20073 (I343931,I2683,I343541,I343957,);
not I_20074 (I343965,I343957);
nor I_20075 (I343527,I343965,I343770);
nand I_20076 (I343996,I343965,I343615);
not I_20077 (I344013,I417052);
nand I_20078 (I344030,I344013,I343719);
nand I_20079 (I344047,I343965,I344030);
nand I_20080 (I343518,I344047,I343996);
nand I_20081 (I343515,I344030,I343914);
not I_20082 (I344119,I2690);
DFFARX1 I_20083 (I262932,I2683,I344119,I344145,);
and I_20084 (I344153,I344145,I262938);
DFFARX1 I_20085 (I344153,I2683,I344119,I344102,);
DFFARX1 I_20086 (I262944,I2683,I344119,I344193,);
not I_20087 (I344201,I262929);
not I_20088 (I344218,I262929);
nand I_20089 (I344235,I344218,I344201);
nor I_20090 (I344090,I344193,I344235);
DFFARX1 I_20091 (I344235,I2683,I344119,I344275,);
not I_20092 (I344111,I344275);
not I_20093 (I344297,I262947);
nand I_20094 (I344314,I344218,I344297);
DFFARX1 I_20095 (I344314,I2683,I344119,I344340,);
not I_20096 (I344348,I344340);
not I_20097 (I344365,I262941);
nand I_20098 (I344382,I344365,I262932);
and I_20099 (I344399,I344201,I344382);
nor I_20100 (I344416,I344314,I344399);
DFFARX1 I_20101 (I344416,I2683,I344119,I344087,);
DFFARX1 I_20102 (I344399,I2683,I344119,I344108,);
nor I_20103 (I344461,I262941,I262950);
nor I_20104 (I344099,I344314,I344461);
or I_20105 (I344492,I262941,I262950);
nor I_20106 (I344509,I262935,I262935);
DFFARX1 I_20107 (I344509,I2683,I344119,I344535,);
not I_20108 (I344543,I344535);
nor I_20109 (I344105,I344543,I344348);
nand I_20110 (I344574,I344543,I344193);
not I_20111 (I344591,I262935);
nand I_20112 (I344608,I344591,I344297);
nand I_20113 (I344625,I344543,I344608);
nand I_20114 (I344096,I344625,I344574);
nand I_20115 (I344093,I344608,I344492);
not I_20116 (I344697,I2690);
DFFARX1 I_20117 (I389433,I2683,I344697,I344723,);
and I_20118 (I344731,I344723,I389415);
DFFARX1 I_20119 (I344731,I2683,I344697,I344680,);
DFFARX1 I_20120 (I389424,I2683,I344697,I344771,);
not I_20121 (I344779,I389409);
not I_20122 (I344796,I389421);
nand I_20123 (I344813,I344796,I344779);
nor I_20124 (I344668,I344771,I344813);
DFFARX1 I_20125 (I344813,I2683,I344697,I344853,);
not I_20126 (I344689,I344853);
not I_20127 (I344875,I389412);
nand I_20128 (I344892,I344796,I344875);
DFFARX1 I_20129 (I344892,I2683,I344697,I344918,);
not I_20130 (I344926,I344918);
not I_20131 (I344943,I389409);
nand I_20132 (I344960,I344943,I389412);
and I_20133 (I344977,I344779,I344960);
nor I_20134 (I344994,I344892,I344977);
DFFARX1 I_20135 (I344994,I2683,I344697,I344665,);
DFFARX1 I_20136 (I344977,I2683,I344697,I344686,);
nor I_20137 (I345039,I389409,I389430);
nor I_20138 (I344677,I344892,I345039);
or I_20139 (I345070,I389409,I389430);
nor I_20140 (I345087,I389418,I389427);
DFFARX1 I_20141 (I345087,I2683,I344697,I345113,);
not I_20142 (I345121,I345113);
nor I_20143 (I344683,I345121,I344926);
nand I_20144 (I345152,I345121,I344771);
not I_20145 (I345169,I389418);
nand I_20146 (I345186,I345169,I344875);
nand I_20147 (I345203,I345121,I345186);
nand I_20148 (I344674,I345203,I345152);
nand I_20149 (I344671,I345186,I345070);
not I_20150 (I345275,I2690);
DFFARX1 I_20151 (I202492,I2683,I345275,I345301,);
and I_20152 (I345309,I345301,I202480);
DFFARX1 I_20153 (I345309,I2683,I345275,I345258,);
DFFARX1 I_20154 (I202483,I2683,I345275,I345349,);
not I_20155 (I345357,I202477);
not I_20156 (I345374,I202501);
nand I_20157 (I345391,I345374,I345357);
nor I_20158 (I345246,I345349,I345391);
DFFARX1 I_20159 (I345391,I2683,I345275,I345431,);
not I_20160 (I345267,I345431);
not I_20161 (I345453,I202489);
nand I_20162 (I345470,I345374,I345453);
DFFARX1 I_20163 (I345470,I2683,I345275,I345496,);
not I_20164 (I345504,I345496);
not I_20165 (I345521,I202498);
nand I_20166 (I345538,I345521,I202495);
and I_20167 (I345555,I345357,I345538);
nor I_20168 (I345572,I345470,I345555);
DFFARX1 I_20169 (I345572,I2683,I345275,I345243,);
DFFARX1 I_20170 (I345555,I2683,I345275,I345264,);
nor I_20171 (I345617,I202498,I202486);
nor I_20172 (I345255,I345470,I345617);
or I_20173 (I345648,I202498,I202486);
nor I_20174 (I345665,I202477,I202480);
DFFARX1 I_20175 (I345665,I2683,I345275,I345691,);
not I_20176 (I345699,I345691);
nor I_20177 (I345261,I345699,I345504);
nand I_20178 (I345730,I345699,I345349);
not I_20179 (I345747,I202477);
nand I_20180 (I345764,I345747,I345453);
nand I_20181 (I345781,I345699,I345764);
nand I_20182 (I345252,I345781,I345730);
nand I_20183 (I345249,I345764,I345648);
not I_20184 (I345853,I2690);
DFFARX1 I_20185 (I270432,I2683,I345853,I345879,);
and I_20186 (I345887,I345879,I270426);
DFFARX1 I_20187 (I345887,I2683,I345853,I345836,);
DFFARX1 I_20188 (I270444,I2683,I345853,I345927,);
not I_20189 (I345935,I270435);
not I_20190 (I345952,I270447);
nand I_20191 (I345969,I345952,I345935);
nor I_20192 (I345824,I345927,I345969);
DFFARX1 I_20193 (I345969,I2683,I345853,I346009,);
not I_20194 (I345845,I346009);
not I_20195 (I346031,I270453);
nand I_20196 (I346048,I345952,I346031);
DFFARX1 I_20197 (I346048,I2683,I345853,I346074,);
not I_20198 (I346082,I346074);
not I_20199 (I346099,I270429);
nand I_20200 (I346116,I346099,I270450);
and I_20201 (I346133,I345935,I346116);
nor I_20202 (I346150,I346048,I346133);
DFFARX1 I_20203 (I346150,I2683,I345853,I345821,);
DFFARX1 I_20204 (I346133,I2683,I345853,I345842,);
nor I_20205 (I346195,I270429,I270441);
nor I_20206 (I345833,I346048,I346195);
or I_20207 (I346226,I270429,I270441);
nor I_20208 (I346243,I270426,I270438);
DFFARX1 I_20209 (I346243,I2683,I345853,I346269,);
not I_20210 (I346277,I346269);
nor I_20211 (I345839,I346277,I346082);
nand I_20212 (I346308,I346277,I345927);
not I_20213 (I346325,I270426);
nand I_20214 (I346342,I346325,I346031);
nand I_20215 (I346359,I346277,I346342);
nand I_20216 (I345830,I346359,I346308);
nand I_20217 (I345827,I346342,I346226);
not I_20218 (I346431,I2690);
DFFARX1 I_20219 (I305962,I2683,I346431,I346457,);
and I_20220 (I346465,I346457,I305956);
DFFARX1 I_20221 (I346465,I2683,I346431,I346414,);
DFFARX1 I_20222 (I305974,I2683,I346431,I346505,);
not I_20223 (I346513,I305965);
not I_20224 (I346530,I305977);
nand I_20225 (I346547,I346530,I346513);
nor I_20226 (I346402,I346505,I346547);
DFFARX1 I_20227 (I346547,I2683,I346431,I346587,);
not I_20228 (I346423,I346587);
not I_20229 (I346609,I305983);
nand I_20230 (I346626,I346530,I346609);
DFFARX1 I_20231 (I346626,I2683,I346431,I346652,);
not I_20232 (I346660,I346652);
not I_20233 (I346677,I305959);
nand I_20234 (I346694,I346677,I305980);
and I_20235 (I346711,I346513,I346694);
nor I_20236 (I346728,I346626,I346711);
DFFARX1 I_20237 (I346728,I2683,I346431,I346399,);
DFFARX1 I_20238 (I346711,I2683,I346431,I346420,);
nor I_20239 (I346773,I305959,I305971);
nor I_20240 (I346411,I346626,I346773);
or I_20241 (I346804,I305959,I305971);
nor I_20242 (I346821,I305956,I305968);
DFFARX1 I_20243 (I346821,I2683,I346431,I346847,);
not I_20244 (I346855,I346847);
nor I_20245 (I346417,I346855,I346660);
nand I_20246 (I346886,I346855,I346505);
not I_20247 (I346903,I305956);
nand I_20248 (I346920,I346903,I346609);
nand I_20249 (I346937,I346855,I346920);
nand I_20250 (I346408,I346937,I346886);
nand I_20251 (I346405,I346920,I346804);
not I_20252 (I347009,I2690);
DFFARX1 I_20253 (I412896,I2683,I347009,I347035,);
and I_20254 (I347043,I347035,I412878);
DFFARX1 I_20255 (I347043,I2683,I347009,I346992,);
DFFARX1 I_20256 (I412869,I2683,I347009,I347083,);
not I_20257 (I347091,I412884);
not I_20258 (I347108,I412872);
nand I_20259 (I347125,I347108,I347091);
nor I_20260 (I346980,I347083,I347125);
DFFARX1 I_20261 (I347125,I2683,I347009,I347165,);
not I_20262 (I347001,I347165);
not I_20263 (I347187,I412881);
nand I_20264 (I347204,I347108,I347187);
DFFARX1 I_20265 (I347204,I2683,I347009,I347230,);
not I_20266 (I347238,I347230);
not I_20267 (I347255,I412890);
nand I_20268 (I347272,I347255,I412869);
and I_20269 (I347289,I347091,I347272);
nor I_20270 (I347306,I347204,I347289);
DFFARX1 I_20271 (I347306,I2683,I347009,I346977,);
DFFARX1 I_20272 (I347289,I2683,I347009,I346998,);
nor I_20273 (I347351,I412890,I412893);
nor I_20274 (I346989,I347204,I347351);
or I_20275 (I347382,I412890,I412893);
nor I_20276 (I347399,I412887,I412875);
DFFARX1 I_20277 (I347399,I2683,I347009,I347425,);
not I_20278 (I347433,I347425);
nor I_20279 (I346995,I347433,I347238);
nand I_20280 (I347464,I347433,I347083);
not I_20281 (I347481,I412887);
nand I_20282 (I347498,I347481,I347187);
nand I_20283 (I347515,I347433,I347498);
nand I_20284 (I346986,I347515,I347464);
nand I_20285 (I346983,I347498,I347382);
not I_20286 (I347587,I2690);
DFFARX1 I_20287 (I398021,I2683,I347587,I347613,);
and I_20288 (I347621,I347613,I398003);
DFFARX1 I_20289 (I347621,I2683,I347587,I347570,);
DFFARX1 I_20290 (I397994,I2683,I347587,I347661,);
not I_20291 (I347669,I398009);
not I_20292 (I347686,I397997);
nand I_20293 (I347703,I347686,I347669);
nor I_20294 (I347558,I347661,I347703);
DFFARX1 I_20295 (I347703,I2683,I347587,I347743,);
not I_20296 (I347579,I347743);
not I_20297 (I347765,I398006);
nand I_20298 (I347782,I347686,I347765);
DFFARX1 I_20299 (I347782,I2683,I347587,I347808,);
not I_20300 (I347816,I347808);
not I_20301 (I347833,I398015);
nand I_20302 (I347850,I347833,I397994);
and I_20303 (I347867,I347669,I347850);
nor I_20304 (I347884,I347782,I347867);
DFFARX1 I_20305 (I347884,I2683,I347587,I347555,);
DFFARX1 I_20306 (I347867,I2683,I347587,I347576,);
nor I_20307 (I347929,I398015,I398018);
nor I_20308 (I347567,I347782,I347929);
or I_20309 (I347960,I398015,I398018);
nor I_20310 (I347977,I398012,I398000);
DFFARX1 I_20311 (I347977,I2683,I347587,I348003,);
not I_20312 (I348011,I348003);
nor I_20313 (I347573,I348011,I347816);
nand I_20314 (I348042,I348011,I347661);
not I_20315 (I348059,I398012);
nand I_20316 (I348076,I348059,I347765);
nand I_20317 (I348093,I348011,I348076);
nand I_20318 (I347564,I348093,I348042);
nand I_20319 (I347561,I348076,I347960);
not I_20320 (I348165,I2690);
DFFARX1 I_20321 (I306608,I2683,I348165,I348191,);
and I_20322 (I348199,I348191,I306602);
DFFARX1 I_20323 (I348199,I2683,I348165,I348148,);
DFFARX1 I_20324 (I306620,I2683,I348165,I348239,);
not I_20325 (I348247,I306611);
not I_20326 (I348264,I306623);
nand I_20327 (I348281,I348264,I348247);
nor I_20328 (I348136,I348239,I348281);
DFFARX1 I_20329 (I348281,I2683,I348165,I348321,);
not I_20330 (I348157,I348321);
not I_20331 (I348343,I306629);
nand I_20332 (I348360,I348264,I348343);
DFFARX1 I_20333 (I348360,I2683,I348165,I348386,);
not I_20334 (I348394,I348386);
not I_20335 (I348411,I306605);
nand I_20336 (I348428,I348411,I306626);
and I_20337 (I348445,I348247,I348428);
nor I_20338 (I348462,I348360,I348445);
DFFARX1 I_20339 (I348462,I2683,I348165,I348133,);
DFFARX1 I_20340 (I348445,I2683,I348165,I348154,);
nor I_20341 (I348507,I306605,I306617);
nor I_20342 (I348145,I348360,I348507);
or I_20343 (I348538,I306605,I306617);
nor I_20344 (I348555,I306602,I306614);
DFFARX1 I_20345 (I348555,I2683,I348165,I348581,);
not I_20346 (I348589,I348581);
nor I_20347 (I348151,I348589,I348394);
nand I_20348 (I348620,I348589,I348239);
not I_20349 (I348637,I306602);
nand I_20350 (I348654,I348637,I348343);
nand I_20351 (I348671,I348589,I348654);
nand I_20352 (I348142,I348671,I348620);
nand I_20353 (I348139,I348654,I348538);
not I_20354 (I348743,I2690);
DFFARX1 I_20355 (I31515,I2683,I348743,I348769,);
and I_20356 (I348777,I348769,I31491);
DFFARX1 I_20357 (I348777,I2683,I348743,I348726,);
DFFARX1 I_20358 (I31509,I2683,I348743,I348817,);
not I_20359 (I348825,I31497);
not I_20360 (I348842,I31494);
nand I_20361 (I348859,I348842,I348825);
nor I_20362 (I348714,I348817,I348859);
DFFARX1 I_20363 (I348859,I2683,I348743,I348899,);
not I_20364 (I348735,I348899);
not I_20365 (I348921,I31503);
nand I_20366 (I348938,I348842,I348921);
DFFARX1 I_20367 (I348938,I2683,I348743,I348964,);
not I_20368 (I348972,I348964);
not I_20369 (I348989,I31494);
nand I_20370 (I349006,I348989,I31512);
and I_20371 (I349023,I348825,I349006);
nor I_20372 (I349040,I348938,I349023);
DFFARX1 I_20373 (I349040,I2683,I348743,I348711,);
DFFARX1 I_20374 (I349023,I2683,I348743,I348732,);
nor I_20375 (I349085,I31494,I31506);
nor I_20376 (I348723,I348938,I349085);
or I_20377 (I349116,I31494,I31506);
nor I_20378 (I349133,I31500,I31491);
DFFARX1 I_20379 (I349133,I2683,I348743,I349159,);
not I_20380 (I349167,I349159);
nor I_20381 (I348729,I349167,I348972);
nand I_20382 (I349198,I349167,I348817);
not I_20383 (I349215,I31500);
nand I_20384 (I349232,I349215,I348921);
nand I_20385 (I349249,I349167,I349232);
nand I_20386 (I348720,I349249,I349198);
nand I_20387 (I348717,I349232,I349116);
not I_20388 (I349321,I2690);
DFFARX1 I_20389 (I37312,I2683,I349321,I349347,);
and I_20390 (I349355,I349347,I37288);
DFFARX1 I_20391 (I349355,I2683,I349321,I349304,);
DFFARX1 I_20392 (I37306,I2683,I349321,I349395,);
not I_20393 (I349403,I37294);
not I_20394 (I349420,I37291);
nand I_20395 (I349437,I349420,I349403);
nor I_20396 (I349292,I349395,I349437);
DFFARX1 I_20397 (I349437,I2683,I349321,I349477,);
not I_20398 (I349313,I349477);
not I_20399 (I349499,I37300);
nand I_20400 (I349516,I349420,I349499);
DFFARX1 I_20401 (I349516,I2683,I349321,I349542,);
not I_20402 (I349550,I349542);
not I_20403 (I349567,I37291);
nand I_20404 (I349584,I349567,I37309);
and I_20405 (I349601,I349403,I349584);
nor I_20406 (I349618,I349516,I349601);
DFFARX1 I_20407 (I349618,I2683,I349321,I349289,);
DFFARX1 I_20408 (I349601,I2683,I349321,I349310,);
nor I_20409 (I349663,I37291,I37303);
nor I_20410 (I349301,I349516,I349663);
or I_20411 (I349694,I37291,I37303);
nor I_20412 (I349711,I37297,I37288);
DFFARX1 I_20413 (I349711,I2683,I349321,I349737,);
not I_20414 (I349745,I349737);
nor I_20415 (I349307,I349745,I349550);
nand I_20416 (I349776,I349745,I349395);
not I_20417 (I349793,I37297);
nand I_20418 (I349810,I349793,I349499);
nand I_20419 (I349827,I349745,I349810);
nand I_20420 (I349298,I349827,I349776);
nand I_20421 (I349295,I349810,I349694);
not I_20422 (I349899,I2690);
DFFARX1 I_20423 (I150831,I2683,I349899,I349925,);
and I_20424 (I349933,I349925,I150846);
DFFARX1 I_20425 (I349933,I2683,I349899,I349882,);
DFFARX1 I_20426 (I150849,I2683,I349899,I349973,);
not I_20427 (I349981,I150843);
not I_20428 (I349998,I150858);
nand I_20429 (I350015,I349998,I349981);
nor I_20430 (I349870,I349973,I350015);
DFFARX1 I_20431 (I350015,I2683,I349899,I350055,);
not I_20432 (I349891,I350055);
not I_20433 (I350077,I150834);
nand I_20434 (I350094,I349998,I350077);
DFFARX1 I_20435 (I350094,I2683,I349899,I350120,);
not I_20436 (I350128,I350120);
not I_20437 (I350145,I150837);
nand I_20438 (I350162,I350145,I150831);
and I_20439 (I350179,I349981,I350162);
nor I_20440 (I350196,I350094,I350179);
DFFARX1 I_20441 (I350196,I2683,I349899,I349867,);
DFFARX1 I_20442 (I350179,I2683,I349899,I349888,);
nor I_20443 (I350241,I150837,I150840);
nor I_20444 (I349879,I350094,I350241);
or I_20445 (I350272,I150837,I150840);
nor I_20446 (I350289,I150855,I150852);
DFFARX1 I_20447 (I350289,I2683,I349899,I350315,);
not I_20448 (I350323,I350315);
nor I_20449 (I349885,I350323,I350128);
nand I_20450 (I350354,I350323,I349973);
not I_20451 (I350371,I150855);
nand I_20452 (I350388,I350371,I350077);
nand I_20453 (I350405,I350323,I350388);
nand I_20454 (I349876,I350405,I350354);
nand I_20455 (I349873,I350388,I350272);
not I_20456 (I350477,I2690);
DFFARX1 I_20457 (I116382,I2683,I350477,I350503,);
and I_20458 (I350511,I350503,I116367);
DFFARX1 I_20459 (I350511,I2683,I350477,I350460,);
DFFARX1 I_20460 (I116373,I2683,I350477,I350551,);
not I_20461 (I350559,I116355);
not I_20462 (I350576,I116376);
nand I_20463 (I350593,I350576,I350559);
nor I_20464 (I350448,I350551,I350593);
DFFARX1 I_20465 (I350593,I2683,I350477,I350633,);
not I_20466 (I350469,I350633);
not I_20467 (I350655,I116379);
nand I_20468 (I350672,I350576,I350655);
DFFARX1 I_20469 (I350672,I2683,I350477,I350698,);
not I_20470 (I350706,I350698);
not I_20471 (I350723,I116370);
nand I_20472 (I350740,I350723,I116358);
and I_20473 (I350757,I350559,I350740);
nor I_20474 (I350774,I350672,I350757);
DFFARX1 I_20475 (I350774,I2683,I350477,I350445,);
DFFARX1 I_20476 (I350757,I2683,I350477,I350466,);
nor I_20477 (I350819,I116370,I116364);
nor I_20478 (I350457,I350672,I350819);
or I_20479 (I350850,I116370,I116364);
nor I_20480 (I350867,I116361,I116355);
DFFARX1 I_20481 (I350867,I2683,I350477,I350893,);
not I_20482 (I350901,I350893);
nor I_20483 (I350463,I350901,I350706);
nand I_20484 (I350932,I350901,I350551);
not I_20485 (I350949,I116361);
nand I_20486 (I350966,I350949,I350655);
nand I_20487 (I350983,I350901,I350966);
nand I_20488 (I350454,I350983,I350932);
nand I_20489 (I350451,I350966,I350850);
not I_20490 (I351055,I2690);
DFFARX1 I_20491 (I26772,I2683,I351055,I351081,);
and I_20492 (I351089,I351081,I26748);
DFFARX1 I_20493 (I351089,I2683,I351055,I351038,);
DFFARX1 I_20494 (I26766,I2683,I351055,I351129,);
not I_20495 (I351137,I26754);
not I_20496 (I351154,I26751);
nand I_20497 (I351171,I351154,I351137);
nor I_20498 (I351026,I351129,I351171);
DFFARX1 I_20499 (I351171,I2683,I351055,I351211,);
not I_20500 (I351047,I351211);
not I_20501 (I351233,I26760);
nand I_20502 (I351250,I351154,I351233);
DFFARX1 I_20503 (I351250,I2683,I351055,I351276,);
not I_20504 (I351284,I351276);
not I_20505 (I351301,I26751);
nand I_20506 (I351318,I351301,I26769);
and I_20507 (I351335,I351137,I351318);
nor I_20508 (I351352,I351250,I351335);
DFFARX1 I_20509 (I351352,I2683,I351055,I351023,);
DFFARX1 I_20510 (I351335,I2683,I351055,I351044,);
nor I_20511 (I351397,I26751,I26763);
nor I_20512 (I351035,I351250,I351397);
or I_20513 (I351428,I26751,I26763);
nor I_20514 (I351445,I26757,I26748);
DFFARX1 I_20515 (I351445,I2683,I351055,I351471,);
not I_20516 (I351479,I351471);
nor I_20517 (I351041,I351479,I351284);
nand I_20518 (I351510,I351479,I351129);
not I_20519 (I351527,I26757);
nand I_20520 (I351544,I351527,I351233);
nand I_20521 (I351561,I351479,I351544);
nand I_20522 (I351032,I351561,I351510);
nand I_20523 (I351029,I351544,I351428);
not I_20524 (I351633,I2690);
DFFARX1 I_20525 (I98464,I2683,I351633,I351659,);
and I_20526 (I351667,I351659,I98449);
DFFARX1 I_20527 (I351667,I2683,I351633,I351616,);
DFFARX1 I_20528 (I98455,I2683,I351633,I351707,);
not I_20529 (I351715,I98437);
not I_20530 (I351732,I98458);
nand I_20531 (I351749,I351732,I351715);
nor I_20532 (I351604,I351707,I351749);
DFFARX1 I_20533 (I351749,I2683,I351633,I351789,);
not I_20534 (I351625,I351789);
not I_20535 (I351811,I98461);
nand I_20536 (I351828,I351732,I351811);
DFFARX1 I_20537 (I351828,I2683,I351633,I351854,);
not I_20538 (I351862,I351854);
not I_20539 (I351879,I98452);
nand I_20540 (I351896,I351879,I98440);
and I_20541 (I351913,I351715,I351896);
nor I_20542 (I351930,I351828,I351913);
DFFARX1 I_20543 (I351930,I2683,I351633,I351601,);
DFFARX1 I_20544 (I351913,I2683,I351633,I351622,);
nor I_20545 (I351975,I98452,I98446);
nor I_20546 (I351613,I351828,I351975);
or I_20547 (I352006,I98452,I98446);
nor I_20548 (I352023,I98443,I98437);
DFFARX1 I_20549 (I352023,I2683,I351633,I352049,);
not I_20550 (I352057,I352049);
nor I_20551 (I351619,I352057,I351862);
nand I_20552 (I352088,I352057,I351707);
not I_20553 (I352105,I98443);
nand I_20554 (I352122,I352105,I351811);
nand I_20555 (I352139,I352057,I352122);
nand I_20556 (I351610,I352139,I352088);
nand I_20557 (I351607,I352122,I352006);
not I_20558 (I352211,I2690);
DFFARX1 I_20559 (I225034,I2683,I352211,I352237,);
and I_20560 (I352245,I352237,I225022);
DFFARX1 I_20561 (I352245,I2683,I352211,I352194,);
DFFARX1 I_20562 (I225025,I2683,I352211,I352285,);
not I_20563 (I352293,I225019);
not I_20564 (I352310,I225043);
nand I_20565 (I352327,I352310,I352293);
nor I_20566 (I352182,I352285,I352327);
DFFARX1 I_20567 (I352327,I2683,I352211,I352367,);
not I_20568 (I352203,I352367);
not I_20569 (I352389,I225031);
nand I_20570 (I352406,I352310,I352389);
DFFARX1 I_20571 (I352406,I2683,I352211,I352432,);
not I_20572 (I352440,I352432);
not I_20573 (I352457,I225040);
nand I_20574 (I352474,I352457,I225037);
and I_20575 (I352491,I352293,I352474);
nor I_20576 (I352508,I352406,I352491);
DFFARX1 I_20577 (I352508,I2683,I352211,I352179,);
DFFARX1 I_20578 (I352491,I2683,I352211,I352200,);
nor I_20579 (I352553,I225040,I225028);
nor I_20580 (I352191,I352406,I352553);
or I_20581 (I352584,I225040,I225028);
nor I_20582 (I352601,I225019,I225022);
DFFARX1 I_20583 (I352601,I2683,I352211,I352627,);
not I_20584 (I352635,I352627);
nor I_20585 (I352197,I352635,I352440);
nand I_20586 (I352666,I352635,I352285);
not I_20587 (I352683,I225019);
nand I_20588 (I352700,I352683,I352389);
nand I_20589 (I352717,I352635,I352700);
nand I_20590 (I352188,I352717,I352666);
nand I_20591 (I352185,I352700,I352584);
not I_20592 (I352789,I2690);
DFFARX1 I_20593 (I380185,I2683,I352789,I352815,);
and I_20594 (I352823,I352815,I380167);
DFFARX1 I_20595 (I352823,I2683,I352789,I352772,);
DFFARX1 I_20596 (I380176,I2683,I352789,I352863,);
not I_20597 (I352871,I380161);
not I_20598 (I352888,I380173);
nand I_20599 (I352905,I352888,I352871);
nor I_20600 (I352760,I352863,I352905);
DFFARX1 I_20601 (I352905,I2683,I352789,I352945,);
not I_20602 (I352781,I352945);
not I_20603 (I352967,I380164);
nand I_20604 (I352984,I352888,I352967);
DFFARX1 I_20605 (I352984,I2683,I352789,I353010,);
not I_20606 (I353018,I353010);
not I_20607 (I353035,I380161);
nand I_20608 (I353052,I353035,I380164);
and I_20609 (I353069,I352871,I353052);
nor I_20610 (I353086,I352984,I353069);
DFFARX1 I_20611 (I353086,I2683,I352789,I352757,);
DFFARX1 I_20612 (I353069,I2683,I352789,I352778,);
nor I_20613 (I353131,I380161,I380182);
nor I_20614 (I352769,I352984,I353131);
or I_20615 (I353162,I380161,I380182);
nor I_20616 (I353179,I380170,I380179);
DFFARX1 I_20617 (I353179,I2683,I352789,I353205,);
not I_20618 (I353213,I353205);
nor I_20619 (I352775,I353213,I353018);
nand I_20620 (I353244,I353213,I352863);
not I_20621 (I353261,I380170);
nand I_20622 (I353278,I353261,I352967);
nand I_20623 (I353295,I353213,I353278);
nand I_20624 (I352766,I353295,I353244);
nand I_20625 (I352763,I353278,I353162);
not I_20626 (I353367,I2690);
DFFARX1 I_20627 (I43109,I2683,I353367,I353393,);
and I_20628 (I353401,I353393,I43085);
DFFARX1 I_20629 (I353401,I2683,I353367,I353350,);
DFFARX1 I_20630 (I43103,I2683,I353367,I353441,);
not I_20631 (I353449,I43091);
not I_20632 (I353466,I43088);
nand I_20633 (I353483,I353466,I353449);
nor I_20634 (I353338,I353441,I353483);
DFFARX1 I_20635 (I353483,I2683,I353367,I353523,);
not I_20636 (I353359,I353523);
not I_20637 (I353545,I43097);
nand I_20638 (I353562,I353466,I353545);
DFFARX1 I_20639 (I353562,I2683,I353367,I353588,);
not I_20640 (I353596,I353588);
not I_20641 (I353613,I43088);
nand I_20642 (I353630,I353613,I43106);
and I_20643 (I353647,I353449,I353630);
nor I_20644 (I353664,I353562,I353647);
DFFARX1 I_20645 (I353664,I2683,I353367,I353335,);
DFFARX1 I_20646 (I353647,I2683,I353367,I353356,);
nor I_20647 (I353709,I43088,I43100);
nor I_20648 (I353347,I353562,I353709);
or I_20649 (I353740,I43088,I43100);
nor I_20650 (I353757,I43094,I43085);
DFFARX1 I_20651 (I353757,I2683,I353367,I353783,);
not I_20652 (I353791,I353783);
nor I_20653 (I353353,I353791,I353596);
nand I_20654 (I353822,I353791,I353441);
not I_20655 (I353839,I43094);
nand I_20656 (I353856,I353839,I353545);
nand I_20657 (I353873,I353791,I353856);
nand I_20658 (I353344,I353873,I353822);
nand I_20659 (I353341,I353856,I353740);
not I_20660 (I353945,I2690);
DFFARX1 I_20661 (I45329,I2683,I353945,I353971,);
and I_20662 (I353979,I353971,I45353);
DFFARX1 I_20663 (I353979,I2683,I353945,I353928,);
DFFARX1 I_20664 (I45329,I2683,I353945,I354019,);
not I_20665 (I354027,I45347);
not I_20666 (I354044,I45332);
nand I_20667 (I354061,I354044,I354027);
nor I_20668 (I353916,I354019,I354061);
DFFARX1 I_20669 (I354061,I2683,I353945,I354101,);
not I_20670 (I353937,I354101);
not I_20671 (I354123,I45341);
nand I_20672 (I354140,I354044,I354123);
DFFARX1 I_20673 (I354140,I2683,I353945,I354166,);
not I_20674 (I354174,I354166);
not I_20675 (I354191,I45338);
nand I_20676 (I354208,I354191,I45335);
and I_20677 (I354225,I354027,I354208);
nor I_20678 (I354242,I354140,I354225);
DFFARX1 I_20679 (I354242,I2683,I353945,I353913,);
DFFARX1 I_20680 (I354225,I2683,I353945,I353934,);
nor I_20681 (I354287,I45338,I45344);
nor I_20682 (I353925,I354140,I354287);
or I_20683 (I354318,I45338,I45344);
nor I_20684 (I354335,I45350,I45356);
DFFARX1 I_20685 (I354335,I2683,I353945,I354361,);
not I_20686 (I354369,I354361);
nor I_20687 (I353931,I354369,I354174);
nand I_20688 (I354400,I354369,I354019);
not I_20689 (I354417,I45350);
nand I_20690 (I354434,I354417,I354123);
nand I_20691 (I354451,I354369,I354434);
nand I_20692 (I353922,I354451,I354400);
nand I_20693 (I353919,I354434,I354318);
not I_20694 (I354523,I2690);
DFFARX1 I_20695 (I254500,I2683,I354523,I354549,);
and I_20696 (I354557,I354549,I254506);
DFFARX1 I_20697 (I354557,I2683,I354523,I354506,);
DFFARX1 I_20698 (I254512,I2683,I354523,I354597,);
not I_20699 (I354605,I254497);
not I_20700 (I354622,I254497);
nand I_20701 (I354639,I354622,I354605);
nor I_20702 (I354494,I354597,I354639);
DFFARX1 I_20703 (I354639,I2683,I354523,I354679,);
not I_20704 (I354515,I354679);
not I_20705 (I354701,I254515);
nand I_20706 (I354718,I354622,I354701);
DFFARX1 I_20707 (I354718,I2683,I354523,I354744,);
not I_20708 (I354752,I354744);
not I_20709 (I354769,I254509);
nand I_20710 (I354786,I354769,I254500);
and I_20711 (I354803,I354605,I354786);
nor I_20712 (I354820,I354718,I354803);
DFFARX1 I_20713 (I354820,I2683,I354523,I354491,);
DFFARX1 I_20714 (I354803,I2683,I354523,I354512,);
nor I_20715 (I354865,I254509,I254518);
nor I_20716 (I354503,I354718,I354865);
or I_20717 (I354896,I254509,I254518);
nor I_20718 (I354913,I254503,I254503);
DFFARX1 I_20719 (I354913,I2683,I354523,I354939,);
not I_20720 (I354947,I354939);
nor I_20721 (I354509,I354947,I354752);
nand I_20722 (I354978,I354947,I354597);
not I_20723 (I354995,I254503);
nand I_20724 (I355012,I354995,I354701);
nand I_20725 (I355029,I354947,I355012);
nand I_20726 (I354500,I355029,I354978);
nand I_20727 (I354497,I355012,I354896);
not I_20728 (I355101,I2690);
DFFARX1 I_20729 (I183418,I2683,I355101,I355127,);
and I_20730 (I355135,I355127,I183406);
DFFARX1 I_20731 (I355135,I2683,I355101,I355084,);
DFFARX1 I_20732 (I183421,I2683,I355101,I355175,);
not I_20733 (I355183,I183412);
not I_20734 (I355200,I183403);
nand I_20735 (I355217,I355200,I355183);
nor I_20736 (I355072,I355175,I355217);
DFFARX1 I_20737 (I355217,I2683,I355101,I355257,);
not I_20738 (I355093,I355257);
not I_20739 (I355279,I183409);
nand I_20740 (I355296,I355200,I355279);
DFFARX1 I_20741 (I355296,I2683,I355101,I355322,);
not I_20742 (I355330,I355322);
not I_20743 (I355347,I183424);
nand I_20744 (I355364,I355347,I183427);
and I_20745 (I355381,I355183,I355364);
nor I_20746 (I355398,I355296,I355381);
DFFARX1 I_20747 (I355398,I2683,I355101,I355069,);
DFFARX1 I_20748 (I355381,I2683,I355101,I355090,);
nor I_20749 (I355443,I183424,I183403);
nor I_20750 (I355081,I355296,I355443);
or I_20751 (I355474,I183424,I183403);
nor I_20752 (I355491,I183415,I183406);
DFFARX1 I_20753 (I355491,I2683,I355101,I355517,);
not I_20754 (I355525,I355517);
nor I_20755 (I355087,I355525,I355330);
nand I_20756 (I355556,I355525,I355175);
not I_20757 (I355573,I183415);
nand I_20758 (I355590,I355573,I355279);
nand I_20759 (I355607,I355525,I355590);
nand I_20760 (I355078,I355607,I355556);
nand I_20761 (I355075,I355590,I355474);
not I_20762 (I355679,I2690);
DFFARX1 I_20763 (I277538,I2683,I355679,I355705,);
and I_20764 (I355713,I355705,I277532);
DFFARX1 I_20765 (I355713,I2683,I355679,I355662,);
DFFARX1 I_20766 (I277550,I2683,I355679,I355753,);
not I_20767 (I355761,I277541);
not I_20768 (I355778,I277553);
nand I_20769 (I355795,I355778,I355761);
nor I_20770 (I355650,I355753,I355795);
DFFARX1 I_20771 (I355795,I2683,I355679,I355835,);
not I_20772 (I355671,I355835);
not I_20773 (I355857,I277559);
nand I_20774 (I355874,I355778,I355857);
DFFARX1 I_20775 (I355874,I2683,I355679,I355900,);
not I_20776 (I355908,I355900);
not I_20777 (I355925,I277535);
nand I_20778 (I355942,I355925,I277556);
and I_20779 (I355959,I355761,I355942);
nor I_20780 (I355976,I355874,I355959);
DFFARX1 I_20781 (I355976,I2683,I355679,I355647,);
DFFARX1 I_20782 (I355959,I2683,I355679,I355668,);
nor I_20783 (I356021,I277535,I277547);
nor I_20784 (I355659,I355874,I356021);
or I_20785 (I356052,I277535,I277547);
nor I_20786 (I356069,I277532,I277544);
DFFARX1 I_20787 (I356069,I2683,I355679,I356095,);
not I_20788 (I356103,I356095);
nor I_20789 (I355665,I356103,I355908);
nand I_20790 (I356134,I356103,I355753);
not I_20791 (I356151,I277532);
nand I_20792 (I356168,I356151,I355857);
nand I_20793 (I356185,I356103,I356168);
nand I_20794 (I355656,I356185,I356134);
nand I_20795 (I355653,I356168,I356052);
not I_20796 (I356257,I2690);
DFFARX1 I_20797 (I397426,I2683,I356257,I356283,);
and I_20798 (I356291,I356283,I397408);
DFFARX1 I_20799 (I356291,I2683,I356257,I356240,);
DFFARX1 I_20800 (I397399,I2683,I356257,I356331,);
not I_20801 (I356339,I397414);
not I_20802 (I356356,I397402);
nand I_20803 (I356373,I356356,I356339);
nor I_20804 (I356228,I356331,I356373);
DFFARX1 I_20805 (I356373,I2683,I356257,I356413,);
not I_20806 (I356249,I356413);
not I_20807 (I356435,I397411);
nand I_20808 (I356452,I356356,I356435);
DFFARX1 I_20809 (I356452,I2683,I356257,I356478,);
not I_20810 (I356486,I356478);
not I_20811 (I356503,I397420);
nand I_20812 (I356520,I356503,I397399);
and I_20813 (I356537,I356339,I356520);
nor I_20814 (I356554,I356452,I356537);
DFFARX1 I_20815 (I356554,I2683,I356257,I356225,);
DFFARX1 I_20816 (I356537,I2683,I356257,I356246,);
nor I_20817 (I356599,I397420,I397423);
nor I_20818 (I356237,I356452,I356599);
or I_20819 (I356630,I397420,I397423);
nor I_20820 (I356647,I397417,I397405);
DFFARX1 I_20821 (I356647,I2683,I356257,I356673,);
not I_20822 (I356681,I356673);
nor I_20823 (I356243,I356681,I356486);
nand I_20824 (I356712,I356681,I356331);
not I_20825 (I356729,I397417);
nand I_20826 (I356746,I356729,I356435);
nand I_20827 (I356763,I356681,I356746);
nand I_20828 (I356234,I356763,I356712);
nand I_20829 (I356231,I356746,I356630);
not I_20830 (I356835,I2690);
DFFARX1 I_20831 (I408731,I2683,I356835,I356861,);
and I_20832 (I356869,I356861,I408713);
DFFARX1 I_20833 (I356869,I2683,I356835,I356818,);
DFFARX1 I_20834 (I408704,I2683,I356835,I356909,);
not I_20835 (I356917,I408719);
not I_20836 (I356934,I408707);
nand I_20837 (I356951,I356934,I356917);
nor I_20838 (I356806,I356909,I356951);
DFFARX1 I_20839 (I356951,I2683,I356835,I356991,);
not I_20840 (I356827,I356991);
not I_20841 (I357013,I408716);
nand I_20842 (I357030,I356934,I357013);
DFFARX1 I_20843 (I357030,I2683,I356835,I357056,);
not I_20844 (I357064,I357056);
not I_20845 (I357081,I408725);
nand I_20846 (I357098,I357081,I408704);
and I_20847 (I357115,I356917,I357098);
nor I_20848 (I357132,I357030,I357115);
DFFARX1 I_20849 (I357132,I2683,I356835,I356803,);
DFFARX1 I_20850 (I357115,I2683,I356835,I356824,);
nor I_20851 (I357177,I408725,I408728);
nor I_20852 (I356815,I357030,I357177);
or I_20853 (I357208,I408725,I408728);
nor I_20854 (I357225,I408722,I408710);
DFFARX1 I_20855 (I357225,I2683,I356835,I357251,);
not I_20856 (I357259,I357251);
nor I_20857 (I356821,I357259,I357064);
nand I_20858 (I357290,I357259,I356909);
not I_20859 (I357307,I408722);
nand I_20860 (I357324,I357307,I357013);
nand I_20861 (I357341,I357259,I357324);
nand I_20862 (I356812,I357341,I357290);
nand I_20863 (I356809,I357324,I357208);
not I_20864 (I357413,I2690);
DFFARX1 I_20865 (I404566,I2683,I357413,I357439,);
and I_20866 (I357447,I357439,I404548);
DFFARX1 I_20867 (I357447,I2683,I357413,I357396,);
DFFARX1 I_20868 (I404539,I2683,I357413,I357487,);
not I_20869 (I357495,I404554);
not I_20870 (I357512,I404542);
nand I_20871 (I357529,I357512,I357495);
nor I_20872 (I357384,I357487,I357529);
DFFARX1 I_20873 (I357529,I2683,I357413,I357569,);
not I_20874 (I357405,I357569);
not I_20875 (I357591,I404551);
nand I_20876 (I357608,I357512,I357591);
DFFARX1 I_20877 (I357608,I2683,I357413,I357634,);
not I_20878 (I357642,I357634);
not I_20879 (I357659,I404560);
nand I_20880 (I357676,I357659,I404539);
and I_20881 (I357693,I357495,I357676);
nor I_20882 (I357710,I357608,I357693);
DFFARX1 I_20883 (I357710,I2683,I357413,I357381,);
DFFARX1 I_20884 (I357693,I2683,I357413,I357402,);
nor I_20885 (I357755,I404560,I404563);
nor I_20886 (I357393,I357608,I357755);
or I_20887 (I357786,I404560,I404563);
nor I_20888 (I357803,I404557,I404545);
DFFARX1 I_20889 (I357803,I2683,I357413,I357829,);
not I_20890 (I357837,I357829);
nor I_20891 (I357399,I357837,I357642);
nand I_20892 (I357868,I357837,I357487);
not I_20893 (I357885,I404557);
nand I_20894 (I357902,I357885,I357591);
nand I_20895 (I357919,I357837,I357902);
nand I_20896 (I357390,I357919,I357868);
nand I_20897 (I357387,I357902,I357786);
not I_20898 (I357991,I2690);
DFFARX1 I_20899 (I278184,I2683,I357991,I358017,);
and I_20900 (I358025,I358017,I278178);
DFFARX1 I_20901 (I358025,I2683,I357991,I357974,);
DFFARX1 I_20902 (I278196,I2683,I357991,I358065,);
not I_20903 (I358073,I278187);
not I_20904 (I358090,I278199);
nand I_20905 (I358107,I358090,I358073);
nor I_20906 (I357962,I358065,I358107);
DFFARX1 I_20907 (I358107,I2683,I357991,I358147,);
not I_20908 (I357983,I358147);
not I_20909 (I358169,I278205);
nand I_20910 (I358186,I358090,I358169);
DFFARX1 I_20911 (I358186,I2683,I357991,I358212,);
not I_20912 (I358220,I358212);
not I_20913 (I358237,I278181);
nand I_20914 (I358254,I358237,I278202);
and I_20915 (I358271,I358073,I358254);
nor I_20916 (I358288,I358186,I358271);
DFFARX1 I_20917 (I358288,I2683,I357991,I357959,);
DFFARX1 I_20918 (I358271,I2683,I357991,I357980,);
nor I_20919 (I358333,I278181,I278193);
nor I_20920 (I357971,I358186,I358333);
or I_20921 (I358364,I278181,I278193);
nor I_20922 (I358381,I278178,I278190);
DFFARX1 I_20923 (I358381,I2683,I357991,I358407,);
not I_20924 (I358415,I358407);
nor I_20925 (I357977,I358415,I358220);
nand I_20926 (I358446,I358415,I358065);
not I_20927 (I358463,I278178);
nand I_20928 (I358480,I358463,I358169);
nand I_20929 (I358497,I358415,I358480);
nand I_20930 (I357968,I358497,I358446);
nand I_20931 (I357965,I358480,I358364);
not I_20932 (I358569,I2690);
DFFARX1 I_20933 (I11992,I2683,I358569,I358595,);
and I_20934 (I358603,I358595,I11995);
DFFARX1 I_20935 (I358603,I2683,I358569,I358552,);
DFFARX1 I_20936 (I11995,I2683,I358569,I358643,);
not I_20937 (I358651,I11998);
not I_20938 (I358668,I12013);
nand I_20939 (I358685,I358668,I358651);
nor I_20940 (I358540,I358643,I358685);
DFFARX1 I_20941 (I358685,I2683,I358569,I358725,);
not I_20942 (I358561,I358725);
not I_20943 (I358747,I12007);
nand I_20944 (I358764,I358668,I358747);
DFFARX1 I_20945 (I358764,I2683,I358569,I358790,);
not I_20946 (I358798,I358790);
not I_20947 (I358815,I12010);
nand I_20948 (I358832,I358815,I11992);
and I_20949 (I358849,I358651,I358832);
nor I_20950 (I358866,I358764,I358849);
DFFARX1 I_20951 (I358866,I2683,I358569,I358537,);
DFFARX1 I_20952 (I358849,I2683,I358569,I358558,);
nor I_20953 (I358911,I12010,I12004);
nor I_20954 (I358549,I358764,I358911);
or I_20955 (I358942,I12010,I12004);
nor I_20956 (I358959,I12001,I12016);
DFFARX1 I_20957 (I358959,I2683,I358569,I358985,);
not I_20958 (I358993,I358985);
nor I_20959 (I358555,I358993,I358798);
nand I_20960 (I359024,I358993,I358643);
not I_20961 (I359041,I12001);
nand I_20962 (I359058,I359041,I358747);
nand I_20963 (I359075,I358993,I359058);
nand I_20964 (I358546,I359075,I359024);
nand I_20965 (I358543,I359058,I358942);
not I_20966 (I359147,I2690);
DFFARX1 I_20967 (I295626,I2683,I359147,I359173,);
and I_20968 (I359181,I359173,I295620);
DFFARX1 I_20969 (I359181,I2683,I359147,I359130,);
DFFARX1 I_20970 (I295638,I2683,I359147,I359221,);
not I_20971 (I359229,I295629);
not I_20972 (I359246,I295641);
nand I_20973 (I359263,I359246,I359229);
nor I_20974 (I359118,I359221,I359263);
DFFARX1 I_20975 (I359263,I2683,I359147,I359303,);
not I_20976 (I359139,I359303);
not I_20977 (I359325,I295647);
nand I_20978 (I359342,I359246,I359325);
DFFARX1 I_20979 (I359342,I2683,I359147,I359368,);
not I_20980 (I359376,I359368);
not I_20981 (I359393,I295623);
nand I_20982 (I359410,I359393,I295644);
and I_20983 (I359427,I359229,I359410);
nor I_20984 (I359444,I359342,I359427);
DFFARX1 I_20985 (I359444,I2683,I359147,I359115,);
DFFARX1 I_20986 (I359427,I2683,I359147,I359136,);
nor I_20987 (I359489,I295623,I295635);
nor I_20988 (I359127,I359342,I359489);
or I_20989 (I359520,I295623,I295635);
nor I_20990 (I359537,I295620,I295632);
DFFARX1 I_20991 (I359537,I2683,I359147,I359563,);
not I_20992 (I359571,I359563);
nor I_20993 (I359133,I359571,I359376);
nand I_20994 (I359602,I359571,I359221);
not I_20995 (I359619,I295620);
nand I_20996 (I359636,I359619,I359325);
nand I_20997 (I359653,I359571,I359636);
nand I_20998 (I359124,I359653,I359602);
nand I_20999 (I359121,I359636,I359520);
not I_21000 (I359725,I2690);
DFFARX1 I_21001 (I383653,I2683,I359725,I359751,);
and I_21002 (I359759,I359751,I383635);
DFFARX1 I_21003 (I359759,I2683,I359725,I359708,);
DFFARX1 I_21004 (I383644,I2683,I359725,I359799,);
not I_21005 (I359807,I383629);
not I_21006 (I359824,I383641);
nand I_21007 (I359841,I359824,I359807);
nor I_21008 (I359696,I359799,I359841);
DFFARX1 I_21009 (I359841,I2683,I359725,I359881,);
not I_21010 (I359717,I359881);
not I_21011 (I359903,I383632);
nand I_21012 (I359920,I359824,I359903);
DFFARX1 I_21013 (I359920,I2683,I359725,I359946,);
not I_21014 (I359954,I359946);
not I_21015 (I359971,I383629);
nand I_21016 (I359988,I359971,I383632);
and I_21017 (I360005,I359807,I359988);
nor I_21018 (I360022,I359920,I360005);
DFFARX1 I_21019 (I360022,I2683,I359725,I359693,);
DFFARX1 I_21020 (I360005,I2683,I359725,I359714,);
nor I_21021 (I360067,I383629,I383650);
nor I_21022 (I359705,I359920,I360067);
or I_21023 (I360098,I383629,I383650);
nor I_21024 (I360115,I383638,I383647);
DFFARX1 I_21025 (I360115,I2683,I359725,I360141,);
not I_21026 (I360149,I360141);
nor I_21027 (I359711,I360149,I359954);
nand I_21028 (I360180,I360149,I359799);
not I_21029 (I360197,I383638);
nand I_21030 (I360214,I360197,I359903);
nand I_21031 (I360231,I360149,I360214);
nand I_21032 (I359702,I360231,I360180);
nand I_21033 (I359699,I360214,I360098);
not I_21034 (I360303,I2690);
DFFARX1 I_21035 (I252392,I2683,I360303,I360329,);
and I_21036 (I360337,I360329,I252398);
DFFARX1 I_21037 (I360337,I2683,I360303,I360286,);
DFFARX1 I_21038 (I252404,I2683,I360303,I360377,);
not I_21039 (I360385,I252389);
not I_21040 (I360402,I252389);
nand I_21041 (I360419,I360402,I360385);
nor I_21042 (I360274,I360377,I360419);
DFFARX1 I_21043 (I360419,I2683,I360303,I360459,);
not I_21044 (I360295,I360459);
not I_21045 (I360481,I252407);
nand I_21046 (I360498,I360402,I360481);
DFFARX1 I_21047 (I360498,I2683,I360303,I360524,);
not I_21048 (I360532,I360524);
not I_21049 (I360549,I252401);
nand I_21050 (I360566,I360549,I252392);
and I_21051 (I360583,I360385,I360566);
nor I_21052 (I360600,I360498,I360583);
DFFARX1 I_21053 (I360600,I2683,I360303,I360271,);
DFFARX1 I_21054 (I360583,I2683,I360303,I360292,);
nor I_21055 (I360645,I252401,I252410);
nor I_21056 (I360283,I360498,I360645);
or I_21057 (I360676,I252401,I252410);
nor I_21058 (I360693,I252395,I252395);
DFFARX1 I_21059 (I360693,I2683,I360303,I360719,);
not I_21060 (I360727,I360719);
nor I_21061 (I360289,I360727,I360532);
nand I_21062 (I360758,I360727,I360377);
not I_21063 (I360775,I252395);
nand I_21064 (I360792,I360775,I360481);
nand I_21065 (I360809,I360727,I360792);
nand I_21066 (I360280,I360809,I360758);
nand I_21067 (I360277,I360792,I360676);
not I_21068 (I360881,I2690);
DFFARX1 I_21069 (I197290,I2683,I360881,I360907,);
and I_21070 (I360915,I360907,I197278);
DFFARX1 I_21071 (I360915,I2683,I360881,I360864,);
DFFARX1 I_21072 (I197281,I2683,I360881,I360955,);
not I_21073 (I360963,I197275);
not I_21074 (I360980,I197299);
nand I_21075 (I360997,I360980,I360963);
nor I_21076 (I360852,I360955,I360997);
DFFARX1 I_21077 (I360997,I2683,I360881,I361037,);
not I_21078 (I360873,I361037);
not I_21079 (I361059,I197287);
nand I_21080 (I361076,I360980,I361059);
DFFARX1 I_21081 (I361076,I2683,I360881,I361102,);
not I_21082 (I361110,I361102);
not I_21083 (I361127,I197296);
nand I_21084 (I361144,I361127,I197293);
and I_21085 (I361161,I360963,I361144);
nor I_21086 (I361178,I361076,I361161);
DFFARX1 I_21087 (I361178,I2683,I360881,I360849,);
DFFARX1 I_21088 (I361161,I2683,I360881,I360870,);
nor I_21089 (I361223,I197296,I197284);
nor I_21090 (I360861,I361076,I361223);
or I_21091 (I361254,I197296,I197284);
nor I_21092 (I361271,I197275,I197278);
DFFARX1 I_21093 (I361271,I2683,I360881,I361297,);
not I_21094 (I361305,I361297);
nor I_21095 (I360867,I361305,I361110);
nand I_21096 (I361336,I361305,I360955);
not I_21097 (I361353,I197275);
nand I_21098 (I361370,I361353,I361059);
nand I_21099 (I361387,I361305,I361370);
nand I_21100 (I360858,I361387,I361336);
nand I_21101 (I360855,I361370,I361254);
not I_21102 (I361459,I2690);
DFFARX1 I_21103 (I210584,I2683,I361459,I361485,);
and I_21104 (I361493,I361485,I210572);
DFFARX1 I_21105 (I361493,I2683,I361459,I361442,);
DFFARX1 I_21106 (I210575,I2683,I361459,I361533,);
not I_21107 (I361541,I210569);
not I_21108 (I361558,I210593);
nand I_21109 (I361575,I361558,I361541);
nor I_21110 (I361430,I361533,I361575);
DFFARX1 I_21111 (I361575,I2683,I361459,I361615,);
not I_21112 (I361451,I361615);
not I_21113 (I361637,I210581);
nand I_21114 (I361654,I361558,I361637);
DFFARX1 I_21115 (I361654,I2683,I361459,I361680,);
not I_21116 (I361688,I361680);
not I_21117 (I361705,I210590);
nand I_21118 (I361722,I361705,I210587);
and I_21119 (I361739,I361541,I361722);
nor I_21120 (I361756,I361654,I361739);
DFFARX1 I_21121 (I361756,I2683,I361459,I361427,);
DFFARX1 I_21122 (I361739,I2683,I361459,I361448,);
nor I_21123 (I361801,I210590,I210578);
nor I_21124 (I361439,I361654,I361801);
or I_21125 (I361832,I210590,I210578);
nor I_21126 (I361849,I210569,I210572);
DFFARX1 I_21127 (I361849,I2683,I361459,I361875,);
not I_21128 (I361883,I361875);
nor I_21129 (I361445,I361883,I361688);
nand I_21130 (I361914,I361883,I361533);
not I_21131 (I361931,I210569);
nand I_21132 (I361948,I361931,I361637);
nand I_21133 (I361965,I361883,I361948);
nand I_21134 (I361436,I361965,I361914);
nand I_21135 (I361433,I361948,I361832);
not I_21136 (I362037,I2690);
DFFARX1 I_21137 (I241852,I2683,I362037,I362063,);
and I_21138 (I362071,I362063,I241858);
DFFARX1 I_21139 (I362071,I2683,I362037,I362020,);
DFFARX1 I_21140 (I241864,I2683,I362037,I362111,);
not I_21141 (I362119,I241849);
not I_21142 (I362136,I241849);
nand I_21143 (I362153,I362136,I362119);
nor I_21144 (I362008,I362111,I362153);
DFFARX1 I_21145 (I362153,I2683,I362037,I362193,);
not I_21146 (I362029,I362193);
not I_21147 (I362215,I241867);
nand I_21148 (I362232,I362136,I362215);
DFFARX1 I_21149 (I362232,I2683,I362037,I362258,);
not I_21150 (I362266,I362258);
not I_21151 (I362283,I241861);
nand I_21152 (I362300,I362283,I241852);
and I_21153 (I362317,I362119,I362300);
nor I_21154 (I362334,I362232,I362317);
DFFARX1 I_21155 (I362334,I2683,I362037,I362005,);
DFFARX1 I_21156 (I362317,I2683,I362037,I362026,);
nor I_21157 (I362379,I241861,I241870);
nor I_21158 (I362017,I362232,I362379);
or I_21159 (I362410,I241861,I241870);
nor I_21160 (I362427,I241855,I241855);
DFFARX1 I_21161 (I362427,I2683,I362037,I362453,);
not I_21162 (I362461,I362453);
nor I_21163 (I362023,I362461,I362266);
nand I_21164 (I362492,I362461,I362111);
not I_21165 (I362509,I241855);
nand I_21166 (I362526,I362509,I362215);
nand I_21167 (I362543,I362461,I362526);
nand I_21168 (I362014,I362543,I362492);
nand I_21169 (I362011,I362526,I362410);
not I_21170 (I362615,I2690);
DFFARX1 I_21171 (I377938,I2683,I362615,I362641,);
and I_21172 (I362649,I362641,I377932);
DFFARX1 I_21173 (I362649,I2683,I362615,I362598,);
DFFARX1 I_21174 (I377917,I2683,I362615,I362689,);
not I_21175 (I362697,I377923);
not I_21176 (I362714,I377935);
nand I_21177 (I362731,I362714,I362697);
nor I_21178 (I362586,I362689,I362731);
DFFARX1 I_21179 (I362731,I2683,I362615,I362771,);
not I_21180 (I362607,I362771);
not I_21181 (I362793,I377917);
nand I_21182 (I362810,I362714,I362793);
DFFARX1 I_21183 (I362810,I2683,I362615,I362836,);
not I_21184 (I362844,I362836);
not I_21185 (I362861,I377941);
nand I_21186 (I362878,I362861,I377929);
and I_21187 (I362895,I362697,I362878);
nor I_21188 (I362912,I362810,I362895);
DFFARX1 I_21189 (I362912,I2683,I362615,I362583,);
DFFARX1 I_21190 (I362895,I2683,I362615,I362604,);
nor I_21191 (I362957,I377941,I377920);
nor I_21192 (I362595,I362810,I362957);
or I_21193 (I362988,I377941,I377920);
nor I_21194 (I363005,I377926,I377920);
DFFARX1 I_21195 (I363005,I2683,I362615,I363031,);
not I_21196 (I363039,I363031);
nor I_21197 (I362601,I363039,I362844);
nand I_21198 (I363070,I363039,I362689);
not I_21199 (I363087,I377926);
nand I_21200 (I363104,I363087,I362793);
nand I_21201 (I363121,I363039,I363104);
nand I_21202 (I362592,I363121,I363070);
nand I_21203 (I362589,I363104,I362988);
not I_21204 (I363193,I2690);
DFFARX1 I_21205 (I401591,I2683,I363193,I363219,);
and I_21206 (I363227,I363219,I401573);
DFFARX1 I_21207 (I363227,I2683,I363193,I363176,);
DFFARX1 I_21208 (I401564,I2683,I363193,I363267,);
not I_21209 (I363275,I401579);
not I_21210 (I363292,I401567);
nand I_21211 (I363309,I363292,I363275);
nor I_21212 (I363164,I363267,I363309);
DFFARX1 I_21213 (I363309,I2683,I363193,I363349,);
not I_21214 (I363185,I363349);
not I_21215 (I363371,I401576);
nand I_21216 (I363388,I363292,I363371);
DFFARX1 I_21217 (I363388,I2683,I363193,I363414,);
not I_21218 (I363422,I363414);
not I_21219 (I363439,I401585);
nand I_21220 (I363456,I363439,I401564);
and I_21221 (I363473,I363275,I363456);
nor I_21222 (I363490,I363388,I363473);
DFFARX1 I_21223 (I363490,I2683,I363193,I363161,);
DFFARX1 I_21224 (I363473,I2683,I363193,I363182,);
nor I_21225 (I363535,I401585,I401588);
nor I_21226 (I363173,I363388,I363535);
or I_21227 (I363566,I401585,I401588);
nor I_21228 (I363583,I401582,I401570);
DFFARX1 I_21229 (I363583,I2683,I363193,I363609,);
not I_21230 (I363617,I363609);
nor I_21231 (I363179,I363617,I363422);
nand I_21232 (I363648,I363617,I363267);
not I_21233 (I363665,I401582);
nand I_21234 (I363682,I363665,I363371);
nand I_21235 (I363699,I363617,I363682);
nand I_21236 (I363170,I363699,I363648);
nand I_21237 (I363167,I363682,I363566);
not I_21238 (I363771,I2690);
DFFARX1 I_21239 (I309835,I2683,I363771,I363797,);
and I_21240 (I363805,I363797,I309832);
DFFARX1 I_21241 (I363805,I2683,I363771,I363754,);
DFFARX1 I_21242 (I309838,I2683,I363771,I363845,);
not I_21243 (I363853,I309841);
not I_21244 (I363870,I309835);
nand I_21245 (I363887,I363870,I363853);
nor I_21246 (I363742,I363845,I363887);
DFFARX1 I_21247 (I363887,I2683,I363771,I363927,);
not I_21248 (I363763,I363927);
not I_21249 (I363949,I309850);
nand I_21250 (I363966,I363870,I363949);
DFFARX1 I_21251 (I363966,I2683,I363771,I363992,);
not I_21252 (I364000,I363992);
not I_21253 (I364017,I309847);
nand I_21254 (I364034,I364017,I309853);
and I_21255 (I364051,I363853,I364034);
nor I_21256 (I364068,I363966,I364051);
DFFARX1 I_21257 (I364068,I2683,I363771,I363739,);
DFFARX1 I_21258 (I364051,I2683,I363771,I363760,);
nor I_21259 (I364113,I309847,I309832);
nor I_21260 (I363751,I363966,I364113);
or I_21261 (I364144,I309847,I309832);
nor I_21262 (I364161,I309844,I309838);
DFFARX1 I_21263 (I364161,I2683,I363771,I364187,);
not I_21264 (I364195,I364187);
nor I_21265 (I363757,I364195,I364000);
nand I_21266 (I364226,I364195,I363845);
not I_21267 (I364243,I309844);
nand I_21268 (I364260,I364243,I363949);
nand I_21269 (I364277,I364195,I364260);
nand I_21270 (I363748,I364277,I364226);
nand I_21271 (I363745,I364260,I364144);
not I_21272 (I364349,I2690);
DFFARX1 I_21273 (I215774,I2683,I364349,I364375,);
nand I_21274 (I364383,I364375,I215789);
DFFARX1 I_21275 (I215783,I2683,I364349,I364409,);
DFFARX1 I_21276 (I364409,I2683,I364349,I364426,);
not I_21277 (I364341,I364426);
not I_21278 (I364448,I215786);
nor I_21279 (I364465,I215786,I215792);
not I_21280 (I364482,I215774);
nand I_21281 (I364499,I364448,I364482);
nor I_21282 (I364516,I215774,I215786);
and I_21283 (I364320,I364516,I364383);
not I_21284 (I364547,I215771);
nand I_21285 (I364564,I364547,I215777);
nor I_21286 (I364581,I215771,I215771);
not I_21287 (I364598,I364581);
nand I_21288 (I364323,I364465,I364598);
DFFARX1 I_21289 (I364581,I2683,I364349,I364338,);
nor I_21290 (I364643,I215780,I215774);
nor I_21291 (I364660,I364643,I215792);
and I_21292 (I364677,I364660,I364564);
DFFARX1 I_21293 (I364677,I2683,I364349,I364335,);
nor I_21294 (I364332,I364643,I364499);
or I_21295 (I364329,I364581,I364643);
nor I_21296 (I364736,I215780,I215795);
DFFARX1 I_21297 (I364736,I2683,I364349,I364762,);
not I_21298 (I364770,I364762);
nand I_21299 (I364787,I364770,I364448);
nor I_21300 (I364804,I364787,I215792);
DFFARX1 I_21301 (I364804,I2683,I364349,I364317,);
nor I_21302 (I364835,I364770,I364499);
nor I_21303 (I364326,I364643,I364835);
not I_21304 (I364893,I2690);
DFFARX1 I_21305 (I317143,I2683,I364893,I364919,);
nand I_21306 (I364927,I364919,I317131);
DFFARX1 I_21307 (I317125,I2683,I364893,I364953,);
DFFARX1 I_21308 (I364953,I2683,I364893,I364970,);
not I_21309 (I364885,I364970);
not I_21310 (I364992,I317125);
nor I_21311 (I365009,I317125,I317137);
not I_21312 (I365026,I317134);
nand I_21313 (I365043,I364992,I365026);
nor I_21314 (I365060,I317134,I317125);
and I_21315 (I364864,I365060,I364927);
not I_21316 (I365091,I317128);
nand I_21317 (I365108,I365091,I317140);
nor I_21318 (I365125,I317128,I317146);
not I_21319 (I365142,I365125);
nand I_21320 (I364867,I365009,I365142);
DFFARX1 I_21321 (I365125,I2683,I364893,I364882,);
nor I_21322 (I365187,I317131,I317134);
nor I_21323 (I365204,I365187,I317137);
and I_21324 (I365221,I365204,I365108);
DFFARX1 I_21325 (I365221,I2683,I364893,I364879,);
nor I_21326 (I364876,I365187,I365043);
or I_21327 (I364873,I365125,I365187);
nor I_21328 (I365280,I317131,I317128);
DFFARX1 I_21329 (I365280,I2683,I364893,I365306,);
not I_21330 (I365314,I365306);
nand I_21331 (I365331,I365314,I364992);
nor I_21332 (I365348,I365331,I317137);
DFFARX1 I_21333 (I365348,I2683,I364893,I364861,);
nor I_21334 (I365379,I365314,I365043);
nor I_21335 (I364870,I365187,I365379);
not I_21336 (I365437,I2690);
DFFARX1 I_21337 (I271718,I2683,I365437,I365463,);
nand I_21338 (I365471,I365463,I271718);
DFFARX1 I_21339 (I271730,I2683,I365437,I365497,);
DFFARX1 I_21340 (I365497,I2683,I365437,I365514,);
not I_21341 (I365429,I365514);
not I_21342 (I365536,I271724);
nor I_21343 (I365553,I271724,I271745);
not I_21344 (I365570,I271733);
nand I_21345 (I365587,I365536,I365570);
nor I_21346 (I365604,I271733,I271724);
and I_21347 (I365408,I365604,I365471);
not I_21348 (I365635,I271727);
nand I_21349 (I365652,I365635,I271742);
nor I_21350 (I365669,I271727,I271736);
not I_21351 (I365686,I365669);
nand I_21352 (I365411,I365553,I365686);
DFFARX1 I_21353 (I365669,I2683,I365437,I365426,);
nor I_21354 (I365731,I271739,I271733);
nor I_21355 (I365748,I365731,I271745);
and I_21356 (I365765,I365748,I365652);
DFFARX1 I_21357 (I365765,I2683,I365437,I365423,);
nor I_21358 (I365420,I365731,I365587);
or I_21359 (I365417,I365669,I365731);
nor I_21360 (I365824,I271739,I271721);
DFFARX1 I_21361 (I365824,I2683,I365437,I365850,);
not I_21362 (I365858,I365850);
nand I_21363 (I365875,I365858,I365536);
nor I_21364 (I365892,I365875,I271745);
DFFARX1 I_21365 (I365892,I2683,I365437,I365405,);
nor I_21366 (I365923,I365858,I365587);
nor I_21367 (I365414,I365731,I365923);
not I_21368 (I365981,I2690);
DFFARX1 I_21369 (I67353,I2683,I365981,I366007,);
nand I_21370 (I366015,I366007,I67368);
DFFARX1 I_21371 (I67365,I2683,I365981,I366041,);
DFFARX1 I_21372 (I366041,I2683,I365981,I366058,);
not I_21373 (I365973,I366058);
not I_21374 (I366080,I67344);
nor I_21375 (I366097,I67344,I67350);
not I_21376 (I366114,I67356);
nand I_21377 (I366131,I366080,I366114);
nor I_21378 (I366148,I67356,I67344);
and I_21379 (I365952,I366148,I366015);
not I_21380 (I366179,I67362);
nand I_21381 (I366196,I366179,I67344);
nor I_21382 (I366213,I67362,I67347);
not I_21383 (I366230,I366213);
nand I_21384 (I365955,I366097,I366230);
DFFARX1 I_21385 (I366213,I2683,I365981,I365970,);
nor I_21386 (I366275,I67347,I67356);
nor I_21387 (I366292,I366275,I67350);
and I_21388 (I366309,I366292,I366196);
DFFARX1 I_21389 (I366309,I2683,I365981,I365967,);
nor I_21390 (I365964,I366275,I366131);
or I_21391 (I365961,I366213,I366275);
nor I_21392 (I366368,I67347,I67359);
DFFARX1 I_21393 (I366368,I2683,I365981,I366394,);
not I_21394 (I366402,I366394);
nand I_21395 (I366419,I366402,I366080);
nor I_21396 (I366436,I366419,I67350);
DFFARX1 I_21397 (I366436,I2683,I365981,I365949,);
nor I_21398 (I366467,I366402,I366131);
nor I_21399 (I365958,I366275,I366467);
not I_21400 (I366525,I2690);
DFFARX1 I_21401 (I94233,I2683,I366525,I366551,);
nand I_21402 (I366559,I366551,I94236);
DFFARX1 I_21403 (I94230,I2683,I366525,I366585,);
DFFARX1 I_21404 (I366585,I2683,I366525,I366602,);
not I_21405 (I366517,I366602);
not I_21406 (I366624,I94239);
nor I_21407 (I366641,I94239,I94224);
not I_21408 (I366658,I94248);
nand I_21409 (I366675,I366624,I366658);
nor I_21410 (I366692,I94248,I94239);
and I_21411 (I366496,I366692,I366559);
not I_21412 (I366723,I94227);
nand I_21413 (I366740,I366723,I94245);
nor I_21414 (I366757,I94227,I94221);
not I_21415 (I366774,I366757);
nand I_21416 (I366499,I366641,I366774);
DFFARX1 I_21417 (I366757,I2683,I366525,I366514,);
nor I_21418 (I366819,I94242,I94248);
nor I_21419 (I366836,I366819,I94224);
and I_21420 (I366853,I366836,I366740);
DFFARX1 I_21421 (I366853,I2683,I366525,I366511,);
nor I_21422 (I366508,I366819,I366675);
or I_21423 (I366505,I366757,I366819);
nor I_21424 (I366912,I94242,I94221);
DFFARX1 I_21425 (I366912,I2683,I366525,I366938,);
not I_21426 (I366946,I366938);
nand I_21427 (I366963,I366946,I366624);
nor I_21428 (I366980,I366963,I94224);
DFFARX1 I_21429 (I366980,I2683,I366525,I366493,);
nor I_21430 (I367011,I366946,I366675);
nor I_21431 (I366502,I366819,I367011);
not I_21432 (I367069,I2690);
DFFARX1 I_21433 (I219820,I2683,I367069,I367095,);
nand I_21434 (I367103,I367095,I219835);
DFFARX1 I_21435 (I219829,I2683,I367069,I367129,);
DFFARX1 I_21436 (I367129,I2683,I367069,I367146,);
not I_21437 (I367061,I367146);
not I_21438 (I367168,I219832);
nor I_21439 (I367185,I219832,I219838);
not I_21440 (I367202,I219820);
nand I_21441 (I367219,I367168,I367202);
nor I_21442 (I367236,I219820,I219832);
and I_21443 (I367040,I367236,I367103);
not I_21444 (I367267,I219817);
nand I_21445 (I367284,I367267,I219823);
nor I_21446 (I367301,I219817,I219817);
not I_21447 (I367318,I367301);
nand I_21448 (I367043,I367185,I367318);
DFFARX1 I_21449 (I367301,I2683,I367069,I367058,);
nor I_21450 (I367363,I219826,I219820);
nor I_21451 (I367380,I367363,I219838);
and I_21452 (I367397,I367380,I367284);
DFFARX1 I_21453 (I367397,I2683,I367069,I367055,);
nor I_21454 (I367052,I367363,I367219);
or I_21455 (I367049,I367301,I367363);
nor I_21456 (I367456,I219826,I219841);
DFFARX1 I_21457 (I367456,I2683,I367069,I367482,);
not I_21458 (I367490,I367482);
nand I_21459 (I367507,I367490,I367168);
nor I_21460 (I367524,I367507,I219838);
DFFARX1 I_21461 (I367524,I2683,I367069,I367037,);
nor I_21462 (I367555,I367490,I367219);
nor I_21463 (I367046,I367363,I367555);
not I_21464 (I367613,I2690);
DFFARX1 I_21465 (I247125,I2683,I367613,I367639,);
nand I_21466 (I367647,I367639,I247119);
DFFARX1 I_21467 (I247122,I2683,I367613,I367673,);
DFFARX1 I_21468 (I367673,I2683,I367613,I367690,);
not I_21469 (I367605,I367690);
not I_21470 (I367712,I247128);
nor I_21471 (I367729,I247128,I247122);
not I_21472 (I367746,I247131);
nand I_21473 (I367763,I367712,I367746);
nor I_21474 (I367780,I247131,I247128);
and I_21475 (I367584,I367780,I367647);
not I_21476 (I367811,I247140);
nand I_21477 (I367828,I367811,I247134);
nor I_21478 (I367845,I247140,I247137);
not I_21479 (I367862,I367845);
nand I_21480 (I367587,I367729,I367862);
DFFARX1 I_21481 (I367845,I2683,I367613,I367602,);
nor I_21482 (I367907,I247119,I247131);
nor I_21483 (I367924,I367907,I247122);
and I_21484 (I367941,I367924,I367828);
DFFARX1 I_21485 (I367941,I2683,I367613,I367599,);
nor I_21486 (I367596,I367907,I367763);
or I_21487 (I367593,I367845,I367907);
nor I_21488 (I368000,I247119,I247125);
DFFARX1 I_21489 (I368000,I2683,I367613,I368026,);
not I_21490 (I368034,I368026);
nand I_21491 (I368051,I368034,I367712);
nor I_21492 (I368068,I368051,I247122);
DFFARX1 I_21493 (I368068,I2683,I367613,I367581,);
nor I_21494 (I368099,I368034,I367763);
nor I_21495 (I367590,I367907,I368099);
not I_21496 (I368157,I2690);
DFFARX1 I_21497 (I7785,I2683,I368157,I368183,);
nand I_21498 (I368191,I368183,I7779);
DFFARX1 I_21499 (I7800,I2683,I368157,I368217,);
DFFARX1 I_21500 (I368217,I2683,I368157,I368234,);
not I_21501 (I368149,I368234);
not I_21502 (I368256,I7788);
nor I_21503 (I368273,I7788,I7797);
not I_21504 (I368290,I7776);
nand I_21505 (I368307,I368256,I368290);
nor I_21506 (I368324,I7776,I7788);
and I_21507 (I368128,I368324,I368191);
not I_21508 (I368355,I7794);
nand I_21509 (I368372,I368355,I7782);
nor I_21510 (I368389,I7794,I7776);
not I_21511 (I368406,I368389);
nand I_21512 (I368131,I368273,I368406);
DFFARX1 I_21513 (I368389,I2683,I368157,I368146,);
nor I_21514 (I368451,I7779,I7776);
nor I_21515 (I368468,I368451,I7797);
and I_21516 (I368485,I368468,I368372);
DFFARX1 I_21517 (I368485,I2683,I368157,I368143,);
nor I_21518 (I368140,I368451,I368307);
or I_21519 (I368137,I368389,I368451);
nor I_21520 (I368544,I7779,I7791);
DFFARX1 I_21521 (I368544,I2683,I368157,I368570,);
not I_21522 (I368578,I368570);
nand I_21523 (I368595,I368578,I368256);
nor I_21524 (I368612,I368595,I7797);
DFFARX1 I_21525 (I368612,I2683,I368157,I368125,);
nor I_21526 (I368643,I368578,I368307);
nor I_21527 (I368134,I368451,I368643);
not I_21528 (I368701,I2690);
DFFARX1 I_21529 (I344111,I2683,I368701,I368727,);
nand I_21530 (I368735,I368727,I344090);
DFFARX1 I_21531 (I344087,I2683,I368701,I368761,);
DFFARX1 I_21532 (I368761,I2683,I368701,I368778,);
not I_21533 (I368693,I368778);
not I_21534 (I368800,I344099);
nor I_21535 (I368817,I344099,I344108);
not I_21536 (I368834,I344096);
nand I_21537 (I368851,I368800,I368834);
nor I_21538 (I368868,I344096,I344099);
and I_21539 (I368672,I368868,I368735);
not I_21540 (I368899,I344105);
nand I_21541 (I368916,I368899,I344102);
nor I_21542 (I368933,I344105,I344087);
not I_21543 (I368950,I368933);
nand I_21544 (I368675,I368817,I368950);
DFFARX1 I_21545 (I368933,I2683,I368701,I368690,);
nor I_21546 (I368995,I344090,I344096);
nor I_21547 (I369012,I368995,I344108);
and I_21548 (I369029,I369012,I368916);
DFFARX1 I_21549 (I369029,I2683,I368701,I368687,);
nor I_21550 (I368684,I368995,I368851);
or I_21551 (I368681,I368933,I368995);
nor I_21552 (I369088,I344090,I344093);
DFFARX1 I_21553 (I369088,I2683,I368701,I369114,);
not I_21554 (I369122,I369114);
nand I_21555 (I369139,I369122,I368800);
nor I_21556 (I369156,I369139,I344108);
DFFARX1 I_21557 (I369156,I2683,I368701,I368669,);
nor I_21558 (I369187,I369122,I368851);
nor I_21559 (I368678,I368995,I369187);
not I_21560 (I369245,I2690);
DFFARX1 I_21561 (I46546,I2683,I369245,I369271,);
nand I_21562 (I369279,I369271,I46519);
DFFARX1 I_21563 (I46537,I2683,I369245,I369305,);
DFFARX1 I_21564 (I369305,I2683,I369245,I369322,);
not I_21565 (I369237,I369322);
not I_21566 (I369344,I46531);
nor I_21567 (I369361,I46531,I46519);
not I_21568 (I369378,I46534);
nand I_21569 (I369395,I369344,I369378);
nor I_21570 (I369412,I46534,I46531);
and I_21571 (I369216,I369412,I369279);
not I_21572 (I369443,I46522);
nand I_21573 (I369460,I369443,I46540);
nor I_21574 (I369477,I46522,I46543);
not I_21575 (I369494,I369477);
nand I_21576 (I369219,I369361,I369494);
DFFARX1 I_21577 (I369477,I2683,I369245,I369234,);
nor I_21578 (I369539,I46525,I46534);
nor I_21579 (I369556,I369539,I46519);
and I_21580 (I369573,I369556,I369460);
DFFARX1 I_21581 (I369573,I2683,I369245,I369231,);
nor I_21582 (I369228,I369539,I369395);
or I_21583 (I369225,I369477,I369539);
nor I_21584 (I369632,I46525,I46528);
DFFARX1 I_21585 (I369632,I2683,I369245,I369658,);
not I_21586 (I369666,I369658);
nand I_21587 (I369683,I369666,I369344);
nor I_21588 (I369700,I369683,I46519);
DFFARX1 I_21589 (I369700,I2683,I369245,I369213,);
nor I_21590 (I369731,I369666,I369395);
nor I_21591 (I369222,I369539,I369731);
not I_21592 (I369789,I2690);
DFFARX1 I_21593 (I194388,I2683,I369789,I369815,);
nand I_21594 (I369823,I369815,I194403);
DFFARX1 I_21595 (I194397,I2683,I369789,I369849,);
DFFARX1 I_21596 (I369849,I2683,I369789,I369866,);
not I_21597 (I369781,I369866);
not I_21598 (I369888,I194400);
nor I_21599 (I369905,I194400,I194406);
not I_21600 (I369922,I194388);
nand I_21601 (I369939,I369888,I369922);
nor I_21602 (I369956,I194388,I194400);
and I_21603 (I369760,I369956,I369823);
not I_21604 (I369987,I194385);
nand I_21605 (I370004,I369987,I194391);
nor I_21606 (I370021,I194385,I194385);
not I_21607 (I370038,I370021);
nand I_21608 (I369763,I369905,I370038);
DFFARX1 I_21609 (I370021,I2683,I369789,I369778,);
nor I_21610 (I370083,I194394,I194388);
nor I_21611 (I370100,I370083,I194406);
and I_21612 (I370117,I370100,I370004);
DFFARX1 I_21613 (I370117,I2683,I369789,I369775,);
nor I_21614 (I369772,I370083,I369939);
or I_21615 (I369769,I370021,I370083);
nor I_21616 (I370176,I194394,I194409);
DFFARX1 I_21617 (I370176,I2683,I369789,I370202,);
not I_21618 (I370210,I370202);
nand I_21619 (I370227,I370210,I369888);
nor I_21620 (I370244,I370227,I194406);
DFFARX1 I_21621 (I370244,I2683,I369789,I369757,);
nor I_21622 (I370275,I370210,I369939);
nor I_21623 (I369766,I370083,I370275);
not I_21624 (I370333,I2690);
DFFARX1 I_21625 (I154119,I2683,I370333,I370359,);
nand I_21626 (I370367,I370359,I154116);
DFFARX1 I_21627 (I154095,I2683,I370333,I370393,);
DFFARX1 I_21628 (I370393,I2683,I370333,I370410,);
not I_21629 (I370325,I370410);
not I_21630 (I370432,I154110);
nor I_21631 (I370449,I154110,I154113);
not I_21632 (I370466,I154104);
nand I_21633 (I370483,I370432,I370466);
nor I_21634 (I370500,I154104,I154110);
and I_21635 (I370304,I370500,I370367);
not I_21636 (I370531,I154101);
nand I_21637 (I370548,I370531,I154122);
nor I_21638 (I370565,I154101,I154098);
not I_21639 (I370582,I370565);
nand I_21640 (I370307,I370449,I370582);
DFFARX1 I_21641 (I370565,I2683,I370333,I370322,);
nor I_21642 (I370627,I154107,I154104);
nor I_21643 (I370644,I370627,I154113);
and I_21644 (I370661,I370644,I370548);
DFFARX1 I_21645 (I370661,I2683,I370333,I370319,);
nor I_21646 (I370316,I370627,I370483);
or I_21647 (I370313,I370565,I370627);
nor I_21648 (I370720,I154107,I154095);
DFFARX1 I_21649 (I370720,I2683,I370333,I370746,);
not I_21650 (I370754,I370746);
nand I_21651 (I370771,I370754,I370432);
nor I_21652 (I370788,I370771,I154113);
DFFARX1 I_21653 (I370788,I2683,I370333,I370301,);
nor I_21654 (I370819,I370754,I370483);
nor I_21655 (I370310,I370627,I370819);
not I_21656 (I370877,I2690);
DFFARX1 I_21657 (I180534,I2683,I370877,I370903,);
nand I_21658 (I370911,I370903,I180522);
DFFARX1 I_21659 (I180528,I2683,I370877,I370937,);
DFFARX1 I_21660 (I370937,I2683,I370877,I370954,);
not I_21661 (I370869,I370954);
not I_21662 (I370976,I180513);
nor I_21663 (I370993,I180513,I180525);
not I_21664 (I371010,I180516);
nand I_21665 (I371027,I370976,I371010);
nor I_21666 (I371044,I180516,I180513);
and I_21667 (I370848,I371044,I370911);
not I_21668 (I371075,I180531);
nand I_21669 (I371092,I371075,I180513);
nor I_21670 (I371109,I180531,I180537);
not I_21671 (I371126,I371109);
nand I_21672 (I370851,I370993,I371126);
DFFARX1 I_21673 (I371109,I2683,I370877,I370866,);
nor I_21674 (I371171,I180519,I180516);
nor I_21675 (I371188,I371171,I180525);
and I_21676 (I371205,I371188,I371092);
DFFARX1 I_21677 (I371205,I2683,I370877,I370863,);
nor I_21678 (I370860,I371171,I371027);
or I_21679 (I370857,I371109,I371171);
nor I_21680 (I371264,I180519,I180516);
DFFARX1 I_21681 (I371264,I2683,I370877,I371290,);
not I_21682 (I371298,I371290);
nand I_21683 (I371315,I371298,I370976);
nor I_21684 (I371332,I371315,I180525);
DFFARX1 I_21685 (I371332,I2683,I370877,I370845,);
nor I_21686 (I371363,I371298,I371027);
nor I_21687 (I370854,I371171,I371363);
not I_21688 (I371421,I2690);
DFFARX1 I_21689 (I25188,I2683,I371421,I371447,);
nand I_21690 (I371455,I371447,I25170);
DFFARX1 I_21691 (I25167,I2683,I371421,I371481,);
DFFARX1 I_21692 (I371481,I2683,I371421,I371498,);
not I_21693 (I371413,I371498);
not I_21694 (I371520,I25185);
nor I_21695 (I371537,I25185,I25179);
not I_21696 (I371554,I25167);
nand I_21697 (I371571,I371520,I371554);
nor I_21698 (I371588,I25167,I25185);
and I_21699 (I371392,I371588,I371455);
not I_21700 (I371619,I25176);
nand I_21701 (I371636,I371619,I25182);
nor I_21702 (I371653,I25176,I25170);
not I_21703 (I371670,I371653);
nand I_21704 (I371395,I371537,I371670);
DFFARX1 I_21705 (I371653,I2683,I371421,I371410,);
nor I_21706 (I371715,I25173,I25167);
nor I_21707 (I371732,I371715,I25179);
and I_21708 (I371749,I371732,I371636);
DFFARX1 I_21709 (I371749,I2683,I371421,I371407,);
nor I_21710 (I371404,I371715,I371571);
or I_21711 (I371401,I371653,I371715);
nor I_21712 (I371808,I25173,I25191);
DFFARX1 I_21713 (I371808,I2683,I371421,I371834,);
not I_21714 (I371842,I371834);
nand I_21715 (I371859,I371842,I371520);
nor I_21716 (I371876,I371859,I25179);
DFFARX1 I_21717 (I371876,I2683,I371421,I371389,);
nor I_21718 (I371907,I371842,I371571);
nor I_21719 (I371398,I371715,I371907);
not I_21720 (I371965,I2690);
DFFARX1 I_21721 (I89490,I2683,I371965,I371991,);
nand I_21722 (I371999,I371991,I89493);
DFFARX1 I_21723 (I89487,I2683,I371965,I372025,);
DFFARX1 I_21724 (I372025,I2683,I371965,I372042,);
not I_21725 (I371957,I372042);
not I_21726 (I372064,I89496);
nor I_21727 (I372081,I89496,I89481);
not I_21728 (I372098,I89505);
nand I_21729 (I372115,I372064,I372098);
nor I_21730 (I372132,I89505,I89496);
and I_21731 (I371936,I372132,I371999);
not I_21732 (I372163,I89484);
nand I_21733 (I372180,I372163,I89502);
nor I_21734 (I372197,I89484,I89478);
not I_21735 (I372214,I372197);
nand I_21736 (I371939,I372081,I372214);
DFFARX1 I_21737 (I372197,I2683,I371965,I371954,);
nor I_21738 (I372259,I89499,I89505);
nor I_21739 (I372276,I372259,I89481);
and I_21740 (I372293,I372276,I372180);
DFFARX1 I_21741 (I372293,I2683,I371965,I371951,);
nor I_21742 (I371948,I372259,I372115);
or I_21743 (I371945,I372197,I372259);
nor I_21744 (I372352,I89499,I89478);
DFFARX1 I_21745 (I372352,I2683,I371965,I372378,);
not I_21746 (I372386,I372378);
nand I_21747 (I372403,I372386,I372064);
nor I_21748 (I372420,I372403,I89481);
DFFARX1 I_21749 (I372420,I2683,I371965,I371933,);
nor I_21750 (I372451,I372386,I372115);
nor I_21751 (I371942,I372259,I372451);
not I_21752 (I372509,I2690);
DFFARX1 I_21753 (I167134,I2683,I372509,I372535,);
nand I_21754 (I372543,I372535,I167158);
DFFARX1 I_21755 (I167137,I2683,I372509,I372569,);
DFFARX1 I_21756 (I372569,I2683,I372509,I372586,);
not I_21757 (I372501,I372586);
not I_21758 (I372608,I167140);
nor I_21759 (I372625,I167140,I167155);
not I_21760 (I372642,I167146);
nand I_21761 (I372659,I372608,I372642);
nor I_21762 (I372676,I167146,I167140);
and I_21763 (I372480,I372676,I372543);
not I_21764 (I372707,I167143);
nand I_21765 (I372724,I372707,I167137);
nor I_21766 (I372741,I167143,I167152);
not I_21767 (I372758,I372741);
nand I_21768 (I372483,I372625,I372758);
DFFARX1 I_21769 (I372741,I2683,I372509,I372498,);
nor I_21770 (I372803,I167149,I167146);
nor I_21771 (I372820,I372803,I167155);
and I_21772 (I372837,I372820,I372724);
DFFARX1 I_21773 (I372837,I2683,I372509,I372495,);
nor I_21774 (I372492,I372803,I372659);
or I_21775 (I372489,I372741,I372803);
nor I_21776 (I372896,I167149,I167134);
DFFARX1 I_21777 (I372896,I2683,I372509,I372922,);
not I_21778 (I372930,I372922);
nand I_21779 (I372947,I372930,I372608);
nor I_21780 (I372964,I372947,I167155);
DFFARX1 I_21781 (I372964,I2683,I372509,I372477,);
nor I_21782 (I372995,I372930,I372659);
nor I_21783 (I372486,I372803,I372995);
not I_21784 (I373053,I2690);
DFFARX1 I_21785 (I326193,I2683,I373053,I373079,);
nand I_21786 (I373087,I373079,I326172);
DFFARX1 I_21787 (I326169,I2683,I373053,I373113,);
DFFARX1 I_21788 (I373113,I2683,I373053,I373130,);
not I_21789 (I373045,I373130);
not I_21790 (I373152,I326181);
nor I_21791 (I373169,I326181,I326190);
not I_21792 (I373186,I326178);
nand I_21793 (I373203,I373152,I373186);
nor I_21794 (I373220,I326178,I326181);
and I_21795 (I373024,I373220,I373087);
not I_21796 (I373251,I326187);
nand I_21797 (I373268,I373251,I326184);
nor I_21798 (I373285,I326187,I326169);
not I_21799 (I373302,I373285);
nand I_21800 (I373027,I373169,I373302);
DFFARX1 I_21801 (I373285,I2683,I373053,I373042,);
nor I_21802 (I373347,I326172,I326178);
nor I_21803 (I373364,I373347,I326190);
and I_21804 (I373381,I373364,I373268);
DFFARX1 I_21805 (I373381,I2683,I373053,I373039,);
nor I_21806 (I373036,I373347,I373203);
or I_21807 (I373033,I373285,I373347);
nor I_21808 (I373440,I326172,I326175);
DFFARX1 I_21809 (I373440,I2683,I373053,I373466,);
not I_21810 (I373474,I373466);
nand I_21811 (I373491,I373474,I373152);
nor I_21812 (I373508,I373491,I326190);
DFFARX1 I_21813 (I373508,I2683,I373053,I373021,);
nor I_21814 (I373539,I373474,I373203);
nor I_21815 (I373030,I373347,I373539);
not I_21816 (I373597,I2690);
DFFARX1 I_21817 (I57833,I2683,I373597,I373623,);
nand I_21818 (I373631,I373623,I57848);
DFFARX1 I_21819 (I57845,I2683,I373597,I373657,);
DFFARX1 I_21820 (I373657,I2683,I373597,I373674,);
not I_21821 (I373589,I373674);
not I_21822 (I373696,I57824);
nor I_21823 (I373713,I57824,I57830);
not I_21824 (I373730,I57836);
nand I_21825 (I373747,I373696,I373730);
nor I_21826 (I373764,I57836,I57824);
and I_21827 (I373568,I373764,I373631);
not I_21828 (I373795,I57842);
nand I_21829 (I373812,I373795,I57824);
nor I_21830 (I373829,I57842,I57827);
not I_21831 (I373846,I373829);
nand I_21832 (I373571,I373713,I373846);
DFFARX1 I_21833 (I373829,I2683,I373597,I373586,);
nor I_21834 (I373891,I57827,I57836);
nor I_21835 (I373908,I373891,I57830);
and I_21836 (I373925,I373908,I373812);
DFFARX1 I_21837 (I373925,I2683,I373597,I373583,);
nor I_21838 (I373580,I373891,I373747);
or I_21839 (I373577,I373829,I373891);
nor I_21840 (I373984,I57827,I57839);
DFFARX1 I_21841 (I373984,I2683,I373597,I374010,);
not I_21842 (I374018,I374010);
nand I_21843 (I374035,I374018,I373696);
nor I_21844 (I374052,I374035,I57830);
DFFARX1 I_21845 (I374052,I2683,I373597,I373565,);
nor I_21846 (I374083,I374018,I373747);
nor I_21847 (I373574,I373891,I374083);
not I_21848 (I374141,I2690);
DFFARX1 I_21849 (I214040,I2683,I374141,I374167,);
nand I_21850 (I374175,I374167,I214055);
DFFARX1 I_21851 (I214049,I2683,I374141,I374201,);
DFFARX1 I_21852 (I374201,I2683,I374141,I374218,);
not I_21853 (I374133,I374218);
not I_21854 (I374240,I214052);
nor I_21855 (I374257,I214052,I214058);
not I_21856 (I374274,I214040);
nand I_21857 (I374291,I374240,I374274);
nor I_21858 (I374308,I214040,I214052);
and I_21859 (I374112,I374308,I374175);
not I_21860 (I374339,I214037);
nand I_21861 (I374356,I374339,I214043);
nor I_21862 (I374373,I214037,I214037);
not I_21863 (I374390,I374373);
nand I_21864 (I374115,I374257,I374390);
DFFARX1 I_21865 (I374373,I2683,I374141,I374130,);
nor I_21866 (I374435,I214046,I214040);
nor I_21867 (I374452,I374435,I214058);
and I_21868 (I374469,I374452,I374356);
DFFARX1 I_21869 (I374469,I2683,I374141,I374127,);
nor I_21870 (I374124,I374435,I374291);
or I_21871 (I374121,I374373,I374435);
nor I_21872 (I374528,I214046,I214061);
DFFARX1 I_21873 (I374528,I2683,I374141,I374554,);
not I_21874 (I374562,I374554);
nand I_21875 (I374579,I374562,I374240);
nor I_21876 (I374596,I374579,I214058);
DFFARX1 I_21877 (I374596,I2683,I374141,I374109,);
nor I_21878 (I374627,I374562,I374291);
nor I_21879 (I374118,I374435,I374627);
not I_21880 (I374685,I2690);
DFFARX1 I_21881 (I331973,I2683,I374685,I374711,);
nand I_21882 (I374719,I374711,I331952);
DFFARX1 I_21883 (I331949,I2683,I374685,I374745,);
DFFARX1 I_21884 (I374745,I2683,I374685,I374762,);
not I_21885 (I374677,I374762);
not I_21886 (I374784,I331961);
nor I_21887 (I374801,I331961,I331970);
not I_21888 (I374818,I331958);
nand I_21889 (I374835,I374784,I374818);
nor I_21890 (I374852,I331958,I331961);
and I_21891 (I374656,I374852,I374719);
not I_21892 (I374883,I331967);
nand I_21893 (I374900,I374883,I331964);
nor I_21894 (I374917,I331967,I331949);
not I_21895 (I374934,I374917);
nand I_21896 (I374659,I374801,I374934);
DFFARX1 I_21897 (I374917,I2683,I374685,I374674,);
nor I_21898 (I374979,I331952,I331958);
nor I_21899 (I374996,I374979,I331970);
and I_21900 (I375013,I374996,I374900);
DFFARX1 I_21901 (I375013,I2683,I374685,I374671,);
nor I_21902 (I374668,I374979,I374835);
or I_21903 (I374665,I374917,I374979);
nor I_21904 (I375072,I331952,I331955);
DFFARX1 I_21905 (I375072,I2683,I374685,I375098,);
not I_21906 (I375106,I375098);
nand I_21907 (I375123,I375106,I374784);
nor I_21908 (I375140,I375123,I331970);
DFFARX1 I_21909 (I375140,I2683,I374685,I374653,);
nor I_21910 (I375171,I375106,I374835);
nor I_21911 (I374662,I374979,I375171);
not I_21912 (I375229,I2690);
DFFARX1 I_21913 (I69138,I2683,I375229,I375255,);
nand I_21914 (I375263,I375255,I69153);
DFFARX1 I_21915 (I69150,I2683,I375229,I375289,);
DFFARX1 I_21916 (I375289,I2683,I375229,I375306,);
not I_21917 (I375221,I375306);
not I_21918 (I375328,I69129);
nor I_21919 (I375345,I69129,I69135);
not I_21920 (I375362,I69141);
nand I_21921 (I375379,I375328,I375362);
nor I_21922 (I375396,I69141,I69129);
and I_21923 (I375200,I375396,I375263);
not I_21924 (I375427,I69147);
nand I_21925 (I375444,I375427,I69129);
nor I_21926 (I375461,I69147,I69132);
not I_21927 (I375478,I375461);
nand I_21928 (I375203,I375345,I375478);
DFFARX1 I_21929 (I375461,I2683,I375229,I375218,);
nor I_21930 (I375523,I69132,I69141);
nor I_21931 (I375540,I375523,I69135);
and I_21932 (I375557,I375540,I375444);
DFFARX1 I_21933 (I375557,I2683,I375229,I375215,);
nor I_21934 (I375212,I375523,I375379);
or I_21935 (I375209,I375461,I375523);
nor I_21936 (I375616,I69132,I69144);
DFFARX1 I_21937 (I375616,I2683,I375229,I375642,);
not I_21938 (I375650,I375642);
nand I_21939 (I375667,I375650,I375328);
nor I_21940 (I375684,I375667,I69135);
DFFARX1 I_21941 (I375684,I2683,I375229,I375197,);
nor I_21942 (I375715,I375650,I375379);
nor I_21943 (I375206,I375523,I375715);
not I_21944 (I375773,I2690);
DFFARX1 I_21945 (I119002,I2683,I375773,I375799,);
nand I_21946 (I375807,I375799,I119005);
DFFARX1 I_21947 (I118999,I2683,I375773,I375833,);
DFFARX1 I_21948 (I375833,I2683,I375773,I375850,);
not I_21949 (I375765,I375850);
not I_21950 (I375872,I119008);
nor I_21951 (I375889,I119008,I118993);
not I_21952 (I375906,I119017);
nand I_21953 (I375923,I375872,I375906);
nor I_21954 (I375940,I119017,I119008);
and I_21955 (I375744,I375940,I375807);
not I_21956 (I375971,I118996);
nand I_21957 (I375988,I375971,I119014);
nor I_21958 (I376005,I118996,I118990);
not I_21959 (I376022,I376005);
nand I_21960 (I375747,I375889,I376022);
DFFARX1 I_21961 (I376005,I2683,I375773,I375762,);
nor I_21962 (I376067,I119011,I119017);
nor I_21963 (I376084,I376067,I118993);
and I_21964 (I376101,I376084,I375988);
DFFARX1 I_21965 (I376101,I2683,I375773,I375759,);
nor I_21966 (I375756,I376067,I375923);
or I_21967 (I375753,I376005,I376067);
nor I_21968 (I376160,I119011,I118990);
DFFARX1 I_21969 (I376160,I2683,I375773,I376186,);
not I_21970 (I376194,I376186);
nand I_21971 (I376211,I376194,I375872);
nor I_21972 (I376228,I376211,I118993);
DFFARX1 I_21973 (I376228,I2683,I375773,I375741,);
nor I_21974 (I376259,I376194,I375923);
nor I_21975 (I375750,I376067,I376259);
not I_21976 (I376317,I2690);
DFFARX1 I_21977 (I349891,I2683,I376317,I376343,);
nand I_21978 (I376351,I376343,I349870);
DFFARX1 I_21979 (I349867,I2683,I376317,I376377,);
DFFARX1 I_21980 (I376377,I2683,I376317,I376394,);
not I_21981 (I376309,I376394);
not I_21982 (I376416,I349879);
nor I_21983 (I376433,I349879,I349888);
not I_21984 (I376450,I349876);
nand I_21985 (I376467,I376416,I376450);
nor I_21986 (I376484,I349876,I349879);
and I_21987 (I376288,I376484,I376351);
not I_21988 (I376515,I349885);
nand I_21989 (I376532,I376515,I349882);
nor I_21990 (I376549,I349885,I349867);
not I_21991 (I376566,I376549);
nand I_21992 (I376291,I376433,I376566);
DFFARX1 I_21993 (I376549,I2683,I376317,I376306,);
nor I_21994 (I376611,I349870,I349876);
nor I_21995 (I376628,I376611,I349888);
and I_21996 (I376645,I376628,I376532);
DFFARX1 I_21997 (I376645,I2683,I376317,I376303,);
nor I_21998 (I376300,I376611,I376467);
or I_21999 (I376297,I376549,I376611);
nor I_22000 (I376704,I349870,I349873);
DFFARX1 I_22001 (I376704,I2683,I376317,I376730,);
not I_22002 (I376738,I376730);
nand I_22003 (I376755,I376738,I376416);
nor I_22004 (I376772,I376755,I349888);
DFFARX1 I_22005 (I376772,I2683,I376317,I376285,);
nor I_22006 (I376803,I376738,I376467);
nor I_22007 (I376294,I376611,I376803);
not I_22008 (I376861,I2690);
DFFARX1 I_22009 (I276886,I2683,I376861,I376887,);
nand I_22010 (I376895,I376887,I276886);
DFFARX1 I_22011 (I276898,I2683,I376861,I376921,);
DFFARX1 I_22012 (I376921,I2683,I376861,I376938,);
not I_22013 (I376853,I376938);
not I_22014 (I376960,I276892);
nor I_22015 (I376977,I276892,I276913);
not I_22016 (I376994,I276901);
nand I_22017 (I377011,I376960,I376994);
nor I_22018 (I377028,I276901,I276892);
and I_22019 (I376832,I377028,I376895);
not I_22020 (I377059,I276895);
nand I_22021 (I377076,I377059,I276910);
nor I_22022 (I377093,I276895,I276904);
not I_22023 (I377110,I377093);
nand I_22024 (I376835,I376977,I377110);
DFFARX1 I_22025 (I377093,I2683,I376861,I376850,);
nor I_22026 (I377155,I276907,I276901);
nor I_22027 (I377172,I377155,I276913);
and I_22028 (I377189,I377172,I377076);
DFFARX1 I_22029 (I377189,I2683,I376861,I376847,);
nor I_22030 (I376844,I377155,I377011);
or I_22031 (I376841,I377093,I377155);
nor I_22032 (I377248,I276907,I276889);
DFFARX1 I_22033 (I377248,I2683,I376861,I377274,);
not I_22034 (I377282,I377274);
nand I_22035 (I377299,I377282,I376960);
nor I_22036 (I377316,I377299,I276913);
DFFARX1 I_22037 (I377316,I2683,I376861,I376829,);
nor I_22038 (I377347,I377282,I377011);
nor I_22039 (I376838,I377155,I377347);
not I_22040 (I377405,I2690);
DFFARX1 I_22041 (I127463,I2683,I377405,I377431,);
nand I_22042 (I377439,I377431,I127460);
DFFARX1 I_22043 (I127439,I2683,I377405,I377465,);
DFFARX1 I_22044 (I377465,I2683,I377405,I377482,);
not I_22045 (I377397,I377482);
not I_22046 (I377504,I127454);
nor I_22047 (I377521,I127454,I127457);
not I_22048 (I377538,I127448);
nand I_22049 (I377555,I377504,I377538);
nor I_22050 (I377572,I127448,I127454);
and I_22051 (I377376,I377572,I377439);
not I_22052 (I377603,I127445);
nand I_22053 (I377620,I377603,I127466);
nor I_22054 (I377637,I127445,I127442);
not I_22055 (I377654,I377637);
nand I_22056 (I377379,I377521,I377654);
DFFARX1 I_22057 (I377637,I2683,I377405,I377394,);
nor I_22058 (I377699,I127451,I127448);
nor I_22059 (I377716,I377699,I127457);
and I_22060 (I377733,I377716,I377620);
DFFARX1 I_22061 (I377733,I2683,I377405,I377391,);
nor I_22062 (I377388,I377699,I377555);
or I_22063 (I377385,I377637,I377699);
nor I_22064 (I377792,I127451,I127439);
DFFARX1 I_22065 (I377792,I2683,I377405,I377818,);
not I_22066 (I377826,I377818);
nand I_22067 (I377843,I377826,I377504);
nor I_22068 (I377860,I377843,I127457);
DFFARX1 I_22069 (I377860,I2683,I377405,I377373,);
nor I_22070 (I377891,I377826,I377555);
nor I_22071 (I377382,I377699,I377891);
not I_22072 (I377949,I2690);
DFFARX1 I_22073 (I338331,I2683,I377949,I377975,);
nand I_22074 (I377983,I377975,I338310);
DFFARX1 I_22075 (I338307,I2683,I377949,I378009,);
DFFARX1 I_22076 (I378009,I2683,I377949,I378026,);
not I_22077 (I377941,I378026);
not I_22078 (I378048,I338319);
nor I_22079 (I378065,I338319,I338328);
not I_22080 (I378082,I338316);
nand I_22081 (I378099,I378048,I378082);
nor I_22082 (I378116,I338316,I338319);
and I_22083 (I377920,I378116,I377983);
not I_22084 (I378147,I338325);
nand I_22085 (I378164,I378147,I338322);
nor I_22086 (I378181,I338325,I338307);
not I_22087 (I378198,I378181);
nand I_22088 (I377923,I378065,I378198);
DFFARX1 I_22089 (I378181,I2683,I377949,I377938,);
nor I_22090 (I378243,I338310,I338316);
nor I_22091 (I378260,I378243,I338328);
and I_22092 (I378277,I378260,I378164);
DFFARX1 I_22093 (I378277,I2683,I377949,I377935,);
nor I_22094 (I377932,I378243,I378099);
or I_22095 (I377929,I378181,I378243);
nor I_22096 (I378336,I338310,I338313);
DFFARX1 I_22097 (I378336,I2683,I377949,I378362,);
not I_22098 (I378370,I378362);
nand I_22099 (I378387,I378370,I378048);
nor I_22100 (I378404,I378387,I338328);
DFFARX1 I_22101 (I378404,I2683,I377949,I377917,);
nor I_22102 (I378435,I378370,I378099);
nor I_22103 (I377926,I378243,I378435);
not I_22104 (I378493,I2690);
DFFARX1 I_22105 (I70328,I2683,I378493,I378519,);
nand I_22106 (I378527,I378519,I70343);
DFFARX1 I_22107 (I70340,I2683,I378493,I378553,);
DFFARX1 I_22108 (I378553,I2683,I378493,I378570,);
not I_22109 (I378485,I378570);
not I_22110 (I378592,I70319);
nor I_22111 (I378609,I70319,I70325);
not I_22112 (I378626,I70331);
nand I_22113 (I378643,I378592,I378626);
nor I_22114 (I378660,I70331,I70319);
and I_22115 (I378464,I378660,I378527);
not I_22116 (I378691,I70337);
nand I_22117 (I378708,I378691,I70319);
nor I_22118 (I378725,I70337,I70322);
not I_22119 (I378742,I378725);
nand I_22120 (I378467,I378609,I378742);
DFFARX1 I_22121 (I378725,I2683,I378493,I378482,);
nor I_22122 (I378787,I70322,I70331);
nor I_22123 (I378804,I378787,I70325);
and I_22124 (I378821,I378804,I378708);
DFFARX1 I_22125 (I378821,I2683,I378493,I378479,);
nor I_22126 (I378476,I378787,I378643);
or I_22127 (I378473,I378725,I378787);
nor I_22128 (I378880,I70322,I70334);
DFFARX1 I_22129 (I378880,I2683,I378493,I378906,);
not I_22130 (I378914,I378906);
nand I_22131 (I378931,I378914,I378592);
nor I_22132 (I378948,I378931,I70325);
DFFARX1 I_22133 (I378948,I2683,I378493,I378461,);
nor I_22134 (I378979,I378914,I378643);
nor I_22135 (I378470,I378787,I378979);
not I_22136 (I379037,I2690);
DFFARX1 I_22137 (I227909,I2683,I379037,I379063,);
nand I_22138 (I379071,I379063,I227912);
not I_22139 (I379088,I379071);
DFFARX1 I_22140 (I227924,I2683,I379037,I379114,);
not I_22141 (I379122,I379114);
not I_22142 (I379139,I227909);
or I_22143 (I379156,I227918,I227909);
nor I_22144 (I379173,I227918,I227909);
or I_22145 (I379190,I227927,I227918);
DFFARX1 I_22146 (I379190,I2683,I379037,I379029,);
not I_22147 (I379221,I227930);
nand I_22148 (I379238,I379221,I227912);
nand I_22149 (I379255,I379139,I379238);
and I_22150 (I379008,I379122,I379255);
nor I_22151 (I379286,I227930,I227915);
and I_22152 (I379303,I379122,I379286);
nor I_22153 (I379014,I379088,I379303);
DFFARX1 I_22154 (I379286,I2683,I379037,I379343,);
not I_22155 (I379351,I379343);
nor I_22156 (I379023,I379122,I379351);
or I_22157 (I379382,I379190,I227921);
nor I_22158 (I379399,I227921,I227927);
nand I_22159 (I379416,I379255,I379399);
nand I_22160 (I379433,I379382,I379416);
DFFARX1 I_22161 (I379433,I2683,I379037,I379026,);
nor I_22162 (I379464,I379399,I379156);
DFFARX1 I_22163 (I379464,I2683,I379037,I379005,);
nor I_22164 (I379495,I227921,I227933);
DFFARX1 I_22165 (I379495,I2683,I379037,I379521,);
DFFARX1 I_22166 (I379521,I2683,I379037,I379020,);
not I_22167 (I379543,I379521);
nand I_22168 (I379017,I379543,I379071);
nand I_22169 (I379011,I379543,I379173);
not I_22170 (I379615,I2690);
DFFARX1 I_22171 (I191498,I2683,I379615,I379641,);
nand I_22172 (I379649,I379641,I191513);
not I_22173 (I379666,I379649);
DFFARX1 I_22174 (I191495,I2683,I379615,I379692,);
not I_22175 (I379700,I379692);
not I_22176 (I379717,I191504);
or I_22177 (I379734,I191498,I191504);
nor I_22178 (I379751,I191498,I191504);
or I_22179 (I379768,I191495,I191498);
DFFARX1 I_22180 (I379768,I2683,I379615,I379607,);
not I_22181 (I379799,I191516);
nand I_22182 (I379816,I379799,I191519);
nand I_22183 (I379833,I379717,I379816);
and I_22184 (I379586,I379700,I379833);
nor I_22185 (I379864,I191516,I191501);
and I_22186 (I379881,I379700,I379864);
nor I_22187 (I379592,I379666,I379881);
DFFARX1 I_22188 (I379864,I2683,I379615,I379921,);
not I_22189 (I379929,I379921);
nor I_22190 (I379601,I379700,I379929);
or I_22191 (I379960,I379768,I191507);
nor I_22192 (I379977,I191507,I191495);
nand I_22193 (I379994,I379833,I379977);
nand I_22194 (I380011,I379960,I379994);
DFFARX1 I_22195 (I380011,I2683,I379615,I379604,);
nor I_22196 (I380042,I379977,I379734);
DFFARX1 I_22197 (I380042,I2683,I379615,I379583,);
nor I_22198 (I380073,I191507,I191510);
DFFARX1 I_22199 (I380073,I2683,I379615,I380099,);
DFFARX1 I_22200 (I380099,I2683,I379615,I379598,);
not I_22201 (I380121,I380099);
nand I_22202 (I379595,I380121,I379649);
nand I_22203 (I379589,I380121,I379751);
not I_22204 (I380193,I2690);
DFFARX1 I_22205 (I395139,I2683,I380193,I380219,);
nand I_22206 (I380227,I380219,I395133);
not I_22207 (I380244,I380227);
DFFARX1 I_22208 (I395148,I2683,I380193,I380270,);
not I_22209 (I380278,I380270);
not I_22210 (I380295,I395124);
or I_22211 (I380312,I395121,I395124);
nor I_22212 (I380329,I395121,I395124);
or I_22213 (I380346,I395127,I395121);
DFFARX1 I_22214 (I380346,I2683,I380193,I380185,);
not I_22215 (I380377,I395121);
nand I_22216 (I380394,I380377,I395136);
nand I_22217 (I380411,I380295,I380394);
and I_22218 (I380164,I380278,I380411);
nor I_22219 (I380442,I395121,I395130);
and I_22220 (I380459,I380278,I380442);
nor I_22221 (I380170,I380244,I380459);
DFFARX1 I_22222 (I380442,I2683,I380193,I380499,);
not I_22223 (I380507,I380499);
nor I_22224 (I380179,I380278,I380507);
or I_22225 (I380538,I380346,I395145);
nor I_22226 (I380555,I395145,I395127);
nand I_22227 (I380572,I380411,I380555);
nand I_22228 (I380589,I380538,I380572);
DFFARX1 I_22229 (I380589,I2683,I380193,I380182,);
nor I_22230 (I380620,I380555,I380312);
DFFARX1 I_22231 (I380620,I2683,I380193,I380161,);
nor I_22232 (I380651,I395145,I395142);
DFFARX1 I_22233 (I380651,I2683,I380193,I380677,);
DFFARX1 I_22234 (I380677,I2683,I380193,I380176,);
not I_22235 (I380699,I380677);
nand I_22236 (I380173,I380699,I380227);
nand I_22237 (I380167,I380699,I380329);
not I_22238 (I380771,I2690);
DFFARX1 I_22239 (I233111,I2683,I380771,I380797,);
nand I_22240 (I380805,I380797,I233114);
not I_22241 (I380822,I380805);
DFFARX1 I_22242 (I233126,I2683,I380771,I380848,);
not I_22243 (I380856,I380848);
not I_22244 (I380873,I233111);
or I_22245 (I380890,I233120,I233111);
nor I_22246 (I380907,I233120,I233111);
or I_22247 (I380924,I233129,I233120);
DFFARX1 I_22248 (I380924,I2683,I380771,I380763,);
not I_22249 (I380955,I233132);
nand I_22250 (I380972,I380955,I233114);
nand I_22251 (I380989,I380873,I380972);
and I_22252 (I380742,I380856,I380989);
nor I_22253 (I381020,I233132,I233117);
and I_22254 (I381037,I380856,I381020);
nor I_22255 (I380748,I380822,I381037);
DFFARX1 I_22256 (I381020,I2683,I380771,I381077,);
not I_22257 (I381085,I381077);
nor I_22258 (I380757,I380856,I381085);
or I_22259 (I381116,I380924,I233123);
nor I_22260 (I381133,I233123,I233129);
nand I_22261 (I381150,I380989,I381133);
nand I_22262 (I381167,I381116,I381150);
DFFARX1 I_22263 (I381167,I2683,I380771,I380760,);
nor I_22264 (I381198,I381133,I380890);
DFFARX1 I_22265 (I381198,I2683,I380771,I380739,);
nor I_22266 (I381229,I233123,I233135);
DFFARX1 I_22267 (I381229,I2683,I380771,I381255,);
DFFARX1 I_22268 (I381255,I2683,I380771,I380754,);
not I_22269 (I381277,I381255);
nand I_22270 (I380751,I381277,I380805);
nand I_22271 (I380745,I381277,I380907);
not I_22272 (I381349,I2690);
DFFARX1 I_22273 (I97916,I2683,I381349,I381375,);
nand I_22274 (I381383,I381375,I97937);
not I_22275 (I381400,I381383);
DFFARX1 I_22276 (I97931,I2683,I381349,I381426,);
not I_22277 (I381434,I381426);
not I_22278 (I381451,I97919);
or I_22279 (I381468,I97934,I97919);
nor I_22280 (I381485,I97934,I97919);
or I_22281 (I381502,I97925,I97934);
DFFARX1 I_22282 (I381502,I2683,I381349,I381341,);
not I_22283 (I381533,I97913);
nand I_22284 (I381550,I381533,I97910);
nand I_22285 (I381567,I381451,I381550);
and I_22286 (I381320,I381434,I381567);
nor I_22287 (I381598,I97913,I97922);
and I_22288 (I381615,I381434,I381598);
nor I_22289 (I381326,I381400,I381615);
DFFARX1 I_22290 (I381598,I2683,I381349,I381655,);
not I_22291 (I381663,I381655);
nor I_22292 (I381335,I381434,I381663);
or I_22293 (I381694,I381502,I97928);
nor I_22294 (I381711,I97928,I97925);
nand I_22295 (I381728,I381567,I381711);
nand I_22296 (I381745,I381694,I381728);
DFFARX1 I_22297 (I381745,I2683,I381349,I381338,);
nor I_22298 (I381776,I381711,I381468);
DFFARX1 I_22299 (I381776,I2683,I381349,I381317,);
nor I_22300 (I381807,I97928,I97910);
DFFARX1 I_22301 (I381807,I2683,I381349,I381833,);
DFFARX1 I_22302 (I381833,I2683,I381349,I381332,);
not I_22303 (I381855,I381833);
nand I_22304 (I381329,I381855,I381383);
nand I_22305 (I381323,I381855,I381485);
not I_22306 (I381927,I2690);
DFFARX1 I_22307 (I48304,I2683,I381927,I381953,);
nand I_22308 (I381961,I381953,I48307);
not I_22309 (I381978,I381961);
DFFARX1 I_22310 (I48316,I2683,I381927,I382004,);
not I_22311 (I382012,I382004);
not I_22312 (I382029,I48319);
or I_22313 (I382046,I48310,I48319);
nor I_22314 (I382063,I48310,I48319);
or I_22315 (I382080,I48322,I48310);
DFFARX1 I_22316 (I382080,I2683,I381927,I381919,);
not I_22317 (I382111,I48307);
nand I_22318 (I382128,I382111,I48313);
nand I_22319 (I382145,I382029,I382128);
and I_22320 (I381898,I382012,I382145);
nor I_22321 (I382176,I48307,I48325);
and I_22322 (I382193,I382012,I382176);
nor I_22323 (I381904,I381978,I382193);
DFFARX1 I_22324 (I382176,I2683,I381927,I382233,);
not I_22325 (I382241,I382233);
nor I_22326 (I381913,I382012,I382241);
or I_22327 (I382272,I382080,I48304);
nor I_22328 (I382289,I48304,I48322);
nand I_22329 (I382306,I382145,I382289);
nand I_22330 (I382323,I382272,I382306);
DFFARX1 I_22331 (I382323,I2683,I381927,I381916,);
nor I_22332 (I382354,I382289,I382046);
DFFARX1 I_22333 (I382354,I2683,I381927,I381895,);
nor I_22334 (I382385,I48304,I48328);
DFFARX1 I_22335 (I382385,I2683,I381927,I382411,);
DFFARX1 I_22336 (I382411,I2683,I381927,I381910,);
not I_22337 (I382433,I382411);
nand I_22338 (I381907,I382433,I381961);
nand I_22339 (I381901,I382433,I382063);
not I_22340 (I382505,I2690);
DFFARX1 I_22341 (I185140,I2683,I382505,I382531,);
nand I_22342 (I382539,I382531,I185155);
not I_22343 (I382556,I382539);
DFFARX1 I_22344 (I185137,I2683,I382505,I382582,);
not I_22345 (I382590,I382582);
not I_22346 (I382607,I185146);
or I_22347 (I382624,I185140,I185146);
nor I_22348 (I382641,I185140,I185146);
or I_22349 (I382658,I185137,I185140);
DFFARX1 I_22350 (I382658,I2683,I382505,I382497,);
not I_22351 (I382689,I185158);
nand I_22352 (I382706,I382689,I185161);
nand I_22353 (I382723,I382607,I382706);
and I_22354 (I382476,I382590,I382723);
nor I_22355 (I382754,I185158,I185143);
and I_22356 (I382771,I382590,I382754);
nor I_22357 (I382482,I382556,I382771);
DFFARX1 I_22358 (I382754,I2683,I382505,I382811,);
not I_22359 (I382819,I382811);
nor I_22360 (I382491,I382590,I382819);
or I_22361 (I382850,I382658,I185149);
nor I_22362 (I382867,I185149,I185137);
nand I_22363 (I382884,I382723,I382867);
nand I_22364 (I382901,I382850,I382884);
DFFARX1 I_22365 (I382901,I2683,I382505,I382494,);
nor I_22366 (I382932,I382867,I382624);
DFFARX1 I_22367 (I382932,I2683,I382505,I382473,);
nor I_22368 (I382963,I185149,I185152);
DFFARX1 I_22369 (I382963,I2683,I382505,I382989,);
DFFARX1 I_22370 (I382989,I2683,I382505,I382488,);
not I_22371 (I383011,I382989);
nand I_22372 (I382485,I383011,I382539);
nand I_22373 (I382479,I383011,I382641);
not I_22374 (I383083,I2690);
DFFARX1 I_22375 (I129074,I2683,I383083,I383109,);
nand I_22376 (I383117,I383109,I129083);
not I_22377 (I383134,I383117);
DFFARX1 I_22378 (I129071,I2683,I383083,I383160,);
not I_22379 (I383168,I383160);
not I_22380 (I383185,I129077);
or I_22381 (I383202,I129071,I129077);
nor I_22382 (I383219,I129071,I129077);
or I_22383 (I383236,I129086,I129071);
DFFARX1 I_22384 (I383236,I2683,I383083,I383075,);
not I_22385 (I383267,I129080);
nand I_22386 (I383284,I383267,I129095);
nand I_22387 (I383301,I383185,I383284);
and I_22388 (I383054,I383168,I383301);
nor I_22389 (I383332,I129080,I129098);
and I_22390 (I383349,I383168,I383332);
nor I_22391 (I383060,I383134,I383349);
DFFARX1 I_22392 (I383332,I2683,I383083,I383389,);
not I_22393 (I383397,I383389);
nor I_22394 (I383069,I383168,I383397);
or I_22395 (I383428,I383236,I129089);
nor I_22396 (I383445,I129089,I129086);
nand I_22397 (I383462,I383301,I383445);
nand I_22398 (I383479,I383428,I383462);
DFFARX1 I_22399 (I383479,I2683,I383083,I383072,);
nor I_22400 (I383510,I383445,I383202);
DFFARX1 I_22401 (I383510,I2683,I383083,I383051,);
nor I_22402 (I383541,I129089,I129092);
DFFARX1 I_22403 (I383541,I2683,I383083,I383567,);
DFFARX1 I_22404 (I383567,I2683,I383083,I383066,);
not I_22405 (I383589,I383567);
nand I_22406 (I383063,I383589,I383117);
nand I_22407 (I383057,I383589,I383219);
not I_22408 (I383661,I2690);
DFFARX1 I_22409 (I179938,I2683,I383661,I383687,);
nand I_22410 (I383695,I383687,I179953);
not I_22411 (I383712,I383695);
DFFARX1 I_22412 (I179935,I2683,I383661,I383738,);
not I_22413 (I383746,I383738);
not I_22414 (I383763,I179944);
or I_22415 (I383780,I179938,I179944);
nor I_22416 (I383797,I179938,I179944);
or I_22417 (I383814,I179935,I179938);
DFFARX1 I_22418 (I383814,I2683,I383661,I383653,);
not I_22419 (I383845,I179956);
nand I_22420 (I383862,I383845,I179959);
nand I_22421 (I383879,I383763,I383862);
and I_22422 (I383632,I383746,I383879);
nor I_22423 (I383910,I179956,I179941);
and I_22424 (I383927,I383746,I383910);
nor I_22425 (I383638,I383712,I383927);
DFFARX1 I_22426 (I383910,I2683,I383661,I383967,);
not I_22427 (I383975,I383967);
nor I_22428 (I383647,I383746,I383975);
or I_22429 (I384006,I383814,I179947);
nor I_22430 (I384023,I179947,I179935);
nand I_22431 (I384040,I383879,I384023);
nand I_22432 (I384057,I384006,I384040);
DFFARX1 I_22433 (I384057,I2683,I383661,I383650,);
nor I_22434 (I384088,I384023,I383780);
DFFARX1 I_22435 (I384088,I2683,I383661,I383629,);
nor I_22436 (I384119,I179947,I179950);
DFFARX1 I_22437 (I384119,I2683,I383661,I384145,);
DFFARX1 I_22438 (I384145,I2683,I383661,I383644,);
not I_22439 (I384167,I384145);
nand I_22440 (I383641,I384167,I383695);
nand I_22441 (I383635,I384167,I383797);
not I_22442 (I384239,I2690);
DFFARX1 I_22443 (I230221,I2683,I384239,I384265,);
nand I_22444 (I384273,I384265,I230224);
not I_22445 (I384290,I384273);
DFFARX1 I_22446 (I230236,I2683,I384239,I384316,);
not I_22447 (I384324,I384316);
not I_22448 (I384341,I230221);
or I_22449 (I384358,I230230,I230221);
nor I_22450 (I384375,I230230,I230221);
or I_22451 (I384392,I230239,I230230);
DFFARX1 I_22452 (I384392,I2683,I384239,I384231,);
not I_22453 (I384423,I230242);
nand I_22454 (I384440,I384423,I230224);
nand I_22455 (I384457,I384341,I384440);
and I_22456 (I384210,I384324,I384457);
nor I_22457 (I384488,I230242,I230227);
and I_22458 (I384505,I384324,I384488);
nor I_22459 (I384216,I384290,I384505);
DFFARX1 I_22460 (I384488,I2683,I384239,I384545,);
not I_22461 (I384553,I384545);
nor I_22462 (I384225,I384324,I384553);
or I_22463 (I384584,I384392,I230233);
nor I_22464 (I384601,I230233,I230239);
nand I_22465 (I384618,I384457,I384601);
nand I_22466 (I384635,I384584,I384618);
DFFARX1 I_22467 (I384635,I2683,I384239,I384228,);
nor I_22468 (I384666,I384601,I384358);
DFFARX1 I_22469 (I384666,I2683,I384239,I384207,);
nor I_22470 (I384697,I230233,I230245);
DFFARX1 I_22471 (I384697,I2683,I384239,I384723,);
DFFARX1 I_22472 (I384723,I2683,I384239,I384222,);
not I_22473 (I384745,I384723);
nand I_22474 (I384219,I384745,I384273);
nand I_22475 (I384213,I384745,I384375);
not I_22476 (I384817,I2690);
DFFARX1 I_22477 (I247649,I2683,I384817,I384843,);
nand I_22478 (I384851,I384843,I247649);
not I_22479 (I384868,I384851);
DFFARX1 I_22480 (I247655,I2683,I384817,I384894,);
not I_22481 (I384902,I384894);
not I_22482 (I384919,I247667);
or I_22483 (I384936,I247652,I247667);
nor I_22484 (I384953,I247652,I247667);
or I_22485 (I384970,I247646,I247652);
DFFARX1 I_22486 (I384970,I2683,I384817,I384809,);
not I_22487 (I385001,I247664);
nand I_22488 (I385018,I385001,I247658);
nand I_22489 (I385035,I384919,I385018);
and I_22490 (I384788,I384902,I385035);
nor I_22491 (I385066,I247664,I247646);
and I_22492 (I385083,I384902,I385066);
nor I_22493 (I384794,I384868,I385083);
DFFARX1 I_22494 (I385066,I2683,I384817,I385123,);
not I_22495 (I385131,I385123);
nor I_22496 (I384803,I384902,I385131);
or I_22497 (I385162,I384970,I247661);
nor I_22498 (I385179,I247661,I247646);
nand I_22499 (I385196,I385035,I385179);
nand I_22500 (I385213,I385162,I385196);
DFFARX1 I_22501 (I385213,I2683,I384817,I384806,);
nor I_22502 (I385244,I385179,I384936);
DFFARX1 I_22503 (I385244,I2683,I384817,I384785,);
nor I_22504 (I385275,I247661,I247652);
DFFARX1 I_22505 (I385275,I2683,I384817,I385301,);
DFFARX1 I_22506 (I385301,I2683,I384817,I384800,);
not I_22507 (I385323,I385301);
nand I_22508 (I384797,I385323,I384851);
nand I_22509 (I384791,I385323,I384953);
not I_22510 (I385395,I2690);
DFFARX1 I_22511 (I342371,I2683,I385395,I385421,);
nand I_22512 (I385429,I385421,I342356);
not I_22513 (I385446,I385429);
DFFARX1 I_22514 (I342359,I2683,I385395,I385472,);
not I_22515 (I385480,I385472);
not I_22516 (I385497,I342374);
or I_22517 (I385514,I342377,I342374);
nor I_22518 (I385531,I342377,I342374);
or I_22519 (I385548,I342353,I342377);
DFFARX1 I_22520 (I385548,I2683,I385395,I385387,);
not I_22521 (I385579,I342365);
nand I_22522 (I385596,I385579,I342368);
nand I_22523 (I385613,I385497,I385596);
and I_22524 (I385366,I385480,I385613);
nor I_22525 (I385644,I342365,I342362);
and I_22526 (I385661,I385480,I385644);
nor I_22527 (I385372,I385446,I385661);
DFFARX1 I_22528 (I385644,I2683,I385395,I385701,);
not I_22529 (I385709,I385701);
nor I_22530 (I385381,I385480,I385709);
or I_22531 (I385740,I385548,I342353);
nor I_22532 (I385757,I342353,I342353);
nand I_22533 (I385774,I385613,I385757);
nand I_22534 (I385791,I385740,I385774);
DFFARX1 I_22535 (I385791,I2683,I385395,I385384,);
nor I_22536 (I385822,I385757,I385514);
DFFARX1 I_22537 (I385822,I2683,I385395,I385363,);
nor I_22538 (I385853,I342353,I342356);
DFFARX1 I_22539 (I385853,I2683,I385395,I385879,);
DFFARX1 I_22540 (I385879,I2683,I385395,I385378,);
not I_22541 (I385901,I385879);
nand I_22542 (I385375,I385901,I385429);
nand I_22543 (I385369,I385901,I385531);
not I_22544 (I385973,I2690);
DFFARX1 I_22545 (I411703,I2683,I385973,I385999,);
nand I_22546 (I386007,I385999,I411694);
not I_22547 (I386024,I386007);
DFFARX1 I_22548 (I411679,I2683,I385973,I386050,);
not I_22549 (I386058,I386050);
not I_22550 (I386075,I411682);
or I_22551 (I386092,I411691,I411682);
nor I_22552 (I386109,I411691,I411682);
or I_22553 (I386126,I411688,I411691);
DFFARX1 I_22554 (I386126,I2683,I385973,I385965,);
not I_22555 (I386157,I411700);
nand I_22556 (I386174,I386157,I411679);
nand I_22557 (I386191,I386075,I386174);
and I_22558 (I385944,I386058,I386191);
nor I_22559 (I386222,I411700,I411685);
and I_22560 (I386239,I386058,I386222);
nor I_22561 (I385950,I386024,I386239);
DFFARX1 I_22562 (I386222,I2683,I385973,I386279,);
not I_22563 (I386287,I386279);
nor I_22564 (I385959,I386058,I386287);
or I_22565 (I386318,I386126,I411706);
nor I_22566 (I386335,I411706,I411688);
nand I_22567 (I386352,I386191,I386335);
nand I_22568 (I386369,I386318,I386352);
DFFARX1 I_22569 (I386369,I2683,I385973,I385962,);
nor I_22570 (I386400,I386335,I386092);
DFFARX1 I_22571 (I386400,I2683,I385973,I385941,);
nor I_22572 (I386431,I411706,I411697);
DFFARX1 I_22573 (I386431,I2683,I385973,I386457,);
DFFARX1 I_22574 (I386457,I2683,I385973,I385956,);
not I_22575 (I386479,I386457);
nand I_22576 (I385953,I386479,I386007);
nand I_22577 (I385947,I386479,I386109);
not I_22578 (I386551,I2690);
DFFARX1 I_22579 (I14633,I2683,I386551,I386577,);
nand I_22580 (I386585,I386577,I14627);
not I_22581 (I386602,I386585);
DFFARX1 I_22582 (I14645,I2683,I386551,I386628,);
not I_22583 (I386636,I386628);
not I_22584 (I386653,I14648);
or I_22585 (I386670,I14651,I14648);
nor I_22586 (I386687,I14651,I14648);
or I_22587 (I386704,I14636,I14651);
DFFARX1 I_22588 (I386704,I2683,I386551,I386543,);
not I_22589 (I386735,I14639);
nand I_22590 (I386752,I386735,I14642);
nand I_22591 (I386769,I386653,I386752);
and I_22592 (I386522,I386636,I386769);
nor I_22593 (I386800,I14639,I14630);
and I_22594 (I386817,I386636,I386800);
nor I_22595 (I386528,I386602,I386817);
DFFARX1 I_22596 (I386800,I2683,I386551,I386857,);
not I_22597 (I386865,I386857);
nor I_22598 (I386537,I386636,I386865);
or I_22599 (I386896,I386704,I14630);
nor I_22600 (I386913,I14630,I14636);
nand I_22601 (I386930,I386769,I386913);
nand I_22602 (I386947,I386896,I386930);
DFFARX1 I_22603 (I386947,I2683,I386551,I386540,);
nor I_22604 (I386978,I386913,I386670);
DFFARX1 I_22605 (I386978,I2683,I386551,I386519,);
nor I_22606 (I387009,I14630,I14627);
DFFARX1 I_22607 (I387009,I2683,I386551,I387035,);
DFFARX1 I_22608 (I387035,I2683,I386551,I386534,);
not I_22609 (I387057,I387035);
nand I_22610 (I386531,I387057,I386585);
nand I_22611 (I386525,I387057,I386687);
not I_22612 (I387129,I2690);
DFFARX1 I_22613 (I235423,I2683,I387129,I387155,);
nand I_22614 (I387163,I387155,I235426);
not I_22615 (I387180,I387163);
DFFARX1 I_22616 (I235438,I2683,I387129,I387206,);
not I_22617 (I387214,I387206);
not I_22618 (I387231,I235423);
or I_22619 (I387248,I235432,I235423);
nor I_22620 (I387265,I235432,I235423);
or I_22621 (I387282,I235441,I235432);
DFFARX1 I_22622 (I387282,I2683,I387129,I387121,);
not I_22623 (I387313,I235444);
nand I_22624 (I387330,I387313,I235426);
nand I_22625 (I387347,I387231,I387330);
and I_22626 (I387100,I387214,I387347);
nor I_22627 (I387378,I235444,I235429);
and I_22628 (I387395,I387214,I387378);
nor I_22629 (I387106,I387180,I387395);
DFFARX1 I_22630 (I387378,I2683,I387129,I387435,);
not I_22631 (I387443,I387435);
nor I_22632 (I387115,I387214,I387443);
or I_22633 (I387474,I387282,I235435);
nor I_22634 (I387491,I235435,I235441);
nand I_22635 (I387508,I387347,I387491);
nand I_22636 (I387525,I387474,I387508);
DFFARX1 I_22637 (I387525,I2683,I387129,I387118,);
nor I_22638 (I387556,I387491,I387248);
DFFARX1 I_22639 (I387556,I2683,I387129,I387097,);
nor I_22640 (I387587,I235435,I235447);
DFFARX1 I_22641 (I387587,I2683,I387129,I387613,);
DFFARX1 I_22642 (I387613,I2683,I387129,I387112,);
not I_22643 (I387635,I387613);
nand I_22644 (I387109,I387635,I387163);
nand I_22645 (I387103,I387635,I387265);
not I_22646 (I387707,I2690);
DFFARX1 I_22647 (I13052,I2683,I387707,I387733,);
nand I_22648 (I387741,I387733,I13046);
not I_22649 (I387758,I387741);
DFFARX1 I_22650 (I13064,I2683,I387707,I387784,);
not I_22651 (I387792,I387784);
not I_22652 (I387809,I13067);
or I_22653 (I387826,I13070,I13067);
nor I_22654 (I387843,I13070,I13067);
or I_22655 (I387860,I13055,I13070);
DFFARX1 I_22656 (I387860,I2683,I387707,I387699,);
not I_22657 (I387891,I13058);
nand I_22658 (I387908,I387891,I13061);
nand I_22659 (I387925,I387809,I387908);
and I_22660 (I387678,I387792,I387925);
nor I_22661 (I387956,I13058,I13049);
and I_22662 (I387973,I387792,I387956);
nor I_22663 (I387684,I387758,I387973);
DFFARX1 I_22664 (I387956,I2683,I387707,I388013,);
not I_22665 (I388021,I388013);
nor I_22666 (I387693,I387792,I388021);
or I_22667 (I388052,I387860,I13049);
nor I_22668 (I388069,I13049,I13055);
nand I_22669 (I388086,I387925,I388069);
nand I_22670 (I388103,I388052,I388086);
DFFARX1 I_22671 (I388103,I2683,I387707,I387696,);
nor I_22672 (I388134,I388069,I387826);
DFFARX1 I_22673 (I388134,I2683,I387707,I387675,);
nor I_22674 (I388165,I13049,I13046);
DFFARX1 I_22675 (I388165,I2683,I387707,I388191,);
DFFARX1 I_22676 (I388191,I2683,I387707,I387690,);
not I_22677 (I388213,I388191);
nand I_22678 (I387687,I388213,I387741);
nand I_22679 (I387681,I388213,I387843);
not I_22680 (I388285,I2690);
DFFARX1 I_22681 (I1628,I2683,I388285,I388311,);
nand I_22682 (I388319,I388311,I1404);
not I_22683 (I388336,I388319);
DFFARX1 I_22684 (I1820,I2683,I388285,I388362,);
not I_22685 (I388370,I388362);
not I_22686 (I388387,I2636);
or I_22687 (I388404,I1868,I2636);
nor I_22688 (I388421,I1868,I2636);
or I_22689 (I388438,I2412,I1868);
DFFARX1 I_22690 (I388438,I2683,I388285,I388277,);
not I_22691 (I388469,I2076);
nand I_22692 (I388486,I388469,I1828);
nand I_22693 (I388503,I388387,I388486);
and I_22694 (I388256,I388370,I388503);
nor I_22695 (I388534,I2076,I1532);
and I_22696 (I388551,I388370,I388534);
nor I_22697 (I388262,I388336,I388551);
DFFARX1 I_22698 (I388534,I2683,I388285,I388591,);
not I_22699 (I388599,I388591);
nor I_22700 (I388271,I388370,I388599);
or I_22701 (I388630,I388438,I1652);
nor I_22702 (I388647,I1652,I2412);
nand I_22703 (I388664,I388503,I388647);
nand I_22704 (I388681,I388630,I388664);
DFFARX1 I_22705 (I388681,I2683,I388285,I388274,);
nor I_22706 (I388712,I388647,I388404);
DFFARX1 I_22707 (I388712,I2683,I388285,I388253,);
nor I_22708 (I388743,I1652,I2092);
DFFARX1 I_22709 (I388743,I2683,I388285,I388769,);
DFFARX1 I_22710 (I388769,I2683,I388285,I388268,);
not I_22711 (I388791,I388769);
nand I_22712 (I388265,I388791,I388319);
nand I_22713 (I388259,I388791,I388421);
not I_22714 (I388863,I2690);
DFFARX1 I_22715 (I175314,I2683,I388863,I388889,);
nand I_22716 (I388897,I388889,I175329);
not I_22717 (I388914,I388897);
DFFARX1 I_22718 (I175311,I2683,I388863,I388940,);
not I_22719 (I388948,I388940);
not I_22720 (I388965,I175320);
or I_22721 (I388982,I175314,I175320);
nor I_22722 (I388999,I175314,I175320);
or I_22723 (I389016,I175311,I175314);
DFFARX1 I_22724 (I389016,I2683,I388863,I388855,);
not I_22725 (I389047,I175332);
nand I_22726 (I389064,I389047,I175335);
nand I_22727 (I389081,I388965,I389064);
and I_22728 (I388834,I388948,I389081);
nor I_22729 (I389112,I175332,I175317);
and I_22730 (I389129,I388948,I389112);
nor I_22731 (I388840,I388914,I389129);
DFFARX1 I_22732 (I389112,I2683,I388863,I389169,);
not I_22733 (I389177,I389169);
nor I_22734 (I388849,I388948,I389177);
or I_22735 (I389208,I389016,I175323);
nor I_22736 (I389225,I175323,I175311);
nand I_22737 (I389242,I389081,I389225);
nand I_22738 (I389259,I389208,I389242);
DFFARX1 I_22739 (I389259,I2683,I388863,I388852,);
nor I_22740 (I389290,I389225,I388982);
DFFARX1 I_22741 (I389290,I2683,I388863,I388831,);
nor I_22742 (I389321,I175323,I175326);
DFFARX1 I_22743 (I389321,I2683,I388863,I389347,);
DFFARX1 I_22744 (I389347,I2683,I388863,I388846,);
not I_22745 (I389369,I389347);
nand I_22746 (I388843,I389369,I388897);
nand I_22747 (I388837,I389369,I388999);
not I_22748 (I389441,I2690);
DFFARX1 I_22749 (I298856,I2683,I389441,I389467,);
nand I_22750 (I389475,I389467,I298877);
not I_22751 (I389492,I389475);
DFFARX1 I_22752 (I298850,I2683,I389441,I389518,);
not I_22753 (I389526,I389518);
not I_22754 (I389543,I298871);
or I_22755 (I389560,I298862,I298871);
nor I_22756 (I389577,I298862,I298871);
or I_22757 (I389594,I298865,I298862);
DFFARX1 I_22758 (I389594,I2683,I389441,I389433,);
not I_22759 (I389625,I298853);
nand I_22760 (I389642,I389625,I298868);
nand I_22761 (I389659,I389543,I389642);
and I_22762 (I389412,I389526,I389659);
nor I_22763 (I389690,I298853,I298850);
and I_22764 (I389707,I389526,I389690);
nor I_22765 (I389418,I389492,I389707);
DFFARX1 I_22766 (I389690,I2683,I389441,I389747,);
not I_22767 (I389755,I389747);
nor I_22768 (I389427,I389526,I389755);
or I_22769 (I389786,I389594,I298874);
nor I_22770 (I389803,I298874,I298865);
nand I_22771 (I389820,I389659,I389803);
nand I_22772 (I389837,I389786,I389820);
DFFARX1 I_22773 (I389837,I2683,I389441,I389430,);
nor I_22774 (I389868,I389803,I389560);
DFFARX1 I_22775 (I389868,I2683,I389441,I389409,);
nor I_22776 (I389899,I298874,I298859);
DFFARX1 I_22777 (I389899,I2683,I389441,I389925,);
DFFARX1 I_22778 (I389925,I2683,I389441,I389424,);
not I_22779 (I389947,I389925);
nand I_22780 (I389421,I389947,I389475);
nand I_22781 (I389415,I389947,I389577);
not I_22782 (I390019,I2690);
DFFARX1 I_22783 (I289166,I2683,I390019,I390045,);
nand I_22784 (I390053,I390045,I289187);
not I_22785 (I390070,I390053);
DFFARX1 I_22786 (I289160,I2683,I390019,I390096,);
not I_22787 (I390104,I390096);
not I_22788 (I390121,I289181);
or I_22789 (I390138,I289172,I289181);
nor I_22790 (I390155,I289172,I289181);
or I_22791 (I390172,I289175,I289172);
DFFARX1 I_22792 (I390172,I2683,I390019,I390011,);
not I_22793 (I390203,I289163);
nand I_22794 (I390220,I390203,I289178);
nand I_22795 (I390237,I390121,I390220);
and I_22796 (I389990,I390104,I390237);
nor I_22797 (I390268,I289163,I289160);
and I_22798 (I390285,I390104,I390268);
nor I_22799 (I389996,I390070,I390285);
DFFARX1 I_22800 (I390268,I2683,I390019,I390325,);
not I_22801 (I390333,I390325);
nor I_22802 (I390005,I390104,I390333);
or I_22803 (I390364,I390172,I289184);
nor I_22804 (I390381,I289184,I289175);
nand I_22805 (I390398,I390237,I390381);
nand I_22806 (I390415,I390364,I390398);
DFFARX1 I_22807 (I390415,I2683,I390019,I390008,);
nor I_22808 (I390446,I390381,I390138);
DFFARX1 I_22809 (I390446,I2683,I390019,I389987,);
nor I_22810 (I390477,I289184,I289169);
DFFARX1 I_22811 (I390477,I2683,I390019,I390503,);
DFFARX1 I_22812 (I390503,I2683,I390019,I390002,);
not I_22813 (I390525,I390503);
nand I_22814 (I389999,I390525,I390053);
nand I_22815 (I389993,I390525,I390155);
not I_22816 (I390597,I2690);
DFFARX1 I_22817 (I293688,I2683,I390597,I390623,);
nand I_22818 (I390631,I390623,I293709);
not I_22819 (I390648,I390631);
DFFARX1 I_22820 (I293682,I2683,I390597,I390674,);
not I_22821 (I390682,I390674);
not I_22822 (I390699,I293703);
or I_22823 (I390716,I293694,I293703);
nor I_22824 (I390733,I293694,I293703);
or I_22825 (I390750,I293697,I293694);
DFFARX1 I_22826 (I390750,I2683,I390597,I390589,);
not I_22827 (I390781,I293685);
nand I_22828 (I390798,I390781,I293700);
nand I_22829 (I390815,I390699,I390798);
and I_22830 (I390568,I390682,I390815);
nor I_22831 (I390846,I293685,I293682);
and I_22832 (I390863,I390682,I390846);
nor I_22833 (I390574,I390648,I390863);
DFFARX1 I_22834 (I390846,I2683,I390597,I390903,);
not I_22835 (I390911,I390903);
nor I_22836 (I390583,I390682,I390911);
or I_22837 (I390942,I390750,I293706);
nor I_22838 (I390959,I293706,I293697);
nand I_22839 (I390976,I390815,I390959);
nand I_22840 (I390993,I390942,I390976);
DFFARX1 I_22841 (I390993,I2683,I390597,I390586,);
nor I_22842 (I391024,I390959,I390716);
DFFARX1 I_22843 (I391024,I2683,I390597,I390565,);
nor I_22844 (I391055,I293706,I293691);
DFFARX1 I_22845 (I391055,I2683,I390597,I391081,);
DFFARX1 I_22846 (I391081,I2683,I390597,I390580,);
not I_22847 (I391103,I391081);
nand I_22848 (I390577,I391103,I390631);
nand I_22849 (I390571,I391103,I390733);
not I_22850 (I391175,I2690);
DFFARX1 I_22851 (I160589,I2683,I391175,I391201,);
nand I_22852 (I391209,I391201,I160598);
not I_22853 (I391226,I391209);
DFFARX1 I_22854 (I160610,I2683,I391175,I391252,);
not I_22855 (I391260,I391252);
not I_22856 (I391277,I160601);
or I_22857 (I391294,I160595,I160601);
nor I_22858 (I391311,I160595,I160601);
or I_22859 (I391328,I160589,I160595);
DFFARX1 I_22860 (I391328,I2683,I391175,I391167,);
not I_22861 (I391359,I160592);
nand I_22862 (I391376,I391359,I160604);
nand I_22863 (I391393,I391277,I391376);
and I_22864 (I391146,I391260,I391393);
nor I_22865 (I391424,I160592,I160613);
and I_22866 (I391441,I391260,I391424);
nor I_22867 (I391152,I391226,I391441);
DFFARX1 I_22868 (I391424,I2683,I391175,I391481,);
not I_22869 (I391489,I391481);
nor I_22870 (I391161,I391260,I391489);
or I_22871 (I391520,I391328,I160607);
nor I_22872 (I391537,I160607,I160589);
nand I_22873 (I391554,I391393,I391537);
nand I_22874 (I391571,I391520,I391554);
DFFARX1 I_22875 (I391571,I2683,I391175,I391164,);
nor I_22876 (I391602,I391537,I391294);
DFFARX1 I_22877 (I391602,I2683,I391175,I391143,);
nor I_22878 (I391633,I160607,I160592);
DFFARX1 I_22879 (I391633,I2683,I391175,I391659,);
DFFARX1 I_22880 (I391659,I2683,I391175,I391158,);
not I_22881 (I391681,I391659);
nand I_22882 (I391155,I391681,I391209);
nand I_22883 (I391149,I391681,I391311);
not I_22884 (I391753,I2690);
DFFARX1 I_22885 (I225597,I2683,I391753,I391779,);
nand I_22886 (I391787,I391779,I225600);
not I_22887 (I391804,I391787);
DFFARX1 I_22888 (I225612,I2683,I391753,I391830,);
not I_22889 (I391838,I391830);
not I_22890 (I391855,I225597);
or I_22891 (I391872,I225606,I225597);
nor I_22892 (I391889,I225606,I225597);
or I_22893 (I391906,I225615,I225606);
DFFARX1 I_22894 (I391906,I2683,I391753,I391745,);
not I_22895 (I391937,I225618);
nand I_22896 (I391954,I391937,I225600);
nand I_22897 (I391971,I391855,I391954);
and I_22898 (I391724,I391838,I391971);
nor I_22899 (I392002,I225618,I225603);
and I_22900 (I392019,I391838,I392002);
nor I_22901 (I391730,I391804,I392019);
DFFARX1 I_22902 (I392002,I2683,I391753,I392059,);
not I_22903 (I392067,I392059);
nor I_22904 (I391739,I391838,I392067);
or I_22905 (I392098,I391906,I225609);
nor I_22906 (I392115,I225609,I225615);
nand I_22907 (I392132,I391971,I392115);
nand I_22908 (I392149,I392098,I392132);
DFFARX1 I_22909 (I392149,I2683,I391753,I391742,);
nor I_22910 (I392180,I392115,I391872);
DFFARX1 I_22911 (I392180,I2683,I391753,I391721,);
nor I_22912 (I392211,I225609,I225621);
DFFARX1 I_22913 (I392211,I2683,I391753,I392237,);
DFFARX1 I_22914 (I392237,I2683,I391753,I391736,);
not I_22915 (I392259,I392237);
nand I_22916 (I391733,I392259,I391787);
nand I_22917 (I391727,I392259,I391889);
not I_22918 (I392331,I2690);
DFFARX1 I_22919 (I245014,I2683,I392331,I392357,);
nand I_22920 (I392365,I392357,I245014);
not I_22921 (I392382,I392365);
DFFARX1 I_22922 (I245020,I2683,I392331,I392408,);
not I_22923 (I392416,I392408);
not I_22924 (I392433,I245032);
or I_22925 (I392450,I245017,I245032);
nor I_22926 (I392467,I245017,I245032);
or I_22927 (I392484,I245011,I245017);
DFFARX1 I_22928 (I392484,I2683,I392331,I392323,);
not I_22929 (I392515,I245029);
nand I_22930 (I392532,I392515,I245023);
nand I_22931 (I392549,I392433,I392532);
and I_22932 (I392302,I392416,I392549);
nor I_22933 (I392580,I245029,I245011);
and I_22934 (I392597,I392416,I392580);
nor I_22935 (I392308,I392382,I392597);
DFFARX1 I_22936 (I392580,I2683,I392331,I392637,);
not I_22937 (I392645,I392637);
nor I_22938 (I392317,I392416,I392645);
or I_22939 (I392676,I392484,I245026);
nor I_22940 (I392693,I245026,I245011);
nand I_22941 (I392710,I392549,I392693);
nand I_22942 (I392727,I392676,I392710);
DFFARX1 I_22943 (I392727,I2683,I392331,I392320,);
nor I_22944 (I392758,I392693,I392450);
DFFARX1 I_22945 (I392758,I2683,I392331,I392299,);
nor I_22946 (I392789,I245026,I245017);
DFFARX1 I_22947 (I392789,I2683,I392331,I392815,);
DFFARX1 I_22948 (I392815,I2683,I392331,I392314,);
not I_22949 (I392837,I392815);
nand I_22950 (I392311,I392837,I392365);
nand I_22951 (I392305,I392837,I392467);
not I_22952 (I392912,I2690);
DFFARX1 I_22953 (I128004,I2683,I392912,I392938,);
nand I_22954 (I392946,I392938,I127986);
not I_22955 (I392963,I392946);
DFFARX1 I_22956 (I127983,I2683,I392912,I392989,);
not I_22957 (I392997,I392989);
nor I_22958 (I393014,I127989,I127983);
not I_22959 (I393031,I393014);
DFFARX1 I_22960 (I393031,I2683,I392912,I392898,);
or I_22961 (I393062,I127992,I127989);
DFFARX1 I_22962 (I393062,I2683,I392912,I392901,);
not I_22963 (I393093,I127998);
nor I_22964 (I393110,I393093,I128010);
nor I_22965 (I393127,I393110,I127983);
nor I_22966 (I393144,I128010,I127995);
nor I_22967 (I393161,I392997,I393144);
nor I_22968 (I392886,I392963,I393161);
not I_22969 (I393192,I393144);
nand I_22970 (I392889,I393192,I392946);
nand I_22971 (I392883,I393192,I393014);
nor I_22972 (I392880,I393144,I393127);
nor I_22973 (I393251,I128001,I127992);
not I_22974 (I393268,I393251);
DFFARX1 I_22975 (I393251,I2683,I392912,I393294,);
not I_22976 (I392904,I393294);
nor I_22977 (I393316,I128001,I128007);
DFFARX1 I_22978 (I393316,I2683,I392912,I393342,);
and I_22979 (I393350,I393342,I127989);
nor I_22980 (I393367,I393350,I393268);
DFFARX1 I_22981 (I393367,I2683,I392912,I392895,);
nor I_22982 (I393398,I393342,I393127);
DFFARX1 I_22983 (I393398,I2683,I392912,I392877,);
nor I_22984 (I392892,I393342,I393031);
not I_22985 (I393473,I2690);
DFFARX1 I_22986 (I192097,I2683,I393473,I393499,);
nand I_22987 (I393507,I393499,I192076);
not I_22988 (I393524,I393507);
DFFARX1 I_22989 (I192088,I2683,I393473,I393550,);
not I_22990 (I393558,I393550);
nor I_22991 (I393575,I192076,I192085);
not I_22992 (I393592,I393575);
DFFARX1 I_22993 (I393592,I2683,I393473,I393459,);
or I_22994 (I393623,I192079,I192076);
DFFARX1 I_22995 (I393623,I2683,I393473,I393462,);
not I_22996 (I393654,I192082);
nor I_22997 (I393671,I393654,I192073);
nor I_22998 (I393688,I393671,I192085);
nor I_22999 (I393705,I192073,I192091);
nor I_23000 (I393722,I393558,I393705);
nor I_23001 (I393447,I393524,I393722);
not I_23002 (I393753,I393705);
nand I_23003 (I393450,I393753,I393507);
nand I_23004 (I393444,I393753,I393575);
nor I_23005 (I393441,I393705,I393688);
nor I_23006 (I393812,I192094,I192079);
not I_23007 (I393829,I393812);
DFFARX1 I_23008 (I393812,I2683,I393473,I393855,);
not I_23009 (I393465,I393855);
nor I_23010 (I393877,I192094,I192073);
DFFARX1 I_23011 (I393877,I2683,I393473,I393903,);
and I_23012 (I393911,I393903,I192076);
nor I_23013 (I393928,I393911,I393829);
DFFARX1 I_23014 (I393928,I2683,I393473,I393456,);
nor I_23015 (I393959,I393903,I393688);
DFFARX1 I_23016 (I393959,I2683,I393473,I393438,);
nor I_23017 (I393453,I393903,I393592);
not I_23018 (I394034,I2690);
DFFARX1 I_23019 (I33623,I2683,I394034,I394060,);
nand I_23020 (I394068,I394060,I33614);
not I_23021 (I394085,I394068);
DFFARX1 I_23022 (I33602,I2683,I394034,I394111,);
not I_23023 (I394119,I394111);
nor I_23024 (I394136,I33605,I33602);
not I_23025 (I394153,I394136);
DFFARX1 I_23026 (I394153,I2683,I394034,I394020,);
or I_23027 (I394184,I33599,I33605);
DFFARX1 I_23028 (I394184,I2683,I394034,I394023,);
not I_23029 (I394215,I33608);
nor I_23030 (I394232,I394215,I33599);
nor I_23031 (I394249,I394232,I33602);
nor I_23032 (I394266,I33599,I33611);
nor I_23033 (I394283,I394119,I394266);
nor I_23034 (I394008,I394085,I394283);
not I_23035 (I394314,I394266);
nand I_23036 (I394011,I394314,I394068);
nand I_23037 (I394005,I394314,I394136);
nor I_23038 (I394002,I394266,I394249);
nor I_23039 (I394373,I33617,I33599);
not I_23040 (I394390,I394373);
DFFARX1 I_23041 (I394373,I2683,I394034,I394416,);
not I_23042 (I394026,I394416);
nor I_23043 (I394438,I33617,I33620);
DFFARX1 I_23044 (I394438,I2683,I394034,I394464,);
and I_23045 (I394472,I394464,I33605);
nor I_23046 (I394489,I394472,I394390);
DFFARX1 I_23047 (I394489,I2683,I394034,I394017,);
nor I_23048 (I394520,I394464,I394249);
DFFARX1 I_23049 (I394520,I2683,I394034,I393999,);
nor I_23050 (I394014,I394464,I394153);
not I_23051 (I394595,I2690);
DFFARX1 I_23052 (I302750,I2683,I394595,I394621,);
nand I_23053 (I394629,I394621,I302732);
not I_23054 (I394646,I394629);
DFFARX1 I_23055 (I302744,I2683,I394595,I394672,);
not I_23056 (I394680,I394672);
nor I_23057 (I394697,I302726,I302726);
not I_23058 (I394714,I394697);
DFFARX1 I_23059 (I394714,I2683,I394595,I394581,);
or I_23060 (I394745,I302738,I302726);
DFFARX1 I_23061 (I394745,I2683,I394595,I394584,);
not I_23062 (I394776,I302753);
nor I_23063 (I394793,I394776,I302741);
nor I_23064 (I394810,I394793,I302726);
nor I_23065 (I394827,I302741,I302729);
nor I_23066 (I394844,I394680,I394827);
nor I_23067 (I394569,I394646,I394844);
not I_23068 (I394875,I394827);
nand I_23069 (I394572,I394875,I394629);
nand I_23070 (I394566,I394875,I394697);
nor I_23071 (I394563,I394827,I394810);
nor I_23072 (I394934,I302735,I302738);
not I_23073 (I394951,I394934);
DFFARX1 I_23074 (I394934,I2683,I394595,I394977,);
not I_23075 (I394587,I394977);
nor I_23076 (I394999,I302735,I302747);
DFFARX1 I_23077 (I394999,I2683,I394595,I395025,);
and I_23078 (I395033,I395025,I302726);
nor I_23079 (I395050,I395033,I394951);
DFFARX1 I_23080 (I395050,I2683,I394595,I394578,);
nor I_23081 (I395081,I395025,I394810);
DFFARX1 I_23082 (I395081,I2683,I394595,I394560,);
nor I_23083 (I394575,I395025,I394714);
not I_23084 (I395156,I2690);
DFFARX1 I_23085 (I95823,I2683,I395156,I395182,);
nand I_23086 (I395190,I395182,I95802);
not I_23087 (I395207,I395190);
DFFARX1 I_23088 (I95811,I2683,I395156,I395233,);
not I_23089 (I395241,I395233);
nor I_23090 (I395258,I95805,I95817);
not I_23091 (I395275,I395258);
DFFARX1 I_23092 (I395275,I2683,I395156,I395142,);
or I_23093 (I395306,I95808,I95805);
DFFARX1 I_23094 (I395306,I2683,I395156,I395145,);
not I_23095 (I395337,I95829);
nor I_23096 (I395354,I395337,I95814);
nor I_23097 (I395371,I395354,I95817);
nor I_23098 (I395388,I95814,I95802);
nor I_23099 (I395405,I395241,I395388);
nor I_23100 (I395130,I395207,I395405);
not I_23101 (I395436,I395388);
nand I_23102 (I395133,I395436,I395190);
nand I_23103 (I395127,I395436,I395258);
nor I_23104 (I395124,I395388,I395371);
nor I_23105 (I395495,I95820,I95808);
not I_23106 (I395512,I395495);
DFFARX1 I_23107 (I395495,I2683,I395156,I395538,);
not I_23108 (I395148,I395538);
nor I_23109 (I395560,I95820,I95826);
DFFARX1 I_23110 (I395560,I2683,I395156,I395586,);
and I_23111 (I395594,I395586,I95805);
nor I_23112 (I395611,I395594,I395512);
DFFARX1 I_23113 (I395611,I2683,I395156,I395139,);
nor I_23114 (I395642,I395586,I395371);
DFFARX1 I_23115 (I395642,I2683,I395156,I395121,);
nor I_23116 (I395136,I395586,I395275);
not I_23117 (I395717,I2690);
DFFARX1 I_23118 (I280786,I2683,I395717,I395743,);
nand I_23119 (I395751,I395743,I280768);
not I_23120 (I395768,I395751);
DFFARX1 I_23121 (I280780,I2683,I395717,I395794,);
not I_23122 (I395802,I395794);
nor I_23123 (I395819,I280762,I280762);
not I_23124 (I395836,I395819);
DFFARX1 I_23125 (I395836,I2683,I395717,I395703,);
or I_23126 (I395867,I280774,I280762);
DFFARX1 I_23127 (I395867,I2683,I395717,I395706,);
not I_23128 (I395898,I280789);
nor I_23129 (I395915,I395898,I280777);
nor I_23130 (I395932,I395915,I280762);
nor I_23131 (I395949,I280777,I280765);
nor I_23132 (I395966,I395802,I395949);
nor I_23133 (I395691,I395768,I395966);
not I_23134 (I395997,I395949);
nand I_23135 (I395694,I395997,I395751);
nand I_23136 (I395688,I395997,I395819);
nor I_23137 (I395685,I395949,I395932);
nor I_23138 (I396056,I280771,I280774);
not I_23139 (I396073,I396056);
DFFARX1 I_23140 (I396056,I2683,I395717,I396099,);
not I_23141 (I395709,I396099);
nor I_23142 (I396121,I280771,I280783);
DFFARX1 I_23143 (I396121,I2683,I395717,I396147,);
and I_23144 (I396155,I396147,I280762);
nor I_23145 (I396172,I396155,I396073);
DFFARX1 I_23146 (I396172,I2683,I395717,I395700,);
nor I_23147 (I396203,I396147,I395932);
DFFARX1 I_23148 (I396203,I2683,I395717,I395682,);
nor I_23149 (I395697,I396147,I395836);
not I_23150 (I396278,I2690);
DFFARX1 I_23151 (I18328,I2683,I396278,I396304,);
nand I_23152 (I396312,I396304,I18322);
not I_23153 (I396329,I396312);
DFFARX1 I_23154 (I18319,I2683,I396278,I396355,);
not I_23155 (I396363,I396355);
nor I_23156 (I396380,I18319,I18325);
not I_23157 (I396397,I396380);
DFFARX1 I_23158 (I396397,I2683,I396278,I396264,);
or I_23159 (I396428,I18334,I18319);
DFFARX1 I_23160 (I396428,I2683,I396278,I396267,);
not I_23161 (I396459,I18316);
nor I_23162 (I396476,I396459,I18340);
nor I_23163 (I396493,I396476,I18325);
nor I_23164 (I396510,I18340,I18316);
nor I_23165 (I396527,I396363,I396510);
nor I_23166 (I396252,I396329,I396527);
not I_23167 (I396558,I396510);
nand I_23168 (I396255,I396558,I396312);
nand I_23169 (I396249,I396558,I396380);
nor I_23170 (I396246,I396510,I396493);
nor I_23171 (I396617,I18337,I18334);
not I_23172 (I396634,I396617);
DFFARX1 I_23173 (I396617,I2683,I396278,I396660,);
not I_23174 (I396270,I396660);
nor I_23175 (I396682,I18337,I18331);
DFFARX1 I_23176 (I396682,I2683,I396278,I396708,);
and I_23177 (I396716,I396708,I18319);
nor I_23178 (I396733,I396716,I396634);
DFFARX1 I_23179 (I396733,I2683,I396278,I396261,);
nor I_23180 (I396764,I396708,I396493);
DFFARX1 I_23181 (I396764,I2683,I396278,I396243,);
nor I_23182 (I396258,I396708,I396397);
not I_23183 (I396839,I2690);
DFFARX1 I_23184 (I283998,I2683,I396839,I396865,);
DFFARX1 I_23185 (I284016,I2683,I396839,I396882,);
not I_23186 (I396890,I396882);
nor I_23187 (I396807,I396865,I396890);
DFFARX1 I_23188 (I396890,I2683,I396839,I396822,);
nor I_23189 (I396935,I283995,I284007);
and I_23190 (I396952,I396935,I283992);
nor I_23191 (I396969,I396952,I283995);
not I_23192 (I396986,I283995);
and I_23193 (I397003,I396986,I284001);
nand I_23194 (I397020,I397003,I284013);
nor I_23195 (I397037,I396986,I397020);
DFFARX1 I_23196 (I397037,I2683,I396839,I396804,);
not I_23197 (I397068,I397020);
nand I_23198 (I397085,I396890,I397068);
nand I_23199 (I396816,I396952,I397068);
DFFARX1 I_23200 (I396986,I2683,I396839,I396831,);
not I_23201 (I397130,I284004);
nor I_23202 (I397147,I397130,I284001);
nor I_23203 (I397164,I397147,I396969);
DFFARX1 I_23204 (I397164,I2683,I396839,I396828,);
not I_23205 (I397195,I397147);
DFFARX1 I_23206 (I397195,I2683,I396839,I397221,);
not I_23207 (I397229,I397221);
nor I_23208 (I396825,I397229,I397147);
nor I_23209 (I397260,I397130,I283992);
and I_23210 (I397277,I397260,I284019);
or I_23211 (I397294,I397277,I284010);
DFFARX1 I_23212 (I397294,I2683,I396839,I397320,);
not I_23213 (I397328,I397320);
nand I_23214 (I397345,I397328,I397068);
not I_23215 (I396819,I397345);
nand I_23216 (I396813,I397345,I397085);
nand I_23217 (I396810,I397328,I396952);
not I_23218 (I397434,I2690);
DFFARX1 I_23219 (I50684,I2683,I397434,I397460,);
DFFARX1 I_23220 (I50687,I2683,I397434,I397477,);
not I_23221 (I397485,I397477);
nor I_23222 (I397402,I397460,I397485);
DFFARX1 I_23223 (I397485,I2683,I397434,I397417,);
nor I_23224 (I397530,I50693,I50687);
and I_23225 (I397547,I397530,I50690);
nor I_23226 (I397564,I397547,I50693);
not I_23227 (I397581,I50693);
and I_23228 (I397598,I397581,I50684);
nand I_23229 (I397615,I397598,I50702);
nor I_23230 (I397632,I397581,I397615);
DFFARX1 I_23231 (I397632,I2683,I397434,I397399,);
not I_23232 (I397663,I397615);
nand I_23233 (I397680,I397485,I397663);
nand I_23234 (I397411,I397547,I397663);
DFFARX1 I_23235 (I397581,I2683,I397434,I397426,);
not I_23236 (I397725,I50696);
nor I_23237 (I397742,I397725,I50684);
nor I_23238 (I397759,I397742,I397564);
DFFARX1 I_23239 (I397759,I2683,I397434,I397423,);
not I_23240 (I397790,I397742);
DFFARX1 I_23241 (I397790,I2683,I397434,I397816,);
not I_23242 (I397824,I397816);
nor I_23243 (I397420,I397824,I397742);
nor I_23244 (I397855,I397725,I50699);
and I_23245 (I397872,I397855,I50705);
or I_23246 (I397889,I397872,I50708);
DFFARX1 I_23247 (I397889,I2683,I397434,I397915,);
not I_23248 (I397923,I397915);
nand I_23249 (I397940,I397923,I397663);
not I_23250 (I397414,I397940);
nand I_23251 (I397408,I397940,I397680);
nand I_23252 (I397405,I397923,I397547);
not I_23253 (I398029,I2690);
DFFARX1 I_23254 (I367037,I2683,I398029,I398055,);
DFFARX1 I_23255 (I367040,I2683,I398029,I398072,);
not I_23256 (I398080,I398072);
nor I_23257 (I397997,I398055,I398080);
DFFARX1 I_23258 (I398080,I2683,I398029,I398012,);
nor I_23259 (I398125,I367040,I367055);
and I_23260 (I398142,I398125,I367049);
nor I_23261 (I398159,I398142,I367040);
not I_23262 (I398176,I367040);
and I_23263 (I398193,I398176,I367058);
nand I_23264 (I398210,I398193,I367046);
nor I_23265 (I398227,I398176,I398210);
DFFARX1 I_23266 (I398227,I2683,I398029,I397994,);
not I_23267 (I398258,I398210);
nand I_23268 (I398275,I398080,I398258);
nand I_23269 (I398006,I398142,I398258);
DFFARX1 I_23270 (I398176,I2683,I398029,I398021,);
not I_23271 (I398320,I367052);
nor I_23272 (I398337,I398320,I367058);
nor I_23273 (I398354,I398337,I398159);
DFFARX1 I_23274 (I398354,I2683,I398029,I398018,);
not I_23275 (I398385,I398337);
DFFARX1 I_23276 (I398385,I2683,I398029,I398411,);
not I_23277 (I398419,I398411);
nor I_23278 (I398015,I398419,I398337);
nor I_23279 (I398450,I398320,I367037);
and I_23280 (I398467,I398450,I367061);
or I_23281 (I398484,I398467,I367043);
DFFARX1 I_23282 (I398484,I2683,I398029,I398510,);
not I_23283 (I398518,I398510);
nand I_23284 (I398535,I398518,I398258);
not I_23285 (I398009,I398535);
nand I_23286 (I398003,I398535,I398275);
nand I_23287 (I398000,I398518,I398142);
not I_23288 (I398624,I2690);
DFFARX1 I_23289 (I8848,I2683,I398624,I398650,);
DFFARX1 I_23290 (I8830,I2683,I398624,I398667,);
not I_23291 (I398675,I398667);
nor I_23292 (I398592,I398650,I398675);
DFFARX1 I_23293 (I398675,I2683,I398624,I398607,);
nor I_23294 (I398720,I8830,I8845);
and I_23295 (I398737,I398720,I8839);
nor I_23296 (I398754,I398737,I8830);
not I_23297 (I398771,I8830);
and I_23298 (I398788,I398771,I8833);
nand I_23299 (I398805,I398788,I8836);
nor I_23300 (I398822,I398771,I398805);
DFFARX1 I_23301 (I398822,I2683,I398624,I398589,);
not I_23302 (I398853,I398805);
nand I_23303 (I398870,I398675,I398853);
nand I_23304 (I398601,I398737,I398853);
DFFARX1 I_23305 (I398771,I2683,I398624,I398616,);
not I_23306 (I398915,I8842);
nor I_23307 (I398932,I398915,I8833);
nor I_23308 (I398949,I398932,I398754);
DFFARX1 I_23309 (I398949,I2683,I398624,I398613,);
not I_23310 (I398980,I398932);
DFFARX1 I_23311 (I398980,I2683,I398624,I399006,);
not I_23312 (I399014,I399006);
nor I_23313 (I398610,I399014,I398932);
nor I_23314 (I399045,I398915,I8854);
and I_23315 (I399062,I399045,I8851);
or I_23316 (I399079,I399062,I8833);
DFFARX1 I_23317 (I399079,I2683,I398624,I399105,);
not I_23318 (I399113,I399105);
nand I_23319 (I399130,I399113,I398853);
not I_23320 (I398604,I399130);
nand I_23321 (I398598,I399130,I398870);
nand I_23322 (I398595,I399113,I398737);
not I_23323 (I399219,I2690);
DFFARX1 I_23324 (I188626,I2683,I399219,I399245,);
DFFARX1 I_23325 (I188620,I2683,I399219,I399262,);
not I_23326 (I399270,I399262);
nor I_23327 (I399187,I399245,I399270);
DFFARX1 I_23328 (I399270,I2683,I399219,I399202,);
nor I_23329 (I399315,I188617,I188608);
and I_23330 (I399332,I399315,I188605);
nor I_23331 (I399349,I399332,I188617);
not I_23332 (I399366,I188617);
and I_23333 (I399383,I399366,I188611);
nand I_23334 (I399400,I399383,I188623);
nor I_23335 (I399417,I399366,I399400);
DFFARX1 I_23336 (I399417,I2683,I399219,I399184,);
not I_23337 (I399448,I399400);
nand I_23338 (I399465,I399270,I399448);
nand I_23339 (I399196,I399332,I399448);
DFFARX1 I_23340 (I399366,I2683,I399219,I399211,);
not I_23341 (I399510,I188629);
nor I_23342 (I399527,I399510,I188611);
nor I_23343 (I399544,I399527,I399349);
DFFARX1 I_23344 (I399544,I2683,I399219,I399208,);
not I_23345 (I399575,I399527);
DFFARX1 I_23346 (I399575,I2683,I399219,I399601,);
not I_23347 (I399609,I399601);
nor I_23348 (I399205,I399609,I399527);
nor I_23349 (I399640,I399510,I188608);
and I_23350 (I399657,I399640,I188614);
or I_23351 (I399674,I399657,I188605);
DFFARX1 I_23352 (I399674,I2683,I399219,I399700,);
not I_23353 (I399708,I399700);
nand I_23354 (I399725,I399708,I399448);
not I_23355 (I399199,I399725);
nand I_23356 (I399193,I399725,I399465);
nand I_23357 (I399190,I399708,I399332);
not I_23358 (I399814,I2690);
DFFARX1 I_23359 (I242385,I2683,I399814,I399840,);
DFFARX1 I_23360 (I242382,I2683,I399814,I399857,);
not I_23361 (I399865,I399857);
nor I_23362 (I399782,I399840,I399865);
DFFARX1 I_23363 (I399865,I2683,I399814,I399797,);
nor I_23364 (I399910,I242397,I242379);
and I_23365 (I399927,I399910,I242376);
nor I_23366 (I399944,I399927,I242397);
not I_23367 (I399961,I242397);
and I_23368 (I399978,I399961,I242382);
nand I_23369 (I399995,I399978,I242394);
nor I_23370 (I400012,I399961,I399995);
DFFARX1 I_23371 (I400012,I2683,I399814,I399779,);
not I_23372 (I400043,I399995);
nand I_23373 (I400060,I399865,I400043);
nand I_23374 (I399791,I399927,I400043);
DFFARX1 I_23375 (I399961,I2683,I399814,I399806,);
not I_23376 (I400105,I242388);
nor I_23377 (I400122,I400105,I242382);
nor I_23378 (I400139,I400122,I399944);
DFFARX1 I_23379 (I400139,I2683,I399814,I399803,);
not I_23380 (I400170,I400122);
DFFARX1 I_23381 (I400170,I2683,I399814,I400196,);
not I_23382 (I400204,I400196);
nor I_23383 (I399800,I400204,I400122);
nor I_23384 (I400235,I400105,I242376);
and I_23385 (I400252,I400235,I242391);
or I_23386 (I400269,I400252,I242379);
DFFARX1 I_23387 (I400269,I2683,I399814,I400295,);
not I_23388 (I400303,I400295);
nand I_23389 (I400320,I400303,I400043);
not I_23390 (I399794,I400320);
nand I_23391 (I399788,I400320,I400060);
nand I_23392 (I399785,I400303,I399927);
not I_23393 (I400409,I2690);
DFFARX1 I_23394 (I319381,I2683,I400409,I400435,);
DFFARX1 I_23395 (I319372,I2683,I400409,I400452,);
not I_23396 (I400460,I400452);
nor I_23397 (I400377,I400435,I400460);
DFFARX1 I_23398 (I400460,I2683,I400409,I400392,);
nor I_23399 (I400505,I319378,I319387);
and I_23400 (I400522,I400505,I319390);
nor I_23401 (I400539,I400522,I319378);
not I_23402 (I400556,I319378);
and I_23403 (I400573,I400556,I319369);
nand I_23404 (I400590,I400573,I319375);
nor I_23405 (I400607,I400556,I400590);
DFFARX1 I_23406 (I400607,I2683,I400409,I400374,);
not I_23407 (I400638,I400590);
nand I_23408 (I400655,I400460,I400638);
nand I_23409 (I400386,I400522,I400638);
DFFARX1 I_23410 (I400556,I2683,I400409,I400401,);
not I_23411 (I400700,I319384);
nor I_23412 (I400717,I400700,I319369);
nor I_23413 (I400734,I400717,I400539);
DFFARX1 I_23414 (I400734,I2683,I400409,I400398,);
not I_23415 (I400765,I400717);
DFFARX1 I_23416 (I400765,I2683,I400409,I400791,);
not I_23417 (I400799,I400791);
nor I_23418 (I400395,I400799,I400717);
nor I_23419 (I400830,I400700,I319369);
and I_23420 (I400847,I400830,I319372);
or I_23421 (I400864,I400847,I319375);
DFFARX1 I_23422 (I400864,I2683,I400409,I400890,);
not I_23423 (I400898,I400890);
nand I_23424 (I400915,I400898,I400638);
not I_23425 (I400389,I400915);
nand I_23426 (I400383,I400915,I400655);
nand I_23427 (I400380,I400898,I400522);
not I_23428 (I401004,I2690);
DFFARX1 I_23429 (I135599,I2683,I401004,I401030,);
DFFARX1 I_23430 (I135605,I2683,I401004,I401047,);
not I_23431 (I401055,I401047);
nor I_23432 (I400972,I401030,I401055);
DFFARX1 I_23433 (I401055,I2683,I401004,I400987,);
nor I_23434 (I401100,I135614,I135599);
and I_23435 (I401117,I401100,I135626);
nor I_23436 (I401134,I401117,I135614);
not I_23437 (I401151,I135614);
and I_23438 (I401168,I401151,I135602);
nand I_23439 (I401185,I401168,I135623);
nor I_23440 (I401202,I401151,I401185);
DFFARX1 I_23441 (I401202,I2683,I401004,I400969,);
not I_23442 (I401233,I401185);
nand I_23443 (I401250,I401055,I401233);
nand I_23444 (I400981,I401117,I401233);
DFFARX1 I_23445 (I401151,I2683,I401004,I400996,);
not I_23446 (I401295,I135611);
nor I_23447 (I401312,I401295,I135602);
nor I_23448 (I401329,I401312,I401134);
DFFARX1 I_23449 (I401329,I2683,I401004,I400993,);
not I_23450 (I401360,I401312);
DFFARX1 I_23451 (I401360,I2683,I401004,I401386,);
not I_23452 (I401394,I401386);
nor I_23453 (I400990,I401394,I401312);
nor I_23454 (I401425,I401295,I135608);
and I_23455 (I401442,I401425,I135620);
or I_23456 (I401459,I401442,I135617);
DFFARX1 I_23457 (I401459,I2683,I401004,I401485,);
not I_23458 (I401493,I401485);
nand I_23459 (I401510,I401493,I401233);
not I_23460 (I400984,I401510);
nand I_23461 (I400978,I401510,I401250);
nand I_23462 (I400975,I401493,I401117);
not I_23463 (I401599,I2690);
DFFARX1 I_23464 (I54254,I2683,I401599,I401625,);
DFFARX1 I_23465 (I54257,I2683,I401599,I401642,);
not I_23466 (I401650,I401642);
nor I_23467 (I401567,I401625,I401650);
DFFARX1 I_23468 (I401650,I2683,I401599,I401582,);
nor I_23469 (I401695,I54263,I54257);
and I_23470 (I401712,I401695,I54260);
nor I_23471 (I401729,I401712,I54263);
not I_23472 (I401746,I54263);
and I_23473 (I401763,I401746,I54254);
nand I_23474 (I401780,I401763,I54272);
nor I_23475 (I401797,I401746,I401780);
DFFARX1 I_23476 (I401797,I2683,I401599,I401564,);
not I_23477 (I401828,I401780);
nand I_23478 (I401845,I401650,I401828);
nand I_23479 (I401576,I401712,I401828);
DFFARX1 I_23480 (I401746,I2683,I401599,I401591,);
not I_23481 (I401890,I54266);
nor I_23482 (I401907,I401890,I54254);
nor I_23483 (I401924,I401907,I401729);
DFFARX1 I_23484 (I401924,I2683,I401599,I401588,);
not I_23485 (I401955,I401907);
DFFARX1 I_23486 (I401955,I2683,I401599,I401981,);
not I_23487 (I401989,I401981);
nor I_23488 (I401585,I401989,I401907);
nor I_23489 (I402020,I401890,I54269);
and I_23490 (I402037,I402020,I54275);
or I_23491 (I402054,I402037,I54278);
DFFARX1 I_23492 (I402054,I2683,I401599,I402080,);
not I_23493 (I402088,I402080);
nand I_23494 (I402105,I402088,I401828);
not I_23495 (I401579,I402105);
nand I_23496 (I401573,I402105,I401845);
nand I_23497 (I401570,I402088,I401712);
not I_23498 (I402194,I2690);
DFFARX1 I_23499 (I117957,I2683,I402194,I402220,);
DFFARX1 I_23500 (I117951,I2683,I402194,I402237,);
not I_23501 (I402245,I402237);
nor I_23502 (I402162,I402220,I402245);
DFFARX1 I_23503 (I402245,I2683,I402194,I402177,);
nor I_23504 (I402290,I117939,I117960);
and I_23505 (I402307,I402290,I117954);
nor I_23506 (I402324,I402307,I117939);
not I_23507 (I402341,I117939);
and I_23508 (I402358,I402341,I117936);
nand I_23509 (I402375,I402358,I117948);
nor I_23510 (I402392,I402341,I402375);
DFFARX1 I_23511 (I402392,I2683,I402194,I402159,);
not I_23512 (I402423,I402375);
nand I_23513 (I402440,I402245,I402423);
nand I_23514 (I402171,I402307,I402423);
DFFARX1 I_23515 (I402341,I2683,I402194,I402186,);
not I_23516 (I402485,I117963);
nor I_23517 (I402502,I402485,I117936);
nor I_23518 (I402519,I402502,I402324);
DFFARX1 I_23519 (I402519,I2683,I402194,I402183,);
not I_23520 (I402550,I402502);
DFFARX1 I_23521 (I402550,I2683,I402194,I402576,);
not I_23522 (I402584,I402576);
nor I_23523 (I402180,I402584,I402502);
nor I_23524 (I402615,I402485,I117945);
and I_23525 (I402632,I402615,I117942);
or I_23526 (I402649,I402632,I117936);
DFFARX1 I_23527 (I402649,I2683,I402194,I402675,);
not I_23528 (I402683,I402675);
nand I_23529 (I402700,I402683,I402423);
not I_23530 (I402174,I402700);
nand I_23531 (I402168,I402700,I402440);
nand I_23532 (I402165,I402683,I402307);
not I_23533 (I402789,I2690);
DFFARX1 I_23534 (I85810,I2683,I402789,I402815,);
DFFARX1 I_23535 (I85804,I2683,I402789,I402832,);
not I_23536 (I402840,I402832);
nor I_23537 (I402757,I402815,I402840);
DFFARX1 I_23538 (I402840,I2683,I402789,I402772,);
nor I_23539 (I402885,I85792,I85813);
and I_23540 (I402902,I402885,I85807);
nor I_23541 (I402919,I402902,I85792);
not I_23542 (I402936,I85792);
and I_23543 (I402953,I402936,I85789);
nand I_23544 (I402970,I402953,I85801);
nor I_23545 (I402987,I402936,I402970);
DFFARX1 I_23546 (I402987,I2683,I402789,I402754,);
not I_23547 (I403018,I402970);
nand I_23548 (I403035,I402840,I403018);
nand I_23549 (I402766,I402902,I403018);
DFFARX1 I_23550 (I402936,I2683,I402789,I402781,);
not I_23551 (I403080,I85816);
nor I_23552 (I403097,I403080,I85789);
nor I_23553 (I403114,I403097,I402919);
DFFARX1 I_23554 (I403114,I2683,I402789,I402778,);
not I_23555 (I403145,I403097);
DFFARX1 I_23556 (I403145,I2683,I402789,I403171,);
not I_23557 (I403179,I403171);
nor I_23558 (I402775,I403179,I403097);
nor I_23559 (I403210,I403080,I85798);
and I_23560 (I403227,I403210,I85795);
or I_23561 (I403244,I403227,I85789);
DFFARX1 I_23562 (I403244,I2683,I402789,I403270,);
not I_23563 (I403278,I403270);
nand I_23564 (I403295,I403278,I403018);
not I_23565 (I402769,I403295);
nand I_23566 (I402763,I403295,I403035);
nand I_23567 (I402760,I403278,I402902);
not I_23568 (I403384,I2690);
DFFARX1 I_23569 (I34674,I2683,I403384,I403410,);
DFFARX1 I_23570 (I34662,I2683,I403384,I403427,);
not I_23571 (I403435,I403427);
nor I_23572 (I403352,I403410,I403435);
DFFARX1 I_23573 (I403435,I2683,I403384,I403367,);
nor I_23574 (I403480,I34653,I34677);
and I_23575 (I403497,I403480,I34656);
nor I_23576 (I403514,I403497,I34653);
not I_23577 (I403531,I34653);
and I_23578 (I403548,I403531,I34659);
nand I_23579 (I403565,I403548,I34671);
nor I_23580 (I403582,I403531,I403565);
DFFARX1 I_23581 (I403582,I2683,I403384,I403349,);
not I_23582 (I403613,I403565);
nand I_23583 (I403630,I403435,I403613);
nand I_23584 (I403361,I403497,I403613);
DFFARX1 I_23585 (I403531,I2683,I403384,I403376,);
not I_23586 (I403675,I34653);
nor I_23587 (I403692,I403675,I34659);
nor I_23588 (I403709,I403692,I403514);
DFFARX1 I_23589 (I403709,I2683,I403384,I403373,);
not I_23590 (I403740,I403692);
DFFARX1 I_23591 (I403740,I2683,I403384,I403766,);
not I_23592 (I403774,I403766);
nor I_23593 (I403370,I403774,I403692);
nor I_23594 (I403805,I403675,I34656);
and I_23595 (I403822,I403805,I34665);
or I_23596 (I403839,I403822,I34668);
DFFARX1 I_23597 (I403839,I2683,I403384,I403865,);
not I_23598 (I403873,I403865);
nand I_23599 (I403890,I403873,I403613);
not I_23600 (I403364,I403890);
nand I_23601 (I403358,I403890,I403630);
nand I_23602 (I403355,I403873,I403497);
not I_23603 (I403979,I2690);
DFFARX1 I_23604 (I116903,I2683,I403979,I404005,);
DFFARX1 I_23605 (I116897,I2683,I403979,I404022,);
not I_23606 (I404030,I404022);
nor I_23607 (I403947,I404005,I404030);
DFFARX1 I_23608 (I404030,I2683,I403979,I403962,);
nor I_23609 (I404075,I116885,I116906);
and I_23610 (I404092,I404075,I116900);
nor I_23611 (I404109,I404092,I116885);
not I_23612 (I404126,I116885);
and I_23613 (I404143,I404126,I116882);
nand I_23614 (I404160,I404143,I116894);
nor I_23615 (I404177,I404126,I404160);
DFFARX1 I_23616 (I404177,I2683,I403979,I403944,);
not I_23617 (I404208,I404160);
nand I_23618 (I404225,I404030,I404208);
nand I_23619 (I403956,I404092,I404208);
DFFARX1 I_23620 (I404126,I2683,I403979,I403971,);
not I_23621 (I404270,I116909);
nor I_23622 (I404287,I404270,I116882);
nor I_23623 (I404304,I404287,I404109);
DFFARX1 I_23624 (I404304,I2683,I403979,I403968,);
not I_23625 (I404335,I404287);
DFFARX1 I_23626 (I404335,I2683,I403979,I404361,);
not I_23627 (I404369,I404361);
nor I_23628 (I403965,I404369,I404287);
nor I_23629 (I404400,I404270,I116891);
and I_23630 (I404417,I404400,I116888);
or I_23631 (I404434,I404417,I116882);
DFFARX1 I_23632 (I404434,I2683,I403979,I404460,);
not I_23633 (I404468,I404460);
nand I_23634 (I404485,I404468,I404208);
not I_23635 (I403959,I404485);
nand I_23636 (I403953,I404485,I404225);
nand I_23637 (I403950,I404468,I404092);
not I_23638 (I404574,I2690);
DFFARX1 I_23639 (I35201,I2683,I404574,I404600,);
DFFARX1 I_23640 (I35189,I2683,I404574,I404617,);
not I_23641 (I404625,I404617);
nor I_23642 (I404542,I404600,I404625);
DFFARX1 I_23643 (I404625,I2683,I404574,I404557,);
nor I_23644 (I404670,I35180,I35204);
and I_23645 (I404687,I404670,I35183);
nor I_23646 (I404704,I404687,I35180);
not I_23647 (I404721,I35180);
and I_23648 (I404738,I404721,I35186);
nand I_23649 (I404755,I404738,I35198);
nor I_23650 (I404772,I404721,I404755);
DFFARX1 I_23651 (I404772,I2683,I404574,I404539,);
not I_23652 (I404803,I404755);
nand I_23653 (I404820,I404625,I404803);
nand I_23654 (I404551,I404687,I404803);
DFFARX1 I_23655 (I404721,I2683,I404574,I404566,);
not I_23656 (I404865,I35180);
nor I_23657 (I404882,I404865,I35186);
nor I_23658 (I404899,I404882,I404704);
DFFARX1 I_23659 (I404899,I2683,I404574,I404563,);
not I_23660 (I404930,I404882);
DFFARX1 I_23661 (I404930,I2683,I404574,I404956,);
not I_23662 (I404964,I404956);
nor I_23663 (I404560,I404964,I404882);
nor I_23664 (I404995,I404865,I35183);
and I_23665 (I405012,I404995,I35192);
or I_23666 (I405029,I405012,I35195);
DFFARX1 I_23667 (I405029,I2683,I404574,I405055,);
not I_23668 (I405063,I405055);
nand I_23669 (I405080,I405063,I404803);
not I_23670 (I404554,I405080);
nand I_23671 (I404548,I405080,I404820);
nand I_23672 (I404545,I405063,I404687);
not I_23673 (I405169,I2690);
DFFARX1 I_23674 (I227352,I2683,I405169,I405195,);
DFFARX1 I_23675 (I227334,I2683,I405169,I405212,);
not I_23676 (I405220,I405212);
nor I_23677 (I405137,I405195,I405220);
DFFARX1 I_23678 (I405220,I2683,I405169,I405152,);
nor I_23679 (I405265,I227340,I227343);
and I_23680 (I405282,I405265,I227331);
nor I_23681 (I405299,I405282,I227340);
not I_23682 (I405316,I227340);
and I_23683 (I405333,I405316,I227349);
nand I_23684 (I405350,I405333,I227337);
nor I_23685 (I405367,I405316,I405350);
DFFARX1 I_23686 (I405367,I2683,I405169,I405134,);
not I_23687 (I405398,I405350);
nand I_23688 (I405415,I405220,I405398);
nand I_23689 (I405146,I405282,I405398);
DFFARX1 I_23690 (I405316,I2683,I405169,I405161,);
not I_23691 (I405460,I227334);
nor I_23692 (I405477,I405460,I227349);
nor I_23693 (I405494,I405477,I405299);
DFFARX1 I_23694 (I405494,I2683,I405169,I405158,);
not I_23695 (I405525,I405477);
DFFARX1 I_23696 (I405525,I2683,I405169,I405551,);
not I_23697 (I405559,I405551);
nor I_23698 (I405155,I405559,I405477);
nor I_23699 (I405590,I405460,I227346);
and I_23700 (I405607,I405590,I227355);
or I_23701 (I405624,I405607,I227331);
DFFARX1 I_23702 (I405624,I2683,I405169,I405650,);
not I_23703 (I405658,I405650);
nand I_23704 (I405675,I405658,I405398);
not I_23705 (I405149,I405675);
nand I_23706 (I405143,I405675,I405415);
nand I_23707 (I405140,I405658,I405282);
not I_23708 (I405764,I2690);
DFFARX1 I_23709 (I173598,I2683,I405764,I405790,);
DFFARX1 I_23710 (I173592,I2683,I405764,I405807,);
not I_23711 (I405815,I405807);
nor I_23712 (I405732,I405790,I405815);
DFFARX1 I_23713 (I405815,I2683,I405764,I405747,);
nor I_23714 (I405860,I173589,I173580);
and I_23715 (I405877,I405860,I173577);
nor I_23716 (I405894,I405877,I173589);
not I_23717 (I405911,I173589);
and I_23718 (I405928,I405911,I173583);
nand I_23719 (I405945,I405928,I173595);
nor I_23720 (I405962,I405911,I405945);
DFFARX1 I_23721 (I405962,I2683,I405764,I405729,);
not I_23722 (I405993,I405945);
nand I_23723 (I406010,I405815,I405993);
nand I_23724 (I405741,I405877,I405993);
DFFARX1 I_23725 (I405911,I2683,I405764,I405756,);
not I_23726 (I406055,I173601);
nor I_23727 (I406072,I406055,I173583);
nor I_23728 (I406089,I406072,I405894);
DFFARX1 I_23729 (I406089,I2683,I405764,I405753,);
not I_23730 (I406120,I406072);
DFFARX1 I_23731 (I406120,I2683,I405764,I406146,);
not I_23732 (I406154,I406146);
nor I_23733 (I405750,I406154,I406072);
nor I_23734 (I406185,I406055,I173580);
and I_23735 (I406202,I406185,I173586);
or I_23736 (I406219,I406202,I173577);
DFFARX1 I_23737 (I406219,I2683,I405764,I406245,);
not I_23738 (I406253,I406245);
nand I_23739 (I406270,I406253,I405993);
not I_23740 (I405744,I406270);
nand I_23741 (I405738,I406270,I406010);
nand I_23742 (I405735,I406253,I405877);
not I_23743 (I406359,I2690);
DFFARX1 I_23744 (I147023,I2683,I406359,I406385,);
DFFARX1 I_23745 (I147029,I2683,I406359,I406402,);
not I_23746 (I406410,I406402);
nor I_23747 (I406327,I406385,I406410);
DFFARX1 I_23748 (I406410,I2683,I406359,I406342,);
nor I_23749 (I406455,I147038,I147023);
and I_23750 (I406472,I406455,I147050);
nor I_23751 (I406489,I406472,I147038);
not I_23752 (I406506,I147038);
and I_23753 (I406523,I406506,I147026);
nand I_23754 (I406540,I406523,I147047);
nor I_23755 (I406557,I406506,I406540);
DFFARX1 I_23756 (I406557,I2683,I406359,I406324,);
not I_23757 (I406588,I406540);
nand I_23758 (I406605,I406410,I406588);
nand I_23759 (I406336,I406472,I406588);
DFFARX1 I_23760 (I406506,I2683,I406359,I406351,);
not I_23761 (I406650,I147035);
nor I_23762 (I406667,I406650,I147026);
nor I_23763 (I406684,I406667,I406489);
DFFARX1 I_23764 (I406684,I2683,I406359,I406348,);
not I_23765 (I406715,I406667);
DFFARX1 I_23766 (I406715,I2683,I406359,I406741,);
not I_23767 (I406749,I406741);
nor I_23768 (I406345,I406749,I406667);
nor I_23769 (I406780,I406650,I147032);
and I_23770 (I406797,I406780,I147044);
or I_23771 (I406814,I406797,I147041);
DFFARX1 I_23772 (I406814,I2683,I406359,I406840,);
not I_23773 (I406848,I406840);
nand I_23774 (I406865,I406848,I406588);
not I_23775 (I406339,I406865);
nand I_23776 (I406333,I406865,I406605);
nand I_23777 (I406330,I406848,I406472);
not I_23778 (I406954,I2690);
DFFARX1 I_23779 (I291104,I2683,I406954,I406980,);
DFFARX1 I_23780 (I291122,I2683,I406954,I406997,);
not I_23781 (I407005,I406997);
nor I_23782 (I406922,I406980,I407005);
DFFARX1 I_23783 (I407005,I2683,I406954,I406937,);
nor I_23784 (I407050,I291101,I291113);
and I_23785 (I407067,I407050,I291098);
nor I_23786 (I407084,I407067,I291101);
not I_23787 (I407101,I291101);
and I_23788 (I407118,I407101,I291107);
nand I_23789 (I407135,I407118,I291119);
nor I_23790 (I407152,I407101,I407135);
DFFARX1 I_23791 (I407152,I2683,I406954,I406919,);
not I_23792 (I407183,I407135);
nand I_23793 (I407200,I407005,I407183);
nand I_23794 (I406931,I407067,I407183);
DFFARX1 I_23795 (I407101,I2683,I406954,I406946,);
not I_23796 (I407245,I291110);
nor I_23797 (I407262,I407245,I291107);
nor I_23798 (I407279,I407262,I407084);
DFFARX1 I_23799 (I407279,I2683,I406954,I406943,);
not I_23800 (I407310,I407262);
DFFARX1 I_23801 (I407310,I2683,I406954,I407336,);
not I_23802 (I407344,I407336);
nor I_23803 (I406940,I407344,I407262);
nor I_23804 (I407375,I407245,I291098);
and I_23805 (I407392,I407375,I291125);
or I_23806 (I407409,I407392,I291116);
DFFARX1 I_23807 (I407409,I2683,I406954,I407435,);
not I_23808 (I407443,I407435);
nand I_23809 (I407460,I407443,I407183);
not I_23810 (I406934,I407460);
nand I_23811 (I406928,I407460,I407200);
nand I_23812 (I406925,I407443,I407067);
not I_23813 (I407549,I2690);
DFFARX1 I_23814 (I374653,I2683,I407549,I407575,);
DFFARX1 I_23815 (I374656,I2683,I407549,I407592,);
not I_23816 (I407600,I407592);
nor I_23817 (I407517,I407575,I407600);
DFFARX1 I_23818 (I407600,I2683,I407549,I407532,);
nor I_23819 (I407645,I374656,I374671);
and I_23820 (I407662,I407645,I374665);
nor I_23821 (I407679,I407662,I374656);
not I_23822 (I407696,I374656);
and I_23823 (I407713,I407696,I374674);
nand I_23824 (I407730,I407713,I374662);
nor I_23825 (I407747,I407696,I407730);
DFFARX1 I_23826 (I407747,I2683,I407549,I407514,);
not I_23827 (I407778,I407730);
nand I_23828 (I407795,I407600,I407778);
nand I_23829 (I407526,I407662,I407778);
DFFARX1 I_23830 (I407696,I2683,I407549,I407541,);
not I_23831 (I407840,I374668);
nor I_23832 (I407857,I407840,I374674);
nor I_23833 (I407874,I407857,I407679);
DFFARX1 I_23834 (I407874,I2683,I407549,I407538,);
not I_23835 (I407905,I407857);
DFFARX1 I_23836 (I407905,I2683,I407549,I407931,);
not I_23837 (I407939,I407931);
nor I_23838 (I407535,I407939,I407857);
nor I_23839 (I407970,I407840,I374653);
and I_23840 (I407987,I407970,I374677);
or I_23841 (I408004,I407987,I374659);
DFFARX1 I_23842 (I408004,I2683,I407549,I408030,);
not I_23843 (I408038,I408030);
nand I_23844 (I408055,I408038,I407778);
not I_23845 (I407529,I408055);
nand I_23846 (I407523,I408055,I407795);
nand I_23847 (I407520,I408038,I407662);
not I_23848 (I408144,I2690);
DFFARX1 I_23849 (I340622,I2683,I408144,I408170,);
DFFARX1 I_23850 (I340634,I2683,I408144,I408187,);
not I_23851 (I408195,I408187);
nor I_23852 (I408112,I408170,I408195);
DFFARX1 I_23853 (I408195,I2683,I408144,I408127,);
nor I_23854 (I408240,I340631,I340625);
and I_23855 (I408257,I408240,I340619);
nor I_23856 (I408274,I408257,I340631);
not I_23857 (I408291,I340631);
and I_23858 (I408308,I408291,I340628);
nand I_23859 (I408325,I408308,I340619);
nor I_23860 (I408342,I408291,I408325);
DFFARX1 I_23861 (I408342,I2683,I408144,I408109,);
not I_23862 (I408373,I408325);
nand I_23863 (I408390,I408195,I408373);
nand I_23864 (I408121,I408257,I408373);
DFFARX1 I_23865 (I408291,I2683,I408144,I408136,);
not I_23866 (I408435,I340643);
nor I_23867 (I408452,I408435,I340628);
nor I_23868 (I408469,I408452,I408274);
DFFARX1 I_23869 (I408469,I2683,I408144,I408133,);
not I_23870 (I408500,I408452);
DFFARX1 I_23871 (I408500,I2683,I408144,I408526,);
not I_23872 (I408534,I408526);
nor I_23873 (I408130,I408534,I408452);
nor I_23874 (I408565,I408435,I340637);
and I_23875 (I408582,I408565,I340640);
or I_23876 (I408599,I408582,I340622);
DFFARX1 I_23877 (I408599,I2683,I408144,I408625,);
not I_23878 (I408633,I408625);
nand I_23879 (I408650,I408633,I408373);
not I_23880 (I408124,I408650);
nand I_23881 (I408118,I408650,I408390);
nand I_23882 (I408115,I408633,I408257);
not I_23883 (I408739,I2690);
DFFARX1 I_23884 (I373565,I2683,I408739,I408765,);
DFFARX1 I_23885 (I373568,I2683,I408739,I408782,);
not I_23886 (I408790,I408782);
nor I_23887 (I408707,I408765,I408790);
DFFARX1 I_23888 (I408790,I2683,I408739,I408722,);
nor I_23889 (I408835,I373568,I373583);
and I_23890 (I408852,I408835,I373577);
nor I_23891 (I408869,I408852,I373568);
not I_23892 (I408886,I373568);
and I_23893 (I408903,I408886,I373586);
nand I_23894 (I408920,I408903,I373574);
nor I_23895 (I408937,I408886,I408920);
DFFARX1 I_23896 (I408937,I2683,I408739,I408704,);
not I_23897 (I408968,I408920);
nand I_23898 (I408985,I408790,I408968);
nand I_23899 (I408716,I408852,I408968);
DFFARX1 I_23900 (I408886,I2683,I408739,I408731,);
not I_23901 (I409030,I373580);
nor I_23902 (I409047,I409030,I373586);
nor I_23903 (I409064,I409047,I408869);
DFFARX1 I_23904 (I409064,I2683,I408739,I408728,);
not I_23905 (I409095,I409047);
DFFARX1 I_23906 (I409095,I2683,I408739,I409121,);
not I_23907 (I409129,I409121);
nor I_23908 (I408725,I409129,I409047);
nor I_23909 (I409160,I409030,I373565);
and I_23910 (I409177,I409160,I373589);
or I_23911 (I409194,I409177,I373571);
DFFARX1 I_23912 (I409194,I2683,I408739,I409220,);
not I_23913 (I409228,I409220);
nand I_23914 (I409245,I409228,I408968);
not I_23915 (I408719,I409245);
nand I_23916 (I408713,I409245,I408985);
nand I_23917 (I408710,I409228,I408852);
not I_23918 (I409334,I2690);
DFFARX1 I_23919 (I348714,I2683,I409334,I409360,);
DFFARX1 I_23920 (I348726,I2683,I409334,I409377,);
not I_23921 (I409385,I409377);
nor I_23922 (I409302,I409360,I409385);
DFFARX1 I_23923 (I409385,I2683,I409334,I409317,);
nor I_23924 (I409430,I348723,I348717);
and I_23925 (I409447,I409430,I348711);
nor I_23926 (I409464,I409447,I348723);
not I_23927 (I409481,I348723);
and I_23928 (I409498,I409481,I348720);
nand I_23929 (I409515,I409498,I348711);
nor I_23930 (I409532,I409481,I409515);
DFFARX1 I_23931 (I409532,I2683,I409334,I409299,);
not I_23932 (I409563,I409515);
nand I_23933 (I409580,I409385,I409563);
nand I_23934 (I409311,I409447,I409563);
DFFARX1 I_23935 (I409481,I2683,I409334,I409326,);
not I_23936 (I409625,I348735);
nor I_23937 (I409642,I409625,I348720);
nor I_23938 (I409659,I409642,I409464);
DFFARX1 I_23939 (I409659,I2683,I409334,I409323,);
not I_23940 (I409690,I409642);
DFFARX1 I_23941 (I409690,I2683,I409334,I409716,);
not I_23942 (I409724,I409716);
nor I_23943 (I409320,I409724,I409642);
nor I_23944 (I409755,I409625,I348729);
and I_23945 (I409772,I409755,I348732);
or I_23946 (I409789,I409772,I348714);
DFFARX1 I_23947 (I409789,I2683,I409334,I409815,);
not I_23948 (I409823,I409815);
nand I_23949 (I409840,I409823,I409563);
not I_23950 (I409314,I409840);
nand I_23951 (I409308,I409840,I409580);
nand I_23952 (I409305,I409823,I409447);
not I_23953 (I409929,I2690);
DFFARX1 I_23954 (I32566,I2683,I409929,I409955,);
DFFARX1 I_23955 (I32554,I2683,I409929,I409972,);
not I_23956 (I409980,I409972);
nor I_23957 (I409897,I409955,I409980);
DFFARX1 I_23958 (I409980,I2683,I409929,I409912,);
nor I_23959 (I410025,I32545,I32569);
and I_23960 (I410042,I410025,I32548);
nor I_23961 (I410059,I410042,I32545);
not I_23962 (I410076,I32545);
and I_23963 (I410093,I410076,I32551);
nand I_23964 (I410110,I410093,I32563);
nor I_23965 (I410127,I410076,I410110);
DFFARX1 I_23966 (I410127,I2683,I409929,I409894,);
not I_23967 (I410158,I410110);
nand I_23968 (I410175,I409980,I410158);
nand I_23969 (I409906,I410042,I410158);
DFFARX1 I_23970 (I410076,I2683,I409929,I409921,);
not I_23971 (I410220,I32545);
nor I_23972 (I410237,I410220,I32551);
nor I_23973 (I410254,I410237,I410059);
DFFARX1 I_23974 (I410254,I2683,I409929,I409918,);
not I_23975 (I410285,I410237);
DFFARX1 I_23976 (I410285,I2683,I409929,I410311,);
not I_23977 (I410319,I410311);
nor I_23978 (I409915,I410319,I410237);
nor I_23979 (I410350,I410220,I32548);
and I_23980 (I410367,I410350,I32557);
or I_23981 (I410384,I410367,I32560);
DFFARX1 I_23982 (I410384,I2683,I409929,I410410,);
not I_23983 (I410418,I410410);
nand I_23984 (I410435,I410418,I410158);
not I_23985 (I409909,I410435);
nand I_23986 (I409903,I410435,I410175);
nand I_23987 (I409900,I410418,I410042);
not I_23988 (I410524,I2690);
DFFARX1 I_23989 (I60204,I2683,I410524,I410550,);
DFFARX1 I_23990 (I60207,I2683,I410524,I410567,);
not I_23991 (I410575,I410567);
nor I_23992 (I410492,I410550,I410575);
DFFARX1 I_23993 (I410575,I2683,I410524,I410507,);
nor I_23994 (I410620,I60213,I60207);
and I_23995 (I410637,I410620,I60210);
nor I_23996 (I410654,I410637,I60213);
not I_23997 (I410671,I60213);
and I_23998 (I410688,I410671,I60204);
nand I_23999 (I410705,I410688,I60222);
nor I_24000 (I410722,I410671,I410705);
DFFARX1 I_24001 (I410722,I2683,I410524,I410489,);
not I_24002 (I410753,I410705);
nand I_24003 (I410770,I410575,I410753);
nand I_24004 (I410501,I410637,I410753);
DFFARX1 I_24005 (I410671,I2683,I410524,I410516,);
not I_24006 (I410815,I60216);
nor I_24007 (I410832,I410815,I60204);
nor I_24008 (I410849,I410832,I410654);
DFFARX1 I_24009 (I410849,I2683,I410524,I410513,);
not I_24010 (I410880,I410832);
DFFARX1 I_24011 (I410880,I2683,I410524,I410906,);
not I_24012 (I410914,I410906);
nor I_24013 (I410510,I410914,I410832);
nor I_24014 (I410945,I410815,I60219);
and I_24015 (I410962,I410945,I60225);
or I_24016 (I410979,I410962,I60228);
DFFARX1 I_24017 (I410979,I2683,I410524,I411005,);
not I_24018 (I411013,I411005);
nand I_24019 (I411030,I411013,I410753);
not I_24020 (I410504,I411030);
nand I_24021 (I410498,I411030,I410770);
nand I_24022 (I410495,I411013,I410637);
not I_24023 (I411119,I2690);
DFFARX1 I_24024 (I245547,I2683,I411119,I411145,);
DFFARX1 I_24025 (I245544,I2683,I411119,I411162,);
not I_24026 (I411170,I411162);
nor I_24027 (I411087,I411145,I411170);
DFFARX1 I_24028 (I411170,I2683,I411119,I411102,);
nor I_24029 (I411215,I245559,I245541);
and I_24030 (I411232,I411215,I245538);
nor I_24031 (I411249,I411232,I245559);
not I_24032 (I411266,I245559);
and I_24033 (I411283,I411266,I245544);
nand I_24034 (I411300,I411283,I245556);
nor I_24035 (I411317,I411266,I411300);
DFFARX1 I_24036 (I411317,I2683,I411119,I411084,);
not I_24037 (I411348,I411300);
nand I_24038 (I411365,I411170,I411348);
nand I_24039 (I411096,I411232,I411348);
DFFARX1 I_24040 (I411266,I2683,I411119,I411111,);
not I_24041 (I411410,I245550);
nor I_24042 (I411427,I411410,I245544);
nor I_24043 (I411444,I411427,I411249);
DFFARX1 I_24044 (I411444,I2683,I411119,I411108,);
not I_24045 (I411475,I411427);
DFFARX1 I_24046 (I411475,I2683,I411119,I411501,);
not I_24047 (I411509,I411501);
nor I_24048 (I411105,I411509,I411427);
nor I_24049 (I411540,I411410,I245538);
and I_24050 (I411557,I411540,I245553);
or I_24051 (I411574,I411557,I245541);
DFFARX1 I_24052 (I411574,I2683,I411119,I411600,);
not I_24053 (I411608,I411600);
nand I_24054 (I411625,I411608,I411348);
not I_24055 (I411099,I411625);
nand I_24056 (I411093,I411625,I411365);
nand I_24057 (I411090,I411608,I411232);
not I_24058 (I411714,I2690);
DFFARX1 I_24059 (I345246,I2683,I411714,I411740,);
DFFARX1 I_24060 (I345258,I2683,I411714,I411757,);
not I_24061 (I411765,I411757);
nor I_24062 (I411682,I411740,I411765);
DFFARX1 I_24063 (I411765,I2683,I411714,I411697,);
nor I_24064 (I411810,I345255,I345249);
and I_24065 (I411827,I411810,I345243);
nor I_24066 (I411844,I411827,I345255);
not I_24067 (I411861,I345255);
and I_24068 (I411878,I411861,I345252);
nand I_24069 (I411895,I411878,I345243);
nor I_24070 (I411912,I411861,I411895);
DFFARX1 I_24071 (I411912,I2683,I411714,I411679,);
not I_24072 (I411943,I411895);
nand I_24073 (I411960,I411765,I411943);
nand I_24074 (I411691,I411827,I411943);
DFFARX1 I_24075 (I411861,I2683,I411714,I411706,);
not I_24076 (I412005,I345267);
nor I_24077 (I412022,I412005,I345252);
nor I_24078 (I412039,I412022,I411844);
DFFARX1 I_24079 (I412039,I2683,I411714,I411703,);
not I_24080 (I412070,I412022);
DFFARX1 I_24081 (I412070,I2683,I411714,I412096,);
not I_24082 (I412104,I412096);
nor I_24083 (I411700,I412104,I412022);
nor I_24084 (I412135,I412005,I345261);
and I_24085 (I412152,I412135,I345264);
or I_24086 (I412169,I412152,I345246);
DFFARX1 I_24087 (I412169,I2683,I411714,I412195,);
not I_24088 (I412203,I412195);
nand I_24089 (I412220,I412203,I411943);
not I_24090 (I411694,I412220);
nand I_24091 (I411688,I412220,I411960);
nand I_24092 (I411685,I412203,I411827);
not I_24093 (I412309,I2690);
DFFARX1 I_24094 (I1940,I2683,I412309,I412335,);
DFFARX1 I_24095 (I2308,I2683,I412309,I412352,);
not I_24096 (I412360,I412352);
nor I_24097 (I412277,I412335,I412360);
DFFARX1 I_24098 (I412360,I2683,I412309,I412292,);
nor I_24099 (I412405,I2276,I1444);
and I_24100 (I412422,I412405,I2108);
nor I_24101 (I412439,I412422,I2276);
not I_24102 (I412456,I2276);
and I_24103 (I412473,I412456,I2220);
nand I_24104 (I412490,I412473,I1956);
nor I_24105 (I412507,I412456,I412490);
DFFARX1 I_24106 (I412507,I2683,I412309,I412274,);
not I_24107 (I412538,I412490);
nand I_24108 (I412555,I412360,I412538);
nand I_24109 (I412286,I412422,I412538);
DFFARX1 I_24110 (I412456,I2683,I412309,I412301,);
not I_24111 (I412600,I2524);
nor I_24112 (I412617,I412600,I2220);
nor I_24113 (I412634,I412617,I412439);
DFFARX1 I_24114 (I412634,I2683,I412309,I412298,);
not I_24115 (I412665,I412617);
DFFARX1 I_24116 (I412665,I2683,I412309,I412691,);
not I_24117 (I412699,I412691);
nor I_24118 (I412295,I412699,I412617);
nor I_24119 (I412730,I412600,I2324);
and I_24120 (I412747,I412730,I1620);
or I_24121 (I412764,I412747,I2084);
DFFARX1 I_24122 (I412764,I2683,I412309,I412790,);
not I_24123 (I412798,I412790);
nand I_24124 (I412815,I412798,I412538);
not I_24125 (I412289,I412815);
nand I_24126 (I412283,I412815,I412555);
nand I_24127 (I412280,I412798,I412422);
not I_24128 (I412904,I2690);
DFFARX1 I_24129 (I275600,I2683,I412904,I412930,);
DFFARX1 I_24130 (I275618,I2683,I412904,I412947,);
not I_24131 (I412955,I412947);
nor I_24132 (I412872,I412930,I412955);
DFFARX1 I_24133 (I412955,I2683,I412904,I412887,);
nor I_24134 (I413000,I275597,I275609);
and I_24135 (I413017,I413000,I275594);
nor I_24136 (I413034,I413017,I275597);
not I_24137 (I413051,I275597);
and I_24138 (I413068,I413051,I275603);
nand I_24139 (I413085,I413068,I275615);
nor I_24140 (I413102,I413051,I413085);
DFFARX1 I_24141 (I413102,I2683,I412904,I412869,);
not I_24142 (I413133,I413085);
nand I_24143 (I413150,I412955,I413133);
nand I_24144 (I412881,I413017,I413133);
DFFARX1 I_24145 (I413051,I2683,I412904,I412896,);
not I_24146 (I413195,I275606);
nor I_24147 (I413212,I413195,I275603);
nor I_24148 (I413229,I413212,I413034);
DFFARX1 I_24149 (I413229,I2683,I412904,I412893,);
not I_24150 (I413260,I413212);
DFFARX1 I_24151 (I413260,I2683,I412904,I413286,);
not I_24152 (I413294,I413286);
nor I_24153 (I412890,I413294,I413212);
nor I_24154 (I413325,I413195,I275594);
and I_24155 (I413342,I413325,I275621);
or I_24156 (I413359,I413342,I275612);
DFFARX1 I_24157 (I413359,I2683,I412904,I413385,);
not I_24158 (I413393,I413385);
nand I_24159 (I413410,I413393,I413133);
not I_24160 (I412884,I413410);
nand I_24161 (I412878,I413410,I413150);
nand I_24162 (I412875,I413393,I413017);
not I_24163 (I413499,I2690);
DFFARX1 I_24164 (I336576,I2683,I413499,I413525,);
DFFARX1 I_24165 (I336588,I2683,I413499,I413542,);
not I_24166 (I413550,I413542);
nor I_24167 (I413467,I413525,I413550);
DFFARX1 I_24168 (I413550,I2683,I413499,I413482,);
nor I_24169 (I413595,I336585,I336579);
and I_24170 (I413612,I413595,I336573);
nor I_24171 (I413629,I413612,I336585);
not I_24172 (I413646,I336585);
and I_24173 (I413663,I413646,I336582);
nand I_24174 (I413680,I413663,I336573);
nor I_24175 (I413697,I413646,I413680);
DFFARX1 I_24176 (I413697,I2683,I413499,I413464,);
not I_24177 (I413728,I413680);
nand I_24178 (I413745,I413550,I413728);
nand I_24179 (I413476,I413612,I413728);
DFFARX1 I_24180 (I413646,I2683,I413499,I413491,);
not I_24181 (I413790,I336597);
nor I_24182 (I413807,I413790,I336582);
nor I_24183 (I413824,I413807,I413629);
DFFARX1 I_24184 (I413824,I2683,I413499,I413488,);
not I_24185 (I413855,I413807);
DFFARX1 I_24186 (I413855,I2683,I413499,I413881,);
not I_24187 (I413889,I413881);
nor I_24188 (I413485,I413889,I413807);
nor I_24189 (I413920,I413790,I336591);
and I_24190 (I413937,I413920,I336594);
or I_24191 (I413954,I413937,I336576);
DFFARX1 I_24192 (I413954,I2683,I413499,I413980,);
not I_24193 (I413988,I413980);
nand I_24194 (I414005,I413988,I413728);
not I_24195 (I413479,I414005);
nand I_24196 (I413473,I414005,I413745);
nand I_24197 (I413470,I413988,I413612);
not I_24198 (I414094,I2690);
DFFARX1 I_24199 (I64964,I2683,I414094,I414120,);
DFFARX1 I_24200 (I64967,I2683,I414094,I414137,);
not I_24201 (I414145,I414137);
nor I_24202 (I414062,I414120,I414145);
DFFARX1 I_24203 (I414145,I2683,I414094,I414077,);
nor I_24204 (I414190,I64973,I64967);
and I_24205 (I414207,I414190,I64970);
nor I_24206 (I414224,I414207,I64973);
not I_24207 (I414241,I64973);
and I_24208 (I414258,I414241,I64964);
nand I_24209 (I414275,I414258,I64982);
nor I_24210 (I414292,I414241,I414275);
DFFARX1 I_24211 (I414292,I2683,I414094,I414059,);
not I_24212 (I414323,I414275);
nand I_24213 (I414340,I414145,I414323);
nand I_24214 (I414071,I414207,I414323);
DFFARX1 I_24215 (I414241,I2683,I414094,I414086,);
not I_24216 (I414385,I64976);
nor I_24217 (I414402,I414385,I64964);
nor I_24218 (I414419,I414402,I414224);
DFFARX1 I_24219 (I414419,I2683,I414094,I414083,);
not I_24220 (I414450,I414402);
DFFARX1 I_24221 (I414450,I2683,I414094,I414476,);
not I_24222 (I414484,I414476);
nor I_24223 (I414080,I414484,I414402);
nor I_24224 (I414515,I414385,I64979);
and I_24225 (I414532,I414515,I64985);
or I_24226 (I414549,I414532,I64988);
DFFARX1 I_24227 (I414549,I2683,I414094,I414575,);
not I_24228 (I414583,I414575);
nand I_24229 (I414600,I414583,I414323);
not I_24230 (I414074,I414600);
nand I_24231 (I414068,I414600,I414340);
nand I_24232 (I414065,I414583,I414207);
not I_24233 (I414689,I2690);
DFFARX1 I_24234 (I262411,I2683,I414689,I414715,);
DFFARX1 I_24235 (I262408,I2683,I414689,I414732,);
not I_24236 (I414740,I414732);
nor I_24237 (I414657,I414715,I414740);
DFFARX1 I_24238 (I414740,I2683,I414689,I414672,);
nor I_24239 (I414785,I262423,I262405);
and I_24240 (I414802,I414785,I262402);
nor I_24241 (I414819,I414802,I262423);
not I_24242 (I414836,I262423);
and I_24243 (I414853,I414836,I262408);
nand I_24244 (I414870,I414853,I262420);
nor I_24245 (I414887,I414836,I414870);
DFFARX1 I_24246 (I414887,I2683,I414689,I414654,);
not I_24247 (I414918,I414870);
nand I_24248 (I414935,I414740,I414918);
nand I_24249 (I414666,I414802,I414918);
DFFARX1 I_24250 (I414836,I2683,I414689,I414681,);
not I_24251 (I414980,I262414);
nor I_24252 (I414997,I414980,I262408);
nor I_24253 (I415014,I414997,I414819);
DFFARX1 I_24254 (I415014,I2683,I414689,I414678,);
not I_24255 (I415045,I414997);
DFFARX1 I_24256 (I415045,I2683,I414689,I415071,);
not I_24257 (I415079,I415071);
nor I_24258 (I414675,I415079,I414997);
nor I_24259 (I415110,I414980,I262402);
and I_24260 (I415127,I415110,I262417);
or I_24261 (I415144,I415127,I262405);
DFFARX1 I_24262 (I415144,I2683,I414689,I415170,);
not I_24263 (I415178,I415170);
nand I_24264 (I415195,I415178,I414918);
not I_24265 (I414669,I415195);
nand I_24266 (I414663,I415195,I414935);
nand I_24267 (I414660,I415178,I414802);
not I_24268 (I415284,I2690);
DFFARX1 I_24269 (I220416,I2683,I415284,I415310,);
DFFARX1 I_24270 (I220398,I2683,I415284,I415327,);
not I_24271 (I415335,I415327);
nor I_24272 (I415252,I415310,I415335);
DFFARX1 I_24273 (I415335,I2683,I415284,I415267,);
nor I_24274 (I415380,I220404,I220407);
and I_24275 (I415397,I415380,I220395);
nor I_24276 (I415414,I415397,I220404);
not I_24277 (I415431,I220404);
and I_24278 (I415448,I415431,I220413);
nand I_24279 (I415465,I415448,I220401);
nor I_24280 (I415482,I415431,I415465);
DFFARX1 I_24281 (I415482,I2683,I415284,I415249,);
not I_24282 (I415513,I415465);
nand I_24283 (I415530,I415335,I415513);
nand I_24284 (I415261,I415397,I415513);
DFFARX1 I_24285 (I415431,I2683,I415284,I415276,);
not I_24286 (I415575,I220398);
nor I_24287 (I415592,I415575,I220413);
nor I_24288 (I415609,I415592,I415414);
DFFARX1 I_24289 (I415609,I2683,I415284,I415273,);
not I_24290 (I415640,I415592);
DFFARX1 I_24291 (I415640,I2683,I415284,I415666,);
not I_24292 (I415674,I415666);
nor I_24293 (I415270,I415674,I415592);
nor I_24294 (I415705,I415575,I220410);
and I_24295 (I415722,I415705,I220419);
or I_24296 (I415739,I415722,I220395);
DFFARX1 I_24297 (I415739,I2683,I415284,I415765,);
not I_24298 (I415773,I415765);
nand I_24299 (I415790,I415773,I415513);
not I_24300 (I415264,I415790);
nand I_24301 (I415258,I415790,I415530);
nand I_24302 (I415255,I415773,I415397);
not I_24303 (I415879,I2690);
DFFARX1 I_24304 (I328484,I2683,I415879,I415905,);
DFFARX1 I_24305 (I328496,I2683,I415879,I415922,);
not I_24306 (I415930,I415922);
nor I_24307 (I415847,I415905,I415930);
DFFARX1 I_24308 (I415930,I2683,I415879,I415862,);
nor I_24309 (I415975,I328493,I328487);
and I_24310 (I415992,I415975,I328481);
nor I_24311 (I416009,I415992,I328493);
not I_24312 (I416026,I328493);
and I_24313 (I416043,I416026,I328490);
nand I_24314 (I416060,I416043,I328481);
nor I_24315 (I416077,I416026,I416060);
DFFARX1 I_24316 (I416077,I2683,I415879,I415844,);
not I_24317 (I416108,I416060);
nand I_24318 (I416125,I415930,I416108);
nand I_24319 (I415856,I415992,I416108);
DFFARX1 I_24320 (I416026,I2683,I415879,I415871,);
not I_24321 (I416170,I328505);
nor I_24322 (I416187,I416170,I328490);
nor I_24323 (I416204,I416187,I416009);
DFFARX1 I_24324 (I416204,I2683,I415879,I415868,);
not I_24325 (I416235,I416187);
DFFARX1 I_24326 (I416235,I2683,I415879,I416261,);
not I_24327 (I416269,I416261);
nor I_24328 (I415865,I416269,I416187);
nor I_24329 (I416300,I416170,I328499);
and I_24330 (I416317,I416300,I328502);
or I_24331 (I416334,I416317,I328484);
DFFARX1 I_24332 (I416334,I2683,I415879,I416360,);
not I_24333 (I416368,I416360);
nand I_24334 (I416385,I416368,I416108);
not I_24335 (I415859,I416385);
nand I_24336 (I415853,I416385,I416125);
nand I_24337 (I415850,I416368,I415992);
not I_24338 (I416474,I2690);
DFFARX1 I_24339 (I312088,I2683,I416474,I416500,);
DFFARX1 I_24340 (I312079,I2683,I416474,I416517,);
not I_24341 (I416525,I416517);
nor I_24342 (I416442,I416500,I416525);
DFFARX1 I_24343 (I416525,I2683,I416474,I416457,);
nor I_24344 (I416570,I312085,I312094);
and I_24345 (I416587,I416570,I312097);
nor I_24346 (I416604,I416587,I312085);
not I_24347 (I416621,I312085);
and I_24348 (I416638,I416621,I312076);
nand I_24349 (I416655,I416638,I312082);
nor I_24350 (I416672,I416621,I416655);
DFFARX1 I_24351 (I416672,I2683,I416474,I416439,);
not I_24352 (I416703,I416655);
nand I_24353 (I416720,I416525,I416703);
nand I_24354 (I416451,I416587,I416703);
DFFARX1 I_24355 (I416621,I2683,I416474,I416466,);
not I_24356 (I416765,I312091);
nor I_24357 (I416782,I416765,I312076);
nor I_24358 (I416799,I416782,I416604);
DFFARX1 I_24359 (I416799,I2683,I416474,I416463,);
not I_24360 (I416830,I416782);
DFFARX1 I_24361 (I416830,I2683,I416474,I416856,);
not I_24362 (I416864,I416856);
nor I_24363 (I416460,I416864,I416782);
nor I_24364 (I416895,I416765,I312076);
and I_24365 (I416912,I416895,I312079);
or I_24366 (I416929,I416912,I312082);
DFFARX1 I_24367 (I416929,I2683,I416474,I416955,);
not I_24368 (I416963,I416955);
nand I_24369 (I416980,I416963,I416703);
not I_24370 (I416454,I416980);
nand I_24371 (I416448,I416980,I416720);
nand I_24372 (I416445,I416963,I416587);
not I_24373 (I417069,I2690);
DFFARX1 I_24374 (I234288,I2683,I417069,I417095,);
DFFARX1 I_24375 (I234270,I2683,I417069,I417112,);
not I_24376 (I417120,I417112);
nor I_24377 (I417037,I417095,I417120);
DFFARX1 I_24378 (I417120,I2683,I417069,I417052,);
nor I_24379 (I417165,I234276,I234279);
and I_24380 (I417182,I417165,I234267);
nor I_24381 (I417199,I417182,I234276);
not I_24382 (I417216,I234276);
and I_24383 (I417233,I417216,I234285);
nand I_24384 (I417250,I417233,I234273);
nor I_24385 (I417267,I417216,I417250);
DFFARX1 I_24386 (I417267,I2683,I417069,I417034,);
not I_24387 (I417298,I417250);
nand I_24388 (I417315,I417120,I417298);
nand I_24389 (I417046,I417182,I417298);
DFFARX1 I_24390 (I417216,I2683,I417069,I417061,);
not I_24391 (I417360,I234270);
nor I_24392 (I417377,I417360,I234285);
nor I_24393 (I417394,I417377,I417199);
DFFARX1 I_24394 (I417394,I2683,I417069,I417058,);
not I_24395 (I417425,I417377);
DFFARX1 I_24396 (I417425,I2683,I417069,I417451,);
not I_24397 (I417459,I417451);
nor I_24398 (I417055,I417459,I417377);
nor I_24399 (I417490,I417360,I234282);
and I_24400 (I417507,I417490,I234291);
or I_24401 (I417524,I417507,I234267);
DFFARX1 I_24402 (I417524,I2683,I417069,I417550,);
not I_24403 (I417558,I417550);
nand I_24404 (I417575,I417558,I417298);
not I_24405 (I417049,I417575);
nand I_24406 (I417043,I417575,I417315);
nand I_24407 (I417040,I417558,I417182);
not I_24408 (I417664,I2690);
DFFARX1 I_24409 (I76864,I2683,I417664,I417690,);
DFFARX1 I_24410 (I76867,I2683,I417664,I417707,);
not I_24411 (I417715,I417707);
nor I_24412 (I417632,I417690,I417715);
DFFARX1 I_24413 (I417715,I2683,I417664,I417647,);
nor I_24414 (I417760,I76873,I76867);
and I_24415 (I417777,I417760,I76870);
nor I_24416 (I417794,I417777,I76873);
not I_24417 (I417811,I76873);
and I_24418 (I417828,I417811,I76864);
nand I_24419 (I417845,I417828,I76882);
nor I_24420 (I417862,I417811,I417845);
DFFARX1 I_24421 (I417862,I2683,I417664,I417629,);
not I_24422 (I417893,I417845);
nand I_24423 (I417910,I417715,I417893);
nand I_24424 (I417641,I417777,I417893);
DFFARX1 I_24425 (I417811,I2683,I417664,I417656,);
not I_24426 (I417955,I76876);
nor I_24427 (I417972,I417955,I76864);
nor I_24428 (I417989,I417972,I417794);
DFFARX1 I_24429 (I417989,I2683,I417664,I417653,);
not I_24430 (I418020,I417972);
DFFARX1 I_24431 (I418020,I2683,I417664,I418046,);
not I_24432 (I418054,I418046);
nor I_24433 (I417650,I418054,I417972);
nor I_24434 (I418085,I417955,I76879);
and I_24435 (I418102,I418085,I76885);
or I_24436 (I418119,I418102,I76888);
DFFARX1 I_24437 (I418119,I2683,I417664,I418145,);
not I_24438 (I418153,I418145);
nand I_24439 (I418170,I418153,I417893);
not I_24440 (I417644,I418170);
nand I_24441 (I417638,I418170,I417910);
nand I_24442 (I417635,I418153,I417777);
not I_24443 (I418259,I2690);
DFFARX1 I_24444 (I137775,I2683,I418259,I418285,);
DFFARX1 I_24445 (I137781,I2683,I418259,I418302,);
not I_24446 (I418310,I418302);
nor I_24447 (I418227,I418285,I418310);
DFFARX1 I_24448 (I418310,I2683,I418259,I418242,);
nor I_24449 (I418355,I137790,I137775);
and I_24450 (I418372,I418355,I137802);
nor I_24451 (I418389,I418372,I137790);
not I_24452 (I418406,I137790);
and I_24453 (I418423,I418406,I137778);
nand I_24454 (I418440,I418423,I137799);
nor I_24455 (I418457,I418406,I418440);
DFFARX1 I_24456 (I418457,I2683,I418259,I418224,);
not I_24457 (I418488,I418440);
nand I_24458 (I418505,I418310,I418488);
nand I_24459 (I418236,I418372,I418488);
DFFARX1 I_24460 (I418406,I2683,I418259,I418251,);
not I_24461 (I418550,I137787);
nor I_24462 (I418567,I418550,I137778);
nor I_24463 (I418584,I418567,I418389);
DFFARX1 I_24464 (I418584,I2683,I418259,I418248,);
not I_24465 (I418615,I418567);
DFFARX1 I_24466 (I418615,I2683,I418259,I418641,);
not I_24467 (I418649,I418641);
nor I_24468 (I418245,I418649,I418567);
nor I_24469 (I418680,I418550,I137784);
and I_24470 (I418697,I418680,I137796);
or I_24471 (I418714,I418697,I137793);
DFFARX1 I_24472 (I418714,I2683,I418259,I418740,);
not I_24473 (I418748,I418740);
nand I_24474 (I418765,I418748,I418488);
not I_24475 (I418239,I418765);
nand I_24476 (I418233,I418765,I418505);
nand I_24477 (I418230,I418748,I418372);
not I_24478 (I418854,I2690);
DFFARX1 I_24479 (I356806,I2683,I418854,I418880,);
DFFARX1 I_24480 (I356818,I2683,I418854,I418897,);
not I_24481 (I418905,I418897);
nor I_24482 (I418822,I418880,I418905);
DFFARX1 I_24483 (I418905,I2683,I418854,I418837,);
nor I_24484 (I418950,I356815,I356809);
and I_24485 (I418967,I418950,I356803);
nor I_24486 (I418984,I418967,I356815);
not I_24487 (I419001,I356815);
and I_24488 (I419018,I419001,I356812);
nand I_24489 (I419035,I419018,I356803);
nor I_24490 (I419052,I419001,I419035);
DFFARX1 I_24491 (I419052,I2683,I418854,I418819,);
not I_24492 (I419083,I419035);
nand I_24493 (I419100,I418905,I419083);
nand I_24494 (I418831,I418967,I419083);
DFFARX1 I_24495 (I419001,I2683,I418854,I418846,);
not I_24496 (I419145,I356827);
nor I_24497 (I419162,I419145,I356812);
nor I_24498 (I419179,I419162,I418984);
DFFARX1 I_24499 (I419179,I2683,I418854,I418843,);
not I_24500 (I419210,I419162);
DFFARX1 I_24501 (I419210,I2683,I418854,I419236,);
not I_24502 (I419244,I419236);
nor I_24503 (I418840,I419244,I419162);
nor I_24504 (I419275,I419145,I356821);
and I_24505 (I419292,I419275,I356824);
or I_24506 (I419309,I419292,I356806);
DFFARX1 I_24507 (I419309,I2683,I418854,I419335,);
not I_24508 (I419343,I419335);
nand I_24509 (I419360,I419343,I419083);
not I_24510 (I418834,I419360);
nand I_24511 (I418828,I419360,I419100);
nand I_24512 (I418825,I419343,I418967);
not I_24513 (I419449,I2690);
DFFARX1 I_24514 (I297564,I2683,I419449,I419475,);
DFFARX1 I_24515 (I297582,I2683,I419449,I419492,);
not I_24516 (I419500,I419492);
nor I_24517 (I419417,I419475,I419500);
DFFARX1 I_24518 (I419500,I2683,I419449,I419432,);
nor I_24519 (I419545,I297561,I297573);
and I_24520 (I419562,I419545,I297558);
nor I_24521 (I419579,I419562,I297561);
not I_24522 (I419596,I297561);
and I_24523 (I419613,I419596,I297567);
nand I_24524 (I419630,I419613,I297579);
nor I_24525 (I419647,I419596,I419630);
DFFARX1 I_24526 (I419647,I2683,I419449,I419414,);
not I_24527 (I419678,I419630);
nand I_24528 (I419695,I419500,I419678);
nand I_24529 (I419426,I419562,I419678);
DFFARX1 I_24530 (I419596,I2683,I419449,I419441,);
not I_24531 (I419740,I297570);
nor I_24532 (I419757,I419740,I297567);
nor I_24533 (I419774,I419757,I419579);
DFFARX1 I_24534 (I419774,I2683,I419449,I419438,);
not I_24535 (I419805,I419757);
DFFARX1 I_24536 (I419805,I2683,I419449,I419831,);
not I_24537 (I419839,I419831);
nor I_24538 (I419435,I419839,I419757);
nor I_24539 (I419870,I419740,I297558);
and I_24540 (I419887,I419870,I297585);
or I_24541 (I419904,I419887,I297576);
DFFARX1 I_24542 (I419904,I2683,I419449,I419930,);
not I_24543 (I419938,I419930);
nand I_24544 (I419955,I419938,I419678);
not I_24545 (I419429,I419955);
nand I_24546 (I419423,I419955,I419695);
nand I_24547 (I419420,I419938,I419562);
endmodule


