module test_I2311(I1231,I1287,I2311);
input I1231,I1287;
output I2311;
wire I2294;
not I_0(I2311,I2294);
nor I_1(I2294,I1287,I1231);
endmodule


