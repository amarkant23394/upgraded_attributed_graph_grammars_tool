module test_I7410(I3368,I1477,I1470,I7410);
input I3368,I1477,I1470;
output I7410;
wire I5594,I6907,I5512,I5082,I5105;
DFFARX1 I_0(I5512,I1470,I5105,,,I5594,);
not I_1(I6907,I1477);
DFFARX1 I_2(I5082,I1470,I6907,,,I7410,);
DFFARX1 I_3(I3368,I1470,I5105,,,I5512,);
not I_4(I5082,I5594);
not I_5(I5105,I1477);
endmodule


