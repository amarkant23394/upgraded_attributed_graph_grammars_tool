module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_7_r_12,n8_12,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_7_r_12,n8_12,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
nor I_40(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_41(N1508_0_r_12,n30_12,n37_12);
nor I_42(N1507_6_r_12,n25_12,n39_12);
nor I_43(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_44(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_45(n_572_7_r_12,n23_12,n24_12);
nand I_46(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_47(n_549_7_r_12,n27_12,n28_12);
nand I_48(n_569_7_r_12,n25_12,n26_12);
nand I_49(n_452_7_r_12,N1508_1_r_8,N1507_6_r_8);
nand I_50(N6147_9_r_12,n30_12,n31_12);
nor I_51(N6134_9_r_12,n35_12,n36_12);
not I_52(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_53(n1_12,n_573_7_r_12);
not I_54(n8_12,blif_reset_net_7_r_12);
not I_55(n23_12,n36_12);
nor I_56(n24_12,n_452_7_r_12,N1371_0_r_8);
nand I_57(n25_12,n23_12,n40_12);
not I_58(n26_12,n35_12);
not I_59(n27_12,N6134_9_r_12);
nand I_60(n28_12,n26_12,n29_12);
not I_61(n29_12,n24_12);
nand I_62(n30_12,n33_12,n41_12);
nand I_63(n31_12,n32_12,n33_12);
nor I_64(n32_12,n26_12,n34_12);
nor I_65(n33_12,N1508_6_r_8,N1508_10_r_8);
nor I_66(n34_12,n42_12,N6134_9_r_8);
nor I_67(n35_12,n38_12,N1507_6_r_8);
nand I_68(n36_12,G199_8_r_8,n_42_8_r_8);
nand I_69(n37_12,n23_12,n35_12);
or I_70(n38_12,N6147_9_r_8,N1508_6_r_8);
not I_71(n39_12,n30_12);
or I_72(n40_12,N1371_0_r_8,N6147_9_r_8);
nor I_73(n41_12,n34_12,n36_12);
nor I_74(n42_12,n_42_8_r_8,G199_8_r_8);
endmodule


