module test_I15519(I12930,I15047,I1477,I1470,I15519);
input I12930,I15047,I1477,I1470;
output I15519;
wire I12602,I13023,I12605,I12947,I15064,I15389,I15406,I12587,I14965,I15423,I15372,I15485,I15502;
not I_0(I12602,I12930);
DFFARX1 I_1(I1470,,,I13023,);
nand I_2(I12605,I13023,I12947);
nor I_3(I12947,I12930);
nand I_4(I15064,I15047,I12587);
not I_5(I15389,I15372);
nor I_6(I15406,I15064,I15389);
DFFARX1 I_7(I1470,,,I12587,);
or I_8(I15519,I15502,I15423);
not I_9(I14965,I1477);
and I_10(I15423,I15372,I15406);
DFFARX1 I_11(I12602,I1470,I14965,,,I15372,);
DFFARX1 I_12(I12605,I1470,I14965,,,I15485,);
not I_13(I15502,I15485);
endmodule


