module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_7_r_1,n9_1,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
and I_34(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_35(N1508_0_r_1,n40_1,n44_1);
nor I_36(N1507_6_r_1,n43_1,n49_1);
nor I_37(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_38(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_39(n_572_7_r_1,n29_1,n30_1);
not I_40(n_573_7_r_1,n_452_7_r_1);
nor I_41(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_42(n_569_7_r_1,n30_1,n31_1);
nor I_43(n_452_7_r_1,n30_1,n32_1);
nor I_44(N6147_9_r_1,n35_1,n36_1);
nand I_45(N6134_9_r_1,n38_1,n39_1);
not I_46(I_BUFF_1_9_r_1,n40_1);
nor I_47(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_48(n9_1,blif_reset_net_7_r_1);
nor I_49(n29_1,n34_1,N1507_6_r_12);
nor I_50(n30_1,n33_1,n34_1);
nor I_51(n31_1,n54_1,n_572_7_r_12);
not I_52(n32_1,n48_1);
nor I_53(n33_1,n_572_7_r_12,N1507_6_r_12);
not I_54(n34_1,n_569_7_r_12);
nor I_55(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_56(n36_1,n29_1);
not I_57(n37_1,n41_1);
nand I_58(n38_1,I_BUFF_1_9_r_1,N1508_6_r_12);
nand I_59(n39_1,n37_1,n40_1);
nand I_60(n40_1,N1371_0_r_12,N1508_0_r_12);
nand I_61(n41_1,n52_1,N6147_9_r_12);
or I_62(n42_1,n36_1,n43_1);
nor I_63(n43_1,n32_1,n49_1);
nand I_64(n44_1,n45_1,n46_1);
nand I_65(n45_1,n47_1,n48_1);
not I_66(n46_1,N1508_6_r_12);
not I_67(n47_1,n31_1);
nand I_68(n48_1,n50_1,n_549_7_r_12);
nor I_69(n49_1,n41_1,n47_1);
and I_70(n50_1,n51_1,G42_7_r_12);
nand I_71(n51_1,n52_1,n53_1);
nand I_72(n52_1,G42_7_r_12,N1508_0_r_12);
not I_73(n53_1,N6147_9_r_12);
or I_74(n54_1,N1508_6_r_12,N1371_0_r_12);
nor I_75(n55_1,n29_1,N1508_6_r_12);
endmodule


