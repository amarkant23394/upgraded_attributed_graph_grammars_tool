module test_I11525(I6992,I6893,I1470,I8862,I9258,I6887,I7057,I11525);
input I6992,I6893,I1470,I8862,I9258,I6887,I7057;
output I11525;
wire I9320,I8824,I11491,I11508,I8827,I8842,I8981,I9303,I6881,I8879,I9083,I8964;
not I_0(I9320,I9303);
nand I_1(I8824,I9083,I8981);
not I_2(I11491,I8827);
nor I_3(I11508,I11491,I8842);
DFFARX1 I_4(I9258,I1470,I8862,,,I8827,);
nor I_5(I8842,I9320,I9083);
and I_6(I11525,I11508,I8824);
not I_7(I8981,I8964);
DFFARX1 I_8(I1470,I8862,,,I9303,);
nand I_9(I6881,I6992,I7057);
not I_10(I8879,I6887);
nand I_11(I9083,I8879,I6881);
not I_12(I8964,I6893);
endmodule


