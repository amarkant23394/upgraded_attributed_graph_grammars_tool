module test_I9015(I1477,I7427,I7026,I1470,I5097,I6924,I9015);
input I1477,I7427,I7026,I1470,I5097,I6924;
output I9015;
wire I8998,I6992,I6975,I7461,I5088,I7057,I6881,I6907,I7221,I6899,I7444;
not I_0(I8998,I6881);
nand I_1(I6992,I6975,I5097);
nor I_2(I6975,I6924);
and I_3(I7461,I7221,I7444);
DFFARX1 I_4(I1470,,,I5088,);
not I_5(I7057,I7026);
nor I_6(I9015,I8998,I6899);
nand I_7(I6881,I6992,I7057);
not I_8(I6907,I1477);
nand I_9(I7221,I6924,I5088);
DFFARX1 I_10(I7461,I1470,I6907,,,I6899,);
nand I_11(I7444,I7427,I6992);
endmodule


