module test_I1937(I1301,I1937);
input I1301;
output I1937;
wire ;
not I_0(I1937,I1301);
endmodule


