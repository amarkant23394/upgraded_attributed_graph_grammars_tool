module test_I11641(I1477,I9148,I8913,I8851,I11525,I1470,I11641);
input I1477,I9148,I8913,I8851,I11525,I1470;
output I11641;
wire I8830,I9179,I11559,I11412,I8827,I11395,I11624,I11576,I11542,I8862,I9258,I11378,I8833,I9227,I11327,I11310;
nand I_0(I8830,I8913,I9227);
DFFARX1 I_1(I1470,I8862,,,I9179,);
DFFARX1 I_2(I11542,I1470,I11310,,,I11559,);
and I_3(I11641,I11624,I11576);
not I_4(I11412,I11395);
DFFARX1 I_5(I9258,I1470,I8862,,,I8827,);
nand I_6(I11395,I11378,I8851);
nand I_7(I11624,I11327,I8827);
nor I_8(I11576,I11559,I11412);
or I_9(I11542,I11525,I8833);
not I_10(I8862,I1477);
or I_11(I9258,I9179,I9148);
nor I_12(I11378,I11327);
not I_13(I8833,I9179);
nor I_14(I9227,I9179);
not I_15(I11327,I8830);
not I_16(I11310,I1477);
endmodule


