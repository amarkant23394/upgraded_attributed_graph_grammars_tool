module test_I15245(I12930,I1477,I15160,I1470,I15245);
input I12930,I1477,I15160,I1470;
output I15245;
wire I12670,I12783,I12584,I13023,I15109,I12608,I15177,I15194,I12593,I15126,I15211,I14965;
DFFARX1 I_0(I1470,,,I12670,);
DFFARX1 I_1(I1470,,,I12783,);
and I_2(I12584,I12670,I12783);
DFFARX1 I_3(I1470,,,I13023,);
not I_4(I15109,I12584);
nor I_5(I12608,I13023,I12930);
and I_6(I15177,I15160,I12593);
or I_7(I15194,I15177,I12608);
nand I_8(I12593,I12670);
not I_9(I15126,I15109);
DFFARX1 I_10(I15194,I1470,I14965,,,I15211,);
not I_11(I14965,I1477);
nor I_12(I15245,I15211,I15126);
endmodule


