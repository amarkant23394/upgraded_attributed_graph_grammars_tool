module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_7_r_3,n10_3,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_7_r_3,n10_3,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
not I_40(N1372_1_r_3,n40_3);
nor I_41(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_42(N1507_6_r_3,n31_3,n42_3);
nor I_43(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_44(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_45(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_46(n_573_7_r_3,n30_3,n31_3);
nor I_47(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_48(n_569_7_r_3,n30_3,n32_3);
nor I_49(n_452_7_r_3,n35_3,G199_8_r_8);
not I_50(N6147_9_r_3,n32_3);
nor I_51(N6134_9_r_3,n36_3,n37_3);
not I_52(I_BUFF_1_9_r_3,n45_3);
nor I_53(n4_7_r_3,I_BUFF_1_9_r_3,G199_8_r_8);
not I_54(n10_3,blif_reset_net_7_r_3);
not I_55(n30_3,n39_3);
not I_56(n31_3,n35_3);
nand I_57(n32_3,n41_3,N1508_1_r_8);
nor I_58(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_59(n34_3,n46_3,N1371_0_r_8);
nor I_60(n35_3,n43_3,n44_3);
not I_61(n36_3,n34_3);
nor I_62(n37_3,N6147_9_r_3,G199_8_r_8);
or I_63(n38_3,n_572_7_r_3,n34_3);
nor I_64(n39_3,n44_3,n_42_8_r_8);
nand I_65(n40_3,n39_3,G199_8_r_8);
nand I_66(n41_3,N1508_1_r_8,N1508_10_r_8);
nor I_67(n42_3,n34_3,n45_3);
not I_68(n43_3,N6147_9_r_8);
nor I_69(n44_3,N1507_6_r_8,N1508_6_r_8);
nand I_70(n45_3,n49_3,n50_3);
and I_71(n46_3,n47_3,n_42_8_r_8);
nand I_72(n47_3,n41_3,n48_3);
not I_73(n48_3,N1508_1_r_8);
nor I_74(n49_3,N1371_0_r_8,G199_8_r_8);
or I_75(n50_3,n51_3,N1508_6_r_8);
nor I_76(n51_3,N6134_9_r_8,N1507_6_r_8);
endmodule


