module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_14,blif_reset_net_1_r_14,G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_14,blif_reset_net_1_r_14;
output G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n_452_1_r_14,n4_1_l_14,n3_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_14,n3_14,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_14,n3_14,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_14,n3_14,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_14,n3_14,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_14,n3_14,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_14,n3_14,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n_452_1_r_14,blif_clk_net_1_r_14,n3_14,G42_1_r_14,);
and I_35(n_572_1_r_14,n18_14,n19_14);
nand I_36(n_573_1_r_14,n16_14,n17_14);
nor I_37(n_549_1_r_14,n20_14,n21_14);
or I_38(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_39(n_452_1_r_14,n23_14,n_573_1_r_4);
nor I_40(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_41(N3_2_r_14,blif_clk_net_1_r_14,n3_14,G199_2_r_14,);
DFFARX1 I_42(n_572_1_l_14,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_14,);
not I_43(P6_5_r_14,P6_5_r_internal_14);
nor I_44(n4_1_l_14,n_572_1_r_4,ACVQN2_3_r_4);
not I_45(n3_14,blif_reset_net_1_r_14);
DFFARX1 I_46(n4_1_l_14,blif_clk_net_1_r_14,n3_14,n15_internal_14,);
not I_47(n15_14,n15_internal_14);
DFFARX1 I_48(ACVQN1_5_r_4,blif_clk_net_1_r_14,n3_14,ACVQN2_3_l_14,);
DFFARX1 I_49(n_549_1_r_4,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_14,);
and I_50(N3_2_r_14,n26_14,n27_14);
nor I_51(n_572_1_l_14,n_266_and_0_3_r_4,n_572_1_r_4);
DFFARX1 I_52(ACVQN2_3_l_14,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_14,);
nor I_53(n16_14,n_573_1_r_4,G42_1_r_4);
not I_54(n17_14,n_572_1_l_14);
nor I_55(n18_14,n_569_1_r_4,G42_1_r_4);
nand I_56(n19_14,ACVQN1_3_l_14,P6_5_r_4);
nor I_57(n20_14,n_572_1_r_4,n_569_1_r_4);
nor I_58(n21_14,n15_14,n22_14);
nand I_59(n22_14,n24_14,n25_14);
nand I_60(n23_14,n15_14,n24_14);
not I_61(n24_14,G42_1_r_4);
not I_62(n25_14,n_569_1_r_4);
nor I_63(n26_14,n20_14,n_573_1_r_4);
nand I_64(n27_14,n28_14,G42_1_r_4);
not I_65(n28_14,n_266_and_0_3_r_4);
endmodule


