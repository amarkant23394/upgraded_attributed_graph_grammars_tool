module test_I11009(I8205,I1477,I1470,I8193,I11009);
input I8205,I1477,I1470,I8193;
output I11009;
wire I10647,I9491,I9816,I9468,I9621,I9864;
not I_0(I10647,I1477);
not I_1(I9491,I1477);
DFFARX1 I_2(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_3(I9864,I1470,I9491,,,I9468,);
DFFARX1 I_4(I9468,I1470,I10647,,,I11009,);
DFFARX1 I_5(I8205,I1470,I9491,,,I9621,);
nor I_6(I9864,I9816,I9621);
endmodule


