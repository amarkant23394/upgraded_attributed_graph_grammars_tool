module test_I7556(I1477,I7782,I6459,I6306,I6843,I1470,I3957,I7556);
input I1477,I7782,I6459,I6306,I6843,I1470,I3957;
output I7556;
wire I6781,I7816,I7850,I6380,I6315,I6294,I6297,I6476,I7621,I6329,I7731,I7714,I6541,I7799,I7570,I7604;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
DFFARX1 I_1(I7799,I1470,I7570,,,I7816,);
nor I_2(I7850,I7816,I7731);
DFFARX1 I_3(I1470,I6329,,,I6380,);
nand I_4(I6315,I6781,I6476);
and I_5(I6294,I6380,I6541);
DFFARX1 I_6(I6843,I1470,I6329,,,I6297,);
nor I_7(I6476,I6380,I6459);
nand I_8(I7621,I7604,I6315);
not I_9(I6329,I1477);
not I_10(I7731,I7714);
not I_11(I7714,I6297);
DFFARX1 I_12(I1470,I6329,,,I6541,);
nand I_13(I7556,I7621,I7850);
or I_14(I7799,I7782,I6306);
not I_15(I7570,I1477);
nor I_16(I7604,I6297,I6294);
endmodule


