module test_I8592(I1477,I4533,I1470,I8592);
input I1477,I4533,I1470;
output I8592;
wire I8527,I8233,I8216,I5751,I5713,I6028,I6110,I6127,I5722;
nand I_0(I8527,I8233,I5713);
not I_1(I8233,I5722);
not I_2(I8216,I1477);
not I_3(I5751,I1477);
DFFARX1 I_4(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_5(I1470,I5751,,,I6028,);
DFFARX1 I_6(I1470,I5751,,,I6110,);
DFFARX1 I_7(I8527,I1470,I8216,,,I8592,);
and I_8(I6127,I6110,I4533);
DFFARX1 I_9(I6028,I1470,I5751,,,I5722,);
endmodule


