module test_I12425(I7556,I10086,I1477,I7731,I1470,I12425);
input I7556,I10086,I1477,I7731,I1470;
output I12425;
wire I10349,I7550,I10038,I10538,I7532,I7977,I11973,I10490,I10052,I10103,I10332;
and I_0(I10349,I10332,I7550);
nand I_1(I7550,I7977,I7731);
nand I_2(I10038,I10349,I10538);
DFFARX1 I_3(I10038,I1470,I11973,,,I12425,);
nor I_4(I10538,I10490,I10103);
DFFARX1 I_5(I1470,,,I7532,);
DFFARX1 I_6(I1470,,,I7977,);
not I_7(I11973,I1477);
DFFARX1 I_8(I7556,I1470,I10052,,,I10490,);
not I_9(I10052,I1477);
DFFARX1 I_10(I10086,I1470,I10052,,,I10103,);
DFFARX1 I_11(I7532,I1470,I10052,,,I10332,);
endmodule


