module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,n_102_5_r_0,n_452_7_r_0,n_431_5_r_0,n6_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_5_r_0,n6_0,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_36(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_37(n_429_or_0_5_r_0,n38_0,N1508_6_r_4);
DFFARX1 I_38(n_431_5_r_0,blif_clk_net_5_r_0,n6_0,G78_5_r_0,);
nand I_39(n_576_5_r_0,n26_0,N1508_6_r_4);
not I_40(n_102_5_r_0,n27_0);
nand I_41(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_42(n4_7_r_0,blif_clk_net_5_r_0,n6_0,G42_7_r_0,);
nor I_43(n_572_7_r_0,n31_0,N1508_6_r_4);
or I_44(n_573_7_r_0,n29_0,n30_0);
nor I_45(n_549_7_r_0,n29_0,n33_0);
nand I_46(n_569_7_r_0,n28_0,n32_0);
nor I_47(n_452_7_r_0,n30_0,n31_0);
nand I_48(n_431_5_r_0,n_102_5_r_0,n35_0);
not I_49(n6_0,blif_reset_net_5_r_0);
nor I_50(n4_7_r_0,n31_0,n37_0);
nor I_51(n26_0,n27_0,n28_0);
nor I_52(n27_0,n28_0,n44_0);
nand I_53(n28_0,G42_7_r_4,n_569_7_r_4);
not I_54(n29_0,n32_0);
nor I_55(n30_0,n39_0,N1371_0_r_4);
not I_56(n31_0,n38_0);
nand I_57(n32_0,n41_0,n42_0);
nor I_58(n33_0,n_102_5_r_0,N1508_6_r_4);
nor I_59(n34_0,n27_0,N1508_6_r_4);
nand I_60(n35_0,n29_0,n36_0);
nor I_61(n36_0,n37_0,n38_0);
not I_62(n37_0,n28_0);
nand I_63(n38_0,n40_0,n_452_7_r_4);
nor I_64(n39_0,n_572_7_r_4,n_549_7_r_4);
or I_65(n40_0,n_572_7_r_4,n_549_7_r_4);
nor I_66(n41_0,N1371_0_r_4,N1507_6_r_4);
or I_67(n42_0,n43_0,G42_7_r_4);
nor I_68(n43_0,N6134_9_r_4,N1508_6_r_4);
nor I_69(n44_0,n45_0,N1507_6_r_4);
and I_70(n45_0,n_549_7_r_4,n_569_7_r_4);
endmodule


