module test_I14066(I10349,I10120,I1477,I1470,I11990,I14066);
input I10349,I10120,I1477,I1470,I11990;
output I14066;
wire I12270,I11956,I10014,I12349,I10041,I14049,I13775,I11973,I11962;
nand I_0(I12270,I11990,I10014);
not I_1(I11956,I12349);
DFFARX1 I_2(I1470,,,I10014,);
DFFARX1 I_3(I10041,I1470,I11973,,,I12349,);
nor I_4(I10041,I10349,I10120);
DFFARX1 I_5(I11962,I1470,I13775,,,I14049,);
not I_6(I13775,I1477);
not I_7(I11973,I1477);
nor I_8(I11962,I12349,I12270);
and I_9(I14066,I14049,I11956);
endmodule


