module test_I9621(I8233,I1477,I1470,I9621);
input I8233,I1477,I1470;
output I9621;
wire I8298,I5719,I5802,I8205,I5740,I8315,I9491;
nor I_0(I8298,I8233,I5719);
DFFARX1 I_1(I1470,,,I5719,);
DFFARX1 I_2(I1470,,,I5802,);
not I_3(I8205,I8315);
DFFARX1 I_4(I8205,I1470,I9491,,,I9621,);
not I_5(I5740,I5802);
nand I_6(I8315,I8298,I5740);
not I_7(I9491,I1477);
endmodule


