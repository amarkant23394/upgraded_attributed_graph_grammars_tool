module test_I13159(I11429,I1477,I1470,I11689,I11751,I13159);
input I11429,I1477,I1470,I11689,I11751;
output I13159;
wire I11559,I11296,I13197,I11768,I11272,I13508,I13491,I11310;
DFFARX1 I_0(I1470,I11310,,,I11559,);
nand I_1(I11296,I11559,I11689);
not I_2(I13197,I1477);
and I_3(I11768,I11429,I11751);
DFFARX1 I_4(I11768,I1470,I11310,,,I11272,);
and I_5(I13508,I13491,I11272);
DFFARX1 I_6(I11296,I1470,I13197,,,I13491,);
not I_7(I11310,I1477);
DFFARX1 I_8(I13508,I1470,I13197,,,I13159,);
endmodule


