module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_5,blif_reset_net_5_r_5,N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_5,blif_reset_net_5_r_5;
output N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5;
wire N1371_0_r_2,N1508_0_r_2,N6147_3_r_2,n_429_or_0_5_r_2,G78_5_r_2,n_576_5_r_2,n_102_5_r_2,n_547_5_r_2,N1372_10_r_2,N1508_10_r_2,n_431_5_r_2,n21_2,n22_2,n23_2,n24_2,n25_2,n26_2,n27_2,n28_2,n29_2,n30_2,n31_2,n32_2,N1508_0_r_5,N1507_6_r_5,n_431_5_r_5,n6_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5;
nor I_0(N1371_0_r_2,n23_2,n24_2);
not I_1(N1508_0_r_2,n24_2);
nor I_2(N6147_3_r_2,n22_2,n26_2);
nand I_3(n_429_or_0_5_r_2,IN_3_1_l_2,n22_2);
DFFARX1 I_4(n_431_5_r_2,blif_clk_net_5_r_5,n6_5,G78_5_r_2,);
nand I_5(n_576_5_r_2,n21_2,n22_2);
not I_6(n_102_5_r_2,n23_2);
nand I_7(n_547_5_r_2,n22_2,n24_2);
not I_8(N1372_10_r_2,n29_2);
nor I_9(N1508_10_r_2,n28_2,n29_2);
nand I_10(n_431_5_r_2,n_102_5_r_2,n25_2);
nor I_11(n21_2,IN_3_1_l_2,n23_2);
and I_12(n22_2,IN_1_1_l_2,IN_2_1_l_2);
nor I_13(n23_2,n24_2,n31_2);
nand I_14(n24_2,IN_1_4_l_2,IN_2_4_l_2);
nand I_15(n25_2,n26_2,n27_2);
nor I_16(n26_2,IN_1_3_l_2,n30_2);
not I_17(n27_2,n_429_or_0_5_r_2);
nor I_18(n28_2,n22_2,n23_2);
nand I_19(n29_2,N1508_0_r_2,n26_2);
or I_20(n30_2,IN_2_3_l_2,IN_3_3_l_2);
nor I_21(n31_2,IN_5_4_l_2,n32_2);
and I_22(n32_2,IN_3_4_l_2,IN_4_4_l_2);
nor I_23(N1371_0_r_5,n28_5,n39_5);
not I_24(N1508_0_r_5,n39_5);
nor I_25(N6147_2_r_5,n28_5,n37_5);
nand I_26(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_27(n_431_5_r_5,blif_clk_net_5_r_5,n6_5,G78_5_r_5,);
nand I_28(n_576_5_r_5,n26_5,n27_5);
not I_29(n_102_5_r_5,n28_5);
nand I_30(n_547_5_r_5,n31_5,n32_5);
nor I_31(N1507_6_r_5,n30_5,n32_5);
nor I_32(N1508_6_r_5,n39_5,n41_5);
nand I_33(n_431_5_r_5,n34_5,n35_5);
not I_34(n6_5,blif_reset_net_5_r_5);
nor I_35(n26_5,n29_5,n30_5);
nor I_36(n27_5,n28_5,N1371_0_r_2);
nor I_37(n28_5,n29_5,n44_5);
not I_38(n29_5,n_547_5_r_2);
nand I_39(n30_5,N1508_0_r_5,n43_5);
nor I_40(n31_5,n28_5,n33_5);
nor I_41(n32_5,n40_5,G78_5_r_2);
nor I_42(n33_5,n29_5,N1371_0_r_2);
or I_43(n34_5,n29_5,N1371_0_r_2);
nand I_44(n35_5,n32_5,n36_5);
not I_45(n36_5,n30_5);
nor I_46(n37_5,N1507_6_r_5,n38_5);
and I_47(n38_5,n39_5,n40_5);
nand I_48(n39_5,n_576_5_r_2,n_547_5_r_2);
nand I_49(n40_5,N1508_10_r_2,N1371_0_r_2);
nand I_50(n41_5,n28_5,n42_5);
or I_51(n42_5,n32_5,n36_5);
or I_52(n43_5,N6147_3_r_2,N1372_10_r_2);
nor I_53(n44_5,N6147_3_r_2,G78_5_r_2);
endmodule


