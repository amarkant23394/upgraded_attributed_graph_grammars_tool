module test_I6924(I1477,I5122,I1470,I6924);
input I1477,I5122,I1470;
output I6924;
wire I5416,I5450,I5351,I5073,I5433,I3356,I5105;
nand I_0(I5416,I5122,I3356);
and I_1(I5450,I5416,I5433);
DFFARX1 I_2(I1470,I5105,,,I5351,);
DFFARX1 I_3(I5450,I1470,I5105,,,I5073,);
nand I_4(I5433,I5416,I5351);
DFFARX1 I_5(I1470,,,I3356,);
not I_6(I5105,I1477);
not I_7(I6924,I5073);
endmodule


