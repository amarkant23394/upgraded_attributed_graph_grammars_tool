module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_17,n6_17,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_17,n6_17,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_17,n6_17,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_17,n6_17,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_17,n6_17,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_34(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_35(n_573_1_r_17,n20_17,n21_17);
nand I_36(n_549_1_r_17,n23_17,n24_17);
nand I_37(n_569_1_r_17,n21_17,n22_17);
not I_38(n_452_1_r_17,n23_17);
DFFARX1 I_39(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_40(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_41(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_42(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_43(n_431_0_l_17,n26_17,n_572_1_r_13);
not I_44(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_45(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_46(n20_17,n20_internal_17);
DFFARX1 I_47(n_572_1_r_13,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_48(ACVQN2_3_r_13,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_49(n19_17,n19_internal_17);
nor I_50(n4_1_r_17,n5_17,n25_17);
not I_51(n2_17,n29_17);
DFFARX1 I_52(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_53(n17_17,n17_internal_17);
nor I_54(N1_4_r_17,n29_17,n31_17);
not I_55(n5_17,n_452_1_r_13);
and I_56(n21_17,n32_17,G42_1_r_13);
not I_57(n22_17,n25_17);
nand I_58(n23_17,n20_17,n22_17);
nand I_59(n24_17,n19_17,n22_17);
nand I_60(n25_17,n30_17,G42_1_r_13);
and I_61(n26_17,n27_17,ACVQN1_5_r_13);
nor I_62(n27_17,n28_17,n_266_and_0_3_r_13);
not I_63(n28_17,P6_5_r_13);
nor I_64(n29_17,n28_17,n_549_1_r_13);
and I_65(n30_17,n5_17,n_549_1_r_13);
nor I_66(n31_17,n21_17,n_452_1_r_13);
nor I_67(n32_17,n_573_1_r_13,n_452_1_r_13);
endmodule


