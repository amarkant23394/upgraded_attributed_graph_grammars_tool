module test_I13891(I1477,I12041,I1470,I10026,I13891);
input I1477,I12041,I1470,I10026;
output I13891;
wire I13775,I12058,I11973,I12075,I11944;
DFFARX1 I_0(I11944,I1470,I13775,,,I13891,);
not I_1(I13775,I1477);
nand I_2(I12058,I12041,I10026);
not I_3(I11973,I1477);
DFFARX1 I_4(I12058,I1470,I11973,,,I12075,);
not I_5(I11944,I12075);
endmodule


