module test_I6907(I1477,I6907);
input I1477;
output I6907;
wire ;
not I_0(I6907,I1477);
endmodule


