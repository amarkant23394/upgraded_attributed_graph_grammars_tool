module test_I2832(I2764,I1294,I1301,I2832);
input I2764,I1294,I1301;
output I2832;
wire I2172,I2815,I2798,I1917,I2781,I2583,I1899,I1905,I1937,I2313,I2505,I2389,I2406,I2488;
DFFARX1 I_0(I1294,I1937,,,I2172,);
or I_1(I2815,I2798,I1917);
and I_2(I2798,I2781,I1899);
nand I_3(I1917,I2406,I2505);
nor I_4(I2781,I2764,I1905);
not I_5(I2583,I1301);
DFFARX1 I_6(I2172,I1294,I1937,,,I1899,);
DFFARX1 I_7(I2172,I1294,I1937,,,I1905,);
not I_8(I1937,I1301);
DFFARX1 I_9(I1294,I1937,,,I2313,);
nor I_10(I2505,I2313,I2488);
DFFARX1 I_11(I1294,I1937,,,I2389,);
not I_12(I2406,I2389);
DFFARX1 I_13(I2815,I1294,I2583,,,I2832,);
not I_14(I2488,I2406);
endmodule


