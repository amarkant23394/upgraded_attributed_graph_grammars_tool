module test_I5785(I2167,I1477,I4708,I2161,I2173,I1470,I2158,I5785);
input I2167,I1477,I4708,I2161,I2173,I1470,I2158;
output I5785;
wire I4629,I4595,I4544,I4524,I4869,I2143,I4561,I4886,I5768,I4530,I4578,I4807,I4515,I4742,I4725,I4824,I4612;
nor I_0(I4629,I2167,I2173);
DFFARX1 I_1(I4578,I1470,I4544,,,I4595,);
not I_2(I4544,I1477);
nor I_3(I4524,I4742,I4595);
DFFARX1 I_4(I1470,I4544,,,I4869,);
and I_5(I5785,I5768,I4524);
DFFARX1 I_6(I1470,,,I2143,);
nand I_7(I4561,I2173);
and I_8(I4886,I4869,I4612);
nand I_9(I5768,I4530,I4515);
nor I_10(I4530,I4824,I4886);
and I_11(I4578,I4561,I2161);
DFFARX1 I_12(I1470,I4544,,,I4807,);
not I_13(I4515,I4629);
DFFARX1 I_14(I4725,I1470,I4544,,,I4742,);
and I_15(I4725,I4708,I2158);
and I_16(I4824,I4807,I2143);
not I_17(I4612,I4595);
endmodule


