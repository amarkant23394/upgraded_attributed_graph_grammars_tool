module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_8_r_10,n11_10,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_8_r_10,n11_10,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
nor I_37(N1371_0_r_10,n37_10,n38_10);
nor I_38(N1508_0_r_10,n37_10,n58_10);
nand I_39(N6147_2_r_10,n39_10,n40_10);
not I_40(N6147_3_r_10,n39_10);
nor I_41(N1372_4_r_10,n46_10,n49_10);
nor I_42(N1508_4_r_10,n51_10,n52_10);
nor I_43(N1507_6_r_10,n49_10,n60_10);
nor I_44(N1508_6_r_10,n49_10,n50_10);
nor I_45(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_46(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_47(N6147_9_r_10,n36_10,n37_10);
nor I_48(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_49(I_BUFF_1_9_r_10,n48_10);
nor I_50(N3_8_r_10,n44_10,n47_10);
not I_51(n11_10,blif_reset_net_8_r_10);
not I_52(n35_10,n49_10);
nor I_53(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_54(n37_10,n_452_7_r_14);
not I_55(n38_10,n46_10);
nand I_56(n39_10,n43_10,n44_10);
nand I_57(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_58(n41_10,n42_10,n_452_7_r_14);
not I_59(n42_10,n44_10);
nor I_60(n43_10,n45_10,n_452_7_r_14);
nand I_61(n44_10,n54_10,N1507_6_r_14);
nor I_62(n45_10,n59_10,N1371_0_r_14);
nand I_63(n46_10,n61_10,n_573_7_r_14);
nor I_64(n47_10,n46_10,n48_10);
nand I_65(n48_10,n62_10,n63_10);
nand I_66(n49_10,n56_10,G42_7_r_14);
not I_67(n50_10,n45_10);
nor I_68(n51_10,n42_10,n53_10);
not I_69(n52_10,N1372_4_r_10);
nor I_70(n53_10,n48_10,n50_10);
and I_71(n54_10,n55_10,N1508_0_r_14);
nand I_72(n55_10,n56_10,n57_10);
nand I_73(n56_10,N1371_0_r_14,N1508_6_r_14);
not I_74(n57_10,G42_7_r_14);
nor I_75(n58_10,n35_10,n45_10);
nor I_76(n59_10,N1508_0_r_14,N1507_6_r_14);
nor I_77(n60_10,n37_10,n46_10);
or I_78(n61_10,N1508_0_r_14,N1507_6_r_14);
nor I_79(n62_10,n_549_7_r_14,N6134_9_r_14);
or I_80(n63_10,n64_10,n_569_7_r_14);
nor I_81(n64_10,n_572_7_r_14,N6147_9_r_14);
endmodule


