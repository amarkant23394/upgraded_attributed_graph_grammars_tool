module test_final(IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_5,blif_reset_net_5_r_5,N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5);
input IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_5_r_5,blif_reset_net_5_r_5;
output N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5;
wire N1371_0_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_102_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4,n_431_5_r_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,N1508_0_r_5,N1507_6_r_5,n_431_5_r_5,n6_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5;
nor I_0(N1371_0_r_4,n25_4,n29_4);
nor I_1(N1508_0_r_4,n25_4,n32_4);
nor I_2(N6147_2_r_4,n24_4,n31_4);
or I_3(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_4(n_431_5_r_4,blif_clk_net_5_r_5,n6_5,G78_5_r_4,);
nand I_5(n_576_5_r_4,n22_4,n23_4);
nand I_6(n_102_5_r_4,n34_4,n35_4);
nand I_7(n_547_5_r_4,n26_4,n27_4);
nor I_8(N1507_6_r_4,n27_4,n30_4);
nor I_9(N1508_6_r_4,n30_4,n33_4);
nand I_10(n_431_5_r_4,n_102_5_r_4,n28_4);
nor I_11(n22_4,n24_4,n25_4);
nor I_12(n23_4,IN_1_3_l_4,n37_4);
not I_13(n24_4,n_102_5_r_4);
nand I_14(n25_4,IN_1_1_l_4,IN_2_1_l_4);
nor I_15(n26_4,n23_4,n24_4);
not I_16(n27_4,n25_4);
nand I_17(n28_4,n23_4,n29_4);
nor I_18(n29_4,IN_3_1_l_4,n25_4);
not I_19(n30_4,n29_4);
nor I_20(n31_4,N1371_0_r_4,n32_4);
nor I_21(n32_4,n23_4,n29_4);
nand I_22(n33_4,n23_4,n24_4);
nor I_23(n34_4,IN_1_2_l_4,IN_2_2_l_4);
or I_24(n35_4,IN_5_2_l_4,n36_4);
nor I_25(n36_4,IN_3_2_l_4,IN_4_2_l_4);
or I_26(n37_4,IN_2_3_l_4,IN_3_3_l_4);
nor I_27(N1371_0_r_5,n28_5,n39_5);
not I_28(N1508_0_r_5,n39_5);
nor I_29(N6147_2_r_5,n28_5,n37_5);
nand I_30(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_31(n_431_5_r_5,blif_clk_net_5_r_5,n6_5,G78_5_r_5,);
nand I_32(n_576_5_r_5,n26_5,n27_5);
not I_33(n_102_5_r_5,n28_5);
nand I_34(n_547_5_r_5,n31_5,n32_5);
nor I_35(N1507_6_r_5,n30_5,n32_5);
nor I_36(N1508_6_r_5,n39_5,n41_5);
nand I_37(n_431_5_r_5,n34_5,n35_5);
not I_38(n6_5,blif_reset_net_5_r_5);
nor I_39(n26_5,n29_5,n30_5);
nor I_40(n27_5,n28_5,n_547_5_r_4);
nor I_41(n28_5,n29_5,n44_5);
not I_42(n29_5,N1507_6_r_4);
nand I_43(n30_5,N1508_0_r_5,n43_5);
nor I_44(n31_5,n28_5,n33_5);
nor I_45(n32_5,n40_5,N6147_2_r_4);
nor I_46(n33_5,n29_5,n_547_5_r_4);
or I_47(n34_5,n29_5,n_547_5_r_4);
nand I_48(n35_5,n32_5,n36_5);
not I_49(n36_5,n30_5);
nor I_50(n37_5,N1507_6_r_5,n38_5);
and I_51(n38_5,n39_5,n40_5);
nand I_52(n39_5,G78_5_r_4,N1508_0_r_4);
nand I_53(n40_5,N1508_0_r_4,n_429_or_0_5_r_4);
nand I_54(n41_5,n28_5,n42_5);
or I_55(n42_5,n32_5,n36_5);
or I_56(n43_5,n_576_5_r_4,N1508_6_r_4);
nor I_57(n44_5,N6147_2_r_4,n_429_or_0_5_r_4);
endmodule


