module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_5_r_9,n10_9,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
nor I_44(N6147_2_r_9,n62_9,n46_9);
not I_45(N1372_4_r_9,n59_9);
nor I_46(N1508_4_r_9,n58_9,n59_9);
nand I_47(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_48(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_49(n_576_5_r_9,n39_9,n40_9);
not I_50(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_51(n_547_5_r_9,n43_9,N6134_9_r_10);
and I_52(n_42_8_r_9,n44_9,N6147_3_r_10);
DFFARX1 I_53(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_54(N6147_9_r_9,n41_9,n45_9);
nor I_55(N6134_9_r_9,n45_9,n51_9);
nor I_56(I_BUFF_1_9_r_9,n41_9,N6134_9_r_10);
nor I_57(n4_7_l_9,N6147_2_r_10,N6147_3_r_10);
not I_58(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_59(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_60(N3_8_l_9,n57_9,N1508_4_r_10);
DFFARX1 I_61(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_62(n38_9,n63_9);
nor I_63(n_431_5_r_9,N6147_3_r_10,N1507_6_r_10);
nor I_64(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_65(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_66(n40_9,n41_9);
nand I_67(n41_9,N1371_0_r_10,N1508_0_r_10);
nor I_68(n42_9,N1508_0_r_10,N1508_6_r_10);
nor I_69(n43_9,n63_9,n41_9);
nor I_70(n44_9,N1508_6_r_10,n_42_8_r_10);
and I_71(n45_9,n52_9,N6147_9_r_10);
nor I_72(n46_9,n47_9,n48_9);
nor I_73(n47_9,n49_9,n50_9);
not I_74(n48_9,n_429_or_0_5_r_9);
not I_75(n49_9,n42_9);
or I_76(n50_9,n63_9,n51_9);
nor I_77(n51_9,N6147_2_r_10,N1371_0_r_10);
nor I_78(n52_9,n49_9,N6147_3_r_10);
nor I_79(n53_9,n54_9,n55_9);
nor I_80(n54_9,n56_9,N6147_3_r_10);
or I_81(n55_9,n44_9,N1508_0_r_10);
not I_82(n56_9,N6147_9_r_10);
nand I_83(n57_9,N6147_2_r_10,G199_8_r_10);
nor I_84(n58_9,n62_9,n60_9);
nand I_85(n59_9,n51_9,n61_9);
nor I_86(n60_9,n38_9,n44_9);
nor I_87(n61_9,n_42_8_r_10,N6147_3_r_10);
endmodule


