module test_I11944(I1477,I10397,I1470,I11990,I11944);
input I1477,I10397,I1470,I11990;
output I11944;
wire I10219,I12041,I10020,I12058,I11973,I12075,I10026;
DFFARX1 I_0(I1470,,,I10219,);
nor I_1(I12041,I11990,I10020);
DFFARX1 I_2(I1470,,,I10020,);
nand I_3(I12058,I12041,I10026);
not I_4(I11973,I1477);
DFFARX1 I_5(I12058,I1470,I11973,,,I12075,);
nand I_6(I10026,I10219,I10397);
not I_7(I11944,I12075);
endmodule


