module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_0,n6_0,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_0,n6_0,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_0,n6_0,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_0,n6_0,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_0,n6_0,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_0,n6_0,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_0,n6_0,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_0,n6_0,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_31(n_572_1_r_0,n23_0,G199_2_r_10);
nand I_32(n_573_1_r_0,n21_0,n22_0);
nand I_33(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_34(n_569_1_r_0,n21_0,n26_0);
nor I_35(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_36(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_37(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_38(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_39(n4_1_l_0,G42_1_r_10,n_572_1_r_10);
not I_40(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_41(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_42(G42_1_r_10,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_43(n20_0,n38_0);
DFFARX1 I_44(n_549_1_r_10,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_45(n4_1_r_0,n23_0,n_42_2_r_10);
nor I_46(N3_2_r_0,n31_0,n32_0);
nor I_47(N1_4_r_0,n29_0,n32_0);
not I_48(n2_0,n31_0);
nor I_49(n21_0,n37_0,ACVQN2_3_r_10);
not I_50(n22_0,G199_2_r_10);
nand I_51(n23_0,n20_0,n30_0);
nand I_52(n24_0,n38_0,n25_0);
nor I_53(n25_0,n_42_2_r_10,ACVQN2_3_r_10);
not I_54(n26_0,n_42_2_r_10);
not I_55(n27_0,n29_0);
nor I_56(n28_0,n_572_1_r_10,n_573_1_r_10);
nand I_57(n29_0,n26_0,n33_0);
not I_58(n30_0,ACVQN2_3_r_10);
nand I_59(n31_0,ACVQN1_3_l_0,n_573_1_r_10);
and I_60(n32_0,n35_0,n36_0);
nand I_61(n33_0,n34_0,n_266_and_0_3_r_10);
not I_62(n34_0,n_573_1_r_10);
nor I_63(n35_0,n_573_1_r_10,n_572_1_r_10);
nor I_64(n36_0,n_572_1_r_10,G199_2_r_10);
endmodule


