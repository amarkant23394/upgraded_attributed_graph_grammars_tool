module test_I13758(I12041,I1477,I10026,I1470,I12024,I12106,I13758);
input I12041,I1477,I10026,I1470,I12024,I12106;
output I13758;
wire I12287,I12304,I12349,I12058,I13843,I11973,I11965,I12380,I11959;
nand I_0(I12287,I12024);
and I_1(I12304,I12106,I12287);
DFFARX1 I_2(I1470,I11973,,,I12349,);
nand I_3(I12058,I12041,I10026);
nor I_4(I13843,I11959,I11965);
not I_5(I11973,I1477);
DFFARX1 I_6(I12304,I1470,I11973,,,I11965,);
nor I_7(I12380,I12349,I12024);
not I_8(I13758,I13843);
nand I_9(I11959,I12058,I12380);
endmodule


