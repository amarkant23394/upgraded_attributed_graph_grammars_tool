module test_I16740(I1477,I16452,I13162,I14777,I14472,I1470,I16740);
input I1477,I16452,I13162,I14777,I14472,I1470;
output I16740;
wire I14338,I16339,I16291,I16469,I16644,I14605,I16486,I14537,I14808,I14370,I16723,I14347,I16240,I14353,I16308;
DFFARX1 I_0(I14605,I1470,I14370,,,I14338,);
nor I_1(I16339,I14353,I14338);
DFFARX1 I_2(I1470,I16240,,,I16291,);
DFFARX1 I_3(I16452,I1470,I16240,,,I16469,);
DFFARX1 I_4(I14347,I1470,I16240,,,I16644,);
and I_5(I14605,I14537,I14472);
or I_6(I16740,I16339,I16723);
nor I_7(I16486,I16469,I16308);
DFFARX1 I_8(I1470,I14370,,,I14537,);
DFFARX1 I_9(I13162,I1470,I14370,,,I14808,);
not I_10(I14370,I1477);
and I_11(I16723,I16644,I16486);
DFFARX1 I_12(I14777,I1470,I14370,,,I14347,);
not I_13(I16240,I1477);
not I_14(I14353,I14808);
not I_15(I16308,I16291);
endmodule


