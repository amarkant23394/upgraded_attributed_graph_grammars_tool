module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_5_r_11,n9_11,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_5_r_11,n9_11,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
not I_40(N1372_1_r_11,n53_11);
nor I_41(N1508_1_r_11,n39_11,n53_11);
nor I_42(N6147_2_r_11,n48_11,n49_11);
nor I_43(N6147_3_r_11,n44_11,n45_11);
nand I_44(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_45(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_46(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_47(n_102_5_r_11,n39_11);
nand I_48(n_547_5_r_11,n36_11,n37_11);
nor I_49(N1507_6_r_11,n52_11,n57_11);
nor I_50(N1508_6_r_11,n46_11,n51_11);
nor I_51(N1372_10_r_11,n43_11,n47_11);
nor I_52(N1508_10_r_11,n55_11,n56_11);
nand I_53(n_431_5_r_11,n40_11,n41_11);
not I_54(n9_11,blif_reset_net_5_r_11);
nor I_55(n36_11,n38_11,n39_11);
not I_56(n37_11,n40_11);
nor I_57(n38_11,n60_11,N1371_0_r_16);
nor I_58(n39_11,n54_11,n_572_7_r_16);
nand I_59(n40_11,N6147_2_r_16,n_569_7_r_16);
nand I_60(n41_11,n_102_5_r_11,n42_11);
and I_61(n42_11,n58_11,n_452_7_r_16);
not I_62(n43_11,n44_11);
nor I_63(n44_11,n40_11,N1508_0_r_16);
nand I_64(n45_11,n46_11,n47_11);
not I_65(n46_11,n38_11);
nand I_66(n47_11,n59_11,n62_11);
and I_67(n48_11,n37_11,n47_11);
or I_68(n49_11,n44_11,n50_11);
nor I_69(n50_11,n60_11,n61_11);
or I_70(n51_11,n_102_5_r_11,n52_11);
nor I_71(n52_11,n42_11,n57_11);
nand I_72(n53_11,n37_11,n50_11);
or I_73(n54_11,N1507_6_r_16,N1508_0_r_16);
nor I_74(n55_11,n38_11,n42_11);
not I_75(n56_11,N1372_10_r_11);
and I_76(n57_11,n38_11,n50_11);
and I_77(n58_11,n59_11,G42_7_r_16);
or I_78(n59_11,n63_11,N1372_1_r_16);
not I_79(n60_11,N1508_1_r_16);
nor I_80(n61_11,N1508_6_r_16,n_573_7_r_16);
nand I_81(n62_11,N1371_0_r_16,N1372_1_r_16);
and I_82(n63_11,N1371_0_r_16,N1372_1_r_16);
endmodule


