module test_I9833(I9508,I1477,I1470,I9833);
input I9508,I1477,I1470;
output I9833;
wire I9542,I8216,I8623,I9816,I9559,I8705,I8184,I9525,I8193,I9491;
DFFARX1 I_0(I9525,I1470,I9491,,,I9542,);
not I_1(I8216,I1477);
DFFARX1 I_2(I1470,I8216,,,I8623,);
DFFARX1 I_3(I8193,I1470,I9491,,,I9816,);
not I_4(I9559,I9542);
DFFARX1 I_5(I8623,I1470,I8216,,,I8705,);
DFFARX1 I_6(I1470,I8216,,,I8184,);
and I_7(I9525,I9508,I8184);
and I_8(I9833,I9816,I9559);
not I_9(I8193,I8705);
not I_10(I9491,I1477);
endmodule


