module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_9,n5_9,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_9,n5_9,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_9,n5_9,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_9,n5_9,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_9,n5_9,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_9,n5_9,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_9,n5_9,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_9,n5_9,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_33(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_34(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_35(n_549_1_r_9,n17_9,n18_9);
or I_36(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_37(n_452_1_r_9,n26_9,n25_9);
nor I_38(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_39(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_40(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_41(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_42(N3_2_l_9,n22_9,G199_4_r_16);
not I_43(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_44(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_45(n16_9,n27_9);
DFFARX1 I_46(ACVQN1_5_r_16,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_47(n15_9,n26_9);
DFFARX1 I_48(G42_1_r_16,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_49(n29_9,n29_internal_9);
and I_50(N1_4_l_9,n24_9,n_569_1_r_16);
DFFARX1 I_51(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_52(n_573_1_r_16,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_53(n28_9,n28_internal_9);
nor I_54(n4_1_r_9,n27_9,n26_9);
nor I_55(N3_2_r_9,n15_9,n21_9);
nor I_56(N1_4_r_9,n16_9,n21_9);
nor I_57(n_42_2_l_9,n_452_1_r_16,P6_5_r_16);
not I_58(n17_9,n_452_1_r_9);
nand I_59(n18_9,n27_9,n15_9);
nor I_60(n19_9,n29_9,n20_9);
not I_61(n20_9,n_572_1_r_16);
and I_62(n21_9,n23_9,n_572_1_r_16);
nand I_63(n22_9,G42_1_r_16,P6_5_r_16);
nor I_64(n23_9,n29_9,n28_9);
nand I_65(n24_9,n_549_1_r_16,G214_4_r_16);
endmodule


