module test_I17390(I17430,I17515,I1477,I15603,I1470,I17390);
input I17430,I17515,I1477,I15603,I1470;
output I17390;
wire I17413,I17916,I17744,I15576,I17998,I17679,I17933,I17727,I17662;
not I_0(I17413,I1477);
DFFARX1 I_1(I15603,I1470,I17413,,,I17916,);
DFFARX1 I_2(I17998,I1470,I17413,,,I17390,);
and I_3(I17744,I17727,I17679);
DFFARX1 I_4(I1470,,,I15576,);
or I_5(I17998,I17933,I17744);
nor I_6(I17679,I17662,I17515);
not I_7(I17933,I17916);
nand I_8(I17727,I17430,I15576);
DFFARX1 I_9(I1470,I17413,,,I17662,);
endmodule


