module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_11,blif_reset_net_1_r_11,G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_11,blif_reset_net_1_r_11;
output G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_431_0_l_11,n9_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_11,n9_11,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_11,n9_11,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_11,n9_11,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_11,n9_11,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_11,n9_11,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_11,n9_11,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_11,n9_11,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_11,n9_11,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_11,n9_11,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_11,n9_11,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_11,blif_clk_net_1_r_11,n9_11,G42_1_r_11,);
nor I_32(n_572_1_r_11,n29_11,n30_11);
nand I_33(n_573_1_r_11,n26_11,n28_11);
nor I_34(n_549_1_r_11,n27_11,n32_11);
nand I_35(n_569_1_r_11,n45_11,n28_11);
nor I_36(n_452_1_r_11,n43_11,n44_11);
nor I_37(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_38(N3_2_r_11,blif_clk_net_1_r_11,n9_11,G199_2_r_11,);
DFFARX1 I_39(n24_11,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_11,);
nor I_40(n_266_and_0_3_r_11,n20_11,n37_11);
or I_41(n_431_0_l_11,n33_11,ACVQN1_5_r_6);
not I_42(n9_11,blif_reset_net_1_r_11);
DFFARX1 I_43(n_431_0_l_11,blif_clk_net_1_r_11,n9_11,n43_11,);
not I_44(n26_11,n43_11);
DFFARX1 I_45(n_573_1_r_6,blif_clk_net_1_r_11,n9_11,n44_11,);
DFFARX1 I_46(n_572_1_r_6,blif_clk_net_1_r_11,n9_11,n45_11,);
not I_47(n27_11,n45_11);
nor I_48(n4_1_r_11,n44_11,n25_11);
nor I_49(N3_2_r_11,n45_11,n40_11);
nand I_50(n24_11,n39_11,G199_4_r_6);
nand I_51(n25_11,n38_11,P6_5_r_6);
DFFARX1 I_52(n25_11,blif_clk_net_1_r_11,n9_11,n20_internal_11,);
not I_53(n20_11,n20_internal_11);
not I_54(n28_11,n25_11);
not I_55(n29_11,G42_1_r_6);
nand I_56(n30_11,n26_11,n31_11);
not I_57(n31_11,n_549_1_r_6);
and I_58(n32_11,n26_11,n44_11);
and I_59(n33_11,n34_11,G42_1_r_6);
nor I_60(n34_11,n29_11,n_569_1_r_6);
not I_61(n35_11,n_452_1_r_6);
nand I_62(n36_11,n31_11,G42_1_r_6);
nor I_63(n37_11,n29_11,n_549_1_r_6);
nor I_64(n38_11,n31_11,n_452_1_r_6);
nor I_65(n39_11,n_452_1_r_6,G214_4_r_6);
nor I_66(n40_11,n41_11,n_452_1_r_6);
nor I_67(n41_11,n42_11,G214_4_r_6);
not I_68(n42_11,G199_4_r_6);
endmodule


