module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_8_r_8,n8_8,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_8,n46_8,n51_8);
not I_43(N1508_0_r_8,n46_8);
nor I_44(N1372_1_r_8,n37_8,n49_8);
and I_45(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_46(N1507_6_r_8,n47_8,n48_8);
nor I_47(N1508_6_r_8,n37_8,n38_8);
nor I_48(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_49(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_50(N6147_9_r_8,n29_8,n30_8);
nor I_51(N6134_9_r_8,n30_8,n31_8);
not I_52(I_BUFF_1_9_r_8,n35_8);
nor I_53(N1372_10_r_8,n46_8,n49_8);
nor I_54(N1508_10_r_8,n40_8,n41_8);
and I_55(N3_8_l_8,n36_8,n_429_or_0_5_r_11);
not I_56(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_57(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_58(n29_8,n53_8);
nor I_59(N3_8_r_8,n33_8,n34_8);
and I_60(n30_8,n32_8,n33_8);
nor I_61(n31_8,N1508_1_r_11,N6147_2_r_11);
nand I_62(n32_8,n42_8,N1372_1_r_11);
or I_63(n33_8,n46_8,N1372_1_r_11);
nor I_64(n34_8,n32_8,n35_8);
nand I_65(n35_8,n44_8,N1508_10_r_11);
nand I_66(n36_8,N1508_1_r_11,n_547_5_r_11);
not I_67(n37_8,n31_8);
nand I_68(n38_8,N1508_0_r_8,n39_8);
nand I_69(n39_8,n33_8,n50_8);
and I_70(n40_8,n32_8,n35_8);
not I_71(n41_8,N1372_10_r_8);
and I_72(n42_8,n43_8,G78_5_r_11);
nand I_73(n43_8,n44_8,n45_8);
nand I_74(n44_8,N6147_3_r_11,N1508_1_r_11);
not I_75(n45_8,N1508_10_r_11);
nand I_76(n46_8,n_576_5_r_11,N1507_6_r_11);
not I_77(n47_8,n39_8);
nor I_78(n48_8,n35_8,n49_8);
not I_79(n49_8,n51_8);
nand I_80(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_81(n51_8,n52_8,N6147_2_r_11);
or I_82(n52_8,N1508_6_r_11,N6147_3_r_11);
endmodule


