module test_I15372(I11105,I10633,I1477,I1470,I15372);
input I11105,I10633,I1477,I1470;
output I15372;
wire I12619,I12602,I12913,I10647,I12930,I14965,I10609;
not I_0(I12619,I1477);
not I_1(I12602,I12930);
DFFARX1 I_2(I10633,I1470,I12619,,,I12913,);
not I_3(I10647,I1477);
and I_4(I12930,I12913,I10609);
not I_5(I14965,I1477);
DFFARX1 I_6(I12602,I1470,I14965,,,I15372,);
DFFARX1 I_7(I11105,I1470,I10647,,,I10609,);
endmodule


