module test_I16886(I12930,I1477,I12590,I15194,I15406,I12584,I1470,I16886);
input I12930,I1477,I12590,I15194,I15406,I12584,I1470;
output I16886;
wire I14948,I14951,I14965,I12581,I15423,I15485,I12619,I15109,I15211,I15372,I15016,I14999,I15126,I15519,I15245,I15502;
DFFARX1 I_0(I15519,I1470,I14965,,,I14948,);
nand I_1(I14951,I15016,I15245);
not I_2(I14965,I1477);
DFFARX1 I_3(I12930,I1470,I12619,,,I12581,);
and I_4(I15423,I15372,I15406);
DFFARX1 I_5(I1470,I14965,,,I15485,);
not I_6(I12619,I1477);
not I_7(I15109,I12584);
DFFARX1 I_8(I15194,I1470,I14965,,,I15211,);
DFFARX1 I_9(I1470,I14965,,,I15372,);
nand I_10(I15016,I14999,I12581);
nor I_11(I14999,I12584,I12590);
not I_12(I15126,I15109);
or I_13(I15519,I15502,I15423);
nor I_14(I15245,I15211,I15126);
nor I_15(I16886,I14951,I14948);
not I_16(I15502,I15485);
endmodule


