module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_7,n8_7,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_7,n8_7,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_7,n8_7,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_7,n8_7,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_7,n8_7,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_7,n8_7,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_7,n8_7,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_7,n8_7,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_7,n8_7,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_34(n_572_1_r_7,n30_7,n31_7);
nand I_35(n_573_1_r_7,n28_7,G42_1_r_9);
nor I_36(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_37(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_38(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_39(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_40(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_41(P6_5_r_7,P6_5_r_internal_7);
or I_42(n_431_0_l_7,n36_7,n_572_1_r_9);
not I_43(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_44(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_45(n27_7,n43_7);
DFFARX1 I_46(n_549_1_r_9,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_47(n_572_1_r_9,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_48(n4_1_r_7,n30_7,n38_7);
nor I_49(N1_4_r_7,n27_7,n40_7);
nand I_50(n26_7,n39_7,G199_2_r_9);
not I_51(n5_7,n_42_2_r_9);
DFFARX1 I_52(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_53(n28_7,n26_7,n29_7);
not I_54(n29_7,n_569_1_r_9);
not I_55(n30_7,n_573_1_r_9);
nand I_56(n31_7,n27_7,n29_7);
nor I_57(n32_7,ACVQN1_5_l_7,n34_7);
nor I_58(n33_7,n29_7,n_42_2_r_9);
not I_59(n34_7,G42_1_r_9);
nor I_60(n35_7,n43_7,n44_7);
and I_61(n36_7,n37_7,G42_1_r_9);
nor I_62(n37_7,n30_7,G199_4_r_9);
nand I_63(n38_7,n29_7,n_42_2_r_9);
nor I_64(n39_7,n_42_2_r_9,G214_4_r_9);
nor I_65(n40_7,n44_7,n41_7);
nor I_66(n41_7,n34_7,n42_7);
nand I_67(n42_7,n5_7,n_569_1_r_9);
endmodule


