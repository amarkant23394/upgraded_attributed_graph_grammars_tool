module test_I4824(I1477,I1303,I1247,I1470,I2215,I4824);
input I1477,I1303,I1247,I1470,I2215;
output I4824;
wire I2540,I2143,I2181,I4544,I2170,I2557,I2232,I4807;
DFFARX1 I_0(I1247,I1470,I2181,,,I2540,);
DFFARX1 I_1(I2557,I1470,I2181,,,I2143,);
not I_2(I2181,I1477);
not I_3(I4544,I1477);
not I_4(I2170,I2232);
and I_5(I2557,I2540,I1303);
DFFARX1 I_6(I2215,I1470,I2181,,,I2232,);
DFFARX1 I_7(I2170,I1470,I4544,,,I4807,);
and I_8(I4824,I4807,I2143);
endmodule


