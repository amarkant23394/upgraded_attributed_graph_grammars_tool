module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_5_r_9,n10_9,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N6147_2_r_9,n62_9,n46_9);
not I_42(N1372_4_r_9,n59_9);
nor I_43(N1508_4_r_9,n58_9,n59_9);
nand I_44(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_45(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_46(n_576_5_r_9,n39_9,n40_9);
not I_47(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_48(n_547_5_r_9,n43_9,N1508_6_r_1);
and I_49(n_42_8_r_9,n44_9,N6147_9_r_1);
DFFARX1 I_50(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_51(N6147_9_r_9,n41_9,n45_9);
nor I_52(N6134_9_r_9,n45_9,n51_9);
nor I_53(I_BUFF_1_9_r_9,n41_9,N1508_6_r_1);
nor I_54(n4_7_l_9,N1507_6_r_1,N6147_9_r_1);
not I_55(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_56(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_57(N3_8_l_9,n57_9,N1508_0_r_1);
DFFARX1 I_58(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_59(n38_9,n63_9);
nor I_60(n_431_5_r_9,n_572_7_r_1,N1508_6_r_1);
nor I_61(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_62(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_63(n40_9,n41_9);
nand I_64(n41_9,N1508_0_r_1,n_569_7_r_1);
nor I_65(n42_9,G42_7_r_1,n_549_7_r_1);
nor I_66(n43_9,n63_9,n41_9);
nor I_67(n44_9,n_573_7_r_1,n_549_7_r_1);
and I_68(n45_9,n52_9,n_572_7_r_1);
nor I_69(n46_9,n47_9,n48_9);
nor I_70(n47_9,n49_9,n50_9);
not I_71(n48_9,n_429_or_0_5_r_9);
not I_72(n49_9,n42_9);
or I_73(n50_9,n63_9,n51_9);
nor I_74(n51_9,N1507_6_r_1,G42_7_r_1);
nor I_75(n52_9,n49_9,N1508_6_r_1);
nor I_76(n53_9,n54_9,n55_9);
nor I_77(n54_9,n56_9,N1508_6_r_1);
or I_78(n55_9,n44_9,G42_7_r_1);
not I_79(n56_9,n_572_7_r_1);
nand I_80(n57_9,N6134_9_r_1,G42_7_r_1);
nor I_81(n58_9,n62_9,n60_9);
nand I_82(n59_9,n51_9,n61_9);
nor I_83(n60_9,n38_9,n44_9);
nor I_84(n61_9,n_573_7_r_1,N6147_9_r_1);
endmodule


