module test_I4325(I2878,I1477,I4000,I1470,I1335,I2793,I4325);
input I2878,I1477,I4000,I1470,I1335,I2793;
output I4325;
wire I2730,I2810,I4017,I3124,I2727,I3076,I4308,I4034,I4051,I3983;
not I_0(I2730,I3076);
nand I_1(I2810,I2793,I1335);
and I_2(I4325,I4308,I4051);
and I_3(I4017,I4000,I2730);
nor I_4(I3124,I3076,I2878);
nand I_5(I2727,I2810,I3124);
DFFARX1 I_6(I1470,,,I3076,);
DFFARX1 I_7(I2727,I1470,I3983,,,I4308,);
DFFARX1 I_8(I4017,I1470,I3983,,,I4034,);
not I_9(I4051,I4034);
not I_10(I3983,I1477);
endmodule


