module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_13,blif_reset_net_1_r_13,G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_13,blif_reset_net_1_r_13;
output G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_569_1_r_13,n4_1_l_13,n7_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_13,n7_13,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_13,n7_13,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_13,n7_13,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_13,n7_13,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_13,n7_13,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_13,blif_clk_net_1_r_13,n7_13,G42_1_r_13,);
nor I_33(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_34(n_573_1_r_13,n18_13,n19_13);
nand I_35(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_36(n_569_1_r_13,n17_13,n18_13);
nor I_37(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_38(n_266_and_0_3_l_13,blif_clk_net_1_r_13,n7_13,ACVQN2_3_r_13,);
nor I_39(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_40(n_549_1_l_13,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_13,);
not I_41(P6_5_r_13,P6_5_r_internal_13);
nor I_42(n4_1_l_13,n_569_1_r_16,P6_5_r_16);
not I_43(n7_13,blif_reset_net_1_r_13);
DFFARX1 I_44(n4_1_l_13,blif_clk_net_1_r_13,n7_13,n17_internal_13,);
not I_45(n17_13,n17_internal_13);
DFFARX1 I_46(G42_1_r_16,blif_clk_net_1_r_13,n7_13,n28_13,);
DFFARX1 I_47(n_572_1_r_16,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_13,);
nor I_48(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_49(n_266_and_0_3_l_13,ACVQN1_3_l_13,ACVQN1_5_r_16);
nand I_50(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_51(n_573_1_l_13,blif_clk_net_1_r_13,n7_13,n14_internal_13,);
not I_52(n14_13,n14_internal_13);
and I_53(n_549_1_l_13,n21_13,n26_13);
nand I_54(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_55(n_569_1_l_13,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_13,);
nand I_56(n18_13,n23_13,n24_13);
or I_57(n19_13,G199_4_r_16,G214_4_r_16);
not I_58(n20_13,G42_1_r_16);
not I_59(n21_13,n_452_1_r_16);
nand I_60(n22_13,n17_13,n28_13);
not I_61(n23_13,n_569_1_r_16);
not I_62(n24_13,n_573_1_r_16);
nor I_63(n25_13,G199_4_r_16,G214_4_r_16);
nand I_64(n26_13,n27_13,n_549_1_r_16);
not I_65(n27_13,G199_4_r_16);
endmodule


