module test_I6941(I1477,I3521,I3846,I1470,I5122,I3453,I6941);
input I1477,I3521,I3846,I1470,I5122,I3453;
output I6941;
wire I5416,I5105,I5187,I3353,I5070,I3380,I3637,I5249,I5094,I3356,I5204,I5481;
nand I_0(I5416,I5122,I3356);
not I_1(I5105,I1477);
nor I_2(I5187,I5122,I3380);
nor I_3(I6941,I5070,I5094);
and I_4(I3353,I3453,I3637);
and I_5(I5070,I5249,I5481);
nand I_6(I3380,I3521,I3846);
DFFARX1 I_7(I1470,,,I3637,);
not I_8(I5249,I3380);
not I_9(I5094,I5204);
DFFARX1 I_10(I1470,,,I3356,);
nand I_11(I5204,I5187,I3353);
DFFARX1 I_12(I5416,I1470,I5105,,,I5481,);
endmodule


