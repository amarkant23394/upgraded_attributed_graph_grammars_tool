module test_I16810(I14930,I1477,I1470,I17013,I16852,I16810);
input I14930,I1477,I1470,I17013,I16852;
output I16810;
wire I14927,I17222,I17047,I17239,I17205,I16869,I16818,I17030;
DFFARX1 I_0(I1470,,,I14927,);
nand I_1(I17222,I17205,I16869);
DFFARX1 I_2(I17030,I1470,I16818,,,I17047,);
and I_3(I17239,I17047,I17222);
DFFARX1 I_4(I14927,I1470,I16818,,,I17205,);
DFFARX1 I_5(I16852,I1470,I16818,,,I16869,);
DFFARX1 I_6(I17239,I1470,I16818,,,I16810,);
not I_7(I16818,I1477);
and I_8(I17030,I17013,I14930);
endmodule


