module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_8_r_6,n9_6,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_8_r_6,n9_6,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_6,n30_6,n33_6);
nor I_36(N1508_0_r_6,n33_6,n44_6);
not I_37(N1372_1_r_6,n41_6);
nor I_38(N1508_1_r_6,n40_6,n41_6);
nor I_39(N1507_6_r_6,n39_6,n45_6);
nor I_40(N1508_6_r_6,n37_6,n38_6);
nor I_41(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_42(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_43(N6147_9_r_6,n32_6,n33_6);
nor I_44(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_45(I_BUFF_1_9_r_6,n37_6);
not I_46(N1372_10_r_6,n43_6);
nor I_47(N1508_10_r_6,n42_6,n43_6);
nor I_48(N3_8_r_6,n36_6,n_429_or_0_5_r_0);
not I_49(n9_6,blif_reset_net_8_r_6);
nor I_50(n30_6,n53_6,G78_5_r_0);
not I_51(n31_6,n36_6);
nor I_52(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_53(n33_6,n_429_or_0_5_r_0);
not I_54(n34_6,n35_6);
nand I_55(n35_6,n49_6,n_569_7_r_0);
nand I_56(n36_6,n51_6,G42_7_r_0);
nand I_57(n37_6,n54_6,n_549_7_r_0);
or I_58(n38_6,n35_6,n39_6);
nor I_59(n39_6,n40_6,n45_6);
and I_60(n40_6,n46_6,n47_6);
nand I_61(n41_6,n30_6,n31_6);
nor I_62(n42_6,n34_6,n40_6);
nand I_63(n43_6,n30_6,n_429_or_0_5_r_0);
nor I_64(n44_6,n31_6,n40_6);
nor I_65(n45_6,n35_6,n36_6);
nor I_66(n46_6,N1371_0_r_0,N1508_0_r_0);
or I_67(n47_6,n48_6,G78_5_r_0);
nor I_68(n48_6,n_576_5_r_0,n_572_7_r_0);
and I_69(n49_6,n50_6,n_573_7_r_0);
nand I_70(n50_6,n51_6,n52_6);
nand I_71(n51_6,N1508_0_r_0,n_576_5_r_0);
not I_72(n52_6,G42_7_r_0);
nor I_73(n53_6,n_547_5_r_0,n_429_or_0_5_r_0);
or I_74(n54_6,n_547_5_r_0,n_429_or_0_5_r_0);
endmodule


