module test_I5743(I2167,I1477,I4524,I5994,I5768,I2173,I1470,I5743);
input I2167,I1477,I4524,I5994,I5768,I2173,I1470;
output I5743;
wire I4629,I6110,I6028,I4544,I5785,I5802,I2143,I6011,I5751,I4521,I6079,I4533,I5013,I4807,I6127,I4824,I4509;
nor I_0(I4629,I2167,I2173);
DFFARX1 I_1(I4509,I1470,I5751,,,I6110,);
DFFARX1 I_2(I6011,I1470,I5751,,,I6028,);
nand I_3(I5743,I6127,I6079);
not I_4(I4544,I1477);
and I_5(I5785,I5768,I4524);
DFFARX1 I_6(I5785,I1470,I5751,,,I5802,);
DFFARX1 I_7(I1470,,,I2143,);
and I_8(I6011,I5994,I4521);
not I_9(I5751,I1477);
DFFARX1 I_10(I1470,I4544,,,I4521,);
nor I_11(I6079,I6028,I5802);
or I_12(I4533,I4824,I4629);
or I_13(I5013,I4824);
DFFARX1 I_14(I1470,I4544,,,I4807,);
and I_15(I6127,I6110,I4533);
and I_16(I4824,I4807,I2143);
DFFARX1 I_17(I5013,I1470,I4544,,,I4509,);
endmodule


