module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_5_r_13,n9_13,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_5_r_13,n9_13,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_13,n59_13,n61_13);
nor I_36(N1508_0_r_13,n59_13,n60_13);
not I_37(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_38(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_39(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_40(n_102_5_r_13,N1371_0_r_0,N1508_0_r_0);
nand I_41(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_42(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_43(n_572_7_r_13,n40_13,n41_13);
nand I_44(n_573_7_r_13,n37_13,n38_13);
nor I_45(n_549_7_r_13,n46_13,n47_13);
nand I_46(n_569_7_r_13,n37_13,n43_13);
nand I_47(n_452_7_r_13,n52_13,n53_13);
nor I_48(n4_7_l_13,n_429_or_0_5_r_0,n_549_7_r_0);
not I_49(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_50(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_51(n33_13,n62_13);
nand I_52(n_431_5_r_13,n54_13,n55_13);
not I_53(n1_13,n52_13);
nor I_54(n34_13,n35_13,n36_13);
nor I_55(n35_13,n42_13,n_576_5_r_0);
nand I_56(n36_13,n50_13,n58_13);
nand I_57(n37_13,n44_13,n45_13);
or I_58(n38_13,n39_13,N1508_0_r_0);
nand I_59(n39_13,n_569_7_r_0,G78_5_r_0);
not I_60(n40_13,n36_13);
nor I_61(n41_13,n35_13,N1371_0_r_0);
not I_62(n42_13,n_429_or_0_5_r_0);
or I_63(n43_13,n_429_or_0_5_r_0,n_547_5_r_0);
not I_64(n44_13,n_576_5_r_0);
not I_65(n45_13,G78_5_r_0);
nor I_66(n46_13,n39_13,n40_13);
nor I_67(n47_13,n_429_or_0_5_r_0,n_547_5_r_0);
nor I_68(n48_13,n50_13,n51_13);
nor I_69(n49_13,G78_5_r_0,n_576_5_r_0);
not I_70(n50_13,n59_13);
not I_71(n51_13,n_102_5_r_13);
nand I_72(n52_13,n33_13,n39_13);
nand I_73(n53_13,n33_13,N1508_0_r_0);
nor I_74(n54_13,n_547_5_r_0,N1508_0_r_0);
nand I_75(n55_13,n62_13,n56_13);
nor I_76(n56_13,n39_13,n57_13);
not I_77(n57_13,n_429_or_0_5_r_0);
or I_78(n58_13,N1371_0_r_0,n_572_7_r_0);
nand I_79(n59_13,G42_7_r_0,n_573_7_r_0);
nor I_80(n60_13,n51_13,n_547_5_r_0);
nor I_81(n61_13,n39_13,N1508_0_r_0);
endmodule


