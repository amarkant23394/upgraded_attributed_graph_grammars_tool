module test_I15696(I12304,I1470,I13775,I12058,I11973,I12380,I11944,I15696);
input I12304,I1470,I13775,I12058,I11973,I12380,I11944;
output I15696;
wire I13826,I13761,I13743,I13860,I15628,I13891,I13843,I13758,I11959,I15679,I11965;
DFFARX1 I_0(I1470,I13775,,,I13826,);
nand I_1(I13761,I13891,I13860);
DFFARX1 I_2(I13891,I1470,I13775,,,I13743,);
nand I_3(I15696,I15679,I13758);
nor I_4(I13860,I13843,I13826);
not I_5(I15628,I13743);
DFFARX1 I_6(I11944,I1470,I13775,,,I13891,);
nor I_7(I13843,I11959,I11965);
not I_8(I13758,I13843);
nand I_9(I11959,I12058,I12380);
nor I_10(I15679,I15628,I13761);
DFFARX1 I_11(I12304,I1470,I11973,,,I11965,);
endmodule


