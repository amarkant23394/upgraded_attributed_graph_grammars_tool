module test_I5751(I1477,I5751);
input I1477;
output I5751;
wire ;
not I_0(I5751,I1477);
endmodule


