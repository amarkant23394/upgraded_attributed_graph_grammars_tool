module test_I1656(I1255,I1247,I1279,I1294,I1271,I1207,I1301,I1656);
input I1255,I1247,I1279,I1294,I1271,I1207,I1301;
output I1656;
wire I1622,I1492,I1342,I1475,I1509,I1639;
DFFARX1 I_0(I1255,I1294,I1342,,,I1622,);
nand I_1(I1656,I1639,I1509);
and I_2(I1492,I1475,I1279);
not I_3(I1342,I1301);
nand I_4(I1475,I1247,I1271);
DFFARX1 I_5(I1492,I1294,I1342,,,I1509,);
and I_6(I1639,I1622,I1207);
endmodule


