module test_I10052_rst(I1477_rst,I10052_rst);
,I10052_rst);
input I1477_rst;
output I10052_rst;
wire ;
not I_0(I10052_rst,I1477_rst);
endmodule


