module Benchmark_testing100(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301,I3217,I3214,I3208,I3238,I3211,I3235,I3232,I3229,I3223,I3226,I3220);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301;
output I3217,I3214,I3208,I3238,I3211,I3235,I3232,I3229,I3223,I3226,I3220;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301,I1342,I1359,I1376,I1393,I1410,I1427,I1444,I1313,I1475,I1492,I1509,I1526,I1543,I1560,I1577,I1310,I1304,I1622,I1639,I1656,I1331,I1687,I1704,I1322,I1316,I1749,I1319,I1780,I1797,I1334,I1828,I1328,I1325,I1873,I1307,I1937,I1954,I1971,I1988,I2005,I2022,I2039,I1908,I2070,I2087,I2104,I2121,I2138,I2155,I2172,I1905,I2203,I1899,I2234,I2251,I2268,I1929,I1902,I2313,I1926,I2344,I1923,I1920,I2389,I2406,I2423,I2440,I2457,I1914,I2488,I2505,I1917,I1911,I2583,I2600,I2617,I2634,I2651,I2668,I2685,I2702,I2572,I2733,I2557,I2764,I2781,I2798,I2815,I2832,I2849,I2866,I2554,I2897,I2914,I2551,I2945,I2962,I2569,I2993,I2566,I3024,I3041,I2545,I2548,I3086,I3103,I3120,I3137,I2575,I3168,I2560,I2563,I3246,I3263,I3280,I3297,I3314,I3331,I3348,I3379,I3396,I3413,I3430,I3447,I3464,I3481,I3512,I3543,I3560,I3577,I3622,I3653,I3698,I3715,I3732,I3749,I3766,I3797,I3814;
not I_0 (I1342,I1301);
nand I_1 (I1359,I1287,I1239);
and I_2 (I1376,I1359,I1231);
DFFARX1 I_3  ( .D(I1376), .CLK(I1294), .RSTB(I1342), .Q(I1393) );
nor I_4 (I1410,I1223,I1239);
DFFARX1 I_5  ( .D(I1263), .CLK(I1294), .RSTB(I1342), .Q(I1427) );
nand I_6 (I1444,I1427,I1410);
DFFARX1 I_7  ( .D(I1427), .CLK(I1294), .RSTB(I1342), .Q(I1313) );
nand I_8 (I1475,I1247,I1271);
and I_9 (I1492,I1475,I1279);
DFFARX1 I_10  ( .D(I1492), .CLK(I1294), .RSTB(I1342), .Q(I1509) );
not I_11 (I1526,I1509);
nor I_12 (I1543,I1393,I1526);
and I_13 (I1560,I1410,I1543);
and I_14 (I1577,I1509,I1444);
DFFARX1 I_15  ( .D(I1577), .CLK(I1294), .RSTB(I1342), .Q(I1310) );
DFFARX1 I_16  ( .D(I1509), .CLK(I1294), .RSTB(I1342), .Q(I1304) );
DFFARX1 I_17  ( .D(I1255), .CLK(I1294), .RSTB(I1342), .Q(I1622) );
and I_18 (I1639,I1622,I1207);
nand I_19 (I1656,I1639,I1509);
nor I_20 (I1331,I1639,I1410);
not I_21 (I1687,I1639);
nor I_22 (I1704,I1393,I1687);
nand I_23 (I1322,I1427,I1704);
nand I_24 (I1316,I1509,I1687);
or I_25 (I1749,I1639,I1560);
DFFARX1 I_26  ( .D(I1749), .CLK(I1294), .RSTB(I1342), .Q(I1319) );
DFFARX1 I_27  ( .D(I1215), .CLK(I1294), .RSTB(I1342), .Q(I1780) );
and I_28 (I1797,I1780,I1656);
DFFARX1 I_29  ( .D(I1797), .CLK(I1294), .RSTB(I1342), .Q(I1334) );
nor I_30 (I1828,I1780,I1393);
nand I_31 (I1328,I1639,I1828);
not I_32 (I1325,I1780);
DFFARX1 I_33  ( .D(I1780), .CLK(I1294), .RSTB(I1342), .Q(I1873) );
and I_34 (I1307,I1780,I1873);
not I_35 (I1937,I1301);
not I_36 (I1954,I1322);
nor I_37 (I1971,I1310,I1319);
nand I_38 (I1988,I1971,I1334);
nor I_39 (I2005,I1954,I1310);
nand I_40 (I2022,I2005,I1316);
DFFARX1 I_41  ( .D(I2022), .CLK(I1294), .RSTB(I1937), .Q(I2039) );
not I_42 (I1908,I2039);
not I_43 (I2070,I1310);
not I_44 (I2087,I2070);
not I_45 (I2104,I1304);
nor I_46 (I2121,I2104,I1325);
and I_47 (I2138,I2121,I1307);
or I_48 (I2155,I2138,I1313);
DFFARX1 I_49  ( .D(I2155), .CLK(I1294), .RSTB(I1937), .Q(I2172) );
DFFARX1 I_50  ( .D(I2172), .CLK(I1294), .RSTB(I1937), .Q(I1905) );
DFFARX1 I_51  ( .D(I2172), .CLK(I1294), .RSTB(I1937), .Q(I2203) );
DFFARX1 I_52  ( .D(I2172), .CLK(I1294), .RSTB(I1937), .Q(I1899) );
nand I_53 (I2234,I1954,I1304);
nand I_54 (I2251,I2234,I1988);
and I_55 (I2268,I2070,I2251);
DFFARX1 I_56  ( .D(I2268), .CLK(I1294), .RSTB(I1937), .Q(I1929) );
and I_57 (I1902,I2234,I2203);
DFFARX1 I_58  ( .D(I1331), .CLK(I1294), .RSTB(I1937), .Q(I2313) );
nor I_59 (I1926,I2313,I2234);
nor I_60 (I2344,I2313,I1988);
nand I_61 (I1923,I2022,I2344);
not I_62 (I1920,I2313);
DFFARX1 I_63  ( .D(I1328), .CLK(I1294), .RSTB(I1937), .Q(I2389) );
not I_64 (I2406,I2389);
nor I_65 (I2423,I2406,I2087);
and I_66 (I2440,I2313,I2423);
or I_67 (I2457,I2234,I2440);
DFFARX1 I_68  ( .D(I2457), .CLK(I1294), .RSTB(I1937), .Q(I1914) );
not I_69 (I2488,I2406);
nor I_70 (I2505,I2313,I2488);
nand I_71 (I1917,I2406,I2505);
nand I_72 (I1911,I2070,I2488);
not I_73 (I2583,I1301);
not I_74 (I2600,I1911);
nor I_75 (I2617,I1908,I1926);
nand I_76 (I2634,I2617,I1929);
nor I_77 (I2651,I2600,I1908);
nand I_78 (I2668,I2651,I1914);
not I_79 (I2685,I2668);
not I_80 (I2702,I1908);
nor I_81 (I2572,I2668,I2702);
not I_82 (I2733,I2702);
nand I_83 (I2557,I2668,I2733);
not I_84 (I2764,I1923);
nor I_85 (I2781,I2764,I1905);
and I_86 (I2798,I2781,I1899);
or I_87 (I2815,I2798,I1917);
DFFARX1 I_88  ( .D(I2815), .CLK(I1294), .RSTB(I2583), .Q(I2832) );
nor I_89 (I2849,I2832,I2685);
DFFARX1 I_90  ( .D(I2832), .CLK(I1294), .RSTB(I2583), .Q(I2866) );
not I_91 (I2554,I2866);
nand I_92 (I2897,I2600,I1923);
and I_93 (I2914,I2897,I2849);
DFFARX1 I_94  ( .D(I2897), .CLK(I1294), .RSTB(I2583), .Q(I2551) );
DFFARX1 I_95  ( .D(I1902), .CLK(I1294), .RSTB(I2583), .Q(I2945) );
nor I_96 (I2962,I2945,I2668);
nand I_97 (I2569,I2832,I2962);
nor I_98 (I2993,I2945,I2733);
not I_99 (I2566,I2945);
nand I_100 (I3024,I2945,I2634);
and I_101 (I3041,I2702,I3024);
DFFARX1 I_102  ( .D(I3041), .CLK(I1294), .RSTB(I2583), .Q(I2545) );
DFFARX1 I_103  ( .D(I2945), .CLK(I1294), .RSTB(I2583), .Q(I2548) );
DFFARX1 I_104  ( .D(I1920), .CLK(I1294), .RSTB(I2583), .Q(I3086) );
not I_105 (I3103,I3086);
nand I_106 (I3120,I3103,I2668);
and I_107 (I3137,I2897,I3120);
DFFARX1 I_108  ( .D(I3137), .CLK(I1294), .RSTB(I2583), .Q(I2575) );
or I_109 (I3168,I3103,I2914);
DFFARX1 I_110  ( .D(I3168), .CLK(I1294), .RSTB(I2583), .Q(I2560) );
nand I_111 (I2563,I3103,I2993);
not I_112 (I3246,I1301);
not I_113 (I3263,I2569);
nor I_114 (I3280,I2548,I2560);
nand I_115 (I3297,I3280,I2563);
nor I_116 (I3314,I3263,I2548);
nand I_117 (I3331,I3314,I2545);
DFFARX1 I_118  ( .D(I3331), .CLK(I1294), .RSTB(I3246), .Q(I3348) );
not I_119 (I3217,I3348);
not I_120 (I3379,I2548);
not I_121 (I3396,I3379);
not I_122 (I3413,I2566);
nor I_123 (I3430,I3413,I2557);
and I_124 (I3447,I3430,I2551);
or I_125 (I3464,I3447,I2575);
DFFARX1 I_126  ( .D(I3464), .CLK(I1294), .RSTB(I3246), .Q(I3481) );
DFFARX1 I_127  ( .D(I3481), .CLK(I1294), .RSTB(I3246), .Q(I3214) );
DFFARX1 I_128  ( .D(I3481), .CLK(I1294), .RSTB(I3246), .Q(I3512) );
DFFARX1 I_129  ( .D(I3481), .CLK(I1294), .RSTB(I3246), .Q(I3208) );
nand I_130 (I3543,I3263,I2566);
nand I_131 (I3560,I3543,I3297);
and I_132 (I3577,I3379,I3560);
DFFARX1 I_133  ( .D(I3577), .CLK(I1294), .RSTB(I3246), .Q(I3238) );
and I_134 (I3211,I3543,I3512);
DFFARX1 I_135  ( .D(I2572), .CLK(I1294), .RSTB(I3246), .Q(I3622) );
nor I_136 (I3235,I3622,I3543);
nor I_137 (I3653,I3622,I3297);
nand I_138 (I3232,I3331,I3653);
not I_139 (I3229,I3622);
DFFARX1 I_140  ( .D(I2554), .CLK(I1294), .RSTB(I3246), .Q(I3698) );
not I_141 (I3715,I3698);
nor I_142 (I3732,I3715,I3396);
and I_143 (I3749,I3622,I3732);
or I_144 (I3766,I3543,I3749);
DFFARX1 I_145  ( .D(I3766), .CLK(I1294), .RSTB(I3246), .Q(I3223) );
not I_146 (I3797,I3715);
nor I_147 (I3814,I3622,I3797);
nand I_148 (I3226,I3715,I3814);
nand I_149 (I3220,I3379,I3797);
endmodule


