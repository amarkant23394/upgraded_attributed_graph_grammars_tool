module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_7_r_2,n10_2,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N1371_0_r_2,n32_2,n35_2);
nor I_42(N1508_0_r_2,n32_2,n55_2);
not I_43(N1372_1_r_2,n54_2);
nor I_44(N1508_1_r_2,n59_2,n54_2);
nor I_45(N6147_2_r_2,n42_2,n43_2);
nor I_46(N1507_6_r_2,n40_2,n53_2);
nor I_47(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_48(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_49(n_572_7_r_2,n36_2,n37_2);
or I_50(n_573_7_r_2,n34_2,n35_2);
nor I_51(n_549_7_r_2,n40_2,n41_2);
nand I_52(n_569_7_r_2,n38_2,n39_2);
nor I_53(n_452_7_r_2,n59_2,n35_2);
nor I_54(n4_7_l_2,N1507_6_r_1,G42_7_r_1);
not I_55(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_56(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_57(n33_2,n59_2);
and I_58(N3_8_l_2,n49_2,n_572_7_r_1);
DFFARX1 I_59(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_60(n32_2,n32_internal_2);
nor I_61(n4_7_r_2,n59_2,n36_2);
not I_62(n34_2,n39_2);
nor I_63(n35_2,N1508_0_r_1,n_569_7_r_1);
nor I_64(n36_2,N1507_6_r_1,G42_7_r_1);
or I_65(n37_2,N1508_6_r_1,n_572_7_r_1);
not I_66(n38_2,n40_2);
nand I_67(n39_2,n45_2,n57_2);
nor I_68(n40_2,n47_2,n_573_7_r_1);
nor I_69(n41_2,n32_2,n36_2);
not I_70(n42_2,n53_2);
nand I_71(n43_2,n44_2,n45_2);
nand I_72(n44_2,n38_2,n46_2);
not I_73(n45_2,N1508_6_r_1);
nand I_74(n46_2,n47_2,n48_2);
nand I_75(n47_2,G42_7_r_1,N6147_9_r_1);
or I_76(n48_2,n_549_7_r_1,N6134_9_r_1);
nand I_77(n49_2,N1508_0_r_1,N1508_6_r_1);
nand I_78(n50_2,n51_2,n52_2);
not I_79(n51_2,n47_2);
nand I_80(n52_2,n38_2,n53_2);
nor I_81(n53_2,N1507_6_r_1,n_572_7_r_1);
nand I_82(n54_2,n42_2,n56_2);
nor I_83(n55_2,n34_2,n56_2);
nor I_84(n56_2,n_549_7_r_1,N6134_9_r_1);
nand I_85(n57_2,n58_2,N1508_0_r_1);
not I_86(n58_2,n_549_7_r_1);
endmodule


