module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_8_r_8,n8_8,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_8,n46_8,n51_8);
not I_37(N1508_0_r_8,n46_8);
nor I_38(N1372_1_r_8,n37_8,n49_8);
and I_39(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_40(N1507_6_r_8,n47_8,n48_8);
nor I_41(N1508_6_r_8,n37_8,n38_8);
nor I_42(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_43(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_44(N6147_9_r_8,n29_8,n30_8);
nor I_45(N6134_9_r_8,n30_8,n31_8);
not I_46(I_BUFF_1_9_r_8,n35_8);
nor I_47(N1372_10_r_8,n46_8,n49_8);
nor I_48(N1508_10_r_8,n40_8,n41_8);
and I_49(N3_8_l_8,n36_8,N1371_0_r_5);
not I_50(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_51(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_52(n29_8,n53_8);
nor I_53(N3_8_r_8,n33_8,n34_8);
and I_54(n30_8,n32_8,n33_8);
nor I_55(n31_8,N1508_0_r_5,N6147_2_r_5);
nand I_56(n32_8,n42_8,n_573_7_r_5);
or I_57(n33_8,n46_8,N1508_1_r_5);
nor I_58(n34_8,n32_8,n35_8);
nand I_59(n35_8,n44_8,N1372_1_r_5);
nand I_60(n36_8,N6147_2_r_5,G42_7_r_5);
not I_61(n37_8,n31_8);
nand I_62(n38_8,N1508_0_r_8,n39_8);
nand I_63(n39_8,n33_8,n50_8);
and I_64(n40_8,n32_8,n35_8);
not I_65(n41_8,N1372_10_r_8);
and I_66(n42_8,n43_8,n_452_7_r_5);
nand I_67(n43_8,n44_8,n45_8);
nand I_68(n44_8,n_572_7_r_5,N1371_0_r_5);
not I_69(n45_8,N1372_1_r_5);
nand I_70(n46_8,N1507_6_r_5,N1508_6_r_5);
not I_71(n47_8,n39_8);
nor I_72(n48_8,n35_8,n49_8);
not I_73(n49_8,n51_8);
nand I_74(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_75(n51_8,n52_8,n_569_7_r_5);
or I_76(n52_8,N1372_1_r_5,N1508_0_r_5);
endmodule


