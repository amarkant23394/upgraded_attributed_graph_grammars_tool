module test_I13601(I1477,I1470,I11327,I9083,I9413,I13601);
input I1477,I1470,I11327,I9083,I9413;
output I13601;
wire I11378,I11429,I9066,I13197,I11299,I11395,I8848,I8851;
nor I_0(I11378,I11327,I8848);
DFFARX1 I_1(I11299,I1470,I13197,,,I13601,);
not I_2(I11429,I8848);
DFFARX1 I_3(I1470,,,I9066,);
not I_4(I13197,I1477);
nor I_5(I11299,I11395,I11429);
nand I_6(I11395,I11378,I8851);
nor I_7(I8848,I9083,I9413);
or I_8(I8851,I9083,I9066);
endmodule


