module test_I10270(I1477,I10202,I7881,I1470,I10270);
input I1477,I10202,I7881,I1470;
output I10270;
wire I10253,I10120,I6297,I7538,I10219,I10052,I7898,I7714,I7946,I10236,I7535,I10069,I10086,I7570,I7544,I7915,I10103;
nor I_0(I10253,I10103,I10236);
nor I_1(I10120,I7538,I7535);
DFFARX1 I_2(I1470,,,I6297,);
DFFARX1 I_3(I7915,I1470,I7570,,,I7538,);
DFFARX1 I_4(I10202,I1470,I10052,,,I10219,);
not I_5(I10052,I1477);
nand I_6(I7898,I7881);
not I_7(I7714,I6297);
DFFARX1 I_8(I7881,I1470,I7570,,,I7946,);
not I_9(I10236,I10219);
and I_10(I7535,I7714,I7946);
nand I_11(I10069,I7535);
and I_12(I10270,I10120,I10253);
and I_13(I10086,I10069,I7544);
not I_14(I7570,I1477);
DFFARX1 I_15(I1470,I7570,,,I7544,);
and I_16(I7915,I7881,I7898);
DFFARX1 I_17(I10086,I1470,I10052,,,I10103,);
endmodule


