module test_I6606(I1477,I1470,I4263,I4212,I6606);
input I1477,I1470,I4263,I4212;
output I6606;
wire I3960,I3951,I3945,I6589,I6329,I4113,I6572,I4308,I4229,I4356,I3983;
DFFARX1 I_0(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_1(I4356,I1470,I3983,,,I3960,);
nand I_2(I3951,I4263,I4229);
nand I_3(I3945,I4308,I4212);
and I_4(I6589,I6572,I3960);
not I_5(I6329,I1477);
DFFARX1 I_6(I1470,I3983,,,I4113,);
nand I_7(I6572,I3951,I3945);
DFFARX1 I_8(I1470,I3983,,,I4308,);
nor I_9(I4229,I4113,I4212);
nor I_10(I4356,I4308,I4113);
not I_11(I3983,I1477);
endmodule


