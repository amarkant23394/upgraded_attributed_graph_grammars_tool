module test_I9258(I5097,I9083,I9049,I7139,I5070,I1470_clk,I1477_rst,I9258);
input I5097,I9083,I9049,I7139,I5070,I1470_clk,I1477_rst;
output I9258;
wire I9131,I7286,I6907_rst,I8964,I6975,I9179,I9066,I6992,I9148,I7026,I7156,I6896,I6893,I9114,I8862_rst;
nor I_0(I9131,I9066,I9114);
nor I_1(I7286,I6992);
not I_2(I6907_rst,I1477_rst);
not I_3(I8964,I6893);
or I_4(I9258,I9179,I9148);
nor I_5(I6975,I5070);
DFFARX1 I_6 (I6896,I1470_clk,I8862_rst,I9179);
DFFARX1 I_7 (I9049,I1470_clk,I8862_rst,I9066);
nand I_8(I6992,I6975,I5097);
and I_9(I9148,I8964,I9131);
not I_10(I7026,I5070);
DFFARX1 I_11 (I7139,I1470_clk,I6907_rst,I7156);
nor I_12(I6896,I6992,I7026);
nand I_13(I6893,I7156,I7286);
not I_14(I9114,I9083);
not I_15(I8862_rst,I1477_rst);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule