module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2,n4_7_l_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_2,n32_2,n35_2);
nor I_1(N1508_0_r_2,n32_2,n55_2);
not I_2(N1372_1_r_2,n54_2);
nor I_3(N1508_1_r_2,n59_2,n54_2);
nor I_4(N6147_2_r_2,n42_2,n43_2);
nor I_5(N1507_6_r_2,n40_2,n53_2);
nor I_6(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_7(n4_7_r_2,blif_clk_net_5_r_13,n9_13,G42_7_r_2,);
nor I_8(n_572_7_r_2,n36_2,n37_2);
or I_9(n_573_7_r_2,n34_2,n35_2);
nor I_10(n_549_7_r_2,n40_2,n41_2);
nand I_11(n_569_7_r_2,n38_2,n39_2);
nor I_12(n_452_7_r_2,n59_2,n35_2);
nor I_13(n4_7_l_2,G18_7_l_2,IN_1_7_l_2);
DFFARX1 I_14(n4_7_l_2,blif_clk_net_5_r_13,n9_13,n59_2,);
not I_15(n33_2,n59_2);
and I_16(N3_8_l_2,IN_6_8_l_2,n49_2);
DFFARX1 I_17(N3_8_l_2,blif_clk_net_5_r_13,n9_13,n32_internal_2,);
not I_18(n32_2,n32_internal_2);
nor I_19(n4_7_r_2,n59_2,n36_2);
not I_20(n34_2,n39_2);
nor I_21(n35_2,IN_1_8_l_2,IN_3_8_l_2);
nor I_22(n36_2,G18_7_l_2,IN_5_7_l_2);
or I_23(n37_2,IN_9_7_l_2,IN_10_7_l_2);
not I_24(n38_2,n40_2);
nand I_25(n39_2,n45_2,n57_2);
nor I_26(n40_2,IN_3_1_l_2,n47_2);
nor I_27(n41_2,n32_2,n36_2);
not I_28(n42_2,n53_2);
nand I_29(n43_2,n44_2,n45_2);
nand I_30(n44_2,n38_2,n46_2);
not I_31(n45_2,IN_10_7_l_2);
nand I_32(n46_2,n47_2,n48_2);
nand I_33(n47_2,IN_1_1_l_2,IN_2_1_l_2);
or I_34(n48_2,G15_7_l_2,IN_7_7_l_2);
nand I_35(n49_2,IN_2_8_l_2,IN_3_8_l_2);
nand I_36(n50_2,n51_2,n52_2);
not I_37(n51_2,n47_2);
nand I_38(n52_2,n38_2,n53_2);
nor I_39(n53_2,IN_5_7_l_2,IN_9_7_l_2);
nand I_40(n54_2,n42_2,n56_2);
nor I_41(n55_2,n34_2,n56_2);
nor I_42(n56_2,G15_7_l_2,IN_7_7_l_2);
nand I_43(n57_2,IN_4_7_l_2,n58_2);
not I_44(n58_2,G15_7_l_2);
nor I_45(N1371_0_r_13,n59_13,n61_13);
nor I_46(N1508_0_r_13,n59_13,n60_13);
not I_47(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_48(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_49(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_50(n_102_5_r_13,N1508_1_r_2,n_452_7_r_2);
nand I_51(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_52(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_53(n_572_7_r_13,n40_13,n41_13);
nand I_54(n_573_7_r_13,n37_13,n38_13);
nor I_55(n_549_7_r_13,n46_13,n47_13);
nand I_56(n_569_7_r_13,n37_13,n43_13);
nand I_57(n_452_7_r_13,n52_13,n53_13);
nor I_58(n4_7_l_13,n_549_7_r_2,N1508_0_r_2);
not I_59(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_60(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_61(n33_13,n62_13);
nand I_62(n_431_5_r_13,n54_13,n55_13);
not I_63(n1_13,n52_13);
nor I_64(n34_13,n35_13,n36_13);
nor I_65(n35_13,n42_13,N1372_1_r_2);
nand I_66(n36_13,n50_13,n58_13);
nand I_67(n37_13,n44_13,n45_13);
or I_68(n38_13,n39_13,n_572_7_r_2);
nand I_69(n39_13,N1371_0_r_2,N6147_2_r_2);
not I_70(n40_13,n36_13);
nor I_71(n41_13,n35_13,N1508_1_r_2);
not I_72(n42_13,N1507_6_r_2);
or I_73(n43_13,N1508_0_r_2,n_549_7_r_2);
not I_74(n44_13,N1372_1_r_2);
not I_75(n45_13,n_573_7_r_2);
nor I_76(n46_13,n39_13,n40_13);
nor I_77(n47_13,N1508_0_r_2,n_549_7_r_2);
nor I_78(n48_13,n50_13,n51_13);
nor I_79(n49_13,N1372_1_r_2,n_573_7_r_2);
not I_80(n50_13,n59_13);
not I_81(n51_13,n_102_5_r_13);
nand I_82(n52_13,n33_13,n39_13);
nand I_83(n53_13,n33_13,n_572_7_r_2);
nor I_84(n54_13,N1508_0_r_2,n_452_7_r_2);
nand I_85(n55_13,n62_13,n56_13);
nor I_86(n56_13,n39_13,n57_13);
not I_87(n57_13,n_549_7_r_2);
or I_88(n58_13,n_569_7_r_2,N1371_0_r_2);
nand I_89(n59_13,N1508_6_r_2,G42_7_r_2);
nor I_90(n60_13,n51_13,N1508_0_r_2);
nor I_91(n61_13,n39_13,n_572_7_r_2);
endmodule


