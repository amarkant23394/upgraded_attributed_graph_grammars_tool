module test_I3310(I1351,I2759,I1431,I1470,I1359,I1407,I3310);
input I1351,I2759,I1431,I1470,I1359,I1407;
output I3310;
wire I3217,I3293,I3200,I2844,I2827,I2776;
not I_0(I3217,I3200);
not I_1(I3293,I3217);
DFFARX1 I_2(I1431,I1470,I2759,,,I3200,);
and I_3(I3310,I2844,I3293);
nand I_4(I2844,I2827,I1359);
nor I_5(I2827,I2776,I1351);
not I_6(I2776,I1407);
endmodule


