module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_7_r_4,n6_4,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_4,n25_4,N6147_2_r_11);
not I_43(N1508_0_r_4,n25_4);
nor I_44(N1507_6_r_4,n32_4,n33_4);
nor I_45(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_46(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_47(n_572_7_r_4,n_573_7_r_4);
nand I_48(n_573_7_r_4,n21_4,n22_4);
nor I_49(n_549_7_r_4,n24_4,N6147_2_r_11);
nand I_50(n_569_7_r_4,n22_4,n23_4);
nor I_51(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_52(N6147_9_r_4,n28_4);
nor I_53(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_54(I_BUFF_1_9_r_4,n21_4);
nor I_55(n4_7_r_4,N6147_9_r_4,N6147_2_r_11);
not I_56(n6_4,blif_reset_net_7_r_4);
nand I_57(n21_4,n39_4,n40_4);
or I_58(n22_4,n31_4,N1508_10_r_11);
not I_59(n23_4,N6147_2_r_11);
nor I_60(n24_4,n25_4,n26_4);
nand I_61(n25_4,N1372_1_r_11,N6147_2_r_11);
nand I_62(n26_4,n21_4,n27_4);
nand I_63(n27_4,n36_4,n37_4);
nand I_64(n28_4,n38_4,N1508_1_r_11);
nand I_65(n29_4,N1508_0_r_4,n30_4);
nand I_66(n30_4,n34_4,n35_4);
nor I_67(n31_4,n_429_or_0_5_r_11,N6147_3_r_11);
not I_68(n32_4,n30_4);
nor I_69(n33_4,n21_4,n28_4);
nand I_70(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_71(n35_4,N1508_0_r_4,n27_4);
not I_72(n36_4,N1508_6_r_11);
nand I_73(n37_4,G78_5_r_11,n_547_5_r_11);
or I_74(n38_4,n_429_or_0_5_r_11,N6147_3_r_11);
nor I_75(n39_4,n_576_5_r_11,N1508_1_r_11);
or I_76(n40_4,n41_4,N1372_1_r_11);
nor I_77(n41_4,N6147_3_r_11,N1507_6_r_11);
endmodule


