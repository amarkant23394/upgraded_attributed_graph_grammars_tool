module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_14,blif_reset_net_1_r_14,G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_14,blif_reset_net_1_r_14;
output G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_452_1_r_14,n4_1_l_14,n3_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_14,n3_14,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_14,n3_14,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_14,n3_14,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_14,n3_14,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_14,n3_14,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n_452_1_r_14,blif_clk_net_1_r_14,n3_14,G42_1_r_14,);
and I_33(n_572_1_r_14,n18_14,n19_14);
nand I_34(n_573_1_r_14,n16_14,n17_14);
nor I_35(n_549_1_r_14,n20_14,n21_14);
or I_36(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_37(n_452_1_r_14,n23_14,n_549_1_r_16);
nor I_38(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_39(N3_2_r_14,blif_clk_net_1_r_14,n3_14,G199_2_r_14,);
DFFARX1 I_40(n_572_1_l_14,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_14,);
not I_41(P6_5_r_14,P6_5_r_internal_14);
nor I_42(n4_1_l_14,n_573_1_r_16,G42_1_r_16);
not I_43(n3_14,blif_reset_net_1_r_14);
DFFARX1 I_44(n4_1_l_14,blif_clk_net_1_r_14,n3_14,n15_internal_14,);
not I_45(n15_14,n15_internal_14);
DFFARX1 I_46(ACVQN1_5_r_16,blif_clk_net_1_r_14,n3_14,ACVQN2_3_l_14,);
DFFARX1 I_47(P6_5_r_16,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_14,);
and I_48(N3_2_r_14,n26_14,n27_14);
nor I_49(n_572_1_l_14,n_452_1_r_16,G214_4_r_16);
DFFARX1 I_50(ACVQN2_3_l_14,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_14,);
nor I_51(n16_14,n_549_1_r_16,G199_4_r_16);
not I_52(n17_14,n_572_1_l_14);
nor I_53(n18_14,n_572_1_r_16,G199_4_r_16);
nand I_54(n19_14,ACVQN1_3_l_14,n_569_1_r_16);
nor I_55(n20_14,n_572_1_r_16,n_573_1_r_16);
nor I_56(n21_14,n15_14,n22_14);
nand I_57(n22_14,n24_14,n25_14);
nand I_58(n23_14,n15_14,n24_14);
not I_59(n24_14,G199_4_r_16);
not I_60(n25_14,n_572_1_r_16);
nor I_61(n26_14,n20_14,n_549_1_r_16);
nand I_62(n27_14,n28_14,G42_1_r_16);
not I_63(n28_14,n_452_1_r_16);
endmodule


