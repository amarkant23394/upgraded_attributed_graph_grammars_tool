module test_I3155(I1351,I1447,I2946,I1477,I1470,I2980,I3155);
input I1351,I1447,I2946,I1477,I1470,I2980;
output I3155;
wire I2759,I3011,I3045,I3076,I3028,I2963,I2861;
not I_0(I2759,I1477);
not I_1(I3011,I2980);
and I_2(I3045,I2861,I3028);
or I_3(I3155,I3076,I3045);
DFFARX1 I_4(I1447,I1470,I2759,,,I3076,);
nor I_5(I3028,I2963,I3011);
DFFARX1 I_6(I2946,I1470,I2759,,,I2963,);
not I_7(I2861,I1351);
endmodule


