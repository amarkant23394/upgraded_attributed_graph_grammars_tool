module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_5_r_15,n9_15,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_5_r_15,n9_15,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_5_r_15,n9_15,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_5_r_15,n9_15,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
and I_43(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_44(N1508_0_r_15,n55_15,n_42_8_r_9);
nor I_45(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_46(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_47(N1372_4_r_15,n39_15);
nor I_48(N1508_4_r_15,n39_15,n43_15);
nand I_49(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_50(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_51(n_576_5_r_15,n31_15,n32_15);
not I_52(n_102_5_r_15,n33_15);
nand I_53(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_54(N1507_6_r_15,n42_15,n46_15);
nand I_55(N1508_6_r_15,n39_15,n40_15);
nand I_56(n_431_5_r_15,n36_15,n37_15);
not I_57(n9_15,blif_reset_net_5_r_15);
nor I_58(n31_15,n33_15,n34_15);
nor I_59(n32_15,n44_15,N6134_9_r_9);
nor I_60(n33_15,n54_15,n55_15);
nand I_61(n34_15,n49_15,N1372_4_r_9);
nand I_62(n35_15,N6147_9_r_9,n_576_5_r_9);
not I_63(n36_15,n32_15);
nand I_64(n37_15,n34_15,n38_15);
not I_65(n38_15,n46_15);
nand I_66(n39_15,n38_15,n41_15);
nand I_67(n40_15,n41_15,n42_15);
and I_68(n41_15,n51_15,G199_8_r_9);
and I_69(n42_15,n47_15,n_576_5_r_9);
and I_70(n43_15,n34_15,n36_15);
or I_71(n44_15,N1372_4_r_9,N1508_4_r_9);
not I_72(n45_15,N1372_1_r_15);
nand I_73(n46_15,n53_15,n_576_5_r_9);
nor I_74(n47_15,n34_15,n48_15);
not I_75(n48_15,N6147_9_r_9);
and I_76(n49_15,n50_15,n_576_5_r_9);
nand I_77(n50_15,n51_15,n52_15);
nand I_78(n51_15,N6147_2_r_9,N1508_4_r_9);
not I_79(n52_15,G199_8_r_9);
nor I_80(n53_15,n48_15,n_547_5_r_9);
nor I_81(n54_15,N6147_2_r_9,G78_5_r_9);
not I_82(n55_15,G78_5_r_9);
endmodule


