module test_I13426(I1477,I11895,I1470,I11395,I11460,I13426);
input I1477,I11895,I1470,I11395,I11460;
output I13426;
wire I11287,I11559,I11281,I11593,I13197,I11284,I13392,I11310,I13409;
DFFARX1 I_0(I11895,I1470,I11310,,,I11287,);
DFFARX1 I_1(I1470,I11310,,,I11559,);
not I_2(I11281,I11593);
DFFARX1 I_3(I11559,I1470,I11310,,,I11593,);
not I_4(I13197,I1477);
DFFARX1 I_5(I13409,I1470,I13197,,,I13426,);
nand I_6(I11284,I11395,I11460);
nand I_7(I13392,I11287,I11284);
not I_8(I11310,I1477);
and I_9(I13409,I13392,I11281);
endmodule


