module test_I3951(I1431,I4164,I1447,I2844,I2980,I1470_clk,I1477_rst,I3951);
input I1431,I4164,I1447,I2844,I2980,I1470_clk,I1477_rst;
output I3951;
wire I3310,I3983_rst,I3076,I4229,I4113,I3217,I3107,I4246,I3200,I2759_rst,I2745,I4263,I4181,I2751,I4212,I2733;
and I_0(I3310,I2844);
not I_1(I3983_rst,I1477_rst);
DFFARX1 I_2 (I1447,I1470_clk,I2759_rst,I3076);
nor I_3(I4229,I4113,I4212);
DFFARX1 I_4 (I2751,I1470_clk,I3983_rst,I4113);
not I_5(I3217,I3200);
nor I_6(I3107,I3076,I2844);
DFFARX1 I_7 (I2745,I1470_clk,I3983_rst,I4246);
DFFARX1 I_8 (I1431,I1470_clk,I2759_rst,I3200);
not I_9(I2759_rst,I1477_rst);
nor I_10(I2745,I2980,I3310);
and I_11(I4263,I4246,I2733);
DFFARX1 I_12 (I4164,I1470_clk,I3983_rst,I4181);
nor I_13(I2751,I3076,I3217);
not I_14(I4212,I4181);
nand I_15(I2733,I3217,I3107);
nand I_16(I3951,I4263,I4229);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule