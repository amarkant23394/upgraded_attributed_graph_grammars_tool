module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_3_r_13,blif_reset_net_3_r_13,n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13);
input IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_3_r_13,blif_reset_net_3_r_13;
output n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13;
wire ACVQN2_0_r_14,n_266_and_0_0_r_14,G199_1_r_14,G214_1_r_14,ACVQN1_2_r_14,P6_2_r_14,n_429_or_0_3_r_14,G78_3_r_14,n_576_3_r_14,n_102_3_r_14,n_547_3_r_14,ACVQN2_0_l_14,n_266_and_0_0_l_14,ACVQN1_0_l_14,N1_1_l_14,G199_1_l_14,G214_1_l_14,n3_1_l_14,n_42_5_l_14,N3_5_l_14,G199_5_l_14,n3_5_l_14,ACVQN1_0_r_14,N1_1_r_14,n3_1_r_14,P6_internal_2_r_14,n12_3_r_14,n_431_3_r_14,n11_3_r_14,n13_3_r_14,n14_3_r_14,n15_3_r_14,n16_3_r_14,n2_3_r_13,ACVQN1_2_l_13,P6_2_l_13,P6_internal_2_l_13,n_429_or_0_3_l_13,n12_3_l_13,n_431_3_l_13,G78_3_l_13,n_576_3_l_13,n11_3_l_13,n_102_3_l_13,n_547_3_l_13,n13_3_l_13,n14_3_l_13,n15_3_l_13,n16_3_l_13,n12_3_r_13,n_431_3_r_13,n11_3_r_13,n13_3_r_13,n14_3_r_13,n15_3_r_13,n16_3_r_13,n4_4_r_13,n_87_4_r_13,n7_4_r_13;
DFFARX1 I_0(n_266_and_0_0_l_14,blif_clk_net_3_r_13,n2_3_r_13,ACVQN2_0_r_14,);
and I_1(n_266_and_0_0_r_14,G199_5_l_14,ACVQN1_0_r_14);
DFFARX1 I_2(N1_1_r_14,blif_clk_net_3_r_13,n2_3_r_13,G199_1_r_14,);
DFFARX1 I_3(G199_1_l_14,blif_clk_net_3_r_13,n2_3_r_13,G214_1_r_14,);
DFFARX1 I_4(ACVQN2_0_l_14,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_r_14,);
not I_5(P6_2_r_14,P6_internal_2_r_14);
nand I_6(n_429_or_0_3_r_14,G214_1_l_14,n12_3_r_14);
DFFARX1 I_7(n_431_3_r_14,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_14,);
nand I_8(n_576_3_r_14,ACVQN2_0_l_14,n11_3_r_14);
not I_9(n_102_3_r_14,G199_5_l_14);
nand I_10(n_547_3_r_14,n_266_and_0_0_l_14,n13_3_r_14);
DFFARX1 I_11(IN_1_0_l_14,blif_clk_net_3_r_13,n2_3_r_13,ACVQN2_0_l_14,);
and I_12(n_266_and_0_0_l_14,IN_4_0_l_14,ACVQN1_0_l_14);
DFFARX1 I_13(IN_2_0_l_14,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_0_l_14,);
and I_14(N1_1_l_14,IN_6_1_l_14,n3_1_l_14);
DFFARX1 I_15(N1_1_l_14,blif_clk_net_3_r_13,n2_3_r_13,G199_1_l_14,);
DFFARX1 I_16(IN_3_1_l_14,blif_clk_net_3_r_13,n2_3_r_13,G214_1_l_14,);
nand I_17(n3_1_l_14,IN_1_1_l_14,IN_2_1_l_14);
nor I_18(n_42_5_l_14,IN_1_5_l_14,IN_3_5_l_14);
and I_19(N3_5_l_14,IN_6_5_l_14,n3_5_l_14);
DFFARX1 I_20(N3_5_l_14,blif_clk_net_3_r_13,n2_3_r_13,G199_5_l_14,);
nand I_21(n3_5_l_14,IN_2_5_l_14,IN_3_5_l_14);
DFFARX1 I_22(G214_1_l_14,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_0_r_14,);
and I_23(N1_1_r_14,G214_1_l_14,n3_1_r_14);
nand I_24(n3_1_r_14,ACVQN2_0_l_14,n_42_5_l_14);
DFFARX1 I_25(G199_5_l_14,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_r_14,);
not I_26(n12_3_r_14,n_42_5_l_14);
or I_27(n_431_3_r_14,n_266_and_0_0_l_14,n14_3_r_14);
nor I_28(n11_3_r_14,G199_5_l_14,n12_3_r_14);
nor I_29(n13_3_r_14,G199_1_l_14,G199_5_l_14);
and I_30(n14_3_r_14,n_42_5_l_14,n15_3_r_14);
nor I_31(n15_3_r_14,G199_1_l_14,n16_3_r_14);
not I_32(n16_3_r_14,G214_1_l_14);
nand I_33(n_429_or_0_3_r_13,n_429_or_0_3_l_13,n12_3_r_13);
DFFARX1 I_34(n_431_3_r_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_13,);
nand I_35(n_576_3_r_13,n_547_3_l_13,n11_3_r_13);
not I_36(n_102_3_r_13,ACVQN1_2_l_13);
nand I_37(n_547_3_r_13,P6_2_l_13,n13_3_r_13);
DFFARX1 I_38(n4_4_r_13,blif_clk_net_3_r_13,n2_3_r_13,G42_4_r_13,);
nor I_39(n_572_4_r_13,P6_2_l_13,n_429_or_0_3_l_13);
or I_40(n_573_4_r_13,ACVQN1_2_l_13,G78_3_l_13);
nor I_41(n_549_4_r_13,n_429_or_0_3_l_13,n7_4_r_13);
or I_42(n_569_4_r_13,n_429_or_0_3_l_13,G78_3_l_13);
nor I_43(n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13);
not I_44(n2_3_r_13,blif_reset_net_3_r_13);
DFFARX1 I_45(G78_3_r_14,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_l_13,);
not I_46(P6_2_l_13,P6_internal_2_l_13);
DFFARX1 I_47(n_429_or_0_3_r_14,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_l_13,);
nand I_48(n_429_or_0_3_l_13,n12_3_l_13,G214_1_r_14);
not I_49(n12_3_l_13,G199_1_r_14);
or I_50(n_431_3_l_13,n14_3_l_13,ACVQN1_2_r_14);
DFFARX1 I_51(n_431_3_l_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_l_13,);
nand I_52(n_576_3_l_13,n11_3_l_13,n_102_3_r_14);
nor I_53(n11_3_l_13,n12_3_l_13,n_547_3_r_14);
not I_54(n_102_3_l_13,n_547_3_r_14);
nand I_55(n_547_3_l_13,n13_3_l_13,ACVQN2_0_r_14);
nor I_56(n13_3_l_13,P6_2_r_14,n_547_3_r_14);
and I_57(n14_3_l_13,n15_3_l_13,n_576_3_r_14);
nor I_58(n15_3_l_13,n16_3_l_13,n_266_and_0_0_r_14);
not I_59(n16_3_l_13,G214_1_r_14);
not I_60(n12_3_r_13,n_102_3_l_13);
or I_61(n_431_3_r_13,ACVQN1_2_l_13,n14_3_r_13);
nor I_62(n11_3_r_13,ACVQN1_2_l_13,n12_3_r_13);
nor I_63(n13_3_r_13,ACVQN1_2_l_13,n_576_3_l_13);
and I_64(n14_3_r_13,n_102_3_l_13,n15_3_r_13);
nor I_65(n15_3_r_13,G78_3_l_13,n16_3_r_13);
not I_66(n16_3_r_13,n_429_or_0_3_l_13);
nor I_67(n4_4_r_13,P6_2_l_13,n_547_3_l_13);
not I_68(n_87_4_r_13,P6_2_l_13);
and I_69(n7_4_r_13,n_576_3_l_13,n_87_4_r_13);
endmodule


