module test_I1750(I1439,I1367,I1279,I1207,I1750);
input I1439,I1367,I1279,I1207;
output I1750;
wire I1733,I1716,I1699;
or I_0(I1750,I1733,I1279);
and I_1(I1733,I1716,I1439);
nor I_2(I1716,I1699,I1367);
not I_3(I1699,I1207);
endmodule


