module test_I15591(I1477,I11938,I1470,I14278,I15591);
input I1477,I11938,I1470,I14278;
output I15591;
wire I13908,I13752,I13743,I15832,I14162,I16052,I15628,I13749,I13775,I15611,I13891,I16069;
not I_0(I13908,I13891);
DFFARX1 I_1(I14278,I1470,I13775,,,I13752,);
DFFARX1 I_2(I13891,I1470,I13775,,,I13743,);
nand I_3(I15832,I15628,I13749);
DFFARX1 I_4(I11938,I1470,I13775,,,I14162,);
DFFARX1 I_5(I13752,I1470,I15611,,,I16052,);
not I_6(I15628,I13743);
nand I_7(I13749,I14162,I13908);
not I_8(I13775,I1477);
not I_9(I15611,I1477);
DFFARX1 I_10(I1470,I13775,,,I13891,);
nor I_11(I15591,I16069,I15832);
not I_12(I16069,I16052);
endmodule


