module test_I6875(I5450,I1477,I1470,I5563,I5642,I6875);
input I5450,I1477,I1470,I5563,I5642;
output I6875;
wire I5659,I5073,I5088,I6907,I7221,I5105,I6924;
or I_0(I5659,I5642,I5563);
DFFARX1 I_1(I7221,I1470,I6907,,,I6875,);
DFFARX1 I_2(I5450,I1470,I5105,,,I5073,);
DFFARX1 I_3(I5659,I1470,I5105,,,I5088,);
not I_4(I6907,I1477);
nand I_5(I7221,I6924,I5088);
not I_6(I5105,I1477);
not I_7(I6924,I5073);
endmodule


