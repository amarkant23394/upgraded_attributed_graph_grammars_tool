module test_I2554(I2798,I1917,I1294,I1301,I2554);
input I2798,I1917,I1294,I1301;
output I2554;
wire I2815,I2866,I2583,I2832;
or I_0(I2815,I2798,I1917);
not I_1(I2554,I2866);
DFFARX1 I_2(I2832,I1294,I2583,,,I2866,);
not I_3(I2583,I1301);
DFFARX1 I_4(I2815,I1294,I2583,,,I2832,);
endmodule


