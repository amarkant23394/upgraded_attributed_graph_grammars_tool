module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_6,blif_reset_net_1_r_6,G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_6,blif_reset_net_1_r_6;
output G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,N3_2_l_6,n4_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_6,n4_6,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_6,n4_6,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_6,n4_6,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_6,n4_6,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_6,n4_6,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_6,n4_6,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_6,blif_clk_net_1_r_6,n4_6,G42_1_r_6,);
nor I_34(n_572_1_r_6,n27_6,n28_6);
nand I_35(n_573_1_r_6,n18_6,n19_6);
nor I_36(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_37(n_569_1_r_6,n19_6,n20_6);
nor I_38(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_39(N1_4_r_6,blif_clk_net_1_r_6,n4_6,G199_4_r_6,);
DFFARX1 I_40(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,G214_4_r_6,);
DFFARX1 I_41(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_6,);
not I_42(P6_5_r_6,P6_5_r_internal_6);
and I_43(N3_2_l_6,n23_6,ACVQN1_5_r_13);
not I_44(n4_6,blif_reset_net_1_r_6);
DFFARX1 I_45(N3_2_l_6,blif_clk_net_1_r_6,n4_6,n27_6,);
not I_46(n17_6,n27_6);
DFFARX1 I_47(n_266_and_0_3_r_13,blif_clk_net_1_r_6,n4_6,n28_6,);
DFFARX1 I_48(P6_5_r_13,blif_clk_net_1_r_6,n4_6,n26_6,);
and I_49(N1_4_l_6,n25_6,n_573_1_r_13);
DFFARX1 I_50(N1_4_l_6,blif_clk_net_1_r_6,n4_6,n29_6,);
not I_51(n18_6,n29_6);
DFFARX1 I_52(n_572_1_r_13,blif_clk_net_1_r_6,n4_6,G214_4_l_6,);
not I_53(n12_6,G214_4_l_6);
nor I_54(n4_1_r_6,n28_6,n22_6);
nor I_55(N1_4_r_6,n12_6,n24_6);
nor I_56(n_42_2_l_6,n_549_1_r_13,G42_1_r_13);
DFFARX1 I_57(G214_4_l_6,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_6,);
nand I_58(n19_6,n26_6,G42_1_r_13);
not I_59(n20_6,n_42_2_l_6);
nor I_60(n21_6,n17_6,n28_6);
and I_61(n22_6,n26_6,G42_1_r_13);
nand I_62(n23_6,n_549_1_r_13,n_452_1_r_13);
nor I_63(n24_6,n17_6,n18_6);
nand I_64(n25_6,ACVQN2_3_r_13,n_572_1_r_13);
endmodule


