module test_I1908(I1687,I1294,I1954,I1301,I1908);
input I1687,I1294,I1954,I1301;
output I1908;
wire I1316,I2005,I1937,I2022,I2039,I1509,I1310;
nand I_0(I1316,I1509,I1687);
nor I_1(I2005,I1954,I1310);
not I_2(I1937,I1301);
nand I_3(I2022,I2005,I1316);
DFFARX1 I_4(I2022,I1294,I1937,,,I2039,);
not I_5(I1908,I2039);
DFFARX1 I_6(I1294,,,I1509,);
DFFARX1 I_7(I1294,,,I1310,);
endmodule


