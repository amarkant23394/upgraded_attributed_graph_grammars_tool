module test_I15126(I12619,I1470,I12653,I15126);
input I12619,I1470,I12653;
output I15126;
wire I12670,I12783,I12584,I15109,I12735;
DFFARX1 I_0(I12653,I1470,I12619,,,I12670,);
DFFARX1 I_1(I12735,I1470,I12619,,,I12783,);
and I_2(I12584,I12670,I12783);
not I_3(I15109,I12584);
DFFARX1 I_4(I1470,I12619,,,I12735,);
not I_5(I15126,I15109);
endmodule


