module test_I3413(I2234,I1294,I1301,I3413);
input I2234,I1294,I1301;
output I3413;
wire I2583,I1902,I2203,I2566,I2945;
not I_0(I2583,I1301);
and I_1(I1902,I2234,I2203);
not I_2(I3413,I2566);
DFFARX1 I_3(I1294,,,I2203,);
not I_4(I2566,I2945);
DFFARX1 I_5(I1902,I1294,I2583,,,I2945,);
endmodule


