module test_I13102(I9477,I9465,I1477,I12814,I10618,I1470,I12653,I13102);
input I9477,I9465,I1477,I12814,I10618,I1470,I12653;
output I13102;
wire I12619,I12670,I10715,I13023,I12831,I12687,I12865,I10766,I10636,I10732,I12848;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
nor I_2(I10715,I9477);
DFFARX1 I_3(I10636,I1470,I12619,,,I13023,);
and I_4(I12831,I12814,I10618);
not I_5(I12687,I12670);
nor I_6(I12865,I12848,I12687);
and I_7(I13102,I13023,I12865);
not I_8(I10766,I9477);
nor I_9(I10636,I10732,I10766);
nand I_10(I10732,I10715,I9465);
DFFARX1 I_11(I12831,I1470,I12619,,,I12848,);
endmodule


