module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_8_r_8,n8_8,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_8_r_8,n8_8,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_8,n46_8,n51_8);
not I_41(N1508_0_r_8,n46_8);
nor I_42(N1372_1_r_8,n37_8,n49_8);
and I_43(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_44(N1507_6_r_8,n47_8,n48_8);
nor I_45(N1508_6_r_8,n37_8,n38_8);
nor I_46(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_47(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_48(N6147_9_r_8,n29_8,n30_8);
nor I_49(N6134_9_r_8,n30_8,n31_8);
not I_50(I_BUFF_1_9_r_8,n35_8);
nor I_51(N1372_10_r_8,n46_8,n49_8);
nor I_52(N1508_10_r_8,n40_8,n41_8);
and I_53(N3_8_l_8,n36_8,n_452_7_r_16);
not I_54(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_55(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_56(n29_8,n53_8);
nor I_57(N3_8_r_8,n33_8,n34_8);
and I_58(n30_8,n32_8,n33_8);
nor I_59(n31_8,N1508_1_r_16,G42_7_r_16);
nand I_60(n32_8,n42_8,n_572_7_r_16);
or I_61(n33_8,n46_8,N1507_6_r_16);
nor I_62(n34_8,n32_8,n35_8);
nand I_63(n35_8,n44_8,N1371_0_r_16);
nand I_64(n36_8,G42_7_r_16,n_573_7_r_16);
not I_65(n37_8,n31_8);
nand I_66(n38_8,N1508_0_r_8,n39_8);
nand I_67(n39_8,n33_8,n50_8);
and I_68(n40_8,n32_8,n35_8);
not I_69(n41_8,N1372_10_r_8);
and I_70(n42_8,n43_8,n_569_7_r_16);
nand I_71(n43_8,n44_8,n45_8);
nand I_72(n44_8,N1371_0_r_16,N1372_1_r_16);
not I_73(n45_8,N1371_0_r_16);
nand I_74(n46_8,N6147_2_r_16,N1508_0_r_16);
not I_75(n47_8,n39_8);
nor I_76(n48_8,n35_8,n49_8);
not I_77(n49_8,n51_8);
nand I_78(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_79(n51_8,n52_8,N1372_1_r_16);
or I_80(n52_8,N1508_0_r_16,N1508_6_r_16);
endmodule


