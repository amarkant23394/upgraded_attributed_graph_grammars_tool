module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9);
input IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9;
wire ACVQN2_0_r_14,n_266_and_0_0_r_14,G199_1_r_14,G214_1_r_14,ACVQN1_2_r_14,P6_2_r_14,n_429_or_0_3_r_14,G78_3_r_14,n_576_3_r_14,n_102_3_r_14,n_547_3_r_14,ACVQN2_0_l_14,n_266_and_0_0_l_14,ACVQN1_0_l_14,N1_1_l_14,G199_1_l_14,G214_1_l_14,n3_1_l_14,n_42_5_l_14,N3_5_l_14,G199_5_l_14,n3_5_l_14,ACVQN1_0_r_14,N1_1_r_14,n3_1_r_14,P6_internal_2_r_14,n12_3_r_14,n_431_3_r_14,n11_3_r_14,n13_3_r_14,n14_3_r_14,n15_3_r_14,n16_3_r_14,n1_1_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9,ACVQN1_0_l_9,n4_4_l_9,G42_4_l_9,n_87_4_l_9,n_572_4_l_9,n_573_4_l_9,n_549_4_l_9,n7_4_l_9,n_569_4_l_9,n_452_4_l_9,N1_1_r_9,n3_1_r_9,P6_internal_2_r_9,n12_3_r_9,n_431_3_r_9,n11_3_r_9,n13_3_r_9,n14_3_r_9,n15_3_r_9,n16_3_r_9,N3_5_r_9,n3_5_r_9;
DFFARX1 I_0(n_266_and_0_0_l_14,blif_clk_net_1_r_9,n1_1_r_9,ACVQN2_0_r_14,);
and I_1(n_266_and_0_0_r_14,G199_5_l_14,ACVQN1_0_r_14);
DFFARX1 I_2(N1_1_r_14,blif_clk_net_1_r_9,n1_1_r_9,G199_1_r_14,);
DFFARX1 I_3(G199_1_l_14,blif_clk_net_1_r_9,n1_1_r_9,G214_1_r_14,);
DFFARX1 I_4(ACVQN2_0_l_14,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_2_r_14,);
not I_5(P6_2_r_14,P6_internal_2_r_14);
nand I_6(n_429_or_0_3_r_14,G214_1_l_14,n12_3_r_14);
DFFARX1 I_7(n_431_3_r_14,blif_clk_net_1_r_9,n1_1_r_9,G78_3_r_14,);
nand I_8(n_576_3_r_14,ACVQN2_0_l_14,n11_3_r_14);
not I_9(n_102_3_r_14,G199_5_l_14);
nand I_10(n_547_3_r_14,n_266_and_0_0_l_14,n13_3_r_14);
DFFARX1 I_11(IN_1_0_l_14,blif_clk_net_1_r_9,n1_1_r_9,ACVQN2_0_l_14,);
and I_12(n_266_and_0_0_l_14,IN_4_0_l_14,ACVQN1_0_l_14);
DFFARX1 I_13(IN_2_0_l_14,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_0_l_14,);
and I_14(N1_1_l_14,IN_6_1_l_14,n3_1_l_14);
DFFARX1 I_15(N1_1_l_14,blif_clk_net_1_r_9,n1_1_r_9,G199_1_l_14,);
DFFARX1 I_16(IN_3_1_l_14,blif_clk_net_1_r_9,n1_1_r_9,G214_1_l_14,);
nand I_17(n3_1_l_14,IN_1_1_l_14,IN_2_1_l_14);
nor I_18(n_42_5_l_14,IN_1_5_l_14,IN_3_5_l_14);
and I_19(N3_5_l_14,IN_6_5_l_14,n3_5_l_14);
DFFARX1 I_20(N3_5_l_14,blif_clk_net_1_r_9,n1_1_r_9,G199_5_l_14,);
nand I_21(n3_5_l_14,IN_2_5_l_14,IN_3_5_l_14);
DFFARX1 I_22(G214_1_l_14,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_0_r_14,);
and I_23(N1_1_r_14,G214_1_l_14,n3_1_r_14);
nand I_24(n3_1_r_14,ACVQN2_0_l_14,n_42_5_l_14);
DFFARX1 I_25(G199_5_l_14,blif_clk_net_1_r_9,n1_1_r_9,P6_internal_2_r_14,);
not I_26(n12_3_r_14,n_42_5_l_14);
or I_27(n_431_3_r_14,n_266_and_0_0_l_14,n14_3_r_14);
nor I_28(n11_3_r_14,G199_5_l_14,n12_3_r_14);
nor I_29(n13_3_r_14,G199_1_l_14,G199_5_l_14);
and I_30(n14_3_r_14,n_42_5_l_14,n15_3_r_14);
nor I_31(n15_3_r_14,G199_1_l_14,n16_3_r_14);
not I_32(n16_3_r_14,G214_1_l_14);
DFFARX1 I_33(N1_1_r_9,blif_clk_net_1_r_9,n1_1_r_9,G199_1_r_9,);
DFFARX1 I_34(G42_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,G214_1_r_9,);
DFFARX1 I_35(n_572_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_2_r_9,);
not I_36(P6_2_r_9,P6_internal_2_r_9);
nand I_37(n_429_or_0_3_r_9,n_572_4_l_9,n12_3_r_9);
DFFARX1 I_38(n_431_3_r_9,blif_clk_net_1_r_9,n1_1_r_9,G78_3_r_9,);
nand I_39(n_576_3_r_9,n_573_4_l_9,n11_3_r_9);
not I_40(n_102_3_r_9,n_266_and_0_0_l_9);
nand I_41(n_547_3_r_9,n_549_4_l_9,n13_3_r_9);
nor I_42(n_42_5_r_9,n_569_4_l_9,n_452_4_l_9);
DFFARX1 I_43(N3_5_r_9,blif_clk_net_1_r_9,n1_1_r_9,G199_5_r_9,);
not I_44(n1_1_r_9,blif_reset_net_1_r_9);
DFFARX1 I_45(n_576_3_r_14,blif_clk_net_1_r_9,n1_1_r_9,ACVQN2_0_l_9,);
and I_46(n_266_and_0_0_l_9,ACVQN1_0_l_9,n_102_3_r_14);
DFFARX1 I_47(n_547_3_r_14,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_0_l_9,);
nor I_48(n4_4_l_9,ACVQN1_2_r_14,n_429_or_0_3_r_14);
DFFARX1 I_49(n4_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,G42_4_l_9,);
not I_50(n_87_4_l_9,G199_1_r_14);
nor I_51(n_572_4_l_9,n_266_and_0_0_r_14,G199_1_r_14);
or I_52(n_573_4_l_9,ACVQN2_0_r_14,G214_1_r_14);
nor I_53(n_549_4_l_9,n7_4_l_9,P6_2_r_14);
and I_54(n7_4_l_9,n_87_4_l_9,G78_3_r_14);
or I_55(n_569_4_l_9,ACVQN2_0_r_14,P6_2_r_14);
nor I_56(n_452_4_l_9,G214_1_r_14,ACVQN1_2_r_14);
and I_57(N1_1_r_9,n_266_and_0_0_l_9,n3_1_r_9);
nand I_58(n3_1_r_9,n_572_4_l_9,n_569_4_l_9);
DFFARX1 I_59(n_266_and_0_0_l_9,blif_clk_net_1_r_9,n1_1_r_9,P6_internal_2_r_9,);
not I_60(n12_3_r_9,G42_4_l_9);
or I_61(n_431_3_r_9,n_549_4_l_9,n14_3_r_9);
nor I_62(n11_3_r_9,ACVQN2_0_l_9,n12_3_r_9);
nor I_63(n13_3_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9);
and I_64(n14_3_r_9,n_452_4_l_9,n15_3_r_9);
nor I_65(n15_3_r_9,G42_4_l_9,n16_3_r_9);
not I_66(n16_3_r_9,n_572_4_l_9);
and I_67(N3_5_r_9,ACVQN2_0_l_9,n3_5_r_9);
nand I_68(n3_5_r_9,n_573_4_l_9,n_452_4_l_9);
endmodule


