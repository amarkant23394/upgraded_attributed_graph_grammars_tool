module test_final(IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_5_r_4,blif_reset_net_5_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4);
input IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_5_r_4,blif_reset_net_5_r_4;
output N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4;
wire N1371_0_r_0,N1508_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0,N3_8_l_0,n40_0,n4_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,N1371_0_r_4,n_102_5_r_4,n_431_5_r_4,n4_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4;
nor I_0(N1371_0_r_0,n24_0,n25_0);
not I_1(N1508_0_r_0,n25_0);
nor I_2(N6147_2_r_0,n28_0,n29_0);
nand I_3(n_429_or_0_5_r_0,n4_0,n25_0);
DFFARX1 I_4(n4_0,blif_clk_net_5_r_4,n4_4,G78_5_r_0,);
nand I_5(n_576_5_r_0,n23_0,n24_0);
not I_6(n_102_5_r_0,n40_0);
nand I_7(n_547_5_r_0,n26_0,n27_0);
nor I_8(N1507_6_r_0,n_102_5_r_0,n37_0);
nor I_9(N1508_6_r_0,n25_0,n33_0);
and I_10(N3_8_l_0,IN_6_8_l_0,n32_0);
DFFARX1 I_11(N3_8_l_0,blif_clk_net_5_r_4,n4_4,n40_0,);
not I_12(n4_0,n31_0);
nor I_13(n23_0,n40_0,n25_0);
and I_14(n24_0,n4_0,n39_0);
nand I_15(n25_0,IN_1_1_l_0,IN_2_1_l_0);
nor I_16(n26_0,n40_0,n24_0);
nor I_17(n27_0,IN_1_8_l_0,IN_3_8_l_0);
nor I_18(n28_0,IN_3_1_l_0,n25_0);
nand I_19(n29_0,n_102_5_r_0,n30_0);
nand I_20(n30_0,n27_0,n31_0);
nand I_21(n31_0,IN_1_10_l_0,IN_2_10_l_0);
nand I_22(n32_0,IN_2_8_l_0,IN_3_8_l_0);
nand I_23(n33_0,n34_0,n35_0);
nand I_24(n34_0,n_102_5_r_0,n36_0);
not I_25(n35_0,IN_3_1_l_0);
not I_26(n36_0,n27_0);
nor I_27(n37_0,n36_0,n38_0);
nand I_28(n38_0,N1508_0_r_0,n35_0);
or I_29(n39_0,IN_3_10_l_0,IN_4_10_l_0);
nor I_30(N1371_0_r_4,n25_4,n29_4);
nor I_31(N1508_0_r_4,n25_4,n32_4);
nor I_32(N6147_2_r_4,n24_4,n31_4);
or I_33(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_34(n_431_5_r_4,blif_clk_net_5_r_4,n4_4,G78_5_r_4,);
nand I_35(n_576_5_r_4,n22_4,n23_4);
nand I_36(n_102_5_r_4,n34_4,n35_4);
nand I_37(n_547_5_r_4,n26_4,n27_4);
nor I_38(N1507_6_r_4,n27_4,n30_4);
nor I_39(N1508_6_r_4,n30_4,n33_4);
nand I_40(n_431_5_r_4,n_102_5_r_4,n28_4);
not I_41(n4_4,blif_reset_net_5_r_4);
nor I_42(n22_4,n24_4,n25_4);
nor I_43(n23_4,n37_4,N1371_0_r_0);
not I_44(n24_4,n_102_5_r_4);
nand I_45(n25_4,G78_5_r_0,N1508_6_r_0);
nor I_46(n26_4,n23_4,n24_4);
not I_47(n27_4,n25_4);
nand I_48(n28_4,n23_4,n29_4);
nor I_49(n29_4,n25_4,n_429_or_0_5_r_0);
not I_50(n30_4,n29_4);
nor I_51(n31_4,N1371_0_r_4,n32_4);
nor I_52(n32_4,n23_4,n29_4);
nand I_53(n33_4,n23_4,n24_4);
nor I_54(n34_4,N6147_2_r_0,n_429_or_0_5_r_0);
or I_55(n35_4,n36_4,N1507_6_r_0);
nor I_56(n36_4,n_576_5_r_0,N1371_0_r_0);
or I_57(n37_4,N6147_2_r_0,n_547_5_r_0);
endmodule


