module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_8_r_8,n8_8,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_8,n46_8,n51_8);
not I_37(N1508_0_r_8,n46_8);
nor I_38(N1372_1_r_8,n37_8,n49_8);
and I_39(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_40(N1507_6_r_8,n47_8,n48_8);
nor I_41(N1508_6_r_8,n37_8,n38_8);
nor I_42(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_43(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_44(N6147_9_r_8,n29_8,n30_8);
nor I_45(N6134_9_r_8,n30_8,n31_8);
not I_46(I_BUFF_1_9_r_8,n35_8);
nor I_47(N1372_10_r_8,n46_8,n49_8);
nor I_48(N1508_10_r_8,n40_8,n41_8);
and I_49(N3_8_l_8,n36_8,G42_7_r_3);
not I_50(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_51(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_52(n29_8,n53_8);
nor I_53(N3_8_r_8,n33_8,n34_8);
and I_54(n30_8,n32_8,n33_8);
nor I_55(n31_8,n_549_7_r_3,N1507_6_r_3);
nand I_56(n32_8,n42_8,N1508_6_r_3);
or I_57(n33_8,n46_8,N1508_1_r_3);
nor I_58(n34_8,n32_8,n35_8);
nand I_59(n35_8,n44_8,n_452_7_r_3);
nand I_60(n36_8,n_549_7_r_3,N1372_1_r_3);
not I_61(n37_8,n31_8);
nand I_62(n38_8,N1508_0_r_8,n39_8);
nand I_63(n39_8,n33_8,n50_8);
and I_64(n40_8,n32_8,n35_8);
not I_65(n41_8,N1372_10_r_8);
and I_66(n42_8,n43_8,N1508_6_r_3);
nand I_67(n43_8,n44_8,n45_8);
nand I_68(n44_8,N1372_1_r_3,n_569_7_r_3);
not I_69(n45_8,n_452_7_r_3);
nand I_70(n46_8,n_573_7_r_3,N6134_9_r_3);
not I_71(n47_8,n39_8);
nor I_72(n48_8,n35_8,n49_8);
not I_73(n49_8,n51_8);
nand I_74(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_75(n51_8,n52_8,G42_7_r_3);
or I_76(n52_8,N1507_6_r_3,N1508_1_r_3);
endmodule


