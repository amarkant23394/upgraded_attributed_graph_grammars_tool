module test_I17402(I15696,I15628,I15579,I13749,I1470,I16145,I15611,I15798,I17402);
input I15696,I15628,I15579,I13749,I1470,I16145,I15611,I15798;
output I17402;
wire I17430,I15597,I15600,I17532,I15832,I15815,I17481,I16162,I17498;
not I_0(I17430,I15579);
nor I_1(I15597,I15832,I16162);
nor I_2(I17402,I17498,I17532);
or I_3(I15600,I15832,I15815);
not I_4(I17532,I15597);
nand I_5(I15832,I15628,I13749);
DFFARX1 I_6(I15798,I1470,I15611,,,I15815,);
nor I_7(I17481,I17430,I15597);
and I_8(I16162,I15696,I16145);
nand I_9(I17498,I17481,I15600);
endmodule


