module test_I14951(I1477,I15177,I1470,I14951);
input I1477,I15177,I1470;
output I14951;
wire I12670,I12783,I12930,I12752,I14965,I12581,I12590,I12608,I15194,I12619,I12913,I15109,I15211,I15016,I12584,I14999,I15126,I15245,I10609;
DFFARX1 I_0(I1470,I12619,,,I12670,);
DFFARX1 I_1(I1470,I12619,,,I12783,);
and I_2(I12930,I12913,I10609);
nand I_3(I14951,I15016,I15245);
DFFARX1 I_4(I1470,I12619,,,I12752,);
not I_5(I14965,I1477);
DFFARX1 I_6(I12930,I1470,I12619,,,I12581,);
not I_7(I12590,I12752);
nor I_8(I12608,I12930);
or I_9(I15194,I15177,I12608);
not I_10(I12619,I1477);
DFFARX1 I_11(I1470,I12619,,,I12913,);
not I_12(I15109,I12584);
DFFARX1 I_13(I15194,I1470,I14965,,,I15211,);
nand I_14(I15016,I14999,I12581);
and I_15(I12584,I12670,I12783);
nor I_16(I14999,I12584,I12590);
not I_17(I15126,I15109);
nor I_18(I15245,I15211,I15126);
DFFARX1 I_19(I1470,,,I10609,);
endmodule


