module test_I1897(I1455,I1477,I1215,I1423,I1470,I1383,I1897);
input I1455,I1477,I1215,I1423,I1470,I1383;
output I1897;
wire I1518,I1880,I1586,I1603,I1535;
not I_0(I1518,I1477);
DFFARX1 I_1(I1383,I1470,I1518,,,I1880,);
nor I_2(I1586,I1535,I1215);
nand I_3(I1603,I1586,I1423);
not I_4(I1535,I1455);
nor I_5(I1897,I1880,I1603);
endmodule


