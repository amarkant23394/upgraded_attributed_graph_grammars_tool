module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_7_r_16,n8_16,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_7_r_16,n8_16,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_7_r_16,n8_16,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_7_r_16,n8_16,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
nor I_43(N1371_0_r_16,n35_16,n39_16);
nor I_44(N1508_0_r_16,n39_16,n46_16);
not I_45(N1372_1_r_16,n45_16);
nor I_46(N1508_1_r_16,n53_16,n45_16);
nor I_47(N6147_2_r_16,n37_16,n38_16);
nor I_48(N1507_6_r_16,n44_16,n49_16);
nor I_49(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_50(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_51(n_572_7_r_16,n32_16,n33_16);
nand I_52(n_573_7_r_16,n30_16,n31_16);
nand I_53(n_549_7_r_16,n47_16,G78_5_r_9);
nand I_54(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_55(n_452_7_r_16,n34_16,n35_16);
and I_56(N3_8_l_16,n41_16,G78_5_r_9);
not I_57(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_58(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_59(n29_16,n53_16);
nor I_60(n4_7_r_16,n35_16,n36_16);
nand I_61(n30_16,n_547_5_r_9,N6147_9_r_9);
not I_62(n31_16,n34_16);
nor I_63(n32_16,n30_16,N1372_4_r_9);
not I_64(n33_16,n_549_7_r_16);
nor I_65(n34_16,n48_16,G199_8_r_9);
and I_66(n35_16,n50_16,N1508_4_r_9);
not I_67(n36_16,n30_16);
nor I_68(n37_16,n31_16,n40_16);
nand I_69(n38_16,n29_16,n39_16);
not I_70(n39_16,n32_16);
nor I_71(n40_16,n_576_5_r_9,n_42_8_r_9);
nand I_72(n41_16,n_42_8_r_9,N6147_2_r_9);
nand I_73(n42_16,n35_16,n43_16);
not I_74(n43_16,n44_16);
nor I_75(n44_16,n32_16,n49_16);
nand I_76(n45_16,n36_16,n40_16);
nor I_77(n46_16,n33_16,n34_16);
nand I_78(n47_16,N1372_4_r_9,N6134_9_r_9);
or I_79(n48_16,N6147_2_r_9,N1508_4_r_9);
and I_80(n49_16,n35_16,n36_16);
and I_81(n50_16,n51_16,n_576_5_r_9);
nand I_82(n51_16,n47_16,n52_16);
not I_83(n52_16,G78_5_r_9);
endmodule


