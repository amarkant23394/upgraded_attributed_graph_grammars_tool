module test_I13119(I10664,I1477,I12831,I10766,I9459,I10732,I1470,I13119);
input I10664,I1477,I12831,I10766,I9459,I10732,I1470;
output I13119;
wire I10647,I12670,I12865,I10961,I13102,I10639,I12848,I13023,I12718,I11184,I10636,I12619,I12687,I10615,I11201;
not I_0(I10647,I1477);
DFFARX1 I_1(I1470,I12619,,,I12670,);
nor I_2(I12865,I12848,I12687);
nand I_3(I10961,I10664,I9459);
and I_4(I13102,I13023,I12865);
DFFARX1 I_5(I11201,I1470,I10647,,,I10639,);
DFFARX1 I_6(I12831,I1470,I12619,,,I12848,);
DFFARX1 I_7(I10636,I1470,I12619,,,I13023,);
nor I_8(I12718,I10615,I10639);
nand I_9(I11184,I10732);
or I_10(I13119,I12718,I13102);
nor I_11(I10636,I10732,I10766);
not I_12(I12619,I1477);
not I_13(I12687,I12670);
DFFARX1 I_14(I10961,I1470,I10647,,,I10615,);
and I_15(I11201,I10961,I11184);
endmodule


