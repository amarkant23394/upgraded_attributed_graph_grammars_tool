module test_I1750(I1367,I1279,I1439,I1207,I1750);
input I1367,I1279,I1439,I1207;
output I1750;
wire I1716,I1733,I1699;
nor I_0(I1716,I1699,I1367);
and I_1(I1733,I1716,I1439);
or I_2(I1750,I1733,I1279);
not I_3(I1699,I1207);
endmodule


