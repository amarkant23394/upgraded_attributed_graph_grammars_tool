module test_final(a_0_ran_l,b_0_ran_l,A0_3_ran_l,A1_3_ran_l,B0_3_ran_l,B1_3_ran_l,sum_0_ran_r,carry_0_ran_r,out_2_ran_r,A_less_B_3_ran_r,A_greater_B_3_ran_r);
input a_0_ran_l,b_0_ran_l,A0_3_ran_l,A1_3_ran_l,B0_3_ran_l,B1_3_ran_l;
output sum_0_ran_r,carry_0_ran_r,out_2_ran_r,A_less_B_3_ran_r,A_greater_B_3_ran_r;
wire sum_0_ran_l,carry_0_ran_l,A_less_B_3_ran_l,A_greater_B_3_ran_l,n34_3_ran_l,n35_3_ran_l,n36_3_ran_l,n37_3_ran_l,n38_3_ran_l,n39_3_ran_l,n40_3_ran_l,n41_3_ran_l,n44_3_ran_l,s0bar_2_ran_r,s1bar_2_ran_r,T1_2_ran_r,T2_2_ran_r,T3_2_ran_r,T4_2_ran_r,n34_3_ran_r,n35_3_ran_r,n36_3_ran_r,n37_3_ran_r,n38_3_ran_r,n39_3_ran_r,n40_3_ran_r,n41_3_ran_r,n44_3_ran_r;
xor I_0(sum_0_ran_l,a_0_ran_l,b_0_ran_l);
and I_1(carry_0_ran_l,a_0_ran_l,b_0_ran_l);
nand I_2(A_less_B_3_ran_l,n34_3_ran_l,n35_3_ran_l);
nand I_3(A_greater_B_3_ran_l,n37_3_ran_l,n38_3_ran_l);
nand I_4(n34_3_ran_l,B1_3_ran_l,n40_3_ran_l);
nand I_5(n35_3_ran_l,n36_3_ran_l,n37_3_ran_l);
nor I_6(n36_3_ran_l,A0_3_ran_l,n44_3_ran_l);
or I_7(n37_3_ran_l,B1_3_ran_l,n40_3_ran_l);
nand I_8(n38_3_ran_l,n34_3_ran_l,n39_3_ran_l);
not I_9(n39_3_ran_l,n41_3_ran_l);
not I_10(n40_3_ran_l,A1_3_ran_l);
nand I_11(n41_3_ran_l,A0_3_ran_l,n44_3_ran_l);
not I_12(n44_3_ran_l,B0_3_ran_l);
xor I_13(sum_0_ran_r,sum_0_ran_l,A_less_B_3_ran_l);
and I_14(carry_0_ran_r,sum_0_ran_l,A_less_B_3_ran_l);
or I_15(out_2_ran_r,T1_2_ran_r,T2_2_ran_r,T3_2_ran_r,T4_2_ran_r);
not I_16(s0bar_2_ran_r,A_greater_B_3_ran_l);
not I_17(s1bar_2_ran_r,carry_0_ran_l);
and I_18(T1_2_ran_r,s0bar_2_ran_r,s1bar_2_ran_r,A_less_B_3_ran_l);
and I_19(T2_2_ran_r,s0bar_2_ran_r,carry_0_ran_l,sum_0_ran_l);
and I_20(T3_2_ran_r,s1bar_2_ran_r,A_greater_B_3_ran_l,sum_0_ran_l);
and I_21(T4_2_ran_r,carry_0_ran_l,A_less_B_3_ran_l,A_greater_B_3_ran_l);
nand I_22(A_less_B_3_ran_r,n34_3_ran_r,n35_3_ran_r);
nand I_23(A_greater_B_3_ran_r,n37_3_ran_r,n38_3_ran_r);
nand I_24(n34_3_ran_r,n40_3_ran_r,A_greater_B_3_ran_l);
nand I_25(n35_3_ran_r,n36_3_ran_r,n37_3_ran_r);
nor I_26(n36_3_ran_r,n44_3_ran_r,sum_0_ran_l);
or I_27(n37_3_ran_r,n40_3_ran_r,A_greater_B_3_ran_l);
nand I_28(n38_3_ran_r,n34_3_ran_r,n39_3_ran_r);
not I_29(n39_3_ran_r,n41_3_ran_r);
not I_30(n40_3_ran_r,carry_0_ran_l);
nand I_31(n41_3_ran_r,n44_3_ran_r,sum_0_ran_l);
not I_32(n44_3_ran_r,A_greater_B_3_ran_l);
endmodule


