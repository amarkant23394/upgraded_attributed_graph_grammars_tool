module test_I9131(I6992,I1477,I7365,I7057,I1470,I9015,I6890,I6887,I9131);
input I6992,I1477,I7365,I7057,I1470,I9015,I6890,I6887;
output I9131;
wire I9066,I9032,I9049,I9114,I8862,I6881,I8879,I6907,I9083,I6869;
nor I_0(I9131,I9066,I9114);
DFFARX1 I_1(I9049,I1470,I8862,,,I9066,);
and I_2(I9032,I9015,I6890);
or I_3(I9049,I9032,I6869);
not I_4(I9114,I9083);
not I_5(I8862,I1477);
nand I_6(I6881,I6992,I7057);
not I_7(I8879,I6887);
not I_8(I6907,I1477);
nand I_9(I9083,I8879,I6881);
DFFARX1 I_10(I7365,I1470,I6907,,,I6869,);
endmodule


