module test_I10023(I8107,I1477,I8028,I1470,I10023);
input I8107,I1477,I8028,I1470;
output I10023;
wire I7570,I10137,I7553,I10052,I8124;
not I_0(I7570,I1477);
DFFARX1 I_1(I10137,I1470,I10052,,,I10023,);
DFFARX1 I_2(I7553,I1470,I10052,,,I10137,);
DFFARX1 I_3(I8124,I1470,I7570,,,I7553,);
not I_4(I10052,I1477);
or I_5(I8124,I8107,I8028);
endmodule


