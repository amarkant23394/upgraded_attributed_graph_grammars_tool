module test_final(IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_2,n_572_1_r_2,n_573_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2,N3_2_l_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_2,blif_clk_net_1_r_15,n4_15,G42_1_r_2,);
nor I_1(n_572_1_r_2,n26_2,n18_2);
nand I_2(n_573_1_r_2,n17_2,n19_2);
nor I_3(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_4(n_569_1_r_2,n13_2,n19_2);
not I_5(n_452_1_r_2,n_573_1_r_2);
nor I_6(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_7(N3_2_r_2,blif_clk_net_1_r_15,n4_15,G199_2_r_2,);
DFFARX1 I_8(ACVQN2_3_l_2,blif_clk_net_1_r_15,n4_15,ACVQN1_5_r_2,);
not I_9(P6_5_r_2,P6_5_r_internal_2);
and I_10(N3_2_l_2,IN_6_2_l_2,n24_2);
DFFARX1 I_11(N3_2_l_2,blif_clk_net_1_r_15,n4_15,G199_2_l_2,);
not I_12(n13_2,G199_2_l_2);
DFFARX1 I_13(IN_1_3_l_2,blif_clk_net_1_r_15,n4_15,ACVQN2_3_l_2,);
DFFARX1 I_14(IN_2_3_l_2,blif_clk_net_1_r_15,n4_15,n16_2,);
and I_15(N1_4_l_2,IN_6_4_l_2,n25_2);
DFFARX1 I_16(N1_4_l_2,blif_clk_net_1_r_15,n4_15,n26_2,);
DFFARX1 I_17(IN_3_4_l_2,blif_clk_net_1_r_15,n4_15,n17_internal_2,);
not I_18(n17_2,n17_internal_2);
nor I_19(n4_1_r_2,n26_2,n22_2);
nor I_20(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_21(G199_2_l_2,blif_clk_net_1_r_15,n4_15,P6_5_r_internal_2,);
nor I_22(n18_2,IN_1_2_l_2,IN_3_2_l_2);
nand I_23(n19_2,IN_4_3_l_2,n16_2);
nor I_24(n20_2,n26_2,n21_2);
not I_25(n21_2,n18_2);
and I_26(n22_2,IN_4_3_l_2,n16_2);
nor I_27(n23_2,n13_2,n21_2);
nand I_28(n24_2,IN_2_2_l_2,IN_3_2_l_2);
nand I_29(n25_2,IN_1_4_l_2,IN_2_4_l_2);
DFFARX1 I_30(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_31(n_572_1_r_15,n17_15,n19_15);
nand I_32(n_573_1_r_15,n15_15,n18_15);
nor I_33(n_549_1_r_15,n21_15,n22_15);
nand I_34(n_569_1_r_15,n15_15,n20_15);
nor I_35(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_36(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_37(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_38(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_39(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_40(n4_1_l_15,ACVQN1_5_r_2,n_572_1_r_2);
not I_41(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_42(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_43(n15_15,G42_1_l_15);
DFFARX1 I_44(G42_1_r_2,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_45(n17_15,n17_internal_15);
DFFARX1 I_46(n_452_1_r_2,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_47(n_572_1_l_15,n_42_2_r_2,G199_2_r_2);
DFFARX1 I_48(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_49(n14_15,n14_internal_15);
nand I_50(N1_4_r_15,n25_15,n26_15);
or I_51(n_573_1_l_15,G42_1_r_2,n_549_1_r_2);
nor I_52(n18_15,G42_1_r_2,n_569_1_r_2);
nand I_53(n19_15,n27_15,n28_15);
nand I_54(n20_15,n30_15,n_572_1_r_2);
not I_55(n21_15,n20_15);
and I_56(n22_15,n17_15,n_572_1_l_15);
nor I_57(n23_15,n_549_1_r_2,n_572_1_r_2);
or I_58(n24_15,G42_1_r_2,n_569_1_r_2);
or I_59(n25_15,n_573_1_l_15,n_572_1_r_2);
nand I_60(n26_15,n19_15,n23_15);
not I_61(n27_15,n_569_1_r_2);
nand I_62(n28_15,n29_15,P6_5_r_2);
not I_63(n29_15,n_42_2_r_2);
endmodule


