module test_I13491(I11378,I8836,I1477,I11525,I8833,I8851,I1470,I13491);
input I11378,I8836,I1477,I11525,I8833,I8851,I1470;
output I13491;
wire I11672,I11559,I11296,I11542,I13197,I11689,I11395,I11310;
DFFARX1 I_0(I8836,I1470,I11310,,,I11672,);
DFFARX1 I_1(I11542,I1470,I11310,,,I11559,);
nand I_2(I11296,I11559,I11689);
or I_3(I11542,I11525,I8833);
not I_4(I13197,I1477);
nor I_5(I11689,I11672,I11395);
nand I_6(I11395,I11378,I8851);
DFFARX1 I_7(I11296,I1470,I13197,,,I13491,);
not I_8(I11310,I1477);
endmodule


