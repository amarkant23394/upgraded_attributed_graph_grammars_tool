module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_11,blif_reset_net_1_r_11,G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_11,blif_reset_net_1_r_11;
output G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_431_0_l_11,n9_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_11,n9_11,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_11,n9_11,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_11,n9_11,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_11,n9_11,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_11,n9_11,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_11,n9_11,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_11,n9_11,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_11,blif_clk_net_1_r_11,n9_11,G42_1_r_11,);
nor I_32(n_572_1_r_11,n29_11,n30_11);
nand I_33(n_573_1_r_11,n26_11,n28_11);
nor I_34(n_549_1_r_11,n27_11,n32_11);
nand I_35(n_569_1_r_11,n45_11,n28_11);
nor I_36(n_452_1_r_11,n43_11,n44_11);
nor I_37(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_38(N3_2_r_11,blif_clk_net_1_r_11,n9_11,G199_2_r_11,);
DFFARX1 I_39(n24_11,blif_clk_net_1_r_11,n9_11,ACVQN2_3_r_11,);
nor I_40(n_266_and_0_3_r_11,n20_11,n37_11);
or I_41(n_431_0_l_11,n33_11,n_42_2_r_14);
not I_42(n9_11,blif_reset_net_1_r_11);
DFFARX1 I_43(n_431_0_l_11,blif_clk_net_1_r_11,n9_11,n43_11,);
not I_44(n26_11,n43_11);
DFFARX1 I_45(G199_2_r_14,blif_clk_net_1_r_11,n9_11,n44_11,);
DFFARX1 I_46(P6_5_r_14,blif_clk_net_1_r_11,n9_11,n45_11,);
not I_47(n27_11,n45_11);
nor I_48(n4_1_r_11,n44_11,n25_11);
nor I_49(N3_2_r_11,n45_11,n40_11);
nand I_50(n24_11,n39_11,ACVQN1_5_r_14);
nand I_51(n25_11,n38_11,n_572_1_r_14);
DFFARX1 I_52(n25_11,blif_clk_net_1_r_11,n9_11,n20_internal_11,);
not I_53(n20_11,n20_internal_11);
not I_54(n28_11,n25_11);
not I_55(n29_11,n_569_1_r_14);
nand I_56(n30_11,n26_11,n31_11);
not I_57(n31_11,n_572_1_r_14);
and I_58(n32_11,n26_11,n44_11);
and I_59(n33_11,n34_11,n_573_1_r_14);
nor I_60(n34_11,n29_11,G42_1_r_14);
not I_61(n35_11,n_549_1_r_14);
nand I_62(n36_11,n31_11,n_569_1_r_14);
nor I_63(n37_11,n29_11,n_572_1_r_14);
nor I_64(n38_11,n31_11,n_549_1_r_14);
nor I_65(n39_11,G42_1_r_14,n_549_1_r_14);
nor I_66(n40_11,n41_11,n_549_1_r_14);
nor I_67(n41_11,n42_11,G42_1_r_14);
not I_68(n42_11,ACVQN1_5_r_14);
endmodule


