module test_I6110(I4629,I4979,I1477,I1470,I6110);
input I4629,I4979,I1477,I1470;
output I6110;
wire I4996,I2143,I5751,I4544,I5013,I4807,I4824,I4509;
and I_0(I4996,I4629,I4979);
DFFARX1 I_1(I1470,,,I2143,);
not I_2(I5751,I1477);
DFFARX1 I_3(I4509,I1470,I5751,,,I6110,);
not I_4(I4544,I1477);
or I_5(I5013,I4824,I4996);
DFFARX1 I_6(I1470,I4544,,,I4807,);
and I_7(I4824,I4807,I2143);
DFFARX1 I_8(I5013,I1470,I4544,,,I4509,);
endmodule


