module test_I6881(I5351,I5073,I5625,I5481,I5249,I5204,I6881);
input I5351,I5073,I5625,I5481,I5249,I5204;
output I6881;
wire I6992,I6975,I5368,I5070,I7026,I7057,I5097,I5642,I6924;
nand I_0(I6992,I6975,I5097);
nor I_1(I6975,I6924,I5070);
nor I_2(I5368,I5351,I5204);
and I_3(I5070,I5249,I5481);
not I_4(I7026,I5070);
not I_5(I7057,I7026);
nand I_6(I6881,I6992,I7057);
nand I_7(I5097,I5642,I5368);
not I_8(I5642,I5625);
not I_9(I6924,I5073);
endmodule


