module test_I16780(I1477,I16835,I1470,I17030,I14957,I16780);
input I1477,I16835,I1470,I17030,I14957;
output I16780;
wire I14933,I17157,I17174,I17047,I16869,I17092,I16818,I16852,I17109;
DFFARX1 I_0(I1470,,,I14933,);
nand I_1(I17157,I17109,I17047);
DFFARX1 I_2(I17174,I1470,I16818,,,I16780,);
and I_3(I17174,I16869,I17157);
DFFARX1 I_4(I17030,I1470,I16818,,,I17047,);
DFFARX1 I_5(I16852,I1470,I16818,,,I16869,);
DFFARX1 I_6(I1470,I16818,,,I17092,);
not I_7(I16818,I1477);
and I_8(I16852,I16835,I14957);
and I_9(I17109,I17092,I14933);
endmodule


