module test_I14455(I1477,I1470,I11624,I14455);
input I1477,I1470,I11624;
output I14455;
wire I13177,I13491,I13542,I13426,I11272,I11302,I11278,I13508,I11864,I13296,I13460,I11310,I14370;
nand I_0(I13177,I13296,I13542);
DFFARX1 I_1(I1470,,,I13491,);
nor I_2(I13542,I13508,I13460);
DFFARX1 I_3(I1470,,,I13426,);
DFFARX1 I_4(I1470,I11310,,,I11272,);
DFFARX1 I_5(I13177,I1470,I14370,,,I14455,);
DFFARX1 I_6(I11864,I1470,I11310,,,I11302,);
DFFARX1 I_7(I11624,I1470,I11310,,,I11278,);
and I_8(I13508,I13491,I11272);
and I_9(I11864,I11624);
nor I_10(I13296,I11278,I11302);
not I_11(I13460,I13426);
not I_12(I11310,I1477);
not I_13(I14370,I1477);
endmodule


