module test_I3293(I1431,I1477,I1470,I3293);
input I1431,I1477,I1470;
output I3293;
wire I3217,I2759,I3200;
not I_0(I3217,I3200);
not I_1(I3293,I3217);
not I_2(I2759,I1477);
DFFARX1 I_3(I1431,I1470,I2759,,,I3200,);
endmodule


