module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_7,n8_7,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_7,n8_7,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_7,n8_7,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_7,n8_7,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_7,n8_7,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_7,n8_7,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_7,n8_7,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_7,n8_7,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_32(n_572_1_r_7,n30_7,n31_7);
nand I_33(n_573_1_r_7,n28_7,G199_4_r_6);
nor I_34(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_35(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_36(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_37(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_38(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_39(P6_5_r_7,P6_5_r_internal_7);
or I_40(n_431_0_l_7,n36_7,n_549_1_r_6);
not I_41(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_42(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_43(n27_7,n43_7);
DFFARX1 I_44(ACVQN1_5_r_6,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_45(G42_1_r_6,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_46(n4_1_r_7,n30_7,n38_7);
nor I_47(N1_4_r_7,n27_7,n40_7);
nand I_48(n26_7,n39_7,P6_5_r_6);
not I_49(n5_7,n_572_1_r_6);
DFFARX1 I_50(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_51(n28_7,n26_7,n29_7);
not I_52(n29_7,G214_4_r_6);
not I_53(n30_7,n_452_1_r_6);
nand I_54(n31_7,n27_7,n29_7);
nor I_55(n32_7,ACVQN1_5_l_7,n34_7);
nor I_56(n33_7,n29_7,n_572_1_r_6);
not I_57(n34_7,G199_4_r_6);
nor I_58(n35_7,n43_7,n44_7);
and I_59(n36_7,n37_7,G42_1_r_6);
nor I_60(n37_7,n30_7,n_569_1_r_6);
nand I_61(n38_7,n29_7,n_572_1_r_6);
nor I_62(n39_7,n_572_1_r_6,n_573_1_r_6);
nor I_63(n40_7,n44_7,n41_7);
nor I_64(n41_7,n34_7,n42_7);
nand I_65(n42_7,n5_7,G214_4_r_6);
endmodule


