module test_I10332(I6309,I1477,I1470,I10332);
input I6309,I1477,I1470;
output I10332;
wire I8107,I8090,I7570,I10052,I7532;
not I_0(I8107,I8090);
DFFARX1 I_1(I6309,I1470,I7570,,,I8090,);
not I_2(I7570,I1477);
not I_3(I10052,I1477);
DFFARX1 I_4(I8107,I1470,I7570,,,I7532,);
DFFARX1 I_5(I7532,I1470,I10052,,,I10332,);
endmodule


