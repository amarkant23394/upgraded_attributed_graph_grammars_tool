module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_5_r_11,n9_11,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
not I_36(N1372_1_r_11,n53_11);
nor I_37(N1508_1_r_11,n39_11,n53_11);
nor I_38(N6147_2_r_11,n48_11,n49_11);
nor I_39(N6147_3_r_11,n44_11,n45_11);
nand I_40(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_41(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_42(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_43(n_102_5_r_11,n39_11);
nand I_44(n_547_5_r_11,n36_11,n37_11);
nor I_45(N1507_6_r_11,n52_11,n57_11);
nor I_46(N1508_6_r_11,n46_11,n51_11);
nor I_47(N1372_10_r_11,n43_11,n47_11);
nor I_48(N1508_10_r_11,n55_11,n56_11);
nand I_49(n_431_5_r_11,n40_11,n41_11);
not I_50(n9_11,blif_reset_net_5_r_11);
nor I_51(n36_11,n38_11,n39_11);
not I_52(n37_11,n40_11);
nor I_53(n38_11,n60_11,N1508_1_r_3);
nor I_54(n39_11,n54_11,N1508_6_r_3);
nand I_55(n40_11,N1507_6_r_3,n_549_7_r_3);
nand I_56(n41_11,n_102_5_r_11,n42_11);
and I_57(n42_11,n58_11,N1372_1_r_3);
not I_58(n43_11,n44_11);
nor I_59(n44_11,n40_11,N1372_1_r_3);
nand I_60(n45_11,n46_11,n47_11);
not I_61(n46_11,n38_11);
nand I_62(n47_11,n59_11,n62_11);
and I_63(n48_11,n37_11,n47_11);
or I_64(n49_11,n44_11,n50_11);
nor I_65(n50_11,n60_11,n61_11);
or I_66(n51_11,n_102_5_r_11,n52_11);
nor I_67(n52_11,n42_11,n57_11);
nand I_68(n53_11,n37_11,n50_11);
or I_69(n54_11,G42_7_r_3,n_452_7_r_3);
nor I_70(n55_11,n38_11,n42_11);
not I_71(n56_11,N1372_10_r_11);
and I_72(n57_11,n38_11,n50_11);
and I_73(n58_11,n59_11,N1508_6_r_3);
or I_74(n59_11,n63_11,n_573_7_r_3);
not I_75(n60_11,n_569_7_r_3);
nor I_76(n61_11,N1507_6_r_3,G42_7_r_3);
nand I_77(n62_11,N1508_1_r_3,N6134_9_r_3);
and I_78(n63_11,N1508_1_r_3,N6134_9_r_3);
endmodule


