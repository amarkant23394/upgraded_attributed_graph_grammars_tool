module test_I7816(I6722,I1477,I1470,I7748,I7816);
input I6722,I1477,I1470,I7748;
output I7816;
wire I7799,I7570,I7765,I6329,I6380,I7782,I6312,I6411,I6303,I6306;
or I_0(I7799,I7782,I6306);
DFFARX1 I_1(I7799,I1470,I7570,,,I7816,);
not I_2(I7570,I1477);
nor I_3(I7765,I7748,I6303);
not I_4(I6329,I1477);
DFFARX1 I_5(I1470,I6329,,,I6380,);
and I_6(I7782,I7765,I6312);
DFFARX1 I_7(I6722,I1470,I6329,,,I6312,);
DFFARX1 I_8(I6380,I1470,I6329,,,I6411,);
DFFARX1 I_9(I1470,I6329,,,I6303,);
not I_10(I6306,I6411);
endmodule


