module test_I2545(I1902,I1294,I1301,I2545);
input I1902,I1294,I1301;
output I2545;
wire I2583,I3024,I2039,I3041,I1908,I2634,I2617,I1929,I2945,I2702;
not I_0(I2583,I1301);
nand I_1(I3024,I2945,I2634);
DFFARX1 I_2(I1294,,,I2039,);
and I_3(I3041,I2702,I3024);
not I_4(I1908,I2039);
DFFARX1 I_5(I3041,I1294,I2583,,,I2545,);
nand I_6(I2634,I2617,I1929);
nor I_7(I2617,I1908);
DFFARX1 I_8(I1294,,,I1929,);
DFFARX1 I_9(I1902,I1294,I2583,,,I2945,);
not I_10(I2702,I1908);
endmodule


