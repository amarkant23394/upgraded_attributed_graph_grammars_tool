module test_I7765(I1477,I1470,I4130,I3972,I7765);
input I1477,I1470,I4130,I3972;
output I7765;
wire I6781,I3957,I6329,I6688,I4308,I6705,I6291,I6303,I7748;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
nand I_1(I3957,I4308,I4130);
nor I_2(I7765,I7748,I6303);
not I_3(I6329,I1477);
DFFARX1 I_4(I1470,I6329,,,I6688,);
DFFARX1 I_5(I1470,,,I4308,);
and I_6(I6705,I6688,I3972);
DFFARX1 I_7(I6705,I1470,I6329,,,I6291,);
DFFARX1 I_8(I6781,I1470,I6329,,,I6303,);
not I_9(I7748,I6291);
endmodule


