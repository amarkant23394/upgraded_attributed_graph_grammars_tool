module test_I12596(I12687,I1477,I10961,I1470,I10636,I12596);
input I12687,I1477,I10961,I1470,I10636;
output I12596;
wire I12619,I10647,I13023,I12718,I10615,I12865,I13119,I13102,I10639,I11201,I12848;
not I_0(I12619,I1477);
not I_1(I10647,I1477);
DFFARX1 I_2(I10636,I1470,I12619,,,I13023,);
nor I_3(I12718,I10615,I10639);
DFFARX1 I_4(I10961,I1470,I10647,,,I10615,);
nor I_5(I12865,I12848,I12687);
DFFARX1 I_6(I13119,I1470,I12619,,,I12596,);
or I_7(I13119,I12718,I13102);
and I_8(I13102,I13023,I12865);
DFFARX1 I_9(I11201,I1470,I10647,,,I10639,);
and I_10(I11201,I10961);
DFFARX1 I_11(I1470,I12619,,,I12848,);
endmodule


