module test_I3983(I1477,I3983);
input I1477;
output I3983;
wire ;
not I_0(I3983,I1477);
endmodule


