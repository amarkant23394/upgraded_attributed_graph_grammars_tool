module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_5_r_11,n9_11,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_5_r_11,n9_11,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_5_r_11,n9_11,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_5_r_11,n9_11,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
not I_43(N1372_1_r_11,n53_11);
nor I_44(N1508_1_r_11,n39_11,n53_11);
nor I_45(N6147_2_r_11,n48_11,n49_11);
nor I_46(N6147_3_r_11,n44_11,n45_11);
nand I_47(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_48(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_49(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_50(n_102_5_r_11,n39_11);
nand I_51(n_547_5_r_11,n36_11,n37_11);
nor I_52(N1507_6_r_11,n52_11,n57_11);
nor I_53(N1508_6_r_11,n46_11,n51_11);
nor I_54(N1372_10_r_11,n43_11,n47_11);
nor I_55(N1508_10_r_11,n55_11,n56_11);
nand I_56(n_431_5_r_11,n40_11,n41_11);
not I_57(n9_11,blif_reset_net_5_r_11);
nor I_58(n36_11,n38_11,n39_11);
not I_59(n37_11,n40_11);
nor I_60(n38_11,n60_11,N6147_2_r_9);
nor I_61(n39_11,n54_11,G78_5_r_9);
nand I_62(n40_11,n_547_5_r_9,N1372_4_r_9);
nand I_63(n41_11,n_102_5_r_11,n42_11);
and I_64(n42_11,n58_11,N1508_4_r_9);
not I_65(n43_11,n44_11);
nor I_66(n44_11,n40_11,G78_5_r_9);
nand I_67(n45_11,n46_11,n47_11);
not I_68(n46_11,n38_11);
nand I_69(n47_11,n59_11,n62_11);
and I_70(n48_11,n37_11,n47_11);
or I_71(n49_11,n44_11,n50_11);
nor I_72(n50_11,n60_11,n61_11);
or I_73(n51_11,n_102_5_r_11,n52_11);
nor I_74(n52_11,n42_11,n57_11);
nand I_75(n53_11,n37_11,n50_11);
or I_76(n54_11,N6147_2_r_9,N1372_4_r_9);
nor I_77(n55_11,n38_11,n42_11);
not I_78(n56_11,N1372_10_r_11);
and I_79(n57_11,n38_11,n50_11);
and I_80(n58_11,n59_11,n_42_8_r_9);
or I_81(n59_11,n63_11,N6147_9_r_9);
not I_82(n60_11,n_576_5_r_9);
nor I_83(n61_11,N1508_4_r_9,N6134_9_r_9);
nand I_84(n62_11,G199_8_r_9,n_576_5_r_9);
and I_85(n63_11,G199_8_r_9,n_576_5_r_9);
endmodule


