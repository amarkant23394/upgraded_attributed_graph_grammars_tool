module test_I5737(I4629,I1477,I4524,I1470,I5737);
input I4629,I1477,I4524,I1470;
output I5737;
wire I4544,I4869,I2149,I5785,I5898,I5802,I4518,I4536,I5881,I5768,I6203,I5751,I4674,I5864,I4515,I4691;
not I_0(I4544,I1477);
DFFARX1 I_1(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_2(I1470,,,I2149,);
and I_3(I5785,I5768,I4524);
nor I_4(I5898,I5802,I5881);
DFFARX1 I_5(I5785,I1470,I5751,,,I5802,);
nand I_6(I4518,I4869,I4691);
nor I_7(I4536,I4869);
not I_8(I5881,I5864);
nand I_9(I5768,I4515);
nand I_10(I5737,I6203,I5898);
DFFARX1 I_11(I4518,I1470,I5751,,,I6203,);
not I_12(I5751,I1477);
DFFARX1 I_13(I1470,I4544,,,I4674,);
nor I_14(I5864,I4536,I4515);
not I_15(I4515,I4629);
nor I_16(I4691,I4674,I4629);
endmodule


