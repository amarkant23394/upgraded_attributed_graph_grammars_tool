module test_I6321(I2733,I1477,I6572,I2742,I6346,I3963,I1470,I6321);
input I2733,I1477,I6572,I2742,I6346,I3963,I1470;
output I6321;
wire I6380,I6705,I3972,I3983,I6329,I6363,I4068,I4263,I2724,I6657,I6688,I4452,I6606,I3960,I6589,I3948,I4246;
DFFARX1 I_0(I6363,I1470,I6329,,,I6380,);
and I_1(I6705,I6688,I3972);
or I_2(I3972,I4263,I4068);
not I_3(I3983,I1477);
not I_4(I6329,I1477);
and I_5(I6363,I6346,I3963);
nor I_6(I4068,I2742,I2724);
and I_7(I4263,I4246,I2733);
DFFARX1 I_8(I1470,,,I2724,);
nor I_9(I6657,I6606,I6380);
nand I_10(I6321,I6705,I6657);
DFFARX1 I_11(I3948,I1470,I6329,,,I6688,);
or I_12(I4452,I4263);
DFFARX1 I_13(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_14(I1470,I3983,,,I3960,);
and I_15(I6589,I6572,I3960);
DFFARX1 I_16(I4452,I1470,I3983,,,I3948,);
DFFARX1 I_17(I1470,I3983,,,I4246,);
endmodule


