module test_final(IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_8_l_1,IN_2_8_l_1,IN_3_8_l_1,IN_6_8_l_1,IN_1_10_l_1,IN_2_10_l_1,IN_3_10_l_1,IN_4_10_l_1,blif_clk_net_5_r_5,blif_reset_net_5_r_5,N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5);
input IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_8_l_1,IN_2_8_l_1,IN_3_8_l_1,IN_6_8_l_1,IN_1_10_l_1,IN_2_10_l_1,IN_3_10_l_1,IN_4_10_l_1,blif_clk_net_5_r_5,blif_reset_net_5_r_5;
output N1371_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1508_6_r_5;
wire N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,N1372_10_r_1,N1508_10_r_1,N3_8_l_1,n38_1,n22_1,N3_8_r_1,n23_1,n24_1,n25_1,n26_1,n27_1,n28_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,N1508_0_r_5,N1507_6_r_5,n_431_5_r_5,n6_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5;
nor I_0(N6147_3_r_1,n26_1,n27_1);
not I_1(N1372_4_r_1,n34_1);
nor I_2(N1508_4_r_1,n30_1,n34_1);
nor I_3(n_42_8_r_1,n23_1,n24_1);
DFFARX1 I_4(N3_8_r_1,blif_clk_net_5_r_5,n6_5,G199_8_r_1,);
nor I_5(N6147_9_r_1,n22_1,n25_1);
nor I_6(N6134_9_r_1,n29_1,n30_1);
not I_7(I_BUFF_1_9_r_1,n32_1);
not I_8(N1372_10_r_1,n36_1);
nor I_9(N1508_10_r_1,n35_1,n36_1);
and I_10(N3_8_l_1,IN_6_8_l_1,n33_1);
DFFARX1 I_11(N3_8_l_1,blif_clk_net_5_r_5,n6_5,n38_1,);
not I_12(n22_1,n38_1);
nor I_13(N3_8_r_1,n31_1,n32_1);
nor I_14(n23_1,IN_3_1_l_1,n28_1);
nor I_15(n24_1,IN_1_8_l_1,IN_3_8_l_1);
nor I_16(n25_1,n23_1,n26_1);
not I_17(n26_1,n30_1);
nand I_18(n27_1,n22_1,n28_1);
nand I_19(n28_1,IN_1_1_l_1,IN_2_1_l_1);
not I_20(n29_1,n28_1);
nand I_21(n30_1,IN_1_10_l_1,IN_2_10_l_1);
and I_22(n31_1,n38_1,n24_1);
nand I_23(n32_1,n26_1,n37_1);
nand I_24(n33_1,IN_2_8_l_1,IN_3_8_l_1);
nand I_25(n34_1,n24_1,n29_1);
nor I_26(n35_1,n38_1,n24_1);
nand I_27(n36_1,I_BUFF_1_9_r_1,n23_1);
or I_28(n37_1,IN_3_10_l_1,IN_4_10_l_1);
nor I_29(N1371_0_r_5,n28_5,n39_5);
not I_30(N1508_0_r_5,n39_5);
nor I_31(N6147_2_r_5,n28_5,n37_5);
nand I_32(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_33(n_431_5_r_5,blif_clk_net_5_r_5,n6_5,G78_5_r_5,);
nand I_34(n_576_5_r_5,n26_5,n27_5);
not I_35(n_102_5_r_5,n28_5);
nand I_36(n_547_5_r_5,n31_5,n32_5);
nor I_37(N1507_6_r_5,n30_5,n32_5);
nor I_38(N1508_6_r_5,n39_5,n41_5);
nand I_39(n_431_5_r_5,n34_5,n35_5);
not I_40(n6_5,blif_reset_net_5_r_5);
nor I_41(n26_5,n29_5,n30_5);
nor I_42(n27_5,n28_5,N6147_3_r_1);
nor I_43(n28_5,n29_5,n44_5);
not I_44(n29_5,N1372_4_r_1);
nand I_45(n30_5,N1508_0_r_5,n43_5);
nor I_46(n31_5,n28_5,n33_5);
nor I_47(n32_5,n40_5,N1372_10_r_1);
nor I_48(n33_5,n29_5,N6147_3_r_1);
or I_49(n34_5,n29_5,N6147_3_r_1);
nand I_50(n35_5,n32_5,n36_5);
not I_51(n36_5,n30_5);
nor I_52(n37_5,N1507_6_r_5,n38_5);
and I_53(n38_5,n39_5,n40_5);
nand I_54(n39_5,N1508_4_r_1,N1508_10_r_1);
nand I_55(n40_5,G199_8_r_1,N1372_4_r_1);
nand I_56(n41_5,n28_5,n42_5);
or I_57(n42_5,n32_5,n36_5);
or I_58(n43_5,n_42_8_r_1,N6147_9_r_1);
nor I_59(n44_5,N6147_3_r_1,N6134_9_r_1);
endmodule


