module test_I17950(I1477,I13749,I15579,I16162,I16069,I15628,I1470,I15798,I17950);
input I1477,I13749,I15579,I16162,I16069,I15628,I1470,I15798;
output I17950;
wire I17413,I15600,I15832,I15815,I15611,I17498,I15928,I15597,I17916,I17430,I15603,I17933,I17481;
not I_0(I17413,I1477);
or I_1(I15600,I15832,I15815);
nand I_2(I15832,I15628,I13749);
DFFARX1 I_3(I15798,I1470,I15611,,,I15815,);
not I_4(I15611,I1477);
nand I_5(I17498,I17481,I15600);
DFFARX1 I_6(I1470,I15611,,,I15928,);
nor I_7(I15597,I15832,I16162);
DFFARX1 I_8(I15603,I1470,I17413,,,I17916,);
not I_9(I17430,I15579);
nand I_10(I17950,I17933,I17498);
nor I_11(I15603,I15928,I16069);
not I_12(I17933,I17916);
nor I_13(I17481,I17430,I15597);
endmodule


