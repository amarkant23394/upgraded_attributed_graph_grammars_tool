module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_7_r_1,n9_1,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
and I_36(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_37(N1508_0_r_1,n40_1,n44_1);
nor I_38(N1507_6_r_1,n43_1,n49_1);
nor I_39(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_40(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_41(n_572_7_r_1,n29_1,n30_1);
not I_42(n_573_7_r_1,n_452_7_r_1);
nor I_43(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_44(n_569_7_r_1,n30_1,n31_1);
nor I_45(n_452_7_r_1,n30_1,n32_1);
nor I_46(N6147_9_r_1,n35_1,n36_1);
nand I_47(N6134_9_r_1,n38_1,n39_1);
not I_48(I_BUFF_1_9_r_1,n40_1);
nor I_49(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_50(n9_1,blif_reset_net_7_r_1);
nor I_51(n29_1,n34_1,N1508_6_r_3);
nor I_52(n30_1,n33_1,n34_1);
nor I_53(n31_1,n54_1,N1508_1_r_3);
not I_54(n32_1,n48_1);
nor I_55(n33_1,N1508_1_r_3,n_569_7_r_3);
not I_56(n34_1,N1372_1_r_3);
nor I_57(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_58(n36_1,n29_1);
not I_59(n37_1,n41_1);
nand I_60(n38_1,I_BUFF_1_9_r_1,N6134_9_r_3);
nand I_61(n39_1,n37_1,n40_1);
nand I_62(n40_1,N1507_6_r_3,G42_7_r_3);
nand I_63(n41_1,n52_1,n_452_7_r_3);
or I_64(n42_1,n36_1,n43_1);
nor I_65(n43_1,n32_1,n49_1);
nand I_66(n44_1,n45_1,n46_1);
nand I_67(n45_1,n47_1,n48_1);
not I_68(n46_1,N6134_9_r_3);
not I_69(n47_1,n31_1);
nand I_70(n48_1,n50_1,N1508_6_r_3);
nor I_71(n49_1,n41_1,n47_1);
and I_72(n50_1,n51_1,n_573_7_r_3);
nand I_73(n51_1,n52_1,n53_1);
nand I_74(n52_1,G42_7_r_3,N1507_6_r_3);
not I_75(n53_1,n_452_7_r_3);
or I_76(n54_1,n_549_7_r_3,N1372_1_r_3);
nor I_77(n55_1,n29_1,N6134_9_r_3);
endmodule


