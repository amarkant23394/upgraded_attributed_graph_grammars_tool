module test_I8753(I5864,I1477,I4527,I1470,I8753);
input I5864,I1477,I4527,I1470;
output I8753;
wire I8216,I5751,I5881,I5915,I5731,I8736;
not I_0(I8216,I1477);
not I_1(I8753,I8736);
not I_2(I5751,I1477);
not I_3(I5881,I5864);
DFFARX1 I_4(I4527,I1470,I5751,,,I5915,);
nand I_5(I5731,I5915,I5881);
DFFARX1 I_6(I5731,I1470,I8216,,,I8736,);
endmodule


