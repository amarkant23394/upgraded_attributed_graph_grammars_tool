module test_I13491(I11378,I8851,I8833,I11525,I8836,I1470_clk,I1477_rst,I13491);
input I11378,I8851,I8833,I11525,I8836,I1470_clk,I1477_rst;
output I13491;
wire I11542,I11689,I11296,I11310_rst,I13197_rst,I11559,I11395,I11672;
or I_0(I11542,I11525,I8833);
nor I_1(I11689,I11672,I11395);
nand I_2(I11296,I11559,I11689);
not I_3(I11310_rst,I1477_rst);
not I_4(I13197_rst,I1477_rst);
DFFARX1 I_5 (I11542,I1470_clk,I11310_rst,I11559);
DFFARX1 I_6 (I11296,I1470_clk,I13197_rst,I13491);
nand I_7(I11395,I11378,I8851);
DFFARX1 I_8 (I8836,I1470_clk,I11310_rst,I11672);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule