module test_I6297(I1477,I1470,I4068,I3957,I6297);
input I1477,I1470,I4068,I3957;
output I6297;
wire I6781,I3966,I3975,I3954,I6826,I6442,I6329,I6493,I6843,I4034;
DFFARX1 I_0(I3957,I1470,I6329,,,I6781,);
DFFARX1 I_1(I6843,I1470,I6329,,,I6297,);
or I_2(I3966,I4068,I4034);
nor I_3(I3975,I4034);
not I_4(I3954,I4068);
nand I_5(I6826,I6781,I6442);
nor I_6(I6442,I3975,I3954);
not I_7(I6329,I1477);
DFFARX1 I_8(I3966,I1470,I6329,,,I6493,);
and I_9(I6843,I6493,I6826);
DFFARX1 I_10(I1470,,,I4034,);
endmodule


