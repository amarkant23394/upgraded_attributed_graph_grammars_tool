module test_I10749(I9576,I9771,I1470,I8193,I9471,I9491,I10749);
input I9576,I9771,I1470,I8193,I9471,I9491;
output I10749;
wire I9477,I10715,I9621,I9465,I9638,I10664,I9816,I9833,I10732;
nor I_0(I9477,I9771,I9833);
nor I_1(I10715,I10664,I9477);
DFFARX1 I_2(I1470,I9491,,,I9621,);
nand I_3(I9465,I9816,I9638);
nor I_4(I9638,I9621,I9576);
not I_5(I10664,I9471);
DFFARX1 I_6(I8193,I1470,I9491,,,I9816,);
not I_7(I10749,I10732);
and I_8(I9833,I9816);
nand I_9(I10732,I10715,I9465);
endmodule


