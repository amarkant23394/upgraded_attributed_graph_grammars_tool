module test_I14942(I12930,I1477,I1470,I14942);
input I12930,I1477,I1470;
output I14942;
wire I12602,I15454,I14965,I15372;
not I_0(I12602,I12930);
not I_1(I14942,I15454);
DFFARX1 I_2(I15372,I1470,I14965,,,I15454,);
not I_3(I14965,I1477);
DFFARX1 I_4(I12602,I1470,I14965,,,I15372,);
endmodule


