module test_I14362(I1477,I14520,I1470,I14362);
input I1477,I14520,I1470;
output I14362;
wire I13361,I14667,I13189,I13162,I14537,I14650,I14825,I14808,I13248,I14370,I14684;
DFFARX1 I_0(I1470,,,I13361,);
DFFARX1 I_1(I14825,I1470,I14370,,,I14362,);
and I_2(I14667,I14650,I13189);
DFFARX1 I_3(I1470,,,I13189,);
and I_4(I13162,I13248,I13361);
DFFARX1 I_5(I14520,I1470,I14370,,,I14537,);
DFFARX1 I_6(I1470,I14370,,,I14650,);
and I_7(I14825,I14808,I14684);
DFFARX1 I_8(I13162,I1470,I14370,,,I14808,);
DFFARX1 I_9(I1470,,,I13248,);
not I_10(I14370,I1477);
nand I_11(I14684,I14667,I14537);
endmodule


