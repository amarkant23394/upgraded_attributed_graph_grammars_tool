module test_final(IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_8_r_1,blif_reset_net_8_r_1,N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1);
input IN_1_1_l_4,IN_2_1_l_4,IN_3_1_l_4,IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_3_l_4,IN_2_3_l_4,IN_3_3_l_4,blif_clk_net_8_r_1,blif_reset_net_8_r_1;
output N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1;
wire N1371_0_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_102_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4,n_431_5_r_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,I_BUFF_1_9_r_1,N3_8_l_1,n7_1,n38_1,n22_1,N3_8_r_1,n23_1,n24_1,n25_1,n26_1,n27_1,n28_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1;
nor I_0(N1371_0_r_4,n25_4,n29_4);
nor I_1(N1508_0_r_4,n25_4,n32_4);
nor I_2(N6147_2_r_4,n24_4,n31_4);
or I_3(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_4(n_431_5_r_4,blif_clk_net_8_r_1,n7_1,G78_5_r_4,);
nand I_5(n_576_5_r_4,n22_4,n23_4);
nand I_6(n_102_5_r_4,n34_4,n35_4);
nand I_7(n_547_5_r_4,n26_4,n27_4);
nor I_8(N1507_6_r_4,n27_4,n30_4);
nor I_9(N1508_6_r_4,n30_4,n33_4);
nand I_10(n_431_5_r_4,n_102_5_r_4,n28_4);
nor I_11(n22_4,n24_4,n25_4);
nor I_12(n23_4,IN_1_3_l_4,n37_4);
not I_13(n24_4,n_102_5_r_4);
nand I_14(n25_4,IN_1_1_l_4,IN_2_1_l_4);
nor I_15(n26_4,n23_4,n24_4);
not I_16(n27_4,n25_4);
nand I_17(n28_4,n23_4,n29_4);
nor I_18(n29_4,IN_3_1_l_4,n25_4);
not I_19(n30_4,n29_4);
nor I_20(n31_4,N1371_0_r_4,n32_4);
nor I_21(n32_4,n23_4,n29_4);
nand I_22(n33_4,n23_4,n24_4);
nor I_23(n34_4,IN_1_2_l_4,IN_2_2_l_4);
or I_24(n35_4,IN_5_2_l_4,n36_4);
nor I_25(n36_4,IN_3_2_l_4,IN_4_2_l_4);
or I_26(n37_4,IN_2_3_l_4,IN_3_3_l_4);
nor I_27(N6147_3_r_1,n26_1,n27_1);
not I_28(N1372_4_r_1,n34_1);
nor I_29(N1508_4_r_1,n30_1,n34_1);
nor I_30(n_42_8_r_1,n23_1,n24_1);
DFFARX1 I_31(N3_8_r_1,blif_clk_net_8_r_1,n7_1,G199_8_r_1,);
nor I_32(N6147_9_r_1,n22_1,n25_1);
nor I_33(N6134_9_r_1,n29_1,n30_1);
not I_34(I_BUFF_1_9_r_1,n32_1);
not I_35(N1372_10_r_1,n36_1);
nor I_36(N1508_10_r_1,n35_1,n36_1);
and I_37(N3_8_l_1,n33_1,N1507_6_r_4);
not I_38(n7_1,blif_reset_net_8_r_1);
DFFARX1 I_39(N3_8_l_1,blif_clk_net_8_r_1,n7_1,n38_1,);
not I_40(n22_1,n38_1);
nor I_41(N3_8_r_1,n31_1,n32_1);
nor I_42(n23_1,n28_1,N6147_2_r_4);
nor I_43(n24_1,G78_5_r_4,N1508_6_r_4);
nor I_44(n25_1,n23_1,n26_1);
not I_45(n26_1,n30_1);
nand I_46(n27_1,n22_1,n28_1);
nand I_47(n28_1,N1508_0_r_4,n_429_or_0_5_r_4);
not I_48(n29_1,n28_1);
nand I_49(n30_1,N6147_2_r_4,n_576_5_r_4);
and I_50(n31_1,n38_1,n24_1);
nand I_51(n32_1,n26_1,n37_1);
nand I_52(n33_1,n_429_or_0_5_r_4,G78_5_r_4);
nand I_53(n34_1,n24_1,n29_1);
nor I_54(n35_1,n38_1,n24_1);
nand I_55(n36_1,I_BUFF_1_9_r_1,n23_1);
or I_56(n37_1,N1508_0_r_4,n_547_5_r_4);
endmodule


