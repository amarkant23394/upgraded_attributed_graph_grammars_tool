module test_I7898(I7765,I1477,I1470,I3972,I7898);
input I7765,I1477,I1470,I3972;
output I7898;
wire I6606,I6300,I7799,I7816,I7881,I7570,I7587,I6329,I6688,I7782,I6312,I6705,I6411,I6291,I6306;
DFFARX1 I_0(I1470,I6329,,,I6606,);
nand I_1(I7898,I7881,I7816);
DFFARX1 I_2(I6606,I1470,I6329,,,I6300,);
or I_3(I7799,I7782,I6306);
DFFARX1 I_4(I7799,I1470,I7570,,,I7816,);
nand I_5(I7881,I7587,I6291);
not I_6(I7570,I1477);
not I_7(I7587,I6300);
not I_8(I6329,I1477);
DFFARX1 I_9(I1470,I6329,,,I6688,);
and I_10(I7782,I7765,I6312);
DFFARX1 I_11(I1470,I6329,,,I6312,);
and I_12(I6705,I6688,I3972);
DFFARX1 I_13(I1470,I6329,,,I6411,);
DFFARX1 I_14(I6705,I1470,I6329,,,I6291,);
not I_15(I6306,I6411);
endmodule


