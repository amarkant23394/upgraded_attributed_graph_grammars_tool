module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_5_r_9,n10_9,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N6147_2_r_9,n62_9,n46_9);
not I_37(N1372_4_r_9,n59_9);
nor I_38(N1508_4_r_9,n58_9,n59_9);
nand I_39(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_40(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_41(n_576_5_r_9,n39_9,n40_9);
not I_42(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_43(n_547_5_r_9,n43_9,N1372_1_r_3);
and I_44(n_42_8_r_9,n44_9,N1507_6_r_3);
DFFARX1 I_45(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_46(N6147_9_r_9,n41_9,n45_9);
nor I_47(N6134_9_r_9,n45_9,n51_9);
nor I_48(I_BUFF_1_9_r_9,n41_9,N1372_1_r_3);
nor I_49(n4_7_l_9,N1372_1_r_3,N1507_6_r_3);
not I_50(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_51(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_52(N3_8_l_9,n57_9,n_573_7_r_3);
DFFARX1 I_53(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_54(n38_9,n63_9);
nor I_55(n_431_5_r_9,N1507_6_r_3,n_549_7_r_3);
nor I_56(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_57(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_58(n40_9,n41_9);
nand I_59(n41_9,N1508_1_r_3,G42_7_r_3);
nor I_60(n42_9,N1508_6_r_3,n_452_7_r_3);
nor I_61(n43_9,n63_9,n41_9);
nor I_62(n44_9,n_452_7_r_3,N6134_9_r_3);
and I_63(n45_9,n52_9,N1508_1_r_3);
nor I_64(n46_9,n47_9,n48_9);
nor I_65(n47_9,n49_9,n50_9);
not I_66(n48_9,n_429_or_0_5_r_9);
not I_67(n49_9,n42_9);
or I_68(n50_9,n63_9,n51_9);
nor I_69(n51_9,G42_7_r_3,N1508_6_r_3);
nor I_70(n52_9,n49_9,n_549_7_r_3);
nor I_71(n53_9,n54_9,n55_9);
nor I_72(n54_9,n56_9,n_549_7_r_3);
or I_73(n55_9,n44_9,N1508_6_r_3);
not I_74(n56_9,N1508_1_r_3);
nand I_75(n57_9,G42_7_r_3,n_569_7_r_3);
nor I_76(n58_9,n62_9,n60_9);
nand I_77(n59_9,n51_9,n61_9);
nor I_78(n60_9,n38_9,n44_9);
nor I_79(n61_9,N6134_9_r_3,N1507_6_r_3);
endmodule


