module test_I11962(I1477,I10202,I10414,I7535,I7550,I1470,I11962);
input I1477,I10202,I10414,I7535,I7550,I1470;
output I11962;
wire I10120,I10032,I7538,I10219,I10014,I10041,I10052,I12270,I10349,I12349,I10332,I11990,I10137,I11973;
nor I_0(I10120,I7538,I7535);
nand I_1(I10032,I10137,I10414);
DFFARX1 I_2(I1470,,,I7538,);
DFFARX1 I_3(I10202,I1470,I10052,,,I10219,);
DFFARX1 I_4(I10219,I1470,I10052,,,I10014,);
nor I_5(I10041,I10349,I10120);
not I_6(I10052,I1477);
nand I_7(I12270,I11990,I10014);
and I_8(I10349,I10332,I7550);
DFFARX1 I_9(I10041,I1470,I11973,,,I12349,);
nor I_10(I11962,I12349,I12270);
DFFARX1 I_11(I1470,I10052,,,I10332,);
not I_12(I11990,I10032);
DFFARX1 I_13(I1470,I10052,,,I10137,);
not I_14(I11973,I1477);
endmodule


