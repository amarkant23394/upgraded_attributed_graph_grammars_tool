module test_I16373(I1477,I1470,I16373);
input I1477,I1470;
output I16373;
wire I16356,I14667,I14856,I13189,I16240,I14650,I14356,I14421,I14808;
DFFARX1 I_0(I14356,I1470,I16240,,,I16356,);
and I_1(I14667,I14650,I13189);
nor I_2(I14856,I14808,I14421);
DFFARX1 I_3(I1470,,,I13189,);
not I_4(I16240,I1477);
DFFARX1 I_5(I1470,,,I14650,);
nand I_6(I14356,I14667,I14856);
DFFARX1 I_7(I1470,,,I14421,);
DFFARX1 I_8(I16356,I1470,I16240,,,I16373,);
DFFARX1 I_9(I1470,,,I14808,);
endmodule


