module test_I3846(I1750,I1668,I1477,I2072,I1470,I1603,I3846);
input I1750,I1668,I1477,I2072,I1470,I1603;
output I3846;
wire I1518,I3388,I1504,I1880,I3555,I3538,I1510,I3747,I1492,I1897,I1767;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
nand I_2(I1504,I1767,I1897);
nor I_3(I3846,I3747,I3555);
DFFARX1 I_4(I1470,I1518,,,I1880,);
DFFARX1 I_5(I3538,I1470,I3388,,,I3555,);
nor I_6(I3538,I1492,I1510);
DFFARX1 I_7(I2072,I1470,I1518,,,I1510,);
DFFARX1 I_8(I1504,I1470,I3388,,,I3747,);
nand I_9(I1492,I1603,I1668);
nor I_10(I1897,I1880,I1603);
DFFARX1 I_11(I1750,I1470,I1518,,,I1767,);
endmodule


