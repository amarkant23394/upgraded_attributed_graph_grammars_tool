module test_I9655(I5716,I1477,I6127,I6079,I1470,I5898,I9655);
input I5716,I1477,I6127,I6079,I1470,I5898;
output I9655;
wire I5737,I8267,I8216,I8360,I6203,I8623,I5743,I8196,I5719,I8377,I8250,I8190;
nand I_0(I5737,I6203,I5898);
nand I_1(I8267,I8250,I5737);
not I_2(I8216,I1477);
not I_3(I8360,I5719);
DFFARX1 I_4(I1470,,,I6203,);
DFFARX1 I_5(I5743,I1470,I8216,,,I8623,);
nand I_6(I5743,I6127,I6079);
nand I_7(I8196,I8623,I8377);
nand I_8(I9655,I8190,I8196);
DFFARX1 I_9(I1470,,,I5719,);
not I_10(I8377,I8360);
nor I_11(I8250,I5719,I5716);
DFFARX1 I_12(I8267,I1470,I8216,,,I8190,);
endmodule


