module test_final(G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7,n_431_0_l_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_7,blif_clk_net_1_r_0,n6_0,G42_1_r_7,);
nor I_1(n_572_1_r_7,n30_7,n31_7);
nand I_2(n_573_1_r_7,IN_7_0_l_7,n28_7);
nor I_3(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_4(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_5(N1_4_r_7,blif_clk_net_1_r_0,n6_0,G199_4_r_7,);
DFFARX1 I_6(n26_7,blif_clk_net_1_r_0,n6_0,G214_4_r_7,);
DFFARX1 I_7(n5_7,blif_clk_net_1_r_0,n6_0,ACVQN1_5_r_7,);
not I_8(P6_5_r_7,P6_5_r_internal_7);
or I_9(n_431_0_l_7,IN_8_0_l_7,n36_7);
DFFARX1 I_10(n_431_0_l_7,blif_clk_net_1_r_0,n6_0,n43_7,);
not I_11(n27_7,n43_7);
DFFARX1 I_12(IN_2_5_l_7,blif_clk_net_1_r_0,n6_0,ACVQN1_5_l_7,);
DFFARX1 I_13(IN_1_5_l_7,blif_clk_net_1_r_0,n6_0,n44_7,);
nor I_14(n4_1_r_7,n30_7,n38_7);
nor I_15(N1_4_r_7,n27_7,n40_7);
nand I_16(n26_7,IN_11_0_l_7,n39_7);
not I_17(n5_7,G2_0_l_7);
DFFARX1 I_18(ACVQN1_5_l_7,blif_clk_net_1_r_0,n6_0,P6_5_r_internal_7,);
nor I_19(n28_7,n26_7,n29_7);
not I_20(n29_7,IN_5_0_l_7);
not I_21(n30_7,G1_0_l_7);
nand I_22(n31_7,n27_7,n29_7);
nor I_23(n32_7,ACVQN1_5_l_7,n34_7);
nor I_24(n33_7,G2_0_l_7,n29_7);
not I_25(n34_7,IN_7_0_l_7);
nor I_26(n35_7,n43_7,n44_7);
and I_27(n36_7,IN_2_0_l_7,n37_7);
nor I_28(n37_7,IN_4_0_l_7,n30_7);
nand I_29(n38_7,G2_0_l_7,n29_7);
nor I_30(n39_7,G2_0_l_7,IN_10_0_l_7);
nor I_31(n40_7,n44_7,n41_7);
nor I_32(n41_7,n34_7,n42_7);
nand I_33(n42_7,IN_5_0_l_7,n5_7);
DFFARX1 I_34(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_35(n_572_1_r_0,n23_0,G199_4_r_7);
nand I_36(n_573_1_r_0,n21_0,n22_0);
nand I_37(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_38(n_569_1_r_0,n21_0,n26_0);
nor I_39(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_40(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_41(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_42(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_43(n4_1_l_0,n_549_1_r_7,n_572_1_r_7);
not I_44(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_45(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_46(G214_4_r_7,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_47(n20_0,n38_0);
DFFARX1 I_48(G42_1_r_7,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_49(n4_1_r_0,n23_0,G42_1_r_7);
nor I_50(N3_2_r_0,n31_0,n32_0);
nor I_51(N1_4_r_0,n29_0,n32_0);
not I_52(n2_0,n31_0);
nor I_53(n21_0,n37_0,n_569_1_r_7);
not I_54(n22_0,G199_4_r_7);
nand I_55(n23_0,n20_0,n30_0);
nand I_56(n24_0,n38_0,n25_0);
nor I_57(n25_0,G42_1_r_7,n_569_1_r_7);
not I_58(n26_0,G42_1_r_7);
not I_59(n27_0,n29_0);
nor I_60(n28_0,n_572_1_r_7,P6_5_r_7);
nand I_61(n29_0,n26_0,n33_0);
not I_62(n30_0,n_569_1_r_7);
nand I_63(n31_0,ACVQN1_3_l_0,ACVQN1_5_r_7);
and I_64(n32_0,n35_0,n36_0);
nand I_65(n33_0,n34_0,n_573_1_r_7);
not I_66(n34_0,n_572_1_r_7);
nor I_67(n35_0,n_572_1_r_7,n_573_1_r_7);
nor I_68(n36_0,G199_4_r_7,P6_5_r_7);
endmodule


