module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_5_r_15,n9_15,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_5_r_15,n9_15,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
and I_40(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_41(N1508_0_r_15,n55_15,N1508_1_r_16);
nor I_42(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_43(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_44(N1372_4_r_15,n39_15);
nor I_45(N1508_4_r_15,n39_15,n43_15);
nand I_46(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_47(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_48(n_576_5_r_15,n31_15,n32_15);
not I_49(n_102_5_r_15,n33_15);
nand I_50(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_51(N1507_6_r_15,n42_15,n46_15);
nand I_52(N1508_6_r_15,n39_15,n40_15);
nand I_53(n_431_5_r_15,n36_15,n37_15);
not I_54(n9_15,blif_reset_net_5_r_15);
nor I_55(n31_15,n33_15,n34_15);
nor I_56(n32_15,n44_15,G42_7_r_16);
nor I_57(n33_15,n54_15,n55_15);
nand I_58(n34_15,n49_15,N6147_2_r_16);
nand I_59(n35_15,n_573_7_r_16,n_569_7_r_16);
not I_60(n36_15,n32_15);
nand I_61(n37_15,n34_15,n38_15);
not I_62(n38_15,n46_15);
nand I_63(n39_15,n38_15,n41_15);
nand I_64(n40_15,n41_15,n42_15);
and I_65(n41_15,n51_15,N1372_1_r_16);
and I_66(n42_15,n47_15,n_569_7_r_16);
and I_67(n43_15,n34_15,n36_15);
or I_68(n44_15,n_572_7_r_16,N1372_1_r_16);
not I_69(n45_15,N1372_1_r_15);
nand I_70(n46_15,n53_15,n_569_7_r_16);
nor I_71(n47_15,n34_15,n48_15);
not I_72(n48_15,n_573_7_r_16);
and I_73(n49_15,n50_15,N1507_6_r_16);
nand I_74(n50_15,n51_15,n52_15);
nand I_75(n51_15,N1371_0_r_16,N1508_0_r_16);
not I_76(n52_15,N1372_1_r_16);
nor I_77(n53_15,n48_15,N1508_6_r_16);
nor I_78(n54_15,n_452_7_r_16,N1371_0_r_16);
not I_79(n55_15,N1508_0_r_16);
endmodule


